//Written by the Majority Logic Package Thu Apr 30 13:06:44 2015
module top (
            pi00, pi01, pi02, pi03, pi04, pi05, pi06, pi07, pi08, pi09, pi10, pi11, pi12, pi13, pi14, pi15, pi16, pi17, pi18, pi19, pi20, pi21, pi22, pi23, pi24, pi25, pi26, pi27, pi28, pi29, pi30, pi31, pi32, pi33, pi34, pi35, pi36, pi37, pi38, pi39, pi40, pi41, pi42, pi43, pi44, pi45, pi46, pi47, pi48, pi49, pi50, pi51, pi52, pi53, pi54, pi55, pi56, pi57, pi58, pi59, pi60, pi61, pi62, pi63, pi64, pi65, pi66, pi67, pi68, pi69, pi70, pi71, pi72, pi73, pi74, pi75, pi76, pi77, pi78, pi79, pi80, pi81, pi82, pi83, pi84, 
            po00, po01, po02, po03, po04, po05, po06, po07, po08, po09, po10, po11, po12, po13, po14, po15, po16, po17, po18, po19, po20, po21, po22, po23, po24, po25, po26, po27, po28, po29, po30, po31, po32, po33, po34, po35, po36, po37, po38, po39, po40, po41, po42, po43, po44, po45, po46, po47, po48, po49, po50, po51, po52, po53, po54, po55, po56, po57, po58, po59, po60, po61, po62, po63, po64, po65, po66, po67, po68, po69, po70, po71, po72, po73, po74, po75);
input pi00, pi01, pi02, pi03, pi04, pi05, pi06, pi07, pi08, pi09, pi10, pi11, pi12, pi13, pi14, pi15, pi16, pi17, pi18, pi19, pi20, pi21, pi22, pi23, pi24, pi25, pi26, pi27, pi28, pi29, pi30, pi31, pi32, pi33, pi34, pi35, pi36, pi37, pi38, pi39, pi40, pi41, pi42, pi43, pi44, pi45, pi46, pi47, pi48, pi49, pi50, pi51, pi52, pi53, pi54, pi55, pi56, pi57, pi58, pi59, pi60, pi61, pi62, pi63, pi64, pi65, pi66, pi67, pi68, pi69, pi70, pi71, pi72, pi73, pi74, pi75, pi76, pi77, pi78, pi79, pi80, pi81, pi82, pi83, pi84;
output po00, po01, po02, po03, po04, po05, po06, po07, po08, po09, po10, po11, po12, po13, po14, po15, po16, po17, po18, po19, po20, po21, po22, po23, po24, po25, po26, po27, po28, po29, po30, po31, po32, po33, po34, po35, po36, po37, po38, po39, po40, po41, po42, po43, po44, po45, po46, po47, po48, po49, po50, po51, po52, po53, po54, po55, po56, po57, po58, po59, po60, po61, po62, po63, po64, po65, po66, po67, po68, po69, po70, po71, po72, po73, po74, po75;
wire one, v0, v1, v2, v3, v4, v5, v6, v7, v8, v9, v10, v11, v12, v13, v14, v15, v16, v17, v18, v19, v20, v21, v22, v23, v24, v25, v26, v27, v28, v29, v30, v31, v32, v33, v34, v35, v36, v37, v38, v39, v40, v41, v42, v43, v44, v45, v46, v47, v48, v49, v50, v51, v52, v53, v54, v55, v56, v57, v58, v59, v60, v61, v62, v63, v64, v65, v66, v67, v68, v69, v70, v71, v72, v73, v74, v75, v76, v77, v78, v79, v80, v81, v82, v83, v84, v85, v86, v87, v88, v89, v90, v91, v92, v93, v94, v95, v96, v97, v98, v99, v100, v101, v102, v103, v104, v105, v106, v107, v108, v109, v110, v111, v112, v113, v114, v115, v116, v117, v118, v119, v120, v121, v122, v123, v124, v125, v126, v127, v128, v129, v130, v131, v132, v133, v134, v135, v136, v137, v138, v139, v140, v141, v142, v143, v144, v145, v146, v147, v148, v149, v150, v151, v152, v153, v154, 
 w0, w1, w2, w3, w4, w5, w6, w7, w8, w9, w10, w11, w12, w13, w14, w15, w16, w17, w18, w19, w20, w21, w22, w23, w24, w25, w26, w27, w28, w29, w30, w31, w32, w33, w34, w35, w36, w37, w38, w39, w40, w41, w42, w43, w44, w45, w46, w47, w48, w49, w50, w51, w52, w53, w54, w55, w56, w57, w58, w59, w60, w61, w62, w63, w64, w65, w66, w67, w68, w69, w70, w71, w72, w73, w74, w75, w76, w77, w78, w79, w80, w81, w82, w83, w84, w85, w86, w87, w88, w89, w90, w91, w92, w93, w94, w95, w96, w97, w98, w99, w100, w101, w102, w103, w104, w105, w106, w107, w108, w109, w110, w111, w112, w113, w114, w115, w116, w117, w118, w119, w120, w121, w122, w123, w124, w125, w126, w127, w128, w129, w130, w131, w132, w133, w134, w135, w136, w137, w138, w139, w140, w141, w142, w143, w144, w145, w146, w147, w148, w149, w150, w151, w152, w153, w154, w155, w156, w157, w158, w159, w160, w161, w162, w163, w164, w165, w166, w167, w168, w169, w170, w171, w172, w173, w174, w175, w176, w177, w178, w179, w180, w181, w182, w183, w184, w185, w186, w187, w188, w189, w190, w191, w192, w193, w194, w195, w196, w197, w198, w199, w200, w201, w202, w203, w204, w205, w206, w207, w208, w209, w210, w211, w212, w213, w214, w215, w216, w217, w218, w219, w220, w221, w222, w223, w224, w225, w226, w227, w228, w229, w230, w231, w232, w233, w234, w235, w236, w237, w238, w239, w240, w241, w242, w243, w244, w245, w246, w247, w248, w249, w250, w251, w252, w253, w254, w255, w256, w257, w258, w259, w260, w261, w262, w263, w264, w265, w266, w267, w268, w269, w270, w271, w272, w273, w274, w275, w276, w277, w278, w279, w280, w281, w282, w283, w284, w285, w286, w287, w288, w289, w290, w291, w292, w293, w294, w295, w296, w297, w298, w299, w300, w301, w302, w303, w304, w305, w306, w307, w308, w309, w310, w311, w312, w313, w314, w315, w316, w317, w318, w319, w320, w321, w322, w323, w324, w325, w326, w327, w328, w329, w330, w331, w332, w333, w334, w335, w336, w337, w338, w339, w340, w341, w342, w343, w344, w345, w346, w347, w348, w349, w350, w351, w352, w353, w354, w355, w356, w357, w358, w359, w360, w361, w362, w363, w364, w365, w366, w367, w368, w369, w370, w371, w372, w373, w374, w375, w376, w377, w378, w379, w380, w381, w382, w383, w384, w385, w386, w387, w388, w389, w390, w391, w392, w393, w394, w395, w396, w397, w398, w399, w400, w401, w402, w403, w404, w405, w406, w407, w408, w409, w410, w411, w412, w413, w414, w415, w416, w417, w418, w419, w420, w421, w422, w423, w424, w425, w426, w427, w428, w429, w430, w431, w432, w433, w434, w435, w436, w437, w438, w439, w440, w441, w442, w443, w444, w445, w446, w447, w448, w449, w450, w451, w452, w453, w454, w455, w456, w457, w458, w459, w460, w461, w462, w463, w464, w465, w466, w467, w468, w469, w470, w471, w472, w473, w474, w475, w476, w477, w478, w479, w480, w481, w482, w483, w484, w485, w486, w487, w488, w489, w490, w491, w492, w493, w494, w495, w496, w497, w498, w499, w500, w501, w502, w503, w504, w505, w506, w507, w508, w509, w510, w511, w512, w513, w514, w515, w516, w517, w518, w519, w520, w521, w522, w523, w524, w525, w526, w527, w528, w529, w530, w531, w532, w533, w534, w535, w536, w537, w538, w539, w540, w541, w542, w543, w544, w545, w546, w547, w548, w549, w550, w551, w552, w553, w554, w555, w556, w557, w558, w559, w560, w561, w562, w563, w564, w565, w566, w567, w568, w569, w570, w571, w572, w573, w574, w575, w576, w577, w578, w579, w580, w581, w582, w583, w584, w585, w586, w587, w588, w589, w590, w591, w592, w593, w594, w595, w596, w597, w598, w599, w600, w601, w602, w603, w604, w605, w606, w607, w608, w609, w610, w611, w612, w613, w614, w615, w616, w617, w618, w619, w620, w621, w622, w623, w624, w625, w626, w627, w628, w629, w630, w631, w632, w633, w634, w635, w636, w637, w638, w639, w640, w641, w642, w643, w644, w645, w646, w647, w648, w649, w650, w651, w652, w653, w654, w655, w656, w657, w658, w659, w660, w661, w662, w663, w664, w665, w666, w667, w668, w669, w670, w671, w672, w673, w674, w675, w676, w677, w678, w679, w680, w681, w682, w683, w684, w685, w686, w687, w688, w689, w690, w691, w692, w693, w694, w695, w696, w697, w698, w699, w700, w701, w702, w703, w704, w705, w706, w707, w708, w709, w710, w711, w712, w713, w714, w715, w716, w717, w718, w719, w720, w721, w722, w723, w724, w725, w726, w727, w728, w729, w730, w731, w732, w733, w734, w735, w736, w737, w738, w739, w740, w741, w742, w743, w744, w745, w746, w747, w748, w749, w750, w751, w752, w753, w754, w755, w756, w757, w758, w759, w760, w761, w762, w763, w764, w765, w766, w767, w768, w769, w770, w771, w772, w773, w774, w775, w776, w777, w778, w779, w780, w781, w782, w783, w784, w785, w786, w787, w788, w789, w790, w791, w792, w793, w794, w795, w796, w797, w798, w799, w800, w801, w802, w803, w804, w805, w806, w807, w808, w809, w810, w811, w812, w813, w814, w815, w816, w817, w818, w819, w820, w821, w822, w823, w824, w825, w826, w827, w828, w829, w830, w831, w832, w833, w834, w835, w836, w837, w838, w839, w840, w841, w842, w843, w844, w845, w846, w847, w848, w849, w850, w851, w852, w853, w854, w855, w856, w857, w858, w859, w860, w861, w862, w863, w864, w865, w866, w867, w868, w869, w870, w871, w872, w873, w874, w875, w876, w877, w878, w879, w880, w881, w882, w883, w884, w885, w886, w887, w888, w889, w890, w891, w892, w893, w894, w895, w896, w897, w898, w899, w900, w901, w902, w903, w904, w905, w906, w907, w908, w909, w910, w911, w912, w913, w914, w915, w916, w917, w918, w919, w920, w921, w922, w923, w924, w925, w926, w927, w928, w929, w930, w931;
assign w0 = ~w793 & w226;
assign w1 = (w747 & ~w116) | (w747 & w240) | (~w116 & w240);
assign w2 = w492 & w600;
assign w3 = w529 & w295;
assign w4 = w134 & pi14;
assign w5 = w218 & w515;
assign w6 = (w422 & w43) | (w422 & w85) | (w43 & w85);
assign w7 = pi03 & ~w324;
assign v0 = ~(w750 | w6);
assign w8 = v0;
assign w9 = w141 & w434;
assign w10 = w587 & w731;
assign w11 = w492 & w707;
assign w12 = (~pi46 & ~w877) | (~pi46 & w888) | (~w877 & w888);
assign v1 = ~(w858 | w120);
assign w13 = v1;
assign w14 = (pi15 & ~w823) | (pi15 & w77) | (~w823 & w77);
assign w15 = pi28 & pi11;
assign w16 = w764 & w243;
assign v2 = ~(pi50 | w518);
assign w17 = v2;
assign w18 = (pi11 & w419) | (pi11 & w674) | (w419 & w674);
assign v3 = ~(pi02 | w684);
assign w19 = v3;
assign w20 = ~w764 & pi57;
assign w21 = ~w588 & w918;
assign w22 = (w337 & w229) | (w337 & w437) | (w229 & w437);
assign w23 = ~w805 & w386;
assign w24 = w134 & w826;
assign v4 = ~(w513 | w64);
assign w25 = v4;
assign w26 = w70 & w851;
assign w27 = w134 & pi12;
assign w28 = pi39 & w315;
assign w29 = ~pi84 & w130;
assign w30 = ~pi28 & w403;
assign w31 = w629 & w527;
assign w32 = w96 & w421;
assign v5 = ~(w295 | pi08);
assign w33 = v5;
assign w34 = w408 & ~pi10;
assign w35 = w64 & w445;
assign w36 = w614 & w817;
assign w37 = (pi52 & ~w492) | (pi52 & w638) | (~w492 & w638);
assign w38 = w643 & w919;
assign w39 = (pi44 & w273) | (pi44 & w755) | (w273 & w755);
assign w40 = w764 & pi51;
assign w41 = (pi19 & ~w703) | (pi19 & w760) | (~w703 & w760);
assign w42 = w30 & w651;
assign w43 = pi28 & pi27;
assign w44 = w311 & w26;
assign w45 = ~pi29 & w414;
assign w46 = w114 & w195;
assign w47 = ~w359 & w514;
assign w48 = (w594 & w822) | (w594 & w802) | (w822 & w802);
assign w49 = w538 & w381;
assign w50 = pi44 & ~w546;
assign w51 = ~w108 & w92;
assign w52 = pi49 & ~pi63;
assign w53 = w70 & w309;
assign w54 = w218 & w232;
assign w55 = ~w271 & w824;
assign w56 = ~w616 & w564;
assign w57 = ~w585 & w157;
assign w58 = ~w239 & w244;
assign w59 = w805 & w386;
assign w60 = ~w771 & w525;
assign v6 = ~(w320 | w859);
assign w61 = v6;
assign w62 = ~pi06 & pi12;
assign v7 = ~(pi10 | w52);
assign w63 = v7;
assign w64 = w84 & w612;
assign w65 = ~w908 & w299;
assign w66 = (~w311 & w395) | (~w311 & w242) | (w395 & w242);
assign w67 = w826 & ~w401;
assign w68 = w210 & w133;
assign w69 = ~w156 & w46;
assign w70 = w154 & w484;
assign w71 = ~pi28 & pi06;
assign w72 = pi27 & ~pi71;
assign v8 = ~(w454 | w916);
assign w73 = v8;
assign w74 = (w218 & w555) | (w218 & w429) | (w555 & w429);
assign w75 = ~w764 & pi48;
assign w76 = w453 & w366;
assign w77 = (pi15 & ~w538) | (pi15 & w427) | (~w538 & w427);
assign w78 = w573 & ~w658;
assign v9 = ~(pi28 | w209);
assign w79 = v9;
assign w80 = w408 & pi10;
assign w81 = (~w659 & ~w48) | (~w659 & w367) | (~w48 & w367);
assign w82 = (w283 & w571) | (w283 & w796) | (w571 & w796);
assign w83 = ~w41 & w107;
assign w84 = w624 & w670;
assign w85 = (pi28 & w783) | (pi28 & w43) | (w783 & w43);
assign w86 = w483 & w3;
assign w87 = (pi37 & w779) | (pi37 & w179) | (w779 & w179);
assign w88 = (w346 & w156) | (w346 & w302) | (w156 & w302);
assign v10 = ~(w651 | w157);
assign w89 = v10;
assign v11 = ~(pi03 | w218);
assign w90 = v11;
assign v12 = ~(w651 | w3);
assign w91 = v12;
assign w92 = (~w124 & w73) | (~w124 & w193) | (w73 & w193);
assign w93 = ~w295 & pi47;
assign w94 = w804 & w679;
assign w95 = ~w915 & w555;
assign w96 = w665 & w593;
assign w97 = w55 & ~w630;
assign w98 = (w794 & w613) | (w794 & w931) | (w613 & w931);
assign w99 = w25 & w106;
assign w100 = w64 & ~w445;
assign w101 = (pi42 & w100) | (pi42 & w223) | (w100 & w223);
assign w102 = ~pi18 & pi22;
assign w103 = (w218 & w695) | (w218 & w745) | (w695 & w745);
assign v13 = ~(w202 | w262);
assign w104 = v13;
assign w105 = pi38 & ~w887;
assign v14 = ~(w314 | w319);
assign w106 = v14;
assign w107 = (w906 & ~w419) | (w906 & w920) | (~w419 & w920);
assign w108 = w651 & ~w440;
assign w109 = w668 & w540;
assign w110 = w492 & w692;
assign w111 = (pi09 & ~w422) | (pi09 & w850) | (~w422 & w850);
assign w112 = pi03 & w810;
assign w113 = ~w209 & pi07;
assign w114 = w689 & w844;
assign w115 = w731 & w285;
assign v15 = ~(w467 | w882);
assign w116 = v15;
assign w117 = ~pi07 & w311;
assign w118 = ~w733 & w362;
assign w119 = pi34 & ~w97;
assign w120 = (~w790 & ~w311) | (~w790 & w503) | (~w311 & w503);
assign w121 = w783 & pi10;
assign w122 = w756 & ~w666;
assign w123 = w764 & ~w740;
assign w124 = (pi03 & w536) | (pi03 & w625) | (w536 & w625);
assign w125 = (~w772 & ~w798) | (~w772 & w523) | (~w798 & w523);
assign w126 = (~w337 & w247) | (~w337 & w261) | (w247 & w261);
assign w127 = w334 & w533;
assign v16 = ~(pi15 | pi36);
assign w128 = v16;
assign w129 = (~w910 & ~w327) | (~w910 & w580) | (~w327 & w580);
assign w130 = w146 & w500;
assign v17 = ~(w434 | w604);
assign w131 = v17;
assign v18 = ~(w443 | w206);
assign w132 = v18;
assign w133 = (pi10 & ~w783) | (pi10 & w768) | (~w783 & w768);
assign w134 = ~pi19 & pi26;
assign w135 = ~w624 & pi42;
assign w136 = ~w383 & w703;
assign v19 = ~(w168 | w626);
assign w137 = v19;
assign v20 = ~(pi12 | w219);
assign w138 = v20;
assign w139 = (pi30 & ~w148) | (pi30 & w185) | (~w148 & w185);
assign w140 = ~w98 & w270;
assign v21 = ~(pi62 | pi64);
assign w141 = v21;
assign w142 = w384 & w586;
assign w143 = (pi26 & ~w136) | (pi26 & w377) | (~w136 & w377);
assign w144 = w492 & w40;
assign v22 = ~(w256 | w304);
assign w145 = v22;
assign w146 = w689 & w595;
assign w147 = w725 & w643;
assign v23 = ~(w918 | w156);
assign w148 = v23;
assign v24 = ~(w522 | w490);
assign w149 = v24;
assign v25 = ~(w668 | pi50);
assign w150 = v25;
assign w151 = ~w116 & w458;
assign w152 = (~pi18 & ~w844) | (~pi18 & w387) | (~w844 & w387);
assign w153 = (pi51 & ~w492) | (pi51 & w781) | (~w492 & w781);
assign v26 = ~(pi19 | pi26);
assign w154 = v26;
assign w155 = (w218 & w609) | (w218 & w394) | (w609 & w394);
assign w156 = w370 & w662;
assign w157 = w665 & w408;
assign w158 = w66 & w422;
assign w159 = ~w157 & w536;
assign w160 = w706 & pi27;
assign w161 = pi79 & w130;
assign w162 = pi28 & ~pi44;
assign v27 = ~(pi27 | pi08);
assign w163 = v27;
assign w164 = ~pi16 & pi17;
assign w165 = (~w3 & ~w439) | (~w3 & w917) | (~w439 & w917);
assign w166 = w3 & ~w483;
assign w167 = w731 & w258;
assign w168 = (pi31 & ~w529) | (pi31 & w169) | (~w529 & w169);
assign w169 = ~w295 & pi31;
assign v28 = ~(pi13 | pi14);
assign w170 = v28;
assign w171 = pi01 & ~w324;
assign v29 = ~(w337 | w248);
assign w172 = v29;
assign w173 = w794 & ~w132;
assign w174 = ~pi10 & pi00;
assign w175 = (w156 & w837) | (w156 & w87) | (w837 & w87);
assign w176 = w218 & w355;
assign w177 = (pi47 & ~w529) | (pi47 & w93) | (~w529 & w93);
assign w178 = ~w764 & pi56;
assign w179 = w588 & pi37;
assign w180 = (w243 & w827) | (w243 & w397) | (w827 & w397);
assign w181 = ~w187 & w297;
assign w182 = pi33 & pi39;
assign w183 = w732 & ~w479;
assign w184 = ~w143 & w231;
assign w185 = ~w344 & pi30;
assign v30 = ~(w810 | w162);
assign w186 = v30;
assign w187 = (~w209 & w254) | (~w209 & w801) | (w254 & w801);
assign w188 = ~w59 & w251;
assign w189 = pi42 & w100;
assign w190 = w156 & w868;
assign w191 = ~w896 & w610;
assign v31 = ~(pi36 | pi42);
assign w192 = v31;
assign w193 = (~w536 & w557) | (~w536 & w834) | (w557 & w834);
assign w194 = w826 & w150;
assign v32 = ~(w878 | w716);
assign w195 = v32;
assign w196 = ~w826 & w643;
assign w197 = ~w637 & w341;
assign w198 = w723 & w823;
assign w199 = ~w295 & pi45;
assign w200 = (w458 & w489) | (w458 & w151) | (w489 & w151);
assign w201 = w632 & w921;
assign w202 = ~w198 & w76;
assign w203 = (w458 & w65) | (w458 & w36) | (w65 & w36);
assign w204 = w665 & w846;
assign w205 = pi34 & ~pi40;
assign w206 = ~w807 & w338;
assign w207 = w408 & pi13;
assign w208 = (~pi22 & ~w844) | (~pi22 & w257) | (~w844 & w257);
assign v33 = ~(w651 | w204);
assign w209 = v33;
assign w210 = w157 & w783;
assign w211 = w573 & w407;
assign w212 = (w556 & ~w156) | (w556 & w701) | (~w156 & w701);
assign w213 = (pi05 & ~w639) | (pi05 & w886) | (~w639 & w886);
assign v34 = ~(w501 | w345);
assign w214 = v34;
assign v35 = ~(w415 | w139);
assign w215 = v35;
assign w216 = pi00 & ~w368;
assign v36 = ~(w678 | w7);
assign w217 = v36;
assign w218 = w146 & w167;
assign w219 = pi03 & pi28;
assign w220 = w509 & ~w198;
assign w221 = w492 & w867;
assign w222 = ~pi15 & w728;
assign w223 = (pi42 & ~w384) | (pi42 & w135) | (~w384 & w135);
assign w224 = ~pi34 & pi40;
assign w225 = (w283 & w317) | (w283 & w447) | (w317 & w447);
assign w226 = ~w559 & w281;
assign w227 = w764 & pi52;
assign w228 = ~w303 & w818;
assign w229 = w665 & w922;
assign w230 = ~w280 & w60;
assign v37 = ~(w771 | w648);
assign w231 = v37;
assign w232 = w643 & w160;
assign w233 = pi24 & ~w156;
assign w234 = w311 & w444;
assign w235 = w214 & w889;
assign w236 = ~w90 & w201;
assign w237 = ~w783 & pi10;
assign w238 = ~pi44 & w545;
assign w239 = (~pi22 & w156) | (~pi22 & w208) | (w156 & w208);
assign w240 = pi12 & w747;
assign w241 = ~w100 & w918;
assign w242 = (pi39 & w791) | (pi39 & w819) | (w791 & w819);
assign w243 = ~pi34 & w182;
assign w244 = w281 & ~w382;
assign w245 = w170 & pi00;
assign w246 = (~pi02 & ~w70) | (~pi02 & w308) | (~w70 & w308);
assign w247 = w154 & w426;
assign w248 = w76 & w445;
assign w249 = pi27 & ~pi66;
assign w250 = w170 & ~w62;
assign v38 = ~(w292 | w198);
assign w251 = v38;
assign w252 = ~w386 & w25;
assign v39 = ~(pi76 | pi06);
assign w253 = v39;
assign v40 = ~(w385 | w491);
assign w254 = v40;
assign w255 = w157 & w532;
assign w256 = (w805 & ~w662) | (w805 & w487) | (~w662 & w487);
assign v41 = ~(w607 | pi22);
assign w257 = v41;
assign w258 = w587 & ~w832;
assign w259 = w281 & ~w870;
assign w260 = (pi53 & ~w492) | (pi53 & w316) | (~w492 & w316);
assign w261 = w529 & w433;
assign w262 = pi49 & w35;
assign w263 = w529 & w373;
assign w264 = w665 & w4;
assign w265 = ~w673 & w693;
assign w266 = ~pi50 & w668;
assign v42 = ~(w59 | w292);
assign w267 = v42;
assign w268 = pi78 & w130;
assign w269 = w632 & ~w776;
assign w270 = (w82 & w901) | (w82 & w225) | (w901 & w225);
assign w271 = ~w477 & w389;
assign w272 = pi02 & w923;
assign w273 = (~w198 & ~w759) | (~w198 & w202) | (~w759 & w202);
assign v43 = ~(w416 | w474);
assign w274 = v43;
assign w275 = w198 & w767;
assign w276 = w614 & w710;
assign w277 = w311 & w726;
assign w278 = pi12 & ~pi10;
assign w279 = ~w156 & w844;
assign w280 = (pi28 & ~w422) | (pi28 & w792) | (~w422 & w792);
assign w281 = (w267 & w370) | (w267 & w188) | (w370 & w188);
assign w282 = ~w766 & w516;
assign v44 = ~(w363 | w234);
assign w283 = v44;
assign w284 = (~w513 & w106) | (~w513 & w831) | (w106 & w831);
assign w285 = w587 & ~w266;
assign v45 = ~(w315 | w419);
assign w286 = v45;
assign w287 = w458 & w924;
assign w288 = w765 & w671;
assign v46 = ~(w472 | w45);
assign w289 = v46;
assign w290 = w492 & w737;
assign w291 = (pi13 & ~w839) | (pi13 & w907) | (~w839 & w907);
assign w292 = w384 & w709;
assign w293 = pi05 & ~w324;
assign w294 = w575 & ~w521;
assign w295 = pi13 & ~pi14;
assign v47 = ~(w782 | w860);
assign w296 = v47;
assign w297 = ~w325 & w589;
assign w298 = (~pi00 & w275) | (~pi00 & w358) | (w275 & w358);
assign w299 = (pi11 & ~w337) | (pi11 & w729) | (~w337 & w729);
assign w300 = w266 & w458;
assign v48 = ~(w100 | w777);
assign w301 = v48;
assign w302 = w918 & w346;
assign w303 = ~w156 & w446;
assign w304 = (w662 & w471) | (w662 & w380) | (w471 & w380);
assign v49 = ~(w449 | w880);
assign w305 = v49;
assign w306 = ~pi20 & pi21;
assign w307 = pi18 & ~pi22;
assign w308 = pi13 & ~pi02;
assign w309 = ~pi13 & w826;
assign w310 = ~w156 & w712;
assign w311 = w732 & w513;
assign w312 = ~pi00 & pi12;
assign w313 = w826 & ~w832;
assign w314 = w765 & w731;
assign w315 = w439 & w89;
assign w316 = ~w764 & pi53;
assign w317 = ~w458 & w796;
assign w318 = (w774 & ~w492) | (w774 & w255) | (~w492 & w255);
assign w319 = w84 & w715;
assign w320 = ~pi12 & w59;
assign w321 = w826 & ~pi77;
assign w322 = pi27 & pi80;
assign w323 = w311 & w856;
assign w324 = w146 & w115;
assign w325 = (w643 & w254) | (w643 & w746) | (w254 & w746);
assign w326 = (pi43 & ~w651) | (pi43 & w734) | (~w651 & w734);
assign v50 = ~(w28 | w431);
assign w327 = v50;
assign w328 = (pi10 & ~w492) | (pi10 & w763) | (~w492 & w763);
assign w329 = ~w425 & w125;
assign v51 = ~(w314 | w64);
assign w330 = v51;
assign w331 = w731 & w365;
assign v52 = ~(w111 | w211);
assign w332 = v52;
assign v53 = ~(w334 | w536);
assign w333 = v53;
assign w334 = w627 & w861;
assign w335 = pi20 & pi16;
assign w336 = w70 & w784;
assign w337 = w509 & w198;
assign w338 = (w218 & w566) | (w218 & w269) | (w566 & w269);
assign v54 = ~(w268 | w293);
assign w339 = v54;
assign v55 = ~(w114 | pi25);
assign w340 = v55;
assign w341 = ~w894 & w165;
assign w342 = (w130 & w264) | (w130 & w356) | (w264 & w356);
assign w343 = w114 & pi23;
assign w344 = w843 & w849;
assign w345 = w810 & w628;
assign w346 = pi15 & ~w292;
assign w347 = w492 & w428;
assign w348 = (~pi16 & ~w848) | (~pi16 & w914) | (~w848 & w914);
assign w349 = pi33 & ~w55;
assign v56 = ~(w76 | w331);
assign w350 = v56;
assign w351 = w337 & w42;
assign w352 = ~w350 & w688;
assign w353 = w845 & w94;
assign w354 = (pi56 & ~w492) | (pi56 & w178) | (~w492 & w178);
assign w355 = pi27 & ~pi69;
assign w356 = (pi14 & w458) | (pi14 & w560) | (w458 & w560);
assign w357 = (w311 & w632) | (w311 & w138) | (w632 & w138);
assign v57 = ~(pi12 | pi00);
assign w358 = v57;
assign w359 = ~w474 & w756;
assign w360 = (pi02 & ~w762) | (pi02 & w478) | (~w762 & w478);
assign w361 = ~w779 & w21;
assign w362 = w281 & ~w310;
assign w363 = ~w311 & w405;
assign v58 = ~(w442 | w277);
assign w364 = v58;
assign w365 = w765 & ~pi28;
assign w366 = w765 & w238;
assign v59 = ~(w809 | w659);
assign w367 = v59;
assign v60 = ~(w275 | w736);
assign w368 = v60;
assign w369 = ~w509 & w759;
assign w370 = w99 & w902;
assign w371 = ~w203 & w872;
assign w372 = ~w548 & w265;
assign w373 = w295 & pi75;
assign w374 = w893 & ~w581;
assign w375 = w157 & ~w334;
assign v61 = ~(w1 | w539);
assign w376 = v61;
assign w377 = w359 & pi26;
assign w378 = w665 & w34;
assign w379 = (~pi07 & ~w311) | (~pi07 & w852) | (~w311 & w852);
assign w380 = pi41 & ~w691;
assign w381 = pi21 & ~pi10;
assign w382 = ~w156 & w114;
assign w383 = w70 & w666;
assign w384 = pi15 & w453;
assign w385 = ~pi05 & w311;
assign w386 = w424 & w462;
assign v62 = ~(pi17 | pi18);
assign w387 = v62;
assign w388 = ~w213 & w413;
assign w389 = ~w826 & w422;
assign v63 = ~(w757 | w452);
assign w390 = v63;
assign v64 = ~(w419 | w359);
assign w391 = v64;
assign w392 = w614 & w53;
assign w393 = (~w439 & ~w337) | (~w439 & w778) | (~w337 & w778);
assign w394 = w794 & ~w876;
assign w395 = (pi39 & w810) | (pi39 & w455) | (w810 & w455);
assign w396 = pi02 & ~w324;
assign w397 = w492 & w16;
assign w398 = w627 & w530;
assign w399 = (w156 & w50) | (w156 & w39) | (w50 & w39);
assign w400 = ~pi32 & pi38;
assign v65 = ~(w775 | w396);
assign w401 = v65;
assign w402 = ~w291 & w511;
assign w403 = pi00 & ~pi27;
assign w404 = (w274 & w342) | (w274 & w468) | (w342 & w468);
assign w405 = pi02 & pi28;
assign w406 = w295 & pi74;
assign w407 = w422 & w606;
assign w408 = pi19 & ~pi26;
assign w409 = pi27 & pi72;
assign w410 = (~w581 & w117) | (~w581 & w374) | (w117 & w374);
assign v66 = ~(w623 | w284);
assign w411 = v66;
assign w412 = (pi39 & w797) | (pi39 & w328) | (w797 & w328);
assign w413 = ~w475 & w329;
assign w414 = ~w864 & w235;
assign w415 = (pi12 & w59) | (pi12 & w718) | (w59 & w718);
assign w416 = w826 & w614;
assign w417 = w334 & pi01;
assign w418 = w469 & ~pi27;
assign w419 = (w157 & ~w337) | (w157 & w57) | (~w337 & w57);
assign w420 = ~w621 & w789;
assign w421 = pi27 & pi08;
assign w422 = (~w334 & ~w439) | (~w334 & w459) | (~w439 & w459);
assign v67 = ~(w153 | w741);
assign w423 = v67;
assign w424 = w769 & w624;
assign w425 = ~w364 & w398;
assign v68 = ~(pi11 | pi13);
assign w426 = v68;
assign w427 = ~pi21 & pi15;
assign w428 = w764 & w738;
assign w429 = (pi27 & w96) | (pi27 & w232) | (w96 & w232);
assign v69 = ~(w643 | w57);
assign w430 = v69;
assign w431 = w492 & w328;
assign v70 = ~(w848 | pi20);
assign w432 = v70;
assign w433 = (~pi13 & ~w403) | (~pi13 & w450) | (~w403 & w450);
assign w434 = w142 & w166;
assign v71 = ~(pi28 | w510);
assign w435 = v71;
assign v72 = ~(w17 | w883);
assign w436 = v72;
assign w437 = w665 & w925;
assign w438 = w170 & pi10;
assign v73 = ~(w458 | w794);
assign w439 = v73;
assign v74 = ~(w454 | w816);
assign w440 = v74;
assign w441 = w218 & w72;
assign w442 = pi05 & ~w311;
assign v75 = ~(w357 | w379);
assign w443 = v75;
assign w444 = pi06 & pi28;
assign w445 = w823 & w49;
assign w446 = w844 & pi17;
assign w447 = ~w458 & w571;
assign w448 = w904 & w641;
assign w449 = pi58 & w330;
assign w450 = pi28 & ~pi13;
assign w451 = w283 & ~w911;
assign w452 = w35 & w464;
assign w453 = w769 & w192;
assign w454 = w311 & w790;
assign w455 = pi39 & pi28;
assign w456 = w492 & w227;
assign w457 = w313 & w643;
assign w458 = w665 & w134;
assign w459 = w651 & ~w334;
assign w460 = ~w334 & pi12;
assign w461 = pi62 & ~pi64;
assign w462 = pi36 & w670;
assign w463 = ~w368 & w298;
assign w464 = pi46 & ~pi49;
assign w465 = pi19 & w656;
assign v76 = ~(w643 | w157);
assign w466 = v76;
assign w467 = w311 & w510;
assign w468 = (w458 & w598) | (w458 & w276) | (w598 & w276);
assign w469 = w538 & w570;
assign w470 = (w794 & w631) | (w794 & w660) | (w631 & w660);
assign w471 = (pi41 & ~w94) | (pi41 & w866) | (~w94 & w866);
assign v77 = ~(w647 | w414);
assign w472 = v77;
assign w473 = w627 & w245;
assign w474 = w337 & w30;
assign w475 = (~w339 & w54) | (~w339 & w74) | (w54 & w74);
assign w476 = pi70 & ~pi12;
assign w477 = pi28 & w311;
assign w478 = pi02 & pi12;
assign v78 = ~(w220 | w605);
assign w479 = v78;
assign w480 = (w156 & w189) | (w156 & w101) | (w189 & w101);
assign w481 = pi44 & w751;
assign v79 = ~(w334 | w393);
assign w482 = v79;
assign w483 = ~pi63 & w141;
assign w484 = ~pi11 & pi14;
assign v80 = ~(w114 | pi23);
assign w485 = v80;
assign v81 = ~(pi28 | w772);
assign w486 = v81;
assign w487 = w76 & w805;
assign v82 = ~(pi27 | pi04);
assign w488 = v82;
assign v83 = ~(pi28 | w296);
assign w489 = v83;
assign w490 = (pi59 & ~w157) | (pi59 & w857) | (~w157 & w857);
assign w491 = (~w510 & ~w311) | (~w510 & w435) | (~w311 & w435);
assign w492 = w146 & w64;
assign w493 = ~w721 & w554;
assign w494 = ~w918 & w156;
assign w495 = w281 & ~w233;
assign w496 = ~w764 & pi54;
assign v84 = ~(pi24 | pi21);
assign w497 = v84;
assign w498 = w493 & w376;
assign w499 = ~w895 & pi36;
assign w500 = w731 & w288;
assign w501 = w319 & w623;
assign w502 = ~w175 & w104;
assign v85 = ~(pi28 | w790);
assign w503 = v85;
assign v86 = ~(w909 | w12);
assign w504 = v86;
assign w505 = ~pi13 & pi04;
assign v87 = ~(pi22 | pi24);
assign w506 = v87;
assign w507 = w295 & pi64;
assign w508 = (w738 & w827) | (w738 & w347) | (w827 & w347);
assign w509 = w865 & w812;
assign w510 = pi01 & pi28;
assign w511 = ~w541 & w743;
assign w512 = ~w156 & w343;
assign w513 = w424 & w892;
assign v88 = ~(w334 | w434);
assign w514 = v88;
assign w515 = w632 & w249;
assign w516 = ~w565 & w517;
assign w517 = (~w909 & ~w78) | (~w909 & w572) | (~w78 & w572);
assign w518 = w529 & w507;
assign w519 = w628 & w186;
assign w520 = w878 & w307;
assign w521 = (pi01 & w417) | (pi01 & w531) | (w417 & w531);
assign w522 = w157 & w121;
assign w523 = (~w772 & w209) | (~w772 & w486) | (w209 & w486);
assign w524 = w172 & w214;
assign v89 = ~(w127 | w598);
assign w525 = v89;
assign w526 = w218 & w730;
assign w527 = w665 & w27;
assign w528 = (~pi12 & w668) | (~pi12 & w761) | (w668 & w761);
assign w529 = ~pi11 & w154;
assign w530 = w170 & pi28;
assign w531 = (w829 & ~w218) | (w829 & w615) | (~w218 & w615);
assign w532 = w780 & ~pi10;
assign w533 = w805 & w319;
assign v90 = ~(w853 | w182);
assign w534 = v90;
assign w535 = pi02 & ~pi28;
assign w536 = w439 & w91;
assign w537 = (~pi12 & ~w73) | (~pi12 & w694) | (~w73 & w694);
assign w538 = ~pi17 & pi20;
assign w539 = ~w176 & w813;
assign v91 = ~(pi50 | pi04);
assign w540 = v91;
assign w541 = (~w666 & w713) | (~w666 & w122) | (w713 & w122);
assign v92 = ~(w349 | w682);
assign w542 = v92;
assign w543 = (pi49 & ~w378) | (pi49 & w926) | (~w378 & w926);
assign w544 = ~pi10 & pi39;
assign w545 = ~pi15 & pi37;
assign w546 = ~w273 & w241;
assign v93 = ~(w129 | w739);
assign w547 = v93;
assign w548 = (~w209 & w13) | (~w209 & w657) | (w13 & w657);
assign v94 = ~(pi10 | w780);
assign w549 = v94;
assign w550 = (pi45 & ~w529) | (pi45 & w199) | (~w529 & w199);
assign w551 = pi46 & w378;
assign w552 = w826 & w668;
assign w553 = pi13 & pi07;
assign w554 = (~w717 & ~w536) | (~w717 & w825) | (~w536 & w825);
assign w555 = pi27 & w96;
assign w556 = w885 & w835;
assign w557 = (~pi03 & ~w665) | (~pi03 & w836) | (~w665 & w836);
assign v95 = ~(w844 | pi17);
assign w558 = v95;
assign w559 = w724 & ~w156;
assign w560 = w665 & w24;
assign w561 = w627 & w438;
assign w562 = w281 & ~w567;
assign w563 = pi10 & pi59;
assign w564 = ~w279 & w281;
assign w565 = (w651 & w748) | (w651 & w392) | (w748 & w392);
assign w566 = w632 & pi07;
assign w567 = (~pi25 & w156) | (~pi25 & w340) | (w156 & w340);
assign w568 = (pi54 & ~w492) | (pi54 & w496) | (~w492 & w496);
assign w569 = (pi07 & ~w70) | (pi07 & w553) | (~w70 & w553);
assign w570 = pi21 & ~pi28;
assign w571 = (~w651 & ~w536) | (~w651 & w246) | (~w536 & w246);
assign w572 = w754 & ~w909;
assign w573 = w826 & ~w614;
assign w574 = (~pi17 & w156) | (~pi17 & w558) | (w156 & w558);
assign w575 = (~w263 & ~w536) | (~w263 & w617) | (~w536 & w617);
assign v96 = ~(w822 | w533);
assign w576 = v96;
assign v97 = ~(w543 | w68);
assign w577 = v97;
assign w578 = (~pi39 & ~w665) | (~pi39 & w644) | (~w665 & w644);
assign w579 = w492 & w123;
assign w580 = w412 & ~w910;
assign w581 = w823 & w418;
assign w582 = (pi57 & ~w492) | (pi57 & w20) | (~w492 & w20);
assign v98 = ~(w699 | w2);
assign w583 = v98;
assign v99 = ~(w260 | w456);
assign w584 = v99;
assign w585 = w780 & w174;
assign w586 = w624 & w266;
assign w587 = ~pi58 & w765;
assign w588 = w513 & ~w623;
assign w589 = ~w95 & w294;
assign v100 = ~(pi46 | pi63);
assign w590 = v100;
assign v101 = ~(w23 | w742);
assign w591 = v101;
assign w592 = pi28 & pi09;
assign w593 = w134 & ~pi28;
assign w594 = ~pi46 & w378;
assign w595 = w878 & w898;
assign w596 = w804 & w520;
assign w597 = w142 & w667;
assign w598 = w130 & w560;
assign v102 = ~(w399 | w519);
assign w599 = v102;
assign w600 = w764 & pi54;
assign w601 = ~pi30 & pi35;
assign w602 = (w555 & w324) | (w555 & w620) | (w324 & w620);
assign w603 = (w527 & w629) | (w527 & w826) | (w629 & w826);
assign w604 = (pi12 & ~w533) | (pi12 & w460) | (~w533 & w460);
assign w605 = w76 & ~w445;
assign w606 = w146 & w314;
assign w607 = pi17 & pi18;
assign w608 = w767 & w732;
assign w609 = w627 & w900;
assign w610 = w281 & ~w830;
assign v103 = ~(w326 | w392);
assign w611 = v103;
assign w612 = ~pi36 & w601;
assign w613 = w794 & w927;
assign w614 = w146 & w10;
assign w615 = w643 & w810;
assign w616 = (~pi16 & w156) | (~pi16 & w348) | (w156 & w348);
assign v104 = ~(pi01 | w263);
assign w617 = v104;
assign v105 = ~(w905 | w216);
assign w618 = v105;
assign w619 = ~w700 & w495;
assign w620 = w96 & w654;
assign w621 = (w794 & w537) | (w794 & w840) | (w537 & w840);
assign w622 = pi30 & ~pi35;
assign w623 = w823 & w469;
assign w624 = w765 & w728;
assign w625 = w334 & pi03;
assign w626 = w614 & w560;
assign w627 = pi11 & w154;
assign w628 = w198 & w513;
assign w629 = w458 & ~w528;
assign w630 = (~w740 & w827) | (~w740 & w579) | (w827 & w579);
assign w631 = ~pi12 & w13;
assign v106 = ~(pi12 | pi28);
assign w632 = v106;
assign v107 = ~(w119 | w180);
assign w633 = v107;
assign w634 = (w458 & ~w130) | (w458 & w881) | (~w130 & w881);
assign w635 = w311 & w903;
assign w636 = (pi04 & w536) | (pi04 & w680) | (w536 & w680);
assign w637 = ~w635 & w690;
assign w638 = ~w764 & pi52;
assign w639 = ~w531 & w333;
assign w640 = w848 & w686;
assign w641 = w524 & ~w463;
assign w642 = ~w803 & pi14;
assign w643 = w627 & w788;
assign v108 = ~(w408 | pi39);
assign w644 = v108;
assign w645 = w764 & pi58;
assign w646 = w643 & w928;
assign v109 = ~(w183 | w410);
assign w647 = v109;
assign w648 = ~w474 & w713;
assign w649 = ~w200 & w498;
assign w650 = (pi36 & w494) | (pi36 & w499) | (w494 & w499);
assign w651 = ~pi13 & w70;
assign w652 = ~w677 & w81;
assign w653 = w588 & pi38;
assign w654 = pi27 & pi07;
assign w655 = ~w441 & w103;
assign w656 = w70 & w433;
assign w657 = w838 & ~w209;
assign v110 = ~(pi00 | w606);
assign w658 = v110;
assign w659 = (pi10 & ~w157) | (pi10 & w237) | (~w157 & w237);
assign w660 = w655 & w794;
assign w661 = w286 & w482;
assign w662 = w369 & w252;
assign w663 = w764 & pi57;
assign w664 = (pi14 & ~w391) | (pi14 & w642) | (~w391 & w642);
assign w665 = ~pi11 & w170;
assign w666 = (~pi13 & ~w337) | (~pi13 & w433) | (~w337 & w433);
assign w667 = w529 & w705;
assign v111 = ~(pi45 | pi47);
assign w668 = v111;
assign w669 = (~pi04 & w109) | (~pi04 & ~w416) | (w109 & ~w416);
assign v112 = ~(pi15 | pi42);
assign w670 = v112;
assign w671 = ~pi58 & pi50;
assign w672 = ~w899 & w131;
assign w673 = ~w681 & w727;
assign w674 = w315 & pi11;
assign w675 = ~w786 & w821;
assign w676 = w614 & w714;
assign w677 = (w614 & w561) | (w614 & w685) | (w561 & w685);
assign w678 = pi83 & w130;
assign w679 = w799 & w506;
assign w680 = w70 & w505;
assign w681 = ~pi82 & w130;
assign w682 = (~pi33 & w827) | (~pi33 & w110) | (w827 & w110);
assign w683 = (~pi08 & ~w529) | (~pi08 & w33) | (~w529 & w33);
assign w684 = w70 & w697;
assign w685 = w794 & ~w912;
assign w686 = w102 & w164;
assign v113 = ~(w704 | w508);
assign w687 = v113;
assign w688 = w823 & w806;
assign w689 = pi22 & w607;
assign w690 = (w311 & w113) | (w311 & w862) | (w113 & w862);
assign w691 = w76 & w353;
assign w692 = w764 & ~pi33;
assign w693 = (~w3 & w422) | (~w3 & w683) | (w422 & w683);
assign w694 = w810 & w875;
assign w695 = w632 & pi08;
assign v114 = ~(w634 | w636);
assign w696 = v114;
assign w697 = ~pi13 & w535;
assign v115 = ~(w354 | w290);
assign w698 = v115;
assign w699 = (pi55 & ~w492) | (pi55 & w811) | (~w492 & w811);
assign w700 = ~pi24 & w156;
assign w701 = w918 & w556;
assign w702 = ~w650 & w591;
assign v116 = ~(w159 | w890);
assign w703 = v116;
assign w704 = pi40 & ~w97;
assign w705 = w295 & w461;
assign w706 = ~pi28 & pi67;
assign w707 = w764 & pi53;
assign w708 = ~w624 & pi35;
assign w709 = w624 & pi12;
assign w710 = w552 & pi14;
assign v117 = ~(w550 | w597);
assign w711 = v117;
assign w712 = w844 & w607;
assign w713 = (w458 & w300) | (w458 & ~w416) | (w300 & ~w416);
assign w714 = w826 & w832;
assign w715 = ~pi36 & w622;
assign w716 = ~pi23 & pi25;
assign w717 = w529 & w720;
assign w718 = w292 & pi12;
assign w719 = pi25 & pi41;
assign w720 = w295 & pi76;
assign w721 = (w651 & w722) | (w651 & w44) | (w722 & w44);
assign w722 = (pi06 & ~w311) | (pi06 & w71) | (~w311 & w71);
assign w723 = pi21 & w538;
assign w724 = pi20 & w848;
assign w725 = w313 & pi68;
assign w726 = pi04 & ~pi12;
assign w727 = (w555 & w324) | (w555 & w32) | (w324 & w32);
assign v118 = ~(pi37 | pi44);
assign w728 = v118;
assign w729 = (pi11 & ~w403) | (pi11 & w15) | (~w403 & w15);
assign w730 = w826 & w476;
assign w731 = w453 & w481;
assign w732 = w845 & w640;
assign w733 = (~pi18 & w156) | (~pi18 & w152) | (w156 & w152);
assign w734 = (pi43 & ~w403) | (pi43 & w874) | (~w403 & w874);
assign w735 = ~w69 & w562;
assign w736 = w445 & w331;
assign w737 = w764 & pi55;
assign w738 = w182 & w205;
assign w739 = (w422 & w323) | (w422 & w158) | (w323 & w158);
assign w740 = pi34 & w182;
assign w741 = w492 & w663;
assign w742 = w736 & w312;
assign v119 = ~(w22 | w351);
assign w743 = v119;
assign v120 = ~(pi20 | pi23);
assign w744 = v120;
assign w745 = w632 & ~w163;
assign w746 = w614 & w147;
assign w747 = w627 & w250;
assign w748 = pi00 & w929;
assign w749 = (pi38 & w273) | (pi38 & w653) | (w273 & w653);
assign w750 = pi27 & ~w407;
assign v121 = ~(pi15 | pi37);
assign w751 = v121;
assign w752 = ~pi28 & pi03;
assign w753 = w198 & ~w100;
assign v122 = ~(w422 | w473);
assign w754 = v122;
assign w755 = w100 & pi44;
assign w756 = (w643 & ~w614) | (w643 & w196) | (~w614 & w196);
assign w757 = (w156 & w105) | (w156 & w749) | (w105 & w749);
assign w758 = pi01 & ~pi28;
assign v123 = ~(w767 | w314);
assign w759 = v123;
assign w760 = (~w337 & w465) | (~w337 & w336) | (w465 & w336);
assign w761 = pi50 & ~pi12;
assign w762 = pi28 & ~pi12;
assign w763 = w534 & pi10;
assign w764 = w665 & w80;
assign v124 = ~(pi32 | pi38);
assign w765 = v124;
assign w766 = pi00 & ~w661;
assign w767 = w865 & w400;
assign w768 = ~pi45 & pi10;
assign v125 = ~(pi30 | pi35);
assign w769 = v125;
assign v126 = ~(w714 | pi19);
assign w770 = v126;
assign w771 = w614 & w457;
assign w772 = w529 & w406;
assign w773 = w863 & w716;
assign w774 = w157 & ~w549;
assign w775 = pi81 & w130;
assign v127 = ~(pi27 | pi07);
assign w776 = v127;
assign w777 = ~w198 & w314;
assign v128 = ~(w30 | w439);
assign w778 = v128;
assign w779 = (~w198 & ~w759) | (~w198 & w220) | (~w759 & w220);
assign v129 = ~(pi46 | pi49);
assign w780 = v129;
assign w781 = ~w764 & pi51;
assign w782 = (pi06 & ~w324) | (pi06 & w820) | (~w324 & w820);
assign w783 = w853 & w224;
assign w784 = ~pi13 & pi19;
assign v130 = ~(w582 | w800);
assign w785 = v130;
assign w786 = ~w5 & w155;
assign w787 = ~w88 & w448;
assign w788 = w170 & ~pi12;
assign w789 = ~w287 & w51;
assign w790 = pi08 & pi28;
assign w791 = w810 & pi39;
assign w792 = ~w783 & pi28;
assign w793 = (~pi20 & w156) | (~pi20 & w432) | (w156 & w432);
assign w794 = w170 & w627;
assign w795 = ~w173 & w197;
assign w796 = (~w684 & ~w536) | (~w684 & w19) | (~w536 & w19);
assign w797 = w780 & w544;
assign w798 = pi04 & w311;
assign v131 = ~(pi18 | pi21);
assign w799 = v131;
assign w800 = w492 & w645;
assign w801 = w758 & ~w209;
assign w802 = w378 & w590;
assign w803 = w839 & ~w126;
assign v132 = ~(pi16 | pi17);
assign w804 = v132;
assign w805 = w724 & w596;
assign w806 = w538 & w891;
assign w807 = w218 & w873;
assign w808 = ~w512 & w259;
assign w809 = pi49 & pi63;
assign v133 = ~(pi27 | pi28);
assign w810 = v133;
assign w811 = ~w764 & pi55;
assign w812 = pi32 & ~pi38;
assign w813 = (w218 & w646) | (w218 & w38) | (w646 & w38);
assign v134 = ~(w177 | w9);
assign w814 = v134;
assign w815 = ~w190 & w855;
assign w816 = (pi03 & ~w311) | (pi03 & w752) | (~w311 & w752);
assign w817 = w194 & w458;
assign w818 = w281 & ~w574;
assign w819 = w534 & pi28;
assign w820 = ~pi27 & pi06;
assign w821 = (~w636 & w669) | (~w636 & w696) | (w669 & w696);
assign w822 = w732 & w76;
assign w823 = w102 & w773;
assign v135 = ~(w315 | w318);
assign w824 = v135;
assign w825 = (~pi06 & w253) | (~pi06 & ~w3) | (w253 & ~w3);
assign w826 = pi27 & ~pi28;
assign w827 = w422 & w477;
assign w828 = (~w209 & ~w311) | (~w209 & w79) | (~w311 & w79);
assign w829 = ~pi28 & w643;
assign w830 = w848 & ~w156;
assign v136 = ~(w198 | w513);
assign w831 = v136;
assign w832 = pi31 & ~pi50;
assign w833 = (~pi19 & ~w614) | (~pi19 & w770) | (~w614 & w770);
assign v137 = ~(w458 | w625);
assign w834 = v137;
assign v138 = ~(w100 | w220);
assign w835 = v138;
assign v139 = ~(w134 | pi03);
assign w836 = v139;
assign w837 = pi37 & ~w361;
assign w838 = pi08 & ~pi28;
assign w839 = (~w334 & ~w536) | (~w334 & w375) | (~w536 & w375);
assign w840 = w236 & w794;
assign v140 = ~(pi28 | pi07);
assign w841 = v140;
assign v141 = ~(w826 | w112);
assign w842 = v141;
assign v142 = ~(w273 | w588);
assign w843 = v142;
assign w844 = w848 & w335;
assign w845 = ~pi25 & w744;
assign w846 = w134 & ~w826;
assign v143 = ~(w480 | w411);
assign w847 = v143;
assign w848 = pi21 & pi24;
assign w849 = (~w100 & w99) | (~w100 & w753) | (w99 & w753);
assign w850 = (pi09 & ~w403) | (pi09 & w592) | (~w403 & w592);
assign w851 = ~pi13 & w510;
assign w852 = pi12 & ~pi07;
assign v144 = ~(pi33 | pi39);
assign w853 = v144;
assign v145 = ~(w568 | w221);
assign w854 = v145;
assign v146 = ~(w100 | w352);
assign w855 = v146;
assign w856 = (pi28 & ~w311) | (pi28 & w819) | (~w311 & w819);
assign w857 = (pi59 & w780) | (pi59 & w563) | (w780 & w563);
assign w858 = ~pi02 & w311;
assign w859 = w780 & w35;
assign w860 = w130 & w322;
assign w861 = w170 & pi12;
assign v147 = ~(w209 | w841);
assign w862 = v147;
assign w863 = pi16 & ~pi24;
assign w864 = w732 & ~w662;
assign w865 = w453 & w222;
assign w866 = (pi41 & ~w744) | (pi41 & w719) | (~w744 & w719);
assign w867 = w764 & pi48;
assign w868 = (pi35 & ~w384) | (pi35 & w708) | (~w384 & w708);
assign v148 = ~(w871 | w11);
assign w869 = v148;
assign w870 = (~pi23 & w156) | (~pi23 & w485) | (w156 & w485);
assign w871 = (pi48 & ~w492) | (pi48 & w75) | (~w492 & w75);
assign w872 = ~w18 & w47;
assign w873 = pi27 & ~pi73;
assign w874 = pi28 & pi43;
assign w875 = pi03 & ~pi12;
assign w876 = (~pi04 & ~w632) | (~pi04 & w488) | (~w632 & w488);
assign w877 = w157 & ~w63;
assign w878 = pi23 & ~pi25;
assign v149 = ~(w664 | w404);
assign w879 = v149;
assign w880 = pi65 & ~w330;
assign w881 = ~w321 & w458;
assign w882 = ~w311 & w444;
assign w883 = w3 & ~w142;
assign v150 = ~(w37 | w144);
assign w884 = v150;
assign v151 = ~(w588 | w202);
assign w885 = v151;
assign w886 = w828 & pi05;
assign w887 = ~w273 & w21;
assign w888 = ~pi46 & w133;
assign w889 = w172 & w576;
assign w890 = (w3 & ~w142) | (w3 & w86) | (~w142 & w86);
assign w891 = pi21 & pi10;
assign w892 = pi42 & w128;
assign w893 = w319 & ~w623;
assign w894 = ~w29 & w602;
assign w895 = w885 & w301;
assign w896 = (~pi21 & w156) | (~pi21 & w497) | (w156 & w497);
assign w897 = ~w470 & w372;
assign w898 = w863 & w306;
assign w899 = (w614 & w31) | (w614 & w603) | (w31 & w603);
assign w900 = w170 & pi04;
assign w901 = ~w67 & w451;
assign w902 = ~w76 & w759;
assign w903 = ~pi03 & pi28;
assign w904 = ~w913 & w61;
assign w905 = pi32 & ~w212;
assign w906 = (w337 & w466) | (w337 & w430) | (w466 & w430);
assign w907 = w890 & pi13;
assign w908 = w826 & w130;
assign w909 = w551 & w608;
assign w910 = (~w157 & ~w315) | (~w157 & w578) | (~w315 & w578);
assign w911 = ~pi27 & w535;
assign w912 = (~pi10 & ~w714) | (~pi10 & w278) | (~w714 & w278);
assign w913 = ~w99 & w14;
assign v152 = ~(pi20 | pi16);
assign w914 = v152;
assign v153 = ~(w161 | w171);
assign w915 = v153;
assign w916 = ~w311 & w219;
assign v154 = ~(w569 | w3);
assign w917 = v154;
assign w918 = w624 & w384;
assign w919 = (w71 & ~pi28) | (w71 & pi27) | (~pi28 & pi27);
assign w920 = (w833 & ~w676) | (w833 & ~w274) | (~w676 & ~w274);
assign w921 = (pi27 & w409) | (pi27 & ~w218) | (w409 & ~w218);
assign w922 = w408 & w207;
assign w923 = (~pi27 & pi12) | (~pi27 & ~w762) | (pi12 & ~w762);
assign w924 = (w112 & ~w842) | (w112 & ~w217) | (~w842 & ~w217);
assign w925 = (w207 & w408) | (w207 & w585) | (w408 & w585);
assign w926 = pi49 & w930;
assign w927 = (w272 & w360) | (w272 & ~w218) | (w360 & ~w218);
assign w928 = ~pi28 & w71;
assign w929 = (pi28 & ~w826) | (pi28 & ~w337) | (~w826 & ~w337);
assign w930 = (~w590 & pi46) | (~w590 & ~w822) | (pi46 & ~w822);
assign w931 = (~pi12 & w526) | (~pi12 & ~w283) | (w526 & ~w283);
assign one = 1;
assign po00 = pi43;// level 0
assign po01 = pi59;// level 0
assign po02 = pi09;// level 0
assign po03 = pi29;// level 0
assign po04 = pi41;// level 0
assign po05 = pi57;// level 0
assign po06 = pi51;// level 0
assign po07 = pi52;// level 0
assign po08 = pi53;// level 0
assign po09 = pi48;// level 0
assign po10 = pi54;// level 0
assign po11 = pi55;// level 0
assign po12 = pi56;// level 0
assign po13 = ~pi60;// level 0
assign po14 = one;// level 0
assign po15 = pi61;// level 0
assign po16 = ~w282;// level 10
assign po17 = ~w181;// level 11
assign po18 = ~w140;// level 11
assign po19 = ~w420;// level 11
assign po20 = ~w675;// level 9
assign po21 = ~w388;// level 11
assign po22 = ~w649;// level 11
assign po23 = ~w795;// level 10
assign po24 = ~w897;// level 10
assign po25 = ~w332;// level 8
assign po26 = ~w652;// level 8
assign po27 = ~w371;// level 10
assign po28 = ~w672;// level 8
assign po29 = ~w402;// level 10
assign po30 = ~w879;// level 10
assign po31 = ~w787;// level 11
assign po32 = w56;// level 11
assign po33 = w228;// level 11
assign po34 = w118;// level 11
assign po35 = ~w83;// level 10
assign po36 = w0;// level 11
assign po37 = w191;// level 11
assign po38 = w58;// level 11
assign po39 = w808;// level 11
assign po40 = w619;// level 11
assign po41 = w735;// level 11
assign po42 = ~w184;// level 10
assign po43 = ~w8;// level 8
assign po44 = ~w230;// level 9
assign po45 = w289;// level 11
assign po46 = ~w215;// level 11
assign po47 = ~w137;// level 7
assign po48 = ~w618;// level 11
assign po49 = ~w542;// level 10
assign po50 = ~w633;// level 11
assign po51 = ~w815;// level 10
assign po52 = ~w702;// level 11
assign po53 = ~w502;// level 10
assign po54 = ~w390;// level 10
assign po55 = ~w547;// level 10
assign po56 = ~w687;// level 11
assign po57 = ~w145;// level 9
assign po58 = ~w847;// level 10
assign po59 = ~w611;// level 7
assign po60 = ~w599;// level 10
assign po61 = ~w711;// level 6
assign po62 = w504;// level 7
assign po63 = ~w814;// level 7
assign po64 = ~w869;// level 7
assign po65 = ~w577;// level 9
assign po66 = w436;// level 6
assign po67 = ~w423;// level 7
assign po68 = ~w884;// level 7
assign po69 = ~w584;// level 7
assign po70 = ~w854;// level 7
assign po71 = ~w583;// level 7
assign po72 = ~w698;// level 7
assign po73 = ~w785;// level 7
assign po74 = ~w305;// level 7
assign po75 = ~w149;// level 5
endmodule
