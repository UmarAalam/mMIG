//Written by the Majority Logic Package Fri May  1 00:06:25 2015
module top (
            pi00, pi01, pi02, pi03, pi04, pi05, pi06, pi07, pi08, pi09, pi10, pi11, pi12, pi13, pi14, pi15, pi16, pi17, pi18, pi19, pi20, pi21, pi22, pi23, pi24, pi25, pi26, pi27, pi28, pi29, pi30, pi31, pi32, pi33, pi34, pi35, pi36, pi37, pi38, pi39, pi40, pi41, pi42, pi43, pi44, pi45, pi46, pi47, pi48, pi49, pi50, pi51, pi52, pi53, pi54, pi55, pi56, pi57, pi58, pi59, pi60, pi61, pi62, pi63, 
            po000, po001, po002, po003, po004, po005, po006, po007, po008, po009, po010, po011, po012, po013, po014, po015, po016, po017, po018, po019, po020, po021, po022, po023, po024, po025, po026, po027, po028, po029, po030, po031, po032, po033, po034, po035, po036, po037, po038, po039, po040, po041, po042, po043, po044, po045, po046, po047, po048, po049, po050, po051, po052, po053, po054, po055, po056, po057, po058, po059, po060, po061, po062, po063, po064, po065, po066, po067, po068, po069, po070, po071, po072, po073, po074, po075, po076, po077, po078, po079, po080, po081, po082, po083, po084, po085, po086, po087, po088, po089, po090, po091, po092, po093, po094, po095, po096, po097, po098, po099, po100, po101, po102, po103, po104, po105, po106, po107, po108, po109, po110, po111, po112, po113, po114, po115, po116, po117, po118, po119, po120, po121, po122, po123, po124, po125, po126);
input pi00, pi01, pi02, pi03, pi04, pi05, pi06, pi07, pi08, pi09, pi10, pi11, pi12, pi13, pi14, pi15, pi16, pi17, pi18, pi19, pi20, pi21, pi22, pi23, pi24, pi25, pi26, pi27, pi28, pi29, pi30, pi31, pi32, pi33, pi34, pi35, pi36, pi37, pi38, pi39, pi40, pi41, pi42, pi43, pi44, pi45, pi46, pi47, pi48, pi49, pi50, pi51, pi52, pi53, pi54, pi55, pi56, pi57, pi58, pi59, pi60, pi61, pi62, pi63;
output po000, po001, po002, po003, po004, po005, po006, po007, po008, po009, po010, po011, po012, po013, po014, po015, po016, po017, po018, po019, po020, po021, po022, po023, po024, po025, po026, po027, po028, po029, po030, po031, po032, po033, po034, po035, po036, po037, po038, po039, po040, po041, po042, po043, po044, po045, po046, po047, po048, po049, po050, po051, po052, po053, po054, po055, po056, po057, po058, po059, po060, po061, po062, po063, po064, po065, po066, po067, po068, po069, po070, po071, po072, po073, po074, po075, po076, po077, po078, po079, po080, po081, po082, po083, po084, po085, po086, po087, po088, po089, po090, po091, po092, po093, po094, po095, po096, po097, po098, po099, po100, po101, po102, po103, po104, po105, po106, po107, po108, po109, po110, po111, po112, po113, po114, po115, po116, po117, po118, po119, po120, po121, po122, po123, po124, po125, po126;
wire one, v0, v1, v2, v3, v4, v5, v6, v7, v8, v9, v10, v11, v12, v13, v14, v15, v16, v17, v18, v19, v20, v21, v22, v23, v24, v25, v26, v27, v28, v29, v30, v31, v32, v33, v34, v35, v36, v37, v38, v39, v40, v41, v42, v43, v44, v45, v46, v47, v48, v49, v50, v51, v52, v53, v54, v55, v56, v57, v58, v59, v60, v61, v62, v63, v64, v65, v66, v67, v68, v69, v70, v71, v72, v73, v74, v75, v76, v77, v78, v79, v80, v81, v82, v83, v84, v85, v86, v87, v88, v89, v90, v91, v92, v93, v94, v95, v96, v97, v98, v99, v100, v101, v102, v103, v104, v105, v106, v107, v108, v109, v110, v111, v112, v113, v114, v115, v116, v117, v118, v119, v120, v121, v122, v123, v124, v125, v126, v127, v128, v129, v130, v131, v132, v133, v134, v135, v136, v137, v138, v139, v140, v141, v142, v143, v144, v145, v146, v147, v148, v149, v150, v151, v152, v153, v154, v155, v156, v157, v158, v159, v160, v161, v162, v163, v164, v165, v166, v167, v168, v169, v170, v171, v172, v173, v174, v175, v176, v177, v178, v179, v180, v181, v182, v183, v184, v185, v186, v187, v188, v189, v190, v191, v192, v193, v194, v195, v196, v197, v198, v199, v200, v201, v202, v203, v204, v205, v206, v207, v208, v209, v210, v211, v212, v213, v214, v215, v216, v217, v218, v219, v220, v221, v222, v223, v224, v225, v226, v227, v228, v229, v230, v231, v232, v233, v234, v235, v236, v237, v238, v239, v240, v241, v242, v243, v244, v245, v246, v247, v248, v249, v250, v251, v252, v253, v254, v255, v256, v257, v258, v259, v260, v261, v262, v263, v264, v265, v266, v267, v268, v269, v270, v271, v272, v273, v274, v275, v276, v277, v278, v279, v280, v281, v282, v283, v284, v285, v286, v287, v288, v289, v290, v291, v292, v293, v294, v295, v296, v297, v298, v299, v300, v301, v302, v303, v304, v305, v306, v307, v308, v309, v310, v311, v312, v313, v314, v315, v316, v317, v318, v319, v320, v321, v322, v323, v324, v325, v326, v327, v328, v329, v330, v331, v332, v333, v334, v335, v336, v337, v338, v339, v340, v341, v342, v343, v344, v345, v346, v347, v348, v349, v350, v351, v352, v353, v354, v355, v356, v357, v358, v359, v360, v361, v362, v363, v364, v365, v366, v367, v368, v369, v370, v371, v372, v373, v374, v375, v376, v377, v378, v379, v380, v381, v382, v383, v384, v385, v386, v387, v388, v389, v390, v391, v392, v393, v394, v395, v396, v397, v398, v399, v400, v401, v402, v403, v404, v405, v406, v407, v408, v409, v410, v411, v412, v413, v414, v415, v416, v417, v418, v419, v420, v421, v422, v423, v424, v425, v426, v427, v428, v429, v430, v431, v432, v433, v434, v435, v436, v437, v438, v439, v440, v441, v442, v443, v444, v445, v446, v447, v448, v449, v450, v451, v452, v453, v454, v455, v456, v457, v458, v459, v460, v461, v462, v463, v464, v465, v466, v467, v468, v469, v470, v471, v472, v473, v474, v475, v476, v477, v478, v479, v480, v481, v482, v483, v484, v485, v486, v487, v488, v489, v490, v491, v492, v493, v494, v495, v496, v497, v498, v499, v500, v501, v502, v503, v504, v505, v506, v507, v508, v509, v510, v511, v512, v513, v514, v515, v516, v517, v518, v519, v520, v521, v522, v523, v524, v525, v526, v527, v528, v529, v530, v531, v532, v533, v534, v535, v536, v537, v538, v539, v540, v541, v542, v543, v544, v545, v546, v547, v548, v549, v550, v551, v552, v553, v554, v555, v556, v557, v558, v559, v560, v561, v562, v563, v564, v565, v566, v567, v568, v569, v570, v571, v572, v573, v574, v575, v576, v577, v578, v579, v580, v581, v582, v583, v584, v585, v586, v587, v588, v589, v590, v591, v592, v593, v594, v595, v596, v597, v598, v599, v600, v601, v602, v603, v604, v605, v606, v607, v608, v609, v610, v611, v612, v613, v614, v615, v616, v617, v618, v619, v620, v621, v622, v623, v624, v625, v626, v627, v628, v629, v630, v631, v632, v633, v634, v635, v636, v637, v638, v639, v640, v641, v642, v643, v644, v645, v646, v647, v648, v649, v650, v651, v652, v653, v654, v655, v656, v657, v658, v659, v660, v661, v662, v663, v664, v665, v666, v667, v668, v669, v670, v671, v672, v673, v674, v675, v676, v677, v678, v679, v680, v681, v682, v683, v684, v685, v686, v687, v688, v689, v690, v691, v692, v693, v694, v695, v696, v697, v698, v699, v700, v701, v702, v703, v704, v705, v706, v707, v708, v709, v710, v711, v712, v713, v714, v715, v716, v717, v718, v719, v720, v721, v722, v723, v724, v725, v726, v727, v728, v729, v730, v731, v732, v733, v734, v735, v736, v737, v738, v739, v740, v741, v742, v743, v744, v745, v746, v747, v748, v749, v750, v751, v752, v753, v754, v755, v756, v757, v758, v759, v760, v761, v762, v763, v764, v765, v766, v767, v768, v769, v770, v771, v772, v773, v774, v775, v776, v777, v778, v779, v780, v781, v782, v783, v784, v785, v786, v787, v788, v789, v790, v791, v792, v793, v794, v795, v796, v797, v798, v799, v800, v801, v802, v803, v804, v805, v806, v807, v808, v809, v810, v811, v812, v813, v814, v815, v816, v817, v818, v819, v820, v821, v822, v823, v824, v825, v826, v827, v828, v829, v830, v831, v832, v833, v834, v835, v836, v837, v838, v839, v840, v841, v842, v843, v844, v845, v846, v847, v848, v849, v850, v851, v852, v853, v854, v855, v856, v857, v858, v859, v860, v861, v862, v863, v864, v865, v866, v867, v868, v869, v870, v871, v872, v873, v874, v875, v876, v877, v878, v879, v880, v881, v882, v883, v884, v885, v886, v887, v888, v889, v890, v891, v892, v893, v894, v895, v896, v897, v898, v899, v900, v901, v902, v903, v904, v905, v906, v907, v908, v909, v910, v911, v912, v913, v914, v915, v916, v917, v918, v919, v920, v921, v922, v923, v924, v925, v926, v927, v928, v929, v930, v931, v932, v933, v934, v935, v936, v937, v938, v939, v940, v941, v942, v943, v944, v945, v946, v947, v948, v949, v950, v951, v952, v953, v954, v955, v956, v957, v958, v959, v960, v961, v962, v963, v964, v965, v966, v967, v968, v969, v970, v971, v972, v973, v974, v975, v976, v977, v978, v979, v980, v981, v982, v983, v984, v985, v986, v987, v988, v989, v990, v991, v992, v993, v994, v995, v996, v997, v998, v999, v1000, v1001, v1002, v1003, v1004, v1005, v1006, v1007, v1008, v1009, v1010, v1011, v1012, v1013, v1014, v1015, v1016, v1017, v1018, v1019, v1020, v1021, v1022, v1023, v1024, v1025, v1026, v1027, v1028, v1029, v1030, v1031, v1032, v1033, v1034, v1035, v1036, v1037, v1038, v1039, v1040, v1041, v1042, v1043, v1044, v1045, v1046, v1047, v1048, v1049, v1050, v1051, v1052, v1053, v1054, v1055, v1056, v1057, v1058, v1059, v1060, v1061, v1062, v1063, v1064, v1065, v1066, v1067, v1068, v1069, v1070, v1071, v1072, v1073, v1074, v1075, v1076, v1077, v1078, v1079, v1080, v1081, v1082, v1083, v1084, v1085, v1086, v1087, v1088, v1089, v1090, v1091, v1092, v1093, v1094, v1095, v1096, v1097, v1098, v1099, v1100, v1101, v1102, v1103, v1104, v1105, v1106, v1107, v1108, v1109, v1110, v1111, v1112, v1113, v1114, v1115, v1116, v1117, v1118, v1119, v1120, v1121, v1122, v1123, v1124, v1125, v1126, v1127, v1128, v1129, v1130, v1131, v1132, v1133, v1134, v1135, v1136, v1137, v1138, v1139, v1140, v1141, v1142, v1143, v1144, v1145, v1146, v1147, v1148, v1149, v1150, v1151, v1152, v1153, v1154, v1155, v1156, v1157, v1158, v1159, v1160, v1161, v1162, v1163, v1164, v1165, v1166, v1167, v1168, v1169, v1170, v1171, v1172, v1173, v1174, v1175, v1176, v1177, v1178, v1179, v1180, v1181, v1182, v1183, v1184, v1185, v1186, v1187, v1188, v1189, v1190, v1191, v1192, v1193, v1194, v1195, v1196, v1197, v1198, v1199, v1200, v1201, v1202, v1203, v1204, v1205, v1206, v1207, v1208, v1209, v1210, v1211, v1212, v1213, v1214, v1215, v1216, v1217, v1218, v1219, v1220, v1221, v1222, v1223, v1224, v1225, v1226, v1227, v1228, v1229, v1230, v1231, v1232, v1233, v1234, v1235, v1236, v1237, v1238, v1239, v1240, v1241, v1242, v1243, v1244, v1245, v1246, v1247, v1248, v1249, v1250, v1251, v1252, v1253, v1254, v1255, v1256, v1257, v1258, v1259, v1260, v1261, v1262, v1263, v1264, v1265, v1266, v1267, v1268, v1269, v1270, v1271, v1272, v1273, v1274, v1275, v1276, v1277, v1278, v1279, v1280, v1281, v1282, v1283, v1284, v1285, v1286, v1287, v1288, v1289, v1290, v1291, v1292, v1293, v1294, v1295, v1296, v1297, v1298, v1299, v1300, v1301, v1302, v1303, v1304, v1305, v1306, v1307, v1308, v1309, v1310, v1311, v1312, v1313, v1314, v1315, v1316, v1317, v1318, v1319, v1320, v1321, v1322, v1323, v1324, v1325, v1326, v1327, v1328, v1329, v1330, v1331, v1332, v1333, v1334, v1335, v1336, v1337, v1338, v1339, v1340, v1341, v1342, v1343, v1344, v1345, v1346, v1347, v1348, v1349, v1350, v1351, v1352, v1353, v1354, v1355, v1356, v1357, v1358, v1359, v1360, v1361, v1362, v1363, v1364, v1365, v1366, v1367, v1368, v1369, v1370, v1371, v1372, v1373, v1374, v1375, v1376, v1377, v1378, v1379, v1380, v1381, v1382, v1383, v1384, v1385, v1386, v1387, v1388, v1389, v1390, v1391, v1392, v1393, v1394, v1395, v1396, v1397, v1398, v1399, v1400, v1401, v1402, v1403, v1404, v1405, v1406, v1407, v1408, v1409, v1410, v1411, v1412, v1413, v1414, v1415, v1416, v1417, v1418, v1419, v1420, v1421, v1422, v1423, v1424, v1425, v1426, v1427, v1428, v1429, v1430, v1431, v1432, v1433, v1434, v1435, v1436, v1437, v1438, v1439, v1440, v1441, v1442, v1443, v1444, v1445, v1446, v1447, v1448, v1449, v1450, v1451, v1452, v1453, v1454, v1455, v1456, v1457, v1458, v1459, v1460, v1461, v1462, v1463, v1464, v1465, v1466, v1467, v1468, v1469, v1470, v1471, v1472, v1473, v1474, v1475, v1476, v1477, v1478, v1479, v1480, v1481, v1482, v1483, v1484, v1485, v1486, v1487, v1488, v1489, v1490, v1491, v1492, v1493, v1494, v1495, v1496, v1497, v1498, v1499, v1500, v1501, v1502, v1503, v1504, v1505, v1506, v1507, v1508, v1509, v1510, v1511, v1512, v1513, v1514, v1515, v1516, v1517, v1518, v1519, v1520, v1521, v1522, v1523, v1524, v1525, v1526, v1527, v1528, v1529, v1530, v1531, v1532, v1533, v1534, v1535, v1536, v1537, v1538, v1539, v1540, v1541, v1542, v1543, v1544, v1545, v1546, v1547, v1548, v1549, v1550, v1551, v1552, v1553, v1554, v1555, v1556, v1557, v1558, v1559, v1560, v1561, v1562, v1563, v1564, v1565, v1566, v1567, v1568, v1569, v1570, v1571, v1572, v1573, v1574, v1575, v1576, v1577, v1578, v1579, v1580, v1581, v1582, v1583, v1584, v1585, v1586, v1587, v1588, v1589, v1590, v1591, v1592, v1593, v1594, v1595, v1596, v1597, v1598, v1599, v1600, v1601, v1602, v1603, v1604, v1605, v1606, v1607, v1608, v1609, v1610, v1611, v1612, v1613, v1614, v1615, v1616, v1617, v1618, v1619, v1620, v1621, v1622, v1623, v1624, v1625, v1626, v1627, v1628, v1629, v1630, v1631, v1632, v1633, v1634, v1635, v1636, v1637, v1638, v1639, v1640, v1641, v1642, v1643, v1644, v1645, v1646, v1647, v1648, v1649, v1650, v1651, v1652, v1653, v1654, v1655, v1656, v1657, v1658, v1659, v1660, v1661, v1662, v1663, v1664, v1665, v1666, v1667, v1668, v1669, v1670, v1671, v1672, v1673, v1674, v1675, v1676, v1677, v1678, v1679, v1680, v1681, v1682, v1683, v1684, v1685, v1686, v1687, v1688, v1689, v1690, v1691, v1692, v1693, v1694, v1695, v1696, v1697, v1698, v1699, v1700, v1701, v1702, v1703, v1704, v1705, v1706, v1707, v1708, v1709, v1710, v1711, v1712, v1713, v1714, v1715, v1716, v1717, v1718, v1719, v1720, v1721, v1722, v1723, v1724, v1725, v1726, v1727, v1728, v1729, v1730, v1731, v1732, v1733, v1734, v1735, v1736, v1737, v1738, v1739, v1740, v1741, v1742, v1743, v1744, v1745, v1746, v1747, v1748, v1749, v1750, v1751, v1752, v1753, v1754, v1755, v1756, v1757, v1758, v1759, v1760, v1761, v1762, v1763, v1764, v1765, v1766, v1767, v1768, v1769, v1770, v1771, v1772, v1773, v1774, v1775, v1776, v1777, v1778, v1779, v1780, v1781, v1782, v1783, v1784, v1785, v1786, v1787, v1788, v1789, v1790, v1791, v1792, v1793, v1794, v1795, v1796, v1797, v1798, v1799, v1800, v1801, v1802, v1803, v1804, v1805, v1806, v1807, v1808, v1809, v1810, v1811, v1812, v1813, v1814, v1815, v1816, v1817, v1818, v1819, v1820, v1821, v1822, v1823, v1824, v1825, v1826, v1827, v1828, v1829, v1830, v1831, v1832, v1833, v1834, v1835, v1836, v1837, v1838, v1839, v1840, v1841, v1842, v1843, v1844, v1845, v1846, v1847, v1848, v1849, v1850, v1851, v1852, v1853, v1854, v1855, v1856, v1857, v1858, v1859, v1860, v1861, v1862, v1863, v1864, v1865, v1866, v1867, v1868, v1869, v1870, v1871, v1872, v1873, v1874, v1875, v1876, v1877, v1878, v1879, v1880, v1881, v1882, v1883, v1884, v1885, v1886, v1887, v1888, v1889, v1890, v1891, v1892, v1893, v1894, v1895, v1896, v1897, v1898, v1899, v1900, v1901, v1902, v1903, v1904, v1905, v1906, v1907, v1908, v1909, v1910, v1911, v1912, v1913, v1914, v1915, v1916, v1917, v1918, v1919, v1920, v1921, v1922, v1923, v1924, v1925, v1926, v1927, v1928, v1929, v1930, v1931, v1932, v1933, v1934, v1935, v1936, v1937, v1938, v1939, v1940, v1941, v1942, v1943, v1944, v1945, v1946, v1947, v1948, v1949, v1950, v1951, v1952, v1953, v1954, v1955, v1956, v1957, v1958, v1959, v1960, v1961, v1962, v1963, v1964, v1965, v1966, v1967, v1968, v1969, v1970, v1971, v1972, v1973, v1974, v1975, v1976, v1977, v1978, v1979, v1980, v1981, v1982, v1983, v1984, v1985, v1986, v1987, v1988, v1989, v1990, v1991, v1992, v1993, v1994, v1995, v1996, v1997, v1998, v1999, v2000, v2001, v2002, v2003, v2004, v2005, v2006, v2007, v2008, v2009, v2010, v2011, v2012, v2013, v2014, v2015, v2016, v2017, v2018, v2019, v2020, v2021, v2022, v2023, v2024, v2025, v2026, v2027, v2028, v2029, v2030, v2031, v2032, v2033, v2034, v2035, v2036, v2037, v2038, v2039, v2040, v2041, v2042, v2043, v2044, v2045, v2046, v2047, v2048, v2049, v2050, v2051, v2052, v2053, v2054, v2055, v2056, v2057, v2058, v2059, v2060, v2061, v2062, v2063, v2064, v2065, v2066, v2067, v2068, v2069, v2070, v2071, v2072, v2073, v2074, v2075, v2076, v2077, v2078, v2079, v2080, v2081, v2082, v2083, v2084, v2085, v2086, v2087, v2088, v2089, v2090, v2091, v2092, v2093, v2094, v2095, v2096, v2097, v2098, v2099, v2100, v2101, v2102, v2103, v2104, v2105, v2106, v2107, v2108, v2109, v2110, v2111, v2112, v2113, v2114, v2115, v2116, v2117, v2118, v2119, v2120, v2121, v2122, v2123, v2124, v2125, v2126, v2127, v2128, v2129, v2130, v2131, v2132, v2133, v2134, v2135, v2136, v2137, v2138, v2139, v2140, v2141, v2142, v2143, v2144, v2145, v2146, v2147, v2148, v2149, v2150, v2151, v2152, v2153, v2154, v2155, v2156, v2157, v2158, v2159, v2160, v2161, v2162, v2163, v2164, v2165, v2166, v2167, v2168, v2169, v2170, v2171, v2172, v2173, v2174, v2175, v2176, v2177, v2178, v2179, v2180, v2181, v2182, v2183, v2184, v2185, v2186, v2187, v2188, v2189, v2190, v2191, v2192, v2193, v2194, v2195, v2196, v2197, v2198, v2199, v2200, v2201, v2202, v2203, v2204, v2205, v2206, v2207, v2208, v2209, v2210, v2211, v2212, v2213, v2214, v2215, v2216, v2217, v2218, v2219, v2220, v2221, v2222, v2223, v2224, v2225, v2226, v2227, v2228, v2229, v2230, v2231, v2232, v2233, v2234, v2235, v2236, v2237, v2238, v2239, v2240, v2241, v2242, v2243, v2244, v2245, v2246, v2247, v2248, v2249, v2250, v2251, v2252, v2253, v2254, v2255, v2256, v2257, v2258, v2259, v2260, v2261, v2262, v2263, v2264, v2265, v2266, v2267, v2268, v2269, v2270, v2271, v2272, v2273, v2274, v2275, v2276, v2277, v2278, v2279, v2280, v2281, v2282, v2283, v2284, v2285, v2286, v2287, v2288, v2289, v2290, v2291, v2292, v2293, v2294, v2295, v2296, v2297, v2298, v2299, v2300, v2301, v2302, v2303, v2304, v2305, v2306, v2307, v2308, v2309, v2310, v2311, v2312, v2313, v2314, v2315, v2316, v2317, v2318, v2319, v2320, v2321, v2322, v2323, v2324, v2325, v2326, v2327, v2328, v2329, v2330, v2331, v2332, v2333, v2334, v2335, v2336, v2337, v2338, v2339, v2340, v2341, v2342, v2343, v2344, v2345, v2346, v2347, v2348, v2349, v2350, v2351, v2352, v2353, v2354, v2355, v2356, v2357, v2358, v2359, v2360, v2361, v2362, v2363, v2364, v2365, v2366, v2367, v2368, v2369, v2370, v2371, v2372, v2373, v2374, v2375, v2376, v2377, v2378, v2379, v2380, v2381, v2382, v2383, v2384, v2385, v2386, v2387, v2388, v2389, v2390, v2391, v2392, v2393, v2394, v2395, v2396, v2397, v2398, v2399, v2400, v2401, v2402, v2403, v2404, v2405, v2406, v2407, v2408, v2409, v2410, v2411, v2412, v2413, v2414, v2415, v2416, v2417, v2418, v2419, v2420, v2421, v2422, v2423, v2424, v2425, v2426, v2427, v2428, v2429, v2430, v2431, v2432, v2433, v2434, v2435, v2436, v2437, v2438, v2439, v2440, v2441, v2442, v2443, v2444, v2445, v2446, v2447, v2448, v2449, v2450, v2451, v2452, v2453, v2454, v2455, v2456, v2457, v2458, v2459, v2460, v2461, v2462, v2463, v2464, v2465, v2466, v2467, v2468, v2469, v2470, v2471, v2472, v2473, v2474, v2475, v2476, v2477, v2478, v2479, v2480, v2481, v2482, v2483, v2484, v2485, v2486, v2487, v2488, v2489, v2490, v2491, v2492, v2493, v2494, v2495, v2496, v2497, v2498, v2499, v2500, v2501, v2502, v2503, v2504, v2505, v2506, v2507, v2508, v2509, v2510, v2511, v2512, v2513, v2514, v2515, v2516, v2517, v2518, v2519, v2520, v2521, v2522, v2523, v2524, v2525, v2526, v2527, v2528, v2529, v2530, v2531, v2532, v2533, v2534, v2535, v2536, v2537, v2538, v2539, v2540, v2541, v2542, v2543, v2544, v2545, v2546, v2547, v2548, v2549, v2550, v2551, v2552, v2553, v2554, v2555, v2556, v2557, v2558, v2559, v2560, v2561, v2562, v2563, v2564, v2565, v2566, v2567, v2568, v2569, v2570, v2571, v2572, v2573, v2574, v2575, v2576, v2577, v2578, v2579, v2580, v2581, v2582, v2583, v2584, v2585, v2586, v2587, v2588, v2589, v2590, v2591, v2592, v2593, v2594, v2595, v2596, v2597, v2598, v2599, v2600, v2601, v2602, v2603, v2604, v2605, v2606, v2607, v2608, v2609, v2610, v2611, v2612, v2613, v2614, v2615, v2616, v2617, v2618, v2619, v2620, v2621, v2622, v2623, v2624, v2625, v2626, v2627, v2628, v2629, v2630, v2631, v2632, v2633, v2634, v2635, v2636, v2637, v2638, v2639, v2640, v2641, v2642, v2643, v2644, v2645, v2646, v2647, v2648, v2649, v2650, v2651, v2652, v2653, v2654, v2655, v2656, v2657, v2658, v2659, v2660, v2661, v2662, v2663, v2664, v2665, v2666, v2667, v2668, v2669, v2670, v2671, v2672, v2673, v2674, v2675, v2676, v2677, v2678, v2679, v2680, v2681, v2682, v2683, v2684, v2685, v2686, v2687, v2688, v2689, v2690, v2691, v2692, v2693, v2694, v2695, v2696, v2697, v2698, v2699, v2700, v2701, v2702, v2703, v2704, v2705, v2706, v2707, v2708, v2709, v2710, v2711, v2712, v2713, v2714, v2715, v2716, v2717, v2718, v2719, v2720, v2721, v2722, v2723, v2724, v2725, v2726, v2727, v2728, v2729, v2730, v2731, v2732, v2733, v2734, v2735, v2736, v2737, v2738, v2739, v2740, v2741, v2742, v2743, v2744, v2745, v2746, v2747, v2748, v2749, v2750, v2751, v2752, v2753, v2754, v2755, v2756, v2757, v2758, v2759, v2760, v2761, v2762, v2763, v2764, v2765, v2766, v2767, v2768, v2769, v2770, v2771, v2772, v2773, v2774, v2775, v2776, v2777, v2778, v2779, v2780, v2781, v2782, v2783, v2784, v2785, v2786, v2787, v2788, v2789, v2790, v2791, v2792, v2793, v2794, v2795, v2796, v2797, v2798, v2799, v2800, v2801, v2802, v2803, v2804, v2805, v2806, v2807, v2808, v2809, v2810, v2811, v2812, v2813, v2814, v2815, v2816, v2817, v2818, v2819, v2820, v2821, v2822, v2823, v2824, v2825, v2826, v2827, v2828, v2829, v2830, v2831, v2832, v2833, v2834, v2835, v2836, v2837, v2838, v2839, v2840, v2841, v2842, v2843, v2844, v2845, v2846, v2847, v2848, v2849, v2850, v2851, v2852, v2853, v2854, v2855, v2856, v2857, v2858, v2859, v2860, v2861, v2862, v2863, v2864, v2865, v2866, v2867, v2868, v2869, v2870, v2871, v2872, v2873, v2874, v2875, v2876, v2877, v2878, v2879, v2880, v2881, v2882, v2883, v2884, v2885, v2886, v2887, v2888, v2889, v2890, v2891, v2892, v2893, v2894, v2895, v2896, v2897, v2898, v2899, v2900, v2901, v2902, v2903, v2904, v2905, v2906, v2907, v2908, v2909, v2910, v2911, v2912, v2913, v2914, v2915, v2916, v2917, v2918, v2919, v2920, v2921, v2922, v2923, v2924, v2925, v2926, v2927, v2928, v2929, v2930, v2931, v2932, v2933, v2934, v2935, v2936, v2937, v2938, v2939, v2940, v2941, v2942, v2943, v2944, v2945, v2946, v2947, v2948, v2949, v2950, v2951, v2952, v2953, v2954, v2955, v2956, v2957, v2958, v2959, v2960, v2961, v2962, v2963, v2964, v2965, v2966, v2967, v2968, v2969, v2970, v2971, v2972, v2973, v2974, v2975, v2976, v2977, v2978, v2979, v2980, v2981, v2982, v2983, v2984, v2985, v2986, v2987, v2988, v2989, v2990, v2991, v2992, v2993, v2994, v2995, v2996, v2997, v2998, v2999, v3000, v3001, v3002, v3003, v3004, v3005, v3006, v3007, v3008, v3009, v3010, v3011, v3012, v3013, v3014, v3015, v3016, v3017, v3018, v3019, v3020, v3021, v3022, v3023, v3024, v3025, v3026, v3027, v3028, v3029, v3030, v3031, v3032, v3033, v3034, v3035, v3036, v3037, v3038, v3039, v3040, v3041, v3042, v3043, v3044, v3045, v3046, v3047, v3048, v3049, v3050, v3051, v3052, v3053, v3054, v3055, v3056, v3057, v3058, v3059, v3060, v3061, v3062, v3063, v3064, v3065, v3066, v3067, v3068, v3069, v3070, v3071, v3072, v3073, v3074, v3075, v3076, v3077, v3078, v3079, v3080, v3081, v3082, v3083, v3084, v3085, v3086, v3087, v3088, v3089, v3090, v3091, v3092, v3093, v3094, v3095, v3096, v3097, v3098, v3099, v3100, v3101, v3102, v3103, v3104, v3105, v3106, v3107, v3108, v3109, v3110, v3111, v3112, v3113, v3114, v3115, v3116, v3117, v3118, v3119, v3120, v3121, v3122, v3123, v3124, v3125, v3126, v3127, v3128, v3129, v3130, v3131, v3132, v3133, v3134, v3135, v3136, v3137, v3138, v3139, v3140, v3141, v3142, v3143, v3144, v3145, v3146, v3147, v3148, v3149, v3150, v3151, v3152, v3153, v3154, v3155, v3156, v3157, v3158, v3159, v3160, v3161, v3162, v3163, v3164, v3165, v3166, v3167, v3168, v3169, v3170, v3171, v3172, v3173, v3174, v3175, v3176, v3177, v3178, v3179, v3180, v3181, v3182, v3183, v3184, v3185, v3186, v3187, v3188, v3189, v3190, v3191, v3192, v3193, v3194, v3195, v3196, v3197, v3198, v3199, v3200, v3201, v3202, v3203, v3204, v3205, v3206, v3207, v3208, v3209, v3210, v3211, v3212, v3213, v3214, v3215, v3216, v3217, v3218, v3219, v3220, v3221, v3222, v3223, v3224, v3225, v3226, v3227, v3228, v3229, v3230, v3231, v3232, v3233, v3234, v3235, v3236, v3237, v3238, v3239, v3240, v3241, v3242, v3243, v3244, v3245, v3246, v3247, v3248, v3249, v3250, v3251, v3252, v3253, v3254, v3255, v3256, v3257, v3258, v3259, v3260, v3261, v3262, v3263, v3264, v3265, v3266, v3267, v3268, v3269, v3270, v3271, v3272, v3273, v3274, v3275, v3276, v3277, v3278, v3279, v3280, v3281, v3282, v3283, v3284, v3285, v3286, v3287, v3288, v3289, v3290, v3291, v3292, v3293, v3294, v3295, v3296, v3297, v3298, v3299, v3300, v3301, v3302, v3303, v3304, v3305, v3306, v3307, v3308, v3309, v3310, v3311, v3312, v3313, v3314, v3315, v3316, v3317, v3318, v3319, v3320, v3321, v3322, v3323, v3324, v3325, v3326, v3327, v3328, v3329, v3330, v3331, v3332, v3333, v3334, v3335, v3336, v3337, v3338, v3339, v3340, v3341, v3342, v3343, v3344, v3345, v3346, v3347, v3348, v3349, v3350, v3351, v3352, v3353, v3354, v3355, v3356, v3357, v3358, v3359, v3360, v3361, v3362, v3363, v3364, v3365, v3366, v3367, v3368, v3369, v3370, v3371, v3372, v3373, v3374, v3375, v3376, v3377, v3378, v3379, v3380, v3381, v3382, v3383, v3384, v3385, v3386, v3387, v3388, v3389, v3390, v3391, v3392, v3393, v3394, v3395, v3396, v3397, v3398, v3399, v3400, v3401, v3402, v3403, v3404, v3405, v3406, v3407, v3408, v3409, v3410, v3411, v3412, v3413, v3414, v3415, v3416, v3417, v3418, v3419, v3420, v3421, v3422, v3423, v3424, v3425, v3426, v3427, v3428, v3429, v3430, v3431, v3432, v3433, v3434, v3435, v3436, v3437, v3438, v3439, v3440, v3441, v3442, v3443, v3444, v3445, v3446, v3447, v3448, v3449, v3450, v3451, v3452, v3453, v3454, v3455, v3456, v3457, v3458, v3459, v3460, v3461, v3462, v3463, v3464, v3465, v3466, v3467, v3468, v3469, v3470, v3471, v3472, v3473, v3474, v3475, v3476, v3477, v3478, v3479, v3480, v3481, v3482, v3483, v3484, v3485, v3486, v3487, v3488, v3489, v3490, v3491, v3492, v3493, v3494, v3495, v3496, v3497, v3498, v3499, v3500, v3501, v3502, v3503, v3504, v3505, v3506, v3507, v3508, v3509, v3510, v3511, v3512, v3513, v3514, v3515, v3516, v3517, v3518, v3519, v3520, v3521, v3522, v3523, v3524, v3525, v3526, v3527, v3528, v3529, v3530, v3531, v3532, v3533, v3534, v3535, v3536, v3537, v3538, v3539, v3540, v3541, v3542, v3543, v3544, v3545, v3546, v3547, v3548, v3549, v3550, v3551, v3552, v3553, v3554, v3555, v3556, v3557, v3558, v3559, v3560, v3561, v3562, v3563, v3564, v3565, v3566, v3567, v3568, v3569, v3570, v3571, v3572, v3573, v3574, v3575, v3576, v3577, v3578, v3579, v3580, v3581, v3582, v3583, v3584, v3585, v3586, v3587, v3588, v3589, v3590, v3591, v3592, v3593, v3594, v3595, v3596, v3597, v3598, v3599, v3600, v3601, v3602, v3603, v3604, v3605, v3606, v3607, v3608, v3609, v3610, v3611, v3612, v3613, v3614, v3615, v3616, v3617, v3618, v3619, v3620, v3621, v3622, v3623, v3624, v3625, v3626, v3627, v3628, v3629, v3630, v3631, v3632, v3633, v3634, v3635, v3636, v3637, v3638, v3639, v3640, v3641, v3642, v3643, v3644, v3645, v3646, v3647, v3648, v3649, v3650, v3651, v3652, v3653, v3654, v3655, v3656, v3657, v3658, v3659, v3660, v3661, v3662, v3663, v3664, v3665, v3666, v3667, v3668, v3669, v3670, v3671, v3672, v3673, v3674, v3675, v3676, v3677, v3678, v3679, v3680, v3681, v3682, v3683, v3684, v3685, v3686, v3687, v3688, v3689, v3690, v3691, v3692, v3693, v3694, v3695, v3696, v3697, v3698, v3699, v3700, v3701, v3702, v3703, v3704, v3705, v3706, v3707, v3708, v3709, v3710, v3711, v3712, v3713, v3714, v3715, v3716, v3717, v3718, v3719, v3720, v3721, v3722, v3723, v3724, v3725, v3726, v3727, v3728, v3729, v3730, v3731, v3732, v3733, v3734, v3735, v3736, v3737, v3738, v3739, v3740, v3741, v3742, v3743, v3744, v3745, v3746, v3747, v3748, v3749, v3750, v3751, v3752, v3753, v3754, v3755, v3756, v3757, v3758, v3759, v3760, v3761, v3762, v3763, v3764, v3765, v3766, v3767, v3768, v3769, v3770, v3771, v3772, v3773, v3774, v3775, v3776, v3777, v3778, v3779, v3780, v3781, v3782, v3783, v3784, v3785, v3786, v3787, v3788, v3789, v3790, v3791, v3792, v3793, v3794, v3795, v3796, v3797, v3798, v3799, v3800, v3801, v3802, v3803, v3804, v3805, v3806, v3807, v3808, v3809, v3810, v3811, v3812, v3813, v3814, v3815, v3816, v3817, v3818, v3819, v3820, v3821, v3822, v3823, v3824, v3825, v3826, v3827, v3828, v3829, v3830, v3831, v3832, v3833, v3834, v3835, v3836, v3837, v3838, v3839, v3840, v3841, v3842, v3843, v3844, v3845, v3846, v3847, v3848, v3849, v3850, v3851, v3852, v3853, v3854, v3855, v3856, v3857, v3858, v3859, v3860, v3861, v3862, v3863, v3864, v3865, v3866, v3867, v3868, v3869, v3870, v3871, v3872, v3873, v3874, v3875, v3876, v3877, v3878, v3879, v3880, v3881, v3882, v3883, v3884, v3885, v3886, v3887, v3888, v3889, v3890, v3891, v3892, v3893, v3894, v3895, v3896, v3897, v3898, v3899, v3900, v3901, v3902, v3903, v3904, v3905, v3906, v3907, v3908, v3909, v3910, v3911, v3912, v3913, v3914, v3915, v3916, v3917, v3918, v3919, v3920, v3921, v3922, v3923, v3924, v3925, v3926, v3927, v3928, v3929, v3930, v3931, v3932, v3933, v3934, v3935, v3936, v3937, v3938, v3939, v3940, v3941, v3942, v3943, v3944, v3945, v3946, v3947, v3948, v3949, v3950, v3951, v3952, v3953, v3954, v3955, v3956, v3957, v3958, v3959, v3960, v3961, v3962, v3963, v3964, v3965, v3966, v3967, v3968, v3969, v3970, v3971, v3972, v3973, v3974, v3975, v3976, v3977, v3978, v3979, v3980, v3981, v3982, v3983, v3984, v3985, v3986, v3987, v3988, v3989, v3990, v3991, v3992, v3993, v3994, v3995, v3996, v3997, v3998, v3999, v4000, v4001, v4002, v4003, v4004, v4005, v4006, v4007, v4008, v4009, v4010, v4011, v4012, v4013, v4014, v4015, v4016, v4017, v4018, v4019, v4020, v4021, v4022, v4023, v4024, v4025, v4026, v4027, v4028, v4029, v4030, v4031, v4032, v4033, v4034, v4035, v4036, v4037, v4038, v4039, v4040, v4041, v4042, v4043, v4044, v4045, v4046, v4047, v4048, v4049, v4050, v4051, v4052, v4053, v4054, v4055, v4056, v4057, v4058, v4059, v4060, v4061, v4062, v4063, v4064, v4065, v4066, v4067, v4068, v4069, v4070, v4071, v4072, v4073, v4074, v4075, v4076, v4077, v4078, v4079, v4080, v4081, v4082, v4083, v4084, v4085, v4086, v4087, v4088, v4089, v4090, v4091, v4092, v4093, v4094, v4095, v4096, v4097, v4098, v4099, v4100, v4101, v4102, v4103, v4104, v4105, v4106, v4107, v4108, v4109, v4110, v4111, v4112, v4113, v4114, v4115, v4116, v4117, v4118, v4119, v4120, v4121, v4122, v4123, v4124, v4125, v4126, v4127, v4128, v4129, v4130, v4131, v4132, v4133, v4134, v4135, v4136, v4137, v4138, v4139, v4140, v4141, v4142, v4143, v4144, v4145, v4146, v4147, v4148, v4149, v4150, v4151, v4152, v4153, v4154, v4155, v4156, v4157, v4158, v4159, v4160, v4161, v4162, v4163, v4164, v4165, v4166, v4167, v4168, v4169, v4170, v4171, v4172, v4173, v4174, v4175, v4176, v4177, v4178, v4179, v4180, v4181, v4182, v4183, v4184, v4185, v4186, v4187, v4188, v4189, v4190, v4191, v4192, v4193, v4194, v4195, v4196, v4197, v4198, v4199, v4200, v4201, v4202, v4203, v4204, v4205, v4206, v4207, v4208, v4209, v4210, v4211, v4212, v4213, v4214, v4215, v4216, v4217, v4218, v4219, v4220, v4221, v4222, v4223, v4224, v4225, v4226, v4227, v4228, v4229, v4230, v4231, v4232, v4233, v4234, v4235, v4236, v4237, v4238, v4239, v4240, v4241, v4242, v4243, v4244, v4245, v4246, v4247, v4248, v4249, v4250, v4251, v4252, v4253, v4254, v4255, v4256, v4257, v4258, v4259, v4260, v4261, v4262, v4263, v4264, v4265, v4266, v4267, v4268, v4269, v4270, v4271, v4272, v4273, v4274, v4275, v4276, v4277, v4278, v4279, v4280, v4281, v4282, v4283, v4284, v4285, v4286, v4287, v4288, v4289, v4290, v4291, v4292, v4293, v4294, v4295, v4296, v4297, v4298, v4299, v4300, v4301, v4302, v4303, v4304, v4305, v4306, v4307, v4308, v4309, v4310, v4311, v4312, v4313, v4314, v4315, v4316, v4317, v4318, v4319, v4320, v4321, v4322, v4323, v4324, v4325, v4326, v4327, v4328, v4329, v4330, v4331, v4332, v4333, v4334, v4335, v4336, v4337, v4338, v4339, v4340, v4341, v4342, v4343, v4344, v4345, v4346, v4347, v4348, v4349, v4350, v4351, v4352, v4353, v4354, v4355, v4356, v4357, v4358, v4359, v4360, v4361, v4362, v4363, v4364, v4365, v4366, v4367, v4368, v4369, v4370, v4371, v4372, v4373, v4374, v4375, v4376, v4377, v4378, v4379, v4380, v4381, v4382, v4383, v4384, v4385, v4386, v4387, v4388, v4389, v4390, v4391, v4392, v4393, v4394, v4395, v4396, v4397, v4398, v4399, v4400, v4401, v4402, v4403, v4404, v4405, v4406, v4407, v4408, v4409, v4410, v4411, v4412, v4413, v4414, v4415, v4416, v4417, v4418, v4419, v4420, v4421, v4422, v4423, v4424, v4425, v4426, v4427, v4428, v4429, v4430, v4431, v4432, v4433, v4434, v4435, v4436, v4437, v4438, v4439, v4440, v4441, v4442, v4443, v4444, v4445, v4446, v4447, v4448, v4449, v4450, v4451, v4452, v4453, v4454, v4455, v4456, v4457, v4458, v4459, v4460, v4461, v4462, v4463, v4464, v4465, v4466, v4467, v4468, v4469, v4470, v4471, v4472, v4473, v4474, v4475, v4476, v4477, v4478, v4479, v4480, v4481, v4482, v4483, v4484, v4485, v4486, v4487, v4488, v4489, v4490, v4491, v4492, v4493, v4494, v4495, v4496, v4497, v4498, v4499, v4500, v4501, v4502, v4503, v4504, v4505, v4506, v4507, v4508, v4509, v4510, v4511, v4512, v4513, v4514, v4515, v4516, v4517, v4518, v4519, v4520, v4521, v4522, v4523, v4524, v4525, v4526, v4527, v4528, v4529, v4530, v4531, v4532, v4533, v4534, v4535, v4536, v4537, v4538, v4539, v4540, v4541, v4542, v4543, v4544, v4545, v4546, v4547, v4548, v4549, v4550, v4551, v4552, v4553, v4554, v4555, v4556, v4557, v4558, v4559, v4560, v4561, v4562, v4563, v4564, v4565, v4566, v4567, v4568, v4569, v4570, v4571, v4572, v4573, v4574, v4575, v4576, v4577, v4578, v4579, v4580, v4581, v4582, v4583, v4584, v4585, v4586, v4587, v4588, v4589, v4590, v4591, v4592, v4593, v4594, v4595, v4596, v4597, v4598, v4599, v4600, v4601, v4602, v4603, v4604, v4605, v4606, v4607, v4608, v4609, v4610, v4611, v4612, v4613, v4614, v4615, v4616, v4617, v4618, v4619, v4620, v4621, v4622, v4623, v4624, v4625, v4626, v4627, v4628, v4629, v4630, v4631, v4632, v4633, v4634, v4635, v4636, v4637, v4638, v4639, v4640, v4641, v4642, v4643, v4644, v4645, v4646, v4647, v4648, v4649, v4650, v4651, v4652, v4653, v4654, v4655, v4656, v4657, v4658, v4659, v4660, v4661, v4662, v4663, v4664, v4665, v4666, v4667, v4668, v4669, v4670, v4671, v4672, v4673, v4674, v4675, v4676, v4677, v4678, v4679, v4680, v4681, v4682, v4683, v4684, v4685, v4686, v4687, v4688, v4689, v4690, v4691, v4692, v4693, v4694, v4695, v4696, v4697, v4698, v4699, v4700, v4701, v4702, v4703, v4704, v4705, v4706, v4707, v4708, v4709, v4710, v4711, v4712, v4713, v4714, v4715, v4716, v4717, v4718, v4719, v4720, v4721, v4722, v4723, v4724, v4725, v4726, v4727, v4728, v4729, v4730, v4731, v4732, v4733, v4734, v4735, v4736, v4737, v4738, v4739, v4740, v4741, v4742, v4743, v4744, v4745, v4746, v4747, v4748, v4749, v4750, v4751, v4752, v4753, v4754, v4755, v4756, v4757, v4758, v4759, v4760, v4761, v4762, v4763, v4764, v4765, v4766, v4767, v4768, v4769, v4770, v4771, v4772, v4773, v4774, v4775, v4776, v4777, v4778, v4779, v4780, v4781, v4782, v4783, v4784, v4785, v4786, v4787, v4788, v4789, v4790, v4791, v4792, v4793, v4794, v4795, v4796, v4797, v4798, v4799, v4800, v4801, v4802, v4803, v4804, v4805, v4806, v4807, v4808, v4809, v4810, v4811, v4812, v4813, v4814, v4815, v4816, v4817, v4818, v4819, v4820, v4821, v4822, v4823, v4824, v4825, v4826, v4827, v4828, v4829, v4830, v4831, v4832, v4833, v4834, v4835, v4836, v4837, v4838, v4839, v4840, v4841, v4842, v4843, v4844, v4845, v4846, v4847, v4848, v4849, v4850, v4851, v4852, v4853, v4854, v4855, v4856, v4857, v4858, v4859, v4860, v4861, v4862, v4863, v4864, v4865, v4866, v4867, v4868, v4869, v4870, v4871, v4872, v4873, v4874, v4875, v4876, v4877, v4878, v4879, v4880, v4881, v4882, v4883, v4884, v4885, v4886, v4887, v4888, v4889, v4890, v4891, v4892, v4893, v4894, v4895, v4896, v4897, v4898, v4899, v4900, v4901, v4902, v4903, v4904, v4905, v4906, v4907, v4908, v4909, v4910, v4911, v4912, v4913, v4914, v4915, v4916, v4917, v4918, v4919, v4920, v4921, v4922, v4923, v4924, v4925, v4926, v4927, v4928, v4929, v4930, v4931, v4932, v4933, v4934, v4935, v4936, v4937, v4938, v4939, v4940, v4941, v4942, v4943, v4944, v4945, v4946, v4947, v4948, v4949, v4950, v4951, v4952, v4953, v4954, v4955, v4956, v4957, v4958, v4959, v4960, v4961, v4962, v4963, v4964, v4965, v4966, v4967, v4968, v4969, v4970, v4971, v4972, v4973, v4974, v4975, v4976, v4977, v4978, v4979, v4980, v4981, v4982, v4983, v4984, v4985, v4986, v4987, v4988, v4989, v4990, v4991, v4992, v4993, v4994, v4995, v4996, v4997, v4998, v4999, v5000, v5001, v5002, v5003, v5004, v5005, v5006, v5007, v5008, v5009, v5010, v5011, v5012, v5013, v5014, v5015, v5016, v5017, v5018, v5019, v5020, v5021, v5022, v5023, v5024, v5025, v5026, v5027, v5028, v5029, v5030, v5031, v5032, v5033, v5034, v5035, v5036, v5037, v5038, v5039, v5040, v5041, v5042, v5043, v5044, v5045, v5046, v5047, v5048, v5049, v5050, v5051, v5052, v5053, v5054, v5055, v5056, v5057, v5058, v5059, v5060, v5061, v5062, v5063, v5064, v5065, v5066, v5067, v5068, v5069, v5070, v5071, v5072, v5073, v5074, v5075, v5076, v5077, v5078, v5079, v5080, v5081, v5082, v5083, v5084, v5085, v5086, v5087, v5088, v5089, v5090, v5091, v5092, v5093, v5094, v5095, v5096, v5097, v5098, v5099, v5100, v5101, v5102, v5103, v5104, v5105, v5106, v5107, v5108, v5109, v5110, v5111, v5112, v5113, v5114, v5115, v5116, v5117, v5118, v5119, v5120, v5121, v5122, v5123, v5124, v5125, v5126, v5127, v5128, v5129, v5130, v5131, v5132, v5133, v5134, v5135, v5136, v5137, v5138, v5139, v5140, v5141, v5142, v5143, v5144, v5145, v5146, v5147, v5148, v5149, v5150, v5151, v5152, v5153, v5154, v5155, v5156, v5157, v5158, v5159, v5160, v5161, v5162, v5163, v5164, v5165, v5166, v5167, v5168, v5169, v5170, v5171, v5172, v5173, v5174, v5175, v5176, v5177, v5178, v5179, v5180, v5181, v5182, v5183, v5184, v5185, v5186, v5187, v5188, v5189, v5190, v5191, v5192, v5193, v5194, v5195, v5196, v5197, v5198, v5199, v5200, v5201, v5202, v5203, v5204, v5205, v5206, v5207, v5208, v5209, v5210, v5211, v5212, v5213, v5214, v5215, v5216, v5217, v5218, v5219, v5220, v5221, v5222, v5223, v5224, v5225, v5226, v5227, v5228, v5229, v5230, v5231, v5232, v5233, v5234, v5235, v5236, v5237, v5238, v5239, v5240, v5241, v5242, v5243, v5244, v5245, v5246, v5247, v5248, v5249, v5250, v5251, v5252, v5253, v5254, v5255, v5256, v5257, v5258, v5259, v5260, v5261, v5262, v5263, v5264, v5265, v5266, v5267, v5268, v5269, v5270, v5271, v5272, v5273, v5274, v5275, v5276, v5277, v5278, v5279, v5280, v5281, v5282, v5283, v5284, v5285, v5286, v5287, v5288, v5289, v5290, v5291, v5292, v5293, v5294, v5295, v5296, v5297, v5298, v5299, v5300, v5301, v5302, v5303, v5304, v5305, v5306, v5307, v5308, v5309, v5310, v5311, v5312, v5313, v5314, v5315, v5316, v5317, v5318, v5319, v5320, v5321, v5322, v5323, v5324, v5325, v5326, v5327, v5328, v5329, v5330, v5331, v5332, v5333, v5334, v5335, v5336, v5337, v5338, v5339, v5340, v5341, v5342, v5343, v5344, v5345, v5346, v5347, v5348, v5349, v5350, v5351, v5352, v5353, v5354, v5355, v5356, v5357, v5358, v5359, v5360, v5361, v5362, v5363, v5364, v5365, v5366, v5367, v5368, v5369, v5370, v5371, v5372, v5373, v5374, v5375, v5376, v5377, v5378, v5379, v5380, v5381, v5382, v5383, v5384, v5385, v5386, v5387, v5388, v5389, v5390, v5391, v5392, v5393, v5394, v5395, v5396, v5397, v5398, v5399, v5400, v5401, v5402, v5403, v5404, v5405, v5406, v5407, v5408, v5409, v5410, v5411, v5412, v5413, v5414, v5415, v5416, v5417, v5418, v5419, v5420, v5421, v5422, v5423, v5424, v5425, v5426, v5427, v5428, v5429, v5430, v5431, v5432, v5433, v5434, v5435, v5436, v5437, v5438, v5439, v5440, v5441, v5442, v5443, v5444, v5445, v5446, v5447, v5448, v5449, v5450, v5451, v5452, v5453, v5454, v5455, v5456, v5457, v5458, v5459, v5460, v5461, v5462, v5463, v5464, v5465, v5466, v5467, v5468, v5469, v5470, v5471, v5472, v5473, v5474, v5475, v5476, v5477, v5478, v5479, v5480, v5481, v5482, v5483, v5484, v5485, v5486, v5487, v5488, v5489, v5490, v5491, v5492, v5493, v5494, v5495, v5496, v5497, v5498, v5499, v5500, v5501, v5502, v5503, v5504, v5505, v5506, v5507, v5508, v5509, v5510, v5511, v5512, v5513, v5514, v5515, v5516, v5517, v5518, v5519, v5520, v5521, v5522, v5523, v5524, v5525, v5526, v5527, v5528, v5529, v5530, v5531, v5532, v5533, v5534, v5535, v5536, v5537, v5538, v5539, v5540, v5541, v5542, v5543, v5544, v5545, v5546, v5547, v5548, v5549, v5550, v5551, v5552, v5553, v5554, v5555, v5556, v5557, v5558, v5559, v5560, v5561, v5562, v5563, v5564, v5565, v5566, v5567, v5568, v5569, v5570, v5571, v5572, v5573, v5574, v5575, v5576, v5577, v5578, v5579, v5580, v5581, v5582, v5583, v5584, v5585, v5586, v5587, v5588, v5589, v5590, v5591, v5592, v5593, v5594, v5595, v5596, v5597, v5598, v5599, v5600, v5601, v5602, v5603, v5604, v5605, v5606, v5607, v5608, v5609, v5610, v5611, v5612, v5613, v5614, v5615, v5616, v5617, v5618, v5619, v5620, v5621, v5622, v5623, v5624, v5625, v5626, v5627, v5628, v5629, v5630, v5631, v5632, v5633, v5634, v5635, v5636, v5637, v5638, v5639, v5640, v5641, v5642, v5643, v5644, v5645, v5646, v5647, v5648, v5649, v5650, v5651, v5652, v5653, v5654, v5655, v5656, v5657, v5658, v5659, v5660, v5661, v5662, v5663, v5664, v5665, v5666, v5667, v5668, v5669, v5670, v5671, v5672, v5673, v5674, v5675, v5676, v5677, v5678, v5679, v5680, v5681, v5682, v5683, v5684, v5685, v5686, v5687, v5688, v5689, v5690, v5691, v5692, v5693, v5694, v5695, v5696, v5697, v5698, v5699, v5700, v5701, v5702, v5703, v5704, v5705, v5706, v5707, v5708, v5709, v5710, v5711, v5712, v5713, v5714, v5715, v5716, v5717, v5718, v5719, v5720, v5721, v5722, v5723, v5724, v5725, v5726, v5727, v5728, v5729, v5730, v5731, v5732, v5733, v5734, v5735, v5736, v5737, v5738, v5739, v5740, v5741, v5742, v5743, v5744, v5745, v5746, v5747, v5748, v5749, v5750, v5751, v5752, v5753, v5754, v5755, v5756, v5757, v5758, v5759, v5760, v5761, v5762, v5763, v5764, v5765, v5766, v5767, v5768, v5769, v5770, v5771, v5772, v5773, v5774, v5775, v5776, v5777, v5778, v5779, v5780, v5781, v5782, v5783, v5784, v5785, v5786, v5787, v5788, v5789, v5790, v5791, v5792, v5793, v5794, v5795, v5796, v5797, v5798, v5799, v5800, v5801, v5802, v5803, v5804, v5805, v5806, v5807, v5808, v5809, v5810, v5811, v5812, v5813, v5814, v5815, v5816, v5817, v5818, v5819, v5820, v5821, v5822, v5823, v5824, v5825, v5826, v5827, v5828, v5829, v5830, v5831, v5832, v5833, v5834, v5835, v5836, v5837, v5838, v5839, v5840, v5841, v5842, v5843, v5844, v5845, v5846, v5847, v5848, v5849, v5850, v5851, v5852, v5853, v5854, v5855, v5856, v5857, v5858, v5859, v5860, v5861, v5862, v5863, v5864, v5865, v5866, v5867, v5868, v5869, v5870, v5871, v5872, v5873, v5874, v5875, v5876, v5877, v5878, v5879, v5880, v5881, v5882, v5883, v5884, v5885, v5886, v5887, v5888, v5889, v5890, v5891, v5892, v5893, v5894, v5895, v5896, v5897, v5898, v5899, v5900, v5901, v5902, v5903, v5904, v5905, v5906, v5907, v5908, v5909, v5910, v5911, v5912, v5913, v5914, v5915, v5916, v5917, v5918, v5919, v5920, v5921, v5922, v5923, v5924, v5925, v5926, v5927, v5928, v5929, v5930, v5931, v5932, v5933, v5934, v5935, v5936, v5937, v5938, v5939, v5940, v5941, v5942, v5943, v5944, v5945, v5946, v5947, v5948, v5949, v5950, v5951, v5952, v5953, v5954, v5955, v5956, v5957, v5958, v5959, v5960, v5961, v5962, v5963, v5964, v5965, v5966, v5967, v5968, v5969, v5970, v5971, v5972, v5973, v5974, v5975, v5976, v5977, v5978, v5979, v5980, v5981, v5982, v5983, v5984, v5985, v5986, v5987, v5988, v5989, v5990, v5991, v5992, v5993, v5994, v5995, v5996, v5997, v5998, v5999, v6000, v6001, v6002, v6003, v6004, v6005, v6006, v6007, v6008, v6009, v6010, v6011, v6012, v6013, v6014, v6015, v6016, v6017, v6018, v6019, v6020, v6021, v6022, v6023, v6024, v6025, v6026, v6027, v6028, v6029, v6030, v6031, v6032, v6033, v6034, v6035, v6036, v6037, v6038, v6039, v6040, v6041, v6042, v6043, v6044, v6045, v6046, v6047, v6048, v6049, v6050, v6051, v6052, v6053, v6054, v6055, v6056, v6057, v6058, v6059, v6060, v6061, v6062, v6063, v6064, v6065, v6066, v6067, v6068, v6069, v6070, v6071, v6072, v6073, v6074, v6075, v6076, v6077, v6078, v6079, v6080, v6081, v6082, v6083, v6084, v6085, v6086, v6087, v6088, v6089, v6090, v6091, v6092, v6093, v6094, v6095, v6096, v6097, v6098, v6099, v6100, v6101, v6102, v6103, v6104, v6105, v6106, v6107, v6108, v6109, v6110, v6111, v6112, v6113, v6114, v6115, v6116, v6117, v6118, v6119, v6120, v6121, v6122, v6123, v6124, v6125, v6126, v6127, v6128, v6129, v6130, v6131, v6132, v6133, v6134, v6135, v6136, v6137, v6138, v6139, v6140, v6141, v6142, v6143, v6144, v6145, v6146, v6147, v6148, v6149, v6150, v6151, v6152, v6153, v6154, v6155, v6156, v6157, v6158, v6159, v6160, v6161, v6162, v6163, v6164, v6165, v6166, v6167, v6168, v6169, v6170, v6171, v6172, v6173, v6174, v6175, v6176, v6177, v6178, v6179, v6180, v6181, v6182, v6183, v6184, v6185, v6186, v6187, v6188, v6189, v6190, v6191, v6192, v6193, v6194, v6195, v6196, v6197, v6198, v6199, v6200, v6201, v6202, v6203, v6204, v6205, v6206, v6207, v6208, v6209, v6210, v6211, v6212, v6213, v6214, v6215, v6216, v6217, v6218, v6219, v6220, v6221, v6222, v6223, v6224, v6225, v6226, v6227, v6228, v6229, v6230, v6231, v6232, v6233, v6234, v6235, v6236, v6237, v6238, v6239, v6240, v6241, v6242, v6243, v6244, v6245, v6246, v6247, v6248, v6249, v6250, v6251, v6252, v6253, v6254, v6255, v6256, v6257, v6258, v6259, v6260, v6261, v6262, v6263, v6264, v6265, v6266, v6267, v6268, v6269, v6270, v6271, v6272, v6273, v6274, v6275, v6276, v6277, v6278, v6279, v6280, v6281, v6282, v6283, v6284, v6285, v6286, v6287, v6288, v6289, v6290, v6291, v6292, v6293, v6294, v6295, v6296, v6297, v6298, v6299, v6300, v6301, v6302, v6303, v6304, v6305, v6306, v6307, v6308, v6309, v6310, v6311, v6312, v6313, v6314, v6315, v6316, v6317, v6318, v6319, v6320, v6321, v6322, v6323, v6324, v6325, v6326, v6327, v6328, v6329, v6330, v6331, v6332, v6333, v6334, v6335, v6336, v6337, v6338, v6339, v6340, v6341, v6342, v6343, v6344, v6345, v6346, v6347, v6348, v6349, v6350, v6351, v6352, v6353, v6354, v6355, v6356, v6357, v6358, v6359, v6360, v6361, v6362, v6363, v6364, v6365, v6366, v6367, v6368, v6369, v6370, v6371, v6372, v6373, v6374, v6375, v6376, v6377, v6378, v6379, v6380, v6381, v6382, v6383, v6384, v6385, v6386, v6387, v6388, v6389, v6390, v6391, v6392, v6393, v6394, v6395, v6396, v6397, v6398, v6399, v6400, v6401, v6402, v6403, v6404, v6405, v6406, v6407, v6408, v6409, v6410, v6411, v6412, v6413, v6414, v6415, v6416, v6417, v6418, v6419, v6420, v6421, v6422, v6423, v6424, v6425, v6426, v6427, v6428, v6429, v6430, v6431, v6432, v6433, v6434, v6435, v6436, v6437, v6438, v6439, v6440, v6441, v6442, v6443, v6444, v6445, v6446, v6447, v6448, v6449, v6450, v6451, v6452, v6453, v6454, v6455, v6456, v6457, v6458, v6459, v6460, v6461, v6462, v6463, v6464, v6465, v6466, v6467, v6468, v6469, v6470, v6471, v6472, v6473, v6474, v6475, v6476, v6477, v6478, v6479, v6480, v6481, v6482, v6483, v6484, v6485, v6486, v6487, v6488, v6489, v6490, v6491, v6492, v6493, v6494, v6495, v6496, v6497, v6498, v6499, v6500, v6501, v6502, v6503, v6504, v6505, v6506, v6507, v6508, v6509, v6510, v6511, v6512, v6513, v6514, v6515, v6516, v6517, v6518, v6519, v6520, v6521, v6522, v6523, v6524, v6525, v6526, v6527, v6528, v6529, v6530, v6531, v6532, v6533, v6534, v6535, v6536, v6537, v6538, v6539, v6540, v6541, v6542, v6543, v6544, v6545, v6546, v6547, v6548, v6549, v6550, v6551, v6552, v6553, v6554, v6555, v6556, v6557, v6558, v6559, v6560, v6561, v6562, v6563, v6564, v6565, v6566, v6567, v6568, v6569, v6570, v6571, v6572, v6573, v6574, v6575, v6576, v6577, v6578, v6579, v6580, v6581, v6582, v6583, v6584, v6585, v6586, v6587, v6588, v6589, v6590, v6591, v6592, v6593, v6594, v6595, v6596, v6597, v6598, v6599, v6600, v6601, v6602, v6603, v6604, v6605, v6606, v6607, v6608, v6609, v6610, v6611, v6612, v6613, v6614, v6615, v6616, v6617, v6618, v6619, v6620, v6621, v6622, v6623, v6624, v6625, v6626, v6627, v6628, v6629, v6630, v6631, v6632, v6633, v6634, v6635, v6636, v6637, v6638, v6639, v6640, v6641, v6642, v6643, v6644, v6645, v6646, v6647, v6648, v6649, v6650, v6651, v6652, v6653, v6654, v6655, v6656, v6657, v6658, v6659, v6660, v6661, v6662, v6663, v6664, v6665, v6666, v6667, v6668, v6669, v6670, v6671, v6672, v6673, v6674, v6675, v6676, v6677, v6678, v6679, v6680, v6681, v6682, v6683, v6684, v6685, v6686, v6687, v6688, v6689, v6690, v6691, v6692, v6693, v6694, v6695, v6696, v6697, v6698, v6699, v6700, v6701, v6702, v6703, v6704, v6705, v6706, v6707, v6708, v6709, v6710, v6711, v6712, v6713, v6714, v6715, v6716, v6717, v6718, v6719, v6720, v6721, v6722, v6723, v6724, v6725, v6726, v6727, v6728, v6729, v6730, v6731, v6732, v6733, v6734, v6735, v6736, v6737, v6738, v6739, v6740, v6741, v6742, v6743, v6744, v6745, v6746, v6747, v6748, v6749, v6750, v6751, v6752, v6753, v6754, v6755, v6756, v6757, v6758, v6759, v6760, v6761, v6762, v6763, v6764, v6765, v6766, v6767, v6768, v6769, v6770, v6771, v6772, v6773, v6774, v6775, v6776, v6777, v6778, v6779, v6780, v6781, v6782, v6783, v6784, v6785, v6786, v6787, v6788, v6789, v6790, v6791, v6792, v6793, v6794, v6795, v6796, v6797, v6798, v6799, v6800, v6801, v6802, v6803, v6804, v6805, v6806, v6807, v6808, v6809, v6810, v6811, v6812, v6813, v6814, v6815, v6816, v6817, v6818, v6819, v6820, v6821, v6822, v6823, v6824, v6825, v6826, v6827, v6828, v6829, v6830, v6831, v6832, v6833, v6834, v6835, v6836, v6837, v6838, v6839, v6840, v6841, v6842, v6843, v6844, v6845, v6846, v6847, v6848, v6849, v6850, v6851, v6852, v6853, v6854, v6855, v6856, v6857, v6858, v6859, v6860, v6861, v6862, v6863, v6864, v6865, v6866, v6867, v6868, v6869, v6870, v6871, v6872, v6873, v6874, v6875, v6876, v6877, v6878, v6879, v6880, v6881, v6882, v6883, v6884, v6885, v6886, v6887, v6888, v6889, v6890, v6891, v6892, v6893, v6894, v6895, v6896, v6897, v6898, v6899, v6900, v6901, v6902, v6903, v6904, v6905, v6906, v6907, v6908, v6909, v6910, v6911, v6912, v6913, v6914, v6915, v6916, v6917, v6918, v6919, v6920, v6921, v6922, v6923, v6924, v6925, v6926, v6927, v6928, v6929, v6930, v6931, v6932, v6933, v6934, v6935, v6936, v6937, v6938, v6939, v6940, v6941, v6942, v6943, v6944, v6945, v6946, v6947, v6948, v6949, v6950, v6951, v6952, v6953, v6954, v6955, v6956, v6957, v6958, v6959, v6960, v6961, v6962, v6963, v6964, v6965, v6966, v6967, v6968, v6969, v6970, v6971, v6972, v6973, v6974, v6975, v6976, v6977, v6978, v6979, v6980, v6981, v6982, v6983, v6984, v6985, v6986, v6987, v6988, v6989, v6990, v6991, v6992, v6993, v6994, v6995, v6996, v6997, v6998, v6999, v7000, v7001, v7002, v7003, v7004, v7005, v7006, v7007, v7008, v7009, v7010, v7011, v7012, v7013, v7014, v7015, v7016, v7017, v7018, v7019, v7020, v7021, v7022, v7023, v7024, v7025, v7026, v7027, v7028, v7029, v7030, v7031, v7032, v7033, v7034, v7035, v7036, v7037, v7038, v7039, v7040, v7041, v7042, v7043, v7044, v7045, v7046, v7047, v7048, v7049, v7050, v7051, v7052, v7053, v7054, v7055, v7056, v7057, v7058, v7059, v7060, v7061, v7062, v7063, v7064, v7065, v7066, v7067, v7068, v7069, v7070, v7071, v7072, v7073, v7074, v7075, v7076, v7077, v7078, v7079, v7080, v7081, v7082, v7083, v7084, v7085, v7086, v7087, v7088, v7089, v7090, v7091, v7092, v7093, v7094, v7095, v7096, v7097, v7098, v7099, v7100, v7101, v7102, v7103, v7104, v7105, v7106, v7107, v7108, v7109, v7110, v7111, v7112, v7113, v7114, v7115, v7116, v7117, v7118, v7119, v7120, v7121, v7122, v7123, v7124, v7125, v7126, v7127, v7128, v7129, v7130, v7131, v7132, v7133, v7134, v7135, v7136, v7137, v7138, v7139, v7140, v7141, v7142, v7143, v7144, v7145, v7146, v7147, v7148, v7149, v7150, v7151, v7152, v7153, v7154, v7155, v7156, v7157, v7158, v7159, v7160, v7161, v7162, v7163, v7164, v7165, v7166, v7167, v7168, v7169, v7170, v7171, v7172, v7173, v7174, v7175, v7176, v7177, v7178, v7179, v7180, v7181, v7182, v7183, v7184, v7185, v7186, v7187, v7188, v7189, v7190, v7191, v7192, v7193, v7194, v7195, v7196, v7197, v7198, v7199, v7200, v7201, v7202, v7203, v7204, v7205, v7206, v7207, v7208, v7209, v7210, v7211, v7212, v7213, v7214, v7215, v7216, v7217, v7218, v7219, v7220, v7221, v7222, v7223, v7224, v7225, v7226, v7227, v7228, v7229, v7230, v7231, v7232, v7233, v7234, v7235, v7236, v7237, v7238, v7239, v7240, v7241, v7242, v7243, v7244, v7245, v7246, v7247, v7248, v7249, v7250, v7251, v7252, v7253, v7254, v7255, v7256, v7257, v7258, v7259, v7260, v7261, v7262, v7263, v7264, v7265, v7266, v7267, v7268, v7269, v7270, v7271, v7272, v7273, v7274, v7275, v7276, v7277, v7278, v7279, v7280, v7281, v7282, v7283, v7284, v7285, v7286, v7287, v7288, v7289, v7290, v7291, v7292, v7293, v7294, v7295, v7296, v7297, v7298, v7299, v7300, v7301, v7302, v7303, v7304, v7305, v7306, v7307, v7308, v7309, v7310, v7311, v7312, v7313, v7314, v7315, v7316, v7317, v7318, v7319, v7320, v7321, v7322, v7323, v7324, v7325, v7326, v7327, v7328, v7329, v7330, v7331, v7332, v7333, v7334, v7335, v7336, v7337, v7338, v7339, v7340, v7341, v7342, v7343, v7344, v7345, v7346, v7347, v7348, v7349, v7350, v7351, v7352, v7353, v7354, v7355, v7356, v7357, v7358, v7359, v7360, v7361, v7362, v7363, v7364, v7365, v7366, v7367, v7368, v7369, v7370, v7371, v7372, v7373, v7374, v7375, v7376, v7377, v7378, v7379, v7380, v7381, v7382, v7383, v7384, v7385, v7386, v7387, v7388, v7389, v7390, v7391, v7392, v7393, v7394, v7395, v7396, v7397, v7398, v7399, v7400, v7401, v7402, v7403, v7404, v7405, v7406, v7407, v7408, v7409, v7410, v7411, v7412, v7413, v7414, v7415, v7416, v7417, v7418, v7419, v7420, v7421, v7422, v7423, v7424, v7425, v7426, v7427, v7428, v7429, v7430, v7431, v7432, v7433, v7434, v7435, v7436, v7437, v7438, v7439, v7440, v7441, v7442, v7443, v7444, v7445, v7446, v7447, v7448, v7449, v7450, v7451, v7452, v7453, v7454, v7455, v7456, v7457, v7458, v7459, v7460, v7461, v7462, v7463, v7464, v7465, v7466, v7467, v7468, v7469, v7470, v7471, v7472, v7473, v7474, v7475, v7476, v7477, v7478, v7479, v7480, v7481, v7482, v7483, v7484, v7485, v7486, v7487, v7488, v7489, v7490, v7491, v7492, v7493, v7494, v7495, v7496, v7497, v7498, v7499, v7500, v7501, v7502, v7503, v7504, v7505, v7506, v7507, v7508, v7509, v7510, v7511, v7512, v7513, v7514, v7515, v7516, v7517, v7518, v7519, v7520, v7521, v7522, v7523, v7524, v7525, v7526, v7527, v7528, v7529, v7530, v7531, v7532, v7533, v7534, v7535, v7536, v7537, v7538, v7539, v7540, v7541, v7542, v7543, v7544, v7545, v7546, v7547, v7548, v7549, v7550, v7551, v7552, v7553, v7554, v7555, v7556, v7557, v7558, v7559, v7560, v7561, v7562, v7563, v7564, v7565, v7566, v7567, v7568, v7569, v7570, v7571, v7572, v7573, v7574, v7575, v7576, v7577, v7578, v7579, v7580, v7581, v7582, v7583, v7584, v7585, v7586, v7587, v7588, v7589, v7590, v7591, v7592, v7593, v7594, v7595, v7596, v7597, v7598, v7599, v7600, v7601, v7602, v7603, v7604, v7605, v7606, v7607, v7608, v7609, v7610, v7611, v7612, v7613, v7614, v7615, v7616, v7617, v7618, v7619, v7620, v7621, v7622, v7623, v7624, v7625, v7626, v7627, v7628, v7629, v7630, v7631, v7632, v7633, v7634, v7635, v7636, v7637, v7638, v7639, v7640, v7641, v7642, v7643, v7644, v7645, v7646, v7647, v7648, v7649, v7650, v7651, v7652, v7653, v7654, v7655, v7656, v7657, v7658, v7659, v7660, v7661, v7662, v7663, v7664, v7665, v7666, v7667, v7668, v7669, v7670, v7671, v7672, v7673, v7674, v7675, v7676, v7677, v7678, v7679, v7680, v7681, v7682, v7683, v7684, v7685, v7686, v7687, v7688, v7689, v7690, v7691, v7692, v7693, v7694, v7695, v7696, v7697, v7698, v7699, v7700, v7701, v7702, v7703, v7704, v7705, v7706, v7707, v7708, v7709, v7710, v7711, v7712, v7713, v7714, v7715, v7716, v7717, v7718, v7719, v7720, v7721, v7722, v7723, v7724, v7725, v7726, v7727, v7728, v7729, v7730, v7731, v7732, v7733, v7734, v7735, v7736, v7737, v7738, v7739, v7740, v7741, v7742, v7743, v7744, v7745, v7746, v7747, v7748, v7749, v7750, v7751, v7752, v7753, v7754, v7755, v7756, v7757, v7758, v7759, v7760, v7761, v7762, v7763, v7764, v7765, v7766, v7767, v7768, v7769, v7770, v7771, v7772, v7773, v7774, v7775, v7776, v7777, v7778, v7779, v7780, v7781, v7782, v7783, v7784, v7785, v7786, v7787, v7788, v7789, v7790, v7791, v7792, v7793, v7794, v7795, v7796, v7797, v7798, v7799, v7800, v7801, v7802, v7803, v7804, v7805, v7806, v7807, v7808, v7809, v7810, v7811, v7812, v7813, v7814, v7815, v7816, v7817, v7818, v7819, v7820, v7821, v7822, v7823, v7824, v7825, v7826, v7827, v7828, v7829, v7830, v7831, v7832, v7833, v7834, v7835, v7836, v7837, v7838, v7839, v7840, v7841, v7842, v7843, v7844, v7845, v7846, v7847, v7848, v7849, v7850, v7851, v7852, v7853, v7854, v7855, v7856, v7857, v7858, v7859, v7860, v7861, v7862, v7863, v7864, v7865, v7866, v7867, v7868, v7869, v7870, v7871, v7872, v7873, v7874, v7875, v7876, v7877, v7878, v7879, v7880, v7881, v7882, v7883, v7884, v7885, v7886, v7887, v7888, v7889, v7890, v7891, v7892, v7893, v7894, v7895, v7896, v7897, v7898, v7899, v7900, v7901, v7902, v7903, v7904, v7905, v7906, v7907, v7908, v7909, v7910, v7911, v7912, v7913, v7914, v7915, v7916, v7917, v7918, v7919, v7920, v7921, v7922, v7923, v7924, v7925, v7926, v7927, v7928, v7929, v7930, v7931, v7932, v7933, v7934, v7935, v7936, v7937, v7938, v7939, v7940, v7941, v7942, v7943, v7944, v7945, v7946, v7947, v7948, v7949, v7950, v7951, v7952, v7953, v7954, v7955, v7956, v7957, v7958, v7959, v7960, v7961, v7962, v7963, v7964, v7965, v7966, v7967, v7968, v7969, v7970, v7971, v7972, v7973, v7974, v7975, v7976, v7977, v7978, v7979, v7980, v7981, v7982, v7983, v7984, v7985, v7986, v7987, v7988, v7989, v7990, v7991, v7992, v7993, v7994, v7995, v7996, v7997, v7998, v7999, v8000, v8001, v8002, v8003, v8004, v8005, v8006, v8007, v8008, v8009, v8010, v8011, v8012, v8013, v8014, v8015, v8016, v8017, v8018, v8019, v8020, v8021, v8022, v8023, v8024, v8025, v8026, v8027, v8028, v8029, v8030, v8031, v8032, v8033, v8034, v8035, v8036, v8037, v8038, v8039, v8040, v8041, v8042, v8043, v8044, v8045, v8046, v8047, v8048, v8049, v8050, v8051, v8052, v8053, v8054, v8055, v8056, v8057, v8058, v8059, v8060, v8061, v8062, v8063, v8064, v8065, v8066, v8067, v8068, v8069, v8070, v8071, v8072, v8073, v8074, v8075, v8076, v8077, v8078, v8079, v8080, v8081, v8082, v8083, v8084, v8085, v8086, v8087, v8088, v8089, v8090, v8091, v8092, v8093, v8094, v8095, v8096, v8097, v8098, v8099, v8100, v8101, v8102, v8103, v8104, v8105, v8106, v8107, v8108, v8109, v8110, v8111, v8112, v8113, v8114, v8115, v8116, v8117, v8118, v8119, v8120, v8121, v8122, v8123, v8124, v8125, v8126, v8127, v8128, v8129, v8130, v8131, v8132, v8133, v8134, v8135, v8136, v8137, v8138, v8139, v8140, v8141, v8142, 
w0, w1, w2, w3, w4, w5, w6, w7, w8, w9, w10, w11, w12, w13, w14, w15, w16, w17, w18, w19, w20, w21, w22, w23, w24, w25, w26, w27, w28, w29, w30, w31, w32, w33, w34, w35, w36, w37, w38, w39, w40, w41, w42, w43, w44, w45, w46, w47, w48, w49, w50, w51, w52, w53, w54, w55, w56, w57, w58, w59, w60, w61, w62, w63, w64, w65, w66, w67, w68, w69, w70, w71, w72, w73, w74, w75, w76, w77, w78, w79, w80, w81, w82, w83, w84, w85, w86, w87, w88, w89, w90, w91, w92, w93, w94, w95, w96, w97, w98, w99, w100, w101, w102, w103, w104, w105, w106, w107, w108, w109, w110, w111, w112, w113, w114, w115, w116, w117, w118, w119, w120, w121, w122, w123, w124, w125, w126, w127, w128, w129, w130, w131, w132, w133, w134, w135, w136, w137, w138, w139, w140, w141, w142, w143, w144, w145, w146, w147, w148, w149, w150, w151, w152, w153, w154, w155, w156, w157, w158, w159, w160, w161, w162, w163, w164, w165, w166, w167, w168, w169, w170, w171, w172, w173, w174, w175, w176, w177, w178, w179, w180, w181, w182, w183, w184, w185, w186, w187, w188, w189, w190, w191, w192, w193, w194, w195, w196, w197, w198, w199, w200, w201, w202, w203, w204, w205, w206, w207, w208, w209, w210, w211, w212, w213, w214, w215, w216, w217, w218, w219, w220, w221, w222, w223, w224, w225, w226, w227, w228, w229, w230, w231, w232, w233, w234, w235, w236, w237, w238, w239, w240, w241, w242, w243, w244, w245, w246, w247, w248, w249, w250, w251, w252, w253, w254, w255, w256, w257, w258, w259, w260, w261, w262, w263, w264, w265, w266, w267, w268, w269, w270, w271, w272, w273, w274, w275, w276, w277, w278, w279, w280, w281, w282, w283, w284, w285, w286, w287, w288, w289, w290, w291, w292, w293, w294, w295, w296, w297, w298, w299, w300, w301, w302, w303, w304, w305, w306, w307, w308, w309, w310, w311, w312, w313, w314, w315, w316, w317, w318, w319, w320, w321, w322, w323, w324, w325, w326, w327, w328, w329, w330, w331, w332, w333, w334, w335, w336, w337, w338, w339, w340, w341, w342, w343, w344, w345, w346, w347, w348, w349, w350, w351, w352, w353, w354, w355, w356, w357, w358, w359, w360, w361, w362, w363, w364, w365, w366, w367, w368, w369, w370, w371, w372, w373, w374, w375, w376, w377, w378, w379, w380, w381, w382, w383, w384, w385, w386, w387, w388, w389, w390, w391, w392, w393, w394, w395, w396, w397, w398, w399, w400, w401, w402, w403, w404, w405, w406, w407, w408, w409, w410, w411, w412, w413, w414, w415, w416, w417, w418, w419, w420, w421, w422, w423, w424, w425, w426, w427, w428, w429, w430, w431, w432, w433, w434, w435, w436, w437, w438, w439, w440, w441, w442, w443, w444, w445, w446, w447, w448, w449, w450, w451, w452, w453, w454, w455, w456, w457, w458, w459, w460, w461, w462, w463, w464, w465, w466, w467, w468, w469, w470, w471, w472, w473, w474, w475, w476, w477, w478, w479, w480, w481, w482, w483, w484, w485, w486, w487, w488, w489, w490, w491, w492, w493, w494, w495, w496, w497, w498, w499, w500, w501, w502, w503, w504, w505, w506, w507, w508, w509, w510, w511, w512, w513, w514, w515, w516, w517, w518, w519, w520, w521, w522, w523, w524, w525, w526, w527, w528, w529, w530, w531, w532, w533, w534, w535, w536, w537, w538, w539, w540, w541, w542, w543, w544, w545, w546, w547, w548, w549, w550, w551, w552, w553, w554, w555, w556, w557, w558, w559, w560, w561, w562, w563, w564, w565, w566, w567, w568, w569, w570, w571, w572, w573, w574, w575, w576, w577, w578, w579, w580, w581, w582, w583, w584, w585, w586, w587, w588, w589, w590, w591, w592, w593, w594, w595, w596, w597, w598, w599, w600, w601, w602, w603, w604, w605, w606, w607, w608, w609, w610, w611, w612, w613, w614, w615, w616, w617, w618, w619, w620, w621, w622, w623, w624, w625, w626, w627, w628, w629, w630, w631, w632, w633, w634, w635, w636, w637, w638, w639, w640, w641, w642, w643, w644, w645, w646, w647, w648, w649, w650, w651, w652, w653, w654, w655, w656, w657, w658, w659, w660, w661, w662, w663, w664, w665, w666, w667, w668, w669, w670, w671, w672, w673, w674, w675, w676, w677, w678, w679, w680, w681, w682, w683, w684, w685, w686, w687, w688, w689, w690, w691, w692, w693, w694, w695, w696, w697, w698, w699, w700, w701, w702, w703, w704, w705, w706, w707, w708, w709, w710, w711, w712, w713, w714, w715, w716, w717, w718, w719, w720, w721, w722, w723, w724, w725, w726, w727, w728, w729, w730, w731, w732, w733, w734, w735, w736, w737, w738, w739, w740, w741, w742, w743, w744, w745, w746, w747, w748, w749, w750, w751, w752, w753, w754, w755, w756, w757, w758, w759, w760, w761, w762, w763, w764, w765, w766, w767, w768, w769, w770, w771, w772, w773, w774, w775, w776, w777, w778, w779, w780, w781, w782, w783, w784, w785, w786, w787, w788, w789, w790, w791, w792, w793, w794, w795, w796, w797, w798, w799, w800, w801, w802, w803, w804, w805, w806, w807, w808, w809, w810, w811, w812, w813, w814, w815, w816, w817, w818, w819, w820, w821, w822, w823, w824, w825, w826, w827, w828, w829, w830, w831, w832, w833, w834, w835, w836, w837, w838, w839, w840, w841, w842, w843, w844, w845, w846, w847, w848, w849, w850, w851, w852, w853, w854, w855, w856, w857, w858, w859, w860, w861, w862, w863, w864, w865, w866, w867, w868, w869, w870, w871, w872, w873, w874, w875, w876, w877, w878, w879, w880, w881, w882, w883, w884, w885, w886, w887, w888, w889, w890, w891, w892, w893, w894, w895, w896, w897, w898, w899, w900, w901, w902, w903, w904, w905, w906, w907, w908, w909, w910, w911, w912, w913, w914, w915, w916, w917, w918, w919, w920, w921, w922, w923, w924, w925, w926, w927, w928, w929, w930, w931, w932, w933, w934, w935, w936, w937, w938, w939, w940, w941, w942, w943, w944, w945, w946, w947, w948, w949, w950, w951, w952, w953, w954, w955, w956, w957, w958, w959, w960, w961, w962, w963, w964, w965, w966, w967, w968, w969, w970, w971, w972, w973, w974, w975, w976, w977, w978, w979, w980, w981, w982, w983, w984, w985, w986, w987, w988, w989, w990, w991, w992, w993, w994, w995, w996, w997, w998, w999, w1000, w1001, w1002, w1003, w1004, w1005, w1006, w1007, w1008, w1009, w1010, w1011, w1012, w1013, w1014, w1015, w1016, w1017, w1018, w1019, w1020, w1021, w1022, w1023, w1024, w1025, w1026, w1027, w1028, w1029, w1030, w1031, w1032, w1033, w1034, w1035, w1036, w1037, w1038, w1039, w1040, w1041, w1042, w1043, w1044, w1045, w1046, w1047, w1048, w1049, w1050, w1051, w1052, w1053, w1054, w1055, w1056, w1057, w1058, w1059, w1060, w1061, w1062, w1063, w1064, w1065, w1066, w1067, w1068, w1069, w1070, w1071, w1072, w1073, w1074, w1075, w1076, w1077, w1078, w1079, w1080, w1081, w1082, w1083, w1084, w1085, w1086, w1087, w1088, w1089, w1090, w1091, w1092, w1093, w1094, w1095, w1096, w1097, w1098, w1099, w1100, w1101, w1102, w1103, w1104, w1105, w1106, w1107, w1108, w1109, w1110, w1111, w1112, w1113, w1114, w1115, w1116, w1117, w1118, w1119, w1120, w1121, w1122, w1123, w1124, w1125, w1126, w1127, w1128, w1129, w1130, w1131, w1132, w1133, w1134, w1135, w1136, w1137, w1138, w1139, w1140, w1141, w1142, w1143, w1144, w1145, w1146, w1147, w1148, w1149, w1150, w1151, w1152, w1153, w1154, w1155, w1156, w1157, w1158, w1159, w1160, w1161, w1162, w1163, w1164, w1165, w1166, w1167, w1168, w1169, w1170, w1171, w1172, w1173, w1174, w1175, w1176, w1177, w1178, w1179, w1180, w1181, w1182, w1183, w1184, w1185, w1186, w1187, w1188, w1189, w1190, w1191, w1192, w1193, w1194, w1195, w1196, w1197, w1198, w1199, w1200, w1201, w1202, w1203, w1204, w1205, w1206, w1207, w1208, w1209, w1210, w1211, w1212, w1213, w1214, w1215, w1216, w1217, w1218, w1219, w1220, w1221, w1222, w1223, w1224, w1225, w1226, w1227, w1228, w1229, w1230, w1231, w1232, w1233, w1234, w1235, w1236, w1237, w1238, w1239, w1240, w1241, w1242, w1243, w1244, w1245, w1246, w1247, w1248, w1249, w1250, w1251, w1252, w1253, w1254, w1255, w1256, w1257, w1258, w1259, w1260, w1261, w1262, w1263, w1264, w1265, w1266, w1267, w1268, w1269, w1270, w1271, w1272, w1273, w1274, w1275, w1276, w1277, w1278, w1279, w1280, w1281, w1282, w1283, w1284, w1285, w1286, w1287, w1288, w1289, w1290, w1291, w1292, w1293, w1294, w1295, w1296, w1297, w1298, w1299, w1300, w1301, w1302, w1303, w1304, w1305, w1306, w1307, w1308, w1309, w1310, w1311, w1312, w1313, w1314, w1315, w1316, w1317, w1318, w1319, w1320, w1321, w1322, w1323, w1324, w1325, w1326, w1327, w1328, w1329, w1330, w1331, w1332, w1333, w1334, w1335, w1336, w1337, w1338, w1339, w1340, w1341, w1342, w1343, w1344, w1345, w1346, w1347, w1348, w1349, w1350, w1351, w1352, w1353, w1354, w1355, w1356, w1357, w1358, w1359, w1360, w1361, w1362, w1363, w1364, w1365, w1366, w1367, w1368, w1369, w1370, w1371, w1372, w1373, w1374, w1375, w1376, w1377, w1378, w1379, w1380, w1381, w1382, w1383, w1384, w1385, w1386, w1387, w1388, w1389, w1390, w1391, w1392, w1393, w1394, w1395, w1396, w1397, w1398, w1399, w1400, w1401, w1402, w1403, w1404, w1405, w1406, w1407, w1408, w1409, w1410, w1411, w1412, w1413, w1414, w1415, w1416, w1417, w1418, w1419, w1420, w1421, w1422, w1423, w1424, w1425, w1426, w1427, w1428, w1429, w1430, w1431, w1432, w1433, w1434, w1435, w1436, w1437, w1438, w1439, w1440, w1441, w1442, w1443, w1444, w1445, w1446, w1447, w1448, w1449, w1450, w1451, w1452, w1453, w1454, w1455, w1456, w1457, w1458, w1459, w1460, w1461, w1462, w1463, w1464, w1465, w1466, w1467, w1468, w1469, w1470, w1471, w1472, w1473, w1474, w1475, w1476, w1477, w1478, w1479, w1480, w1481, w1482, w1483, w1484, w1485, w1486, w1487, w1488, w1489, w1490, w1491, w1492, w1493, w1494, w1495, w1496, w1497, w1498, w1499, w1500, w1501, w1502, w1503, w1504, w1505, w1506, w1507, w1508, w1509, w1510, w1511, w1512, w1513, w1514, w1515, w1516, w1517, w1518, w1519, w1520, w1521, w1522, w1523, w1524, w1525, w1526, w1527, w1528, w1529, w1530, w1531, w1532, w1533, w1534, w1535, w1536, w1537, w1538, w1539, w1540, w1541, w1542, w1543, w1544, w1545, w1546, w1547, w1548, w1549, w1550, w1551, w1552, w1553, w1554, w1555, w1556, w1557, w1558, w1559, w1560, w1561, w1562, w1563, w1564, w1565, w1566, w1567, w1568, w1569, w1570, w1571, w1572, w1573, w1574, w1575, w1576, w1577, w1578, w1579, w1580, w1581, w1582, w1583, w1584, w1585, w1586, w1587, w1588, w1589, w1590, w1591, w1592, w1593, w1594, w1595, w1596, w1597, w1598, w1599, w1600, w1601, w1602, w1603, w1604, w1605, w1606, w1607, w1608, w1609, w1610, w1611, w1612, w1613, w1614, w1615, w1616, w1617, w1618, w1619, w1620, w1621, w1622, w1623, w1624, w1625, w1626, w1627, w1628, w1629, w1630, w1631, w1632, w1633, w1634, w1635, w1636, w1637, w1638, w1639, w1640, w1641, w1642, w1643, w1644, w1645, w1646, w1647, w1648, w1649, w1650, w1651, w1652, w1653, w1654, w1655, w1656, w1657, w1658, w1659, w1660, w1661, w1662, w1663, w1664, w1665, w1666, w1667, w1668, w1669, w1670, w1671, w1672, w1673, w1674, w1675, w1676, w1677, w1678, w1679, w1680, w1681, w1682, w1683, w1684, w1685, w1686, w1687, w1688, w1689, w1690, w1691, w1692, w1693, w1694, w1695, w1696, w1697, w1698, w1699, w1700, w1701, w1702, w1703, w1704, w1705, w1706, w1707, w1708, w1709, w1710, w1711, w1712, w1713, w1714, w1715, w1716, w1717, w1718, w1719, w1720, w1721, w1722, w1723, w1724, w1725, w1726, w1727, w1728, w1729, w1730, w1731, w1732, w1733, w1734, w1735, w1736, w1737, w1738, w1739, w1740, w1741, w1742, w1743, w1744, w1745, w1746, w1747, w1748, w1749, w1750, w1751, w1752, w1753, w1754, w1755, w1756, w1757, w1758, w1759, w1760, w1761, w1762, w1763, w1764, w1765, w1766, w1767, w1768, w1769, w1770, w1771, w1772, w1773, w1774, w1775, w1776, w1777, w1778, w1779, w1780, w1781, w1782, w1783, w1784, w1785, w1786, w1787, w1788, w1789, w1790, w1791, w1792, w1793, w1794, w1795, w1796, w1797, w1798, w1799, w1800, w1801, w1802, w1803, w1804, w1805, w1806, w1807, w1808, w1809, w1810, w1811, w1812, w1813, w1814, w1815, w1816, w1817, w1818, w1819, w1820, w1821, w1822, w1823, w1824, w1825, w1826, w1827, w1828, w1829, w1830, w1831, w1832, w1833, w1834, w1835, w1836, w1837, w1838, w1839, w1840, w1841, w1842, w1843, w1844, w1845, w1846, w1847, w1848, w1849, w1850, w1851, w1852, w1853, w1854, w1855, w1856, w1857, w1858, w1859, w1860, w1861, w1862, w1863, w1864, w1865, w1866, w1867, w1868, w1869, w1870, w1871, w1872, w1873, w1874, w1875, w1876, w1877, w1878, w1879, w1880, w1881, w1882, w1883, w1884, w1885, w1886, w1887, w1888, w1889, w1890, w1891, w1892, w1893, w1894, w1895, w1896, w1897, w1898, w1899, w1900, w1901, w1902, w1903, w1904, w1905, w1906, w1907, w1908, w1909, w1910, w1911, w1912, w1913, w1914, w1915, w1916, w1917, w1918, w1919, w1920, w1921, w1922, w1923, w1924, w1925, w1926, w1927, w1928, w1929, w1930, w1931, w1932, w1933, w1934, w1935, w1936, w1937, w1938, w1939, w1940, w1941, w1942, w1943, w1944, w1945, w1946, w1947, w1948, w1949, w1950, w1951, w1952, w1953, w1954, w1955, w1956, w1957, w1958, w1959, w1960, w1961, w1962, w1963, w1964, w1965, w1966, w1967, w1968, w1969, w1970, w1971, w1972, w1973, w1974, w1975, w1976, w1977, w1978, w1979, w1980, w1981, w1982, w1983, w1984, w1985, w1986, w1987, w1988, w1989, w1990, w1991, w1992, w1993, w1994, w1995, w1996, w1997, w1998, w1999, w2000, w2001, w2002, w2003, w2004, w2005, w2006, w2007, w2008, w2009, w2010, w2011, w2012, w2013, w2014, w2015, w2016, w2017, w2018, w2019, w2020, w2021, w2022, w2023, w2024, w2025, w2026, w2027, w2028, w2029, w2030, w2031, w2032, w2033, w2034, w2035, w2036, w2037, w2038, w2039, w2040, w2041, w2042, w2043, w2044, w2045, w2046, w2047, w2048, w2049, w2050, w2051, w2052, w2053, w2054, w2055, w2056, w2057, w2058, w2059, w2060, w2061, w2062, w2063, w2064, w2065, w2066, w2067, w2068, w2069, w2070, w2071, w2072, w2073, w2074, w2075, w2076, w2077, w2078, w2079, w2080, w2081, w2082, w2083, w2084, w2085, w2086, w2087, w2088, w2089, w2090, w2091, w2092, w2093, w2094, w2095, w2096, w2097, w2098, w2099, w2100, w2101, w2102, w2103, w2104, w2105, w2106, w2107, w2108, w2109, w2110, w2111, w2112, w2113, w2114, w2115, w2116, w2117, w2118, w2119, w2120, w2121, w2122, w2123, w2124, w2125, w2126, w2127, w2128, w2129, w2130, w2131, w2132, w2133, w2134, w2135, w2136, w2137, w2138, w2139, w2140, w2141, w2142, w2143, w2144, w2145, w2146, w2147, w2148, w2149, w2150, w2151, w2152, w2153, w2154, w2155, w2156, w2157, w2158, w2159, w2160, w2161, w2162, w2163, w2164, w2165, w2166, w2167, w2168, w2169, w2170, w2171, w2172, w2173, w2174, w2175, w2176, w2177, w2178, w2179, w2180, w2181, w2182, w2183, w2184, w2185, w2186, w2187, w2188, w2189, w2190, w2191, w2192, w2193, w2194, w2195, w2196, w2197, w2198, w2199, w2200, w2201, w2202, w2203, w2204, w2205, w2206, w2207, w2208, w2209, w2210, w2211, w2212, w2213, w2214, w2215, w2216, w2217, w2218, w2219, w2220, w2221, w2222, w2223, w2224, w2225, w2226, w2227, w2228, w2229, w2230, w2231, w2232, w2233, w2234, w2235, w2236, w2237, w2238, w2239, w2240, w2241, w2242, w2243, w2244, w2245, w2246, w2247, w2248, w2249, w2250, w2251, w2252, w2253, w2254, w2255, w2256, w2257, w2258, w2259, w2260, w2261, w2262, w2263, w2264, w2265, w2266, w2267, w2268, w2269, w2270, w2271, w2272, w2273, w2274, w2275, w2276, w2277, w2278, w2279, w2280, w2281, w2282, w2283, w2284, w2285, w2286, w2287, w2288, w2289, w2290, w2291, w2292, w2293, w2294, w2295, w2296, w2297, w2298, w2299, w2300, w2301, w2302, w2303, w2304, w2305, w2306, w2307, w2308, w2309, w2310, w2311, w2312, w2313, w2314, w2315, w2316, w2317, w2318, w2319, w2320, w2321, w2322, w2323, w2324, w2325, w2326, w2327, w2328, w2329, w2330, w2331, w2332, w2333, w2334, w2335, w2336, w2337, w2338, w2339, w2340, w2341, w2342, w2343, w2344, w2345, w2346, w2347, w2348, w2349, w2350, w2351, w2352, w2353, w2354, w2355, w2356, w2357, w2358, w2359, w2360, w2361, w2362, w2363, w2364, w2365, w2366, w2367, w2368, w2369, w2370, w2371, w2372, w2373, w2374, w2375, w2376, w2377, w2378, w2379, w2380, w2381, w2382, w2383, w2384, w2385, w2386, w2387, w2388, w2389, w2390, w2391, w2392, w2393, w2394, w2395, w2396, w2397, w2398, w2399, w2400, w2401, w2402, w2403, w2404, w2405, w2406, w2407, w2408, w2409, w2410, w2411, w2412, w2413, w2414, w2415, w2416, w2417, w2418, w2419, w2420, w2421, w2422, w2423, w2424, w2425, w2426, w2427, w2428, w2429, w2430, w2431, w2432, w2433, w2434, w2435, w2436, w2437, w2438, w2439, w2440, w2441, w2442, w2443, w2444, w2445, w2446, w2447, w2448, w2449, w2450, w2451, w2452, w2453, w2454, w2455, w2456, w2457, w2458, w2459, w2460, w2461, w2462, w2463, w2464, w2465, w2466, w2467, w2468, w2469, w2470, w2471, w2472, w2473, w2474, w2475, w2476, w2477, w2478, w2479, w2480, w2481, w2482, w2483, w2484, w2485, w2486, w2487, w2488, w2489, w2490, w2491, w2492, w2493, w2494, w2495, w2496, w2497, w2498, w2499, w2500, w2501, w2502, w2503, w2504, w2505, w2506, w2507, w2508, w2509, w2510, w2511, w2512, w2513, w2514, w2515, w2516, w2517, w2518, w2519, w2520, w2521, w2522, w2523, w2524, w2525, w2526, w2527, w2528, w2529, w2530, w2531, w2532, w2533, w2534, w2535, w2536, w2537, w2538, w2539, w2540, w2541, w2542, w2543, w2544, w2545, w2546, w2547, w2548, w2549, w2550, w2551, w2552, w2553, w2554, w2555, w2556, w2557, w2558, w2559, w2560, w2561, w2562, w2563, w2564, w2565, w2566, w2567, w2568, w2569, w2570, w2571, w2572, w2573, w2574, w2575, w2576, w2577, w2578, w2579, w2580, w2581, w2582, w2583, w2584, w2585, w2586, w2587, w2588, w2589, w2590, w2591, w2592, w2593, w2594, w2595, w2596, w2597, w2598, w2599, w2600, w2601, w2602, w2603, w2604, w2605, w2606, w2607, w2608, w2609, w2610, w2611, w2612, w2613, w2614, w2615, w2616, w2617, w2618, w2619, w2620, w2621, w2622, w2623, w2624, w2625, w2626, w2627, w2628, w2629, w2630, w2631, w2632, w2633, w2634, w2635, w2636, w2637, w2638, w2639, w2640, w2641, w2642, w2643, w2644, w2645, w2646, w2647, w2648, w2649, w2650, w2651, w2652, w2653, w2654, w2655, w2656, w2657, w2658, w2659, w2660, w2661, w2662, w2663, w2664, w2665, w2666, w2667, w2668, w2669, w2670, w2671, w2672, w2673, w2674, w2675, w2676, w2677, w2678, w2679, w2680, w2681, w2682, w2683, w2684, w2685, w2686, w2687, w2688, w2689, w2690, w2691, w2692, w2693, w2694, w2695, w2696, w2697, w2698, w2699, w2700, w2701, w2702, w2703, w2704, w2705, w2706, w2707, w2708, w2709, w2710, w2711, w2712, w2713, w2714, w2715, w2716, w2717, w2718, w2719, w2720, w2721, w2722, w2723, w2724, w2725, w2726, w2727, w2728, w2729, w2730, w2731, w2732, w2733, w2734, w2735, w2736, w2737, w2738, w2739, w2740, w2741, w2742, w2743, w2744, w2745, w2746, w2747, w2748, w2749, w2750, w2751, w2752, w2753, w2754, w2755, w2756, w2757, w2758, w2759, w2760, w2761, w2762, w2763, w2764, w2765, w2766, w2767, w2768, w2769, w2770, w2771, w2772, w2773, w2774, w2775, w2776, w2777, w2778, w2779, w2780, w2781, w2782, w2783, w2784, w2785, w2786, w2787, w2788, w2789, w2790, w2791, w2792, w2793, w2794, w2795, w2796, w2797, w2798, w2799, w2800, w2801, w2802, w2803, w2804, w2805, w2806, w2807, w2808, w2809, w2810, w2811, w2812, w2813, w2814, w2815, w2816, w2817, w2818, w2819, w2820, w2821, w2822, w2823, w2824, w2825, w2826, w2827, w2828, w2829, w2830, w2831, w2832, w2833, w2834, w2835, w2836, w2837, w2838, w2839, w2840, w2841, w2842, w2843, w2844, w2845, w2846, w2847, w2848, w2849, w2850, w2851, w2852, w2853, w2854, w2855, w2856, w2857, w2858, w2859, w2860, w2861, w2862, w2863, w2864, w2865, w2866, w2867, w2868, w2869, w2870, w2871, w2872, w2873, w2874, w2875, w2876, w2877, w2878, w2879, w2880, w2881, w2882, w2883, w2884, w2885, w2886, w2887, w2888, w2889, w2890, w2891, w2892, w2893, w2894, w2895, w2896, w2897, w2898, w2899, w2900, w2901, w2902, w2903, w2904, w2905, w2906, w2907, w2908, w2909, w2910, w2911, w2912, w2913, w2914, w2915, w2916, w2917, w2918, w2919, w2920, w2921, w2922, w2923, w2924, w2925, w2926, w2927, w2928, w2929, w2930, w2931, w2932, w2933, w2934, w2935, w2936, w2937, w2938, w2939, w2940, w2941, w2942, w2943, w2944, w2945, w2946, w2947, w2948, w2949, w2950, w2951, w2952, w2953, w2954, w2955, w2956, w2957, w2958, w2959, w2960, w2961, w2962, w2963, w2964, w2965, w2966, w2967, w2968, w2969, w2970, w2971, w2972, w2973, w2974, w2975, w2976, w2977, w2978, w2979, w2980, w2981, w2982, w2983, w2984, w2985, w2986, w2987, w2988, w2989, w2990, w2991, w2992, w2993, w2994, w2995, w2996, w2997, w2998, w2999, w3000, w3001, w3002, w3003, w3004, w3005, w3006, w3007, w3008, w3009, w3010, w3011, w3012, w3013, w3014, w3015, w3016, w3017, w3018, w3019, w3020, w3021, w3022, w3023, w3024, w3025, w3026, w3027, w3028, w3029, w3030, w3031, w3032, w3033, w3034, w3035, w3036, w3037, w3038, w3039, w3040, w3041, w3042, w3043, w3044, w3045, w3046, w3047, w3048, w3049, w3050, w3051, w3052, w3053, w3054, w3055, w3056, w3057, w3058, w3059, w3060, w3061, w3062, w3063, w3064, w3065, w3066, w3067, w3068, w3069, w3070, w3071, w3072, w3073, w3074, w3075, w3076, w3077, w3078, w3079, w3080, w3081, w3082, w3083, w3084, w3085, w3086, w3087, w3088, w3089, w3090, w3091, w3092, w3093, w3094, w3095, w3096, w3097, w3098, w3099, w3100, w3101, w3102, w3103, w3104, w3105, w3106, w3107, w3108, w3109, w3110, w3111, w3112, w3113, w3114, w3115, w3116, w3117, w3118, w3119, w3120, w3121, w3122, w3123, w3124, w3125, w3126, w3127, w3128, w3129, w3130, w3131, w3132, w3133, w3134, w3135, w3136, w3137, w3138, w3139, w3140, w3141, w3142, w3143, w3144, w3145, w3146, w3147, w3148, w3149, w3150, w3151, w3152, w3153, w3154, w3155, w3156, w3157, w3158, w3159, w3160, w3161, w3162, w3163, w3164, w3165, w3166, w3167, w3168, w3169, w3170, w3171, w3172, w3173, w3174, w3175, w3176, w3177, w3178, w3179, w3180, w3181, w3182, w3183, w3184, w3185, w3186, w3187, w3188, w3189, w3190, w3191, w3192, w3193, w3194, w3195, w3196, w3197, w3198, w3199, w3200, w3201, w3202, w3203, w3204, w3205, w3206, w3207, w3208, w3209, w3210, w3211, w3212, w3213, w3214, w3215, w3216, w3217, w3218, w3219, w3220, w3221, w3222, w3223, w3224, w3225, w3226, w3227, w3228, w3229, w3230, w3231, w3232, w3233, w3234, w3235, w3236, w3237, w3238, w3239, w3240, w3241, w3242, w3243, w3244, w3245, w3246, w3247, w3248, w3249, w3250, w3251, w3252, w3253, w3254, w3255, w3256, w3257, w3258, w3259, w3260, w3261, w3262, w3263, w3264, w3265, w3266, w3267, w3268, w3269, w3270, w3271, w3272, w3273, w3274, w3275, w3276, w3277, w3278, w3279, w3280, w3281, w3282, w3283, w3284, w3285, w3286, w3287, w3288, w3289, w3290, w3291, w3292, w3293, w3294, w3295, w3296, w3297, w3298, w3299, w3300, w3301, w3302, w3303, w3304, w3305, w3306, w3307, w3308, w3309, w3310, w3311, w3312, w3313, w3314, w3315, w3316, w3317, w3318, w3319, w3320, w3321, w3322, w3323, w3324, w3325, w3326, w3327, w3328, w3329, w3330, w3331, w3332, w3333, w3334, w3335, w3336, w3337, w3338, w3339, w3340, w3341, w3342, w3343, w3344, w3345, w3346, w3347, w3348, w3349, w3350, w3351, w3352, w3353, w3354, w3355, w3356, w3357, w3358, w3359, w3360, w3361, w3362, w3363, w3364, w3365, w3366, w3367, w3368, w3369, w3370, w3371, w3372, w3373, w3374, w3375, w3376, w3377, w3378, w3379, w3380, w3381, w3382, w3383, w3384, w3385, w3386, w3387, w3388, w3389, w3390, w3391, w3392, w3393, w3394, w3395, w3396, w3397, w3398, w3399, w3400, w3401, w3402, w3403, w3404, w3405, w3406, w3407, w3408, w3409, w3410, w3411, w3412, w3413, w3414, w3415, w3416, w3417, w3418, w3419, w3420, w3421, w3422, w3423, w3424, w3425, w3426, w3427, w3428, w3429, w3430, w3431, w3432, w3433, w3434, w3435, w3436, w3437, w3438, w3439, w3440, w3441, w3442, w3443, w3444, w3445, w3446, w3447, w3448, w3449, w3450, w3451, w3452, w3453, w3454, w3455, w3456, w3457, w3458, w3459, w3460, w3461, w3462, w3463, w3464, w3465, w3466, w3467, w3468, w3469, w3470, w3471, w3472, w3473, w3474, w3475, w3476, w3477, w3478, w3479, w3480, w3481, w3482, w3483, w3484, w3485, w3486, w3487, w3488, w3489, w3490, w3491, w3492, w3493, w3494, w3495, w3496, w3497, w3498, w3499, w3500, w3501, w3502, w3503, w3504, w3505, w3506, w3507, w3508, w3509, w3510, w3511, w3512, w3513, w3514, w3515, w3516, w3517, w3518, w3519, w3520, w3521, w3522, w3523, w3524, w3525, w3526, w3527, w3528, w3529, w3530, w3531, w3532, w3533, w3534, w3535, w3536, w3537, w3538, w3539, w3540, w3541, w3542, w3543, w3544, w3545, w3546, w3547, w3548, w3549, w3550, w3551, w3552, w3553, w3554, w3555, w3556, w3557, w3558, w3559, w3560, w3561, w3562, w3563, w3564, w3565, w3566, w3567, w3568, w3569, w3570, w3571, w3572, w3573, w3574, w3575, w3576, w3577, w3578, w3579, w3580, w3581, w3582, w3583, w3584, w3585, w3586, w3587, w3588, w3589, w3590, w3591, w3592, w3593, w3594, w3595, w3596, w3597, w3598, w3599, w3600, w3601, w3602, w3603, w3604, w3605, w3606, w3607, w3608, w3609, w3610, w3611, w3612, w3613, w3614, w3615, w3616, w3617, w3618, w3619, w3620, w3621, w3622, w3623, w3624, w3625, w3626, w3627, w3628, w3629, w3630, w3631, w3632, w3633, w3634, w3635, w3636, w3637, w3638, w3639, w3640, w3641, w3642, w3643, w3644, w3645, w3646, w3647, w3648, w3649, w3650, w3651, w3652, w3653, w3654, w3655, w3656, w3657, w3658, w3659, w3660, w3661, w3662, w3663, w3664, w3665, w3666, w3667, w3668, w3669, w3670, w3671, w3672, w3673, w3674, w3675, w3676, w3677, w3678, w3679, w3680, w3681, w3682, w3683, w3684, w3685, w3686, w3687, w3688, w3689, w3690, w3691, w3692, w3693, w3694, w3695, w3696, w3697, w3698, w3699, w3700, w3701, w3702, w3703, w3704, w3705, w3706, w3707, w3708, w3709, w3710, w3711, w3712, w3713, w3714, w3715, w3716, w3717, w3718, w3719, w3720, w3721, w3722, w3723, w3724, w3725, w3726, w3727, w3728, w3729, w3730, w3731, w3732, w3733, w3734, w3735, w3736, w3737, w3738, w3739, w3740, w3741, w3742, w3743, w3744, w3745, w3746, w3747, w3748, w3749, w3750, w3751, w3752, w3753, w3754, w3755, w3756, w3757, w3758, w3759, w3760, w3761, w3762, w3763, w3764, w3765, w3766, w3767, w3768, w3769, w3770, w3771, w3772, w3773, w3774, w3775, w3776, w3777, w3778, w3779, w3780, w3781, w3782, w3783, w3784, w3785, w3786, w3787, w3788, w3789, w3790, w3791, w3792, w3793, w3794, w3795, w3796, w3797, w3798, w3799, w3800, w3801, w3802, w3803, w3804, w3805, w3806, w3807, w3808, w3809, w3810, w3811, w3812, w3813, w3814, w3815, w3816, w3817, w3818, w3819, w3820, w3821, w3822, w3823, w3824, w3825, w3826, w3827, w3828, w3829, w3830, w3831, w3832, w3833, w3834, w3835, w3836, w3837, w3838, w3839, w3840, w3841, w3842, w3843, w3844, w3845, w3846, w3847, w3848, w3849, w3850, w3851, w3852, w3853, w3854, w3855, w3856, w3857, w3858, w3859, w3860, w3861, w3862, w3863, w3864, w3865, w3866, w3867, w3868, w3869, w3870, w3871, w3872, w3873, w3874, w3875, w3876, w3877, w3878, w3879, w3880, w3881, w3882, w3883, w3884, w3885, w3886, w3887, w3888, w3889, w3890, w3891, w3892, w3893, w3894, w3895, w3896, w3897, w3898, w3899, w3900, w3901, w3902, w3903, w3904, w3905, w3906, w3907, w3908, w3909, w3910, w3911, w3912, w3913, w3914, w3915, w3916, w3917, w3918, w3919, w3920, w3921, w3922, w3923, w3924, w3925, w3926, w3927, w3928, w3929, w3930, w3931, w3932, w3933, w3934, w3935, w3936, w3937, w3938, w3939, w3940, w3941, w3942, w3943, w3944, w3945, w3946, w3947, w3948, w3949, w3950, w3951, w3952, w3953, w3954, w3955, w3956, w3957, w3958, w3959, w3960, w3961, w3962, w3963, w3964, w3965, w3966, w3967, w3968, w3969, w3970, w3971, w3972, w3973, w3974, w3975, w3976, w3977, w3978, w3979, w3980, w3981, w3982, w3983, w3984, w3985, w3986, w3987, w3988, w3989, w3990, w3991, w3992, w3993, w3994, w3995, w3996, w3997, w3998, w3999, w4000, w4001, w4002, w4003, w4004, w4005, w4006, w4007, w4008, w4009, w4010, w4011, w4012, w4013, w4014, w4015, w4016, w4017, w4018, w4019, w4020, w4021, w4022, w4023, w4024, w4025, w4026, w4027, w4028, w4029, w4030, w4031, w4032, w4033, w4034, w4035, w4036, w4037, w4038, w4039, w4040, w4041, w4042, w4043, w4044, w4045, w4046, w4047, w4048, w4049, w4050, w4051, w4052, w4053, w4054, w4055, w4056, w4057, w4058, w4059, w4060, w4061, w4062, w4063, w4064, w4065, w4066, w4067, w4068, w4069, w4070, w4071, w4072, w4073, w4074, w4075, w4076, w4077, w4078, w4079, w4080, w4081, w4082, w4083, w4084, w4085, w4086, w4087, w4088, w4089, w4090, w4091, w4092, w4093, w4094, w4095, w4096, w4097, w4098, w4099, w4100, w4101, w4102, w4103, w4104, w4105, w4106, w4107, w4108, w4109, w4110, w4111, w4112, w4113, w4114, w4115, w4116, w4117, w4118, w4119, w4120, w4121, w4122, w4123, w4124, w4125, w4126, w4127, w4128, w4129, w4130, w4131, w4132, w4133, w4134, w4135, w4136, w4137, w4138, w4139, w4140, w4141, w4142, w4143, w4144, w4145, w4146, w4147, w4148, w4149, w4150, w4151, w4152, w4153, w4154, w4155, w4156, w4157, w4158, w4159, w4160, w4161, w4162, w4163, w4164, w4165, w4166, w4167, w4168, w4169, w4170, w4171, w4172, w4173, w4174, w4175, w4176, w4177, w4178, w4179, w4180, w4181, w4182, w4183, w4184, w4185, w4186, w4187, w4188, w4189, w4190, w4191, w4192, w4193, w4194, w4195, w4196, w4197, w4198, w4199, w4200, w4201, w4202, w4203, w4204, w4205, w4206, w4207, w4208, w4209, w4210, w4211, w4212, w4213, w4214, w4215, w4216, w4217, w4218, w4219, w4220, w4221, w4222, w4223, w4224, w4225, w4226, w4227, w4228, w4229, w4230, w4231, w4232, w4233, w4234, w4235, w4236, w4237, w4238, w4239, w4240, w4241, w4242, w4243, w4244, w4245, w4246, w4247, w4248, w4249, w4250, w4251, w4252, w4253, w4254, w4255, w4256, w4257, w4258, w4259, w4260, w4261, w4262, w4263, w4264, w4265, w4266, w4267, w4268, w4269, w4270, w4271, w4272, w4273, w4274, w4275, w4276, w4277, w4278, w4279, w4280, w4281, w4282, w4283, w4284, w4285, w4286, w4287, w4288, w4289, w4290, w4291, w4292, w4293, w4294, w4295, w4296, w4297, w4298, w4299, w4300, w4301, w4302, w4303, w4304, w4305, w4306, w4307, w4308, w4309, w4310, w4311, w4312, w4313, w4314, w4315, w4316, w4317, w4318, w4319, w4320, w4321, w4322, w4323, w4324, w4325, w4326, w4327, w4328, w4329, w4330, w4331, w4332, w4333, w4334, w4335, w4336, w4337, w4338, w4339, w4340, w4341, w4342, w4343, w4344, w4345, w4346, w4347, w4348, w4349, w4350, w4351, w4352, w4353, w4354, w4355, w4356, w4357, w4358, w4359, w4360, w4361, w4362, w4363, w4364, w4365, w4366, w4367, w4368, w4369, w4370, w4371, w4372, w4373, w4374, w4375, w4376, w4377, w4378, w4379, w4380, w4381, w4382, w4383, w4384, w4385, w4386, w4387, w4388, w4389, w4390, w4391, w4392, w4393, w4394, w4395, w4396, w4397, w4398, w4399, w4400, w4401, w4402, w4403, w4404, w4405, w4406, w4407, w4408, w4409, w4410, w4411, w4412, w4413, w4414, w4415, w4416, w4417, w4418, w4419, w4420, w4421, w4422, w4423, w4424, w4425, w4426, w4427, w4428, w4429, w4430, w4431, w4432, w4433, w4434, w4435, w4436, w4437, w4438, w4439, w4440, w4441, w4442, w4443, w4444, w4445, w4446, w4447, w4448, w4449, w4450, w4451, w4452, w4453, w4454, w4455, w4456, w4457, w4458, w4459, w4460, w4461, w4462, w4463, w4464, w4465, w4466, w4467, w4468, w4469, w4470, w4471, w4472, w4473, w4474, w4475, w4476, w4477, w4478, w4479, w4480, w4481, w4482, w4483, w4484, w4485, w4486, w4487, w4488, w4489, w4490, w4491, w4492, w4493, w4494, w4495, w4496, w4497, w4498, w4499, w4500, w4501, w4502, w4503, w4504, w4505, w4506, w4507, w4508, w4509, w4510, w4511, w4512, w4513, w4514, w4515, w4516, w4517, w4518, w4519, w4520, w4521, w4522, w4523, w4524, w4525, w4526, w4527, w4528, w4529, w4530, w4531, w4532, w4533, w4534, w4535, w4536, w4537, w4538, w4539, w4540, w4541, w4542, w4543, w4544, w4545, w4546, w4547, w4548, w4549, w4550, w4551, w4552, w4553, w4554, w4555, w4556, w4557, w4558, w4559, w4560, w4561, w4562, w4563, w4564, w4565, w4566, w4567, w4568, w4569, w4570, w4571, w4572, w4573, w4574, w4575, w4576, w4577, w4578, w4579, w4580, w4581, w4582, w4583, w4584, w4585, w4586, w4587, w4588, w4589, w4590, w4591, w4592, w4593, w4594, w4595, w4596, w4597, w4598, w4599, w4600, w4601, w4602, w4603, w4604, w4605, w4606, w4607, w4608, w4609, w4610, w4611, w4612, w4613, w4614, w4615, w4616, w4617, w4618, w4619, w4620, w4621, w4622, w4623, w4624, w4625, w4626, w4627, w4628, w4629, w4630, w4631, w4632, w4633, w4634, w4635, w4636, w4637, w4638, w4639, w4640, w4641, w4642, w4643, w4644, w4645, w4646, w4647, w4648, w4649, w4650, w4651, w4652, w4653, w4654, w4655, w4656, w4657, w4658, w4659, w4660, w4661, w4662, w4663, w4664, w4665, w4666, w4667, w4668, w4669, w4670, w4671, w4672, w4673, w4674, w4675, w4676, w4677, w4678, w4679, w4680, w4681, w4682, w4683, w4684, w4685, w4686, w4687, w4688, w4689, w4690, w4691, w4692, w4693, w4694, w4695, w4696, w4697, w4698, w4699, w4700, w4701, w4702, w4703, w4704, w4705, w4706, w4707, w4708, w4709, w4710, w4711, w4712, w4713, w4714, w4715, w4716, w4717, w4718, w4719, w4720, w4721, w4722, w4723, w4724, w4725, w4726, w4727, w4728, w4729, w4730, w4731, w4732, w4733, w4734, w4735, w4736, w4737, w4738, w4739, w4740, w4741, w4742, w4743, w4744, w4745, w4746, w4747, w4748, w4749, w4750, w4751, w4752, w4753, w4754, w4755, w4756, w4757, w4758, w4759, w4760, w4761, w4762, w4763, w4764, w4765, w4766, w4767, w4768, w4769, w4770, w4771, w4772, w4773, w4774, w4775, w4776, w4777, w4778, w4779, w4780, w4781, w4782, w4783, w4784, w4785, w4786, w4787, w4788, w4789, w4790, w4791, w4792, w4793, w4794, w4795, w4796, w4797, w4798, w4799, w4800, w4801, w4802, w4803, w4804, w4805, w4806, w4807, w4808, w4809, w4810, w4811, w4812, w4813, w4814, w4815, w4816, w4817, w4818, w4819, w4820, w4821, w4822, w4823, w4824, w4825, w4826, w4827, w4828, w4829, w4830, w4831, w4832, w4833, w4834, w4835, w4836, w4837, w4838, w4839, w4840, w4841, w4842, w4843, w4844, w4845, w4846, w4847, w4848, w4849, w4850, w4851, w4852, w4853, w4854, w4855, w4856, w4857, w4858, w4859, w4860, w4861, w4862, w4863, w4864, w4865, w4866, w4867, w4868, w4869, w4870, w4871, w4872, w4873, w4874, w4875, w4876, w4877, w4878, w4879, w4880, w4881, w4882, w4883, w4884, w4885, w4886, w4887, w4888, w4889, w4890, w4891, w4892, w4893, w4894, w4895, w4896, w4897, w4898, w4899, w4900, w4901, w4902, w4903, w4904, w4905, w4906, w4907, w4908, w4909, w4910, w4911, w4912, w4913, w4914, w4915, w4916, w4917, w4918, w4919, w4920, w4921, w4922, w4923, w4924, w4925, w4926, w4927, w4928, w4929, w4930, w4931, w4932, w4933, w4934, w4935, w4936, w4937, w4938, w4939, w4940, w4941, w4942, w4943, w4944, w4945, w4946, w4947, w4948, w4949, w4950, w4951, w4952, w4953, w4954, w4955, w4956, w4957, w4958, w4959, w4960, w4961, w4962, w4963, w4964, w4965, w4966, w4967, w4968, w4969, w4970, w4971, w4972, w4973, w4974, w4975, w4976, w4977, w4978, w4979, w4980, w4981, w4982, w4983, w4984, w4985, w4986, w4987, w4988, w4989, w4990, w4991, w4992, w4993, w4994, w4995, w4996, w4997, w4998, w4999, w5000, w5001, w5002, w5003, w5004, w5005, w5006, w5007, w5008, w5009, w5010, w5011, w5012, w5013, w5014, w5015, w5016, w5017, w5018, w5019, w5020, w5021, w5022, w5023, w5024, w5025, w5026, w5027, w5028, w5029, w5030, w5031, w5032, w5033, w5034, w5035, w5036, w5037, w5038, w5039, w5040, w5041, w5042, w5043, w5044, w5045, w5046, w5047, w5048, w5049, w5050, w5051, w5052, w5053, w5054, w5055, w5056, w5057, w5058, w5059, w5060, w5061, w5062, w5063, w5064, w5065, w5066, w5067, w5068, w5069, w5070, w5071, w5072, w5073, w5074, w5075, w5076, w5077, w5078, w5079, w5080, w5081, w5082, w5083, w5084, w5085, w5086, w5087, w5088, w5089, w5090, w5091, w5092, w5093, w5094, w5095, w5096, w5097, w5098, w5099, w5100, w5101, w5102, w5103, w5104, w5105, w5106, w5107, w5108, w5109, w5110, w5111, w5112, w5113, w5114, w5115, w5116, w5117, w5118, w5119, w5120, w5121, w5122, w5123, w5124, w5125, w5126, w5127, w5128, w5129, w5130, w5131, w5132, w5133, w5134, w5135, w5136, w5137, w5138, w5139, w5140, w5141, w5142, w5143, w5144, w5145, w5146, w5147, w5148, w5149, w5150, w5151, w5152, w5153, w5154, w5155, w5156, w5157, w5158, w5159, w5160, w5161, w5162, w5163, w5164, w5165, w5166, w5167, w5168, w5169, w5170, w5171, w5172, w5173, w5174, w5175, w5176, w5177, w5178, w5179, w5180, w5181, w5182, w5183, w5184, w5185, w5186, w5187, w5188, w5189, w5190, w5191, w5192, w5193, w5194, w5195, w5196, w5197, w5198, w5199, w5200, w5201, w5202, w5203, w5204, w5205, w5206, w5207, w5208, w5209, w5210, w5211, w5212, w5213, w5214, w5215, w5216, w5217, w5218, w5219, w5220, w5221, w5222, w5223, w5224, w5225, w5226, w5227, w5228, w5229, w5230, w5231, w5232, w5233, w5234, w5235, w5236, w5237, w5238, w5239, w5240, w5241, w5242, w5243, w5244, w5245, w5246, w5247, w5248, w5249, w5250, w5251, w5252, w5253, w5254, w5255, w5256, w5257, w5258, w5259, w5260, w5261, w5262, w5263, w5264, w5265, w5266, w5267, w5268, w5269, w5270, w5271, w5272, w5273, w5274, w5275, w5276, w5277, w5278, w5279, w5280, w5281, w5282, w5283, w5284, w5285, w5286, w5287, w5288, w5289, w5290, w5291, w5292, w5293, w5294, w5295, w5296, w5297, w5298, w5299, w5300, w5301, w5302, w5303, w5304, w5305, w5306, w5307, w5308, w5309, w5310, w5311, w5312, w5313, w5314, w5315, w5316, w5317, w5318, w5319, w5320, w5321, w5322, w5323, w5324, w5325, w5326, w5327, w5328, w5329, w5330, w5331, w5332, w5333, w5334, w5335, w5336, w5337, w5338, w5339, w5340, w5341, w5342, w5343, w5344, w5345, w5346, w5347, w5348, w5349, w5350, w5351, w5352, w5353, w5354, w5355, w5356, w5357, w5358, w5359, w5360, w5361, w5362, w5363, w5364, w5365, w5366, w5367, w5368, w5369, w5370, w5371, w5372, w5373, w5374, w5375, w5376, w5377, w5378, w5379, w5380, w5381, w5382, w5383, w5384, w5385, w5386, w5387, w5388, w5389, w5390, w5391, w5392, w5393, w5394, w5395, w5396, w5397, w5398, w5399, w5400, w5401, w5402, w5403, w5404, w5405, w5406, w5407, w5408, w5409, w5410, w5411, w5412, w5413, w5414, w5415, w5416, w5417, w5418, w5419, w5420, w5421, w5422, w5423, w5424, w5425, w5426, w5427, w5428, w5429, w5430, w5431, w5432, w5433, w5434, w5435, w5436, w5437, w5438, w5439, w5440, w5441, w5442, w5443, w5444, w5445, w5446, w5447, w5448, w5449, w5450, w5451, w5452, w5453, w5454, w5455, w5456, w5457, w5458, w5459, w5460, w5461, w5462, w5463, w5464, w5465, w5466, w5467, w5468, w5469, w5470, w5471, w5472, w5473, w5474, w5475, w5476, w5477, w5478, w5479, w5480, w5481, w5482, w5483, w5484, w5485, w5486, w5487, w5488, w5489, w5490, w5491, w5492, w5493, w5494, w5495, w5496, w5497, w5498, w5499, w5500, w5501, w5502, w5503, w5504, w5505, w5506, w5507, w5508, w5509, w5510, w5511, w5512, w5513, w5514, w5515, w5516, w5517, w5518, w5519, w5520, w5521, w5522, w5523, w5524, w5525, w5526, w5527, w5528, w5529, w5530, w5531, w5532, w5533, w5534, w5535, w5536, w5537, w5538, w5539, w5540, w5541, w5542, w5543, w5544, w5545, w5546, w5547, w5548, w5549, w5550, w5551, w5552, w5553, w5554, w5555, w5556, w5557, w5558, w5559, w5560, w5561, w5562, w5563, w5564, w5565, w5566, w5567, w5568, w5569, w5570, w5571, w5572, w5573, w5574, w5575, w5576, w5577, w5578, w5579, w5580, w5581, w5582, w5583, w5584, w5585, w5586, w5587, w5588, w5589, w5590, w5591, w5592, w5593, w5594, w5595, w5596, w5597, w5598, w5599, w5600, w5601, w5602, w5603, w5604, w5605, w5606, w5607, w5608, w5609, w5610, w5611, w5612, w5613, w5614, w5615, w5616, w5617, w5618, w5619, w5620, w5621, w5622, w5623, w5624, w5625, w5626, w5627, w5628, w5629, w5630, w5631, w5632, w5633, w5634, w5635, w5636, w5637, w5638, w5639, w5640, w5641, w5642, w5643, w5644, w5645, w5646, w5647, w5648, w5649, w5650, w5651, w5652, w5653, w5654, w5655, w5656, w5657, w5658, w5659, w5660, w5661, w5662, w5663, w5664, w5665, w5666, w5667, w5668, w5669, w5670, w5671, w5672, w5673, w5674, w5675, w5676, w5677, w5678, w5679, w5680, w5681, w5682, w5683, w5684, w5685, w5686, w5687, w5688, w5689, w5690, w5691, w5692, w5693, w5694, w5695, w5696, w5697, w5698, w5699, w5700, w5701, w5702, w5703, w5704, w5705, w5706, w5707, w5708, w5709, w5710, w5711, w5712, w5713, w5714, w5715, w5716, w5717, w5718, w5719, w5720, w5721, w5722, w5723, w5724, w5725, w5726, w5727, w5728, w5729, w5730, w5731, w5732, w5733, w5734, w5735, w5736, w5737, w5738, w5739, w5740, w5741, w5742, w5743, w5744, w5745, w5746, w5747, w5748, w5749, w5750, w5751, w5752, w5753, w5754, w5755, w5756, w5757, w5758, w5759, w5760, w5761, w5762, w5763, w5764, w5765, w5766, w5767, w5768, w5769, w5770, w5771, w5772, w5773, w5774, w5775, w5776, w5777, w5778, w5779, w5780, w5781, w5782, w5783, w5784, w5785, w5786, w5787, w5788, w5789, w5790, w5791, w5792, w5793, w5794, w5795, w5796, w5797, w5798, w5799, w5800, w5801, w5802, w5803, w5804, w5805, w5806, w5807, w5808, w5809, w5810, w5811, w5812, w5813, w5814, w5815, w5816, w5817, w5818, w5819, w5820, w5821, w5822, w5823, w5824, w5825, w5826, w5827, w5828, w5829, w5830, w5831, w5832, w5833, w5834, w5835, w5836, w5837, w5838, w5839, w5840, w5841, w5842, w5843, w5844, w5845, w5846, w5847, w5848, w5849, w5850, w5851, w5852, w5853, w5854, w5855, w5856, w5857, w5858, w5859, w5860, w5861, w5862, w5863, w5864, w5865, w5866, w5867, w5868, w5869, w5870, w5871, w5872, w5873, w5874, w5875, w5876, w5877, w5878, w5879, w5880, w5881, w5882, w5883, w5884, w5885, w5886, w5887, w5888, w5889, w5890, w5891, w5892, w5893, w5894, w5895, w5896, w5897, w5898, w5899, w5900, w5901, w5902, w5903, w5904, w5905, w5906, w5907, w5908, w5909, w5910, w5911, w5912, w5913, w5914, w5915, w5916, w5917, w5918, w5919, w5920, w5921, w5922, w5923, w5924, w5925, w5926, w5927, w5928, w5929, w5930, w5931, w5932, w5933, w5934, w5935, w5936, w5937, w5938, w5939, w5940, w5941, w5942, w5943, w5944, w5945, w5946, w5947, w5948, w5949, w5950, w5951, w5952, w5953, w5954, w5955, w5956, w5957, w5958, w5959, w5960, w5961, w5962, w5963, w5964, w5965, w5966, w5967, w5968, w5969, w5970, w5971, w5972, w5973, w5974, w5975, w5976, w5977, w5978, w5979, w5980, w5981, w5982, w5983, w5984, w5985, w5986, w5987, w5988, w5989, w5990, w5991, w5992, w5993, w5994, w5995, w5996, w5997, w5998, w5999, w6000, w6001, w6002, w6003, w6004, w6005, w6006, w6007, w6008, w6009, w6010, w6011, w6012, w6013, w6014, w6015, w6016, w6017, w6018, w6019, w6020, w6021, w6022, w6023, w6024, w6025, w6026, w6027, w6028, w6029, w6030, w6031, w6032, w6033, w6034, w6035, w6036, w6037, w6038, w6039, w6040, w6041, w6042, w6043, w6044, w6045, w6046, w6047, w6048, w6049, w6050, w6051, w6052, w6053, w6054, w6055, w6056, w6057, w6058, w6059, w6060, w6061, w6062, w6063, w6064, w6065, w6066, w6067, w6068, w6069, w6070, w6071, w6072, w6073, w6074, w6075, w6076, w6077, w6078, w6079, w6080, w6081, w6082, w6083, w6084, w6085, w6086, w6087, w6088, w6089, w6090, w6091, w6092, w6093, w6094, w6095, w6096, w6097, w6098, w6099, w6100, w6101, w6102, w6103, w6104, w6105, w6106, w6107, w6108, w6109, w6110, w6111, w6112, w6113, w6114, w6115, w6116, w6117, w6118, w6119, w6120, w6121, w6122, w6123, w6124, w6125, w6126, w6127, w6128, w6129, w6130, w6131, w6132, w6133, w6134, w6135, w6136, w6137, w6138, w6139, w6140, w6141, w6142, w6143, w6144, w6145, w6146, w6147, w6148, w6149, w6150, w6151, w6152, w6153, w6154, w6155, w6156, w6157, w6158, w6159, w6160, w6161, w6162, w6163, w6164, w6165, w6166, w6167, w6168, w6169, w6170, w6171, w6172, w6173, w6174, w6175, w6176, w6177, w6178, w6179, w6180, w6181, w6182, w6183, w6184, w6185, w6186, w6187, w6188, w6189, w6190, w6191, w6192, w6193, w6194, w6195, w6196, w6197, w6198, w6199, w6200, w6201, w6202, w6203, w6204, w6205, w6206, w6207, w6208, w6209, w6210, w6211, w6212, w6213, w6214, w6215, w6216, w6217, w6218, w6219, w6220, w6221, w6222, w6223, w6224, w6225, w6226, w6227, w6228, w6229, w6230, w6231, w6232, w6233, w6234, w6235, w6236, w6237, w6238, w6239, w6240, w6241, w6242, w6243, w6244, w6245, w6246, w6247, w6248, w6249, w6250, w6251, w6252, w6253, w6254, w6255, w6256, w6257, w6258, w6259, w6260, w6261, w6262, w6263, w6264, w6265, w6266, w6267, w6268, w6269, w6270, w6271, w6272, w6273, w6274, w6275, w6276, w6277, w6278, w6279, w6280, w6281, w6282, w6283, w6284, w6285, w6286, w6287, w6288, w6289, w6290, w6291, w6292, w6293, w6294, w6295, w6296, w6297, w6298, w6299, w6300, w6301, w6302, w6303, w6304, w6305, w6306, w6307, w6308, w6309, w6310, w6311, w6312, w6313, w6314, w6315, w6316, w6317, w6318, w6319, w6320, w6321, w6322, w6323, w6324, w6325, w6326, w6327, w6328, w6329, w6330, w6331, w6332, w6333, w6334, w6335, w6336, w6337, w6338, w6339, w6340, w6341, w6342, w6343, w6344, w6345, w6346, w6347, w6348, w6349, w6350, w6351, w6352, w6353, w6354, w6355, w6356, w6357, w6358, w6359, w6360, w6361, w6362, w6363, w6364, w6365, w6366, w6367, w6368, w6369, w6370, w6371, w6372, w6373, w6374, w6375, w6376, w6377, w6378, w6379, w6380, w6381, w6382, w6383, w6384, w6385, w6386, w6387, w6388, w6389, w6390, w6391, w6392, w6393, w6394, w6395, w6396, w6397, w6398, w6399, w6400, w6401, w6402, w6403, w6404, w6405, w6406, w6407, w6408, w6409, w6410, w6411, w6412, w6413, w6414, w6415, w6416, w6417, w6418, w6419, w6420, w6421, w6422, w6423, w6424, w6425, w6426, w6427, w6428, w6429, w6430, w6431, w6432, w6433, w6434, w6435, w6436, w6437, w6438, w6439, w6440, w6441, w6442, w6443, w6444, w6445, w6446, w6447, w6448, w6449, w6450, w6451, w6452, w6453, w6454, w6455, w6456, w6457, w6458, w6459, w6460, w6461, w6462, w6463, w6464, w6465, w6466, w6467, w6468, w6469, w6470, w6471, w6472, w6473, w6474, w6475, w6476, w6477, w6478, w6479, w6480, w6481, w6482, w6483, w6484, w6485, w6486, w6487, w6488, w6489, w6490, w6491, w6492, w6493, w6494, w6495, w6496, w6497, w6498, w6499, w6500, w6501, w6502, w6503, w6504, w6505, w6506, w6507, w6508, w6509, w6510, w6511, w6512, w6513, w6514, w6515, w6516, w6517, w6518, w6519, w6520, w6521, w6522, w6523, w6524, w6525, w6526, w6527, w6528, w6529, w6530, w6531, w6532, w6533, w6534, w6535, w6536, w6537, w6538, w6539, w6540, w6541, w6542, w6543, w6544, w6545, w6546, w6547, w6548, w6549, w6550, w6551, w6552, w6553, w6554, w6555, w6556, w6557, w6558, w6559, w6560, w6561, w6562, w6563, w6564, w6565, w6566, w6567, w6568, w6569, w6570, w6571, w6572, w6573, w6574, w6575, w6576, w6577, w6578, w6579, w6580, w6581, w6582, w6583, w6584, w6585, w6586, w6587, w6588, w6589, w6590, w6591, w6592, w6593, w6594, w6595, w6596, w6597, w6598, w6599, w6600, w6601, w6602, w6603, w6604, w6605, w6606, w6607, w6608, w6609, w6610, w6611, w6612, w6613, w6614, w6615, w6616, w6617, w6618, w6619, w6620, w6621, w6622, w6623, w6624, w6625, w6626, w6627, w6628, w6629, w6630, w6631, w6632, w6633, w6634, w6635, w6636, w6637, w6638, w6639, w6640, w6641, w6642, w6643, w6644, w6645, w6646, w6647, w6648, w6649, w6650, w6651, w6652, w6653, w6654, w6655, w6656, w6657, w6658, w6659, w6660, w6661, w6662, w6663, w6664, w6665, w6666, w6667, w6668, w6669, w6670, w6671, w6672, w6673, w6674, w6675, w6676, w6677, w6678, w6679, w6680, w6681, w6682, w6683, w6684, w6685, w6686, w6687, w6688, w6689, w6690, w6691, w6692, w6693, w6694, w6695, w6696, w6697, w6698, w6699, w6700, w6701, w6702, w6703, w6704, w6705, w6706, w6707, w6708, w6709, w6710, w6711, w6712, w6713, w6714, w6715, w6716, w6717, w6718, w6719, w6720, w6721, w6722, w6723, w6724, w6725, w6726, w6727, w6728, w6729, w6730, w6731, w6732, w6733, w6734, w6735, w6736, w6737, w6738, w6739, w6740, w6741, w6742, w6743, w6744, w6745, w6746, w6747, w6748, w6749, w6750, w6751, w6752, w6753, w6754, w6755, w6756, w6757, w6758, w6759, w6760, w6761, w6762, w6763, w6764, w6765, w6766, w6767, w6768, w6769, w6770, w6771, w6772, w6773, w6774, w6775, w6776, w6777, w6778, w6779, w6780, w6781, w6782, w6783, w6784, w6785, w6786, w6787, w6788, w6789, w6790, w6791, w6792, w6793, w6794, w6795, w6796, w6797, w6798, w6799, w6800, w6801, w6802, w6803, w6804, w6805, w6806, w6807, w6808, w6809, w6810, w6811, w6812, w6813, w6814, w6815, w6816, w6817, w6818, w6819, w6820, w6821, w6822, w6823, w6824, w6825, w6826, w6827, w6828, w6829, w6830, w6831, w6832, w6833, w6834, w6835, w6836, w6837, w6838, w6839, w6840, w6841, w6842, w6843, w6844, w6845, w6846, w6847, w6848, w6849, w6850, w6851, w6852, w6853, w6854, w6855, w6856, w6857, w6858, w6859, w6860, w6861, w6862, w6863, w6864, w6865, w6866, w6867, w6868, w6869, w6870, w6871, w6872, w6873, w6874, w6875, w6876, w6877, w6878, w6879, w6880, w6881, w6882, w6883, w6884, w6885, w6886, w6887, w6888, w6889, w6890, w6891, w6892, w6893, w6894, w6895, w6896, w6897, w6898, w6899, w6900, w6901, w6902, w6903, w6904, w6905, w6906, w6907, w6908, w6909, w6910, w6911, w6912, w6913, w6914, w6915, w6916, w6917, w6918, w6919, w6920, w6921, w6922, w6923, w6924, w6925, w6926, w6927, w6928, w6929, w6930, w6931, w6932, w6933, w6934, w6935, w6936, w6937, w6938, w6939, w6940, w6941, w6942, w6943, w6944, w6945, w6946, w6947, w6948, w6949, w6950, w6951, w6952, w6953, w6954, w6955, w6956, w6957, w6958, w6959, w6960, w6961, w6962, w6963, w6964, w6965, w6966, w6967, w6968, w6969, w6970, w6971, w6972, w6973, w6974, w6975, w6976, w6977, w6978, w6979, w6980, w6981, w6982, w6983, w6984, w6985, w6986, w6987, w6988, w6989, w6990, w6991, w6992, w6993, w6994, w6995, w6996, w6997, w6998, w6999, w7000, w7001, w7002, w7003, w7004, w7005, w7006, w7007, w7008, w7009, w7010, w7011, w7012, w7013, w7014, w7015, w7016, w7017, w7018, w7019, w7020, w7021, w7022, w7023, w7024, w7025, w7026, w7027, w7028, w7029, w7030, w7031, w7032, w7033, w7034, w7035, w7036, w7037, w7038, w7039, w7040, w7041, w7042, w7043, w7044, w7045, w7046, w7047, w7048, w7049, w7050, w7051, w7052, w7053, w7054, w7055, w7056, w7057, w7058, w7059, w7060, w7061, w7062, w7063, w7064, w7065, w7066, w7067, w7068, w7069, w7070, w7071, w7072, w7073, w7074, w7075, w7076, w7077, w7078, w7079, w7080, w7081, w7082, w7083, w7084, w7085, w7086, w7087, w7088, w7089, w7090, w7091, w7092, w7093, w7094, w7095, w7096, w7097, w7098, w7099, w7100, w7101, w7102, w7103, w7104, w7105, w7106, w7107, w7108, w7109, w7110, w7111, w7112, w7113, w7114, w7115, w7116, w7117, w7118, w7119, w7120, w7121, w7122, w7123, w7124, w7125, w7126, w7127, w7128, w7129, w7130, w7131, w7132, w7133, w7134, w7135, w7136, w7137, w7138, w7139, w7140, w7141, w7142, w7143, w7144, w7145, w7146, w7147, w7148, w7149, w7150, w7151, w7152, w7153, w7154, w7155, w7156, w7157, w7158, w7159, w7160, w7161, w7162, w7163, w7164, w7165, w7166, w7167, w7168, w7169, w7170, w7171, w7172, w7173, w7174, w7175, w7176, w7177, w7178, w7179, w7180, w7181, w7182, w7183, w7184, w7185, w7186, w7187, w7188, w7189, w7190, w7191, w7192, w7193, w7194, w7195, w7196, w7197, w7198, w7199, w7200, w7201, w7202, w7203, w7204, w7205, w7206, w7207, w7208, w7209, w7210, w7211, w7212, w7213, w7214, w7215, w7216, w7217, w7218, w7219, w7220, w7221, w7222, w7223, w7224, w7225, w7226, w7227, w7228, w7229, w7230, w7231, w7232, w7233, w7234, w7235, w7236, w7237, w7238, w7239, w7240, w7241, w7242, w7243, w7244, w7245, w7246, w7247, w7248, w7249, w7250, w7251, w7252, w7253, w7254, w7255, w7256, w7257, w7258, w7259, w7260, w7261, w7262, w7263, w7264, w7265, w7266, w7267, w7268, w7269, w7270, w7271, w7272, w7273, w7274, w7275, w7276, w7277, w7278, w7279, w7280, w7281, w7282, w7283, w7284, w7285, w7286, w7287, w7288, w7289, w7290, w7291, w7292, w7293, w7294, w7295, w7296, w7297, w7298, w7299, w7300, w7301, w7302, w7303, w7304, w7305, w7306, w7307, w7308, w7309, w7310, w7311, w7312, w7313, w7314, w7315, w7316, w7317, w7318, w7319, w7320, w7321, w7322, w7323, w7324, w7325, w7326, w7327, w7328, w7329, w7330, w7331, w7332, w7333, w7334, w7335, w7336, w7337, w7338, w7339, w7340, w7341, w7342, w7343, w7344, w7345, w7346, w7347, w7348, w7349, w7350, w7351, w7352, w7353, w7354, w7355, w7356, w7357, w7358, w7359, w7360, w7361, w7362, w7363, w7364, w7365, w7366, w7367, w7368, w7369, w7370, w7371, w7372, w7373, w7374, w7375, w7376, w7377, w7378, w7379, w7380, w7381, w7382, w7383, w7384, w7385, w7386, w7387, w7388, w7389, w7390, w7391, w7392, w7393, w7394, w7395, w7396, w7397, w7398, w7399, w7400, w7401, w7402, w7403, w7404, w7405, w7406, w7407, w7408, w7409, w7410, w7411, w7412, w7413, w7414, w7415, w7416, w7417, w7418, w7419, w7420, w7421, w7422, w7423, w7424, w7425, w7426, w7427, w7428, w7429, w7430, w7431, w7432, w7433, w7434, w7435, w7436, w7437, w7438, w7439, w7440, w7441, w7442, w7443, w7444, w7445, w7446, w7447, w7448, w7449, w7450, w7451, w7452, w7453, w7454, w7455, w7456, w7457, w7458, w7459, w7460, w7461, w7462, w7463, w7464, w7465, w7466, w7467, w7468, w7469, w7470, w7471, w7472, w7473, w7474, w7475, w7476, w7477, w7478, w7479, w7480, w7481, w7482, w7483, w7484, w7485, w7486, w7487, w7488, w7489, w7490, w7491, w7492, w7493, w7494, w7495, w7496, w7497, w7498, w7499, w7500, w7501, w7502, w7503, w7504, w7505, w7506, w7507, w7508, w7509, w7510, w7511, w7512, w7513, w7514, w7515, w7516, w7517, w7518, w7519, w7520, w7521, w7522, w7523, w7524, w7525, w7526, w7527, w7528, w7529, w7530, w7531, w7532, w7533, w7534, w7535, w7536, w7537, w7538, w7539, w7540, w7541, w7542, w7543, w7544, w7545, w7546, w7547, w7548, w7549, w7550, w7551, w7552, w7553, w7554, w7555, w7556, w7557, w7558, w7559, w7560, w7561, w7562, w7563, w7564, w7565, w7566, w7567, w7568, w7569, w7570, w7571, w7572, w7573, w7574, w7575, w7576, w7577, w7578, w7579, w7580, w7581, w7582, w7583, w7584, w7585, w7586, w7587, w7588, w7589, w7590, w7591, w7592, w7593, w7594, w7595, w7596, w7597, w7598, w7599, w7600, w7601, w7602, w7603, w7604, w7605, w7606, w7607, w7608, w7609, w7610, w7611, w7612, w7613, w7614, w7615, w7616, w7617, w7618, w7619, w7620, w7621, w7622, w7623, w7624, w7625, w7626, w7627, w7628, w7629, w7630, w7631, w7632, w7633, w7634, w7635, w7636, w7637, w7638, w7639, w7640, w7641, w7642, w7643, w7644, w7645, w7646, w7647, w7648, w7649, w7650, w7651, w7652, w7653, w7654, w7655, w7656, w7657, w7658, w7659, w7660, w7661, w7662, w7663, w7664, w7665, w7666, w7667, w7668, w7669, w7670, w7671, w7672, w7673, w7674, w7675, w7676, w7677, w7678, w7679, w7680, w7681, w7682, w7683, w7684, w7685, w7686, w7687, w7688, w7689, w7690, w7691, w7692, w7693, w7694, w7695, w7696, w7697, w7698, w7699, w7700, w7701, w7702, w7703, w7704, w7705, w7706, w7707, w7708, w7709, w7710, w7711, w7712, w7713, w7714, w7715, w7716, w7717, w7718, w7719, w7720, w7721, w7722, w7723, w7724, w7725, w7726, w7727, w7728, w7729, w7730, w7731, w7732, w7733, w7734, w7735, w7736, w7737, w7738, w7739, w7740, w7741, w7742, w7743, w7744, w7745, w7746, w7747, w7748, w7749, w7750, w7751, w7752, w7753, w7754, w7755, w7756, w7757, w7758, w7759, w7760, w7761, w7762, w7763, w7764, w7765, w7766, w7767, w7768, w7769, w7770, w7771, w7772, w7773, w7774, w7775, w7776, w7777, w7778, w7779, w7780, w7781, w7782, w7783, w7784, w7785, w7786, w7787, w7788, w7789, w7790, w7791, w7792, w7793, w7794, w7795, w7796, w7797, w7798, w7799, w7800, w7801, w7802, w7803, w7804, w7805, w7806, w7807, w7808, w7809, w7810, w7811, w7812, w7813, w7814, w7815, w7816, w7817, w7818, w7819, w7820, w7821, w7822, w7823, w7824, w7825, w7826, w7827, w7828, w7829, w7830, w7831, w7832, w7833, w7834, w7835, w7836, w7837, w7838, w7839, w7840, w7841, w7842, w7843, w7844, w7845, w7846, w7847, w7848, w7849, w7850, w7851, w7852, w7853, w7854, w7855, w7856, w7857, w7858, w7859, w7860, w7861, w7862, w7863, w7864, w7865, w7866, w7867, w7868, w7869, w7870, w7871, w7872, w7873, w7874, w7875, w7876, w7877, w7878, w7879, w7880, w7881, w7882, w7883, w7884, w7885, w7886, w7887, w7888, w7889, w7890, w7891, w7892, w7893, w7894, w7895, w7896, w7897, w7898, w7899, w7900, w7901, w7902, w7903, w7904, w7905, w7906, w7907, w7908, w7909, w7910, w7911, w7912, w7913, w7914, w7915, w7916, w7917, w7918, w7919, w7920, w7921, w7922, w7923, w7924, w7925, w7926, w7927, w7928, w7929, w7930, w7931, w7932, w7933, w7934, w7935, w7936, w7937, w7938, w7939, w7940, w7941, w7942, w7943, w7944, w7945, w7946, w7947, w7948, w7949, w7950, w7951, w7952, w7953, w7954, w7955, w7956, w7957, w7958, w7959, w7960, w7961, w7962, w7963, w7964, w7965, w7966, w7967, w7968, w7969, w7970, w7971, w7972, w7973, w7974, w7975, w7976, w7977, w7978, w7979, w7980, w7981, w7982, w7983, w7984, w7985, w7986, w7987, w7988, w7989, w7990, w7991, w7992, w7993, w7994, w7995, w7996, w7997, w7998, w7999, w8000, w8001, w8002, w8003, w8004, w8005, w8006, w8007, w8008, w8009, w8010, w8011, w8012, w8013, w8014, w8015, w8016, w8017, w8018, w8019, w8020, w8021, w8022, w8023, w8024, w8025, w8026, w8027, w8028, w8029, w8030, w8031, w8032, w8033, w8034, w8035, w8036, w8037, w8038, w8039, w8040, w8041, w8042, w8043, w8044, w8045, w8046, w8047, w8048, w8049, w8050, w8051, w8052, w8053, w8054, w8055, w8056, w8057, w8058, w8059, w8060, w8061, w8062, w8063, w8064, w8065, w8066, w8067, w8068, w8069, w8070, w8071, w8072, w8073, w8074, w8075, w8076, w8077, w8078, w8079, w8080, w8081, w8082, w8083, w8084, w8085, w8086, w8087, w8088, w8089, w8090, w8091, w8092, w8093, w8094, w8095, w8096, w8097, w8098, w8099, w8100, w8101, w8102, w8103, w8104, w8105, w8106, w8107, w8108, w8109, w8110, w8111, w8112, w8113, w8114, w8115, w8116, w8117, w8118, w8119, w8120, w8121, w8122, w8123, w8124, w8125, w8126, w8127, w8128, w8129, w8130, w8131, w8132, w8133, w8134, w8135, w8136, w8137, w8138, w8139, w8140, w8141, w8142, w8143, w8144, w8145, w8146, w8147, w8148, w8149, w8150, w8151, w8152, w8153, w8154, w8155, w8156, w8157, w8158, w8159, w8160, w8161, w8162, w8163, w8164, w8165, w8166, w8167, w8168, w8169, w8170, w8171, w8172, w8173, w8174, w8175, w8176, w8177, w8178, w8179, w8180, w8181, w8182, w8183, w8184, w8185, w8186, w8187, w8188, w8189, w8190, w8191, w8192, w8193, w8194, w8195, w8196, w8197, w8198, w8199, w8200, w8201, w8202, w8203, w8204, w8205, w8206, w8207, w8208, w8209, w8210, w8211, w8212, w8213, w8214, w8215, w8216, w8217, w8218, w8219, w8220, w8221, w8222, w8223, w8224, w8225, w8226, w8227, w8228, w8229, w8230, w8231, w8232, w8233, w8234, w8235, w8236, w8237, w8238, w8239, w8240, w8241, w8242, w8243, w8244, w8245, w8246, w8247, w8248, w8249, w8250, w8251, w8252, w8253, w8254, w8255, w8256, w8257, w8258, w8259, w8260, w8261, w8262, w8263, w8264, w8265, w8266, w8267, w8268, w8269, w8270, w8271, w8272, w8273, w8274, w8275, w8276, w8277, w8278, w8279, w8280, w8281, w8282, w8283, w8284, w8285, w8286, w8287, w8288, w8289, w8290, w8291, w8292, w8293, w8294, w8295, w8296, w8297, w8298, w8299, w8300, w8301, w8302, w8303, w8304, w8305, w8306, w8307, w8308, w8309, w8310, w8311, w8312, w8313, w8314, w8315, w8316, w8317, w8318, w8319, w8320, w8321, w8322, w8323, w8324, w8325, w8326, w8327, w8328, w8329, w8330, w8331, w8332, w8333, w8334, w8335, w8336, w8337, w8338, w8339, w8340, w8341, w8342, w8343, w8344, w8345, w8346, w8347, w8348, w8349, w8350, w8351, w8352, w8353, w8354, w8355, w8356, w8357, w8358, w8359, w8360, w8361, w8362, w8363, w8364, w8365, w8366, w8367, w8368, w8369, w8370, w8371, w8372, w8373, w8374, w8375, w8376, w8377, w8378, w8379, w8380, w8381, w8382, w8383, w8384, w8385, w8386, w8387, w8388, w8389, w8390, w8391, w8392, w8393, w8394, w8395, w8396, w8397, w8398, w8399, w8400, w8401, w8402, w8403, w8404, w8405, w8406, w8407, w8408, w8409, w8410, w8411, w8412, w8413, w8414, w8415, w8416, w8417, w8418, w8419, w8420, w8421, w8422, w8423, w8424, w8425, w8426, w8427, w8428, w8429, w8430, w8431, w8432, w8433, w8434, w8435, w8436, w8437, w8438, w8439, w8440, w8441, w8442, w8443, w8444, w8445, w8446, w8447, w8448, w8449, w8450, w8451, w8452, w8453, w8454, w8455, w8456, w8457, w8458, w8459, w8460, w8461, w8462, w8463, w8464, w8465, w8466, w8467, w8468, w8469, w8470, w8471, w8472, w8473, w8474, w8475, w8476, w8477, w8478, w8479, w8480, w8481, w8482, w8483, w8484, w8485, w8486, w8487, w8488, w8489, w8490, w8491, w8492, w8493, w8494, w8495, w8496, w8497, w8498, w8499, w8500, w8501, w8502, w8503, w8504, w8505, w8506, w8507, w8508, w8509, w8510, w8511, w8512, w8513, w8514, w8515, w8516, w8517, w8518, w8519, w8520, w8521, w8522, w8523, w8524, w8525, w8526, w8527, w8528, w8529, w8530, w8531, w8532, w8533, w8534, w8535, w8536, w8537, w8538, w8539, w8540, w8541, w8542, w8543, w8544, w8545, w8546, w8547, w8548, w8549, w8550, w8551, w8552, w8553, w8554, w8555, w8556, w8557, w8558, w8559, w8560, w8561, w8562, w8563, w8564, w8565, w8566, w8567, w8568, w8569, w8570, w8571, w8572, w8573, w8574, w8575, w8576, w8577, w8578, w8579, w8580, w8581, w8582, w8583, w8584, w8585, w8586, w8587, w8588, w8589, w8590, w8591, w8592, w8593, w8594, w8595, w8596, w8597, w8598, w8599, w8600, w8601, w8602, w8603, w8604, w8605, w8606, w8607, w8608, w8609, w8610, w8611, w8612, w8613, w8614, w8615, w8616, w8617, w8618, w8619, w8620, w8621, w8622, w8623, w8624, w8625, w8626, w8627, w8628, w8629, w8630, w8631, w8632, w8633, w8634, w8635, w8636, w8637, w8638, w8639, w8640, w8641, w8642, w8643, w8644, w8645, w8646, w8647, w8648, w8649, w8650, w8651, w8652, w8653, w8654, w8655, w8656, w8657, w8658, w8659, w8660, w8661, w8662, w8663, w8664, w8665, w8666, w8667, w8668, w8669, w8670, w8671, w8672, w8673, w8674, w8675, w8676, w8677, w8678, w8679, w8680, w8681, w8682, w8683, w8684, w8685, w8686, w8687, w8688, w8689, w8690, w8691, w8692, w8693, w8694, w8695, w8696, w8697, w8698, w8699, w8700, w8701, w8702, w8703, w8704, w8705, w8706, w8707, w8708, w8709, w8710, w8711, w8712, w8713, w8714, w8715, w8716, w8717, w8718, w8719, w8720, w8721, w8722, w8723, w8724, w8725, w8726, w8727, w8728, w8729, w8730, w8731, w8732, w8733, w8734, w8735, w8736, w8737, w8738, w8739, w8740, w8741, w8742, w8743, w8744, w8745, w8746, w8747, w8748, w8749, w8750, w8751, w8752, w8753, w8754, w8755, w8756, w8757, w8758, w8759, w8760, w8761, w8762, w8763, w8764, w8765, w8766, w8767, w8768, w8769, w8770, w8771, w8772, w8773, w8774, w8775, w8776, w8777, w8778, w8779, w8780, w8781, w8782, w8783, w8784, w8785, w8786, w8787, w8788, w8789, w8790, w8791, w8792, w8793, w8794, w8795, w8796, w8797, w8798, w8799, w8800, w8801, w8802, w8803, w8804, w8805, w8806, w8807, w8808, w8809, w8810, w8811, w8812, w8813, w8814, w8815, w8816, w8817, w8818, w8819, w8820, w8821, w8822, w8823, w8824, w8825, w8826, w8827, w8828, w8829, w8830, w8831, w8832, w8833, w8834, w8835, w8836, w8837, w8838, w8839, w8840, w8841, w8842, w8843, w8844, w8845, w8846, w8847, w8848, w8849, w8850, w8851, w8852, w8853, w8854, w8855, w8856, w8857, w8858, w8859, w8860, w8861, w8862, w8863, w8864, w8865, w8866, w8867, w8868, w8869, w8870, w8871, w8872, w8873, w8874, w8875, w8876, w8877, w8878, w8879, w8880, w8881, w8882, w8883, w8884, w8885, w8886, w8887, w8888, w8889, w8890, w8891, w8892, w8893, w8894, w8895, w8896, w8897, w8898, w8899, w8900, w8901, w8902, w8903, w8904, w8905, w8906, w8907, w8908, w8909, w8910, w8911, w8912, w8913, w8914, w8915, w8916, w8917, w8918, w8919, w8920, w8921, w8922, w8923, w8924, w8925, w8926, w8927, w8928, w8929, w8930, w8931, w8932, w8933, w8934, w8935, w8936, w8937, w8938, w8939, w8940, w8941, w8942, w8943, w8944, w8945, w8946, w8947, w8948, w8949, w8950, w8951, w8952, w8953, w8954, w8955, w8956, w8957, w8958, w8959, w8960, w8961, w8962, w8963, w8964, w8965, w8966, w8967, w8968, w8969, w8970, w8971, w8972, w8973, w8974, w8975, w8976, w8977, w8978, w8979, w8980, w8981, w8982, w8983, w8984, w8985, w8986, w8987, w8988, w8989, w8990, w8991, w8992, w8993, w8994, w8995, w8996, w8997, w8998, w8999, w9000, w9001, w9002, w9003, w9004, w9005, w9006, w9007, w9008, w9009, w9010, w9011, w9012, w9013, w9014, w9015, w9016, w9017, w9018, w9019, w9020, w9021, w9022, w9023, w9024, w9025, w9026, w9027, w9028, w9029, w9030, w9031, w9032, w9033, w9034, w9035, w9036, w9037, w9038, w9039, w9040, w9041, w9042, w9043, w9044, w9045, w9046, w9047, w9048, w9049, w9050, w9051, w9052, w9053, w9054, w9055, w9056, w9057, w9058, w9059, w9060, w9061, w9062, w9063, w9064, w9065, w9066, w9067, w9068, w9069, w9070, w9071, w9072, w9073, w9074, w9075, w9076, w9077, w9078, w9079, w9080, w9081, w9082, w9083, w9084, w9085, w9086, w9087, w9088, w9089, w9090, w9091, w9092, w9093, w9094, w9095, w9096, w9097, w9098, w9099, w9100, w9101, w9102, w9103, w9104, w9105, w9106, w9107, w9108, w9109, w9110, w9111, w9112, w9113, w9114, w9115, w9116, w9117, w9118, w9119, w9120, w9121, w9122, w9123, w9124, w9125, w9126, w9127, w9128, w9129, w9130, w9131, w9132, w9133, w9134, w9135, w9136, w9137, w9138, w9139, w9140, w9141, w9142, w9143, w9144, w9145, w9146, w9147, w9148, w9149, w9150, w9151, w9152, w9153, w9154, w9155, w9156, w9157, w9158, w9159, w9160, w9161, w9162, w9163, w9164, w9165, w9166, w9167, w9168, w9169, w9170, w9171, w9172, w9173, w9174, w9175, w9176, w9177, w9178, w9179, w9180, w9181, w9182, w9183, w9184, w9185, w9186, w9187, w9188, w9189, w9190, w9191, w9192, w9193, w9194, w9195, w9196, w9197, w9198, w9199, w9200, w9201, w9202, w9203, w9204, w9205, w9206, w9207, w9208, w9209, w9210, w9211, w9212, w9213, w9214, w9215, w9216, w9217, w9218, w9219, w9220, w9221, w9222, w9223, w9224, w9225, w9226, w9227, w9228, w9229, w9230, w9231, w9232, w9233, w9234, w9235, w9236, w9237, w9238, w9239, w9240, w9241, w9242, w9243, w9244, w9245, w9246, w9247, w9248, w9249, w9250, w9251, w9252, w9253, w9254, w9255, w9256, w9257, w9258, w9259, w9260, w9261, w9262, w9263, w9264, w9265, w9266, w9267, w9268, w9269, w9270, w9271, w9272, w9273, w9274, w9275, w9276, w9277, w9278, w9279, w9280, w9281, w9282, w9283, w9284, w9285, w9286, w9287, w9288, w9289, w9290, w9291, w9292, w9293, w9294, w9295, w9296, w9297, w9298, w9299, w9300, w9301, w9302, w9303, w9304, w9305, w9306, w9307, w9308, w9309, w9310, w9311, w9312, w9313, w9314, w9315, w9316, w9317, w9318, w9319, w9320, w9321, w9322, w9323, w9324, w9325, w9326, w9327, w9328, w9329, w9330, w9331, w9332, w9333, w9334, w9335, w9336, w9337, w9338, w9339, w9340, w9341, w9342, w9343, w9344, w9345, w9346, w9347, w9348, w9349, w9350, w9351, w9352, w9353, w9354, w9355, w9356, w9357, w9358, w9359, w9360, w9361, w9362, w9363, w9364, w9365, w9366, w9367, w9368, w9369, w9370, w9371, w9372, w9373, w9374, w9375, w9376, w9377, w9378, w9379, w9380, w9381, w9382, w9383, w9384, w9385, w9386, w9387, w9388, w9389, w9390, w9391, w9392, w9393, w9394, w9395, w9396, w9397, w9398, w9399, w9400, w9401, w9402, w9403, w9404, w9405, w9406, w9407, w9408, w9409, w9410, w9411, w9412, w9413, w9414, w9415, w9416, w9417, w9418, w9419, w9420, w9421, w9422, w9423, w9424, w9425, w9426, w9427, w9428, w9429, w9430, w9431, w9432, w9433, w9434, w9435, w9436, w9437, w9438, w9439, w9440, w9441, w9442, w9443, w9444, w9445, w9446, w9447, w9448, w9449, w9450, w9451, w9452, w9453, w9454, w9455, w9456, w9457, w9458, w9459, w9460, w9461, w9462, w9463, w9464, w9465, w9466, w9467, w9468, w9469, w9470, w9471, w9472, w9473, w9474, w9475, w9476, w9477, w9478, w9479, w9480, w9481, w9482, w9483, w9484, w9485, w9486, w9487, w9488, w9489, w9490, w9491, w9492, w9493, w9494, w9495, w9496, w9497, w9498, w9499, w9500, w9501, w9502, w9503, w9504, w9505, w9506, w9507, w9508, w9509, w9510, w9511, w9512, w9513, w9514, w9515, w9516, w9517, w9518, w9519, w9520, w9521, w9522, w9523, w9524, w9525, w9526, w9527, w9528, w9529, w9530, w9531, w9532, w9533, w9534, w9535, w9536, w9537, w9538, w9539, w9540, w9541, w9542, w9543, w9544, w9545, w9546, w9547, w9548, w9549, w9550, w9551, w9552, w9553, w9554, w9555, w9556, w9557, w9558, w9559, w9560, w9561, w9562, w9563, w9564, w9565, w9566, w9567, w9568, w9569, w9570, w9571, w9572, w9573, w9574, w9575, w9576, w9577, w9578, w9579, w9580, w9581, w9582, w9583, w9584, w9585, w9586, w9587, w9588, w9589, w9590, w9591, w9592, w9593, w9594, w9595, w9596, w9597, w9598, w9599, w9600, w9601, w9602, w9603, w9604, w9605, w9606, w9607, w9608, w9609, w9610, w9611, w9612, w9613, w9614, w9615, w9616, w9617, w9618, w9619, w9620, w9621, w9622, w9623, w9624, w9625, w9626, w9627, w9628, w9629, w9630, w9631, w9632, w9633, w9634, w9635, w9636, w9637, w9638, w9639, w9640, w9641, w9642, w9643, w9644, w9645, w9646, w9647, w9648, w9649, w9650, w9651, w9652, w9653, w9654, w9655, w9656, w9657, w9658, w9659, w9660, w9661, w9662, w9663, w9664, w9665, w9666, w9667, w9668, w9669, w9670, w9671, w9672, w9673, w9674, w9675, w9676, w9677, w9678, w9679, w9680, w9681, w9682, w9683, w9684, w9685, w9686, w9687, w9688, w9689, w9690, w9691, w9692, w9693, w9694, w9695, w9696, w9697, w9698, w9699, w9700, w9701, w9702, w9703, w9704, w9705, w9706, w9707, w9708, w9709, w9710, w9711, w9712, w9713, w9714, w9715, w9716, w9717, w9718, w9719, w9720, w9721, w9722, w9723, w9724, w9725, w9726, w9727, w9728, w9729, w9730, w9731, w9732, w9733, w9734, w9735, w9736, w9737, w9738, w9739, w9740, w9741, w9742, w9743, w9744, w9745, w9746, w9747, w9748, w9749, w9750, w9751, w9752, w9753, w9754, w9755, w9756, w9757, w9758, w9759, w9760, w9761, w9762, w9763, w9764, w9765, w9766, w9767, w9768, w9769, w9770, w9771, w9772, w9773, w9774, w9775, w9776, w9777, w9778, w9779, w9780, w9781, w9782, w9783, w9784, w9785, w9786, w9787, w9788, w9789, w9790, w9791, w9792, w9793, w9794, w9795, w9796, w9797, w9798, w9799, w9800, w9801, w9802, w9803, w9804, w9805, w9806, w9807, w9808, w9809, w9810, w9811, w9812, w9813, w9814, w9815, w9816, w9817, w9818, w9819, w9820, w9821, w9822, w9823, w9824, w9825, w9826, w9827, w9828, w9829, w9830, w9831, w9832, w9833, w9834, w9835, w9836, w9837, w9838, w9839, w9840, w9841, w9842, w9843, w9844, w9845, w9846, w9847, w9848, w9849, w9850, w9851, w9852, w9853, w9854, w9855, w9856, w9857, w9858, w9859, w9860, w9861, w9862, w9863, w9864, w9865, w9866, w9867, w9868, w9869, w9870, w9871, w9872, w9873, w9874, w9875, w9876, w9877, w9878, w9879, w9880, w9881, w9882, w9883, w9884, w9885, w9886, w9887, w9888, w9889, w9890, w9891, w9892, w9893, w9894, w9895, w9896, w9897, w9898, w9899, w9900, w9901, w9902, w9903, w9904, w9905, w9906, w9907, w9908, w9909, w9910, w9911, w9912, w9913, w9914, w9915, w9916, w9917, w9918, w9919, w9920, w9921, w9922, w9923, w9924, w9925, w9926, w9927, w9928, w9929, w9930, w9931, w9932, w9933, w9934, w9935, w9936, w9937, w9938, w9939, w9940, w9941, w9942, w9943, w9944, w9945, w9946, w9947, w9948, w9949, w9950, w9951, w9952, w9953, w9954, w9955, w9956, w9957, w9958, w9959, w9960, w9961, w9962, w9963, w9964, w9965, w9966, w9967, w9968, w9969, w9970, w9971, w9972, w9973, w9974, w9975, w9976, w9977, w9978, w9979, w9980, w9981, w9982, w9983, w9984, w9985, w9986, w9987, w9988, w9989, w9990, w9991, w9992, w9993, w9994, w9995, w9996, w9997, w9998, w9999, w10000, w10001, w10002, w10003, w10004, w10005, w10006, w10007, w10008, w10009, w10010, w10011, w10012, w10013, w10014, w10015, w10016, w10017, w10018, w10019, w10020, w10021, w10022, w10023, w10024, w10025, w10026, w10027, w10028, w10029, w10030, w10031, w10032, w10033, w10034, w10035, w10036, w10037, w10038, w10039, w10040, w10041, w10042, w10043, w10044, w10045, w10046, w10047, w10048, w10049, w10050, w10051, w10052, w10053, w10054, w10055, w10056, w10057, w10058, w10059, w10060, w10061, w10062, w10063, w10064, w10065, w10066, w10067, w10068, w10069, w10070, w10071, w10072, w10073, w10074, w10075, w10076, w10077, w10078, w10079, w10080, w10081, w10082, w10083, w10084, w10085, w10086, w10087, w10088, w10089, w10090, w10091, w10092, w10093, w10094, w10095, w10096, w10097, w10098, w10099, w10100, w10101, w10102, w10103, w10104, w10105, w10106, w10107, w10108, w10109, w10110, w10111, w10112, w10113, w10114, w10115, w10116, w10117, w10118, w10119, w10120, w10121, w10122, w10123, w10124, w10125, w10126, w10127, w10128, w10129, w10130, w10131, w10132, w10133, w10134, w10135, w10136, w10137, w10138, w10139, w10140, w10141, w10142, w10143, w10144, w10145, w10146, w10147, w10148, w10149, w10150, w10151, w10152, w10153, w10154, w10155, w10156, w10157, w10158, w10159, w10160, w10161, w10162, w10163, w10164, w10165, w10166, w10167, w10168, w10169, w10170, w10171, w10172, w10173, w10174, w10175, w10176, w10177, w10178, w10179, w10180, w10181, w10182, w10183, w10184, w10185, w10186, w10187, w10188, w10189, w10190, w10191, w10192, w10193, w10194, w10195, w10196, w10197, w10198, w10199, w10200, w10201, w10202, w10203, w10204, w10205, w10206, w10207, w10208, w10209, w10210, w10211, w10212, w10213, w10214, w10215, w10216, w10217, w10218, w10219, w10220, w10221, w10222, w10223, w10224, w10225, w10226, w10227, w10228, w10229, w10230, w10231, w10232, w10233, w10234, w10235, w10236, w10237, w10238, w10239, w10240, w10241, w10242, w10243, w10244, w10245, w10246, w10247, w10248, w10249, w10250, w10251, w10252, w10253, w10254, w10255, w10256, w10257, w10258, w10259, w10260, w10261, w10262, w10263, w10264, w10265, w10266, w10267, w10268, w10269, w10270, w10271, w10272, w10273, w10274, w10275, w10276, w10277, w10278, w10279, w10280, w10281, w10282, w10283, w10284, w10285, w10286, w10287, w10288, w10289, w10290, w10291, w10292, w10293, w10294, w10295, w10296, w10297, w10298, w10299, w10300, w10301, w10302, w10303, w10304, w10305, w10306, w10307, w10308, w10309, w10310, w10311, w10312, w10313, w10314, w10315, w10316, w10317, w10318, w10319, w10320, w10321, w10322, w10323, w10324, w10325, w10326, w10327, w10328, w10329, w10330, w10331, w10332, w10333, w10334, w10335, w10336, w10337, w10338, w10339, w10340, w10341, w10342, w10343, w10344, w10345, w10346, w10347, w10348, w10349, w10350, w10351, w10352, w10353, w10354, w10355, w10356, w10357, w10358, w10359, w10360, w10361, w10362, w10363, w10364, w10365, w10366, w10367, w10368, w10369, w10370, w10371, w10372, w10373, w10374, w10375, w10376, w10377, w10378, w10379, w10380, w10381, w10382, w10383, w10384, w10385, w10386, w10387, w10388, w10389, w10390, w10391, w10392, w10393, w10394, w10395, w10396, w10397, w10398, w10399, w10400, w10401, w10402, w10403, w10404, w10405, w10406, w10407, w10408, w10409, w10410, w10411, w10412, w10413, w10414, w10415, w10416, w10417, w10418, w10419, w10420, w10421, w10422, w10423, w10424, w10425, w10426, w10427, w10428, w10429, w10430, w10431, w10432, w10433, w10434, w10435, w10436, w10437, w10438, w10439, w10440, w10441, w10442, w10443, w10444, w10445, w10446, w10447, w10448, w10449, w10450, w10451, w10452, w10453, w10454, w10455, w10456, w10457, w10458, w10459, w10460, w10461, w10462, w10463, w10464, w10465, w10466, w10467, w10468, w10469, w10470, w10471, w10472, w10473, w10474, w10475, w10476, w10477, w10478, w10479, w10480, w10481, w10482, w10483, w10484, w10485, w10486, w10487, w10488, w10489, w10490, w10491, w10492, w10493, w10494, w10495, w10496, w10497, w10498, w10499, w10500, w10501, w10502, w10503, w10504, w10505, w10506, w10507, w10508, w10509, w10510, w10511, w10512, w10513, w10514, w10515, w10516, w10517, w10518, w10519, w10520, w10521, w10522, w10523, w10524, w10525, w10526, w10527, w10528, w10529, w10530, w10531, w10532, w10533, w10534, w10535, w10536, w10537, w10538, w10539, w10540, w10541, w10542, w10543, w10544, w10545, w10546, w10547, w10548, w10549, w10550, w10551, w10552, w10553, w10554, w10555, w10556, w10557, w10558, w10559, w10560, w10561, w10562, w10563, w10564, w10565, w10566, w10567, w10568, w10569, w10570, w10571, w10572, w10573, w10574, w10575, w10576, w10577, w10578, w10579, w10580, w10581, w10582, w10583, w10584, w10585, w10586, w10587, w10588, w10589, w10590, w10591, w10592, w10593, w10594, w10595, w10596, w10597, w10598, w10599, w10600, w10601, w10602, w10603, w10604, w10605, w10606, w10607, w10608, w10609, w10610, w10611, w10612, w10613, w10614, w10615, w10616, w10617, w10618, w10619, w10620, w10621, w10622, w10623, w10624, w10625, w10626, w10627, w10628, w10629, w10630, w10631, w10632, w10633, w10634, w10635, w10636, w10637, w10638, w10639, w10640, w10641, w10642, w10643, w10644, w10645, w10646, w10647, w10648, w10649, w10650, w10651, w10652, w10653, w10654, w10655, w10656, w10657, w10658, w10659, w10660, w10661, w10662, w10663, w10664, w10665, w10666, w10667, w10668, w10669, w10670, w10671, w10672, w10673, w10674, w10675, w10676, w10677, w10678, w10679, w10680, w10681, w10682, w10683, w10684, w10685, w10686, w10687, w10688, w10689, w10690, w10691, w10692, w10693, w10694, w10695, w10696, w10697, w10698, w10699, w10700, w10701, w10702, w10703, w10704, w10705, w10706, w10707, w10708, w10709, w10710, w10711, w10712, w10713, w10714, w10715, w10716, w10717, w10718, w10719, w10720, w10721, w10722, w10723, w10724, w10725, w10726, w10727, w10728, w10729, w10730, w10731, w10732, w10733, w10734, w10735, w10736, w10737, w10738, w10739, w10740, w10741, w10742, w10743, w10744, w10745, w10746, w10747, w10748, w10749, w10750, w10751, w10752, w10753, w10754, w10755, w10756, w10757, w10758, w10759, w10760, w10761, w10762, w10763, w10764, w10765, w10766, w10767, w10768, w10769, w10770, w10771, w10772, w10773, w10774, w10775, w10776, w10777, w10778, w10779, w10780, w10781, w10782, w10783, w10784, w10785, w10786, w10787, w10788, w10789, w10790, w10791, w10792, w10793, w10794, w10795, w10796, w10797, w10798, w10799, w10800, w10801, w10802, w10803, w10804, w10805, w10806, w10807, w10808, w10809, w10810, w10811, w10812, w10813, w10814, w10815, w10816, w10817, w10818, w10819, w10820, w10821, w10822, w10823, w10824, w10825, w10826, w10827, w10828, w10829, w10830, w10831, w10832, w10833, w10834, w10835, w10836, w10837, w10838, w10839, w10840, w10841, w10842, w10843, w10844, w10845, w10846, w10847, w10848, w10849, w10850, w10851, w10852, w10853, w10854, w10855, w10856, w10857, w10858, w10859, w10860, w10861, w10862, w10863, w10864, w10865, w10866, w10867, w10868, w10869, w10870, w10871, w10872, w10873, w10874, w10875, w10876, w10877, w10878, w10879, w10880, w10881, w10882, w10883, w10884, w10885, w10886, w10887, w10888, w10889, w10890, w10891, w10892, w10893, w10894, w10895, w10896, w10897, w10898, w10899, w10900, w10901, w10902, w10903, w10904, w10905, w10906, w10907, w10908, w10909, w10910, w10911, w10912, w10913, w10914, w10915, w10916, w10917, w10918, w10919, w10920, w10921, w10922, w10923, w10924, w10925, w10926, w10927, w10928, w10929, w10930, w10931, w10932, w10933, w10934, w10935, w10936, w10937, w10938, w10939, w10940, w10941, w10942, w10943, w10944, w10945, w10946, w10947, w10948, w10949, w10950, w10951, w10952, w10953, w10954, w10955, w10956, w10957, w10958, w10959, w10960, w10961, w10962, w10963, w10964, w10965, w10966, w10967, w10968, w10969, w10970, w10971, w10972, w10973, w10974, w10975, w10976, w10977, w10978, w10979, w10980, w10981, w10982, w10983, w10984, w10985, w10986, w10987, w10988, w10989, w10990, w10991, w10992, w10993, w10994, w10995, w10996, w10997, w10998, w10999, w11000, w11001, w11002, w11003, w11004, w11005, w11006, w11007, w11008, w11009, w11010, w11011, w11012, w11013, w11014, w11015, w11016, w11017, w11018, w11019, w11020, w11021, w11022, w11023, w11024, w11025, w11026, w11027, w11028, w11029, w11030, w11031, w11032, w11033, w11034, w11035, w11036, w11037, w11038, w11039, w11040, w11041, w11042, w11043, w11044, w11045, w11046, w11047, w11048, w11049, w11050, w11051, w11052, w11053, w11054, w11055, w11056, w11057, w11058, w11059, w11060, w11061, w11062, w11063, w11064, w11065, w11066, w11067, w11068, w11069, w11070, w11071, w11072, w11073, w11074, w11075, w11076, w11077, w11078, w11079, w11080, w11081, w11082, w11083, w11084, w11085, w11086, w11087, w11088, w11089, w11090, w11091, w11092, w11093, w11094, w11095, w11096, w11097, w11098, w11099, w11100, w11101, w11102, w11103, w11104, w11105, w11106, w11107, w11108, w11109, w11110, w11111, w11112, w11113, w11114, w11115, w11116, w11117, w11118, w11119, w11120, w11121, w11122, w11123, w11124, w11125, w11126, w11127, w11128, w11129, w11130, w11131, w11132, w11133, w11134, w11135, w11136, w11137, w11138, w11139, w11140, w11141, w11142, w11143, w11144, w11145, w11146, w11147, w11148, w11149, w11150, w11151, w11152, w11153, w11154, w11155, w11156, w11157, w11158, w11159, w11160, w11161, w11162, w11163, w11164, w11165, w11166, w11167, w11168, w11169, w11170, w11171, w11172, w11173, w11174, w11175, w11176, w11177, w11178, w11179, w11180, w11181, w11182, w11183, w11184, w11185, w11186, w11187, w11188, w11189, w11190, w11191, w11192, w11193, w11194, w11195, w11196, w11197, w11198, w11199, w11200, w11201, w11202, w11203, w11204, w11205, w11206, w11207, w11208, w11209, w11210, w11211, w11212, w11213, w11214, w11215, w11216, w11217, w11218, w11219, w11220, w11221, w11222, w11223, w11224, w11225, w11226, w11227, w11228, w11229, w11230, w11231, w11232, w11233, w11234, w11235, w11236, w11237, w11238, w11239, w11240, w11241, w11242, w11243, w11244, w11245, w11246, w11247, w11248, w11249, w11250, w11251, w11252, w11253, w11254, w11255, w11256, w11257, w11258, w11259, w11260, w11261, w11262, w11263, w11264, w11265, w11266, w11267, w11268, w11269, w11270, w11271, w11272, w11273, w11274, w11275, w11276, w11277, w11278, w11279, w11280, w11281, w11282, w11283, w11284, w11285, w11286, w11287, w11288, w11289, w11290, w11291, w11292, w11293, w11294, w11295, w11296, w11297, w11298, w11299, w11300, w11301, w11302, w11303, w11304, w11305, w11306, w11307, w11308, w11309, w11310, w11311, w11312, w11313, w11314, w11315, w11316, w11317, w11318, w11319, w11320, w11321, w11322, w11323, w11324, w11325, w11326, w11327, w11328, w11329, w11330, w11331, w11332, w11333, w11334, w11335, w11336, w11337, w11338, w11339, w11340, w11341, w11342, w11343, w11344, w11345, w11346, w11347, w11348, w11349, w11350, w11351, w11352, w11353, w11354, w11355, w11356, w11357, w11358, w11359, w11360, w11361, w11362, w11363, w11364, w11365, w11366, w11367, w11368, w11369, w11370, w11371, w11372, w11373, w11374, w11375, w11376, w11377, w11378, w11379, w11380, w11381, w11382, w11383, w11384, w11385, w11386, w11387, w11388, w11389, w11390, w11391, w11392, w11393, w11394, w11395, w11396, w11397, w11398, w11399, w11400, w11401, w11402, w11403, w11404, w11405, w11406, w11407, w11408, w11409, w11410, w11411, w11412, w11413, w11414, w11415, w11416, w11417, w11418, w11419, w11420, w11421, w11422, w11423, w11424, w11425, w11426, w11427, w11428, w11429, w11430, w11431, w11432, w11433, w11434, w11435, w11436, w11437, w11438, w11439, w11440, w11441, w11442, w11443, w11444, w11445, w11446, w11447, w11448, w11449, w11450, w11451, w11452, w11453, w11454, w11455, w11456, w11457, w11458, w11459, w11460, w11461, w11462, w11463, w11464, w11465, w11466, w11467, w11468, w11469, w11470, w11471, w11472, w11473, w11474, w11475, w11476, w11477, w11478, w11479, w11480, w11481, w11482, w11483, w11484, w11485, w11486, w11487, w11488, w11489, w11490, w11491, w11492, w11493, w11494, w11495, w11496, w11497, w11498, w11499, w11500, w11501, w11502, w11503, w11504, w11505, w11506, w11507, w11508, w11509, w11510, w11511, w11512, w11513, w11514, w11515, w11516, w11517, w11518, w11519, w11520, w11521, w11522, w11523, w11524, w11525, w11526, w11527, w11528, w11529, w11530, w11531, w11532, w11533, w11534, w11535, w11536, w11537, w11538, w11539, w11540, w11541, w11542, w11543, w11544, w11545, w11546, w11547, w11548, w11549, w11550, w11551, w11552, w11553, w11554, w11555, w11556, w11557, w11558, w11559, w11560, w11561, w11562, w11563, w11564, w11565, w11566, w11567, w11568, w11569, w11570, w11571, w11572, w11573, w11574, w11575, w11576, w11577, w11578, w11579, w11580, w11581, w11582, w11583, w11584, w11585, w11586, w11587, w11588, w11589, w11590, w11591, w11592, w11593, w11594, w11595, w11596, w11597, w11598, w11599, w11600, w11601, w11602, w11603, w11604, w11605, w11606, w11607, w11608, w11609, w11610, w11611, w11612, w11613, w11614, w11615, w11616, w11617, w11618, w11619, w11620, w11621, w11622, w11623, w11624, w11625, w11626, w11627, w11628, w11629, w11630, w11631, w11632, w11633, w11634, w11635, w11636, w11637, w11638, w11639, w11640, w11641, w11642, w11643, w11644, w11645, w11646, w11647, w11648, w11649, w11650, w11651, w11652, w11653, w11654, w11655, w11656, w11657, w11658, w11659, w11660, w11661, w11662, w11663, w11664, w11665, w11666, w11667, w11668, w11669, w11670, w11671, w11672, w11673, w11674, w11675, w11676, w11677, w11678, w11679, w11680, w11681, w11682, w11683, w11684, w11685, w11686, w11687, w11688, w11689, w11690, w11691, w11692, w11693, w11694, w11695, w11696, w11697, w11698, w11699, w11700, w11701, w11702, w11703, w11704, w11705, w11706, w11707, w11708, w11709, w11710, w11711, w11712, w11713, w11714, w11715, w11716, w11717, w11718, w11719, w11720, w11721, w11722, w11723, w11724, w11725, w11726, w11727, w11728, w11729, w11730, w11731, w11732, w11733, w11734, w11735, w11736, w11737, w11738, w11739, w11740, w11741, w11742, w11743, w11744, w11745, w11746, w11747, w11748, w11749, w11750, w11751, w11752, w11753, w11754, w11755, w11756, w11757, w11758, w11759, w11760, w11761, w11762, w11763, w11764, w11765, w11766, w11767, w11768, w11769, w11770, w11771, w11772, w11773, w11774, w11775, w11776, w11777, w11778, w11779, w11780, w11781, w11782, w11783, w11784, w11785, w11786, w11787, w11788, w11789, w11790, w11791, w11792, w11793, w11794, w11795, w11796, w11797, w11798, w11799, w11800, w11801, w11802, w11803, w11804, w11805, w11806, w11807, w11808, w11809, w11810, w11811, w11812, w11813, w11814, w11815, w11816, w11817, w11818, w11819, w11820, w11821, w11822, w11823, w11824, w11825, w11826, w11827, w11828, w11829, w11830, w11831, w11832, w11833, w11834, w11835, w11836, w11837, w11838, w11839, w11840, w11841, w11842, w11843, w11844, w11845, w11846, w11847, w11848, w11849, w11850, w11851, w11852, w11853, w11854, w11855, w11856, w11857, w11858, w11859, w11860, w11861, w11862, w11863, w11864, w11865, w11866, w11867, w11868, w11869, w11870, w11871, w11872, w11873, w11874, w11875, w11876, w11877, w11878, w11879, w11880, w11881, w11882, w11883, w11884, w11885, w11886, w11887, w11888, w11889, w11890, w11891, w11892, w11893, w11894, w11895, w11896, w11897, w11898, w11899, w11900, w11901, w11902, w11903, w11904, w11905, w11906, w11907, w11908, w11909, w11910, w11911, w11912, w11913, w11914, w11915, w11916, w11917, w11918, w11919, w11920, w11921, w11922, w11923, w11924, w11925, w11926, w11927, w11928, w11929, w11930, w11931, w11932, w11933, w11934, w11935, w11936, w11937, w11938, w11939, w11940, w11941, w11942, w11943, w11944, w11945, w11946, w11947, w11948, w11949, w11950, w11951, w11952, w11953, w11954, w11955, w11956, w11957, w11958, w11959, w11960, w11961, w11962, w11963, w11964, w11965, w11966, w11967, w11968, w11969, w11970, w11971, w11972, w11973, w11974, w11975, w11976, w11977, w11978, w11979, w11980, w11981, w11982, w11983, w11984, w11985, w11986, w11987, w11988, w11989, w11990, w11991, w11992, w11993, w11994, w11995, w11996, w11997, w11998, w11999, w12000, w12001, w12002, w12003, w12004, w12005, w12006, w12007, w12008, w12009, w12010, w12011, w12012, w12013, w12014, w12015, w12016, w12017, w12018, w12019, w12020, w12021, w12022, w12023, w12024, w12025, w12026, w12027, w12028, w12029, w12030, w12031, w12032, w12033, w12034, w12035, w12036, w12037, w12038, w12039, w12040, w12041, w12042, w12043, w12044, w12045, w12046, w12047, w12048, w12049, w12050, w12051, w12052, w12053, w12054, w12055, w12056, w12057, w12058, w12059, w12060, w12061, w12062, w12063, w12064, w12065, w12066, w12067, w12068, w12069, w12070, w12071, w12072, w12073, w12074, w12075, w12076, w12077, w12078, w12079, w12080, w12081, w12082, w12083, w12084, w12085, w12086, w12087, w12088, w12089, w12090, w12091, w12092, w12093, w12094, w12095, w12096, w12097, w12098, w12099, w12100, w12101, w12102, w12103, w12104, w12105, w12106, w12107, w12108, w12109, w12110, w12111, w12112, w12113, w12114, w12115, w12116, w12117, w12118, w12119, w12120, w12121, w12122, w12123, w12124, w12125, w12126, w12127, w12128, w12129, w12130, w12131, w12132, w12133, w12134, w12135, w12136, w12137, w12138, w12139, w12140, w12141, w12142, w12143, w12144, w12145, w12146, w12147, w12148, w12149, w12150, w12151, w12152, w12153, w12154, w12155, w12156, w12157, w12158, w12159, w12160, w12161, w12162, w12163, w12164, w12165, w12166, w12167, w12168, w12169, w12170, w12171, w12172, w12173, w12174, w12175, w12176, w12177, w12178, w12179, w12180, w12181, w12182, w12183, w12184, w12185, w12186, w12187, w12188, w12189, w12190, w12191, w12192, w12193, w12194, w12195, w12196, w12197, w12198, w12199, w12200, w12201, w12202, w12203, w12204, w12205, w12206, w12207, w12208, w12209, w12210, w12211, w12212, w12213, w12214, w12215, w12216, w12217, w12218, w12219, w12220, w12221, w12222, w12223, w12224, w12225, w12226, w12227, w12228, w12229, w12230, w12231, w12232, w12233, w12234, w12235, w12236, w12237, w12238, w12239, w12240, w12241, w12242, w12243, w12244, w12245, w12246, w12247, w12248, w12249, w12250, w12251, w12252, w12253, w12254, w12255, w12256, w12257, w12258, w12259, w12260, w12261, w12262, w12263, w12264, w12265, w12266, w12267, w12268, w12269, w12270, w12271, w12272, w12273, w12274, w12275, w12276, w12277, w12278, w12279, w12280, w12281, w12282, w12283, w12284, w12285, w12286, w12287, w12288, w12289, w12290, w12291, w12292, w12293, w12294, w12295, w12296, w12297, w12298, w12299, w12300, w12301, w12302, w12303, w12304, w12305, w12306, w12307, w12308, w12309, w12310, w12311, w12312, w12313, w12314, w12315, w12316, w12317, w12318, w12319, w12320, w12321, w12322, w12323, w12324, w12325, w12326, w12327, w12328, w12329, w12330, w12331, w12332, w12333, w12334, w12335, w12336, w12337, w12338, w12339, w12340, w12341, w12342, w12343, w12344, w12345, w12346, w12347, w12348, w12349, w12350, w12351, w12352, w12353, w12354, w12355, w12356, w12357, w12358, w12359, w12360, w12361, w12362, w12363, w12364, w12365, w12366, w12367, w12368, w12369, w12370, w12371, w12372, w12373, w12374, w12375, w12376, w12377, w12378, w12379, w12380, w12381, w12382, w12383, w12384, w12385, w12386, w12387, w12388, w12389, w12390, w12391, w12392, w12393, w12394, w12395, w12396, w12397, w12398, w12399, w12400, w12401, w12402, w12403, w12404, w12405, w12406, w12407, w12408, w12409, w12410, w12411, w12412, w12413, w12414, w12415, w12416, w12417, w12418, w12419, w12420, w12421, w12422, w12423, w12424, w12425, w12426, w12427, w12428, w12429, w12430, w12431, w12432, w12433, w12434, w12435, w12436, w12437, w12438, w12439, w12440, w12441, w12442, w12443, w12444, w12445, w12446, w12447, w12448, w12449, w12450, w12451, w12452, w12453, w12454, w12455, w12456, w12457, w12458, w12459, w12460, w12461, w12462, w12463, w12464, w12465, w12466, w12467, w12468, w12469, w12470, w12471, w12472, w12473, w12474, w12475, w12476, w12477, w12478, w12479, w12480, w12481, w12482, w12483, w12484, w12485, w12486, w12487, w12488, w12489, w12490, w12491, w12492, w12493, w12494, w12495, w12496, w12497, w12498, w12499, w12500, w12501, w12502, w12503, w12504, w12505, w12506, w12507, w12508, w12509, w12510, w12511, w12512, w12513, w12514, w12515, w12516, w12517, w12518, w12519, w12520, w12521, w12522, w12523, w12524, w12525, w12526, w12527, w12528, w12529, w12530, w12531, w12532, w12533, w12534, w12535, w12536, w12537, w12538, w12539, w12540, w12541, w12542, w12543, w12544, w12545, w12546, w12547, w12548, w12549, w12550, w12551, w12552, w12553, w12554, w12555, w12556, w12557, w12558, w12559, w12560, w12561, w12562, w12563, w12564, w12565, w12566, w12567, w12568, w12569, w12570, w12571, w12572, w12573, w12574, w12575, w12576, w12577, w12578, w12579, w12580, w12581, w12582, w12583, w12584, w12585, w12586, w12587, w12588, w12589, w12590, w12591, w12592, w12593, w12594, w12595, w12596, w12597, w12598, w12599, w12600, w12601, w12602, w12603, w12604, w12605, w12606, w12607, w12608, w12609, w12610, w12611, w12612, w12613, w12614, w12615, w12616, w12617, w12618, w12619, w12620, w12621, w12622, w12623, w12624, w12625, w12626, w12627, w12628, w12629, w12630, w12631, w12632, w12633, w12634, w12635, w12636, w12637, w12638, w12639, w12640, w12641, w12642, w12643, w12644, w12645, w12646, w12647, w12648, w12649, w12650, w12651, w12652, w12653, w12654, w12655, w12656, w12657, w12658, w12659, w12660, w12661, w12662, w12663, w12664, w12665, w12666, w12667, w12668, w12669, w12670, w12671, w12672, w12673, w12674, w12675, w12676, w12677, w12678, w12679, w12680, w12681, w12682, w12683, w12684, w12685, w12686, w12687, w12688, w12689, w12690, w12691, w12692, w12693, w12694, w12695, w12696, w12697, w12698, w12699, w12700, w12701, w12702, w12703, w12704, w12705, w12706, w12707, w12708, w12709, w12710, w12711, w12712, w12713, w12714, w12715, w12716, w12717, w12718, w12719, w12720, w12721, w12722, w12723, w12724, w12725, w12726, w12727, w12728, w12729, w12730, w12731, w12732, w12733, w12734, w12735, w12736, w12737, w12738, w12739, w12740, w12741, w12742, w12743, w12744, w12745, w12746, w12747, w12748, w12749, w12750, w12751, w12752, w12753, w12754, w12755, w12756, w12757, w12758, w12759, w12760, w12761, w12762, w12763, w12764, w12765, w12766, w12767, w12768, w12769, w12770, w12771, w12772, w12773, w12774, w12775, w12776, w12777, w12778, w12779, w12780, w12781, w12782, w12783, w12784, w12785, w12786, w12787, w12788, w12789, w12790, w12791, w12792, w12793, w12794, w12795, w12796, w12797, w12798, w12799, w12800, w12801, w12802, w12803, w12804, w12805, w12806, w12807, w12808, w12809, w12810, w12811, w12812, w12813, w12814, w12815, w12816, w12817, w12818, w12819, w12820, w12821, w12822, w12823, w12824, w12825, w12826, w12827, w12828, w12829, w12830, w12831, w12832, w12833, w12834, w12835, w12836, w12837, w12838, w12839, w12840, w12841, w12842, w12843, w12844, w12845, w12846, w12847, w12848, w12849, w12850, w12851, w12852, w12853, w12854, w12855, w12856, w12857, w12858, w12859, w12860, w12861, w12862, w12863, w12864, w12865, w12866, w12867, w12868, w12869, w12870, w12871, w12872, w12873, w12874, w12875, w12876, w12877, w12878, w12879, w12880, w12881, w12882, w12883, w12884, w12885, w12886, w12887, w12888, w12889, w12890, w12891, w12892, w12893, w12894, w12895, w12896, w12897, w12898, w12899, w12900, w12901, w12902, w12903, w12904, w12905, w12906, w12907, w12908, w12909, w12910, w12911, w12912, w12913, w12914, w12915, w12916, w12917, w12918, w12919, w12920, w12921, w12922, w12923, w12924, w12925, w12926, w12927, w12928, w12929, w12930, w12931, w12932, w12933, w12934, w12935, w12936, w12937, w12938, w12939, w12940, w12941, w12942, w12943, w12944, w12945, w12946, w12947, w12948, w12949, w12950, w12951, w12952, w12953, w12954, w12955, w12956, w12957, w12958, w12959, w12960, w12961, w12962, w12963, w12964, w12965, w12966, w12967, w12968, w12969, w12970, w12971, w12972, w12973, w12974, w12975, w12976, w12977, w12978, w12979, w12980, w12981, w12982, w12983, w12984, w12985, w12986, w12987, w12988, w12989, w12990, w12991, w12992, w12993, w12994, w12995, w12996, w12997, w12998, w12999, w13000, w13001, w13002, w13003, w13004, w13005, w13006, w13007, w13008, w13009, w13010, w13011, w13012, w13013, w13014, w13015, w13016, w13017, w13018, w13019, w13020, w13021, w13022, w13023, w13024, w13025, w13026, w13027, w13028, w13029, w13030, w13031, w13032, w13033, w13034, w13035, w13036, w13037, w13038, w13039, w13040, w13041, w13042, w13043, w13044, w13045, w13046, w13047, w13048, w13049, w13050, w13051, w13052, w13053, w13054, w13055, w13056, w13057, w13058, w13059, w13060, w13061, w13062, w13063, w13064, w13065, w13066, w13067, w13068, w13069, w13070, w13071, w13072, w13073, w13074, w13075, w13076, w13077, w13078, w13079, w13080, w13081, w13082, w13083, w13084, w13085, w13086, w13087, w13088, w13089, w13090, w13091, w13092, w13093, w13094, w13095, w13096, w13097, w13098, w13099, w13100, w13101, w13102, w13103, w13104, w13105, w13106, w13107, w13108, w13109, w13110, w13111, w13112, w13113, w13114, w13115, w13116, w13117, w13118, w13119, w13120, w13121, w13122, w13123, w13124, w13125, w13126, w13127, w13128, w13129, w13130, w13131, w13132, w13133, w13134, w13135, w13136, w13137, w13138, w13139, w13140, w13141, w13142, w13143, w13144, w13145, w13146, w13147, w13148, w13149, w13150, w13151, w13152, w13153, w13154, w13155, w13156, w13157, w13158, w13159, w13160, w13161, w13162, w13163, w13164, w13165, w13166, w13167, w13168, w13169, w13170, w13171, w13172, w13173, w13174, w13175, w13176, w13177, w13178, w13179, w13180, w13181, w13182, w13183, w13184, w13185, w13186, w13187, w13188, w13189, w13190, w13191, w13192, w13193, w13194, w13195, w13196, w13197, w13198, w13199, w13200, w13201, w13202, w13203, w13204, w13205, w13206, w13207, w13208, w13209, w13210, w13211, w13212, w13213, w13214, w13215, w13216, w13217, w13218, w13219, w13220, w13221, w13222, w13223, w13224, w13225, w13226, w13227, w13228, w13229, w13230, w13231, w13232, w13233, w13234, w13235, w13236, w13237, w13238, w13239, w13240, w13241, w13242, w13243, w13244, w13245, w13246, w13247, w13248, w13249, w13250, w13251, w13252, w13253, w13254, w13255, w13256, w13257, w13258, w13259, w13260, w13261, w13262, w13263, w13264, w13265, w13266, w13267, w13268, w13269, w13270, w13271, w13272, w13273, w13274, w13275, w13276, w13277, w13278, w13279, w13280, w13281, w13282, w13283, w13284, w13285, w13286, w13287, w13288, w13289, w13290, w13291, w13292, w13293, w13294, w13295, w13296, w13297, w13298, w13299, w13300, w13301, w13302, w13303, w13304, w13305, w13306, w13307, w13308, w13309, w13310, w13311, w13312, w13313, w13314, w13315, w13316, w13317, w13318, w13319, w13320, w13321, w13322, w13323, w13324, w13325, w13326, w13327, w13328, w13329, w13330, w13331, w13332, w13333, w13334, w13335, w13336, w13337, w13338, w13339, w13340, w13341, w13342, w13343, w13344, w13345, w13346, w13347, w13348, w13349, w13350, w13351, w13352, w13353, w13354, w13355, w13356, w13357, w13358, w13359, w13360, w13361, w13362, w13363, w13364, w13365, w13366, w13367, w13368, w13369, w13370, w13371, w13372, w13373, w13374, w13375, w13376, w13377, w13378, w13379, w13380, w13381, w13382, w13383, w13384, w13385, w13386, w13387, w13388, w13389, w13390, w13391, w13392, w13393, w13394, w13395, w13396, w13397, w13398, w13399, w13400, w13401, w13402, w13403, w13404, w13405, w13406, w13407, w13408, w13409, w13410, w13411, w13412, w13413, w13414, w13415, w13416, w13417, w13418, w13419, w13420, w13421, w13422, w13423, w13424, w13425, w13426, w13427, w13428, w13429, w13430, w13431, w13432, w13433, w13434, w13435, w13436, w13437, w13438, w13439, w13440, w13441, w13442, w13443, w13444, w13445, w13446, w13447, w13448, w13449, w13450, w13451, w13452, w13453, w13454, w13455, w13456, w13457, w13458, w13459, w13460, w13461, w13462, w13463, w13464, w13465, w13466, w13467, w13468, w13469, w13470, w13471, w13472, w13473, w13474, w13475, w13476, w13477, w13478, w13479, w13480, w13481, w13482, w13483, w13484, w13485, w13486, w13487, w13488, w13489, w13490, w13491, w13492, w13493, w13494, w13495, w13496, w13497, w13498, w13499, w13500, w13501, w13502, w13503, w13504, w13505, w13506, w13507, w13508, w13509, w13510, w13511, w13512, w13513, w13514, w13515, w13516, w13517, w13518, w13519, w13520, w13521, w13522, w13523, w13524, w13525, w13526, w13527, w13528, w13529, w13530, w13531, w13532, w13533, w13534, w13535, w13536, w13537, w13538, w13539, w13540, w13541, w13542, w13543, w13544, w13545, w13546, w13547, w13548, w13549, w13550, w13551, w13552, w13553, w13554, w13555, w13556, w13557, w13558, w13559, w13560, w13561, w13562, w13563, w13564, w13565, w13566, w13567, w13568, w13569, w13570, w13571, w13572, w13573, w13574, w13575, w13576, w13577, w13578, w13579, w13580, w13581, w13582, w13583, w13584, w13585, w13586, w13587, w13588, w13589, w13590, w13591, w13592, w13593, w13594, w13595, w13596, w13597, w13598, w13599, w13600, w13601, w13602, w13603, w13604, w13605, w13606, w13607, w13608, w13609, w13610, w13611, w13612, w13613, w13614, w13615, w13616, w13617, w13618, w13619, w13620, w13621, w13622, w13623, w13624, w13625, w13626, w13627, w13628, w13629, w13630, w13631, w13632, w13633, w13634, w13635, w13636, w13637, w13638, w13639, w13640, w13641, w13642, w13643, w13644, w13645, w13646, w13647, w13648, w13649, w13650, w13651, w13652, w13653, w13654, w13655, w13656, w13657, w13658, w13659, w13660, w13661, w13662, w13663, w13664, w13665, w13666, w13667, w13668, w13669, w13670, w13671, w13672, w13673, w13674, w13675, w13676, w13677, w13678, w13679, w13680, w13681, w13682, w13683, w13684, w13685, w13686, w13687, w13688, w13689, w13690, w13691, w13692, w13693, w13694, w13695, w13696, w13697, w13698, w13699, w13700, w13701, w13702, w13703, w13704, w13705, w13706, w13707, w13708, w13709, w13710, w13711, w13712, w13713, w13714, w13715, w13716, w13717, w13718, w13719, w13720, w13721, w13722, w13723, w13724, w13725, w13726, w13727, w13728, w13729, w13730, w13731, w13732, w13733, w13734, w13735, w13736, w13737, w13738, w13739, w13740, w13741, w13742, w13743, w13744, w13745, w13746, w13747, w13748, w13749, w13750, w13751, w13752, w13753, w13754, w13755, w13756, w13757, w13758, w13759, w13760, w13761, w13762, w13763, w13764, w13765, w13766, w13767, w13768, w13769, w13770, w13771, w13772, w13773, w13774, w13775, w13776, w13777, w13778, w13779, w13780, w13781, w13782, w13783, w13784, w13785, w13786, w13787, w13788, w13789, w13790, w13791, w13792, w13793, w13794, w13795, w13796, w13797, w13798, w13799, w13800, w13801, w13802, w13803, w13804, w13805, w13806, w13807, w13808, w13809, w13810, w13811, w13812, w13813, w13814, w13815, w13816, w13817, w13818, w13819, w13820, w13821, w13822, w13823, w13824, w13825, w13826, w13827, w13828, w13829, w13830, w13831, w13832, w13833, w13834, w13835, w13836, w13837, w13838, w13839, w13840, w13841, w13842, w13843, w13844, w13845, w13846, w13847, w13848, w13849, w13850, w13851, w13852, w13853, w13854, w13855, w13856, w13857, w13858, w13859, w13860, w13861, w13862, w13863, w13864, w13865, w13866, w13867, w13868, w13869, w13870, w13871, w13872, w13873, w13874, w13875, w13876, w13877, w13878, w13879, w13880, w13881, w13882, w13883, w13884, w13885, w13886, w13887, w13888, w13889, w13890, w13891, w13892, w13893, w13894, w13895, w13896, w13897, w13898, w13899, w13900, w13901, w13902, w13903, w13904, w13905, w13906, w13907, w13908, w13909, w13910, w13911, w13912, w13913, w13914, w13915, w13916, w13917, w13918, w13919, w13920, w13921, w13922, w13923, w13924, w13925, w13926, w13927, w13928, w13929, w13930, w13931, w13932, w13933, w13934, w13935, w13936, w13937, w13938, w13939, w13940, w13941, w13942, w13943, w13944, w13945, w13946, w13947, w13948, w13949, w13950, w13951, w13952, w13953, w13954, w13955, w13956, w13957, w13958, w13959, w13960, w13961, w13962, w13963, w13964, w13965, w13966, w13967, w13968, w13969, w13970, w13971, w13972, w13973, w13974, w13975, w13976, w13977, w13978, w13979, w13980, w13981, w13982, w13983, w13984, w13985, w13986, w13987, w13988, w13989, w13990, w13991, w13992, w13993, w13994, w13995, w13996, w13997, w13998, w13999, w14000, w14001, w14002, w14003, w14004, w14005, w14006, w14007, w14008, w14009, w14010, w14011, w14012, w14013, w14014, w14015, w14016, w14017, w14018, w14019, w14020, w14021, w14022, w14023, w14024, w14025, w14026, w14027, w14028, w14029, w14030, w14031, w14032, w14033, w14034, w14035, w14036, w14037, w14038, w14039, w14040, w14041, w14042, w14043, w14044, w14045, w14046, w14047, w14048, w14049, w14050, w14051, w14052, w14053, w14054, w14055, w14056, w14057, w14058, w14059, w14060, w14061, w14062, w14063, w14064, w14065, w14066, w14067, w14068, w14069, w14070, w14071, w14072, w14073, w14074, w14075, w14076, w14077, w14078, w14079, w14080, w14081, w14082, w14083, w14084, w14085, w14086, w14087, w14088, w14089, w14090, w14091, w14092, w14093, w14094, w14095, w14096, w14097, w14098, w14099, w14100, w14101, w14102, w14103, w14104, w14105, w14106, w14107, w14108, w14109, w14110, w14111, w14112, w14113, w14114, w14115, w14116, w14117, w14118, w14119, w14120, w14121, w14122, w14123, w14124, w14125, w14126, w14127, w14128, w14129, w14130, w14131, w14132, w14133, w14134, w14135, w14136, w14137, w14138, w14139, w14140, w14141, w14142, w14143, w14144, w14145, w14146, w14147, w14148, w14149, w14150, w14151, w14152, w14153, w14154, w14155, w14156, w14157, w14158, w14159, w14160, w14161, w14162, w14163, w14164, w14165, w14166, w14167, w14168, w14169, w14170, w14171, w14172, w14173, w14174, w14175, w14176, w14177, w14178, w14179, w14180, w14181, w14182, w14183, w14184, w14185, w14186, w14187, w14188, w14189, w14190, w14191, w14192, w14193, w14194, w14195, w14196, w14197, w14198, w14199, w14200, w14201, w14202, w14203, w14204, w14205, w14206, w14207, w14208, w14209, w14210, w14211, w14212, w14213, w14214, w14215, w14216, w14217, w14218, w14219, w14220, w14221, w14222, w14223, w14224, w14225, w14226, w14227, w14228, w14229, w14230, w14231, w14232, w14233, w14234, w14235, w14236, w14237, w14238, w14239, w14240, w14241, w14242, w14243, w14244, w14245, w14246, w14247, w14248, w14249, w14250, w14251, w14252, w14253, w14254, w14255, w14256, w14257, w14258, w14259, w14260, w14261, w14262, w14263, w14264, w14265, w14266, w14267, w14268, w14269, w14270, w14271, w14272, w14273, w14274, w14275, w14276, w14277, w14278, w14279, w14280, w14281, w14282, w14283, w14284, w14285, w14286, w14287, w14288, w14289, w14290, w14291, w14292, w14293, w14294, w14295, w14296, w14297, w14298, w14299, w14300, w14301, w14302, w14303, w14304, w14305, w14306, w14307, w14308, w14309, w14310, w14311, w14312, w14313, w14314, w14315, w14316, w14317, w14318, w14319, w14320, w14321, w14322, w14323, w14324, w14325, w14326, w14327, w14328, w14329, w14330, w14331, w14332, w14333, w14334, w14335, w14336, w14337, w14338, w14339, w14340, w14341, w14342, w14343, w14344, w14345, w14346, w14347, w14348, w14349, w14350, w14351, w14352, w14353, w14354, w14355, w14356, w14357, w14358, w14359, w14360, w14361, w14362, w14363, w14364, w14365, w14366, w14367, w14368, w14369, w14370, w14371, w14372, w14373, w14374, w14375, w14376, w14377, w14378, w14379, w14380, w14381, w14382, w14383, w14384, w14385, w14386, w14387, w14388, w14389, w14390, w14391, w14392, w14393, w14394, w14395, w14396, w14397, w14398, w14399, w14400, w14401, w14402, w14403, w14404, w14405, w14406, w14407, w14408, w14409, w14410, w14411, w14412, w14413, w14414, w14415, w14416, w14417, w14418, w14419, w14420, w14421, w14422, w14423, w14424, w14425, w14426, w14427, w14428, w14429, w14430, w14431, w14432, w14433, w14434, w14435, w14436, w14437, w14438, w14439, w14440, w14441, w14442, w14443, w14444, w14445, w14446, w14447, w14448, w14449, w14450, w14451, w14452, w14453, w14454, w14455, w14456, w14457, w14458, w14459, w14460, w14461, w14462, w14463, w14464, w14465, w14466, w14467, w14468, w14469, w14470, w14471, w14472, w14473, w14474, w14475, w14476, w14477, w14478, w14479, w14480, w14481, w14482, w14483, w14484, w14485, w14486, w14487, w14488, w14489, w14490, w14491, w14492, w14493, w14494, w14495, w14496, w14497, w14498, w14499, w14500, w14501, w14502, w14503, w14504, w14505, w14506, w14507, w14508, w14509, w14510, w14511, w14512, w14513, w14514, w14515, w14516, w14517, w14518, w14519, w14520, w14521, w14522, w14523, w14524, w14525, w14526, w14527, w14528, w14529, w14530, w14531, w14532, w14533, w14534, w14535, w14536, w14537, w14538, w14539, w14540, w14541, w14542, w14543, w14544, w14545, w14546, w14547, w14548, w14549, w14550, w14551, w14552, w14553, w14554, w14555, w14556, w14557, w14558, w14559, w14560, w14561, w14562, w14563, w14564, w14565, w14566, w14567, w14568, w14569, w14570, w14571, w14572, w14573, w14574, w14575, w14576, w14577, w14578, w14579, w14580, w14581, w14582, w14583, w14584, w14585, w14586, w14587, w14588, w14589, w14590, w14591, w14592, w14593, w14594, w14595, w14596, w14597, w14598, w14599, w14600, w14601, w14602, w14603, w14604, w14605, w14606, w14607, w14608, w14609, w14610, w14611, w14612, w14613, w14614, w14615, w14616, w14617, w14618, w14619, w14620, w14621, w14622, w14623, w14624, w14625, w14626, w14627, w14628, w14629, w14630, w14631, w14632, w14633, w14634, w14635, w14636, w14637, w14638, w14639, w14640, w14641, w14642, w14643, w14644, w14645, w14646, w14647, w14648, w14649, w14650, w14651, w14652, w14653, w14654, w14655, w14656, w14657, w14658, w14659, w14660, w14661, w14662, w14663, w14664, w14665, w14666, w14667, w14668, w14669, w14670, w14671, w14672, w14673, w14674, w14675, w14676, w14677, w14678, w14679, w14680, w14681, w14682, w14683, w14684, w14685, w14686, w14687, w14688, w14689, w14690, w14691, w14692, w14693, w14694, w14695, w14696, w14697, w14698, w14699, w14700, w14701, w14702, w14703, w14704, w14705, w14706, w14707, w14708, w14709, w14710, w14711, w14712, w14713, w14714, w14715, w14716, w14717, w14718, w14719, w14720, w14721, w14722, w14723, w14724, w14725, w14726, w14727, w14728, w14729, w14730, w14731, w14732, w14733, w14734, w14735, w14736, w14737, w14738, w14739, w14740, w14741, w14742, w14743, w14744, w14745, w14746, w14747, w14748, w14749, w14750, w14751, w14752, w14753, w14754, w14755, w14756, w14757, w14758, w14759, w14760, w14761, w14762, w14763, w14764, w14765, w14766, w14767, w14768, w14769, w14770, w14771, w14772, w14773, w14774, w14775, w14776, w14777, w14778, w14779, w14780, w14781, w14782, w14783, w14784, w14785, w14786, w14787, w14788, w14789, w14790, w14791, w14792, w14793, w14794, w14795, w14796, w14797, w14798, w14799, w14800, w14801, w14802, w14803, w14804, w14805, w14806, w14807, w14808, w14809, w14810, w14811, w14812, w14813, w14814, w14815, w14816, w14817, w14818, w14819, w14820, w14821, w14822, w14823, w14824, w14825, w14826, w14827, w14828, w14829, w14830, w14831, w14832, w14833, w14834, w14835, w14836, w14837, w14838, w14839, w14840, w14841, w14842, w14843, w14844, w14845, w14846, w14847, w14848, w14849, w14850, w14851, w14852, w14853, w14854, w14855, w14856, w14857, w14858, w14859, w14860, w14861, w14862, w14863, w14864, w14865, w14866, w14867, w14868, w14869, w14870, w14871, w14872, w14873, w14874, w14875, w14876, w14877, w14878, w14879, w14880, w14881, w14882, w14883, w14884, w14885, w14886, w14887, w14888, w14889, w14890, w14891, w14892, w14893, w14894, w14895, w14896, w14897, w14898, w14899, w14900, w14901, w14902, w14903, w14904, w14905, w14906, w14907, w14908, w14909, w14910, w14911, w14912, w14913, w14914, w14915, w14916, w14917, w14918, w14919, w14920, w14921, w14922, w14923, w14924, w14925, w14926, w14927, w14928, w14929, w14930, w14931, w14932, w14933, w14934, w14935, w14936, w14937, w14938, w14939, w14940, w14941, w14942, w14943, w14944, w14945, w14946, w14947, w14948, w14949, w14950, w14951, w14952, w14953, w14954, w14955, w14956, w14957, w14958, w14959, w14960, w14961, w14962, w14963, w14964, w14965, w14966, w14967, w14968, w14969, w14970, w14971, w14972, w14973, w14974, w14975, w14976, w14977, w14978, w14979, w14980, w14981, w14982, w14983, w14984, w14985, w14986, w14987, w14988, w14989, w14990, w14991, w14992, w14993, w14994, w14995, w14996, w14997, w14998, w14999, w15000, w15001, w15002, w15003, w15004, w15005, w15006, w15007, w15008, w15009, w15010, w15011, w15012, w15013, w15014, w15015, w15016, w15017, w15018, w15019, w15020, w15021, w15022, w15023, w15024, w15025, w15026, w15027, w15028, w15029, w15030, w15031, w15032, w15033, w15034, w15035, w15036, w15037, w15038, w15039, w15040, w15041, w15042, w15043, w15044, w15045, w15046, w15047, w15048, w15049, w15050, w15051, w15052, w15053, w15054, w15055, w15056, w15057, w15058, w15059, w15060, w15061, w15062, w15063, w15064, w15065, w15066, w15067, w15068, w15069, w15070, w15071, w15072, w15073, w15074, w15075, w15076, w15077, w15078, w15079, w15080, w15081, w15082, w15083, w15084, w15085, w15086, w15087, w15088, w15089, w15090, w15091, w15092, w15093, w15094, w15095, w15096, w15097, w15098, w15099, w15100, w15101, w15102, w15103, w15104, w15105, w15106, w15107, w15108, w15109, w15110, w15111, w15112, w15113, w15114, w15115, w15116, w15117, w15118, w15119, w15120, w15121, w15122, w15123, w15124, w15125, w15126, w15127, w15128, w15129, w15130, w15131, w15132, w15133, w15134, w15135, w15136, w15137, w15138, w15139, w15140, w15141, w15142, w15143, w15144, w15145, w15146, w15147, w15148, w15149, w15150, w15151, w15152, w15153, w15154, w15155, w15156, w15157, w15158, w15159, w15160, w15161, w15162, w15163, w15164, w15165, w15166, w15167, w15168, w15169, w15170, w15171, w15172, w15173, w15174, w15175, w15176, w15177, w15178, w15179, w15180, w15181, w15182, w15183, w15184, w15185, w15186, w15187, w15188, w15189, w15190, w15191, w15192, w15193, w15194, w15195, w15196, w15197, w15198, w15199, w15200, w15201, w15202, w15203, w15204, w15205, w15206, w15207, w15208, w15209, w15210, w15211, w15212, w15213, w15214, w15215, w15216, w15217, w15218, w15219, w15220, w15221, w15222, w15223, w15224, w15225, w15226, w15227, w15228, w15229, w15230, w15231, w15232, w15233, w15234, w15235, w15236, w15237, w15238, w15239, w15240, w15241, w15242, w15243, w15244, w15245, w15246, w15247, w15248, w15249, w15250, w15251, w15252, w15253, w15254, w15255, w15256, w15257, w15258, w15259, w15260, w15261, w15262, w15263, w15264, w15265, w15266, w15267, w15268, w15269, w15270, w15271, w15272, w15273, w15274, w15275, w15276, w15277, w15278, w15279, w15280, w15281, w15282, w15283, w15284, w15285, w15286, w15287, w15288, w15289, w15290, w15291, w15292, w15293, w15294, w15295, w15296, w15297, w15298, w15299, w15300, w15301, w15302, w15303, w15304, w15305, w15306, w15307, w15308, w15309, w15310, w15311, w15312, w15313, w15314, w15315, w15316, w15317, w15318, w15319, w15320, w15321, w15322, w15323, w15324, w15325, w15326, w15327, w15328, w15329, w15330, w15331, w15332, w15333, w15334, w15335, w15336, w15337, w15338, w15339, w15340, w15341, w15342, w15343, w15344, w15345, w15346, w15347, w15348, w15349, w15350, w15351, w15352, w15353, w15354, w15355, w15356, w15357, w15358, w15359, w15360, w15361, w15362, w15363, w15364, w15365, w15366, w15367, w15368, w15369, w15370, w15371, w15372, w15373, w15374, w15375, w15376, w15377, w15378, w15379, w15380, w15381, w15382, w15383, w15384, w15385, w15386, w15387, w15388, w15389, w15390, w15391, w15392, w15393, w15394, w15395, w15396, w15397, w15398, w15399, w15400, w15401, w15402, w15403, w15404, w15405, w15406, w15407, w15408, w15409, w15410, w15411, w15412, w15413, w15414, w15415, w15416, w15417, w15418, w15419, w15420, w15421, w15422, w15423, w15424, w15425, w15426, w15427, w15428, w15429, w15430, w15431, w15432, w15433, w15434, w15435, w15436, w15437, w15438, w15439, w15440, w15441, w15442, w15443, w15444, w15445, w15446, w15447, w15448, w15449, w15450, w15451, w15452, w15453, w15454, w15455, w15456, w15457, w15458, w15459, w15460, w15461, w15462, w15463, w15464, w15465, w15466, w15467, w15468, w15469, w15470, w15471, w15472, w15473, w15474, w15475, w15476, w15477, w15478, w15479, w15480, w15481, w15482, w15483, w15484, w15485, w15486, w15487, w15488, w15489, w15490, w15491, w15492, w15493, w15494, w15495, w15496, w15497, w15498, w15499, w15500, w15501, w15502, w15503, w15504, w15505, w15506, w15507, w15508, w15509, w15510, w15511, w15512, w15513, w15514, w15515, w15516, w15517, w15518, w15519, w15520, w15521, w15522, w15523, w15524, w15525, w15526, w15527, w15528, w15529, w15530, w15531, w15532, w15533, w15534, w15535, w15536, w15537, w15538, w15539, w15540, w15541, w15542, w15543, w15544, w15545, w15546, w15547, w15548, w15549, w15550, w15551, w15552, w15553, w15554, w15555, w15556, w15557, w15558, w15559, w15560, w15561, w15562, w15563, w15564, w15565, w15566, w15567, w15568, w15569, w15570, w15571, w15572, w15573, w15574, w15575, w15576, w15577, w15578, w15579, w15580, w15581, w15582, w15583, w15584, w15585, w15586, w15587, w15588, w15589, w15590, w15591, w15592, w15593, w15594, w15595, w15596, w15597, w15598, w15599, w15600, w15601, w15602, w15603, w15604, w15605, w15606, w15607, w15608, w15609, w15610, w15611, w15612, w15613, w15614, w15615, w15616, w15617, w15618, w15619, w15620, w15621, w15622, w15623, w15624, w15625, w15626, w15627, w15628, w15629, w15630, w15631, w15632, w15633, w15634, w15635, w15636, w15637, w15638, w15639, w15640, w15641, w15642, w15643, w15644, w15645, w15646, w15647, w15648, w15649, w15650, w15651, w15652, w15653, w15654, w15655, w15656, w15657, w15658, w15659, w15660, w15661, w15662, w15663, w15664, w15665, w15666, w15667, w15668, w15669, w15670, w15671, w15672, w15673, w15674, w15675, w15676, w15677, w15678, w15679, w15680, w15681, w15682, w15683, w15684, w15685, w15686, w15687, w15688, w15689, w15690, w15691, w15692, w15693, w15694, w15695, w15696, w15697, w15698, w15699, w15700, w15701, w15702, w15703, w15704, w15705, w15706, w15707, w15708, w15709, w15710, w15711, w15712, w15713, w15714, w15715, w15716, w15717, w15718, w15719, w15720, w15721, w15722, w15723, w15724, w15725, w15726, w15727, w15728, w15729, w15730, w15731, w15732, w15733, w15734, w15735, w15736, w15737, w15738, w15739, w15740, w15741, w15742, w15743, w15744, w15745, w15746, w15747, w15748, w15749, w15750, w15751, w15752, w15753, w15754, w15755, w15756, w15757, w15758, w15759, w15760, w15761, w15762, w15763, w15764, w15765, w15766, w15767, w15768, w15769, w15770, w15771, w15772, w15773, w15774, w15775, w15776, w15777, w15778, w15779, w15780, w15781, w15782, w15783, w15784, w15785, w15786, w15787, w15788, w15789, w15790, w15791, w15792, w15793, w15794, w15795, w15796, w15797, w15798, w15799, w15800, w15801, w15802, w15803, w15804, w15805, w15806, w15807, w15808, w15809, w15810, w15811, w15812, w15813, w15814, w15815, w15816, w15817, w15818, w15819, w15820, w15821, w15822, w15823, w15824, w15825, w15826, w15827, w15828, w15829, w15830, w15831, w15832, w15833, w15834, w15835, w15836, w15837, w15838, w15839, w15840, w15841, w15842, w15843, w15844, w15845, w15846, w15847, w15848, w15849, w15850, w15851, w15852, w15853, w15854, w15855, w15856, w15857, w15858, w15859, w15860, w15861, w15862, w15863, w15864, w15865, w15866, w15867, w15868, w15869, w15870, w15871, w15872, w15873, w15874, w15875, w15876, w15877, w15878, w15879, w15880, w15881, w15882, w15883, w15884, w15885, w15886, w15887, w15888, w15889, w15890, w15891, w15892, w15893, w15894, w15895, w15896, w15897, w15898, w15899, w15900, w15901, w15902, w15903, w15904, w15905, w15906, w15907, w15908, w15909, w15910, w15911, w15912, w15913, w15914, w15915, w15916, w15917, w15918, w15919, w15920, w15921, w15922, w15923, w15924, w15925, w15926, w15927, w15928, w15929, w15930, w15931, w15932, w15933, w15934, w15935, w15936, w15937, w15938, w15939, w15940, w15941, w15942, w15943, w15944, w15945, w15946, w15947, w15948, w15949, w15950, w15951, w15952, w15953, w15954, w15955, w15956, w15957, w15958, w15959, w15960, w15961, w15962, w15963, w15964, w15965, w15966, w15967, w15968, w15969, w15970, w15971, w15972, w15973, w15974, w15975, w15976, w15977, w15978, w15979, w15980, w15981, w15982, w15983, w15984, w15985, w15986, w15987, w15988, w15989, w15990, w15991, w15992, w15993, w15994, w15995, w15996, w15997, w15998, w15999, w16000, w16001, w16002, w16003, w16004, w16005, w16006, w16007, w16008, w16009, w16010, w16011, w16012, w16013, w16014, w16015, w16016, w16017, w16018, w16019, w16020, w16021, w16022, w16023, w16024, w16025, w16026, w16027, w16028, w16029, w16030, w16031, w16032, w16033, w16034, w16035, w16036, w16037, w16038, w16039, w16040, w16041, w16042, w16043, w16044, w16045, w16046, w16047, w16048, w16049, w16050, w16051, w16052, w16053, w16054, w16055, w16056, w16057, w16058, w16059, w16060, w16061, w16062, w16063, w16064, w16065, w16066, w16067, w16068, w16069, w16070, w16071, w16072, w16073, w16074, w16075, w16076, w16077, w16078, w16079, w16080, w16081, w16082, w16083, w16084, w16085, w16086, w16087, w16088, w16089, w16090, w16091, w16092, w16093, w16094, w16095, w16096, w16097, w16098, w16099, w16100, w16101, w16102, w16103, w16104, w16105, w16106, w16107, w16108, w16109, w16110, w16111, w16112, w16113, w16114, w16115, w16116, w16117, w16118, w16119, w16120, w16121, w16122, w16123, w16124, w16125, w16126, w16127, w16128, w16129, w16130, w16131, w16132, w16133, w16134, w16135, w16136, w16137, w16138, w16139, w16140, w16141, w16142, w16143, w16144, w16145, w16146, w16147, w16148, w16149, w16150, w16151, w16152, w16153, w16154, w16155, w16156, w16157, w16158, w16159, w16160, w16161, w16162, w16163, w16164, w16165, w16166, w16167, w16168, w16169, w16170, w16171, w16172, w16173, w16174, w16175, w16176, w16177, w16178, w16179, w16180, w16181, w16182, w16183, w16184, w16185, w16186, w16187, w16188, w16189, w16190, w16191, w16192, w16193, w16194, w16195, w16196, w16197, w16198, w16199, w16200, w16201, w16202, w16203, w16204, w16205, w16206, w16207, w16208, w16209, w16210, w16211, w16212, w16213, w16214, w16215, w16216, w16217, w16218, w16219, w16220, w16221, w16222, w16223, w16224, w16225, w16226, w16227, w16228, w16229, w16230, w16231, w16232, w16233, w16234, w16235, w16236, w16237, w16238, w16239, w16240, w16241, w16242, w16243, w16244, w16245, w16246, w16247, w16248, w16249, w16250, w16251, w16252, w16253, w16254, w16255, w16256, w16257, w16258, w16259, w16260, w16261, w16262, w16263, w16264, w16265, w16266, w16267, w16268, w16269, w16270, w16271, w16272, w16273, w16274, w16275, w16276, w16277, w16278, w16279, w16280, w16281, w16282, w16283, w16284, w16285, w16286, w16287, w16288, w16289, w16290, w16291, w16292, w16293, w16294, w16295, w16296, w16297, w16298, w16299, w16300, w16301, w16302, w16303, w16304, w16305, w16306, w16307, w16308, w16309, w16310, w16311, w16312, w16313, w16314, w16315, w16316, w16317, w16318, w16319, w16320, w16321, w16322, w16323, w16324, w16325, w16326, w16327, w16328, w16329, w16330, w16331, w16332, w16333, w16334, w16335, w16336, w16337, w16338, w16339, w16340, w16341, w16342, w16343, w16344, w16345, w16346, w16347, w16348, w16349, w16350, w16351, w16352, w16353, w16354, w16355, w16356, w16357, w16358, w16359, w16360, w16361, w16362, w16363, w16364, w16365, w16366, w16367, w16368, w16369, w16370, w16371, w16372, w16373, w16374, w16375, w16376, w16377, w16378, w16379, w16380, w16381, w16382, w16383, w16384, w16385, w16386, w16387, w16388, w16389, w16390, w16391, w16392, w16393, w16394, w16395, w16396, w16397, w16398, w16399, w16400, w16401, w16402, w16403, w16404, w16405, w16406, w16407, w16408, w16409, w16410, w16411, w16412, w16413, w16414, w16415, w16416, w16417, w16418, w16419, w16420, w16421, w16422, w16423, w16424, w16425, w16426, w16427, w16428, w16429, w16430, w16431, w16432, w16433, w16434, w16435, w16436, w16437, w16438, w16439, w16440, w16441, w16442, w16443, w16444, w16445, w16446, w16447, w16448, w16449, w16450, w16451, w16452, w16453, w16454, w16455, w16456, w16457, w16458, w16459, w16460, w16461, w16462, w16463, w16464, w16465, w16466, w16467, w16468, w16469, w16470, w16471, w16472, w16473, w16474, w16475, w16476, w16477, w16478, w16479, w16480, w16481, w16482, w16483, w16484, w16485, w16486, w16487, w16488, w16489, w16490, w16491, w16492, w16493, w16494, w16495, w16496, w16497, w16498, w16499, w16500, w16501, w16502, w16503, w16504, w16505, w16506, w16507, w16508, w16509, w16510, w16511, w16512, w16513, w16514, w16515, w16516, w16517, w16518, w16519, w16520, w16521, w16522, w16523, w16524, w16525, w16526, w16527, w16528, w16529, w16530, w16531, w16532, w16533, w16534, w16535, w16536, w16537, w16538, w16539, w16540, w16541, w16542, w16543, w16544, w16545, w16546, w16547, w16548, w16549, w16550, w16551, w16552, w16553, w16554, w16555, w16556, w16557, w16558, w16559, w16560, w16561, w16562, w16563, w16564, w16565, w16566, w16567, w16568, w16569, w16570, w16571, w16572, w16573, w16574, w16575, w16576, w16577, w16578, w16579, w16580, w16581, w16582, w16583, w16584, w16585, w16586, w16587, w16588, w16589, w16590, w16591, w16592, w16593, w16594, w16595, w16596, w16597, w16598, w16599, w16600, w16601, w16602, w16603, w16604, w16605, w16606, w16607, w16608, w16609, w16610, w16611, w16612, w16613, w16614, w16615, w16616, w16617, w16618, w16619, w16620, w16621, w16622, w16623, w16624, w16625, w16626, w16627, w16628, w16629, w16630, w16631, w16632, w16633, w16634, w16635, w16636, w16637, w16638, w16639, w16640, w16641, w16642, w16643, w16644, w16645, w16646, w16647, w16648, w16649, w16650, w16651, w16652, w16653, w16654, w16655, w16656, w16657, w16658, w16659, w16660, w16661, w16662, w16663, w16664, w16665, w16666, w16667, w16668, w16669, w16670, w16671, w16672, w16673, w16674, w16675, w16676, w16677, w16678, w16679, w16680, w16681, w16682, w16683, w16684, w16685, w16686, w16687, w16688, w16689, w16690, w16691, w16692, w16693, w16694, w16695, w16696, w16697, w16698, w16699, w16700, w16701, w16702, w16703, w16704, w16705, w16706, w16707, w16708, w16709, w16710, w16711, w16712, w16713, w16714, w16715, w16716, w16717, w16718, w16719, w16720, w16721, w16722, w16723, w16724, w16725, w16726, w16727, w16728, w16729, w16730, w16731, w16732, w16733, w16734, w16735, w16736, w16737, w16738, w16739, w16740, w16741, w16742, w16743, w16744, w16745, w16746, w16747, w16748, w16749, w16750, w16751, w16752, w16753, w16754, w16755, w16756, w16757, w16758, w16759, w16760, w16761, w16762, w16763, w16764, w16765, w16766, w16767, w16768, w16769, w16770, w16771, w16772, w16773, w16774, w16775, w16776, w16777, w16778, w16779, w16780, w16781, w16782, w16783, w16784, w16785, w16786, w16787, w16788, w16789, w16790, w16791, w16792, w16793, w16794, w16795, w16796, w16797, w16798, w16799, w16800, w16801, w16802, w16803, w16804, w16805, w16806, w16807, w16808, w16809, w16810, w16811, w16812, w16813, w16814, w16815, w16816, w16817, w16818, w16819, w16820, w16821, w16822, w16823, w16824, w16825, w16826, w16827, w16828, w16829, w16830, w16831, w16832, w16833, w16834, w16835, w16836, w16837, w16838, w16839, w16840, w16841, w16842, w16843, w16844, w16845, w16846, w16847, w16848, w16849, w16850, w16851, w16852, w16853, w16854, w16855, w16856, w16857, w16858, w16859, w16860, w16861, w16862, w16863, w16864, w16865, w16866, w16867, w16868, w16869, w16870, w16871, w16872, w16873, w16874, w16875, w16876, w16877, w16878, w16879, w16880, w16881, w16882, w16883, w16884, w16885, w16886, w16887, w16888, w16889, w16890, w16891, w16892, w16893, w16894, w16895, w16896, w16897, w16898, w16899, w16900, w16901, w16902, w16903, w16904, w16905, w16906, w16907, w16908, w16909, w16910, w16911, w16912, w16913, w16914, w16915, w16916, w16917, w16918, w16919, w16920, w16921, w16922, w16923, w16924, w16925, w16926, w16927, w16928, w16929, w16930, w16931, w16932, w16933, w16934, w16935, w16936, w16937, w16938, w16939, w16940, w16941, w16942, w16943, w16944, w16945, w16946, w16947, w16948, w16949, w16950, w16951, w16952, w16953, w16954, w16955, w16956, w16957, w16958, w16959, w16960, w16961, w16962, w16963, w16964, w16965, w16966, w16967, w16968, w16969, w16970, w16971, w16972, w16973, w16974, w16975, w16976, w16977, w16978, w16979, w16980, w16981, w16982, w16983, w16984, w16985, w16986, w16987, w16988, w16989, w16990, w16991, w16992, w16993, w16994, w16995, w16996, w16997, w16998, w16999, w17000, w17001, w17002, w17003, w17004, w17005, w17006, w17007, w17008, w17009, w17010, w17011, w17012, w17013, w17014, w17015, w17016, w17017, w17018, w17019, w17020, w17021, w17022, w17023, w17024, w17025, w17026, w17027, w17028, w17029, w17030, w17031, w17032, w17033, w17034, w17035, w17036, w17037, w17038, w17039, w17040, w17041, w17042, w17043, w17044, w17045, w17046, w17047, w17048, w17049, w17050, w17051, w17052, w17053, w17054, w17055, w17056, w17057, w17058, w17059, w17060, w17061, w17062, w17063, w17064, w17065, w17066, w17067, w17068, w17069, w17070, w17071, w17072, w17073, w17074, w17075, w17076, w17077, w17078, w17079, w17080, w17081, w17082, w17083, w17084, w17085, w17086, w17087, w17088, w17089, w17090, w17091, w17092, w17093, w17094, w17095, w17096, w17097, w17098, w17099, w17100, w17101, w17102, w17103, w17104, w17105, w17106, w17107, w17108, w17109, w17110, w17111, w17112, w17113, w17114, w17115, w17116, w17117, w17118, w17119, w17120, w17121, w17122, w17123, w17124, w17125, w17126, w17127, w17128, w17129, w17130, w17131, w17132, w17133, w17134, w17135, w17136, w17137, w17138, w17139, w17140, w17141, w17142, w17143, w17144, w17145, w17146, w17147, w17148, w17149, w17150, w17151, w17152, w17153, w17154, w17155, w17156, w17157, w17158, w17159, w17160, w17161, w17162, w17163, w17164, w17165, w17166, w17167, w17168, w17169, w17170, w17171, w17172, w17173, w17174, w17175, w17176, w17177, w17178, w17179, w17180, w17181, w17182, w17183, w17184, w17185, w17186, w17187, w17188, w17189, w17190, w17191, w17192, w17193, w17194, w17195, w17196, w17197, w17198, w17199, w17200, w17201, w17202, w17203, w17204, w17205, w17206, w17207, w17208, w17209, w17210, w17211, w17212, w17213, w17214, w17215, w17216, w17217, w17218, w17219, w17220, w17221, w17222, w17223, w17224, w17225, w17226, w17227, w17228, w17229, w17230, w17231, w17232, w17233, w17234, w17235, w17236, w17237, w17238, w17239, w17240, w17241, w17242, w17243, w17244, w17245, w17246, w17247, w17248, w17249, w17250, w17251, w17252, w17253, w17254, w17255, w17256, w17257, w17258, w17259, w17260, w17261, w17262, w17263, w17264, w17265, w17266, w17267, w17268, w17269, w17270, w17271, w17272, w17273, w17274, w17275, w17276, w17277, w17278, w17279, w17280, w17281, w17282, w17283, w17284, w17285, w17286, w17287, w17288, w17289, w17290, w17291, w17292, w17293, w17294, w17295, w17296, w17297, w17298, w17299, w17300, w17301, w17302, w17303, w17304, w17305, w17306, w17307, w17308, w17309, w17310, w17311, w17312, w17313, w17314, w17315, w17316, w17317, w17318, w17319, w17320, w17321, w17322, w17323, w17324, w17325, w17326, w17327, w17328, w17329, w17330, w17331, w17332, w17333, w17334, w17335, w17336, w17337, w17338, w17339, w17340, w17341, w17342, w17343, w17344, w17345, w17346, w17347, w17348, w17349, w17350, w17351, w17352, w17353, w17354, w17355, w17356, w17357, w17358, w17359, w17360, w17361, w17362, w17363, w17364, w17365, w17366, w17367, w17368, w17369, w17370, w17371, w17372, w17373, w17374, w17375, w17376, w17377, w17378, w17379, w17380, w17381, w17382, w17383, w17384, w17385, w17386, w17387, w17388, w17389, w17390, w17391, w17392, w17393, w17394, w17395, w17396, w17397, w17398, w17399, w17400, w17401, w17402, w17403, w17404, w17405, w17406, w17407, w17408, w17409, w17410, w17411, w17412, w17413, w17414, w17415, w17416, w17417, w17418, w17419, w17420, w17421, w17422, w17423, w17424, w17425, w17426, w17427, w17428, w17429, w17430, w17431, w17432, w17433, w17434, w17435, w17436, w17437, w17438, w17439, w17440, w17441, w17442, w17443, w17444, w17445, w17446, w17447, w17448, w17449, w17450, w17451, w17452, w17453, w17454, w17455, w17456, w17457, w17458, w17459, w17460, w17461, w17462, w17463, w17464, w17465, w17466, w17467, w17468, w17469, w17470, w17471, w17472, w17473, w17474, w17475, w17476, w17477, w17478, w17479, w17480, w17481, w17482, w17483, w17484, w17485, w17486, w17487, w17488, w17489, w17490, w17491, w17492, w17493, w17494, w17495, w17496, w17497, w17498, w17499, w17500, w17501, w17502, w17503, w17504, w17505, w17506, w17507, w17508, w17509, w17510, w17511, w17512, w17513, w17514, w17515, w17516, w17517, w17518, w17519, w17520, w17521, w17522, w17523, w17524, w17525, w17526, w17527, w17528, w17529, w17530, w17531, w17532, w17533, w17534, w17535, w17536, w17537, w17538, w17539, w17540, w17541, w17542, w17543, w17544, w17545, w17546, w17547, w17548, w17549, w17550, w17551, w17552, w17553, w17554, w17555, w17556, w17557, w17558, w17559, w17560, w17561, w17562, w17563, w17564, w17565, w17566, w17567, w17568, w17569, w17570, w17571, w17572, w17573, w17574, w17575, w17576, w17577, w17578, w17579, w17580, w17581, w17582, w17583, w17584, w17585, w17586, w17587, w17588, w17589, w17590, w17591, w17592, w17593, w17594, w17595, w17596, w17597, w17598, w17599, w17600, w17601, w17602, w17603, w17604, w17605, w17606, w17607, w17608, w17609, w17610, w17611, w17612, w17613, w17614, w17615, w17616, w17617, w17618, w17619, w17620, w17621, w17622, w17623, w17624, w17625, w17626, w17627, w17628, w17629, w17630, w17631, w17632, w17633, w17634, w17635, w17636, w17637, w17638, w17639, w17640, w17641, w17642, w17643, w17644, w17645, w17646, w17647, w17648, w17649, w17650, w17651, w17652, w17653, w17654, w17655, w17656, w17657, w17658, w17659, w17660, w17661, w17662, w17663, w17664, w17665, w17666, w17667, w17668, w17669, w17670, w17671, w17672, w17673, w17674, w17675, w17676, w17677, w17678, w17679, w17680, w17681, w17682, w17683, w17684, w17685, w17686, w17687, w17688, w17689, w17690, w17691, w17692, w17693, w17694, w17695, w17696, w17697, w17698, w17699, w17700, w17701, w17702, w17703, w17704, w17705, w17706, w17707, w17708, w17709, w17710, w17711, w17712, w17713, w17714, w17715, w17716, w17717, w17718, w17719, w17720, w17721, w17722, w17723, w17724, w17725, w17726, w17727, w17728, w17729, w17730, w17731, w17732, w17733, w17734, w17735, w17736, w17737, w17738, w17739, w17740, w17741, w17742, w17743, w17744, w17745, w17746, w17747, w17748, w17749, w17750, w17751, w17752, w17753, w17754, w17755, w17756, w17757, w17758, w17759, w17760, w17761, w17762, w17763, w17764, w17765, w17766, w17767, w17768, w17769, w17770, w17771, w17772, w17773, w17774, w17775, w17776, w17777, w17778, w17779, w17780, w17781, w17782, w17783, w17784, w17785, w17786, w17787, w17788, w17789, w17790, w17791, w17792, w17793, w17794, w17795, w17796, w17797, w17798, w17799, w17800, w17801, w17802, w17803, w17804, w17805, w17806, w17807, w17808, w17809, w17810, w17811, w17812, w17813, w17814, w17815, w17816, w17817, w17818, w17819, w17820, w17821, w17822, w17823, w17824, w17825, w17826, w17827, w17828, w17829, w17830, w17831, w17832, w17833, w17834, w17835, w17836, w17837, w17838, w17839, w17840, w17841, w17842, w17843, w17844, w17845, w17846, w17847, w17848, w17849, w17850, w17851, w17852, w17853, w17854, w17855, w17856, w17857, w17858, w17859, w17860, w17861, w17862, w17863, w17864, w17865, w17866, w17867, w17868, w17869, w17870, w17871, w17872, w17873, w17874, w17875, w17876, w17877, w17878, w17879, w17880, w17881, w17882, w17883, w17884, w17885, w17886;
assign w0 = ~pi00 & pi01;
assign v0 = ~(pi01 | pi02);
assign w1 = v0;
assign w2 = pi01 & pi02;
assign w3 = pi00 & ~w1;
assign w4 = ~w2 & w3;
assign w5 = pi02 & pi03;
assign w6 = pi00 & w5;
assign w7 = pi00 & pi03;
assign w8 = pi02 & ~w0;
assign v1 = ~(w7 | w8);
assign w9 = v1;
assign v2 = ~(w6 | w9);
assign w10 = v2;
assign w11 = pi00 & pi04;
assign w12 = pi01 & pi03;
assign v3 = ~(w11 | w12);
assign w13 = v3;
assign w14 = pi01 & pi04;
assign w15 = w7 & w14;
assign v4 = ~(w13 | w15);
assign w16 = v4;
assign v5 = ~(w2 | w16);
assign w17 = v5;
assign w18 = w2 & w16;
assign v6 = ~(w17 | w18);
assign w19 = v6;
assign w20 = w6 & ~w19;
assign w21 = ~w6 & w19;
assign v7 = ~(w20 | w21);
assign w22 = v7;
assign w23 = ~pi02 & pi03;
assign w24 = pi01 & pi05;
assign w25 = w11 & w24;
assign w26 = w15 & w25;
assign w27 = pi00 & pi05;
assign v8 = ~(w14 | w27);
assign w28 = v8;
assign v9 = ~(w15 | w25);
assign w29 = v9;
assign w30 = ~w28 & w29;
assign w31 = ~w30 & w16482;
assign w32 = (~w6 & ~w16) | (~w6 & w16483) | (~w16 & w16483);
assign v10 = ~(w17 | w32);
assign w33 = v10;
assign w34 = w31 & ~w33;
assign w35 = (w23 & w30) | (w23 & w16484) | (w30 & w16484);
assign w36 = ~w31 & w33;
assign v11 = ~(w35 | w36);
assign w37 = v11;
assign w38 = ~w34 & w37;
assign w39 = pi00 & pi06;
assign v12 = ~(w5 | w39);
assign w40 = v12;
assign w41 = w5 & w39;
assign v13 = ~(w40 | w41);
assign w42 = v13;
assign w43 = pi02 & pi04;
assign v14 = ~(w24 | w43);
assign w44 = v14;
assign w45 = w24 & w43;
assign v15 = ~(w44 | w45);
assign w46 = v15;
assign w47 = w42 & w46;
assign v16 = ~(w42 | w46);
assign w48 = v16;
assign v17 = ~(w47 | w48);
assign w49 = v17;
assign w50 = w29 & ~w49;
assign w51 = ~w29 & w49;
assign v18 = ~(w50 | w51);
assign w52 = v18;
assign w53 = w37 & w52;
assign v19 = ~(w37 | w52);
assign w54 = v19;
assign v20 = ~(w53 | w54);
assign w55 = v20;
assign v21 = ~(w41 | w47);
assign w56 = v21;
assign w57 = ~pi06 & w45;
assign w58 = pi01 & pi06;
assign v22 = ~(pi04 | w58);
assign w59 = v22;
assign w60 = pi04 & w58;
assign v23 = ~(w59 | w60);
assign w61 = v23;
assign v24 = ~(w45 | w61);
assign w62 = v24;
assign v25 = ~(w57 | w62);
assign w63 = v25;
assign w64 = ~w56 & w63;
assign w65 = w56 & ~w63;
assign v26 = ~(w64 | w65);
assign w66 = v26;
assign w67 = pi00 & pi07;
assign w68 = pi02 & pi05;
assign w69 = pi03 & pi04;
assign v27 = ~(w68 | w69);
assign w70 = v27;
assign w71 = w68 & w69;
assign v28 = ~(w70 | w71);
assign w72 = v28;
assign w73 = w67 & ~w72;
assign w74 = ~w67 & w72;
assign v29 = ~(w73 | w74);
assign w75 = v29;
assign w76 = ~w66 & w75;
assign w77 = w66 & ~w75;
assign v30 = ~(w76 | w77);
assign w78 = v30;
assign v31 = ~(w35 | w51);
assign w79 = v31;
assign w80 = (~w50 & ~w79) | (~w50 & w16485) | (~w79 & w16485);
assign w81 = w78 & w80;
assign v32 = ~(w78 | w80);
assign w82 = v32;
assign v33 = ~(w81 | w82);
assign w83 = v33;
assign v34 = ~(w57 | w64);
assign w84 = v34;
assign w85 = pi03 & pi05;
assign w86 = pi01 & pi07;
assign v35 = ~(w85 | w86);
assign w87 = v35;
assign w88 = w85 & w86;
assign v36 = ~(w87 | w88);
assign w89 = v36;
assign v37 = ~(w67 | w71);
assign w90 = v37;
assign v38 = ~(w70 | w90);
assign w91 = v38;
assign w92 = w89 & w91;
assign v39 = ~(w89 | w91);
assign w93 = v39;
assign v40 = ~(w92 | w93);
assign w94 = v40;
assign w95 = pi02 & pi06;
assign w96 = pi00 & pi08;
assign v41 = ~(w95 | w96);
assign w97 = v41;
assign w98 = pi02 & pi08;
assign w99 = w39 & w98;
assign v42 = ~(w97 | w99);
assign w100 = v42;
assign w101 = w60 & ~w100;
assign w102 = ~w60 & w100;
assign v43 = ~(w101 | w102);
assign w103 = v43;
assign w104 = w94 & ~w103;
assign w105 = ~w94 & w103;
assign v44 = ~(w104 | w105);
assign w106 = v44;
assign w107 = w84 & ~w106;
assign w108 = ~w84 & w106;
assign v45 = ~(w107 | w108);
assign w109 = v45;
assign w110 = ~w76 & w80;
assign v46 = ~(w77 | w110);
assign w111 = v46;
assign w112 = w109 & w111;
assign v47 = ~(w109 | w111);
assign w113 = v47;
assign v48 = ~(w112 | w113);
assign w114 = v48;
assign v49 = ~(w92 | w104);
assign w115 = v49;
assign w116 = pi08 & w24;
assign w117 = pi01 & pi08;
assign v50 = ~(pi05 | w117);
assign w118 = v50;
assign v51 = ~(w116 | w118);
assign w119 = v51;
assign w120 = pi00 & pi09;
assign w121 = w88 & w120;
assign v52 = ~(w88 | w120);
assign w122 = v52;
assign v53 = ~(w121 | w122);
assign w123 = v53;
assign w124 = w119 & w123;
assign v54 = ~(w119 | w123);
assign w125 = v54;
assign v55 = ~(w124 | w125);
assign w126 = v55;
assign w127 = w60 & ~w97;
assign v56 = ~(w99 | w127);
assign w128 = v56;
assign w129 = pi02 & pi07;
assign w130 = pi04 & pi05;
assign w131 = pi03 & pi06;
assign v57 = ~(w130 | w131);
assign w132 = v57;
assign w133 = w130 & w131;
assign v58 = ~(w132 | w133);
assign w134 = v58;
assign w135 = w129 & ~w134;
assign w136 = ~w129 & w134;
assign v59 = ~(w135 | w136);
assign w137 = v59;
assign v60 = ~(w128 | w137);
assign w138 = v60;
assign w139 = w128 & w137;
assign v61 = ~(w138 | w139);
assign w140 = v61;
assign w141 = w126 & w140;
assign v62 = ~(w126 | w140);
assign w142 = v62;
assign v63 = ~(w141 | w142);
assign w143 = v63;
assign w144 = ~w115 & w143;
assign w145 = w115 & ~w143;
assign v64 = ~(w144 | w145);
assign w146 = v64;
assign v65 = ~(w77 | w108);
assign w147 = v65;
assign w148 = (~w107 & ~w147) | (~w107 & w16486) | (~w147 & w16486);
assign w149 = w146 & w148;
assign v66 = ~(w146 | w148);
assign w150 = v66;
assign v67 = ~(w149 | w150);
assign w151 = v67;
assign v68 = ~(w138 | w141);
assign w152 = v68;
assign w153 = pi04 & pi06;
assign w154 = pi01 & pi09;
assign v69 = ~(w153 | w154);
assign w155 = v69;
assign w156 = w153 & w154;
assign v70 = ~(w155 | w156);
assign w157 = v70;
assign w158 = w116 & w157;
assign v71 = ~(w116 | w157);
assign w159 = v71;
assign v72 = ~(w158 | w159);
assign w160 = v72;
assign v73 = ~(w129 | w133);
assign w161 = v73;
assign v74 = ~(w132 | w161);
assign w162 = v74;
assign w163 = w160 & w162;
assign v75 = ~(w160 | w162);
assign w164 = v75;
assign v76 = ~(w163 | w164);
assign w165 = v76;
assign w166 = (~w121 & ~w123) | (~w121 & w16487) | (~w123 & w16487);
assign w167 = pi03 & pi07;
assign w168 = pi00 & pi10;
assign v77 = ~(w167 | w168);
assign w169 = v77;
assign w170 = w167 & w168;
assign v78 = ~(w169 | w170);
assign w171 = v78;
assign w172 = w98 & ~w171;
assign w173 = ~w98 & w171;
assign v79 = ~(w172 | w173);
assign w174 = v79;
assign v80 = ~(w166 | w174);
assign w175 = v80;
assign w176 = w166 & w174;
assign v81 = ~(w175 | w176);
assign w177 = v81;
assign w178 = w165 & w177;
assign v82 = ~(w165 | w177);
assign w179 = v82;
assign v83 = ~(w178 | w179);
assign w180 = v83;
assign w181 = ~w152 & w180;
assign w182 = w152 & ~w180;
assign v84 = ~(w181 | w182);
assign w183 = v84;
assign v85 = ~(w144 | w148);
assign w184 = v85;
assign v86 = ~(w145 | w184);
assign w185 = v86;
assign w186 = w183 & w185;
assign v87 = ~(w183 | w185);
assign w187 = v87;
assign v88 = ~(w186 | w187);
assign w188 = v88;
assign v89 = ~(w175 | w178);
assign w189 = v89;
assign w190 = pi10 & w58;
assign w191 = pi01 & pi10;
assign v90 = ~(pi06 | w191);
assign w192 = v90;
assign v91 = ~(w190 | w192);
assign w193 = v91;
assign v92 = ~(w98 | w170);
assign w194 = v92;
assign v93 = ~(w169 | w194);
assign w195 = v93;
assign w196 = w193 & w195;
assign v94 = ~(w193 | w195);
assign w197 = v94;
assign v95 = ~(w196 | w197);
assign w198 = v95;
assign w199 = pi03 & pi08;
assign w200 = pi02 & pi09;
assign v96 = ~(w199 | w200);
assign w201 = v96;
assign w202 = w199 & w200;
assign v97 = ~(w201 | w202);
assign w203 = v97;
assign w204 = w156 & ~w203;
assign w205 = ~w156 & w203;
assign v98 = ~(w204 | w205);
assign w206 = v98;
assign w207 = w198 & ~w206;
assign w208 = ~w198 & w206;
assign v99 = ~(w207 | w208);
assign w209 = v99;
assign w210 = (~w158 & ~w160) | (~w158 & w16488) | (~w160 & w16488);
assign w211 = pi00 & pi11;
assign w212 = pi05 & pi06;
assign w213 = pi04 & pi07;
assign v100 = ~(w212 | w213);
assign w214 = v100;
assign w215 = w212 & w213;
assign v101 = ~(w214 | w215);
assign w216 = v101;
assign w217 = w211 & ~w216;
assign w218 = ~w211 & w216;
assign v102 = ~(w217 | w218);
assign w219 = v102;
assign v103 = ~(w210 | w219);
assign w220 = v103;
assign w221 = w210 & w219;
assign v104 = ~(w220 | w221);
assign w222 = v104;
assign w223 = w209 & w222;
assign v105 = ~(w209 | w222);
assign w224 = v105;
assign v106 = ~(w223 | w224);
assign w225 = v106;
assign w226 = w189 & ~w225;
assign w227 = ~w189 & w225;
assign v107 = ~(w226 | w227);
assign w228 = v107;
assign v108 = ~(w145 | w182);
assign w229 = v108;
assign w230 = ~w184 & w229;
assign v109 = ~(w181 | w230);
assign w231 = v109;
assign w232 = w228 & w231;
assign v110 = ~(w228 | w231);
assign w233 = v110;
assign v111 = ~(w232 | w233);
assign w234 = v111;
assign v112 = ~(w181 | w227);
assign w235 = v112;
assign w236 = (~w226 & w230) | (~w226 & w16489) | (w230 & w16489);
assign v113 = ~(w220 | w223);
assign w237 = v113;
assign v114 = ~(w211 | w215);
assign w238 = v114;
assign v115 = ~(w214 | w238);
assign w239 = v115;
assign v116 = ~(w156 | w202);
assign w240 = v116;
assign v117 = ~(w201 | w240);
assign w241 = v117;
assign w242 = w239 & w241;
assign v118 = ~(w239 | w241);
assign w243 = v118;
assign v119 = ~(w242 | w243);
assign w244 = v119;
assign w245 = pi03 & pi09;
assign w246 = pi00 & pi12;
assign w247 = pi02 & pi10;
assign v120 = ~(w246 | w247);
assign w248 = v120;
assign w249 = pi02 & pi12;
assign w250 = w168 & w249;
assign v121 = ~(w248 | w250);
assign w251 = v121;
assign w252 = w245 & ~w251;
assign w253 = ~w245 & w251;
assign v122 = ~(w252 | w253);
assign w254 = v122;
assign w255 = ~w244 & w254;
assign w256 = w244 & ~w254;
assign v123 = ~(w255 | w256);
assign w257 = v123;
assign w258 = (~w196 & ~w198) | (~w196 & w16490) | (~w198 & w16490);
assign w259 = pi05 & pi07;
assign w260 = pi01 & pi11;
assign v124 = ~(w259 | w260);
assign w261 = v124;
assign w262 = w259 & w260;
assign v125 = ~(w261 | w262);
assign w263 = v125;
assign w264 = pi04 & pi08;
assign v126 = ~(w190 | w264);
assign w265 = v126;
assign w266 = w190 & w264;
assign v127 = ~(w265 | w266);
assign w267 = v127;
assign w268 = w263 & ~w267;
assign w269 = ~w263 & w267;
assign v128 = ~(w268 | w269);
assign w270 = v128;
assign v129 = ~(w258 | w270);
assign w271 = v129;
assign w272 = w258 & w270;
assign v130 = ~(w271 | w272);
assign w273 = v130;
assign w274 = w257 & w273;
assign v131 = ~(w257 | w273);
assign w275 = v131;
assign v132 = ~(w274 | w275);
assign w276 = v132;
assign w277 = w237 & ~w276;
assign w278 = ~w237 & w276;
assign v133 = ~(w277 | w278);
assign w279 = v133;
assign w280 = w236 & ~w279;
assign w281 = ~w236 & w279;
assign v134 = ~(w280 | w281);
assign w282 = v134;
assign v135 = ~(w236 | w278);
assign w283 = v135;
assign v136 = ~(w277 | w283);
assign w284 = v136;
assign v137 = ~(w242 | w256);
assign w285 = v137;
assign w286 = ~pi12 & w262;
assign w287 = pi12 & w86;
assign w288 = pi01 & pi12;
assign v138 = ~(pi07 | w288);
assign w289 = v138;
assign v139 = ~(w287 | w289);
assign w290 = v139;
assign v140 = ~(w262 | w290);
assign w291 = v140;
assign v141 = ~(w286 | w291);
assign w292 = v141;
assign w293 = w245 & ~w248;
assign v142 = ~(w250 | w293);
assign w294 = v142;
assign w295 = ~w292 & w294;
assign w296 = w292 & ~w294;
assign v143 = ~(w295 | w296);
assign w297 = v143;
assign w298 = ~w285 & w297;
assign w299 = w285 & ~w297;
assign v144 = ~(w298 | w299);
assign w300 = v144;
assign w301 = (~w271 & ~w273) | (~w271 & w16491) | (~w273 & w16491);
assign w302 = ~w300 & w301;
assign w303 = w300 & ~w301;
assign v145 = ~(w302 | w303);
assign w304 = v145;
assign w305 = pi03 & pi10;
assign w306 = pi04 & pi09;
assign w307 = pi00 & pi13;
assign v146 = ~(w306 | w307);
assign w308 = v146;
assign w309 = w306 & w307;
assign v147 = ~(w308 | w309);
assign w310 = v147;
assign w311 = w305 & ~w310;
assign w312 = ~w305 & w310;
assign v148 = ~(w311 | w312);
assign w313 = v148;
assign w314 = w263 & ~w265;
assign v149 = ~(w266 | w314);
assign w315 = v149;
assign v150 = ~(w313 | w315);
assign w316 = v150;
assign w317 = w313 & w315;
assign v151 = ~(w316 | w317);
assign w318 = v151;
assign w319 = pi02 & pi11;
assign w320 = pi06 & pi07;
assign w321 = pi05 & pi08;
assign v152 = ~(w320 | w321);
assign w322 = v152;
assign w323 = w320 & w321;
assign v153 = ~(w322 | w323);
assign w324 = v153;
assign w325 = w319 & ~w324;
assign w326 = ~w319 & w324;
assign v154 = ~(w325 | w326);
assign w327 = v154;
assign w328 = w318 & ~w327;
assign w329 = ~w318 & w327;
assign v155 = ~(w328 | w329);
assign w330 = v155;
assign v156 = ~(w304 | w330);
assign w331 = v156;
assign w332 = w304 & w330;
assign v157 = ~(w331 | w332);
assign w333 = v157;
assign w334 = w284 & w333;
assign v158 = ~(w284 | w333);
assign w335 = v158;
assign v159 = ~(w334 | w335);
assign w336 = v159;
assign v160 = ~(w277 | w331);
assign w337 = v160;
assign w338 = ~w283 & w337;
assign v161 = ~(w332 | w338);
assign w339 = v161;
assign v162 = ~(w298 | w303);
assign w340 = v162;
assign w341 = pi04 & pi10;
assign w342 = pi05 & pi09;
assign v163 = ~(w341 | w342);
assign w343 = v163;
assign w344 = w341 & w342;
assign v164 = ~(w343 | w344);
assign w345 = v164;
assign w346 = w287 & ~w345;
assign w347 = ~w287 & w345;
assign v165 = ~(w346 | w347);
assign w348 = v165;
assign w349 = pi00 & pi14;
assign w350 = pi03 & pi11;
assign v166 = ~(w249 | w350);
assign w351 = v166;
assign w352 = w249 & w350;
assign v167 = ~(w351 | w352);
assign w353 = v167;
assign w354 = w349 & ~w353;
assign w355 = ~w349 & w353;
assign v168 = ~(w354 | w355);
assign w356 = v168;
assign v169 = ~(w348 | w356);
assign w357 = v169;
assign w358 = w348 & w356;
assign v170 = ~(w357 | w358);
assign w359 = v170;
assign w360 = (~w286 & ~w292) | (~w286 & w16807) | (~w292 & w16807);
assign w361 = ~w359 & w360;
assign w362 = w359 & ~w360;
assign v171 = ~(w361 | w362);
assign w363 = v171;
assign w364 = (~w316 & ~w318) | (~w316 & w16697) | (~w318 & w16697);
assign w365 = pi06 & pi08;
assign w366 = pi01 & pi13;
assign v172 = ~(w365 | w366);
assign w367 = v172;
assign w368 = w365 & w366;
assign v173 = ~(w367 | w368);
assign w369 = v173;
assign v174 = ~(w319 | w323);
assign w370 = v174;
assign v175 = ~(w322 | w370);
assign w371 = v175;
assign w372 = w369 & w371;
assign v176 = ~(w369 | w371);
assign w373 = v176;
assign v177 = ~(w372 | w373);
assign w374 = v177;
assign v178 = ~(w305 | w309);
assign w375 = v178;
assign v179 = ~(w308 | w375);
assign w376 = v179;
assign w377 = w374 & w376;
assign v180 = ~(w374 | w376);
assign w378 = v180;
assign v181 = ~(w377 | w378);
assign w379 = v181;
assign w380 = ~w364 & w379;
assign w381 = w364 & ~w379;
assign v182 = ~(w380 | w381);
assign w382 = v182;
assign w383 = w363 & w382;
assign v183 = ~(w363 | w382);
assign w384 = v183;
assign v184 = ~(w383 | w384);
assign w385 = v184;
assign w386 = ~w340 & w385;
assign w387 = w340 & ~w385;
assign v185 = ~(w386 | w387);
assign w388 = v185;
assign w389 = w339 & w388;
assign v186 = ~(w339 | w388);
assign w390 = v186;
assign v187 = ~(w389 | w390);
assign w391 = v187;
assign v188 = ~(w332 | w386);
assign w392 = v188;
assign w393 = (~w387 & w338) | (~w387 & w16492) | (w338 & w16492);
assign v189 = ~(w380 | w383);
assign w394 = v189;
assign w395 = (~w372 & ~w374) | (~w372 & w16698) | (~w374 & w16698);
assign w396 = pi04 & pi11;
assign v190 = ~(w368 | w396);
assign w397 = v190;
assign w398 = w368 & w396;
assign v191 = ~(w397 | w398);
assign w399 = v191;
assign w400 = pi01 & pi14;
assign w401 = pi08 & w400;
assign v192 = ~(pi08 | w400);
assign w402 = v192;
assign v193 = ~(w401 | w402);
assign w403 = v193;
assign w404 = ~w399 & w403;
assign w405 = w399 & ~w403;
assign v194 = ~(w404 | w405);
assign w406 = v194;
assign w407 = pi02 & pi13;
assign w408 = pi06 & pi09;
assign w409 = pi07 & pi08;
assign v195 = ~(w408 | w409);
assign w410 = v195;
assign w411 = w408 & w409;
assign v196 = ~(w410 | w411);
assign w412 = v196;
assign w413 = w407 & ~w412;
assign w414 = ~w407 & w412;
assign v197 = ~(w413 | w414);
assign w415 = v197;
assign v198 = ~(w406 | w415);
assign w416 = v198;
assign w417 = w406 & w415;
assign v199 = ~(w416 | w417);
assign w418 = v199;
assign w419 = w395 & ~w418;
assign w420 = ~w395 & w418;
assign v200 = ~(w419 | w420);
assign w421 = v200;
assign v201 = ~(w349 | w352);
assign w422 = v201;
assign v202 = ~(w351 | w422);
assign w423 = v202;
assign v203 = ~(w287 | w344);
assign w424 = v203;
assign v204 = ~(w343 | w424);
assign w425 = v204;
assign w426 = w423 & w425;
assign v205 = ~(w423 | w425);
assign w427 = v205;
assign v206 = ~(w426 | w427);
assign w428 = v206;
assign w429 = pi05 & pi10;
assign w430 = pi03 & pi12;
assign w431 = pi00 & pi15;
assign v207 = ~(w430 | w431);
assign w432 = v207;
assign w433 = w430 & w431;
assign v208 = ~(w432 | w433);
assign w434 = v208;
assign w435 = w429 & ~w434;
assign w436 = ~w429 & w434;
assign v209 = ~(w435 | w436);
assign w437 = v209;
assign w438 = ~w428 & w437;
assign w439 = w428 & ~w437;
assign v210 = ~(w438 | w439);
assign w440 = v210;
assign w441 = (~w357 & ~w359) | (~w357 & w16808) | (~w359 & w16808);
assign w442 = w440 & ~w441;
assign w443 = ~w440 & w441;
assign v211 = ~(w442 | w443);
assign w444 = v211;
assign w445 = w421 & w444;
assign v212 = ~(w421 | w444);
assign w446 = v212;
assign v213 = ~(w445 | w446);
assign w447 = v213;
assign w448 = ~w394 & w447;
assign w449 = w394 & ~w447;
assign v214 = ~(w448 | w449);
assign w450 = v214;
assign w451 = w393 & ~w450;
assign w452 = ~w393 & w450;
assign v215 = ~(w451 | w452);
assign w453 = v215;
assign v216 = ~(w442 | w445);
assign w454 = v216;
assign v217 = ~(w429 | w433);
assign w455 = v217;
assign v218 = ~(w432 | w455);
assign w456 = v218;
assign v219 = ~(w398 | w403);
assign w457 = v219;
assign v220 = ~(w397 | w457);
assign w458 = v220;
assign w459 = w456 & w458;
assign v221 = ~(w456 | w458);
assign w460 = v221;
assign v222 = ~(w459 | w460);
assign w461 = v222;
assign w462 = pi05 & pi11;
assign w463 = pi00 & pi16;
assign w464 = pi06 & pi10;
assign v223 = ~(w463 | w464);
assign w465 = v223;
assign w466 = w463 & w464;
assign v224 = ~(w465 | w466);
assign w467 = v224;
assign w468 = w462 & ~w467;
assign w469 = ~w462 & w467;
assign v225 = ~(w468 | w469);
assign w470 = v225;
assign w471 = ~w461 & w470;
assign w472 = w461 & ~w470;
assign v226 = ~(w471 | w472);
assign w473 = v226;
assign w474 = (~w416 & ~w418) | (~w416 & w16699) | (~w418 & w16699);
assign w475 = w473 & ~w474;
assign w476 = ~w473 & w474;
assign v227 = ~(w475 | w476);
assign w477 = v227;
assign w478 = pi07 & pi09;
assign w479 = pi01 & pi15;
assign v228 = ~(w478 | w479);
assign w480 = v228;
assign w481 = w478 & w479;
assign v229 = ~(w480 | w481);
assign w482 = v229;
assign w483 = w401 & w482;
assign v230 = ~(w401 | w482);
assign w484 = v230;
assign v231 = ~(w483 | w484);
assign w485 = v231;
assign v232 = ~(w407 | w411);
assign w486 = v232;
assign v233 = ~(w410 | w486);
assign w487 = v233;
assign w488 = w485 & w487;
assign v234 = ~(w485 | w487);
assign w489 = v234;
assign v235 = ~(w488 | w489);
assign w490 = v235;
assign w491 = (~w426 & ~w428) | (~w426 & w16700) | (~w428 & w16700);
assign w492 = pi04 & pi12;
assign w493 = pi03 & pi13;
assign w494 = pi02 & pi14;
assign v236 = ~(w493 | w494);
assign w495 = v236;
assign w496 = w493 & w494;
assign v237 = ~(w495 | w496);
assign w497 = v237;
assign w498 = w492 & ~w497;
assign w499 = ~w492 & w497;
assign v238 = ~(w498 | w499);
assign w500 = v238;
assign v239 = ~(w491 | w500);
assign w501 = v239;
assign w502 = w491 & w500;
assign v240 = ~(w501 | w502);
assign w503 = v240;
assign w504 = w490 & w503;
assign v241 = ~(w490 | w503);
assign w505 = v241;
assign v242 = ~(w504 | w505);
assign w506 = v242;
assign v243 = ~(w477 | w506);
assign w507 = v243;
assign w508 = w477 & w506;
assign v244 = ~(w507 | w508);
assign w509 = v244;
assign w510 = ~w454 & w509;
assign w511 = w454 & ~w509;
assign v245 = ~(w510 | w511);
assign w512 = v245;
assign v246 = ~(w393 | w448);
assign w513 = v246;
assign v247 = ~(w449 | w513);
assign w514 = v247;
assign w515 = w512 & w514;
assign v248 = ~(w512 | w514);
assign w516 = v248;
assign v249 = ~(w515 | w516);
assign w517 = v249;
assign v250 = ~(w475 | w508);
assign w518 = v250;
assign w519 = pi01 & pi16;
assign v251 = ~(pi09 | w519);
assign w520 = v251;
assign w521 = pi16 & w154;
assign v252 = ~(w520 | w521);
assign w522 = v252;
assign v253 = ~(w492 | w496);
assign w523 = v253;
assign v254 = ~(w495 | w523);
assign w524 = v254;
assign w525 = w522 & w524;
assign v255 = ~(w522 | w524);
assign w526 = v255;
assign v256 = ~(w525 | w526);
assign w527 = v256;
assign v257 = ~(w462 | w466);
assign w528 = v257;
assign v258 = ~(w465 | w528);
assign w529 = v258;
assign w530 = w527 & w529;
assign v259 = ~(w527 | w529);
assign w531 = v259;
assign v260 = ~(w530 | w531);
assign w532 = v260;
assign v261 = ~(w483 | w488);
assign w533 = v261;
assign w534 = (~w459 & ~w461) | (~w459 & w16701) | (~w461 & w16701);
assign v262 = ~(w533 | w534);
assign w535 = v262;
assign w536 = w533 & w534;
assign v263 = ~(w535 | w536);
assign w537 = v263;
assign v264 = ~(w532 | w537);
assign w538 = v264;
assign w539 = w532 & w537;
assign v265 = ~(w538 | w539);
assign w540 = v265;
assign w541 = (~w501 & ~w503) | (~w501 & w16809) | (~w503 & w16809);
assign w542 = pi05 & pi12;
assign w543 = pi00 & pi17;
assign v266 = ~(w542 | w543);
assign w544 = v266;
assign w545 = w542 & w543;
assign v267 = ~(w544 | w545);
assign w546 = v267;
assign w547 = w481 & ~w546;
assign w548 = ~w481 & w546;
assign v268 = ~(w547 | w548);
assign w549 = v268;
assign w550 = pi03 & pi14;
assign w551 = pi07 & pi10;
assign w552 = pi08 & pi09;
assign v269 = ~(w551 | w552);
assign w553 = v269;
assign w554 = w551 & w552;
assign v270 = ~(w553 | w554);
assign w555 = v270;
assign w556 = w550 & ~w555;
assign w557 = ~w550 & w555;
assign v271 = ~(w556 | w557);
assign w558 = v271;
assign v272 = ~(w549 | w558);
assign w559 = v272;
assign w560 = w549 & w558;
assign v273 = ~(w559 | w560);
assign w561 = v273;
assign w562 = pi06 & pi11;
assign w563 = pi04 & pi13;
assign w564 = pi02 & pi15;
assign v274 = ~(w563 | w564);
assign w565 = v274;
assign w566 = w563 & w564;
assign v275 = ~(w565 | w566);
assign w567 = v275;
assign w568 = w562 & ~w567;
assign w569 = ~w562 & w567;
assign v276 = ~(w568 | w569);
assign w570 = v276;
assign w571 = w561 & ~w570;
assign w572 = ~w561 & w570;
assign v277 = ~(w571 | w572);
assign w573 = v277;
assign w574 = ~w541 & w573;
assign w575 = w541 & ~w573;
assign v278 = ~(w574 | w575);
assign w576 = v278;
assign w577 = w540 & w576;
assign v279 = ~(w540 | w576);
assign w578 = v279;
assign v280 = ~(w577 | w578);
assign w579 = v280;
assign w580 = ~w518 & w579;
assign w581 = w518 & ~w579;
assign v281 = ~(w580 | w581);
assign w582 = v281;
assign v282 = ~(w449 | w511);
assign w583 = v282;
assign w584 = (w338 & w16810) | (w338 & w16811) | (w16810 & w16811);
assign v283 = ~(w510 | w584);
assign w585 = v283;
assign w586 = w582 & w585;
assign v284 = ~(w582 | w585);
assign w587 = v284;
assign v285 = ~(w586 | w587);
assign w588 = v285;
assign w589 = (~w510 & ~w579) | (~w510 & w16494) | (~w579 & w16494);
assign w590 = (~w581 & w584) | (~w581 & w16495) | (w584 & w16495);
assign v286 = ~(w574 | w577);
assign w591 = v286;
assign v287 = ~(w481 | w545);
assign w592 = v287;
assign v288 = ~(w544 | w592);
assign w593 = v288;
assign v289 = ~(w550 | w554);
assign w594 = v289;
assign v290 = ~(w553 | w594);
assign w595 = v290;
assign v291 = ~(w562 | w566);
assign w596 = v291;
assign v292 = ~(w565 | w596);
assign w597 = v292;
assign w598 = w595 & w597;
assign v293 = ~(w595 | w597);
assign w599 = v293;
assign v294 = ~(w598 | w599);
assign w600 = v294;
assign v295 = ~(w593 | w600);
assign w601 = v295;
assign w602 = w593 & w600;
assign v296 = ~(w601 | w602);
assign w603 = v296;
assign w604 = (~w525 & ~w527) | (~w525 & w16812) | (~w527 & w16812);
assign w605 = (~w559 & ~w561) | (~w559 & w16702) | (~w561 & w16702);
assign v297 = ~(w604 | w605);
assign w606 = v297;
assign w607 = w604 & w605;
assign v298 = ~(w606 | w607);
assign w608 = v298;
assign w609 = w603 & w608;
assign v299 = ~(w603 | w608);
assign w610 = v299;
assign v300 = ~(w609 | w610);
assign w611 = v300;
assign w612 = (~w535 & ~w537) | (~w535 & w16813) | (~w537 & w16813);
assign w613 = pi07 & pi11;
assign w614 = pi00 & pi18;
assign w615 = pi05 & pi13;
assign v301 = ~(w614 | w615);
assign w616 = v301;
assign w617 = w614 & w615;
assign v302 = ~(w616 | w617);
assign w618 = v302;
assign w619 = w613 & ~w618;
assign w620 = ~w613 & w618;
assign v303 = ~(w619 | w620);
assign w621 = v303;
assign w622 = pi04 & pi14;
assign w623 = pi03 & pi15;
assign w624 = pi02 & pi16;
assign v304 = ~(w623 | w624);
assign w625 = v304;
assign w626 = w623 & w624;
assign v305 = ~(w625 | w626);
assign w627 = v305;
assign w628 = w622 & ~w627;
assign w629 = ~w622 & w627;
assign v306 = ~(w628 | w629);
assign w630 = v306;
assign v307 = ~(w621 | w630);
assign w631 = v307;
assign w632 = w621 & w630;
assign v308 = ~(w631 | w632);
assign w633 = v308;
assign w634 = pi06 & pi12;
assign v309 = ~(w521 | w634);
assign w635 = v309;
assign w636 = w521 & w634;
assign v310 = ~(w635 | w636);
assign w637 = v310;
assign w638 = pi08 & pi10;
assign w639 = pi01 & pi17;
assign v311 = ~(w638 | w639);
assign w640 = v311;
assign w641 = w638 & w639;
assign v312 = ~(w640 | w641);
assign w642 = v312;
assign w643 = ~w637 & w642;
assign w644 = w637 & ~w642;
assign v313 = ~(w643 | w644);
assign w645 = v313;
assign w646 = w633 & ~w645;
assign w647 = ~w633 & w645;
assign v314 = ~(w646 | w647);
assign w648 = v314;
assign w649 = ~w612 & w648;
assign w650 = w612 & ~w648;
assign v315 = ~(w649 | w650);
assign w651 = v315;
assign w652 = w611 & w651;
assign v316 = ~(w611 | w651);
assign w653 = v316;
assign v317 = ~(w652 | w653);
assign w654 = v317;
assign w655 = w591 & ~w654;
assign w656 = ~w591 & w654;
assign v318 = ~(w655 | w656);
assign w657 = v318;
assign w658 = w590 & ~w657;
assign w659 = ~w590 & w657;
assign v319 = ~(w658 | w659);
assign w660 = v319;
assign w661 = (~w584 & w16703) | (~w584 & w16704) | (w16703 & w16704);
assign v320 = ~(w655 | w661);
assign w662 = v320;
assign v321 = ~(w613 | w617);
assign w663 = v321;
assign v322 = ~(w616 | w663);
assign w664 = v322;
assign v323 = ~(w636 | w642);
assign w665 = v323;
assign v324 = ~(w635 | w665);
assign w666 = v324;
assign w667 = w664 & w666;
assign v325 = ~(w664 | w666);
assign w668 = v325;
assign v326 = ~(w667 | w668);
assign w669 = v326;
assign w670 = pi03 & pi16;
assign w671 = pi09 & pi10;
assign w672 = pi08 & pi11;
assign v327 = ~(w671 | w672);
assign w673 = v327;
assign w674 = w671 & w672;
assign v328 = ~(w673 | w674);
assign w675 = v328;
assign w676 = w670 & ~w675;
assign w677 = ~w670 & w675;
assign v329 = ~(w676 | w677);
assign w678 = v329;
assign w679 = ~w669 & w678;
assign w680 = w669 & ~w678;
assign v330 = ~(w679 | w680);
assign w681 = v330;
assign w682 = (~w631 & ~w633) | (~w631 & w16705) | (~w633 & w16705);
assign w683 = ~pi18 & w641;
assign w684 = pi01 & pi18;
assign v331 = ~(pi10 | w684);
assign w685 = v331;
assign w686 = pi10 & w684;
assign v332 = ~(w685 | w686);
assign w687 = v332;
assign v333 = ~(w641 | w687);
assign w688 = v333;
assign v334 = ~(w683 | w688);
assign w689 = v334;
assign v335 = ~(w622 | w626);
assign w690 = v335;
assign v336 = ~(w625 | w690);
assign w691 = v336;
assign w692 = w689 & w691;
assign v337 = ~(w689 | w691);
assign w693 = v337;
assign v338 = ~(w692 | w693);
assign w694 = v338;
assign w695 = ~w682 & w694;
assign w696 = w682 & ~w694;
assign v339 = ~(w695 | w696);
assign w697 = v339;
assign w698 = w681 & w697;
assign v340 = ~(w681 | w697);
assign w699 = v340;
assign v341 = ~(w698 | w699);
assign w700 = v341;
assign w701 = (~w598 & ~w600) | (~w598 & w16814) | (~w600 & w16814);
assign w702 = pi00 & pi19;
assign w703 = pi04 & pi15;
assign w704 = pi02 & pi17;
assign v342 = ~(w703 | w704);
assign w705 = v342;
assign w706 = w703 & w704;
assign v343 = ~(w705 | w706);
assign w707 = v343;
assign w708 = w702 & ~w707;
assign w709 = ~w702 & w707;
assign v344 = ~(w708 | w709);
assign w710 = v344;
assign w711 = pi05 & pi14;
assign w712 = pi06 & pi13;
assign w713 = pi07 & pi12;
assign v345 = ~(w712 | w713);
assign w714 = v345;
assign w715 = w712 & w713;
assign v346 = ~(w714 | w715);
assign w716 = v346;
assign w717 = w711 & ~w716;
assign w718 = ~w711 & w716;
assign v347 = ~(w717 | w718);
assign w719 = v347;
assign v348 = ~(w710 | w719);
assign w720 = v348;
assign w721 = w710 & w719;
assign v349 = ~(w720 | w721);
assign w722 = v349;
assign w723 = w701 & ~w722;
assign w724 = ~w701 & w722;
assign v350 = ~(w723 | w724);
assign w725 = v350;
assign w726 = (~w606 & ~w608) | (~w606 & w16815) | (~w608 & w16815);
assign w727 = ~w725 & w726;
assign w728 = w725 & ~w726;
assign v351 = ~(w727 | w728);
assign w729 = v351;
assign w730 = w700 & w729;
assign v352 = ~(w700 | w729);
assign w731 = v352;
assign v353 = ~(w730 | w731);
assign w732 = v353;
assign w733 = (~w649 & ~w651) | (~w649 & w17025) | (~w651 & w17025);
assign w734 = ~w732 & w733;
assign w735 = w732 & ~w733;
assign v354 = ~(w734 | w735);
assign w736 = v354;
assign w737 = w662 & w736;
assign v355 = ~(w662 | w736);
assign w738 = v355;
assign v356 = ~(w737 | w738);
assign w739 = v356;
assign v357 = ~(w655 | w734);
assign w740 = v357;
assign w741 = ~w661 & w740;
assign v358 = ~(w735 | w741);
assign w742 = v358;
assign w743 = (~w728 & ~w729) | (~w728 & w17026) | (~w729 & w17026);
assign w744 = (~w667 & ~w669) | (~w667 & w16816) | (~w669 & w16816);
assign w745 = (~w683 & ~w689) | (~w683 & w16817) | (~w689 & w16817);
assign w746 = pi02 & pi18;
assign w747 = pi03 & pi17;
assign w748 = pi04 & pi16;
assign v359 = ~(w747 | w748);
assign w749 = v359;
assign w750 = w747 & w748;
assign v360 = ~(w749 | w750);
assign w751 = v360;
assign w752 = w746 & ~w751;
assign w753 = ~w746 & w751;
assign v361 = ~(w752 | w753);
assign w754 = v361;
assign v362 = ~(w745 | w754);
assign w755 = v362;
assign w756 = w745 & w754;
assign v363 = ~(w755 | w756);
assign w757 = v363;
assign w758 = w744 & ~w757;
assign w759 = ~w744 & w757;
assign v364 = ~(w758 | w759);
assign w760 = v364;
assign w761 = (~w695 & ~w697) | (~w695 & w16818) | (~w697 & w16818);
assign w762 = ~w760 & w761;
assign w763 = w760 & ~w761;
assign v365 = ~(w762 | w763);
assign w764 = v365;
assign v366 = ~(w711 | w715);
assign w765 = v366;
assign v367 = ~(w714 | w765);
assign w766 = v367;
assign w767 = pi07 & pi13;
assign w768 = pi00 & pi20;
assign v368 = ~(w767 | w768);
assign w769 = v368;
assign w770 = w767 & w768;
assign v369 = ~(w769 | w770);
assign w771 = v369;
assign w772 = w686 & ~w771;
assign w773 = ~w686 & w771;
assign v370 = ~(w772 | w773);
assign w774 = v370;
assign w775 = w766 & ~w774;
assign w776 = ~w766 & w774;
assign v371 = ~(w775 | w776);
assign w777 = v371;
assign w778 = pi08 & pi12;
assign w779 = pi05 & pi15;
assign w780 = pi06 & pi14;
assign v372 = ~(w779 | w780);
assign w781 = v372;
assign w782 = w779 & w780;
assign v373 = ~(w781 | w782);
assign w783 = v373;
assign w784 = w778 & ~w783;
assign w785 = ~w778 & w783;
assign v374 = ~(w784 | w785);
assign w786 = v374;
assign w787 = ~w777 & w786;
assign w788 = w777 & ~w786;
assign v375 = ~(w787 | w788);
assign w789 = v375;
assign v376 = ~(w720 | w724);
assign w790 = v376;
assign w791 = pi09 & pi11;
assign w792 = pi01 & pi19;
assign v377 = ~(w791 | w792);
assign w793 = v377;
assign w794 = w791 & w792;
assign v378 = ~(w793 | w794);
assign w795 = v378;
assign v379 = ~(w670 | w674);
assign w796 = v379;
assign v380 = ~(w673 | w796);
assign w797 = v380;
assign w798 = w795 & w797;
assign v381 = ~(w795 | w797);
assign w799 = v381;
assign v382 = ~(w798 | w799);
assign w800 = v382;
assign v383 = ~(w702 | w706);
assign w801 = v383;
assign v384 = ~(w705 | w801);
assign w802 = v384;
assign w803 = w800 & w802;
assign v385 = ~(w800 | w802);
assign w804 = v385;
assign v386 = ~(w803 | w804);
assign w805 = v386;
assign w806 = ~w790 & w805;
assign w807 = w790 & ~w805;
assign v387 = ~(w806 | w807);
assign w808 = v387;
assign w809 = w789 & w808;
assign v388 = ~(w789 | w808);
assign w810 = v388;
assign v389 = ~(w809 | w810);
assign w811 = v389;
assign w812 = w764 & w811;
assign v390 = ~(w764 | w811);
assign w813 = v390;
assign v391 = ~(w812 | w813);
assign w814 = v391;
assign w815 = ~w743 & w814;
assign w816 = w743 & ~w814;
assign v392 = ~(w815 | w816);
assign w817 = v392;
assign w818 = w742 & w817;
assign v393 = ~(w742 | w817);
assign w819 = v393;
assign v394 = ~(w818 | w819);
assign w820 = v394;
assign v395 = ~(w763 | w812);
assign w821 = v395;
assign v396 = ~(w746 | w750);
assign w822 = v396;
assign v397 = ~(w749 | w822);
assign w823 = v397;
assign v398 = ~(w778 | w782);
assign w824 = v398;
assign v399 = ~(w781 | w824);
assign w825 = v399;
assign w826 = w823 & w825;
assign v400 = ~(w823 | w825);
assign w827 = v400;
assign v401 = ~(w826 | w827);
assign w828 = v401;
assign v402 = ~(w686 | w770);
assign w829 = v402;
assign v403 = ~(w769 | w829);
assign w830 = v403;
assign v404 = ~(w828 | w830);
assign w831 = v404;
assign w832 = w828 & w830;
assign v405 = ~(w831 | w832);
assign w833 = v405;
assign w834 = ~w759 & w17027;
assign w835 = (w833 & w759) | (w833 & w17028) | (w759 & w17028);
assign v406 = ~(w834 | w835);
assign w836 = v406;
assign w837 = pi06 & pi15;
assign w838 = pi08 & pi13;
assign w839 = pi07 & pi14;
assign v407 = ~(w838 | w839);
assign w840 = v407;
assign w841 = w838 & w839;
assign v408 = ~(w840 | w841);
assign w842 = v408;
assign w843 = w837 & ~w842;
assign w844 = ~w837 & w842;
assign v409 = ~(w843 | w844);
assign w845 = v409;
assign w846 = pi05 & pi16;
assign w847 = pi02 & pi19;
assign w848 = pi03 & pi18;
assign v410 = ~(w847 | w848);
assign w849 = v410;
assign w850 = w847 & w848;
assign v411 = ~(w849 | w850);
assign w851 = v411;
assign w852 = w846 & ~w851;
assign w853 = ~w846 & w851;
assign v412 = ~(w852 | w853);
assign w854 = v412;
assign v413 = ~(w845 | w854);
assign w855 = v413;
assign w856 = w845 & w854;
assign v414 = ~(w855 | w856);
assign w857 = v414;
assign w858 = pi04 & pi17;
assign w859 = pi10 & pi11;
assign w860 = pi09 & pi12;
assign v415 = ~(w859 | w860);
assign w861 = v415;
assign w862 = w859 & w860;
assign v416 = ~(w861 | w862);
assign w863 = v416;
assign w864 = w858 & ~w863;
assign w865 = ~w858 & w863;
assign v417 = ~(w864 | w865);
assign w866 = v417;
assign w867 = w857 & ~w866;
assign w868 = ~w857 & w866;
assign v418 = ~(w867 | w868);
assign w869 = v418;
assign v419 = ~(w836 | w869);
assign w870 = v419;
assign w871 = w836 & w869;
assign v420 = ~(w870 | w871);
assign w872 = v420;
assign w873 = (~w798 & ~w800) | (~w798 & w16706) | (~w800 & w16706);
assign w874 = pi00 & pi21;
assign w875 = w794 & w874;
assign v421 = ~(w794 | w874);
assign w876 = v421;
assign v422 = ~(w875 | w876);
assign w877 = v422;
assign w878 = pi01 & pi20;
assign w879 = pi11 & w878;
assign v423 = ~(pi11 | w878);
assign w880 = v423;
assign v424 = ~(w879 | w880);
assign w881 = v424;
assign w882 = w877 & w881;
assign v425 = ~(w877 | w881);
assign w883 = v425;
assign v426 = ~(w882 | w883);
assign w884 = v426;
assign w885 = ~w873 & w884;
assign w886 = w873 & ~w884;
assign v427 = ~(w885 | w886);
assign w887 = v427;
assign w888 = (~w775 & ~w777) | (~w775 & w16819) | (~w777 & w16819);
assign w889 = ~w887 & w888;
assign w890 = w887 & ~w888;
assign v428 = ~(w889 | w890);
assign w891 = v428;
assign w892 = (~w806 & ~w808) | (~w806 & w17029) | (~w808 & w17029);
assign w893 = ~w891 & w892;
assign w894 = w891 & ~w892;
assign v429 = ~(w893 | w894);
assign w895 = v429;
assign w896 = w872 & w895;
assign v430 = ~(w872 | w895);
assign w897 = v430;
assign v431 = ~(w896 | w897);
assign w898 = v431;
assign w899 = ~w821 & w898;
assign w900 = w821 & ~w898;
assign v432 = ~(w899 | w900);
assign w901 = v432;
assign v433 = ~(w735 | w815);
assign w902 = v433;
assign w903 = (w902 & w661) | (w902 & w16496) | (w661 & w16496);
assign v434 = ~(w816 | w903);
assign w904 = v434;
assign w905 = w901 & w904;
assign v435 = ~(w901 | w904);
assign w906 = v435;
assign v436 = ~(w905 | w906);
assign w907 = v436;
assign v437 = ~(w894 | w896);
assign w908 = v437;
assign w909 = (~w875 & ~w877) | (~w875 & w17030) | (~w877 & w17030);
assign v438 = ~(w837 | w841);
assign w910 = v438;
assign v439 = ~(w840 | w910);
assign w911 = v439;
assign v440 = ~(w846 | w850);
assign w912 = v440;
assign v441 = ~(w849 | w912);
assign w913 = v441;
assign w914 = w911 & w913;
assign v442 = ~(w911 | w913);
assign w915 = v442;
assign v443 = ~(w914 | w915);
assign w916 = v443;
assign w917 = w909 & ~w916;
assign w918 = ~w909 & w916;
assign v444 = ~(w917 | w918);
assign w919 = v444;
assign w920 = (~w885 & ~w887) | (~w885 & w16820) | (~w887 & w16820);
assign w921 = ~w919 & w920;
assign w922 = w919 & ~w920;
assign v445 = ~(w921 | w922);
assign w923 = v445;
assign w924 = pi09 & pi13;
assign w925 = pi06 & pi16;
assign w926 = pi02 & pi20;
assign v446 = ~(w925 | w926);
assign w927 = v446;
assign w928 = w925 & w926;
assign v447 = ~(w927 | w928);
assign w929 = v447;
assign w930 = w924 & ~w929;
assign w931 = ~w924 & w929;
assign v448 = ~(w930 | w931);
assign w932 = v448;
assign w933 = pi00 & pi22;
assign w934 = pi07 & pi15;
assign w935 = pi08 & pi14;
assign v449 = ~(w934 | w935);
assign w936 = v449;
assign w937 = w934 & w935;
assign v450 = ~(w936 | w937);
assign w938 = v450;
assign w939 = w933 & ~w938;
assign w940 = ~w933 & w938;
assign v451 = ~(w939 | w940);
assign w941 = v451;
assign v452 = ~(w932 | w941);
assign w942 = v452;
assign w943 = w932 & w941;
assign v453 = ~(w942 | w943);
assign w944 = v453;
assign w945 = pi03 & pi19;
assign w946 = pi05 & pi17;
assign w947 = pi04 & pi18;
assign v454 = ~(w946 | w947);
assign w948 = v454;
assign w949 = w946 & w947;
assign v455 = ~(w948 | w949);
assign w950 = v455;
assign w951 = w945 & ~w950;
assign w952 = ~w945 & w950;
assign v456 = ~(w951 | w952);
assign w953 = v456;
assign w954 = w944 & ~w953;
assign w955 = ~w944 & w953;
assign v457 = ~(w954 | w955);
assign w956 = v457;
assign v458 = ~(w923 | w956);
assign w957 = v458;
assign w958 = w923 & w956;
assign v459 = ~(w957 | w958);
assign w959 = v459;
assign v460 = ~(w835 | w871);
assign w960 = v460;
assign w961 = (~w855 & ~w857) | (~w855 & w17282) | (~w857 & w17282);
assign w962 = (~w826 & ~w828) | (~w826 & w17031) | (~w828 & w17031);
assign w963 = pi10 & pi12;
assign w964 = pi01 & pi21;
assign v461 = ~(w963 | w964);
assign w965 = v461;
assign w966 = w963 & w964;
assign v462 = ~(w965 | w966);
assign w967 = v462;
assign w968 = w879 & w967;
assign v463 = ~(w879 | w967);
assign w969 = v463;
assign v464 = ~(w968 | w969);
assign w970 = v464;
assign v465 = ~(w858 | w862);
assign w971 = v465;
assign v466 = ~(w861 | w971);
assign w972 = v466;
assign w973 = w970 & w972;
assign v467 = ~(w970 | w972);
assign w974 = v467;
assign v468 = ~(w973 | w974);
assign w975 = v468;
assign w976 = ~w962 & w975;
assign w977 = w962 & ~w975;
assign v469 = ~(w976 | w977);
assign w978 = v469;
assign w979 = ~w961 & w978;
assign w980 = w961 & ~w978;
assign v470 = ~(w979 | w980);
assign w981 = v470;
assign w982 = ~w960 & w981;
assign w983 = w960 & ~w981;
assign v471 = ~(w982 | w983);
assign w984 = v471;
assign w985 = w959 & w984;
assign v472 = ~(w959 | w984);
assign w986 = v472;
assign v473 = ~(w985 | w986);
assign w987 = v473;
assign w988 = ~w908 & w987;
assign w989 = w908 & ~w987;
assign v474 = ~(w988 | w989);
assign w990 = v474;
assign w991 = (w661 & w16821) | (w661 & w16822) | (w16821 & w16822);
assign v475 = ~(w900 | w991);
assign w992 = v475;
assign w993 = w990 & w992;
assign v476 = ~(w990 | w992);
assign w994 = v476;
assign v477 = ~(w993 | w994);
assign w995 = v477;
assign v478 = ~(w982 | w985);
assign w996 = v478;
assign w997 = (~w976 & ~w978) | (~w976 & w17283) | (~w978 & w17283);
assign w998 = (~w968 & ~w970) | (~w968 & w16707) | (~w970 & w16707);
assign w999 = pi04 & pi19;
assign w1000 = pi11 & pi12;
assign w1001 = pi10 & pi13;
assign v479 = ~(w1000 | w1001);
assign w1002 = v479;
assign w1003 = w1000 & w1001;
assign v480 = ~(w1002 | w1003);
assign w1004 = v480;
assign w1005 = w999 & ~w1004;
assign w1006 = ~w999 & w1004;
assign v481 = ~(w1005 | w1006);
assign w1007 = v481;
assign w1008 = pi06 & pi17;
assign w1009 = pi05 & pi18;
assign w1010 = pi03 & pi20;
assign v482 = ~(w1009 | w1010);
assign w1011 = v482;
assign w1012 = w1009 & w1010;
assign v483 = ~(w1011 | w1012);
assign w1013 = v483;
assign w1014 = w1008 & ~w1013;
assign w1015 = ~w1008 & w1013;
assign v484 = ~(w1014 | w1015);
assign w1016 = v484;
assign v485 = ~(w1007 | w1016);
assign w1017 = v485;
assign w1018 = w1007 & w1016;
assign v486 = ~(w1017 | w1018);
assign w1019 = v486;
assign w1020 = w998 & ~w1019;
assign w1021 = ~w998 & w1019;
assign v487 = ~(w1020 | w1021);
assign w1022 = v487;
assign v488 = ~(w933 | w937);
assign w1023 = v488;
assign v489 = ~(w936 | w1023);
assign w1024 = v489;
assign w1025 = pi00 & pi23;
assign w1026 = pi02 & pi21;
assign v490 = ~(w1025 | w1026);
assign w1027 = v490;
assign w1028 = pi02 & pi23;
assign w1029 = w874 & w1028;
assign v491 = ~(w1027 | w1029);
assign w1030 = v491;
assign w1031 = w966 & ~w1030;
assign w1032 = ~w966 & w1030;
assign v492 = ~(w1031 | w1032);
assign w1033 = v492;
assign w1034 = w1024 & ~w1033;
assign w1035 = ~w1024 & w1033;
assign v493 = ~(w1034 | w1035);
assign w1036 = v493;
assign w1037 = pi07 & pi16;
assign w1038 = pi08 & pi15;
assign w1039 = pi09 & pi14;
assign v494 = ~(w1038 | w1039);
assign w1040 = v494;
assign w1041 = w1038 & w1039;
assign v495 = ~(w1040 | w1041);
assign w1042 = v495;
assign w1043 = w1037 & ~w1042;
assign w1044 = ~w1037 & w1042;
assign v496 = ~(w1043 | w1044);
assign w1045 = v496;
assign w1046 = w1036 & ~w1045;
assign w1047 = ~w1036 & w1045;
assign v497 = ~(w1046 | w1047);
assign w1048 = v497;
assign w1049 = w1022 & w1048;
assign v498 = ~(w1022 | w1048);
assign w1050 = v498;
assign v499 = ~(w1049 | w1050);
assign w1051 = v499;
assign w1052 = ~w997 & w1051;
assign w1053 = w997 & ~w1051;
assign v500 = ~(w1052 | w1053);
assign w1054 = v500;
assign w1055 = (~w922 & ~w923) | (~w922 & w17032) | (~w923 & w17032);
assign w1056 = pi01 & pi22;
assign w1057 = pi12 & w1056;
assign v501 = ~(pi12 | w1056);
assign w1058 = v501;
assign v502 = ~(w1057 | w1058);
assign w1059 = v502;
assign v503 = ~(w945 | w949);
assign w1060 = v503;
assign v504 = ~(w948 | w1060);
assign w1061 = v504;
assign w1062 = w1059 & w1061;
assign v505 = ~(w1059 | w1061);
assign w1063 = v505;
assign v506 = ~(w1062 | w1063);
assign w1064 = v506;
assign v507 = ~(w924 | w928);
assign w1065 = v507;
assign v508 = ~(w927 | w1065);
assign w1066 = v508;
assign w1067 = w1064 & w1066;
assign v509 = ~(w1064 | w1066);
assign w1068 = v509;
assign v510 = ~(w1067 | w1068);
assign w1069 = v510;
assign w1070 = (~w914 & ~w916) | (~w914 & w17033) | (~w916 & w17033);
assign w1071 = (~w942 & ~w944) | (~w942 & w16823) | (~w944 & w16823);
assign v511 = ~(w1070 | w1071);
assign w1072 = v511;
assign w1073 = w1070 & w1071;
assign v512 = ~(w1072 | w1073);
assign w1074 = v512;
assign w1075 = w1069 & w1074;
assign v513 = ~(w1069 | w1074);
assign w1076 = v513;
assign v514 = ~(w1075 | w1076);
assign w1077 = v514;
assign w1078 = ~w1055 & w1077;
assign w1079 = w1055 & ~w1077;
assign v515 = ~(w1078 | w1079);
assign w1080 = v515;
assign w1081 = w1054 & w1080;
assign v516 = ~(w1054 | w1080);
assign w1082 = v516;
assign v517 = ~(w1081 | w1082);
assign w1083 = v517;
assign w1084 = w996 & ~w1083;
assign w1085 = ~w996 & w1083;
assign v518 = ~(w1084 | w1085);
assign w1086 = v518;
assign v519 = ~(w900 | w989);
assign w1087 = v519;
assign w1088 = ~w991 & w1087;
assign v520 = ~(w988 | w1088);
assign w1089 = v520;
assign w1090 = w1086 & w1089;
assign v521 = ~(w1086 | w1089);
assign w1091 = v521;
assign v522 = ~(w1090 | w1091);
assign w1092 = v522;
assign v523 = ~(w988 | w1085);
assign w1093 = v523;
assign w1094 = (~w1084 & w1088) | (~w1084 & w16498) | (w1088 & w16498);
assign w1095 = (~w1078 & ~w1080) | (~w1078 & w17284) | (~w1080 & w17284);
assign w1096 = (~w1049 & ~w1051) | (~w1049 & w17285) | (~w1051 & w17285);
assign v524 = ~(w1008 | w1012);
assign w1097 = v524;
assign v525 = ~(w1011 | w1097);
assign w1098 = v525;
assign v526 = ~(w999 | w1003);
assign w1099 = v526;
assign v527 = ~(w1002 | w1099);
assign w1100 = v527;
assign w1101 = w1098 & w1100;
assign v528 = ~(w1098 | w1100);
assign w1102 = v528;
assign v529 = ~(w1101 | w1102);
assign w1103 = v529;
assign v530 = ~(w1037 | w1041);
assign w1104 = v530;
assign v531 = ~(w1040 | w1104);
assign w1105 = v531;
assign v532 = ~(w1103 | w1105);
assign w1106 = v532;
assign w1107 = w1103 & w1105;
assign v533 = ~(w1106 | w1107);
assign w1108 = v533;
assign w1109 = (~w1017 & ~w1019) | (~w1017 & w16708) | (~w1019 & w16708);
assign w1110 = (~w1034 & ~w1036) | (~w1034 & w16709) | (~w1036 & w16709);
assign v534 = ~(w1109 | w1110);
assign w1111 = v534;
assign w1112 = w1109 & w1110;
assign v535 = ~(w1111 | w1112);
assign w1113 = v535;
assign w1114 = w1108 & w1113;
assign v536 = ~(w1108 | w1113);
assign w1115 = v536;
assign v537 = ~(w1114 | w1115);
assign w1116 = v537;
assign w1117 = ~w1096 & w1116;
assign w1118 = w1096 & ~w1116;
assign v538 = ~(w1117 | w1118);
assign w1119 = v538;
assign w1120 = (~w1072 & ~w1074) | (~w1072 & w17034) | (~w1074 & w17034);
assign w1121 = (~w1062 & ~w1064) | (~w1062 & w17035) | (~w1064 & w17035);
assign w1122 = pi00 & pi24;
assign w1123 = w1057 & w1122;
assign v539 = ~(w1057 | w1122);
assign w1124 = v539;
assign v540 = ~(w1123 | w1124);
assign w1125 = v540;
assign w1126 = pi11 & pi13;
assign w1127 = pi01 & pi23;
assign v541 = ~(w1126 | w1127);
assign w1128 = v541;
assign w1129 = pi11 & pi23;
assign w1130 = w366 & w1129;
assign v542 = ~(w1128 | w1130);
assign w1131 = v542;
assign w1132 = w1125 & w1131;
assign v543 = ~(w1125 | w1131);
assign w1133 = v543;
assign v544 = ~(w1132 | w1133);
assign w1134 = v544;
assign w1135 = pi07 & pi17;
assign w1136 = pi02 & pi22;
assign w1137 = pi06 & pi18;
assign v545 = ~(w1136 | w1137);
assign w1138 = v545;
assign w1139 = w1136 & w1137;
assign v546 = ~(w1138 | w1139);
assign w1140 = v546;
assign w1141 = w1135 & ~w1140;
assign w1142 = ~w1135 & w1140;
assign v547 = ~(w1141 | w1142);
assign w1143 = v547;
assign w1144 = w1134 & ~w1143;
assign w1145 = ~w1134 & w1143;
assign v548 = ~(w1144 | w1145);
assign w1146 = v548;
assign w1147 = w1121 & ~w1146;
assign w1148 = ~w1121 & w1146;
assign v549 = ~(w1147 | w1148);
assign w1149 = v549;
assign w1150 = w966 & ~w1027;
assign v550 = ~(w1029 | w1150);
assign w1151 = v550;
assign w1152 = pi03 & pi21;
assign w1153 = pi05 & pi19;
assign w1154 = pi04 & pi20;
assign v551 = ~(w1153 | w1154);
assign w1155 = v551;
assign w1156 = w1153 & w1154;
assign v552 = ~(w1155 | w1156);
assign w1157 = v552;
assign w1158 = w1152 & ~w1157;
assign w1159 = ~w1152 & w1157;
assign v553 = ~(w1158 | w1159);
assign w1160 = v553;
assign v554 = ~(w1151 | w1160);
assign w1161 = v554;
assign w1162 = w1151 & w1160;
assign v555 = ~(w1161 | w1162);
assign w1163 = v555;
assign w1164 = pi08 & pi16;
assign w1165 = pi09 & pi15;
assign w1166 = pi10 & pi14;
assign v556 = ~(w1165 | w1166);
assign w1167 = v556;
assign w1168 = w1165 & w1166;
assign v557 = ~(w1167 | w1168);
assign w1169 = v557;
assign w1170 = w1164 & ~w1169;
assign w1171 = ~w1164 & w1169;
assign v558 = ~(w1170 | w1171);
assign w1172 = v558;
assign w1173 = w1163 & ~w1172;
assign w1174 = ~w1163 & w1172;
assign v559 = ~(w1173 | w1174);
assign w1175 = v559;
assign w1176 = w1149 & w1175;
assign v560 = ~(w1149 | w1175);
assign w1177 = v560;
assign v561 = ~(w1176 | w1177);
assign w1178 = v561;
assign w1179 = ~w1120 & w1178;
assign w1180 = w1120 & ~w1178;
assign v562 = ~(w1179 | w1180);
assign w1181 = v562;
assign w1182 = w1119 & w1181;
assign v563 = ~(w1119 | w1181);
assign w1183 = v563;
assign v564 = ~(w1182 | w1183);
assign w1184 = v564;
assign w1185 = ~w1095 & w1184;
assign w1186 = w1095 & ~w1184;
assign v565 = ~(w1185 | w1186);
assign w1187 = v565;
assign w1188 = w1094 & ~w1187;
assign w1189 = ~w1094 & w1187;
assign v566 = ~(w1188 | w1189);
assign w1190 = v566;
assign v567 = ~(w1117 | w1182);
assign w1191 = v567;
assign w1192 = (~w1123 & ~w1125) | (~w1123 & w16710) | (~w1125 & w16710);
assign v568 = ~(w1164 | w1168);
assign w1193 = v568;
assign v569 = ~(w1167 | w1193);
assign w1194 = v569;
assign v570 = ~(w1135 | w1139);
assign w1195 = v570;
assign v571 = ~(w1138 | w1195);
assign w1196 = v571;
assign w1197 = w1194 & w1196;
assign v572 = ~(w1194 | w1196);
assign w1198 = v572;
assign v573 = ~(w1197 | w1198);
assign w1199 = v573;
assign w1200 = w1192 & ~w1199;
assign w1201 = ~w1192 & w1199;
assign v574 = ~(w1200 | w1201);
assign w1202 = v574;
assign w1203 = (~w1161 & ~w1163) | (~w1161 & w16824) | (~w1163 & w16824);
assign w1204 = ~w1202 & w1203;
assign w1205 = w1202 & ~w1203;
assign v575 = ~(w1204 | w1205);
assign w1206 = v575;
assign w1207 = (~w1144 & ~w1146) | (~w1144 & w17036) | (~w1146 & w17036);
assign w1208 = ~w1206 & w1207;
assign w1209 = w1206 & ~w1207;
assign v576 = ~(w1208 | w1209);
assign w1210 = v576;
assign w1211 = (~w1176 & ~w1178) | (~w1176 & w17037) | (~w1178 & w17037);
assign w1212 = ~w1210 & w1211;
assign w1213 = w1210 & ~w1211;
assign v577 = ~(w1212 | w1213);
assign w1214 = v577;
assign w1215 = pi01 & pi24;
assign w1216 = (w1215 & w1130) | (w1215 & w16825) | (w1130 & w16825);
assign w1217 = ~w1130 & w16826;
assign v578 = ~(w1216 | w1217);
assign w1218 = v578;
assign v579 = ~(w1152 | w1156);
assign w1219 = v579;
assign v580 = ~(w1155 | w1219);
assign w1220 = v580;
assign w1221 = ~w1218 & w1220;
assign w1222 = w1218 & ~w1220;
assign v581 = ~(w1221 | w1222);
assign w1223 = v581;
assign w1224 = (~w1101 & ~w1103) | (~w1101 & w17038) | (~w1103 & w17038);
assign w1225 = pi05 & pi20;
assign w1226 = pi12 & pi13;
assign w1227 = pi11 & pi14;
assign v582 = ~(w1226 | w1227);
assign w1228 = v582;
assign w1229 = w1226 & w1227;
assign v583 = ~(w1228 | w1229);
assign w1230 = v583;
assign w1231 = w1225 & ~w1230;
assign w1232 = ~w1225 & w1230;
assign v584 = ~(w1231 | w1232);
assign w1233 = v584;
assign v585 = ~(w1224 | w1233);
assign w1234 = v585;
assign w1235 = w1224 & w1233;
assign v586 = ~(w1234 | w1235);
assign w1236 = v586;
assign v587 = ~(w1223 | w1236);
assign w1237 = v587;
assign w1238 = w1223 & w1236;
assign v588 = ~(w1237 | w1238);
assign w1239 = v588;
assign w1240 = (~w1111 & ~w1113) | (~w1111 & w16827) | (~w1113 & w16827);
assign w1241 = pi10 & pi15;
assign w1242 = pi00 & pi25;
assign v589 = ~(w1028 | w1242);
assign w1243 = v589;
assign w1244 = pi02 & pi25;
assign w1245 = w1025 & w1244;
assign v590 = ~(w1243 | w1245);
assign w1246 = v590;
assign w1247 = w1241 & ~w1246;
assign w1248 = ~w1241 & w1246;
assign v591 = ~(w1247 | w1248);
assign w1249 = v591;
assign w1250 = pi07 & pi18;
assign w1251 = pi08 & pi17;
assign w1252 = pi09 & pi16;
assign v592 = ~(w1251 | w1252);
assign w1253 = v592;
assign w1254 = w1251 & w1252;
assign v593 = ~(w1253 | w1254);
assign w1255 = v593;
assign w1256 = w1250 & ~w1255;
assign w1257 = ~w1250 & w1255;
assign v594 = ~(w1256 | w1257);
assign w1258 = v594;
assign v595 = ~(w1249 | w1258);
assign w1259 = v595;
assign w1260 = w1249 & w1258;
assign v596 = ~(w1259 | w1260);
assign w1261 = v596;
assign w1262 = pi06 & pi19;
assign w1263 = pi03 & pi22;
assign w1264 = pi04 & pi21;
assign v597 = ~(w1263 | w1264);
assign w1265 = v597;
assign w1266 = w1263 & w1264;
assign v598 = ~(w1265 | w1266);
assign w1267 = v598;
assign w1268 = w1262 & ~w1267;
assign w1269 = ~w1262 & w1267;
assign v599 = ~(w1268 | w1269);
assign w1270 = v599;
assign w1271 = w1261 & ~w1270;
assign w1272 = ~w1261 & w1270;
assign v600 = ~(w1271 | w1272);
assign w1273 = v600;
assign w1274 = ~w1240 & w1273;
assign w1275 = w1240 & ~w1273;
assign v601 = ~(w1274 | w1275);
assign w1276 = v601;
assign w1277 = w1239 & w1276;
assign v602 = ~(w1239 | w1276);
assign w1278 = v602;
assign v603 = ~(w1277 | w1278);
assign w1279 = v603;
assign w1280 = w1214 & w1279;
assign v604 = ~(w1214 | w1279);
assign w1281 = v604;
assign v605 = ~(w1280 | w1281);
assign w1282 = v605;
assign w1283 = w1191 & ~w1282;
assign w1284 = ~w1191 & w1282;
assign v606 = ~(w1283 | w1284);
assign w1285 = v606;
assign v607 = ~(w1094 | w1185);
assign w1286 = v607;
assign v608 = ~(w1186 | w1286);
assign w1287 = v608;
assign w1288 = w1285 & w1287;
assign v609 = ~(w1285 | w1287);
assign w1289 = v609;
assign v610 = ~(w1288 | w1289);
assign w1290 = v610;
assign v611 = ~(w1213 | w1280);
assign w1291 = v611;
assign w1292 = (~w1274 & ~w1276) | (~w1274 & w17039) | (~w1276 & w17039);
assign w1293 = (~w1234 & ~w1236) | (~w1234 & w17286) | (~w1236 & w17286);
assign w1294 = (~w1259 & ~w1261) | (~w1259 & w17287) | (~w1261 & w17287);
assign w1295 = pi12 & pi14;
assign w1296 = pi01 & pi25;
assign v612 = ~(w1295 | w1296);
assign w1297 = v612;
assign w1298 = w1295 & w1296;
assign v613 = ~(w1297 | w1298);
assign w1299 = v613;
assign v614 = ~(w1225 | w1229);
assign w1300 = v614;
assign v615 = ~(w1228 | w1300);
assign w1301 = v615;
assign w1302 = w1299 & w1301;
assign v616 = ~(w1299 | w1301);
assign w1303 = v616;
assign v617 = ~(w1302 | w1303);
assign w1304 = v617;
assign v618 = ~(w1262 | w1266);
assign w1305 = v618;
assign v619 = ~(w1265 | w1305);
assign w1306 = v619;
assign w1307 = w1304 & w1306;
assign v620 = ~(w1304 | w1306);
assign w1308 = v620;
assign v621 = ~(w1307 | w1308);
assign w1309 = v621;
assign w1310 = ~w1294 & w1309;
assign w1311 = w1294 & ~w1309;
assign v622 = ~(w1310 | w1311);
assign w1312 = v622;
assign w1313 = ~w1293 & w1312;
assign w1314 = w1293 & ~w1312;
assign v623 = ~(w1313 | w1314);
assign w1315 = v623;
assign w1316 = ~w1292 & w1315;
assign w1317 = w1292 & ~w1315;
assign v624 = ~(w1316 | w1317);
assign w1318 = v624;
assign v625 = ~(w1250 | w1254);
assign w1319 = v625;
assign v626 = ~(w1253 | w1319);
assign w1320 = v626;
assign w1321 = w1241 & ~w1243;
assign v627 = ~(w1245 | w1321);
assign w1322 = v627;
assign w1323 = w1320 & ~w1322;
assign w1324 = ~w1320 & w1322;
assign v628 = ~(w1323 | w1324);
assign w1325 = v628;
assign w1326 = pi13 & w1215;
assign w1327 = pi00 & pi26;
assign w1328 = pi08 & pi18;
assign v629 = ~(w1327 | w1328);
assign w1329 = v629;
assign w1330 = w1327 & w1328;
assign v630 = ~(w1329 | w1330);
assign w1331 = v630;
assign w1332 = w1326 & ~w1331;
assign w1333 = ~w1326 & w1331;
assign v631 = ~(w1332 | w1333);
assign w1334 = v631;
assign w1335 = ~w1325 & w1334;
assign w1336 = w1325 & ~w1334;
assign v632 = ~(w1335 | w1336);
assign w1337 = v632;
assign w1338 = (~w1197 & ~w1199) | (~w1197 & w16711) | (~w1199 & w16711);
assign w1339 = ~pi24 & w1130;
assign v633 = ~(w1221 | w1339);
assign w1340 = v633;
assign v634 = ~(w1338 | w1340);
assign w1341 = v634;
assign w1342 = w1338 & w1340;
assign v635 = ~(w1341 | w1342);
assign w1343 = v635;
assign w1344 = w1337 & w1343;
assign v636 = ~(w1337 | w1343);
assign w1345 = v636;
assign v637 = ~(w1344 | w1345);
assign w1346 = v637;
assign w1347 = (~w1205 & ~w1206) | (~w1205 & w17040) | (~w1206 & w17040);
assign w1348 = pi02 & pi24;
assign w1349 = pi03 & pi23;
assign w1350 = pi07 & pi19;
assign v638 = ~(w1349 | w1350);
assign w1351 = v638;
assign w1352 = w1349 & w1350;
assign v639 = ~(w1351 | w1352);
assign w1353 = v639;
assign w1354 = w1348 & ~w1353;
assign w1355 = ~w1348 & w1353;
assign v640 = ~(w1354 | w1355);
assign w1356 = v640;
assign w1357 = pi09 & pi17;
assign w1358 = pi10 & pi16;
assign w1359 = pi11 & pi15;
assign v641 = ~(w1358 | w1359);
assign w1360 = v641;
assign w1361 = w1358 & w1359;
assign v642 = ~(w1360 | w1361);
assign w1362 = v642;
assign w1363 = w1357 & ~w1362;
assign w1364 = ~w1357 & w1362;
assign v643 = ~(w1363 | w1364);
assign w1365 = v643;
assign v644 = ~(w1356 | w1365);
assign w1366 = v644;
assign w1367 = w1356 & w1365;
assign v645 = ~(w1366 | w1367);
assign w1368 = v645;
assign w1369 = pi04 & pi22;
assign w1370 = pi06 & pi20;
assign w1371 = pi05 & pi21;
assign v646 = ~(w1370 | w1371);
assign w1372 = v646;
assign w1373 = w1370 & w1371;
assign v647 = ~(w1372 | w1373);
assign w1374 = v647;
assign w1375 = w1369 & ~w1374;
assign w1376 = ~w1369 & w1374;
assign v648 = ~(w1375 | w1376);
assign w1377 = v648;
assign w1378 = w1368 & ~w1377;
assign w1379 = ~w1368 & w1377;
assign v649 = ~(w1378 | w1379);
assign w1380 = v649;
assign w1381 = ~w1347 & w1380;
assign w1382 = w1347 & ~w1380;
assign v650 = ~(w1381 | w1382);
assign w1383 = v650;
assign w1384 = w1346 & w1383;
assign v651 = ~(w1346 | w1383);
assign w1385 = v651;
assign v652 = ~(w1384 | w1385);
assign w1386 = v652;
assign w1387 = w1318 & w1386;
assign v653 = ~(w1318 | w1386);
assign w1388 = v653;
assign v654 = ~(w1387 | w1388);
assign w1389 = v654;
assign w1390 = ~w1291 & w1389;
assign w1391 = w1291 & ~w1389;
assign v655 = ~(w1390 | w1391);
assign w1392 = v655;
assign v656 = ~(w1186 | w1283);
assign w1393 = v656;
assign w1394 = (w1393 & w1094) | (w1393 & w16499) | (w1094 & w16499);
assign v657 = ~(w1284 | w1394);
assign w1395 = v657;
assign w1396 = w1392 & w1395;
assign v658 = ~(w1392 | w1395);
assign w1397 = v658;
assign v659 = ~(w1396 | w1397);
assign w1398 = v659;
assign v660 = ~(w1316 | w1387);
assign w1399 = v660;
assign w1400 = (~w1381 & ~w1383) | (~w1381 & w17288) | (~w1383 & w17288);
assign w1401 = pi26 & w400;
assign w1402 = pi01 & pi26;
assign v661 = ~(pi14 | w1402);
assign w1403 = v661;
assign v662 = ~(w1401 | w1403);
assign w1404 = v662;
assign w1405 = pi00 & pi27;
assign w1406 = w1298 & w1405;
assign v663 = ~(w1298 | w1405);
assign w1407 = v663;
assign v664 = ~(w1406 | w1407);
assign w1408 = v664;
assign w1409 = w1404 & w1408;
assign v665 = ~(w1404 | w1408);
assign w1410 = v665;
assign v666 = ~(w1409 | w1410);
assign w1411 = v666;
assign w1412 = pi03 & pi24;
assign w1413 = pi06 & pi21;
assign w1414 = pi04 & pi23;
assign v667 = ~(w1413 | w1414);
assign w1415 = v667;
assign w1416 = w1413 & w1414;
assign v668 = ~(w1415 | w1416);
assign w1417 = v668;
assign w1418 = w1412 & ~w1417;
assign w1419 = ~w1412 & w1417;
assign v669 = ~(w1418 | w1419);
assign w1420 = v669;
assign w1421 = pi05 & pi22;
assign w1422 = pi12 & pi15;
assign w1423 = pi13 & pi14;
assign v670 = ~(w1422 | w1423);
assign w1424 = v670;
assign w1425 = w1422 & w1423;
assign v671 = ~(w1424 | w1425);
assign w1426 = v671;
assign w1427 = w1421 & ~w1426;
assign w1428 = ~w1421 & w1426;
assign v672 = ~(w1427 | w1428);
assign w1429 = v672;
assign v673 = ~(w1420 | w1429);
assign w1430 = v673;
assign w1431 = w1420 & w1429;
assign v674 = ~(w1430 | w1431);
assign w1432 = v674;
assign w1433 = w1411 & w1432;
assign v675 = ~(w1411 | w1432);
assign w1434 = v675;
assign v676 = ~(w1433 | w1434);
assign w1435 = v676;
assign v677 = ~(w1369 | w1373);
assign w1436 = v677;
assign v678 = ~(w1372 | w1436);
assign w1437 = v678;
assign v679 = ~(w1357 | w1361);
assign w1438 = v679;
assign v680 = ~(w1360 | w1438);
assign w1439 = v680;
assign w1440 = w1437 & w1439;
assign v681 = ~(w1437 | w1439);
assign w1441 = v681;
assign v682 = ~(w1440 | w1441);
assign w1442 = v682;
assign v683 = ~(w1348 | w1352);
assign w1443 = v683;
assign v684 = ~(w1351 | w1443);
assign w1444 = v684;
assign v685 = ~(w1442 | w1444);
assign w1445 = v685;
assign w1446 = w1442 & w1444;
assign v686 = ~(w1445 | w1446);
assign w1447 = v686;
assign w1448 = (~w1341 & ~w1343) | (~w1341 & w16828) | (~w1343 & w16828);
assign w1449 = ~w1447 & w1448;
assign w1450 = w1447 & ~w1448;
assign v687 = ~(w1449 | w1450);
assign w1451 = v687;
assign w1452 = w1435 & w1451;
assign v688 = ~(w1435 | w1451);
assign w1453 = v688;
assign v689 = ~(w1452 | w1453);
assign w1454 = v689;
assign w1455 = ~w1400 & w1454;
assign w1456 = w1400 & ~w1454;
assign v690 = ~(w1455 | w1456);
assign w1457 = v690;
assign w1458 = (~w1366 & ~w1368) | (~w1366 & w16829) | (~w1368 & w16829);
assign w1459 = (~w1302 & ~w1304) | (~w1302 & w16712) | (~w1304 & w16712);
assign w1460 = (~w1323 & ~w1325) | (~w1323 & w16713) | (~w1325 & w16713);
assign v691 = ~(w1459 | w1460);
assign w1461 = v691;
assign w1462 = w1459 & w1460;
assign v692 = ~(w1461 | w1462);
assign w1463 = v692;
assign w1464 = w1458 & ~w1463;
assign w1465 = ~w1458 & w1463;
assign v693 = ~(w1464 | w1465);
assign w1466 = v693;
assign v694 = ~(w1326 | w1330);
assign w1467 = v694;
assign v695 = ~(w1329 | w1467);
assign w1468 = v695;
assign w1469 = pi11 & pi16;
assign w1470 = pi07 & pi20;
assign v696 = ~(w1244 | w1470);
assign w1471 = v696;
assign w1472 = w1244 & w1470;
assign v697 = ~(w1471 | w1472);
assign w1473 = v697;
assign w1474 = w1469 & ~w1473;
assign w1475 = ~w1469 & w1473;
assign v698 = ~(w1474 | w1475);
assign w1476 = v698;
assign w1477 = w1468 & ~w1476;
assign w1478 = ~w1468 & w1476;
assign v699 = ~(w1477 | w1478);
assign w1479 = v699;
assign w1480 = pi08 & pi19;
assign w1481 = pi10 & pi17;
assign w1482 = pi09 & pi18;
assign v700 = ~(w1481 | w1482);
assign w1483 = v700;
assign w1484 = w1481 & w1482;
assign v701 = ~(w1483 | w1484);
assign w1485 = v701;
assign w1486 = w1480 & ~w1485;
assign w1487 = ~w1480 & w1485;
assign v702 = ~(w1486 | w1487);
assign w1488 = v702;
assign w1489 = ~w1479 & w1488;
assign w1490 = w1479 & ~w1488;
assign v703 = ~(w1489 | w1490);
assign w1491 = v703;
assign v704 = ~(w1310 | w1313);
assign w1492 = v704;
assign w1493 = w1491 & ~w1492;
assign w1494 = ~w1491 & w1492;
assign v705 = ~(w1493 | w1494);
assign w1495 = v705;
assign w1496 = w1466 & w1495;
assign v706 = ~(w1466 | w1495);
assign w1497 = v706;
assign v707 = ~(w1496 | w1497);
assign w1498 = v707;
assign w1499 = w1457 & w1498;
assign v708 = ~(w1457 | w1498);
assign w1500 = v708;
assign v709 = ~(w1499 | w1500);
assign w1501 = v709;
assign w1502 = ~w1399 & w1501;
assign w1503 = w1399 & ~w1501;
assign v710 = ~(w1502 | w1503);
assign w1504 = v710;
assign v711 = ~(w1284 | w1390);
assign w1505 = v711;
assign w1506 = (~w1094 & w16500) | (~w1094 & w16501) | (w16500 & w16501);
assign v712 = ~(w1391 | w1506);
assign w1507 = v712;
assign w1508 = w1504 & w1507;
assign v713 = ~(w1504 | w1507);
assign w1509 = v713;
assign v714 = ~(w1508 | w1509);
assign w1510 = v714;
assign w1511 = (~w1406 & ~w1408) | (~w1406 & w16714) | (~w1408 & w16714);
assign w1512 = pi08 & pi20;
assign w1513 = pi03 & pi25;
assign w1514 = pi04 & pi24;
assign v715 = ~(w1513 | w1514);
assign w1515 = v715;
assign w1516 = w1513 & w1514;
assign v716 = ~(w1515 | w1516);
assign w1517 = v716;
assign w1518 = w1512 & ~w1517;
assign w1519 = ~w1512 & w1517;
assign v717 = ~(w1518 | w1519);
assign w1520 = v717;
assign v718 = ~(w1511 | w1520);
assign w1521 = v718;
assign w1522 = w1511 & w1520;
assign v719 = ~(w1521 | w1522);
assign w1523 = v719;
assign w1524 = pi07 & pi21;
assign w1525 = pi06 & pi22;
assign w1526 = pi05 & pi23;
assign v720 = ~(w1525 | w1526);
assign w1527 = v720;
assign w1528 = w1525 & w1526;
assign v721 = ~(w1527 | w1528);
assign w1529 = v721;
assign w1530 = w1524 & ~w1529;
assign w1531 = ~w1524 & w1529;
assign v722 = ~(w1530 | w1531);
assign w1532 = v722;
assign w1533 = w1523 & ~w1532;
assign w1534 = ~w1523 & w1532;
assign v723 = ~(w1533 | w1534);
assign w1535 = v723;
assign w1536 = (w1451 & w17289) | (w1451 & w17290) | (w17289 & w17290);
assign w1537 = (~w1451 & w17291) | (~w1451 & w17292) | (w17291 & w17292);
assign v724 = ~(w1536 | w1537);
assign w1538 = v724;
assign v725 = ~(w1430 | w1433);
assign w1539 = v725;
assign w1540 = (~w1477 & ~w1479) | (~w1477 & w17293) | (~w1479 & w17293);
assign w1541 = pi13 & pi15;
assign w1542 = pi01 & pi27;
assign v726 = ~(w1541 | w1542);
assign w1543 = v726;
assign w1544 = w1541 & w1542;
assign v727 = ~(w1543 | w1544);
assign w1545 = v727;
assign w1546 = w1401 & w1545;
assign v728 = ~(w1401 | w1545);
assign w1547 = v728;
assign v729 = ~(w1546 | w1547);
assign w1548 = v729;
assign v730 = ~(w1421 | w1425);
assign w1549 = v730;
assign v731 = ~(w1424 | w1549);
assign w1550 = v731;
assign w1551 = w1548 & w1550;
assign v732 = ~(w1548 | w1550);
assign w1552 = v732;
assign v733 = ~(w1551 | w1552);
assign w1553 = v733;
assign w1554 = ~w1540 & w1553;
assign w1555 = w1540 & ~w1553;
assign v734 = ~(w1554 | w1555);
assign w1556 = v734;
assign w1557 = ~w1539 & w1556;
assign w1558 = w1539 & ~w1556;
assign v735 = ~(w1557 | w1558);
assign w1559 = v735;
assign w1560 = w1538 & w1559;
assign v736 = ~(w1538 | w1559);
assign w1561 = v736;
assign v737 = ~(w1560 | w1561);
assign w1562 = v737;
assign v738 = ~(w1455 | w1499);
assign w1563 = v738;
assign v739 = ~(w1493 | w1496);
assign w1564 = v739;
assign v740 = ~(w1480 | w1484);
assign w1565 = v740;
assign v741 = ~(w1483 | w1565);
assign w1566 = v741;
assign v742 = ~(w1412 | w1416);
assign w1567 = v742;
assign v743 = ~(w1415 | w1567);
assign w1568 = v743;
assign w1569 = w1566 & w1568;
assign v744 = ~(w1566 | w1568);
assign w1570 = v744;
assign v745 = ~(w1569 | w1570);
assign w1571 = v745;
assign v746 = ~(w1469 | w1472);
assign w1572 = v746;
assign v747 = ~(w1471 | w1572);
assign w1573 = v747;
assign v748 = ~(w1571 | w1573);
assign w1574 = v748;
assign w1575 = w1571 & w1573;
assign v749 = ~(w1574 | w1575);
assign w1576 = v749;
assign w1577 = (~w1461 & ~w1463) | (~w1461 & w16830) | (~w1463 & w16830);
assign w1578 = ~w1576 & w1577;
assign w1579 = w1576 & ~w1577;
assign v750 = ~(w1578 | w1579);
assign w1580 = v750;
assign w1581 = (~w1440 & ~w1442) | (~w1440 & w16715) | (~w1442 & w16715);
assign w1582 = pi11 & pi17;
assign w1583 = pi00 & pi28;
assign w1584 = pi12 & pi16;
assign v751 = ~(w1583 | w1584);
assign w1585 = v751;
assign w1586 = w1583 & w1584;
assign v752 = ~(w1585 | w1586);
assign w1587 = v752;
assign w1588 = w1582 & ~w1587;
assign w1589 = ~w1582 & w1587;
assign v753 = ~(w1588 | w1589);
assign w1590 = v753;
assign w1591 = pi02 & pi26;
assign w1592 = pi09 & pi19;
assign w1593 = pi10 & pi18;
assign v754 = ~(w1592 | w1593);
assign w1594 = v754;
assign w1595 = w1592 & w1593;
assign v755 = ~(w1594 | w1595);
assign w1596 = v755;
assign w1597 = w1591 & ~w1596;
assign w1598 = ~w1591 & w1596;
assign v756 = ~(w1597 | w1598);
assign w1599 = v756;
assign v757 = ~(w1590 | w1599);
assign w1600 = v757;
assign w1601 = w1590 & w1599;
assign v758 = ~(w1600 | w1601);
assign w1602 = v758;
assign w1603 = w1581 & ~w1602;
assign w1604 = ~w1581 & w1602;
assign v759 = ~(w1603 | w1604);
assign w1605 = v759;
assign w1606 = w1580 & w1605;
assign v760 = ~(w1580 | w1605);
assign w1607 = v760;
assign v761 = ~(w1606 | w1607);
assign w1608 = v761;
assign w1609 = ~w1564 & w1608;
assign w1610 = w1564 & ~w1608;
assign v762 = ~(w1609 | w1610);
assign w1611 = v762;
assign w1612 = ~w1563 & w1611;
assign w1613 = w1563 & ~w1611;
assign v763 = ~(w1612 | w1613);
assign w1614 = v763;
assign v764 = ~(w1562 | w1614);
assign w1615 = v764;
assign w1616 = w1562 & w1614;
assign v765 = ~(w1615 | w1616);
assign w1617 = v765;
assign w1618 = (~w1094 & w17042) | (~w1094 & w17043) | (w17042 & w17043);
assign v766 = ~(w1503 | w1618);
assign w1619 = v766;
assign w1620 = w1617 & w1619;
assign v767 = ~(w1617 | w1619);
assign w1621 = v767;
assign v768 = ~(w1620 | w1621);
assign w1622 = v768;
assign v769 = ~(w1609 | w1612);
assign w1623 = v769;
assign v770 = ~(w1591 | w1595);
assign w1624 = v770;
assign v771 = ~(w1594 | w1624);
assign w1625 = v771;
assign v772 = ~(w1582 | w1586);
assign w1626 = v772;
assign v773 = ~(w1585 | w1626);
assign w1627 = v773;
assign w1628 = w1625 & w1627;
assign v774 = ~(w1625 | w1627);
assign w1629 = v774;
assign v775 = ~(w1628 | w1629);
assign w1630 = v775;
assign w1631 = pi00 & pi29;
assign w1632 = pi02 & pi27;
assign v776 = ~(w1631 | w1632);
assign w1633 = v776;
assign w1634 = pi02 & pi29;
assign w1635 = w1405 & w1634;
assign v777 = ~(w1633 | w1635);
assign w1636 = v777;
assign w1637 = w1544 & ~w1636;
assign w1638 = ~w1544 & w1636;
assign v778 = ~(w1637 | w1638);
assign w1639 = v778;
assign w1640 = ~w1630 & w1639;
assign w1641 = w1630 & ~w1639;
assign v779 = ~(w1640 | w1641);
assign w1642 = v779;
assign v780 = ~(w1600 | w1604);
assign w1643 = v780;
assign w1644 = (~w1521 & ~w1523) | (~w1521 & w16831) | (~w1523 & w16831);
assign v781 = ~(w1643 | w1644);
assign w1645 = v781;
assign w1646 = w1643 & w1644;
assign v782 = ~(w1645 | w1646);
assign w1647 = v782;
assign w1648 = w1642 & w1647;
assign v783 = ~(w1642 | w1647);
assign w1649 = v783;
assign v784 = ~(w1648 | w1649);
assign w1650 = v784;
assign w1651 = (~w1579 & ~w1580) | (~w1579 & w17044) | (~w1580 & w17044);
assign v785 = ~(w1554 | w1557);
assign w1652 = v785;
assign v786 = ~(w1651 | w1652);
assign w1653 = v786;
assign w1654 = w1651 & w1652;
assign v787 = ~(w1653 | w1654);
assign w1655 = v787;
assign w1656 = w1650 & w1655;
assign v788 = ~(w1650 | w1655);
assign w1657 = v788;
assign v789 = ~(w1656 | w1657);
assign w1658 = v789;
assign v790 = ~(w1536 | w1560);
assign w1659 = v790;
assign w1660 = (~w1569 & ~w1571) | (~w1569 & w17045) | (~w1571 & w17045);
assign w1661 = (~w1546 & ~w1548) | (~w1546 & w16832) | (~w1548 & w16832);
assign w1662 = pi06 & pi23;
assign w1663 = pi14 & pi15;
assign w1664 = pi13 & pi16;
assign v791 = ~(w1663 | w1664);
assign w1665 = v791;
assign w1666 = w1663 & w1664;
assign v792 = ~(w1665 | w1666);
assign w1667 = v792;
assign w1668 = w1662 & ~w1667;
assign w1669 = ~w1662 & w1667;
assign v793 = ~(w1668 | w1669);
assign w1670 = v793;
assign v794 = ~(w1661 | w1670);
assign w1671 = v794;
assign w1672 = w1661 & w1670;
assign v795 = ~(w1671 | w1672);
assign w1673 = v795;
assign w1674 = w1660 & ~w1673;
assign w1675 = ~w1660 & w1673;
assign v796 = ~(w1674 | w1675);
assign w1676 = v796;
assign w1677 = pi28 & w479;
assign w1678 = pi01 & pi28;
assign v797 = ~(pi15 | w1678);
assign w1679 = v797;
assign v798 = ~(w1677 | w1679);
assign w1680 = v798;
assign v799 = ~(w1524 | w1528);
assign w1681 = v799;
assign v800 = ~(w1527 | w1681);
assign w1682 = v800;
assign w1683 = w1680 & w1682;
assign v801 = ~(w1680 | w1682);
assign w1684 = v801;
assign v802 = ~(w1683 | w1684);
assign w1685 = v802;
assign v803 = ~(w1512 | w1516);
assign w1686 = v803;
assign v804 = ~(w1515 | w1686);
assign w1687 = v804;
assign w1688 = w1685 & w1687;
assign v805 = ~(w1685 | w1687);
assign w1689 = v805;
assign v806 = ~(w1688 | w1689);
assign w1690 = v806;
assign w1691 = pi12 & pi17;
assign w1692 = pi03 & pi26;
assign w1693 = pi08 & pi21;
assign v807 = ~(w1692 | w1693);
assign w1694 = v807;
assign w1695 = w1692 & w1693;
assign v808 = ~(w1694 | w1695);
assign w1696 = v808;
assign w1697 = w1691 & ~w1696;
assign w1698 = ~w1691 & w1696;
assign v809 = ~(w1697 | w1698);
assign w1699 = v809;
assign w1700 = pi09 & pi20;
assign w1701 = pi10 & pi19;
assign w1702 = pi11 & pi18;
assign v810 = ~(w1701 | w1702);
assign w1703 = v810;
assign w1704 = w1701 & w1702;
assign v811 = ~(w1703 | w1704);
assign w1705 = v811;
assign w1706 = w1700 & ~w1705;
assign w1707 = ~w1700 & w1705;
assign v812 = ~(w1706 | w1707);
assign w1708 = v812;
assign v813 = ~(w1699 | w1708);
assign w1709 = v813;
assign w1710 = w1699 & w1708;
assign v814 = ~(w1709 | w1710);
assign w1711 = v814;
assign w1712 = pi04 & pi25;
assign w1713 = pi07 & pi22;
assign w1714 = pi05 & pi24;
assign v815 = ~(w1713 | w1714);
assign w1715 = v815;
assign w1716 = w1713 & w1714;
assign v816 = ~(w1715 | w1716);
assign w1717 = v816;
assign w1718 = w1712 & ~w1717;
assign w1719 = ~w1712 & w1717;
assign v817 = ~(w1718 | w1719);
assign w1720 = v817;
assign w1721 = w1711 & ~w1720;
assign w1722 = ~w1711 & w1720;
assign v818 = ~(w1721 | w1722);
assign w1723 = v818;
assign w1724 = w1690 & w1723;
assign v819 = ~(w1690 | w1723);
assign w1725 = v819;
assign v820 = ~(w1724 | w1725);
assign w1726 = v820;
assign w1727 = w1676 & w1726;
assign v821 = ~(w1676 | w1726);
assign w1728 = v821;
assign v822 = ~(w1727 | w1728);
assign w1729 = v822;
assign w1730 = ~w1659 & w1729;
assign w1731 = w1659 & ~w1729;
assign v823 = ~(w1730 | w1731);
assign w1732 = v823;
assign w1733 = w1658 & w1732;
assign v824 = ~(w1658 | w1732);
assign w1734 = v824;
assign v825 = ~(w1733 | w1734);
assign w1735 = v825;
assign w1736 = ~w1623 & w1735;
assign w1737 = w1623 & ~w1735;
assign v826 = ~(w1736 | w1737);
assign w1738 = v826;
assign v827 = ~(w1503 | w1615);
assign w1739 = v827;
assign w1740 = ~w1618 & w1739;
assign v828 = ~(w1616 | w1740);
assign w1741 = v828;
assign w1742 = w1738 & w1741;
assign v829 = ~(w1738 | w1741);
assign w1743 = v829;
assign v830 = ~(w1742 | w1743);
assign w1744 = v830;
assign v831 = ~(w1730 | w1733);
assign w1745 = v831;
assign w1746 = (~w1628 & ~w1630) | (~w1628 & w17046) | (~w1630 & w17046);
assign w1747 = (~w1683 & ~w1685) | (~w1683 & w16716) | (~w1685 & w16716);
assign w1748 = pi00 & pi30;
assign w1749 = w1677 & w1748;
assign v832 = ~(w1677 | w1748);
assign w1750 = v832;
assign v833 = ~(w1749 | w1750);
assign w1751 = v833;
assign w1752 = pi14 & pi16;
assign w1753 = pi01 & pi29;
assign v834 = ~(w1752 | w1753);
assign w1754 = v834;
assign w1755 = pi14 & pi29;
assign w1756 = w519 & w1755;
assign v835 = ~(w1754 | w1756);
assign w1757 = v835;
assign w1758 = w1751 & w1757;
assign v836 = ~(w1751 | w1757);
assign w1759 = v836;
assign v837 = ~(w1758 | w1759);
assign w1760 = v837;
assign w1761 = ~w1747 & w1760;
assign w1762 = w1747 & ~w1760;
assign v838 = ~(w1761 | w1762);
assign w1763 = v838;
assign w1764 = w1746 & ~w1763;
assign w1765 = ~w1746 & w1763;
assign v839 = ~(w1764 | w1765);
assign w1766 = v839;
assign w1767 = (~w1724 & ~w1726) | (~w1724 & w17294) | (~w1726 & w17294);
assign w1768 = ~w1766 & w1767;
assign w1769 = w1766 & ~w1767;
assign v840 = ~(w1768 | w1769);
assign w1770 = v840;
assign v841 = ~(w1691 | w1695);
assign w1771 = v841;
assign v842 = ~(w1694 | w1771);
assign w1772 = v842;
assign v843 = ~(w1700 | w1704);
assign w1773 = v843;
assign v844 = ~(w1703 | w1773);
assign w1774 = v844;
assign w1775 = w1772 & w1774;
assign v845 = ~(w1772 | w1774);
assign w1776 = v845;
assign v846 = ~(w1775 | w1776);
assign w1777 = v846;
assign w1778 = w1544 & ~w1633;
assign v847 = ~(w1635 | w1778);
assign w1779 = v847;
assign w1780 = ~w1777 & w1779;
assign w1781 = w1777 & ~w1779;
assign v848 = ~(w1780 | w1781);
assign w1782 = v848;
assign v849 = ~(w1712 | w1716);
assign w1783 = v849;
assign v850 = ~(w1715 | w1783);
assign w1784 = v850;
assign v851 = ~(w1662 | w1666);
assign w1785 = v851;
assign v852 = ~(w1665 | w1785);
assign w1786 = v852;
assign w1787 = w1784 & w1786;
assign v853 = ~(w1784 | w1786);
assign w1788 = v853;
assign v854 = ~(w1787 | w1788);
assign w1789 = v854;
assign w1790 = pi13 & pi17;
assign w1791 = pi02 & pi28;
assign w1792 = pi09 & pi21;
assign v855 = ~(w1791 | w1792);
assign w1793 = v855;
assign w1794 = w1791 & w1792;
assign v856 = ~(w1793 | w1794);
assign w1795 = v856;
assign w1796 = w1790 & ~w1795;
assign w1797 = ~w1790 & w1795;
assign v857 = ~(w1796 | w1797);
assign w1798 = v857;
assign w1799 = ~w1789 & w1798;
assign w1800 = w1789 & ~w1798;
assign v858 = ~(w1799 | w1800);
assign w1801 = v858;
assign w1802 = (~w1709 & ~w1711) | (~w1709 & w16833) | (~w1711 & w16833);
assign w1803 = w1801 & ~w1802;
assign w1804 = ~w1801 & w1802;
assign v859 = ~(w1803 | w1804);
assign w1805 = v859;
assign w1806 = w1782 & w1805;
assign v860 = ~(w1782 | w1805);
assign w1807 = v860;
assign v861 = ~(w1806 | w1807);
assign w1808 = v861;
assign w1809 = w1770 & w1808;
assign v862 = ~(w1770 | w1808);
assign w1810 = v862;
assign v863 = ~(w1809 | w1810);
assign w1811 = v863;
assign w1812 = (~w1653 & ~w1655) | (~w1653 & w17295) | (~w1655 & w17295);
assign w1813 = (~w1645 & ~w1647) | (~w1645 & w16834) | (~w1647 & w16834);
assign w1814 = (~w1671 & ~w1673) | (~w1671 & w17047) | (~w1673 & w17047);
assign w1815 = pi03 & pi27;
assign w1816 = pi04 & pi26;
assign w1817 = pi08 & pi22;
assign v864 = ~(w1816 | w1817);
assign w1818 = v864;
assign w1819 = w1816 & w1817;
assign v865 = ~(w1818 | w1819);
assign w1820 = v865;
assign w1821 = w1815 & ~w1820;
assign w1822 = ~w1815 & w1820;
assign v866 = ~(w1821 | w1822);
assign w1823 = v866;
assign w1824 = pi05 & pi25;
assign w1825 = pi07 & pi23;
assign w1826 = pi06 & pi24;
assign v867 = ~(w1825 | w1826);
assign w1827 = v867;
assign w1828 = w1825 & w1826;
assign v868 = ~(w1827 | w1828);
assign w1829 = v868;
assign w1830 = w1824 & ~w1829;
assign w1831 = ~w1824 & w1829;
assign v869 = ~(w1830 | w1831);
assign w1832 = v869;
assign v870 = ~(w1823 | w1832);
assign w1833 = v870;
assign w1834 = w1823 & w1832;
assign v871 = ~(w1833 | w1834);
assign w1835 = v871;
assign w1836 = pi10 & pi20;
assign w1837 = pi11 & pi19;
assign w1838 = pi12 & pi18;
assign v872 = ~(w1837 | w1838);
assign w1839 = v872;
assign w1840 = w1837 & w1838;
assign v873 = ~(w1839 | w1840);
assign w1841 = v873;
assign w1842 = w1836 & ~w1841;
assign w1843 = ~w1836 & w1841;
assign v874 = ~(w1842 | w1843);
assign w1844 = v874;
assign w1845 = w1835 & ~w1844;
assign w1846 = ~w1835 & w1844;
assign v875 = ~(w1845 | w1846);
assign w1847 = v875;
assign w1848 = ~w1814 & w1847;
assign w1849 = w1814 & ~w1847;
assign v876 = ~(w1848 | w1849);
assign w1850 = v876;
assign w1851 = ~w1813 & w1850;
assign w1852 = w1813 & ~w1850;
assign v877 = ~(w1851 | w1852);
assign w1853 = v877;
assign w1854 = ~w1812 & w1853;
assign w1855 = w1812 & ~w1853;
assign v878 = ~(w1854 | w1855);
assign w1856 = v878;
assign w1857 = w1811 & w1856;
assign v879 = ~(w1811 | w1856);
assign w1858 = v879;
assign v880 = ~(w1857 | w1858);
assign w1859 = v880;
assign w1860 = ~w1745 & w1859;
assign w1861 = w1745 & ~w1859;
assign v881 = ~(w1860 | w1861);
assign w1862 = v881;
assign v882 = ~(w1616 | w1736);
assign w1863 = v882;
assign w1864 = (~w1737 & w1740) | (~w1737 & w16503) | (w1740 & w16503);
assign w1865 = w1862 & w1864;
assign v883 = ~(w1862 | w1864);
assign w1866 = v883;
assign v884 = ~(w1865 | w1866);
assign w1867 = v884;
assign v885 = ~(w1854 | w1857);
assign w1868 = v885;
assign v886 = ~(w1769 | w1809);
assign w1869 = v886;
assign w1870 = (~w1803 & ~w1805) | (~w1803 & w17048) | (~w1805 & w17048);
assign w1871 = (~w1749 & ~w1751) | (~w1749 & w16835) | (~w1751 & w16835);
assign w1872 = pi11 & pi20;
assign w1873 = pi12 & pi19;
assign w1874 = pi13 & pi18;
assign v887 = ~(w1873 | w1874);
assign w1875 = v887;
assign w1876 = w1873 & w1874;
assign v888 = ~(w1875 | w1876);
assign w1877 = v888;
assign w1878 = w1872 & ~w1877;
assign w1879 = ~w1872 & w1877;
assign v889 = ~(w1878 | w1879);
assign w1880 = v889;
assign v890 = ~(w1871 | w1880);
assign w1881 = v890;
assign w1882 = w1871 & w1880;
assign v891 = ~(w1881 | w1882);
assign w1883 = v891;
assign w1884 = pi10 & pi21;
assign w1885 = pi00 & pi31;
assign w1886 = pi09 & pi22;
assign v892 = ~(w1885 | w1886);
assign w1887 = v892;
assign w1888 = w1885 & w1886;
assign v893 = ~(w1887 | w1888);
assign w1889 = v893;
assign w1890 = w1884 & ~w1889;
assign w1891 = ~w1884 & w1889;
assign v894 = ~(w1890 | w1891);
assign w1892 = v894;
assign w1893 = w1883 & ~w1892;
assign w1894 = ~w1883 & w1892;
assign v895 = ~(w1893 | w1894);
assign w1895 = v895;
assign w1896 = pi06 & pi25;
assign w1897 = pi15 & pi16;
assign w1898 = pi14 & pi17;
assign v896 = ~(w1897 | w1898);
assign w1899 = v896;
assign w1900 = w1897 & w1898;
assign v897 = ~(w1899 | w1900);
assign w1901 = v897;
assign w1902 = w1896 & ~w1901;
assign w1903 = ~w1896 & w1901;
assign v898 = ~(w1902 | w1903);
assign w1904 = v898;
assign w1905 = pi08 & pi23;
assign w1906 = pi07 & pi24;
assign w1907 = pi05 & pi26;
assign v899 = ~(w1906 | w1907);
assign w1908 = v899;
assign w1909 = w1906 & w1907;
assign v900 = ~(w1908 | w1909);
assign w1910 = v900;
assign w1911 = w1905 & ~w1910;
assign w1912 = ~w1905 & w1910;
assign v901 = ~(w1911 | w1912);
assign w1913 = v901;
assign v902 = ~(w1904 | w1913);
assign w1914 = v902;
assign w1915 = w1904 & w1913;
assign v903 = ~(w1914 | w1915);
assign w1916 = v903;
assign w1917 = pi04 & pi27;
assign w1918 = pi03 & pi28;
assign v904 = ~(w1917 | w1918);
assign w1919 = v904;
assign w1920 = w1917 & w1918;
assign v905 = ~(w1919 | w1920);
assign w1921 = v905;
assign w1922 = w1634 & ~w1921;
assign w1923 = ~w1634 & w1921;
assign v906 = ~(w1922 | w1923);
assign w1924 = v906;
assign w1925 = w1916 & ~w1924;
assign w1926 = ~w1916 & w1924;
assign v907 = ~(w1925 | w1926);
assign w1927 = v907;
assign w1928 = w1895 & w1927;
assign v908 = ~(w1895 | w1927);
assign w1929 = v908;
assign v909 = ~(w1928 | w1929);
assign w1930 = v909;
assign w1931 = ~w1870 & w1930;
assign w1932 = w1870 & ~w1930;
assign v910 = ~(w1931 | w1932);
assign w1933 = v910;
assign w1934 = ~w1869 & w1933;
assign w1935 = w1869 & ~w1933;
assign v911 = ~(w1934 | w1935);
assign w1936 = v911;
assign w1937 = (~w1848 & w1813) | (~w1848 & w17049) | (w1813 & w17049);
assign w1938 = pi16 & ~w1756;
assign w1939 = pi01 & pi30;
assign w1940 = ~w1938 & w1939;
assign w1941 = w1938 & ~w1939;
assign v912 = ~(w1940 | w1941);
assign w1942 = v912;
assign v913 = ~(w1824 | w1828);
assign w1943 = v913;
assign v914 = ~(w1827 | w1943);
assign w1944 = v914;
assign w1945 = ~w1942 & w1944;
assign w1946 = w1942 & ~w1944;
assign v915 = ~(w1945 | w1946);
assign w1947 = v915;
assign v916 = ~(w1787 | w1800);
assign w1948 = v916;
assign v917 = ~(w1775 | w1781);
assign w1949 = v917;
assign v918 = ~(w1948 | w1949);
assign w1950 = v918;
assign w1951 = w1948 & w1949;
assign v919 = ~(w1950 | w1951);
assign w1952 = v919;
assign w1953 = w1947 & w1952;
assign v920 = ~(w1947 | w1952);
assign w1954 = v920;
assign v921 = ~(w1953 | w1954);
assign w1955 = v921;
assign w1956 = ~w1937 & w1955;
assign w1957 = w1937 & ~w1955;
assign v922 = ~(w1956 | w1957);
assign w1958 = v922;
assign v923 = ~(w1815 | w1819);
assign w1959 = v923;
assign v924 = ~(w1818 | w1959);
assign w1960 = v924;
assign v925 = ~(w1790 | w1794);
assign w1961 = v925;
assign v926 = ~(w1793 | w1961);
assign w1962 = v926;
assign w1963 = w1960 & w1962;
assign v927 = ~(w1960 | w1962);
assign w1964 = v927;
assign v928 = ~(w1963 | w1964);
assign w1965 = v928;
assign v929 = ~(w1836 | w1840);
assign w1966 = v929;
assign v930 = ~(w1839 | w1966);
assign w1967 = v930;
assign v931 = ~(w1965 | w1967);
assign w1968 = v931;
assign w1969 = w1965 & w1967;
assign v932 = ~(w1968 | w1969);
assign w1970 = v932;
assign w1971 = (~w1833 & ~w1835) | (~w1833 & w16836) | (~w1835 & w16836);
assign w1972 = ~w1970 & w1971;
assign w1973 = w1970 & ~w1971;
assign v933 = ~(w1972 | w1973);
assign w1974 = v933;
assign w1975 = (~w1761 & ~w1763) | (~w1761 & w16837) | (~w1763 & w16837);
assign w1976 = ~w1974 & w1975;
assign w1977 = w1974 & ~w1975;
assign v934 = ~(w1976 | w1977);
assign w1978 = v934;
assign w1979 = w1958 & w1978;
assign v935 = ~(w1958 | w1978);
assign w1980 = v935;
assign v936 = ~(w1979 | w1980);
assign w1981 = v936;
assign w1982 = w1936 & w1981;
assign v937 = ~(w1936 | w1981);
assign w1983 = v937;
assign v938 = ~(w1982 | w1983);
assign w1984 = v938;
assign w1985 = ~w1868 & w1984;
assign w1986 = w1868 & ~w1984;
assign v939 = ~(w1985 | w1986);
assign w1987 = v939;
assign v940 = ~(w1860 | w1864);
assign w1988 = v940;
assign v941 = ~(w1861 | w1988);
assign w1989 = v941;
assign w1990 = w1987 & w1989;
assign v942 = ~(w1987 | w1989);
assign w1991 = v942;
assign v943 = ~(w1990 | w1991);
assign w1992 = v943;
assign v944 = ~(w1861 | w1986);
assign w1993 = v944;
assign w1994 = (w1993 & w1864) | (w1993 & w16504) | (w1864 & w16504);
assign v945 = ~(w1985 | w1994);
assign w1995 = v945;
assign v946 = ~(w1934 | w1982);
assign w1996 = v946;
assign v947 = ~(w1956 | w1979);
assign w1997 = v947;
assign v948 = ~(w1973 | w1977);
assign w1998 = v948;
assign w1999 = ~pi30 & w1756;
assign v949 = ~(w1945 | w1999);
assign w2000 = v949;
assign w2001 = pi09 & pi23;
assign w2002 = pi04 & pi28;
assign w2003 = pi05 & pi27;
assign v950 = ~(w2002 | w2003);
assign w2004 = v950;
assign w2005 = w2002 & w2003;
assign v951 = ~(w2004 | w2005);
assign w2006 = v951;
assign w2007 = w2001 & ~w2006;
assign w2008 = ~w2001 & w2006;
assign v952 = ~(w2007 | w2008);
assign w2009 = v952;
assign w2010 = pi08 & pi24;
assign w2011 = pi07 & pi25;
assign w2012 = pi06 & pi26;
assign v953 = ~(w2011 | w2012);
assign w2013 = v953;
assign w2014 = w2011 & w2012;
assign v954 = ~(w2013 | w2014);
assign w2015 = v954;
assign w2016 = w2010 & ~w2015;
assign w2017 = ~w2010 & w2015;
assign v955 = ~(w2016 | w2017);
assign w2018 = v955;
assign v956 = ~(w2009 | w2018);
assign w2019 = v956;
assign w2020 = w2009 & w2018;
assign v957 = ~(w2019 | w2020);
assign w2021 = v957;
assign w2022 = w2000 & ~w2021;
assign w2023 = ~w2000 & w2021;
assign v958 = ~(w2022 | w2023);
assign w2024 = v958;
assign w2025 = pi16 & w1939;
assign w2026 = pi00 & pi32;
assign w2027 = pi02 & pi30;
assign v959 = ~(w2026 | w2027);
assign w2028 = v959;
assign w2029 = pi02 & pi32;
assign w2030 = w1748 & w2029;
assign v960 = ~(w2028 | w2030);
assign w2031 = v960;
assign w2032 = w2025 & ~w2031;
assign w2033 = ~w2025 & w2031;
assign v961 = ~(w2032 | w2033);
assign w2034 = v961;
assign w2035 = pi11 & pi21;
assign w2036 = pi13 & pi19;
assign w2037 = pi12 & pi20;
assign v962 = ~(w2036 | w2037);
assign w2038 = v962;
assign w2039 = w2036 & w2037;
assign v963 = ~(w2038 | w2039);
assign w2040 = v963;
assign w2041 = w2035 & ~w2040;
assign w2042 = ~w2035 & w2040;
assign v964 = ~(w2041 | w2042);
assign w2043 = v964;
assign v965 = ~(w2034 | w2043);
assign w2044 = v965;
assign w2045 = w2034 & w2043;
assign v966 = ~(w2044 | w2045);
assign w2046 = v966;
assign w2047 = pi14 & pi18;
assign w2048 = pi03 & pi29;
assign w2049 = pi10 & pi22;
assign v967 = ~(w2048 | w2049);
assign w2050 = v967;
assign w2051 = w2048 & w2049;
assign v968 = ~(w2050 | w2051);
assign w2052 = v968;
assign w2053 = w2047 & ~w2052;
assign w2054 = ~w2047 & w2052;
assign v969 = ~(w2053 | w2054);
assign w2055 = v969;
assign w2056 = w2046 & ~w2055;
assign w2057 = ~w2046 & w2055;
assign v970 = ~(w2056 | w2057);
assign w2058 = v970;
assign v971 = ~(w2024 | w2058);
assign w2059 = v971;
assign w2060 = w2024 & w2058;
assign v972 = ~(w2059 | w2060);
assign w2061 = v972;
assign w2062 = ~w1998 & w2061;
assign w2063 = w1998 & ~w2061;
assign v973 = ~(w2062 | w2063);
assign w2064 = v973;
assign w2065 = ~w1997 & w2064;
assign w2066 = w1997 & ~w2064;
assign v974 = ~(w2065 | w2066);
assign w2067 = v974;
assign v975 = ~(w1950 | w1953);
assign w2068 = v975;
assign v976 = ~(w1884 | w1888);
assign w2069 = v976;
assign v977 = ~(w1887 | w2069);
assign w2070 = v977;
assign v978 = ~(w1872 | w1876);
assign w2071 = v978;
assign v979 = ~(w1875 | w2071);
assign w2072 = v979;
assign w2073 = w2070 & w2072;
assign v980 = ~(w2070 | w2072);
assign w2074 = v980;
assign v981 = ~(w2073 | w2074);
assign w2075 = v981;
assign v982 = ~(w1634 | w1920);
assign w2076 = v982;
assign v983 = ~(w1919 | w2076);
assign w2077 = v983;
assign v984 = ~(w2075 | w2077);
assign w2078 = v984;
assign w2079 = w2075 & w2077;
assign v985 = ~(w2078 | w2079);
assign w2080 = v985;
assign w2081 = pi15 & pi17;
assign w2082 = pi01 & pi31;
assign v986 = ~(w2081 | w2082);
assign w2083 = v986;
assign w2084 = w2081 & w2082;
assign v987 = ~(w2083 | w2084);
assign w2085 = v987;
assign v988 = ~(w1896 | w1900);
assign w2086 = v988;
assign v989 = ~(w1899 | w2086);
assign w2087 = v989;
assign w2088 = w2085 & w2087;
assign v990 = ~(w2085 | w2087);
assign w2089 = v990;
assign v991 = ~(w2088 | w2089);
assign w2090 = v991;
assign v992 = ~(w1905 | w1909);
assign w2091 = v992;
assign v993 = ~(w1908 | w2091);
assign w2092 = v993;
assign w2093 = w2090 & w2092;
assign v994 = ~(w2090 | w2092);
assign w2094 = v994;
assign v995 = ~(w2093 | w2094);
assign w2095 = v995;
assign w2096 = w2080 & w2095;
assign v996 = ~(w2080 | w2095);
assign w2097 = v996;
assign v997 = ~(w2096 | w2097);
assign w2098 = v997;
assign w2099 = w2068 & ~w2098;
assign w2100 = ~w2068 & w2098;
assign v998 = ~(w2099 | w2100);
assign w2101 = v998;
assign v999 = ~(w1914 | w1925);
assign w2102 = v999;
assign w2103 = (~w1881 & ~w1883) | (~w1881 & w17050) | (~w1883 & w17050);
assign v1000 = ~(w1963 | w1969);
assign w2104 = v1000;
assign v1001 = ~(w2103 | w2104);
assign w2105 = v1001;
assign w2106 = w2103 & w2104;
assign v1002 = ~(w2105 | w2106);
assign w2107 = v1002;
assign w2108 = w2102 & ~w2107;
assign w2109 = ~w2102 & w2107;
assign v1003 = ~(w2108 | w2109);
assign w2110 = v1003;
assign v1004 = ~(w1928 | w1931);
assign w2111 = v1004;
assign w2112 = ~w2110 & w2111;
assign w2113 = w2110 & ~w2111;
assign v1005 = ~(w2112 | w2113);
assign w2114 = v1005;
assign w2115 = w2101 & w2114;
assign v1006 = ~(w2101 | w2114);
assign w2116 = v1006;
assign v1007 = ~(w2115 | w2116);
assign w2117 = v1007;
assign w2118 = w2067 & w2117;
assign v1008 = ~(w2067 | w2117);
assign w2119 = v1008;
assign v1009 = ~(w2118 | w2119);
assign w2120 = v1009;
assign w2121 = ~w1996 & w2120;
assign w2122 = w1996 & ~w2120;
assign v1010 = ~(w2121 | w2122);
assign w2123 = v1010;
assign w2124 = w1995 & w2123;
assign v1011 = ~(w1995 | w2123);
assign w2125 = v1011;
assign v1012 = ~(w2124 | w2125);
assign w2126 = v1012;
assign v1013 = ~(w2035 | w2039);
assign w2127 = v1013;
assign v1014 = ~(w2038 | w2127);
assign w2128 = v1014;
assign w2129 = w2025 & ~w2028;
assign v1015 = ~(w2030 | w2129);
assign w2130 = v1015;
assign w2131 = w2128 & ~w2130;
assign w2132 = ~w2128 & w2130;
assign v1016 = ~(w2131 | w2132);
assign w2133 = v1016;
assign v1017 = ~(w2047 | w2051);
assign w2134 = v1017;
assign v1018 = ~(w2050 | w2134);
assign w2135 = v1018;
assign v1019 = ~(w2133 | w2135);
assign w2136 = v1019;
assign w2137 = w2133 & w2135;
assign v1020 = ~(w2136 | w2137);
assign w2138 = v1020;
assign v1021 = ~(w2010 | w2014);
assign w2139 = v1021;
assign v1022 = ~(w2013 | w2139);
assign w2140 = v1022;
assign v1023 = ~(w2001 | w2005);
assign w2141 = v1023;
assign v1024 = ~(w2004 | w2141);
assign w2142 = v1024;
assign w2143 = w2140 & w2142;
assign v1025 = ~(w2140 | w2142);
assign w2144 = v1025;
assign v1026 = ~(w2143 | w2144);
assign w2145 = v1026;
assign w2146 = pi02 & pi31;
assign w2147 = pi00 & pi33;
assign w2148 = pi11 & pi22;
assign v1027 = ~(w2147 | w2148);
assign w2149 = v1027;
assign w2150 = w2147 & w2148;
assign v1028 = ~(w2149 | w2150);
assign w2151 = v1028;
assign w2152 = w2146 & ~w2151;
assign w2153 = ~w2146 & w2151;
assign v1029 = ~(w2152 | w2153);
assign w2154 = v1029;
assign w2155 = ~w2145 & w2154;
assign w2156 = w2145 & ~w2154;
assign v1030 = ~(w2155 | w2156);
assign w2157 = v1030;
assign v1031 = ~(w2138 | w2157);
assign w2158 = v1031;
assign w2159 = w2138 & w2157;
assign v1032 = ~(w2158 | w2159);
assign w2160 = v1032;
assign w2161 = pi03 & pi30;
assign w2162 = pi04 & pi29;
assign w2163 = pi09 & pi24;
assign v1033 = ~(w2162 | w2163);
assign w2164 = v1033;
assign w2165 = w2162 & w2163;
assign v1034 = ~(w2164 | w2165);
assign w2166 = v1034;
assign w2167 = w2161 & ~w2166;
assign w2168 = ~w2161 & w2166;
assign v1035 = ~(w2167 | w2168);
assign w2169 = v1035;
assign w2170 = pi05 & pi28;
assign w2171 = pi08 & pi25;
assign w2172 = pi06 & pi27;
assign v1036 = ~(w2171 | w2172);
assign w2173 = v1036;
assign w2174 = w2171 & w2172;
assign v1037 = ~(w2173 | w2174);
assign w2175 = v1037;
assign w2176 = w2170 & ~w2175;
assign w2177 = ~w2170 & w2175;
assign v1038 = ~(w2176 | w2177);
assign w2178 = v1038;
assign v1039 = ~(w2169 | w2178);
assign w2179 = v1039;
assign w2180 = w2169 & w2178;
assign v1040 = ~(w2179 | w2180);
assign w2181 = v1040;
assign w2182 = pi07 & pi26;
assign w2183 = pi16 & pi17;
assign w2184 = pi15 & pi18;
assign v1041 = ~(w2183 | w2184);
assign w2185 = v1041;
assign w2186 = w2183 & w2184;
assign v1042 = ~(w2185 | w2186);
assign w2187 = v1042;
assign w2188 = w2182 & ~w2187;
assign w2189 = ~w2182 & w2187;
assign v1043 = ~(w2188 | w2189);
assign w2190 = v1043;
assign w2191 = w2181 & ~w2190;
assign w2192 = ~w2181 & w2190;
assign v1044 = ~(w2191 | w2192);
assign w2193 = v1044;
assign v1045 = ~(w2160 | w2193);
assign w2194 = v1045;
assign w2195 = w2160 & w2193;
assign v1046 = ~(w2194 | w2195);
assign w2196 = v1046;
assign v1047 = ~(w2019 | w2023);
assign w2197 = v1047;
assign w2198 = (~w2073 & ~w2075) | (~w2073 & w16838) | (~w2075 & w16838);
assign w2199 = (~w2044 & ~w2046) | (~w2044 & w16717) | (~w2046 & w16717);
assign v1048 = ~(w2198 | w2199);
assign w2200 = v1048;
assign w2201 = w2198 & w2199;
assign v1049 = ~(w2200 | w2201);
assign w2202 = v1049;
assign w2203 = w2197 & ~w2202;
assign w2204 = ~w2197 & w2202;
assign v1050 = ~(w2203 | w2204);
assign w2205 = v1050;
assign w2206 = (~w2060 & w1998) | (~w2060 & w17051) | (w1998 & w17051);
assign w2207 = ~w2205 & w2206;
assign w2208 = w2205 & ~w2206;
assign v1051 = ~(w2207 | w2208);
assign w2209 = v1051;
assign w2210 = w2196 & w2209;
assign v1052 = ~(w2196 | w2209);
assign w2211 = v1052;
assign v1053 = ~(w2210 | w2211);
assign w2212 = v1053;
assign w2213 = (~w2088 & ~w2090) | (~w2088 & w16839) | (~w2090 & w16839);
assign w2214 = pi10 & pi23;
assign v1054 = ~(w2084 | w2214);
assign w2215 = v1054;
assign w2216 = w2084 & w2214;
assign v1055 = ~(w2215 | w2216);
assign w2217 = v1055;
assign w2218 = pi01 & pi32;
assign w2219 = pi17 & w2218;
assign v1056 = ~(pi17 | w2218);
assign w2220 = v1056;
assign v1057 = ~(w2219 | w2220);
assign w2221 = v1057;
assign w2222 = ~w2217 & w2221;
assign w2223 = w2217 & ~w2221;
assign v1058 = ~(w2222 | w2223);
assign w2224 = v1058;
assign w2225 = pi12 & pi21;
assign w2226 = pi13 & pi20;
assign w2227 = pi14 & pi19;
assign v1059 = ~(w2226 | w2227);
assign w2228 = v1059;
assign w2229 = w2226 & w2227;
assign v1060 = ~(w2228 | w2229);
assign w2230 = v1060;
assign w2231 = w2225 & ~w2230;
assign w2232 = ~w2225 & w2230;
assign v1061 = ~(w2231 | w2232);
assign w2233 = v1061;
assign v1062 = ~(w2224 | w2233);
assign w2234 = v1062;
assign w2235 = w2224 & w2233;
assign v1063 = ~(w2234 | w2235);
assign w2236 = v1063;
assign w2237 = w2213 & ~w2236;
assign w2238 = ~w2213 & w2236;
assign v1064 = ~(w2237 | w2238);
assign w2239 = v1064;
assign w2240 = (~w2105 & ~w2107) | (~w2105 & w17052) | (~w2107 & w17052);
assign w2241 = ~w2239 & w2240;
assign w2242 = w2239 & ~w2240;
assign v1065 = ~(w2241 | w2242);
assign w2243 = v1065;
assign w2244 = (~w2096 & w2068) | (~w2096 & w17053) | (w2068 & w17053);
assign w2245 = ~w2243 & w2244;
assign w2246 = w2243 & ~w2244;
assign v1066 = ~(w2245 | w2246);
assign w2247 = v1066;
assign w2248 = (~w2113 & ~w2114) | (~w2113 & w17054) | (~w2114 & w17054);
assign w2249 = ~w2247 & w2248;
assign w2250 = w2247 & ~w2248;
assign v1067 = ~(w2249 | w2250);
assign w2251 = v1067;
assign w2252 = w2212 & w2251;
assign v1068 = ~(w2212 | w2251);
assign w2253 = v1068;
assign v1069 = ~(w2252 | w2253);
assign w2254 = v1069;
assign w2255 = (~w2065 & ~w2067) | (~w2065 & w17055) | (~w2067 & w17055);
assign w2256 = ~w2254 & w2255;
assign w2257 = w2254 & ~w2255;
assign v1070 = ~(w2256 | w2257);
assign w2258 = v1070;
assign v1071 = ~(w1985 | w2121);
assign w2259 = v1071;
assign w2260 = (~w1864 & w16505) | (~w1864 & w16506) | (w16505 & w16506);
assign v1072 = ~(w2122 | w2260);
assign w2261 = v1072;
assign w2262 = w2258 & w2261;
assign v1073 = ~(w2258 | w2261);
assign w2263 = v1073;
assign v1074 = ~(w2262 | w2263);
assign w2264 = v1074;
assign v1075 = ~(w2250 | w2252);
assign w2265 = v1075;
assign w2266 = (~w2208 & ~w2209) | (~w2208 & w17056) | (~w2209 & w17056);
assign w2267 = (~w2143 & ~w2145) | (~w2143 & w17057) | (~w2145 & w17057);
assign w2268 = (~w2131 & ~w2133) | (~w2131 & w16718) | (~w2133 & w16718);
assign w2269 = pi00 & pi34;
assign w2270 = pi03 & pi31;
assign w2271 = pi04 & pi30;
assign v1076 = ~(w2270 | w2271);
assign w2272 = v1076;
assign w2273 = w2270 & w2271;
assign v1077 = ~(w2272 | w2273);
assign w2274 = v1077;
assign w2275 = w2269 & ~w2274;
assign w2276 = ~w2269 & w2274;
assign v1078 = ~(w2275 | w2276);
assign w2277 = v1078;
assign v1079 = ~(w2268 | w2277);
assign w2278 = v1079;
assign w2279 = w2268 & w2277;
assign v1080 = ~(w2278 | w2279);
assign w2280 = v1080;
assign w2281 = ~w2267 & w2280;
assign w2282 = w2267 & ~w2280;
assign v1081 = ~(w2281 | w2282);
assign w2283 = v1081;
assign w2284 = (~w2159 & ~w2160) | (~w2159 & w16840) | (~w2160 & w16840);
assign w2285 = (~w2200 & ~w2202) | (~w2200 & w16841) | (~w2202 & w16841);
assign v1082 = ~(w2284 | w2285);
assign w2286 = v1082;
assign w2287 = w2284 & w2285;
assign v1083 = ~(w2286 | w2287);
assign w2288 = v1083;
assign w2289 = w2283 & w2288;
assign v1084 = ~(w2283 | w2288);
assign w2290 = v1084;
assign v1085 = ~(w2289 | w2290);
assign w2291 = v1085;
assign w2292 = ~w2266 & w2291;
assign w2293 = w2266 & ~w2291;
assign v1086 = ~(w2292 | w2293);
assign w2294 = v1086;
assign v1087 = ~(w2146 | w2150);
assign w2295 = v1087;
assign v1088 = ~(w2149 | w2295);
assign w2296 = v1088;
assign v1089 = ~(w2161 | w2165);
assign w2297 = v1089;
assign v1090 = ~(w2164 | w2297);
assign w2298 = v1090;
assign w2299 = w2296 & w2298;
assign v1091 = ~(w2296 | w2298);
assign w2300 = v1091;
assign v1092 = ~(w2299 | w2300);
assign w2301 = v1092;
assign v1093 = ~(w2170 | w2174);
assign w2302 = v1093;
assign v1094 = ~(w2173 | w2302);
assign w2303 = v1094;
assign v1095 = ~(w2301 | w2303);
assign w2304 = v1095;
assign w2305 = w2301 & w2303;
assign v1096 = ~(w2304 | w2305);
assign w2306 = v1096;
assign w2307 = (~w2179 & ~w2181) | (~w2179 & w16719) | (~w2181 & w16719);
assign w2308 = pi16 & pi18;
assign w2309 = pi01 & pi33;
assign v1097 = ~(w2308 | w2309);
assign w2310 = v1097;
assign w2311 = w2308 & w2309;
assign v1098 = ~(w2310 | w2311);
assign w2312 = v1098;
assign w2313 = w2219 & w2312;
assign v1099 = ~(w2219 | w2312);
assign w2314 = v1099;
assign v1100 = ~(w2313 | w2314);
assign w2315 = v1100;
assign v1101 = ~(w2182 | w2186);
assign w2316 = v1101;
assign v1102 = ~(w2185 | w2316);
assign w2317 = v1102;
assign w2318 = w2315 & w2317;
assign v1103 = ~(w2315 | w2317);
assign w2319 = v1103;
assign v1104 = ~(w2318 | w2319);
assign w2320 = v1104;
assign w2321 = ~w2307 & w2320;
assign w2322 = w2307 & ~w2320;
assign v1105 = ~(w2321 | w2322);
assign w2323 = v1105;
assign w2324 = w2306 & w2323;
assign v1106 = ~(w2306 | w2323);
assign w2325 = v1106;
assign v1107 = ~(w2324 | w2325);
assign w2326 = v1107;
assign v1108 = ~(w2225 | w2229);
assign w2327 = v1108;
assign v1109 = ~(w2228 | w2327);
assign w2328 = v1109;
assign v1110 = ~(w2216 | w2221);
assign w2329 = v1110;
assign v1111 = ~(w2215 | w2329);
assign w2330 = v1111;
assign w2331 = w2328 & w2330;
assign v1112 = ~(w2328 | w2330);
assign w2332 = v1112;
assign v1113 = ~(w2331 | w2332);
assign w2333 = v1113;
assign w2334 = pi12 & pi22;
assign v1114 = ~(w1129 | w2334);
assign w2335 = v1114;
assign w2336 = w1129 & w2334;
assign v1115 = ~(w2335 | w2336);
assign w2337 = v1115;
assign w2338 = w2029 & ~w2337;
assign w2339 = ~w2029 & w2337;
assign v1116 = ~(w2338 | w2339);
assign w2340 = v1116;
assign w2341 = ~w2333 & w2340;
assign w2342 = w2333 & ~w2340;
assign v1117 = ~(w2341 | w2342);
assign w2343 = v1117;
assign w2344 = (~w2234 & ~w2236) | (~w2234 & w16842) | (~w2236 & w16842);
assign w2345 = w2343 & ~w2344;
assign w2346 = ~w2343 & w2344;
assign v1118 = ~(w2345 | w2346);
assign w2347 = v1118;
assign w2348 = pi10 & pi24;
assign w2349 = pi05 & pi29;
assign w2350 = pi09 & pi25;
assign v1119 = ~(w2349 | w2350);
assign w2351 = v1119;
assign w2352 = w2349 & w2350;
assign v1120 = ~(w2351 | w2352);
assign w2353 = v1120;
assign w2354 = w2348 & ~w2353;
assign w2355 = ~w2348 & w2353;
assign v1121 = ~(w2354 | w2355);
assign w2356 = v1121;
assign w2357 = pi13 & pi21;
assign w2358 = pi14 & pi20;
assign w2359 = pi15 & pi19;
assign v1122 = ~(w2358 | w2359);
assign w2360 = v1122;
assign w2361 = w2358 & w2359;
assign v1123 = ~(w2360 | w2361);
assign w2362 = v1123;
assign w2363 = w2357 & ~w2362;
assign w2364 = ~w2357 & w2362;
assign v1124 = ~(w2363 | w2364);
assign w2365 = v1124;
assign v1125 = ~(w2356 | w2365);
assign w2366 = v1125;
assign w2367 = w2356 & w2365;
assign v1126 = ~(w2366 | w2367);
assign w2368 = v1126;
assign w2369 = pi06 & pi28;
assign w2370 = pi08 & pi26;
assign w2371 = pi07 & pi27;
assign v1127 = ~(w2370 | w2371);
assign w2372 = v1127;
assign w2373 = w2370 & w2371;
assign v1128 = ~(w2372 | w2373);
assign w2374 = v1128;
assign w2375 = w2369 & ~w2374;
assign w2376 = ~w2369 & w2374;
assign v1129 = ~(w2375 | w2376);
assign w2377 = v1129;
assign w2378 = w2368 & ~w2377;
assign w2379 = ~w2368 & w2377;
assign v1130 = ~(w2378 | w2379);
assign w2380 = v1130;
assign w2381 = w2347 & w2380;
assign v1131 = ~(w2347 | w2380);
assign w2382 = v1131;
assign v1132 = ~(w2381 | w2382);
assign w2383 = v1132;
assign w2384 = w2326 & w2383;
assign v1133 = ~(w2326 | w2383);
assign w2385 = v1133;
assign v1134 = ~(w2384 | w2385);
assign w2386 = v1134;
assign v1135 = ~(w2242 | w2246);
assign w2387 = v1135;
assign w2388 = w2386 & ~w2387;
assign w2389 = ~w2386 & w2387;
assign v1136 = ~(w2388 | w2389);
assign w2390 = v1136;
assign w2391 = w2294 & w2390;
assign v1137 = ~(w2294 | w2390);
assign w2392 = v1137;
assign v1138 = ~(w2391 | w2392);
assign w2393 = v1138;
assign w2394 = ~w2265 & w2393;
assign w2395 = w2265 & ~w2393;
assign v1139 = ~(w2394 | w2395);
assign w2396 = v1139;
assign w2397 = (~w2257 & w2260) | (~w2257 & w16507) | (w2260 & w16507);
assign v1140 = ~(w2256 | w2397);
assign w2398 = v1140;
assign w2399 = w2396 & w2398;
assign v1141 = ~(w2396 | w2398);
assign w2400 = v1141;
assign v1142 = ~(w2399 | w2400);
assign w2401 = v1142;
assign v1143 = ~(w2256 | w2395);
assign w2402 = v1143;
assign w2403 = (~w2260 & w16508) | (~w2260 & w16509) | (w16508 & w16509);
assign v1144 = ~(w2394 | w2403);
assign w2404 = v1144;
assign v1145 = ~(w2292 | w2391);
assign w2405 = v1145;
assign v1146 = ~(w2384 | w2388);
assign w2406 = v1146;
assign w2407 = (~w2331 & ~w2333) | (~w2331 & w17058) | (~w2333 & w17058);
assign w2408 = (~w2299 & ~w2301) | (~w2299 & w16843) | (~w2301 & w16843);
assign w2409 = (~w2313 & ~w2315) | (~w2313 & w17059) | (~w2315 & w17059);
assign v1147 = ~(w2408 | w2409);
assign w2410 = v1147;
assign w2411 = w2408 & w2409;
assign v1148 = ~(w2410 | w2411);
assign w2412 = v1148;
assign w2413 = w2407 & ~w2412;
assign w2414 = ~w2407 & w2412;
assign v1149 = ~(w2413 | w2414);
assign w2415 = v1149;
assign w2416 = (~w2321 & ~w2323) | (~w2321 & w16844) | (~w2323 & w16844);
assign w2417 = ~w2415 & w2416;
assign w2418 = w2415 & ~w2416;
assign v1150 = ~(w2417 | w2418);
assign w2419 = v1150;
assign w2420 = (~w2345 & ~w2347) | (~w2345 & w17060) | (~w2347 & w17060);
assign w2421 = w2419 & ~w2420;
assign w2422 = ~w2419 & w2420;
assign v1151 = ~(w2421 | w2422);
assign w2423 = v1151;
assign w2424 = ~w2406 & w2423;
assign w2425 = w2406 & ~w2423;
assign v1152 = ~(w2424 | w2425);
assign w2426 = v1152;
assign w2427 = (~w2286 & ~w2288) | (~w2286 & w17061) | (~w2288 & w17061);
assign v1153 = ~(w2029 | w2336);
assign w2428 = v1153;
assign v1154 = ~(w2335 | w2428);
assign w2429 = v1154;
assign v1155 = ~(w2357 | w2361);
assign w2430 = v1155;
assign v1156 = ~(w2360 | w2430);
assign w2431 = v1156;
assign w2432 = w2429 & w2431;
assign v1157 = ~(w2429 | w2431);
assign w2433 = v1157;
assign v1158 = ~(w2432 | w2433);
assign w2434 = v1158;
assign v1159 = ~(w2269 | w2273);
assign w2435 = v1159;
assign v1160 = ~(w2272 | w2435);
assign w2436 = v1160;
assign v1161 = ~(w2434 | w2436);
assign w2437 = v1161;
assign w2438 = w2434 & w2436;
assign v1162 = ~(w2437 | w2438);
assign w2439 = v1162;
assign w2440 = (~w2366 & ~w2368) | (~w2366 & w16845) | (~w2368 & w16845);
assign w2441 = pi34 & w684;
assign w2442 = pi01 & pi34;
assign v1163 = ~(pi18 | w2442);
assign w2443 = v1163;
assign v1164 = ~(w2441 | w2443);
assign w2444 = v1164;
assign v1165 = ~(w2369 | w2373);
assign w2445 = v1165;
assign v1166 = ~(w2372 | w2445);
assign w2446 = v1166;
assign w2447 = w2444 & w2446;
assign v1167 = ~(w2444 | w2446);
assign w2448 = v1167;
assign v1168 = ~(w2447 | w2448);
assign w2449 = v1168;
assign v1169 = ~(w2348 | w2352);
assign w2450 = v1169;
assign v1170 = ~(w2351 | w2450);
assign w2451 = v1170;
assign w2452 = w2449 & w2451;
assign v1171 = ~(w2449 | w2451);
assign w2453 = v1171;
assign v1172 = ~(w2452 | w2453);
assign w2454 = v1172;
assign w2455 = ~w2440 & w2454;
assign w2456 = w2440 & ~w2454;
assign v1173 = ~(w2455 | w2456);
assign w2457 = v1173;
assign w2458 = w2439 & w2457;
assign v1174 = ~(w2439 | w2457);
assign w2459 = v1174;
assign v1175 = ~(w2458 | w2459);
assign w2460 = v1175;
assign w2461 = ~w2427 & w2460;
assign w2462 = w2427 & ~w2460;
assign v1176 = ~(w2461 | w2462);
assign w2463 = v1176;
assign w2464 = (~w2278 & ~w2280) | (~w2278 & w16846) | (~w2280 & w16846);
assign w2465 = pi07 & pi28;
assign w2466 = pi17 & pi18;
assign w2467 = pi16 & pi19;
assign v1177 = ~(w2466 | w2467);
assign w2468 = v1177;
assign w2469 = w2466 & w2467;
assign v1178 = ~(w2468 | w2469);
assign w2470 = v1178;
assign w2471 = w2465 & ~w2470;
assign w2472 = ~w2465 & w2470;
assign v1179 = ~(w2471 | w2472);
assign w2473 = v1179;
assign w2474 = pi05 & pi30;
assign w2475 = pi08 & pi27;
assign w2476 = pi06 & pi29;
assign v1180 = ~(w2475 | w2476);
assign w2477 = v1180;
assign w2478 = w2475 & w2476;
assign v1181 = ~(w2477 | w2478);
assign w2479 = v1181;
assign w2480 = w2474 & ~w2479;
assign w2481 = ~w2474 & w2479;
assign v1182 = ~(w2480 | w2481);
assign w2482 = v1182;
assign v1183 = ~(w2473 | w2482);
assign w2483 = v1183;
assign w2484 = w2473 & w2482;
assign v1184 = ~(w2483 | w2484);
assign w2485 = v1184;
assign w2486 = pi04 & pi31;
assign w2487 = pi09 & pi26;
assign w2488 = pi10 & pi25;
assign v1185 = ~(w2487 | w2488);
assign w2489 = v1185;
assign w2490 = w2487 & w2488;
assign v1186 = ~(w2489 | w2490);
assign w2491 = v1186;
assign w2492 = w2486 & ~w2491;
assign w2493 = ~w2486 & w2491;
assign v1187 = ~(w2492 | w2493);
assign w2494 = v1187;
assign w2495 = w2485 & ~w2494;
assign w2496 = ~w2485 & w2494;
assign v1188 = ~(w2495 | w2496);
assign w2497 = v1188;
assign w2498 = ~w2464 & w2497;
assign w2499 = w2464 & ~w2497;
assign v1189 = ~(w2498 | w2499);
assign w2500 = v1189;
assign w2501 = pi00 & pi35;
assign w2502 = pi02 & pi33;
assign v1190 = ~(w2501 | w2502);
assign w2503 = v1190;
assign w2504 = pi02 & pi35;
assign w2505 = w2147 & w2504;
assign v1191 = ~(w2503 | w2505);
assign w2506 = v1191;
assign w2507 = w2311 & ~w2506;
assign w2508 = ~w2311 & w2506;
assign v1192 = ~(w2507 | w2508);
assign w2509 = v1192;
assign w2510 = pi03 & pi32;
assign w2511 = pi12 & pi23;
assign w2512 = pi11 & pi24;
assign v1193 = ~(w2511 | w2512);
assign w2513 = v1193;
assign w2514 = w2511 & w2512;
assign v1194 = ~(w2513 | w2514);
assign w2515 = v1194;
assign w2516 = w2510 & ~w2515;
assign w2517 = ~w2510 & w2515;
assign v1195 = ~(w2516 | w2517);
assign w2518 = v1195;
assign v1196 = ~(w2509 | w2518);
assign w2519 = v1196;
assign w2520 = w2509 & w2518;
assign v1197 = ~(w2519 | w2520);
assign w2521 = v1197;
assign w2522 = pi13 & pi22;
assign w2523 = pi15 & pi20;
assign w2524 = pi14 & pi21;
assign v1198 = ~(w2523 | w2524);
assign w2525 = v1198;
assign w2526 = w2523 & w2524;
assign v1199 = ~(w2525 | w2526);
assign w2527 = v1199;
assign w2528 = w2522 & ~w2527;
assign w2529 = ~w2522 & w2527;
assign v1200 = ~(w2528 | w2529);
assign w2530 = v1200;
assign w2531 = w2521 & ~w2530;
assign w2532 = ~w2521 & w2530;
assign v1201 = ~(w2531 | w2532);
assign w2533 = v1201;
assign w2534 = w2500 & w2533;
assign v1202 = ~(w2500 | w2533);
assign w2535 = v1202;
assign v1203 = ~(w2534 | w2535);
assign w2536 = v1203;
assign w2537 = w2463 & w2536;
assign v1204 = ~(w2463 | w2536);
assign w2538 = v1204;
assign v1205 = ~(w2537 | w2538);
assign w2539 = v1205;
assign v1206 = ~(w2426 | w2539);
assign w2540 = v1206;
assign w2541 = w2426 & w2539;
assign v1207 = ~(w2540 | w2541);
assign w2542 = v1207;
assign w2543 = w2405 & ~w2542;
assign w2544 = ~w2405 & w2542;
assign v1208 = ~(w2543 | w2544);
assign w2545 = v1208;
assign w2546 = w2404 & w2545;
assign v1209 = ~(w2404 | w2545);
assign w2547 = v1209;
assign v1210 = ~(w2546 | w2547);
assign w2548 = v1210;
assign w2549 = (~w2424 & ~w2426) | (~w2424 & w16847) | (~w2426 & w16847);
assign w2550 = (~w2461 & ~w2463) | (~w2461 & w16848) | (~w2463 & w16848);
assign w2551 = (~w2519 & ~w2521) | (~w2519 & w16849) | (~w2521 & w16849);
assign w2552 = (~w2432 & ~w2434) | (~w2432 & w16720) | (~w2434 & w16720);
assign w2553 = (~w2447 & ~w2449) | (~w2447 & w16721) | (~w2449 & w16721);
assign v1211 = ~(w2552 | w2553);
assign w2554 = v1211;
assign w2555 = w2552 & w2553;
assign v1212 = ~(w2554 | w2555);
assign w2556 = v1212;
assign w2557 = w2551 & ~w2556;
assign w2558 = ~w2551 & w2556;
assign v1213 = ~(w2557 | w2558);
assign w2559 = v1213;
assign w2560 = (~w2455 & ~w2457) | (~w2455 & w16850) | (~w2457 & w16850);
assign w2561 = ~w2559 & w2560;
assign w2562 = w2559 & ~w2560;
assign v1214 = ~(w2561 | w2562);
assign w2563 = v1214;
assign w2564 = (~w2498 & ~w2500) | (~w2498 & w16851) | (~w2500 & w16851);
assign w2565 = w2563 & ~w2564;
assign w2566 = ~w2563 & w2564;
assign v1215 = ~(w2565 | w2566);
assign w2567 = v1215;
assign w2568 = ~w2550 & w2567;
assign w2569 = w2550 & ~w2567;
assign v1216 = ~(w2568 | w2569);
assign w2570 = v1216;
assign w2571 = pi02 & pi34;
assign w2572 = pi12 & pi24;
assign w2573 = pi13 & pi23;
assign v1217 = ~(w2572 | w2573);
assign w2574 = v1217;
assign w2575 = w2572 & w2573;
assign v1218 = ~(w2574 | w2575);
assign w2576 = v1218;
assign w2577 = w2571 & ~w2576;
assign w2578 = ~w2571 & w2576;
assign v1219 = ~(w2577 | w2578);
assign w2579 = v1219;
assign w2580 = pi10 & pi26;
assign w2581 = pi05 & pi31;
assign w2582 = pi09 & pi27;
assign v1220 = ~(w2581 | w2582);
assign w2583 = v1220;
assign w2584 = w2581 & w2582;
assign v1221 = ~(w2583 | w2584);
assign w2585 = v1221;
assign w2586 = w2580 & ~w2585;
assign w2587 = ~w2580 & w2585;
assign v1222 = ~(w2586 | w2587);
assign w2588 = v1222;
assign v1223 = ~(w2579 | w2588);
assign w2589 = v1223;
assign w2590 = w2579 & w2588;
assign v1224 = ~(w2589 | w2590);
assign w2591 = v1224;
assign w2592 = pi06 & pi30;
assign w2593 = pi08 & pi28;
assign w2594 = pi07 & pi29;
assign v1225 = ~(w2593 | w2594);
assign w2595 = v1225;
assign w2596 = w2593 & w2594;
assign v1226 = ~(w2595 | w2596);
assign w2597 = v1226;
assign w2598 = w2592 & ~w2597;
assign w2599 = ~w2592 & w2597;
assign v1227 = ~(w2598 | w2599);
assign w2600 = v1227;
assign w2601 = w2591 & ~w2600;
assign w2602 = ~w2591 & w2600;
assign v1228 = ~(w2601 | w2602);
assign w2603 = v1228;
assign w2604 = (~w2410 & ~w2412) | (~w2410 & w17062) | (~w2412 & w17062);
assign w2605 = pi00 & pi36;
assign w2606 = w2441 & w2605;
assign v1229 = ~(w2441 | w2605);
assign w2607 = v1229;
assign v1230 = ~(w2606 | w2607);
assign w2608 = v1230;
assign w2609 = pi17 & pi19;
assign w2610 = pi01 & pi35;
assign v1231 = ~(w2609 | w2610);
assign w2611 = v1231;
assign w2612 = w2609 & w2610;
assign v1232 = ~(w2611 | w2612);
assign w2613 = v1232;
assign w2614 = w2608 & w2613;
assign v1233 = ~(w2608 | w2613);
assign w2615 = v1233;
assign v1234 = ~(w2614 | w2615);
assign w2616 = v1234;
assign w2617 = pi03 & pi33;
assign w2618 = pi04 & pi32;
assign w2619 = pi11 & pi25;
assign v1235 = ~(w2618 | w2619);
assign w2620 = v1235;
assign w2621 = w2618 & w2619;
assign v1236 = ~(w2620 | w2621);
assign w2622 = v1236;
assign w2623 = w2617 & ~w2622;
assign w2624 = ~w2617 & w2622;
assign v1237 = ~(w2623 | w2624);
assign w2625 = v1237;
assign w2626 = pi14 & pi22;
assign w2627 = pi15 & pi21;
assign w2628 = pi16 & pi20;
assign v1238 = ~(w2627 | w2628);
assign w2629 = v1238;
assign w2630 = w2627 & w2628;
assign v1239 = ~(w2629 | w2630);
assign w2631 = v1239;
assign w2632 = w2626 & ~w2631;
assign w2633 = ~w2626 & w2631;
assign v1240 = ~(w2632 | w2633);
assign w2634 = v1240;
assign v1241 = ~(w2625 | w2634);
assign w2635 = v1241;
assign w2636 = w2625 & w2634;
assign v1242 = ~(w2635 | w2636);
assign w2637 = v1242;
assign w2638 = w2616 & w2637;
assign v1243 = ~(w2616 | w2637);
assign w2639 = v1243;
assign v1244 = ~(w2638 | w2639);
assign w2640 = v1244;
assign w2641 = ~w2604 & w2640;
assign w2642 = w2604 & ~w2640;
assign v1245 = ~(w2641 | w2642);
assign w2643 = v1245;
assign w2644 = w2603 & w2643;
assign v1246 = ~(w2603 | w2643);
assign w2645 = v1246;
assign v1247 = ~(w2644 | w2645);
assign w2646 = v1247;
assign v1248 = ~(w2486 | w2490);
assign w2647 = v1248;
assign v1249 = ~(w2489 | w2647);
assign w2648 = v1249;
assign v1250 = ~(w2474 | w2478);
assign w2649 = v1250;
assign v1251 = ~(w2477 | w2649);
assign w2650 = v1251;
assign w2651 = w2648 & w2650;
assign v1252 = ~(w2648 | w2650);
assign w2652 = v1252;
assign v1253 = ~(w2651 | w2652);
assign w2653 = v1253;
assign v1254 = ~(w2465 | w2469);
assign w2654 = v1254;
assign v1255 = ~(w2468 | w2654);
assign w2655 = v1255;
assign v1256 = ~(w2653 | w2655);
assign w2656 = v1256;
assign w2657 = w2653 & w2655;
assign v1257 = ~(w2656 | w2657);
assign w2658 = v1257;
assign v1258 = ~(w2522 | w2526);
assign w2659 = v1258;
assign v1259 = ~(w2525 | w2659);
assign w2660 = v1259;
assign v1260 = ~(w2510 | w2514);
assign w2661 = v1260;
assign v1261 = ~(w2513 | w2661);
assign w2662 = v1261;
assign w2663 = w2660 & w2662;
assign v1262 = ~(w2660 | w2662);
assign w2664 = v1262;
assign v1263 = ~(w2663 | w2664);
assign w2665 = v1263;
assign w2666 = w2311 & ~w2503;
assign v1264 = ~(w2505 | w2666);
assign w2667 = v1264;
assign w2668 = ~w2665 & w2667;
assign w2669 = w2665 & ~w2667;
assign v1265 = ~(w2668 | w2669);
assign w2670 = v1265;
assign w2671 = (~w2483 & ~w2485) | (~w2483 & w17063) | (~w2485 & w17063);
assign w2672 = ~w2670 & w2671;
assign w2673 = w2670 & ~w2671;
assign v1266 = ~(w2672 | w2673);
assign w2674 = v1266;
assign w2675 = w2658 & w2674;
assign v1267 = ~(w2658 | w2674);
assign w2676 = v1267;
assign v1268 = ~(w2675 | w2676);
assign w2677 = v1268;
assign w2678 = (w2677 & w2421) | (w2677 & w16852) | (w2421 & w16852);
assign w2679 = ~w2421 & w16853;
assign v1269 = ~(w2678 | w2679);
assign w2680 = v1269;
assign w2681 = w2646 & w2680;
assign v1270 = ~(w2646 | w2680);
assign w2682 = v1270;
assign v1271 = ~(w2681 | w2682);
assign w2683 = v1271;
assign w2684 = w2570 & w2683;
assign v1272 = ~(w2570 | w2683);
assign w2685 = v1272;
assign v1273 = ~(w2684 | w2685);
assign w2686 = v1273;
assign w2687 = w2549 & ~w2686;
assign w2688 = ~w2549 & w2686;
assign v1274 = ~(w2687 | w2688);
assign w2689 = v1274;
assign v1275 = ~(w2394 | w2544);
assign w2690 = v1275;
assign w2691 = (~w2260 & w16510) | (~w2260 & w16511) | (w16510 & w16511);
assign w2692 = w2689 & w2691;
assign v1276 = ~(w2689 | w2691);
assign w2693 = v1276;
assign v1277 = ~(w2692 | w2693);
assign w2694 = v1277;
assign v1278 = ~(w2568 | w2684);
assign w2695 = v1278;
assign w2696 = (~w2663 & ~w2665) | (~w2663 & w17064) | (~w2665 & w17064);
assign w2697 = pi08 & pi29;
assign w2698 = pi18 & pi19;
assign w2699 = pi17 & pi20;
assign v1279 = ~(w2698 | w2699);
assign w2700 = v1279;
assign w2701 = w2698 & w2699;
assign v1280 = ~(w2700 | w2701);
assign w2702 = v1280;
assign w2703 = w2697 & ~w2702;
assign w2704 = ~w2697 & w2702;
assign v1281 = ~(w2703 | w2704);
assign w2705 = v1281;
assign w2706 = pi11 & pi26;
assign w2707 = pi05 & pi32;
assign w2708 = pi10 & pi27;
assign v1282 = ~(w2707 | w2708);
assign w2709 = v1282;
assign w2710 = w2707 & w2708;
assign v1283 = ~(w2709 | w2710);
assign w2711 = v1283;
assign w2712 = w2706 & ~w2711;
assign w2713 = ~w2706 & w2711;
assign v1284 = ~(w2712 | w2713);
assign w2714 = v1284;
assign v1285 = ~(w2705 | w2714);
assign w2715 = v1285;
assign w2716 = w2705 & w2714;
assign v1286 = ~(w2715 | w2716);
assign w2717 = v1286;
assign w2718 = w2696 & ~w2717;
assign w2719 = ~w2696 & w2717;
assign v1287 = ~(w2718 | w2719);
assign w2720 = v1287;
assign w2721 = (~w2554 & ~w2556) | (~w2554 & w16854) | (~w2556 & w16854);
assign w2722 = ~w2720 & w2721;
assign w2723 = w2720 & ~w2721;
assign v1288 = ~(w2722 | w2723);
assign w2724 = v1288;
assign w2725 = pi16 & pi21;
assign w2726 = pi03 & pi34;
assign v1289 = ~(w2504 | w2726);
assign w2727 = v1289;
assign w2728 = pi03 & pi35;
assign w2729 = w2571 & w2728;
assign v1290 = ~(w2727 | w2729);
assign w2730 = v1290;
assign w2731 = w2725 & ~w2730;
assign w2732 = ~w2725 & w2730;
assign v1291 = ~(w2731 | w2732);
assign w2733 = v1291;
assign w2734 = pi00 & pi37;
assign w2735 = pi12 & pi25;
assign w2736 = pi04 & pi33;
assign v1292 = ~(w2735 | w2736);
assign w2737 = v1292;
assign w2738 = w2735 & w2736;
assign v1293 = ~(w2737 | w2738);
assign w2739 = v1293;
assign w2740 = w2734 & ~w2739;
assign w2741 = ~w2734 & w2739;
assign v1294 = ~(w2740 | w2741);
assign w2742 = v1294;
assign v1295 = ~(w2733 | w2742);
assign w2743 = v1295;
assign w2744 = w2733 & w2742;
assign v1296 = ~(w2743 | w2744);
assign w2745 = v1296;
assign w2746 = pi09 & pi28;
assign w2747 = pi06 & pi31;
assign w2748 = pi07 & pi30;
assign v1297 = ~(w2747 | w2748);
assign w2749 = v1297;
assign w2750 = w2747 & w2748;
assign v1298 = ~(w2749 | w2750);
assign w2751 = v1298;
assign w2752 = w2746 & ~w2751;
assign w2753 = ~w2746 & w2751;
assign v1299 = ~(w2752 | w2753);
assign w2754 = v1299;
assign w2755 = w2745 & ~w2754;
assign w2756 = ~w2745 & w2754;
assign v1300 = ~(w2755 | w2756);
assign w2757 = v1300;
assign v1301 = ~(w2724 | w2757);
assign w2758 = v1301;
assign w2759 = w2724 & w2757;
assign v1302 = ~(w2758 | w2759);
assign w2760 = v1302;
assign w2761 = (~w2606 & ~w2608) | (~w2606 & w16855) | (~w2608 & w16855);
assign v1303 = ~(w2580 | w2584);
assign w2762 = v1303;
assign v1304 = ~(w2583 | w2762);
assign w2763 = v1304;
assign w2764 = ~w2761 & w2763;
assign w2765 = w2761 & ~w2763;
assign v1305 = ~(w2764 | w2765);
assign w2766 = v1305;
assign w2767 = pi13 & pi24;
assign w2768 = pi14 & pi23;
assign w2769 = pi15 & pi22;
assign v1306 = ~(w2768 | w2769);
assign w2770 = v1306;
assign w2771 = w2768 & w2769;
assign v1307 = ~(w2770 | w2771);
assign w2772 = v1307;
assign w2773 = w2767 & ~w2772;
assign w2774 = ~w2767 & w2772;
assign v1308 = ~(w2773 | w2774);
assign w2775 = v1308;
assign w2776 = ~w2766 & w2775;
assign w2777 = w2766 & ~w2775;
assign v1309 = ~(w2776 | w2777);
assign w2778 = v1309;
assign v1310 = ~(w2626 | w2630);
assign w2779 = v1310;
assign v1311 = ~(w2629 | w2779);
assign w2780 = v1311;
assign v1312 = ~(w2617 | w2621);
assign w2781 = v1312;
assign v1313 = ~(w2620 | w2781);
assign w2782 = v1313;
assign w2783 = w2780 & w2782;
assign v1314 = ~(w2780 | w2782);
assign w2784 = v1314;
assign v1315 = ~(w2783 | w2784);
assign w2785 = v1315;
assign v1316 = ~(w2571 | w2575);
assign w2786 = v1316;
assign v1317 = ~(w2574 | w2786);
assign w2787 = v1317;
assign v1318 = ~(w2785 | w2787);
assign w2788 = v1318;
assign w2789 = w2785 & w2787;
assign v1319 = ~(w2788 | w2789);
assign w2790 = v1319;
assign v1320 = ~(w2635 | w2638);
assign w2791 = v1320;
assign w2792 = ~w2790 & w2791;
assign w2793 = w2790 & ~w2791;
assign v1321 = ~(w2792 | w2793);
assign w2794 = v1321;
assign w2795 = w2778 & w2794;
assign v1322 = ~(w2778 | w2794);
assign w2796 = v1322;
assign v1323 = ~(w2795 | w2796);
assign w2797 = v1323;
assign w2798 = (w2797 & w2565) | (w2797 & w17065) | (w2565 & w17065);
assign w2799 = ~w2565 & w17066;
assign v1324 = ~(w2798 | w2799);
assign w2800 = v1324;
assign w2801 = w2760 & w2800;
assign v1325 = ~(w2760 | w2800);
assign w2802 = v1325;
assign v1326 = ~(w2801 | w2802);
assign w2803 = v1326;
assign w2804 = (~w2678 & ~w2680) | (~w2678 & w17067) | (~w2680 & w17067);
assign v1327 = ~(w2641 | w2644);
assign w2805 = v1327;
assign v1328 = ~(w2673 | w2675);
assign w2806 = v1328;
assign v1329 = ~(w2589 | w2601);
assign w2807 = v1329;
assign w2808 = (~w2651 & ~w2653) | (~w2651 & w17068) | (~w2653 & w17068);
assign w2809 = ~pi36 & w2612;
assign w2810 = pi36 & w792;
assign w2811 = pi01 & pi36;
assign v1330 = ~(pi19 | w2811);
assign w2812 = v1330;
assign v1331 = ~(w2810 | w2812);
assign w2813 = v1331;
assign v1332 = ~(w2612 | w2813);
assign w2814 = v1332;
assign v1333 = ~(w2809 | w2814);
assign w2815 = v1333;
assign v1334 = ~(w2592 | w2596);
assign w2816 = v1334;
assign v1335 = ~(w2595 | w2816);
assign w2817 = v1335;
assign w2818 = w2815 & w2817;
assign v1336 = ~(w2815 | w2817);
assign w2819 = v1336;
assign v1337 = ~(w2818 | w2819);
assign w2820 = v1337;
assign w2821 = ~w2808 & w2820;
assign w2822 = w2808 & ~w2820;
assign v1338 = ~(w2821 | w2822);
assign w2823 = v1338;
assign w2824 = ~w2807 & w2823;
assign w2825 = w2807 & ~w2823;
assign v1339 = ~(w2824 | w2825);
assign w2826 = v1339;
assign w2827 = ~w2806 & w2826;
assign w2828 = w2806 & ~w2826;
assign v1340 = ~(w2827 | w2828);
assign w2829 = v1340;
assign w2830 = ~w2805 & w2829;
assign w2831 = w2805 & ~w2829;
assign v1341 = ~(w2830 | w2831);
assign w2832 = v1341;
assign w2833 = ~w2804 & w2832;
assign w2834 = w2804 & ~w2832;
assign v1342 = ~(w2833 | w2834);
assign w2835 = v1342;
assign w2836 = w2803 & w2835;
assign v1343 = ~(w2803 | w2835);
assign w2837 = v1343;
assign v1344 = ~(w2836 | w2837);
assign w2838 = v1344;
assign w2839 = ~w2695 & w2838;
assign w2840 = w2695 & ~w2838;
assign v1345 = ~(w2839 | w2840);
assign w2841 = v1345;
assign v1346 = ~(w2688 | w2691);
assign w2842 = v1346;
assign v1347 = ~(w2687 | w2842);
assign w2843 = v1347;
assign w2844 = w2841 & w2843;
assign v1348 = ~(w2841 | w2843);
assign w2845 = v1348;
assign v1349 = ~(w2844 | w2845);
assign w2846 = v1349;
assign v1350 = ~(w2833 | w2836);
assign w2847 = v1350;
assign v1351 = ~(w2827 | w2830);
assign w2848 = v1351;
assign w2849 = pi18 & pi20;
assign w2850 = pi01 & pi37;
assign v1352 = ~(w2849 | w2850);
assign w2851 = v1352;
assign w2852 = w2849 & w2850;
assign v1353 = ~(w2851 | w2852);
assign w2853 = v1353;
assign v1354 = ~(w2697 | w2701);
assign w2854 = v1354;
assign v1355 = ~(w2700 | w2854);
assign w2855 = v1355;
assign w2856 = w2853 & w2855;
assign v1356 = ~(w2853 | w2855);
assign w2857 = v1356;
assign v1357 = ~(w2856 | w2857);
assign w2858 = v1357;
assign v1358 = ~(w2746 | w2750);
assign w2859 = v1358;
assign v1359 = ~(w2749 | w2859);
assign w2860 = v1359;
assign w2861 = w2858 & w2860;
assign v1360 = ~(w2858 | w2860);
assign w2862 = v1360;
assign v1361 = ~(w2861 | w2862);
assign w2863 = v1361;
assign w2864 = (~w2764 & ~w2766) | (~w2764 & w17069) | (~w2766 & w17069);
assign w2865 = (~w2743 & ~w2745) | (~w2743 & w17070) | (~w2745 & w17070);
assign v1362 = ~(w2864 | w2865);
assign w2866 = v1362;
assign w2867 = w2864 & w2865;
assign v1363 = ~(w2866 | w2867);
assign w2868 = v1363;
assign w2869 = w2863 & w2868;
assign v1364 = ~(w2863 | w2868);
assign w2870 = v1364;
assign v1365 = ~(w2869 | w2870);
assign w2871 = v1365;
assign w2872 = ~w2848 & w2871;
assign w2873 = w2848 & ~w2871;
assign v1366 = ~(w2872 | w2873);
assign w2874 = v1366;
assign w2875 = (~w2783 & ~w2785) | (~w2783 & w17071) | (~w2785 & w17071);
assign w2876 = (~w2809 & ~w2815) | (~w2809 & w16856) | (~w2815 & w16856);
assign w2877 = pi12 & pi26;
assign w2878 = pi04 & pi34;
assign w2879 = pi11 & pi27;
assign v1367 = ~(w2878 | w2879);
assign w2880 = v1367;
assign w2881 = w2878 & w2879;
assign v1368 = ~(w2880 | w2881);
assign w2882 = v1368;
assign w2883 = w2877 & ~w2882;
assign w2884 = ~w2877 & w2882;
assign v1369 = ~(w2883 | w2884);
assign w2885 = v1369;
assign v1370 = ~(w2876 | w2885);
assign w2886 = v1370;
assign w2887 = w2876 & w2885;
assign v1371 = ~(w2886 | w2887);
assign w2888 = v1371;
assign w2889 = w2875 & ~w2888;
assign w2890 = ~w2875 & w2888;
assign v1372 = ~(w2889 | w2890);
assign w2891 = v1372;
assign v1373 = ~(w2821 | w2824);
assign w2892 = v1373;
assign v1374 = ~(w2706 | w2710);
assign w2893 = v1374;
assign v1375 = ~(w2709 | w2893);
assign w2894 = v1375;
assign w2895 = pi00 & pi38;
assign w2896 = pi02 & pi36;
assign v1376 = ~(w2895 | w2896);
assign w2897 = v1376;
assign w2898 = pi02 & pi38;
assign w2899 = w2605 & w2898;
assign v1377 = ~(w2897 | w2899);
assign w2900 = v1377;
assign w2901 = w2810 & ~w2900;
assign w2902 = ~w2810 & w2900;
assign v1378 = ~(w2901 | w2902);
assign w2903 = v1378;
assign w2904 = w2894 & ~w2903;
assign w2905 = ~w2894 & w2903;
assign v1379 = ~(w2904 | w2905);
assign w2906 = v1379;
assign w2907 = pi13 & pi25;
assign w2908 = pi14 & pi24;
assign v1380 = ~(w2907 | w2908);
assign w2909 = v1380;
assign w2910 = w2907 & w2908;
assign v1381 = ~(w2909 | w2910);
assign w2911 = v1381;
assign w2912 = w2728 & ~w2911;
assign w2913 = ~w2728 & w2911;
assign v1382 = ~(w2912 | w2913);
assign w2914 = v1382;
assign w2915 = w2906 & ~w2914;
assign w2916 = ~w2906 & w2914;
assign v1383 = ~(w2915 | w2916);
assign w2917 = v1383;
assign w2918 = ~w2892 & w2917;
assign w2919 = w2892 & ~w2917;
assign v1384 = ~(w2918 | w2919);
assign w2920 = v1384;
assign w2921 = w2891 & w2920;
assign v1385 = ~(w2891 | w2920);
assign w2922 = v1385;
assign v1386 = ~(w2921 | w2922);
assign w2923 = v1386;
assign w2924 = w2874 & w2923;
assign v1387 = ~(w2874 | w2923);
assign w2925 = v1387;
assign v1388 = ~(w2924 | w2925);
assign w2926 = v1388;
assign v1389 = ~(w2734 | w2738);
assign w2927 = v1389;
assign v1390 = ~(w2737 | w2927);
assign w2928 = v1390;
assign w2929 = w2725 & ~w2727;
assign v1391 = ~(w2729 | w2929);
assign w2930 = v1391;
assign w2931 = w2928 & ~w2930;
assign w2932 = ~w2928 & w2930;
assign v1392 = ~(w2931 | w2932);
assign w2933 = v1392;
assign v1393 = ~(w2767 | w2771);
assign w2934 = v1393;
assign v1394 = ~(w2770 | w2934);
assign w2935 = v1394;
assign v1395 = ~(w2933 | w2935);
assign w2936 = v1395;
assign w2937 = w2933 & w2935;
assign v1396 = ~(w2936 | w2937);
assign w2938 = v1396;
assign v1397 = ~(w2715 | w2719);
assign w2939 = v1397;
assign w2940 = ~w2938 & w2939;
assign w2941 = w2938 & ~w2939;
assign v1398 = ~(w2940 | w2941);
assign w2942 = v1398;
assign w2943 = pi05 & pi33;
assign w2944 = pi06 & pi32;
assign w2945 = pi10 & pi28;
assign v1399 = ~(w2944 | w2945);
assign w2946 = v1399;
assign w2947 = w2944 & w2945;
assign v1400 = ~(w2946 | w2947);
assign w2948 = v1400;
assign w2949 = w2943 & ~w2948;
assign w2950 = ~w2943 & w2948;
assign v1401 = ~(w2949 | w2950);
assign w2951 = v1401;
assign w2952 = pi15 & pi23;
assign w2953 = pi16 & pi22;
assign w2954 = pi17 & pi21;
assign v1402 = ~(w2953 | w2954);
assign w2955 = v1402;
assign w2956 = w2953 & w2954;
assign v1403 = ~(w2955 | w2956);
assign w2957 = v1403;
assign w2958 = w2952 & ~w2957;
assign w2959 = ~w2952 & w2957;
assign v1404 = ~(w2958 | w2959);
assign w2960 = v1404;
assign v1405 = ~(w2951 | w2960);
assign w2961 = v1405;
assign w2962 = w2951 & w2960;
assign v1406 = ~(w2961 | w2962);
assign w2963 = v1406;
assign w2964 = pi09 & pi29;
assign w2965 = pi07 & pi31;
assign w2966 = pi08 & pi30;
assign v1407 = ~(w2965 | w2966);
assign w2967 = v1407;
assign w2968 = w2965 & w2966;
assign v1408 = ~(w2967 | w2968);
assign w2969 = v1408;
assign w2970 = w2964 & ~w2969;
assign w2971 = ~w2964 & w2969;
assign v1409 = ~(w2970 | w2971);
assign w2972 = v1409;
assign w2973 = w2963 & ~w2972;
assign w2974 = ~w2963 & w2972;
assign v1410 = ~(w2973 | w2974);
assign w2975 = v1410;
assign w2976 = w2942 & w2975;
assign v1411 = ~(w2942 | w2975);
assign w2977 = v1411;
assign v1412 = ~(w2976 | w2977);
assign w2978 = v1412;
assign w2979 = (~w2723 & ~w2724) | (~w2723 & w17072) | (~w2724 & w17072);
assign v1413 = ~(w2793 | w2795);
assign w2980 = v1413;
assign v1414 = ~(w2979 | w2980);
assign w2981 = v1414;
assign w2982 = w2979 & w2980;
assign v1415 = ~(w2981 | w2982);
assign w2983 = v1415;
assign w2984 = w2978 & w2983;
assign v1416 = ~(w2978 | w2983);
assign w2985 = v1416;
assign v1417 = ~(w2984 | w2985);
assign w2986 = v1417;
assign v1418 = ~(w2798 | w2801);
assign w2987 = v1418;
assign w2988 = w2986 & ~w2987;
assign w2989 = ~w2986 & w2987;
assign v1419 = ~(w2988 | w2989);
assign w2990 = v1419;
assign v1420 = ~(w2926 | w2990);
assign w2991 = v1420;
assign w2992 = w2926 & w2990;
assign v1421 = ~(w2991 | w2992);
assign w2993 = v1421;
assign w2994 = ~w2847 & w2993;
assign w2995 = w2847 & ~w2993;
assign v1422 = ~(w2994 | w2995);
assign w2996 = v1422;
assign v1423 = ~(w2687 | w2840);
assign w2997 = v1423;
assign w2998 = (w2997 & w2691) | (w2997 & w16512) | (w2691 & w16512);
assign v1424 = ~(w2839 | w2998);
assign w2999 = v1424;
assign w3000 = w2996 & w2999;
assign v1425 = ~(w2996 | w2999);
assign w3001 = v1425;
assign v1426 = ~(w3000 | w3001);
assign w3002 = v1426;
assign v1427 = ~(w2988 | w2992);
assign w3003 = v1427;
assign v1428 = ~(w2872 | w2924);
assign w3004 = v1428;
assign v1429 = ~(w2918 | w2921);
assign w3005 = v1429;
assign v1430 = ~(w2931 | w2937);
assign w3006 = v1430;
assign w3007 = (~w2856 & ~w2858) | (~w2856 & w16857) | (~w2858 & w16857);
assign w3008 = pi38 & w878;
assign w3009 = pi01 & pi38;
assign v1431 = ~(pi20 | w3009);
assign w3010 = v1431;
assign v1432 = ~(w3008 | w3010);
assign w3011 = v1432;
assign w3012 = pi00 & pi39;
assign w3013 = w2852 & w3012;
assign v1433 = ~(w2852 | w3012);
assign w3014 = v1433;
assign v1434 = ~(w3013 | w3014);
assign w3015 = v1434;
assign w3016 = w3011 & w3015;
assign v1435 = ~(w3011 | w3015);
assign w3017 = v1435;
assign v1436 = ~(w3016 | w3017);
assign w3018 = v1436;
assign w3019 = ~w3007 & w3018;
assign w3020 = w3007 & ~w3018;
assign v1437 = ~(w3019 | w3020);
assign w3021 = v1437;
assign w3022 = w3006 & ~w3021;
assign w3023 = ~w3006 & w3021;
assign v1438 = ~(w3022 | w3023);
assign w3024 = v1438;
assign v1439 = ~(w2728 | w2910);
assign w3025 = v1439;
assign v1440 = ~(w2909 | w3025);
assign w3026 = v1440;
assign v1441 = ~(w2810 | w2899);
assign w3027 = v1441;
assign v1442 = ~(w2897 | w3027);
assign w3028 = v1442;
assign w3029 = w3026 & w3028;
assign v1443 = ~(w3026 | w3028);
assign w3030 = v1443;
assign v1444 = ~(w3029 | w3030);
assign w3031 = v1444;
assign v1445 = ~(w2952 | w2956);
assign w3032 = v1445;
assign v1446 = ~(w2955 | w3032);
assign w3033 = v1446;
assign v1447 = ~(w3031 | w3033);
assign w3034 = v1447;
assign w3035 = w3031 & w3033;
assign v1448 = ~(w3034 | w3035);
assign w3036 = v1448;
assign w3037 = (~w2961 & ~w2963) | (~w2961 & w16858) | (~w2963 & w16858);
assign w3038 = (~w2904 & ~w2906) | (~w2904 & w16859) | (~w2906 & w16859);
assign v1449 = ~(w3037 | w3038);
assign w3039 = v1449;
assign w3040 = w3037 & w3038;
assign v1450 = ~(w3039 | w3040);
assign w3041 = v1450;
assign w3042 = w3036 & w3041;
assign v1451 = ~(w3036 | w3041);
assign w3043 = v1451;
assign v1452 = ~(w3042 | w3043);
assign w3044 = v1452;
assign w3045 = w3024 & w3044;
assign v1453 = ~(w3024 | w3044);
assign w3046 = v1453;
assign v1454 = ~(w3045 | w3046);
assign w3047 = v1454;
assign w3048 = ~w3005 & w3047;
assign w3049 = w3005 & ~w3047;
assign v1455 = ~(w3048 | w3049);
assign w3050 = v1455;
assign w3051 = ~w3004 & w3050;
assign w3052 = w3004 & ~w3050;
assign v1456 = ~(w3051 | w3052);
assign w3053 = v1456;
assign v1457 = ~(w2981 | w2984);
assign w3054 = v1457;
assign v1458 = ~(w2877 | w2881);
assign w3055 = v1458;
assign v1459 = ~(w2880 | w3055);
assign w3056 = v1459;
assign v1460 = ~(w2964 | w2968);
assign w3057 = v1460;
assign v1461 = ~(w2967 | w3057);
assign w3058 = v1461;
assign w3059 = w3056 & w3058;
assign v1462 = ~(w3056 | w3058);
assign w3060 = v1462;
assign v1463 = ~(w3059 | w3060);
assign w3061 = v1463;
assign v1464 = ~(w2943 | w2947);
assign w3062 = v1464;
assign v1465 = ~(w2946 | w3062);
assign w3063 = v1465;
assign v1466 = ~(w3061 | w3063);
assign w3064 = v1466;
assign w3065 = w3061 & w3063;
assign v1467 = ~(w3064 | w3065);
assign w3066 = v1467;
assign w3067 = (~w2886 & ~w2888) | (~w2886 & w17073) | (~w2888 & w17073);
assign w3068 = ~w3066 & w3067;
assign w3069 = w3066 & ~w3067;
assign v1468 = ~(w3068 | w3069);
assign w3070 = v1468;
assign w3071 = pi17 & pi22;
assign w3072 = pi04 & pi35;
assign w3073 = pi12 & pi27;
assign v1469 = ~(w3072 | w3073);
assign w3074 = v1469;
assign w3075 = w3072 & w3073;
assign v1470 = ~(w3074 | w3075);
assign w3076 = v1470;
assign w3077 = w3071 & ~w3076;
assign w3078 = ~w3071 & w3076;
assign v1471 = ~(w3077 | w3078);
assign w3079 = v1471;
assign w3080 = pi08 & pi31;
assign w3081 = pi19 & pi20;
assign w3082 = pi18 & pi21;
assign v1472 = ~(w3081 | w3082);
assign w3083 = v1472;
assign w3084 = w3081 & w3082;
assign v1473 = ~(w3083 | w3084);
assign w3085 = v1473;
assign w3086 = w3080 & ~w3085;
assign w3087 = ~w3080 & w3085;
assign v1474 = ~(w3086 | w3087);
assign w3088 = v1474;
assign v1475 = ~(w3079 | w3088);
assign w3089 = v1475;
assign w3090 = w3079 & w3088;
assign v1476 = ~(w3089 | w3090);
assign w3091 = v1476;
assign w3092 = pi11 & pi28;
assign w3093 = pi10 & pi29;
assign w3094 = pi05 & pi34;
assign v1477 = ~(w3093 | w3094);
assign w3095 = v1477;
assign w3096 = w3093 & w3094;
assign v1478 = ~(w3095 | w3096);
assign w3097 = v1478;
assign w3098 = w3092 & ~w3097;
assign w3099 = ~w3092 & w3097;
assign v1479 = ~(w3098 | w3099);
assign w3100 = v1479;
assign w3101 = w3091 & ~w3100;
assign w3102 = ~w3091 & w3100;
assign v1480 = ~(w3101 | w3102);
assign w3103 = v1480;
assign w3104 = w3070 & w3103;
assign v1481 = ~(w3070 | w3103);
assign w3105 = v1481;
assign v1482 = ~(w3104 | w3105);
assign w3106 = v1482;
assign w3107 = ~w3054 & w3106;
assign w3108 = w3054 & ~w3106;
assign v1483 = ~(w3107 | w3108);
assign w3109 = v1483;
assign v1484 = ~(w2941 | w2976);
assign w3110 = v1484;
assign v1485 = ~(w2866 | w2869);
assign w3111 = v1485;
assign w3112 = pi02 & pi37;
assign w3113 = pi03 & pi36;
assign w3114 = pi13 & pi26;
assign v1486 = ~(w3113 | w3114);
assign w3115 = v1486;
assign w3116 = w3113 & w3114;
assign v1487 = ~(w3115 | w3116);
assign w3117 = v1487;
assign w3118 = w3112 & ~w3117;
assign w3119 = ~w3112 & w3117;
assign v1488 = ~(w3118 | w3119);
assign w3120 = v1488;
assign w3121 = pi14 & pi25;
assign w3122 = pi15 & pi24;
assign w3123 = pi16 & pi23;
assign v1489 = ~(w3122 | w3123);
assign w3124 = v1489;
assign w3125 = w3122 & w3123;
assign v1490 = ~(w3124 | w3125);
assign w3126 = v1490;
assign w3127 = w3121 & ~w3126;
assign w3128 = ~w3121 & w3126;
assign v1491 = ~(w3127 | w3128);
assign w3129 = v1491;
assign v1492 = ~(w3120 | w3129);
assign w3130 = v1492;
assign w3131 = w3120 & w3129;
assign v1493 = ~(w3130 | w3131);
assign w3132 = v1493;
assign w3133 = pi06 & pi33;
assign w3134 = pi09 & pi30;
assign w3135 = pi07 & pi32;
assign v1494 = ~(w3134 | w3135);
assign w3136 = v1494;
assign w3137 = w3134 & w3135;
assign v1495 = ~(w3136 | w3137);
assign w3138 = v1495;
assign w3139 = w3133 & ~w3138;
assign w3140 = ~w3133 & w3138;
assign v1496 = ~(w3139 | w3140);
assign w3141 = v1496;
assign w3142 = w3132 & ~w3141;
assign w3143 = ~w3132 & w3141;
assign v1497 = ~(w3142 | w3143);
assign w3144 = v1497;
assign w3145 = ~w3111 & w3144;
assign w3146 = w3111 & ~w3144;
assign v1498 = ~(w3145 | w3146);
assign w3147 = v1498;
assign w3148 = ~w3110 & w3147;
assign w3149 = w3110 & ~w3147;
assign v1499 = ~(w3148 | w3149);
assign w3150 = v1499;
assign w3151 = w3109 & w3150;
assign v1500 = ~(w3109 | w3150);
assign w3152 = v1500;
assign v1501 = ~(w3151 | w3152);
assign w3153 = v1501;
assign w3154 = w3053 & w3153;
assign v1502 = ~(w3053 | w3153);
assign w3155 = v1502;
assign v1503 = ~(w3154 | w3155);
assign w3156 = v1503;
assign w3157 = ~w3003 & w3156;
assign w3158 = w3003 & ~w3156;
assign v1504 = ~(w3157 | w3158);
assign w3159 = v1504;
assign v1505 = ~(w2839 | w2994);
assign w3160 = v1505;
assign w3161 = (w2691 & w16514) | (w2691 & w16515) | (w16514 & w16515);
assign w3162 = w3159 & w3161;
assign v1506 = ~(w3159 | w3161);
assign w3163 = v1506;
assign v1507 = ~(w3162 | w3163);
assign w3164 = v1507;
assign v1508 = ~(w3051 | w3154);
assign w3165 = v1508;
assign w3166 = (~w3013 & ~w3015) | (~w3013 & w16722) | (~w3015 & w16722);
assign v1509 = ~(w3121 | w3125);
assign w3167 = v1509;
assign v1510 = ~(w3124 | w3167);
assign w3168 = v1510;
assign v1511 = ~(w3133 | w3137);
assign w3169 = v1511;
assign v1512 = ~(w3136 | w3169);
assign w3170 = v1512;
assign w3171 = w3168 & w3170;
assign v1513 = ~(w3168 | w3170);
assign w3172 = v1513;
assign v1514 = ~(w3171 | w3172);
assign w3173 = v1514;
assign w3174 = w3166 & ~w3173;
assign w3175 = ~w3166 & w3173;
assign v1515 = ~(w3174 | w3175);
assign w3176 = v1515;
assign w3177 = (~w3019 & ~w3021) | (~w3019 & w17074) | (~w3021 & w17074);
assign w3178 = ~w3176 & w3177;
assign w3179 = w3176 & ~w3177;
assign v1516 = ~(w3178 | w3179);
assign w3180 = v1516;
assign w3181 = pi18 & pi22;
assign w3182 = pi00 & pi40;
assign v1517 = ~(w2898 | w3182);
assign w3183 = v1517;
assign w3184 = pi02 & pi40;
assign w3185 = w2895 & w3184;
assign v1518 = ~(w3183 | w3185);
assign w3186 = v1518;
assign w3187 = w3181 & ~w3186;
assign w3188 = ~w3181 & w3186;
assign v1519 = ~(w3187 | w3188);
assign w3189 = v1519;
assign w3190 = pi07 & pi33;
assign w3191 = pi09 & pi31;
assign w3192 = pi08 & pi32;
assign v1520 = ~(w3191 | w3192);
assign w3193 = v1520;
assign w3194 = w3191 & w3192;
assign v1521 = ~(w3193 | w3194);
assign w3195 = v1521;
assign w3196 = w3190 & ~w3195;
assign w3197 = ~w3190 & w3195;
assign v1522 = ~(w3196 | w3197);
assign w3198 = v1522;
assign v1523 = ~(w3189 | w3198);
assign w3199 = v1523;
assign w3200 = w3189 & w3198;
assign v1524 = ~(w3199 | w3200);
assign w3201 = v1524;
assign w3202 = pi04 & pi36;
assign w3203 = pi12 & pi28;
assign w3204 = pi05 & pi35;
assign v1525 = ~(w3203 | w3204);
assign w3205 = v1525;
assign w3206 = w3203 & w3204;
assign v1526 = ~(w3205 | w3206);
assign w3207 = v1526;
assign w3208 = w3202 & ~w3207;
assign w3209 = ~w3202 & w3207;
assign v1527 = ~(w3208 | w3209);
assign w3210 = v1527;
assign w3211 = w3201 & ~w3210;
assign w3212 = ~w3201 & w3210;
assign v1528 = ~(w3211 | w3212);
assign w3213 = v1528;
assign v1529 = ~(w3180 | w3213);
assign w3214 = v1529;
assign w3215 = w3180 & w3213;
assign v1530 = ~(w3214 | w3215);
assign w3216 = v1530;
assign v1531 = ~(w3045 | w3048);
assign w3217 = v1531;
assign w3218 = ~w3216 & w3217;
assign w3219 = w3216 & ~w3217;
assign v1532 = ~(w3218 | w3219);
assign w3220 = v1532;
assign w3221 = pi19 & pi21;
assign w3222 = pi01 & pi39;
assign v1533 = ~(w3221 | w3222);
assign w3223 = v1533;
assign w3224 = w3221 & w3222;
assign v1534 = ~(w3223 | w3224);
assign w3225 = v1534;
assign w3226 = w3008 & w3225;
assign v1535 = ~(w3008 | w3225);
assign w3227 = v1535;
assign v1536 = ~(w3226 | w3227);
assign w3228 = v1536;
assign v1537 = ~(w3080 | w3084);
assign w3229 = v1537;
assign v1538 = ~(w3083 | w3229);
assign w3230 = v1538;
assign w3231 = w3228 & w3230;
assign v1539 = ~(w3228 | w3230);
assign w3232 = v1539;
assign v1540 = ~(w3231 | w3232);
assign w3233 = v1540;
assign w3234 = (~w3059 & ~w3061) | (~w3059 & w16860) | (~w3061 & w16860);
assign w3235 = (~w3029 & ~w3031) | (~w3029 & w16861) | (~w3031 & w16861);
assign v1541 = ~(w3234 | w3235);
assign w3236 = v1541;
assign w3237 = w3234 & w3235;
assign v1542 = ~(w3236 | w3237);
assign w3238 = v1542;
assign w3239 = w3233 & w3238;
assign v1543 = ~(w3233 | w3238);
assign w3240 = v1543;
assign v1544 = ~(w3239 | w3240);
assign w3241 = v1544;
assign w3242 = (~w3039 & ~w3041) | (~w3039 & w17075) | (~w3041 & w17075);
assign w3243 = pi03 & pi37;
assign w3244 = pi13 & pi27;
assign w3245 = pi14 & pi26;
assign v1545 = ~(w3244 | w3245);
assign w3246 = v1545;
assign w3247 = w3244 & w3245;
assign v1546 = ~(w3246 | w3247);
assign w3248 = v1546;
assign w3249 = w3243 & ~w3248;
assign w3250 = ~w3243 & w3248;
assign v1547 = ~(w3249 | w3250);
assign w3251 = v1547;
assign w3252 = pi15 & pi25;
assign w3253 = pi16 & pi24;
assign w3254 = pi17 & pi23;
assign v1548 = ~(w3253 | w3254);
assign w3255 = v1548;
assign w3256 = w3253 & w3254;
assign v1549 = ~(w3255 | w3256);
assign w3257 = v1549;
assign w3258 = w3252 & ~w3257;
assign w3259 = ~w3252 & w3257;
assign v1550 = ~(w3258 | w3259);
assign w3260 = v1550;
assign v1551 = ~(w3251 | w3260);
assign w3261 = v1551;
assign w3262 = w3251 & w3260;
assign v1552 = ~(w3261 | w3262);
assign w3263 = v1552;
assign w3264 = pi11 & pi29;
assign w3265 = pi06 & pi34;
assign w3266 = pi10 & pi30;
assign v1553 = ~(w3265 | w3266);
assign w3267 = v1553;
assign w3268 = w3265 & w3266;
assign v1554 = ~(w3267 | w3268);
assign w3269 = v1554;
assign w3270 = w3264 & ~w3269;
assign w3271 = ~w3264 & w3269;
assign v1555 = ~(w3270 | w3271);
assign w3272 = v1555;
assign w3273 = w3263 & ~w3272;
assign w3274 = ~w3263 & w3272;
assign v1556 = ~(w3273 | w3274);
assign w3275 = v1556;
assign w3276 = ~w3242 & w3275;
assign w3277 = w3242 & ~w3275;
assign v1557 = ~(w3276 | w3277);
assign w3278 = v1557;
assign w3279 = w3241 & w3278;
assign v1558 = ~(w3241 | w3278);
assign w3280 = v1558;
assign v1559 = ~(w3279 | w3280);
assign w3281 = v1559;
assign w3282 = w3220 & w3281;
assign v1560 = ~(w3220 | w3281);
assign w3283 = v1560;
assign v1561 = ~(w3282 | w3283);
assign w3284 = v1561;
assign v1562 = ~(w3145 | w3148);
assign w3285 = v1562;
assign v1563 = ~(w3069 | w3104);
assign w3286 = v1563;
assign v1564 = ~(w3092 | w3096);
assign w3287 = v1564;
assign v1565 = ~(w3095 | w3287);
assign w3288 = v1565;
assign v1566 = ~(w3112 | w3116);
assign w3289 = v1566;
assign v1567 = ~(w3115 | w3289);
assign w3290 = v1567;
assign w3291 = w3288 & w3290;
assign v1568 = ~(w3288 | w3290);
assign w3292 = v1568;
assign v1569 = ~(w3291 | w3292);
assign w3293 = v1569;
assign v1570 = ~(w3071 | w3075);
assign w3294 = v1570;
assign v1571 = ~(w3074 | w3294);
assign w3295 = v1571;
assign v1572 = ~(w3293 | w3295);
assign w3296 = v1572;
assign w3297 = w3293 & w3295;
assign v1573 = ~(w3296 | w3297);
assign w3298 = v1573;
assign w3299 = (~w3089 & ~w3091) | (~w3089 & w16862) | (~w3091 & w16862);
assign w3300 = (~w3130 & ~w3132) | (~w3130 & w16863) | (~w3132 & w16863);
assign v1574 = ~(w3299 | w3300);
assign w3301 = v1574;
assign w3302 = w3299 & w3300;
assign v1575 = ~(w3301 | w3302);
assign w3303 = v1575;
assign w3304 = w3298 & w3303;
assign v1576 = ~(w3298 | w3303);
assign w3305 = v1576;
assign v1577 = ~(w3304 | w3305);
assign w3306 = v1577;
assign w3307 = ~w3286 & w3306;
assign w3308 = w3286 & ~w3306;
assign v1578 = ~(w3307 | w3308);
assign w3309 = v1578;
assign w3310 = ~w3285 & w3309;
assign w3311 = w3285 & ~w3309;
assign v1579 = ~(w3310 | w3311);
assign w3312 = v1579;
assign v1580 = ~(w3107 | w3151);
assign w3313 = v1580;
assign w3314 = w3312 & ~w3313;
assign w3315 = ~w3312 & w3313;
assign v1581 = ~(w3314 | w3315);
assign w3316 = v1581;
assign w3317 = w3284 & w3316;
assign v1582 = ~(w3284 | w3316);
assign w3318 = v1582;
assign v1583 = ~(w3317 | w3318);
assign w3319 = v1583;
assign w3320 = ~w3165 & w3319;
assign w3321 = w3165 & ~w3319;
assign v1584 = ~(w3320 | w3321);
assign w3322 = v1584;
assign v1585 = ~(w3157 | w3161);
assign w3323 = v1585;
assign v1586 = ~(w3158 | w3323);
assign w3324 = v1586;
assign w3325 = w3322 & w3324;
assign v1587 = ~(w3322 | w3324);
assign w3326 = v1587;
assign v1588 = ~(w3325 | w3326);
assign w3327 = v1588;
assign v1589 = ~(w3314 | w3317);
assign w3328 = v1589;
assign v1590 = ~(w3276 | w3279);
assign w3329 = v1590;
assign v1591 = ~(w3179 | w3215);
assign w3330 = v1591;
assign v1592 = ~(w3252 | w3256);
assign w3331 = v1592;
assign v1593 = ~(w3255 | w3331);
assign w3332 = v1593;
assign w3333 = w3181 & ~w3183;
assign v1594 = ~(w3185 | w3333);
assign w3334 = v1594;
assign w3335 = w3332 & ~w3334;
assign w3336 = ~w3332 & w3334;
assign v1595 = ~(w3335 | w3336);
assign w3337 = v1595;
assign v1596 = ~(w3243 | w3247);
assign w3338 = v1596;
assign v1597 = ~(w3246 | w3338);
assign w3339 = v1597;
assign v1598 = ~(w3337 | w3339);
assign w3340 = v1598;
assign w3341 = w3337 & w3339;
assign v1599 = ~(w3340 | w3341);
assign w3342 = v1599;
assign w3343 = (~w3199 & ~w3201) | (~w3199 & w16864) | (~w3201 & w16864);
assign w3344 = ~w3342 & w3343;
assign w3345 = w3342 & ~w3343;
assign v1600 = ~(w3344 | w3345);
assign w3346 = v1600;
assign w3347 = pi40 & w964;
assign w3348 = pi01 & pi40;
assign v1601 = ~(pi21 | w3348);
assign w3349 = v1601;
assign v1602 = ~(w3347 | w3349);
assign w3350 = v1602;
assign v1603 = ~(w3190 | w3194);
assign w3351 = v1603;
assign v1604 = ~(w3193 | w3351);
assign w3352 = v1604;
assign w3353 = w3350 & w3352;
assign v1605 = ~(w3350 | w3352);
assign w3354 = v1605;
assign v1606 = ~(w3353 | w3354);
assign w3355 = v1606;
assign v1607 = ~(w3264 | w3268);
assign w3356 = v1607;
assign v1608 = ~(w3267 | w3356);
assign w3357 = v1608;
assign w3358 = w3355 & w3357;
assign v1609 = ~(w3355 | w3357);
assign w3359 = v1609;
assign v1610 = ~(w3358 | w3359);
assign w3360 = v1610;
assign w3361 = w3346 & w3360;
assign v1611 = ~(w3346 | w3360);
assign w3362 = v1611;
assign v1612 = ~(w3361 | w3362);
assign w3363 = v1612;
assign w3364 = ~w3330 & w3363;
assign w3365 = w3330 & ~w3363;
assign v1613 = ~(w3364 | w3365);
assign w3366 = v1613;
assign w3367 = w3329 & ~w3366;
assign w3368 = ~w3329 & w3366;
assign v1614 = ~(w3367 | w3368);
assign w3369 = v1614;
assign v1615 = ~(w3219 | w3282);
assign w3370 = v1615;
assign w3371 = ~w3369 & w3370;
assign w3372 = w3369 & ~w3370;
assign v1616 = ~(w3371 | w3372);
assign w3373 = v1616;
assign w3374 = (~w3261 & ~w3263) | (~w3261 & w16865) | (~w3263 & w16865);
assign w3375 = (~w3171 & ~w3173) | (~w3171 & w16723) | (~w3173 & w16723);
assign w3376 = (~w3291 & ~w3293) | (~w3291 & w16724) | (~w3293 & w16724);
assign v1617 = ~(w3375 | w3376);
assign w3377 = v1617;
assign w3378 = w3375 & w3376;
assign v1618 = ~(w3377 | w3378);
assign w3379 = v1618;
assign w3380 = w3374 & ~w3379;
assign w3381 = ~w3374 & w3379;
assign v1619 = ~(w3380 | w3381);
assign w3382 = v1619;
assign v1620 = ~(w3202 | w3206);
assign w3383 = v1620;
assign v1621 = ~(w3205 | w3383);
assign w3384 = v1621;
assign w3385 = pi00 & pi41;
assign w3386 = pi02 & pi39;
assign v1622 = ~(w3385 | w3386);
assign w3387 = v1622;
assign w3388 = pi02 & pi41;
assign w3389 = w3012 & w3388;
assign v1623 = ~(w3387 | w3389);
assign w3390 = v1623;
assign w3391 = w3224 & ~w3390;
assign w3392 = ~w3224 & w3390;
assign v1624 = ~(w3391 | w3392);
assign w3393 = v1624;
assign w3394 = w3384 & ~w3393;
assign w3395 = ~w3384 & w3393;
assign v1625 = ~(w3394 | w3395);
assign w3396 = v1625;
assign w3397 = pi03 & pi38;
assign w3398 = pi13 & pi28;
assign w3399 = pi15 & pi26;
assign v1626 = ~(w3398 | w3399);
assign w3400 = v1626;
assign w3401 = w3398 & w3399;
assign v1627 = ~(w3400 | w3401);
assign w3402 = v1627;
assign w3403 = w3397 & ~w3402;
assign w3404 = ~w3397 & w3402;
assign v1628 = ~(w3403 | w3404);
assign w3405 = v1628;
assign w3406 = ~w3396 & w3405;
assign w3407 = w3396 & ~w3405;
assign v1629 = ~(w3406 | w3407);
assign w3408 = v1629;
assign w3409 = (~w3301 & ~w3303) | (~w3301 & w17076) | (~w3303 & w17076);
assign w3410 = w3408 & ~w3409;
assign w3411 = ~w3408 & w3409;
assign v1630 = ~(w3410 | w3411);
assign w3412 = v1630;
assign v1631 = ~(w3382 | w3412);
assign w3413 = v1631;
assign w3414 = w3382 & w3412;
assign v1632 = ~(w3413 | w3414);
assign w3415 = v1632;
assign w3416 = (~w3307 & w3285) | (~w3307 & w16725) | (w3285 & w16725);
assign w3417 = (~w3226 & ~w3228) | (~w3226 & w17077) | (~w3228 & w17077);
assign w3418 = pi08 & pi33;
assign w3419 = pi20 & pi21;
assign w3420 = pi19 & pi22;
assign v1633 = ~(w3419 | w3420);
assign w3421 = v1633;
assign w3422 = w3419 & w3420;
assign v1634 = ~(w3421 | w3422);
assign w3423 = v1634;
assign w3424 = w3418 & ~w3423;
assign w3425 = ~w3418 & w3423;
assign v1635 = ~(w3424 | w3425);
assign w3426 = v1635;
assign w3427 = pi05 & pi36;
assign w3428 = pi06 & pi35;
assign w3429 = pi11 & pi30;
assign v1636 = ~(w3428 | w3429);
assign w3430 = v1636;
assign w3431 = w3428 & w3429;
assign v1637 = ~(w3430 | w3431);
assign w3432 = v1637;
assign w3433 = w3427 & ~w3432;
assign w3434 = ~w3427 & w3432;
assign v1638 = ~(w3433 | w3434);
assign w3435 = v1638;
assign v1639 = ~(w3426 | w3435);
assign w3436 = v1639;
assign w3437 = w3426 & w3435;
assign v1640 = ~(w3436 | w3437);
assign w3438 = v1640;
assign w3439 = w3417 & ~w3438;
assign w3440 = ~w3417 & w3438;
assign v1641 = ~(w3439 | w3440);
assign w3441 = v1641;
assign w3442 = (~w3236 & ~w3238) | (~w3236 & w16726) | (~w3238 & w16726);
assign w3443 = ~w3441 & w3442;
assign w3444 = w3441 & ~w3442;
assign v1642 = ~(w3443 | w3444);
assign w3445 = v1642;
assign w3446 = pi14 & pi27;
assign w3447 = pi04 & pi37;
assign w3448 = pi12 & pi29;
assign v1643 = ~(w3447 | w3448);
assign w3449 = v1643;
assign w3450 = w3447 & w3448;
assign v1644 = ~(w3449 | w3450);
assign w3451 = v1644;
assign w3452 = w3446 & ~w3451;
assign w3453 = ~w3446 & w3451;
assign v1645 = ~(w3452 | w3453);
assign w3454 = v1645;
assign w3455 = pi16 & pi25;
assign w3456 = pi17 & pi24;
assign w3457 = pi18 & pi23;
assign v1646 = ~(w3456 | w3457);
assign w3458 = v1646;
assign w3459 = w3456 & w3457;
assign v1647 = ~(w3458 | w3459);
assign w3460 = v1647;
assign w3461 = w3455 & ~w3460;
assign w3462 = ~w3455 & w3460;
assign v1648 = ~(w3461 | w3462);
assign w3463 = v1648;
assign v1649 = ~(w3454 | w3463);
assign w3464 = v1649;
assign w3465 = w3454 & w3463;
assign v1650 = ~(w3464 | w3465);
assign w3466 = v1650;
assign w3467 = pi10 & pi31;
assign w3468 = pi09 & pi32;
assign w3469 = pi07 & pi34;
assign v1651 = ~(w3468 | w3469);
assign w3470 = v1651;
assign w3471 = w3468 & w3469;
assign v1652 = ~(w3470 | w3471);
assign w3472 = v1652;
assign w3473 = w3467 & ~w3472;
assign w3474 = ~w3467 & w3472;
assign v1653 = ~(w3473 | w3474);
assign w3475 = v1653;
assign w3476 = w3466 & ~w3475;
assign w3477 = ~w3466 & w3475;
assign v1654 = ~(w3476 | w3477);
assign w3478 = v1654;
assign v1655 = ~(w3445 | w3478);
assign w3479 = v1655;
assign w3480 = w3445 & w3478;
assign v1656 = ~(w3479 | w3480);
assign w3481 = v1656;
assign w3482 = ~w3416 & w3481;
assign w3483 = w3416 & ~w3481;
assign v1657 = ~(w3482 | w3483);
assign w3484 = v1657;
assign w3485 = w3415 & w3484;
assign v1658 = ~(w3415 | w3484);
assign w3486 = v1658;
assign v1659 = ~(w3485 | w3486);
assign w3487 = v1659;
assign w3488 = w3373 & w3487;
assign v1660 = ~(w3373 | w3487);
assign w3489 = v1660;
assign v1661 = ~(w3488 | w3489);
assign w3490 = v1661;
assign w3491 = w3328 & ~w3490;
assign w3492 = ~w3328 & w3490;
assign v1662 = ~(w3491 | w3492);
assign w3493 = v1662;
assign v1663 = ~(w3158 | w3321);
assign w3494 = v1663;
assign w3495 = (w3494 & w3161) | (w3494 & w16516) | (w3161 & w16516);
assign v1664 = ~(w3320 | w3495);
assign w3496 = v1664;
assign w3497 = w3493 & w3496;
assign v1665 = ~(w3493 | w3496);
assign w3498 = v1665;
assign v1666 = ~(w3497 | w3498);
assign w3499 = v1666;
assign v1667 = ~(w3320 | w3492);
assign w3500 = v1667;
assign w3501 = (~w3491 & w3495) | (~w3491 & w16517) | (w3495 & w16517);
assign v1668 = ~(w3372 | w3488);
assign w3502 = v1668;
assign v1669 = ~(w3482 | w3485);
assign w3503 = v1669;
assign v1670 = ~(w3410 | w3414);
assign w3504 = v1670;
assign v1671 = ~(w3464 | w3476);
assign w3505 = v1671;
assign v1672 = ~(w3335 | w3341);
assign w3506 = v1672;
assign w3507 = (~w3394 & ~w3396) | (~w3394 & w17078) | (~w3396 & w17078);
assign v1673 = ~(w3506 | w3507);
assign w3508 = v1673;
assign w3509 = w3506 & w3507;
assign v1674 = ~(w3508 | w3509);
assign w3510 = v1674;
assign w3511 = w3505 & ~w3510;
assign w3512 = ~w3505 & w3510;
assign v1675 = ~(w3511 | w3512);
assign w3513 = v1675;
assign w3514 = (~w3444 & ~w3445) | (~w3444 & w17079) | (~w3445 & w17079);
assign w3515 = ~w3513 & w3514;
assign w3516 = w3513 & ~w3514;
assign v1676 = ~(w3515 | w3516);
assign w3517 = v1676;
assign w3518 = ~w3504 & w3517;
assign w3519 = w3504 & ~w3517;
assign v1677 = ~(w3518 | w3519);
assign w3520 = v1677;
assign w3521 = ~w3503 & w3520;
assign w3522 = w3503 & ~w3520;
assign v1678 = ~(w3521 | w3522);
assign w3523 = v1678;
assign w3524 = (~w3364 & ~w3366) | (~w3364 & w16727) | (~w3366 & w16727);
assign v1679 = ~(w3467 | w3471);
assign w3525 = v1679;
assign v1680 = ~(w3470 | w3525);
assign w3526 = v1680;
assign w3527 = pi06 & pi36;
assign w3528 = pi07 & pi35;
assign w3529 = pi11 & pi31;
assign v1681 = ~(w3528 | w3529);
assign w3530 = v1681;
assign w3531 = w3528 & w3529;
assign v1682 = ~(w3530 | w3531);
assign w3532 = v1682;
assign w3533 = w3527 & ~w3532;
assign w3534 = ~w3527 & w3532;
assign v1683 = ~(w3533 | w3534);
assign w3535 = v1683;
assign w3536 = w3526 & ~w3535;
assign w3537 = ~w3526 & w3535;
assign v1684 = ~(w3536 | w3537);
assign w3538 = v1684;
assign w3539 = pi10 & pi32;
assign w3540 = pi09 & pi33;
assign w3541 = pi08 & pi34;
assign v1685 = ~(w3540 | w3541);
assign w3542 = v1685;
assign w3543 = w3540 & w3541;
assign v1686 = ~(w3542 | w3543);
assign w3544 = v1686;
assign w3545 = w3539 & ~w3544;
assign w3546 = ~w3539 & w3544;
assign v1687 = ~(w3545 | w3546);
assign w3547 = v1687;
assign w3548 = w3538 & ~w3547;
assign w3549 = ~w3538 & w3547;
assign v1688 = ~(w3548 | w3549);
assign w3550 = v1688;
assign w3551 = (w3550 & w3381) | (w3550 & w16728) | (w3381 & w16728);
assign w3552 = ~w3381 & w16729;
assign v1689 = ~(w3551 | w3552);
assign w3553 = v1689;
assign w3554 = pi03 & pi39;
assign w3555 = pi16 & pi26;
assign v1690 = ~(w3554 | w3555);
assign w3556 = v1690;
assign w3557 = w3554 & w3555;
assign v1691 = ~(w3556 | w3557);
assign w3558 = v1691;
assign w3559 = w3184 & ~w3558;
assign w3560 = ~w3184 & w3558;
assign v1692 = ~(w3559 | w3560);
assign w3561 = v1692;
assign w3562 = pi17 & pi25;
assign w3563 = pi18 & pi24;
assign w3564 = pi19 & pi23;
assign v1693 = ~(w3563 | w3564);
assign w3565 = v1693;
assign w3566 = w3563 & w3564;
assign v1694 = ~(w3565 | w3566);
assign w3567 = v1694;
assign w3568 = w3562 & ~w3567;
assign w3569 = ~w3562 & w3567;
assign v1695 = ~(w3568 | w3569);
assign w3570 = v1695;
assign v1696 = ~(w3561 | w3570);
assign w3571 = v1696;
assign w3572 = w3561 & w3570;
assign v1697 = ~(w3571 | w3572);
assign w3573 = v1697;
assign w3574 = pi15 & pi27;
assign w3575 = pi04 & pi38;
assign w3576 = pi14 & pi28;
assign v1698 = ~(w3575 | w3576);
assign w3577 = v1698;
assign w3578 = w3575 & w3576;
assign v1699 = ~(w3577 | w3578);
assign w3579 = v1699;
assign w3580 = w3574 & ~w3579;
assign w3581 = ~w3574 & w3579;
assign v1700 = ~(w3580 | w3581);
assign w3582 = v1700;
assign w3583 = w3573 & ~w3582;
assign w3584 = ~w3573 & w3582;
assign v1701 = ~(w3583 | w3584);
assign w3585 = v1701;
assign w3586 = w3553 & w3585;
assign v1702 = ~(w3553 | w3585);
assign w3587 = v1702;
assign v1703 = ~(w3586 | w3587);
assign w3588 = v1703;
assign w3589 = ~w3524 & w3588;
assign w3590 = w3524 & ~w3588;
assign v1704 = ~(w3589 | w3590);
assign w3591 = v1704;
assign w3592 = (~w3353 & ~w3355) | (~w3353 & w16866) | (~w3355 & w16866);
assign w3593 = pi00 & pi42;
assign w3594 = w3347 & w3593;
assign v1705 = ~(w3347 | w3593);
assign w3595 = v1705;
assign v1706 = ~(w3594 | w3595);
assign w3596 = v1706;
assign w3597 = pi20 & pi22;
assign w3598 = pi01 & pi41;
assign v1707 = ~(w3597 | w3598);
assign w3599 = v1707;
assign w3600 = w3597 & w3598;
assign v1708 = ~(w3599 | w3600);
assign w3601 = v1708;
assign w3602 = w3596 & w3601;
assign v1709 = ~(w3596 | w3601);
assign w3603 = v1709;
assign v1710 = ~(w3602 | w3603);
assign w3604 = v1710;
assign w3605 = pi13 & pi29;
assign w3606 = pi05 & pi37;
assign w3607 = pi12 & pi30;
assign v1711 = ~(w3606 | w3607);
assign w3608 = v1711;
assign w3609 = w3606 & w3607;
assign v1712 = ~(w3608 | w3609);
assign w3610 = v1712;
assign w3611 = w3605 & ~w3610;
assign w3612 = ~w3605 & w3610;
assign v1713 = ~(w3611 | w3612);
assign w3613 = v1713;
assign w3614 = w3604 & ~w3613;
assign w3615 = ~w3604 & w3613;
assign v1714 = ~(w3614 | w3615);
assign w3616 = v1714;
assign w3617 = w3592 & ~w3616;
assign w3618 = ~w3592 & w3616;
assign v1715 = ~(w3617 | w3618);
assign w3619 = v1715;
assign w3620 = (~w3345 & ~w3346) | (~w3345 & w16730) | (~w3346 & w16730);
assign w3621 = ~w3619 & w3620;
assign w3622 = w3619 & ~w3620;
assign v1716 = ~(w3621 | w3622);
assign w3623 = v1716;
assign v1717 = ~(w3446 | w3450);
assign w3624 = v1717;
assign v1718 = ~(w3449 | w3624);
assign w3625 = v1718;
assign v1719 = ~(w3418 | w3422);
assign w3626 = v1719;
assign v1720 = ~(w3421 | w3626);
assign w3627 = v1720;
assign w3628 = w3625 & w3627;
assign v1721 = ~(w3625 | w3627);
assign w3629 = v1721;
assign v1722 = ~(w3628 | w3629);
assign w3630 = v1722;
assign v1723 = ~(w3427 | w3431);
assign w3631 = v1723;
assign v1724 = ~(w3430 | w3631);
assign w3632 = v1724;
assign v1725 = ~(w3630 | w3632);
assign w3633 = v1725;
assign w3634 = w3630 & w3632;
assign v1726 = ~(w3633 | w3634);
assign w3635 = v1726;
assign w3636 = (~w3436 & ~w3438) | (~w3436 & w17080) | (~w3438 & w17080);
assign w3637 = ~w3635 & w3636;
assign w3638 = w3635 & ~w3636;
assign v1727 = ~(w3637 | w3638);
assign w3639 = v1727;
assign v1728 = ~(w3397 | w3401);
assign w3640 = v1728;
assign v1729 = ~(w3400 | w3640);
assign w3641 = v1729;
assign v1730 = ~(w3455 | w3459);
assign w3642 = v1730;
assign v1731 = ~(w3458 | w3642);
assign w3643 = v1731;
assign w3644 = w3641 & w3643;
assign v1732 = ~(w3641 | w3643);
assign w3645 = v1732;
assign v1733 = ~(w3644 | w3645);
assign w3646 = v1733;
assign w3647 = w3224 & ~w3387;
assign v1734 = ~(w3389 | w3647);
assign w3648 = v1734;
assign w3649 = ~w3646 & w3648;
assign w3650 = w3646 & ~w3648;
assign v1735 = ~(w3649 | w3650);
assign w3651 = v1735;
assign w3652 = w3639 & w3651;
assign v1736 = ~(w3639 | w3651);
assign w3653 = v1736;
assign v1737 = ~(w3652 | w3653);
assign w3654 = v1737;
assign w3655 = w3623 & w3654;
assign v1738 = ~(w3623 | w3654);
assign w3656 = v1738;
assign v1739 = ~(w3655 | w3656);
assign w3657 = v1739;
assign w3658 = w3591 & w3657;
assign v1740 = ~(w3591 | w3657);
assign w3659 = v1740;
assign v1741 = ~(w3658 | w3659);
assign w3660 = v1741;
assign v1742 = ~(w3523 | w3660);
assign w3661 = v1742;
assign w3662 = w3523 & w3660;
assign v1743 = ~(w3661 | w3662);
assign w3663 = v1743;
assign w3664 = w3502 & ~w3663;
assign w3665 = ~w3502 & w3663;
assign v1744 = ~(w3664 | w3665);
assign w3666 = v1744;
assign w3667 = w3501 & ~w3666;
assign w3668 = ~w3501 & w3666;
assign v1745 = ~(w3667 | w3668);
assign w3669 = v1745;
assign w3670 = (~w3495 & w16518) | (~w3495 & w16519) | (w16518 & w16519);
assign v1746 = ~(w3664 | w3670);
assign w3671 = v1746;
assign v1747 = ~(w3521 | w3662);
assign w3672 = v1747;
assign v1748 = ~(w3516 | w3518);
assign w3673 = v1748;
assign v1749 = ~(w3508 | w3512);
assign w3674 = v1749;
assign w3675 = pi04 & pi39;
assign w3676 = pi00 & pi43;
assign w3677 = pi03 & pi40;
assign v1750 = ~(w3676 | w3677);
assign w3678 = v1750;
assign w3679 = w3676 & w3677;
assign v1751 = ~(w3678 | w3679);
assign w3680 = v1751;
assign w3681 = w3675 & ~w3680;
assign w3682 = ~w3675 & w3680;
assign v1752 = ~(w3681 | w3682);
assign w3683 = v1752;
assign w3684 = pi15 & pi28;
assign w3685 = pi16 & pi27;
assign v1753 = ~(w3684 | w3685);
assign w3686 = v1753;
assign w3687 = w3684 & w3685;
assign v1754 = ~(w3686 | w3687);
assign w3688 = v1754;
assign w3689 = w1755 & ~w3688;
assign w3690 = ~w1755 & w3688;
assign v1755 = ~(w3689 | w3690);
assign w3691 = v1755;
assign v1756 = ~(w3683 | w3691);
assign w3692 = v1756;
assign w3693 = w3683 & w3691;
assign v1757 = ~(w3692 | w3693);
assign w3694 = v1757;
assign w3695 = pi17 & pi26;
assign w3696 = pi19 & pi24;
assign w3697 = pi18 & pi25;
assign v1758 = ~(w3696 | w3697);
assign w3698 = v1758;
assign w3699 = w3696 & w3697;
assign v1759 = ~(w3698 | w3699);
assign w3700 = v1759;
assign w3701 = w3695 & ~w3700;
assign w3702 = ~w3695 & w3700;
assign v1760 = ~(w3701 | w3702);
assign w3703 = v1760;
assign w3704 = w3694 & ~w3703;
assign w3705 = ~w3694 & w3703;
assign v1761 = ~(w3704 | w3705);
assign w3706 = v1761;
assign w3707 = pi09 & pi34;
assign w3708 = pi21 & pi22;
assign w3709 = pi20 & pi23;
assign v1762 = ~(w3708 | w3709);
assign w3710 = v1762;
assign w3711 = w3708 & w3709;
assign v1763 = ~(w3710 | w3711);
assign w3712 = v1763;
assign w3713 = w3707 & ~w3712;
assign w3714 = ~w3707 & w3712;
assign v1764 = ~(w3713 | w3714);
assign w3715 = v1764;
assign w3716 = pi07 & pi36;
assign w3717 = pi10 & pi33;
assign w3718 = pi08 & pi35;
assign v1765 = ~(w3717 | w3718);
assign w3719 = v1765;
assign w3720 = w3717 & w3718;
assign v1766 = ~(w3719 | w3720);
assign w3721 = v1766;
assign w3722 = w3716 & ~w3721;
assign w3723 = ~w3716 & w3721;
assign v1767 = ~(w3722 | w3723);
assign w3724 = v1767;
assign v1768 = ~(w3715 | w3724);
assign w3725 = v1768;
assign w3726 = w3715 & w3724;
assign v1769 = ~(w3725 | w3726);
assign w3727 = v1769;
assign w3728 = pi05 & pi38;
assign w3729 = pi13 & pi30;
assign v1770 = ~(w3728 | w3729);
assign w3730 = v1770;
assign w3731 = w3728 & w3729;
assign v1771 = ~(w3730 | w3731);
assign w3732 = v1771;
assign w3733 = w3388 & ~w3732;
assign w3734 = ~w3388 & w3732;
assign v1772 = ~(w3733 | w3734);
assign w3735 = v1772;
assign w3736 = w3727 & ~w3735;
assign w3737 = ~w3727 & w3735;
assign v1773 = ~(w3736 | w3737);
assign w3738 = v1773;
assign w3739 = w3706 & w3738;
assign v1774 = ~(w3706 | w3738);
assign w3740 = v1774;
assign v1775 = ~(w3739 | w3740);
assign w3741 = v1775;
assign w3742 = ~w3674 & w3741;
assign w3743 = w3674 & ~w3741;
assign v1776 = ~(w3742 | w3743);
assign w3744 = v1776;
assign w3745 = ~w3673 & w3744;
assign w3746 = w3673 & ~w3744;
assign v1777 = ~(w3745 | w3746);
assign w3747 = v1777;
assign w3748 = (~w3614 & ~w3616) | (~w3614 & w16867) | (~w3616 & w16867);
assign v1778 = ~(w3574 | w3578);
assign w3749 = v1778;
assign v1779 = ~(w3577 | w3749);
assign w3750 = v1779;
assign v1780 = ~(w3527 | w3531);
assign w3751 = v1780;
assign v1781 = ~(w3530 | w3751);
assign w3752 = v1781;
assign w3753 = w3750 & w3752;
assign v1782 = ~(w3750 | w3752);
assign w3754 = v1782;
assign v1783 = ~(w3753 | w3754);
assign w3755 = v1783;
assign v1784 = ~(w3562 | w3566);
assign w3756 = v1784;
assign v1785 = ~(w3565 | w3756);
assign w3757 = v1785;
assign v1786 = ~(w3755 | w3757);
assign w3758 = v1786;
assign w3759 = w3755 & w3757;
assign v1787 = ~(w3758 | w3759);
assign w3760 = v1787;
assign w3761 = (~w3594 & ~w3596) | (~w3594 & w16868) | (~w3596 & w16868);
assign v1788 = ~(w3184 | w3557);
assign w3762 = v1788;
assign v1789 = ~(w3556 | w3762);
assign w3763 = v1789;
assign v1790 = ~(w3605 | w3609);
assign w3764 = v1790;
assign v1791 = ~(w3608 | w3764);
assign w3765 = v1791;
assign w3766 = w3763 & w3765;
assign v1792 = ~(w3763 | w3765);
assign w3767 = v1792;
assign v1793 = ~(w3766 | w3767);
assign w3768 = v1793;
assign w3769 = w3761 & ~w3768;
assign w3770 = ~w3761 & w3768;
assign v1794 = ~(w3769 | w3770);
assign w3771 = v1794;
assign w3772 = w3760 & w3771;
assign v1795 = ~(w3760 | w3771);
assign w3773 = v1795;
assign v1796 = ~(w3772 | w3773);
assign w3774 = v1796;
assign w3775 = ~w3748 & w3774;
assign w3776 = w3748 & ~w3774;
assign v1797 = ~(w3775 | w3776);
assign w3777 = v1797;
assign w3778 = (~w3644 & ~w3646) | (~w3644 & w17081) | (~w3646 & w17081);
assign w3779 = (~w3628 & ~w3630) | (~w3628 & w16731) | (~w3630 & w16731);
assign w3780 = pi12 & pi31;
assign w3781 = pi11 & pi32;
assign w3782 = pi06 & pi37;
assign v1798 = ~(w3781 | w3782);
assign w3783 = v1798;
assign w3784 = w3781 & w3782;
assign v1799 = ~(w3783 | w3784);
assign w3785 = v1799;
assign w3786 = w3780 & ~w3785;
assign w3787 = ~w3780 & w3785;
assign v1800 = ~(w3786 | w3787);
assign w3788 = v1800;
assign v1801 = ~(w3779 | w3788);
assign w3789 = v1801;
assign w3790 = w3779 & w3788;
assign v1802 = ~(w3789 | w3790);
assign w3791 = v1802;
assign w3792 = w3778 & ~w3791;
assign w3793 = ~w3778 & w3791;
assign v1803 = ~(w3792 | w3793);
assign w3794 = v1803;
assign v1804 = ~(w3638 | w3652);
assign w3795 = v1804;
assign w3796 = ~w3794 & w3795;
assign w3797 = w3794 & ~w3795;
assign v1805 = ~(w3796 | w3797);
assign w3798 = v1805;
assign w3799 = w3777 & w3798;
assign v1806 = ~(w3777 | w3798);
assign w3800 = v1806;
assign v1807 = ~(w3799 | w3800);
assign w3801 = v1807;
assign w3802 = w3747 & w3801;
assign v1808 = ~(w3747 | w3801);
assign w3803 = v1808;
assign v1809 = ~(w3802 | w3803);
assign w3804 = v1809;
assign v1810 = ~(w3589 | w3658);
assign w3805 = v1810;
assign w3806 = (~w3622 & ~w3623) | (~w3622 & w17082) | (~w3623 & w17082);
assign w3807 = (~w3551 & ~w3553) | (~w3551 & w16869) | (~w3553 & w16869);
assign v1811 = ~(w3571 | w3583);
assign w3808 = v1811;
assign w3809 = (~w3536 & ~w3538) | (~w3536 & w17083) | (~w3538 & w17083);
assign w3810 = ~pi42 & w3600;
assign w3811 = pi42 & w1056;
assign w3812 = pi01 & pi42;
assign v1812 = ~(pi22 | w3812);
assign w3813 = v1812;
assign v1813 = ~(w3811 | w3813);
assign w3814 = v1813;
assign v1814 = ~(w3600 | w3814);
assign w3815 = v1814;
assign v1815 = ~(w3810 | w3815);
assign w3816 = v1815;
assign v1816 = ~(w3539 | w3543);
assign w3817 = v1816;
assign v1817 = ~(w3542 | w3817);
assign w3818 = v1817;
assign w3819 = w3816 & w3818;
assign v1818 = ~(w3816 | w3818);
assign w3820 = v1818;
assign v1819 = ~(w3819 | w3820);
assign w3821 = v1819;
assign w3822 = ~w3809 & w3821;
assign w3823 = w3809 & ~w3821;
assign v1820 = ~(w3822 | w3823);
assign w3824 = v1820;
assign w3825 = ~w3808 & w3824;
assign w3826 = w3808 & ~w3824;
assign v1821 = ~(w3825 | w3826);
assign w3827 = v1821;
assign w3828 = ~w3807 & w3827;
assign w3829 = w3807 & ~w3827;
assign v1822 = ~(w3828 | w3829);
assign w3830 = v1822;
assign w3831 = ~w3806 & w3830;
assign w3832 = w3806 & ~w3830;
assign v1823 = ~(w3831 | w3832);
assign w3833 = v1823;
assign w3834 = ~w3805 & w3833;
assign w3835 = w3805 & ~w3833;
assign v1824 = ~(w3834 | w3835);
assign w3836 = v1824;
assign w3837 = w3804 & w3836;
assign v1825 = ~(w3804 | w3836);
assign w3838 = v1825;
assign v1826 = ~(w3837 | w3838);
assign w3839 = v1826;
assign w3840 = ~w3672 & w3839;
assign w3841 = w3672 & ~w3839;
assign v1827 = ~(w3840 | w3841);
assign w3842 = v1827;
assign w3843 = w3671 & w3842;
assign v1828 = ~(w3671 | w3842);
assign w3844 = v1828;
assign v1829 = ~(w3843 | w3844);
assign w3845 = v1829;
assign v1830 = ~(w3834 | w3837);
assign w3846 = v1830;
assign v1831 = ~(w3745 | w3802);
assign w3847 = v1831;
assign v1832 = ~(w3797 | w3799);
assign w3848 = v1832;
assign v1833 = ~(w3739 | w3742);
assign w3849 = v1833;
assign v1834 = ~(w3675 | w3679);
assign w3850 = v1834;
assign v1835 = ~(w3678 | w3850);
assign w3851 = v1835;
assign v1836 = ~(w3388 | w3731);
assign w3852 = v1836;
assign v1837 = ~(w3730 | w3852);
assign w3853 = v1837;
assign w3854 = w3851 & w3853;
assign v1838 = ~(w3851 | w3853);
assign w3855 = v1838;
assign v1839 = ~(w3854 | w3855);
assign w3856 = v1839;
assign v1840 = ~(w3695 | w3699);
assign w3857 = v1840;
assign v1841 = ~(w3698 | w3857);
assign w3858 = v1841;
assign v1842 = ~(w3856 | w3858);
assign w3859 = v1842;
assign w3860 = w3856 & w3858;
assign v1843 = ~(w3859 | w3860);
assign w3861 = v1843;
assign v1844 = ~(w3725 | w3736);
assign w3862 = v1844;
assign v1845 = ~(w3692 | w3704);
assign w3863 = v1845;
assign v1846 = ~(w3862 | w3863);
assign w3864 = v1846;
assign w3865 = w3862 & w3863;
assign v1847 = ~(w3864 | w3865);
assign w3866 = v1847;
assign w3867 = w3861 & w3866;
assign v1848 = ~(w3861 | w3866);
assign w3868 = v1848;
assign v1849 = ~(w3867 | w3868);
assign w3869 = v1849;
assign w3870 = ~w3849 & w3869;
assign w3871 = w3849 & ~w3869;
assign v1850 = ~(w3870 | w3871);
assign w3872 = v1850;
assign w3873 = ~w3848 & w3872;
assign w3874 = w3848 & ~w3872;
assign v1851 = ~(w3873 | w3874);
assign w3875 = v1851;
assign w3876 = ~w3847 & w3875;
assign w3877 = w3847 & ~w3875;
assign v1852 = ~(w3876 | w3877);
assign w3878 = v1852;
assign w3879 = (~w3828 & ~w3830) | (~w3828 & w17084) | (~w3830 & w17084);
assign v1853 = ~(w3822 | w3825);
assign w3880 = v1853;
assign w3881 = pi03 & pi41;
assign w3882 = pi15 & pi29;
assign w3883 = pi17 & pi27;
assign v1854 = ~(w3882 | w3883);
assign w3884 = v1854;
assign w3885 = w3882 & w3883;
assign v1855 = ~(w3884 | w3885);
assign w3886 = v1855;
assign w3887 = w3881 & ~w3886;
assign w3888 = ~w3881 & w3886;
assign v1856 = ~(w3887 | w3888);
assign w3889 = v1856;
assign w3890 = pi18 & pi26;
assign w3891 = pi19 & pi25;
assign w3892 = pi20 & pi24;
assign v1857 = ~(w3891 | w3892);
assign w3893 = v1857;
assign w3894 = w3891 & w3892;
assign v1858 = ~(w3893 | w3894);
assign w3895 = v1858;
assign w3896 = w3890 & ~w3895;
assign w3897 = ~w3890 & w3895;
assign v1859 = ~(w3896 | w3897);
assign w3898 = v1859;
assign v1860 = ~(w3889 | w3898);
assign w3899 = v1860;
assign w3900 = w3889 & w3898;
assign v1861 = ~(w3899 | w3900);
assign w3901 = v1861;
assign w3902 = pi06 & pi38;
assign w3903 = pi11 & pi33;
assign w3904 = pi07 & pi37;
assign v1862 = ~(w3903 | w3904);
assign w3905 = v1862;
assign w3906 = w3903 & w3904;
assign v1863 = ~(w3905 | w3906);
assign w3907 = v1863;
assign w3908 = w3902 & ~w3907;
assign w3909 = ~w3902 & w3907;
assign v1864 = ~(w3908 | w3909);
assign w3910 = v1864;
assign w3911 = w3901 & ~w3910;
assign w3912 = ~w3901 & w3910;
assign v1865 = ~(w3911 | w3912);
assign w3913 = v1865;
assign w3914 = pi08 & pi36;
assign w3915 = pi10 & pi34;
assign w3916 = pi09 & pi35;
assign v1866 = ~(w3915 | w3916);
assign w3917 = v1866;
assign w3918 = pi10 & pi35;
assign w3919 = w3707 & w3918;
assign v1867 = ~(w3917 | w3919);
assign w3920 = v1867;
assign w3921 = w3914 & ~w3920;
assign w3922 = ~w3914 & w3920;
assign v1868 = ~(w3921 | w3922);
assign w3923 = v1868;
assign w3924 = pi16 & pi28;
assign w3925 = pi04 & pi40;
assign w3926 = pi14 & pi30;
assign v1869 = ~(w3925 | w3926);
assign w3927 = v1869;
assign w3928 = w3925 & w3926;
assign v1870 = ~(w3927 | w3928);
assign w3929 = v1870;
assign w3930 = w3924 & ~w3929;
assign w3931 = ~w3924 & w3929;
assign v1871 = ~(w3930 | w3931);
assign w3932 = v1871;
assign v1872 = ~(w3923 | w3932);
assign w3933 = v1872;
assign w3934 = w3923 & w3932;
assign v1873 = ~(w3933 | w3934);
assign w3935 = v1873;
assign w3936 = pi05 & pi39;
assign w3937 = pi12 & pi32;
assign w3938 = pi13 & pi31;
assign v1874 = ~(w3937 | w3938);
assign w3939 = v1874;
assign w3940 = w3937 & w3938;
assign v1875 = ~(w3939 | w3940);
assign w3941 = v1875;
assign w3942 = w3936 & ~w3941;
assign w3943 = ~w3936 & w3941;
assign v1876 = ~(w3942 | w3943);
assign w3944 = v1876;
assign w3945 = w3935 & ~w3944;
assign w3946 = ~w3935 & w3944;
assign v1877 = ~(w3945 | w3946);
assign w3947 = v1877;
assign w3948 = w3913 & w3947;
assign v1878 = ~(w3913 | w3947);
assign w3949 = v1878;
assign v1879 = ~(w3948 | w3949);
assign w3950 = v1879;
assign w3951 = ~w3880 & w3950;
assign w3952 = w3880 & ~w3950;
assign v1880 = ~(w3951 | w3952);
assign w3953 = v1880;
assign w3954 = ~w3879 & w3953;
assign w3955 = w3879 & ~w3953;
assign v1881 = ~(w3954 | w3955);
assign w3956 = v1881;
assign v1882 = ~(w1755 | w3687);
assign w3957 = v1882;
assign v1883 = ~(w3686 | w3957);
assign w3958 = v1883;
assign v1884 = ~(w3780 | w3784);
assign w3959 = v1884;
assign v1885 = ~(w3783 | w3959);
assign w3960 = v1885;
assign w3961 = w3958 & w3960;
assign v1886 = ~(w3958 | w3960);
assign w3962 = v1886;
assign v1887 = ~(w3961 | w3962);
assign w3963 = v1887;
assign w3964 = pi00 & pi44;
assign w3965 = pi02 & pi42;
assign v1888 = ~(w3964 | w3965);
assign w3966 = v1888;
assign w3967 = pi02 & pi44;
assign w3968 = w3593 & w3967;
assign v1889 = ~(w3966 | w3968);
assign w3969 = v1889;
assign w3970 = w3811 & ~w3969;
assign w3971 = ~w3811 & w3969;
assign v1890 = ~(w3970 | w3971);
assign w3972 = v1890;
assign w3973 = ~w3963 & w3972;
assign w3974 = w3963 & ~w3972;
assign v1891 = ~(w3973 | w3974);
assign w3975 = v1891;
assign w3976 = pi21 & pi23;
assign w3977 = pi01 & pi43;
assign v1892 = ~(w3976 | w3977);
assign w3978 = v1892;
assign w3979 = w3976 & w3977;
assign v1893 = ~(w3978 | w3979);
assign w3980 = v1893;
assign v1894 = ~(w3707 | w3711);
assign w3981 = v1894;
assign v1895 = ~(w3710 | w3981);
assign w3982 = v1895;
assign w3983 = w3980 & w3982;
assign v1896 = ~(w3980 | w3982);
assign w3984 = v1896;
assign v1897 = ~(w3983 | w3984);
assign w3985 = v1897;
assign v1898 = ~(w3716 | w3720);
assign w3986 = v1898;
assign v1899 = ~(w3719 | w3986);
assign w3987 = v1899;
assign w3988 = w3985 & w3987;
assign v1900 = ~(w3985 | w3987);
assign w3989 = v1900;
assign v1901 = ~(w3988 | w3989);
assign w3990 = v1901;
assign w3991 = w3975 & w3990;
assign v1902 = ~(w3975 | w3990);
assign w3992 = v1902;
assign v1903 = ~(w3991 | w3992);
assign w3993 = v1903;
assign w3994 = (~w3789 & ~w3791) | (~w3789 & w16870) | (~w3791 & w16870);
assign w3995 = ~w3993 & w3994;
assign w3996 = w3993 & ~w3994;
assign v1904 = ~(w3995 | w3996);
assign w3997 = v1904;
assign w3998 = (~w3772 & ~w3774) | (~w3772 & w16871) | (~w3774 & w16871);
assign v1905 = ~(w3753 | w3759);
assign w3999 = v1905;
assign w4000 = (~w3766 & ~w3768) | (~w3766 & w16872) | (~w3768 & w16872);
assign w4001 = (~w3810 & ~w3816) | (~w3810 & w17085) | (~w3816 & w17085);
assign v1906 = ~(w4000 | w4001);
assign w4002 = v1906;
assign w4003 = w4000 & w4001;
assign v1907 = ~(w4002 | w4003);
assign w4004 = v1907;
assign w4005 = w3999 & ~w4004;
assign w4006 = ~w3999 & w4004;
assign v1908 = ~(w4005 | w4006);
assign w4007 = v1908;
assign w4008 = ~w3998 & w4007;
assign w4009 = w3998 & ~w4007;
assign v1909 = ~(w4008 | w4009);
assign w4010 = v1909;
assign v1910 = ~(w3997 | w4010);
assign w4011 = v1910;
assign w4012 = w3997 & w4010;
assign v1911 = ~(w4011 | w4012);
assign w4013 = v1911;
assign w4014 = w3956 & w4013;
assign v1912 = ~(w3956 | w4013);
assign w4015 = v1912;
assign v1913 = ~(w4014 | w4015);
assign w4016 = v1913;
assign w4017 = w3878 & w4016;
assign v1914 = ~(w3878 | w4016);
assign w4018 = v1914;
assign v1915 = ~(w4017 | w4018);
assign w4019 = v1915;
assign w4020 = ~w3846 & w4019;
assign w4021 = w3846 & ~w4019;
assign v1916 = ~(w4020 | w4021);
assign w4022 = v1916;
assign v1917 = ~(w3664 | w3841);
assign w4023 = v1917;
assign w4024 = ~w3670 & w4023;
assign v1918 = ~(w3840 | w4024);
assign w4025 = v1918;
assign w4026 = w4022 & w4025;
assign v1919 = ~(w4022 | w4025);
assign w4027 = v1919;
assign v1920 = ~(w4026 | w4027);
assign w4028 = v1920;
assign v1921 = ~(w3840 | w4020);
assign w4029 = v1921;
assign w4030 = (~w3670 & w16521) | (~w3670 & w16522) | (w16521 & w16522);
assign v1922 = ~(w3876 | w4017);
assign w4031 = v1922;
assign w4032 = (~w3983 & ~w3985) | (~w3983 & w17086) | (~w3985 & w17086);
assign w4033 = (~w3961 & ~w3963) | (~w3961 & w16732) | (~w3963 & w16732);
assign w4034 = (~w3854 & ~w3856) | (~w3854 & w16733) | (~w3856 & w16733);
assign v1923 = ~(w4033 | w4034);
assign w4035 = v1923;
assign w4036 = w4033 & w4034;
assign v1924 = ~(w4035 | w4036);
assign w4037 = v1924;
assign w4038 = w4032 & ~w4037;
assign w4039 = ~w4032 & w4037;
assign v1925 = ~(w4038 | w4039);
assign w4040 = v1925;
assign v1926 = ~(w3991 | w3996);
assign w4041 = v1926;
assign w4042 = ~w4040 & w4041;
assign w4043 = w4040 & ~w4041;
assign v1927 = ~(w4042 | w4043);
assign w4044 = v1927;
assign v1928 = ~(w3902 | w3906);
assign w4045 = v1928;
assign v1929 = ~(w3905 | w4045);
assign w4046 = v1929;
assign v1930 = ~(w3924 | w3928);
assign w4047 = v1930;
assign v1931 = ~(w3927 | w4047);
assign w4048 = v1931;
assign w4049 = w4046 & w4048;
assign v1932 = ~(w4046 | w4048);
assign w4050 = v1932;
assign v1933 = ~(w4049 | w4050);
assign w4051 = v1933;
assign v1934 = ~(w3936 | w3940);
assign w4052 = v1934;
assign v1935 = ~(w3939 | w4052);
assign w4053 = v1935;
assign v1936 = ~(w4051 | w4053);
assign w4054 = v1936;
assign w4055 = w4051 & w4053;
assign v1937 = ~(w4054 | w4055);
assign w4056 = v1937;
assign w4057 = (~w3933 & ~w3935) | (~w3933 & w16873) | (~w3935 & w16873);
assign w4058 = (~w3899 & ~w3901) | (~w3899 & w16874) | (~w3901 & w16874);
assign v1938 = ~(w4057 | w4058);
assign w4059 = v1938;
assign w4060 = w4057 & w4058;
assign v1939 = ~(w4059 | w4060);
assign w4061 = v1939;
assign w4062 = w4056 & w4061;
assign v1940 = ~(w4056 | w4061);
assign w4063 = v1940;
assign v1941 = ~(w4062 | w4063);
assign w4064 = v1941;
assign w4065 = w4044 & w4064;
assign v1942 = ~(w4044 | w4064);
assign w4066 = v1942;
assign v1943 = ~(w4065 | w4066);
assign w4067 = v1943;
assign v1944 = ~(w3870 | w3873);
assign w4068 = v1944;
assign v1945 = ~(w3864 | w3867);
assign w4069 = v1945;
assign w4070 = pi00 & pi45;
assign w4071 = pi02 & pi43;
assign w4072 = pi04 & pi41;
assign v1946 = ~(w4071 | w4072);
assign w4073 = v1946;
assign w4074 = w4071 & w4072;
assign v1947 = ~(w4073 | w4074);
assign w4075 = v1947;
assign w4076 = w4070 & ~w4075;
assign w4077 = ~w4070 & w4075;
assign v1948 = ~(w4076 | w4077);
assign w4078 = v1948;
assign w4079 = pi07 & pi38;
assign w4080 = pi08 & pi37;
assign w4081 = pi09 & pi36;
assign v1949 = ~(w4080 | w4081);
assign w4082 = v1949;
assign w4083 = w4080 & w4081;
assign v1950 = ~(w4082 | w4083);
assign w4084 = v1950;
assign w4085 = w4079 & ~w4084;
assign w4086 = ~w4079 & w4084;
assign v1951 = ~(w4085 | w4086);
assign w4087 = v1951;
assign v1952 = ~(w4078 | w4087);
assign w4088 = v1952;
assign w4089 = w4078 & w4087;
assign v1953 = ~(w4088 | w4089);
assign w4090 = v1953;
assign w4091 = pi22 & pi23;
assign w4092 = pi21 & pi24;
assign v1954 = ~(w4091 | w4092);
assign w4093 = v1954;
assign w4094 = w4091 & w4092;
assign v1955 = ~(w4093 | w4094);
assign w4095 = v1955;
assign w4096 = w3918 & ~w4095;
assign w4097 = ~w3918 & w4095;
assign v1956 = ~(w4096 | w4097);
assign w4098 = v1956;
assign w4099 = w4090 & ~w4098;
assign w4100 = ~w4090 & w4098;
assign v1957 = ~(w4099 | w4100);
assign w4101 = v1957;
assign w4102 = w3914 & ~w3917;
assign v1958 = ~(w3919 | w4102);
assign w4103 = v1958;
assign w4104 = pi18 & pi27;
assign w4105 = pi20 & pi25;
assign w4106 = pi19 & pi26;
assign v1959 = ~(w4105 | w4106);
assign w4107 = v1959;
assign w4108 = w4105 & w4106;
assign v1960 = ~(w4107 | w4108);
assign w4109 = v1960;
assign w4110 = w4104 & ~w4109;
assign w4111 = ~w4104 & w4109;
assign v1961 = ~(w4110 | w4111);
assign w4112 = v1961;
assign v1962 = ~(w4103 | w4112);
assign w4113 = v1962;
assign w4114 = w4103 & w4112;
assign v1963 = ~(w4113 | w4114);
assign w4115 = v1963;
assign w4116 = pi14 & pi31;
assign w4117 = pi13 & pi32;
assign w4118 = pi05 & pi40;
assign v1964 = ~(w4117 | w4118);
assign w4119 = v1964;
assign w4120 = w4117 & w4118;
assign v1965 = ~(w4119 | w4120);
assign w4121 = v1965;
assign w4122 = w4116 & ~w4121;
assign w4123 = ~w4116 & w4121;
assign v1966 = ~(w4122 | w4123);
assign w4124 = v1966;
assign w4125 = w4115 & ~w4124;
assign w4126 = ~w4115 & w4124;
assign v1967 = ~(w4125 | w4126);
assign w4127 = v1967;
assign w4128 = w4101 & w4127;
assign v1968 = ~(w4101 | w4127);
assign w4129 = v1968;
assign v1969 = ~(w4128 | w4129);
assign w4130 = v1969;
assign w4131 = ~w4069 & w4130;
assign w4132 = w4069 & ~w4130;
assign v1970 = ~(w4131 | w4132);
assign w4133 = v1970;
assign w4134 = ~w4068 & w4133;
assign w4135 = w4068 & ~w4133;
assign v1971 = ~(w4134 | w4135);
assign w4136 = v1971;
assign w4137 = w4067 & w4136;
assign v1972 = ~(w4067 | w4136);
assign w4138 = v1972;
assign v1973 = ~(w4137 | w4138);
assign w4139 = v1973;
assign v1974 = ~(w3811 | w3968);
assign w4140 = v1974;
assign v1975 = ~(w3966 | w4140);
assign w4141 = v1975;
assign v1976 = ~(w3881 | w3885);
assign w4142 = v1976;
assign v1977 = ~(w3884 | w4142);
assign w4143 = v1977;
assign w4144 = w4141 & w4143;
assign v1978 = ~(w4141 | w4143);
assign w4145 = v1978;
assign v1979 = ~(w4144 | w4145);
assign w4146 = v1979;
assign v1980 = ~(w3890 | w3894);
assign w4147 = v1980;
assign v1981 = ~(w3893 | w4147);
assign w4148 = v1981;
assign v1982 = ~(w4146 | w4148);
assign w4149 = v1982;
assign w4150 = w4146 & w4148;
assign v1983 = ~(w4149 | w4150);
assign w4151 = v1983;
assign v1984 = ~(w4002 | w4006);
assign w4152 = v1984;
assign w4153 = ~w4151 & w4152;
assign w4154 = w4151 & ~w4152;
assign v1985 = ~(w4153 | w4154);
assign w4155 = v1985;
assign w4156 = pi12 & pi33;
assign w4157 = pi11 & pi34;
assign w4158 = pi06 & pi39;
assign v1986 = ~(w4157 | w4158);
assign w4159 = v1986;
assign w4160 = w4157 & w4158;
assign v1987 = ~(w4159 | w4160);
assign w4161 = v1987;
assign w4162 = w4156 & ~w4161;
assign w4163 = ~w4156 & w4161;
assign v1988 = ~(w4162 | w4163);
assign w4164 = v1988;
assign w4165 = pi15 & pi30;
assign w4166 = pi16 & pi29;
assign w4167 = pi17 & pi28;
assign v1989 = ~(w4166 | w4167);
assign w4168 = v1989;
assign w4169 = w4166 & w4167;
assign v1990 = ~(w4168 | w4169);
assign w4170 = v1990;
assign w4171 = w4165 & ~w4170;
assign w4172 = ~w4165 & w4170;
assign v1991 = ~(w4171 | w4172);
assign w4173 = v1991;
assign v1992 = ~(w4164 | w4173);
assign w4174 = v1992;
assign w4175 = w4164 & w4173;
assign v1993 = ~(w4174 | w4175);
assign w4176 = v1993;
assign w4177 = pi44 & w1127;
assign w4178 = pi01 & pi44;
assign v1994 = ~(pi23 | w4178);
assign w4179 = v1994;
assign v1995 = ~(w4177 | w4179);
assign w4180 = v1995;
assign w4181 = pi03 & pi42;
assign v1996 = ~(w3979 | w4181);
assign w4182 = v1996;
assign w4183 = w3979 & w4181;
assign v1997 = ~(w4182 | w4183);
assign w4184 = v1997;
assign w4185 = w4180 & ~w4184;
assign w4186 = ~w4180 & w4184;
assign v1998 = ~(w4185 | w4186);
assign w4187 = v1998;
assign w4188 = w4176 & ~w4187;
assign w4189 = ~w4176 & w4187;
assign v1999 = ~(w4188 | w4189);
assign w4190 = v1999;
assign w4191 = w4155 & w4190;
assign v2000 = ~(w4155 | w4190);
assign w4192 = v2000;
assign v2001 = ~(w4191 | w4192);
assign w4193 = v2001;
assign v2002 = ~(w3948 | w3951);
assign w4194 = v2002;
assign w4195 = (~w4008 & ~w4010) | (~w4008 & w17087) | (~w4010 & w17087);
assign v2003 = ~(w4194 | w4195);
assign w4196 = v2003;
assign w4197 = w4194 & w4195;
assign v2004 = ~(w4196 | w4197);
assign w4198 = v2004;
assign w4199 = w4193 & w4198;
assign v2005 = ~(w4193 | w4198);
assign w4200 = v2005;
assign v2006 = ~(w4199 | w4200);
assign w4201 = v2006;
assign v2007 = ~(w3954 | w4014);
assign w4202 = v2007;
assign w4203 = w4201 & ~w4202;
assign w4204 = ~w4201 & w4202;
assign v2008 = ~(w4203 | w4204);
assign w4205 = v2008;
assign w4206 = w4139 & w4205;
assign v2009 = ~(w4139 | w4205);
assign w4207 = v2009;
assign v2010 = ~(w4206 | w4207);
assign w4208 = v2010;
assign w4209 = ~w4031 & w4208;
assign w4210 = w4031 & ~w4208;
assign v2011 = ~(w4209 | w4210);
assign w4211 = v2011;
assign w4212 = w4030 & ~w4211;
assign w4213 = ~w4030 & w4211;
assign v2012 = ~(w4212 | w4213);
assign w4214 = v2012;
assign w4215 = (w3670 & w16523) | (w3670 & w16524) | (w16523 & w16524);
assign v2013 = ~(w4210 | w4215);
assign w4216 = v2013;
assign v2014 = ~(w4203 | w4206);
assign w4217 = v2014;
assign v2015 = ~(w4134 | w4137);
assign w4218 = v2015;
assign w4219 = (~w4049 & ~w4051) | (~w4049 & w17088) | (~w4051 & w17088);
assign w4220 = pi14 & pi32;
assign w4221 = pi06 & pi40;
assign w4222 = pi13 & pi33;
assign v2016 = ~(w4221 | w4222);
assign w4223 = v2016;
assign w4224 = w4221 & w4222;
assign v2017 = ~(w4223 | w4224);
assign w4225 = v2017;
assign w4226 = w4220 & ~w4225;
assign w4227 = ~w4220 & w4225;
assign v2018 = ~(w4226 | w4227);
assign w4228 = v2018;
assign w4229 = pi15 & pi31;
assign w4230 = pi05 & pi41;
assign v2019 = ~(w4229 | w4230);
assign w4231 = v2019;
assign w4232 = w4229 & w4230;
assign v2020 = ~(w4231 | w4232);
assign w4233 = v2020;
assign w4234 = w3967 & ~w4233;
assign w4235 = ~w3967 & w4233;
assign v2021 = ~(w4234 | w4235);
assign w4236 = v2021;
assign v2022 = ~(w4228 | w4236);
assign w4237 = v2022;
assign w4238 = w4228 & w4236;
assign v2023 = ~(w4237 | w4238);
assign w4239 = v2023;
assign w4240 = w4219 & ~w4239;
assign w4241 = ~w4219 & w4239;
assign v2024 = ~(w4240 | w4241);
assign w4242 = v2024;
assign v2025 = ~(w4104 | w4108);
assign w4243 = v2025;
assign v2026 = ~(w4107 | w4243);
assign w4244 = v2026;
assign v2027 = ~(w4165 | w4169);
assign w4245 = v2027;
assign v2028 = ~(w4168 | w4245);
assign w4246 = v2028;
assign w4247 = w4244 & w4246;
assign v2029 = ~(w4244 | w4246);
assign w4248 = v2029;
assign v2030 = ~(w4247 | w4248);
assign w4249 = v2030;
assign v2031 = ~(w4156 | w4160);
assign w4250 = v2031;
assign v2032 = ~(w4159 | w4250);
assign w4251 = v2032;
assign v2033 = ~(w4249 | w4251);
assign w4252 = v2033;
assign w4253 = w4249 & w4251;
assign v2034 = ~(w4252 | w4253);
assign w4254 = v2034;
assign w4255 = (~w4035 & ~w4037) | (~w4035 & w16875) | (~w4037 & w16875);
assign w4256 = ~w4254 & w4255;
assign w4257 = w4254 & ~w4255;
assign v2035 = ~(w4256 | w4257);
assign w4258 = v2035;
assign w4259 = w4242 & w4258;
assign v2036 = ~(w4242 | w4258);
assign w4260 = v2036;
assign v2037 = ~(w4259 | w4260);
assign w4261 = v2037;
assign w4262 = (~w4043 & ~w4044) | (~w4043 & w17089) | (~w4044 & w17089);
assign v2038 = ~(w4128 | w4131);
assign w4263 = v2038;
assign v2039 = ~(w4262 | w4263);
assign w4264 = v2039;
assign w4265 = w4262 & w4263;
assign v2040 = ~(w4264 | w4265);
assign w4266 = v2040;
assign w4267 = w4261 & w4266;
assign v2041 = ~(w4261 | w4266);
assign w4268 = v2041;
assign v2042 = ~(w4267 | w4268);
assign w4269 = v2042;
assign w4270 = ~w4218 & w4269;
assign w4271 = w4218 & ~w4269;
assign v2043 = ~(w4270 | w4271);
assign w4272 = v2043;
assign w4273 = w4217 & ~w4272;
assign w4274 = ~w4217 & w4272;
assign v2044 = ~(w4273 | w4274);
assign w4275 = v2044;
assign v2045 = ~(w4196 | w4199);
assign w4276 = v2045;
assign w4277 = (~w4059 & ~w4061) | (~w4059 & w17090) | (~w4061 & w17090);
assign w4278 = pi03 & pi43;
assign w4279 = pi00 & pi46;
assign w4280 = pi04 & pi42;
assign v2046 = ~(w4279 | w4280);
assign w4281 = v2046;
assign w4282 = w4279 & w4280;
assign v2047 = ~(w4281 | w4282);
assign w4283 = v2047;
assign w4284 = w4278 & ~w4283;
assign w4285 = ~w4278 & w4283;
assign v2048 = ~(w4284 | w4285);
assign w4286 = v2048;
assign w4287 = pi09 & pi37;
assign w4288 = pi11 & pi35;
assign w4289 = pi10 & pi36;
assign v2049 = ~(w4288 | w4289);
assign w4290 = v2049;
assign w4291 = w4288 & w4289;
assign v2050 = ~(w4290 | w4291);
assign w4292 = v2050;
assign w4293 = w4287 & ~w4292;
assign w4294 = ~w4287 & w4292;
assign v2051 = ~(w4293 | w4294);
assign w4295 = v2051;
assign v2052 = ~(w4286 | w4295);
assign w4296 = v2052;
assign w4297 = w4286 & w4295;
assign v2053 = ~(w4296 | w4297);
assign w4298 = v2053;
assign w4299 = pi19 & pi27;
assign w4300 = pi20 & pi26;
assign w4301 = pi21 & pi25;
assign v2054 = ~(w4300 | w4301);
assign w4302 = v2054;
assign w4303 = w4300 & w4301;
assign v2055 = ~(w4302 | w4303);
assign w4304 = v2055;
assign w4305 = w4299 & ~w4304;
assign w4306 = ~w4299 & w4304;
assign v2056 = ~(w4305 | w4306);
assign w4307 = v2056;
assign w4308 = w4298 & ~w4307;
assign w4309 = ~w4298 & w4307;
assign v2057 = ~(w4308 | w4309);
assign w4310 = v2057;
assign w4311 = pi16 & pi30;
assign w4312 = pi17 & pi29;
assign w4313 = pi18 & pi28;
assign v2058 = ~(w4312 | w4313);
assign w4314 = v2058;
assign w4315 = w4312 & w4313;
assign v2059 = ~(w4314 | w4315);
assign w4316 = v2059;
assign w4317 = w4311 & ~w4316;
assign w4318 = ~w4311 & w4316;
assign v2060 = ~(w4317 | w4318);
assign w4319 = v2060;
assign v2061 = ~(w4180 | w4183);
assign w4320 = v2061;
assign v2062 = ~(w4182 | w4320);
assign w4321 = v2062;
assign w4322 = ~w4319 & w4321;
assign w4323 = w4319 & ~w4321;
assign v2063 = ~(w4322 | w4323);
assign w4324 = v2063;
assign w4325 = pi12 & pi34;
assign w4326 = pi08 & pi38;
assign w4327 = pi07 & pi39;
assign v2064 = ~(w4326 | w4327);
assign w4328 = v2064;
assign w4329 = pi08 & pi39;
assign w4330 = w4079 & w4329;
assign v2065 = ~(w4328 | w4330);
assign w4331 = v2065;
assign w4332 = w4325 & ~w4331;
assign w4333 = ~w4325 & w4331;
assign v2066 = ~(w4332 | w4333);
assign w4334 = v2066;
assign w4335 = w4324 & ~w4334;
assign w4336 = ~w4324 & w4334;
assign v2067 = ~(w4335 | w4336);
assign w4337 = v2067;
assign w4338 = w4310 & w4337;
assign v2068 = ~(w4310 | w4337);
assign w4339 = v2068;
assign v2069 = ~(w4338 | w4339);
assign w4340 = v2069;
assign w4341 = ~w4277 & w4340;
assign w4342 = w4277 & ~w4340;
assign v2070 = ~(w4341 | w4342);
assign w4343 = v2070;
assign w4344 = ~w4276 & w4343;
assign w4345 = w4276 & ~w4343;
assign v2071 = ~(w4344 | w4345);
assign w4346 = v2071;
assign v2072 = ~(w4174 | w4188);
assign w4347 = v2072;
assign v2073 = ~(w4113 | w4125);
assign w4348 = v2073;
assign v2074 = ~(w4088 | w4099);
assign w4349 = v2074;
assign v2075 = ~(w4348 | w4349);
assign w4350 = v2075;
assign w4351 = w4348 & w4349;
assign v2076 = ~(w4350 | w4351);
assign w4352 = v2076;
assign w4353 = w4347 & ~w4352;
assign w4354 = ~w4347 & w4352;
assign v2077 = ~(w4353 | w4354);
assign w4355 = v2077;
assign v2078 = ~(w4154 | w4191);
assign w4356 = v2078;
assign v2079 = ~(w4116 | w4120);
assign w4357 = v2079;
assign v2080 = ~(w4119 | w4357);
assign w4358 = v2080;
assign v2081 = ~(w4070 | w4074);
assign w4359 = v2081;
assign v2082 = ~(w4073 | w4359);
assign w4360 = v2082;
assign w4361 = w4358 & w4360;
assign v2083 = ~(w4358 | w4360);
assign w4362 = v2083;
assign v2084 = ~(w4361 | w4362);
assign w4363 = v2084;
assign v2085 = ~(w4079 | w4083);
assign w4364 = v2085;
assign v2086 = ~(w4082 | w4364);
assign w4365 = v2086;
assign v2087 = ~(w4363 | w4365);
assign w4366 = v2087;
assign w4367 = w4363 & w4365;
assign v2088 = ~(w4366 | w4367);
assign w4368 = v2088;
assign w4369 = (~w4144 & ~w4146) | (~w4144 & w17091) | (~w4146 & w17091);
assign w4370 = pi22 & pi24;
assign w4371 = pi01 & pi45;
assign v2089 = ~(w4370 | w4371);
assign w4372 = v2089;
assign w4373 = w4370 & w4371;
assign v2090 = ~(w4372 | w4373);
assign w4374 = v2090;
assign w4375 = w4177 & w4374;
assign v2091 = ~(w4177 | w4374);
assign w4376 = v2091;
assign v2092 = ~(w4375 | w4376);
assign w4377 = v2092;
assign v2093 = ~(w3918 | w4094);
assign w4378 = v2093;
assign v2094 = ~(w4093 | w4378);
assign w4379 = v2094;
assign w4380 = w4377 & w4379;
assign v2095 = ~(w4377 | w4379);
assign w4381 = v2095;
assign v2096 = ~(w4380 | w4381);
assign w4382 = v2096;
assign w4383 = ~w4369 & w4382;
assign w4384 = w4369 & ~w4382;
assign v2097 = ~(w4383 | w4384);
assign w4385 = v2097;
assign w4386 = w4368 & w4385;
assign v2098 = ~(w4368 | w4385);
assign w4387 = v2098;
assign v2099 = ~(w4386 | w4387);
assign w4388 = v2099;
assign w4389 = ~w4356 & w4388;
assign w4390 = w4356 & ~w4388;
assign v2100 = ~(w4389 | w4390);
assign w4391 = v2100;
assign w4392 = w4355 & w4391;
assign v2101 = ~(w4355 | w4391);
assign w4393 = v2101;
assign v2102 = ~(w4392 | w4393);
assign w4394 = v2102;
assign w4395 = w4346 & w4394;
assign v2103 = ~(w4346 | w4394);
assign w4396 = v2103;
assign v2104 = ~(w4395 | w4396);
assign w4397 = v2104;
assign v2105 = ~(w4275 | w4397);
assign w4398 = v2105;
assign w4399 = w4275 & w4397;
assign v2106 = ~(w4398 | w4399);
assign w4400 = v2106;
assign w4401 = w4216 & ~w4400;
assign w4402 = ~w4216 & w4400;
assign v2107 = ~(w4401 | w4402);
assign w4403 = v2107;
assign v2108 = ~(w4270 | w4274);
assign w4404 = v2108;
assign v2109 = ~(w3967 | w4232);
assign w4405 = v2109;
assign v2110 = ~(w4231 | w4405);
assign w4406 = v2110;
assign v2111 = ~(w4299 | w4303);
assign w4407 = v2111;
assign v2112 = ~(w4302 | w4407);
assign w4408 = v2112;
assign w4409 = w4406 & w4408;
assign v2113 = ~(w4406 | w4408);
assign w4410 = v2113;
assign v2114 = ~(w4409 | w4410);
assign w4411 = v2114;
assign v2115 = ~(w4278 | w4282);
assign w4412 = v2115;
assign v2116 = ~(w4281 | w4412);
assign w4413 = v2116;
assign v2117 = ~(w4411 | w4413);
assign w4414 = v2117;
assign w4415 = w4411 & w4413;
assign v2118 = ~(w4414 | w4415);
assign w4416 = v2118;
assign w4417 = (~w4296 & ~w4298) | (~w4296 & w16876) | (~w4298 & w16876);
assign w4418 = ~w4416 & w4417;
assign w4419 = w4416 & ~w4417;
assign v2119 = ~(w4418 | w4419);
assign w4420 = v2119;
assign v2120 = ~(w4237 | w4241);
assign w4421 = v2120;
assign w4422 = ~w4420 & w4421;
assign w4423 = w4420 & ~w4421;
assign v2121 = ~(w4422 | w4423);
assign w4424 = v2121;
assign v2122 = ~(w4338 | w4341);
assign w4425 = v2122;
assign w4426 = (~w4257 & ~w4258) | (~w4257 & w17092) | (~w4258 & w17092);
assign v2123 = ~(w4425 | w4426);
assign w4427 = v2123;
assign w4428 = w4425 & w4426;
assign v2124 = ~(w4427 | w4428);
assign w4429 = v2124;
assign w4430 = w4424 & w4429;
assign v2125 = ~(w4424 | w4429);
assign w4431 = v2125;
assign v2126 = ~(w4430 | w4431);
assign w4432 = v2126;
assign v2127 = ~(w4264 | w4267);
assign w4433 = v2127;
assign v2128 = ~(w4389 | w4392);
assign w4434 = v2128;
assign v2129 = ~(w4433 | w4434);
assign w4435 = v2129;
assign w4436 = w4433 & w4434;
assign v2130 = ~(w4435 | w4436);
assign w4437 = v2130;
assign w4438 = w4432 & w4437;
assign v2131 = ~(w4432 | w4437);
assign w4439 = v2131;
assign v2132 = ~(w4438 | w4439);
assign w4440 = v2132;
assign v2133 = ~(w4344 | w4395);
assign w4441 = v2133;
assign w4442 = (~w4247 & ~w4249) | (~w4247 & w17093) | (~w4249 & w17093);
assign w4443 = (~w4375 & ~w4377) | (~w4375 & w16877) | (~w4377 & w16877);
assign w4444 = pi13 & pi34;
assign w4445 = pi12 & pi35;
assign w4446 = pi07 & pi40;
assign v2134 = ~(w4445 | w4446);
assign w4447 = v2134;
assign w4448 = w4445 & w4446;
assign v2135 = ~(w4447 | w4448);
assign w4449 = v2135;
assign w4450 = w4444 & ~w4449;
assign w4451 = ~w4444 & w4449;
assign v2136 = ~(w4450 | w4451);
assign w4452 = v2136;
assign v2137 = ~(w4443 | w4452);
assign w4453 = v2137;
assign w4454 = w4443 & w4452;
assign v2138 = ~(w4453 | w4454);
assign w4455 = v2138;
assign w4456 = w4442 & ~w4455;
assign w4457 = ~w4442 & w4455;
assign v2139 = ~(w4456 | w4457);
assign w4458 = v2139;
assign v2140 = ~(w4383 | w4386);
assign w4459 = v2140;
assign w4460 = ~w4458 & w4459;
assign w4461 = w4458 & ~w4459;
assign v2141 = ~(w4460 | w4461);
assign w4462 = v2141;
assign v2142 = ~(w4350 | w4354);
assign w4463 = v2142;
assign w4464 = ~w4462 & w4463;
assign w4465 = w4462 & ~w4463;
assign v2143 = ~(w4464 | w4465);
assign w4466 = v2143;
assign w4467 = pi01 & pi46;
assign v2144 = ~(pi24 | w4467);
assign w4468 = v2144;
assign w4469 = pi46 & w1215;
assign v2145 = ~(w4468 | w4469);
assign w4470 = v2145;
assign v2146 = ~(w4287 | w4291);
assign w4471 = v2146;
assign v2147 = ~(w4290 | w4471);
assign w4472 = v2147;
assign w4473 = w4470 & w4472;
assign v2148 = ~(w4470 | w4472);
assign w4474 = v2148;
assign v2149 = ~(w4473 | w4474);
assign w4475 = v2149;
assign w4476 = w4325 & ~w4328;
assign v2150 = ~(w4330 | w4476);
assign w4477 = v2150;
assign w4478 = w4475 & ~w4477;
assign w4479 = ~w4475 & w4477;
assign v2151 = ~(w4478 | w4479);
assign w4480 = v2151;
assign w4481 = (~w4322 & ~w4324) | (~w4322 & w16878) | (~w4324 & w16878);
assign w4482 = (~w4361 & ~w4363) | (~w4361 & w17094) | (~w4363 & w17094);
assign v2152 = ~(w4481 | w4482);
assign w4483 = v2152;
assign w4484 = w4481 & w4482;
assign v2153 = ~(w4483 | w4484);
assign w4485 = v2153;
assign v2154 = ~(w4480 | w4485);
assign w4486 = v2154;
assign w4487 = w4480 & w4485;
assign v2155 = ~(w4486 | w4487);
assign w4488 = v2155;
assign w4489 = pi00 & pi47;
assign w4490 = pi02 & pi45;
assign v2156 = ~(w4489 | w4490);
assign w4491 = v2156;
assign w4492 = pi02 & pi47;
assign w4493 = w4070 & w4492;
assign v2157 = ~(w4491 | w4493);
assign w4494 = v2157;
assign w4495 = w4373 & ~w4494;
assign w4496 = ~w4373 & w4494;
assign v2158 = ~(w4495 | w4496);
assign w4497 = v2158;
assign w4498 = pi16 & pi31;
assign w4499 = pi18 & pi29;
assign w4500 = pi17 & pi30;
assign v2159 = ~(w4499 | w4500);
assign w4501 = v2159;
assign w4502 = w4499 & w4500;
assign v2160 = ~(w4501 | w4502);
assign w4503 = v2160;
assign w4504 = w4498 & ~w4503;
assign w4505 = ~w4498 & w4503;
assign v2161 = ~(w4504 | w4505);
assign w4506 = v2161;
assign v2162 = ~(w4497 | w4506);
assign w4507 = v2162;
assign w4508 = w4497 & w4506;
assign v2163 = ~(w4507 | w4508);
assign w4509 = v2163;
assign w4510 = pi19 & pi28;
assign w4511 = pi21 & pi26;
assign w4512 = pi20 & pi27;
assign v2164 = ~(w4511 | w4512);
assign w4513 = v2164;
assign w4514 = w4511 & w4512;
assign v2165 = ~(w4513 | w4514);
assign w4515 = v2165;
assign w4516 = w4510 & ~w4515;
assign w4517 = ~w4510 & w4515;
assign v2166 = ~(w4516 | w4517);
assign w4518 = v2166;
assign w4519 = w4509 & ~w4518;
assign w4520 = ~w4509 & w4518;
assign v2167 = ~(w4519 | w4520);
assign w4521 = v2167;
assign v2168 = ~(w4311 | w4315);
assign w4522 = v2168;
assign v2169 = ~(w4314 | w4522);
assign w4523 = v2169;
assign v2170 = ~(w4220 | w4224);
assign w4524 = v2170;
assign v2171 = ~(w4223 | w4524);
assign w4525 = v2171;
assign w4526 = w4523 & w4525;
assign v2172 = ~(w4523 | w4525);
assign w4527 = v2172;
assign v2173 = ~(w4526 | w4527);
assign w4528 = v2173;
assign w4529 = pi03 & pi44;
assign w4530 = pi04 & pi43;
assign w4531 = pi15 & pi32;
assign v2174 = ~(w4530 | w4531);
assign w4532 = v2174;
assign w4533 = w4530 & w4531;
assign v2175 = ~(w4532 | w4533);
assign w4534 = v2175;
assign w4535 = w4529 & ~w4534;
assign w4536 = ~w4529 & w4534;
assign v2176 = ~(w4535 | w4536);
assign w4537 = v2176;
assign w4538 = ~w4528 & w4537;
assign w4539 = w4528 & ~w4537;
assign v2177 = ~(w4538 | w4539);
assign w4540 = v2177;
assign w4541 = pi10 & pi37;
assign w4542 = pi23 & pi24;
assign w4543 = pi22 & pi25;
assign v2178 = ~(w4542 | w4543);
assign w4544 = v2178;
assign w4545 = w4542 & w4543;
assign v2179 = ~(w4544 | w4545);
assign w4546 = v2179;
assign w4547 = w4541 & ~w4546;
assign w4548 = ~w4541 & w4546;
assign v2180 = ~(w4547 | w4548);
assign w4549 = v2180;
assign w4550 = pi11 & pi36;
assign w4551 = pi09 & pi38;
assign v2181 = ~(w4550 | w4551);
assign w4552 = v2181;
assign w4553 = w4550 & w4551;
assign v2182 = ~(w4552 | w4553);
assign w4554 = v2182;
assign w4555 = w4329 & ~w4554;
assign w4556 = ~w4329 & w4554;
assign v2183 = ~(w4555 | w4556);
assign w4557 = v2183;
assign v2184 = ~(w4549 | w4557);
assign w4558 = v2184;
assign w4559 = w4549 & w4557;
assign v2185 = ~(w4558 | w4559);
assign w4560 = v2185;
assign w4561 = pi05 & pi42;
assign w4562 = pi06 & pi41;
assign w4563 = pi14 & pi33;
assign v2186 = ~(w4562 | w4563);
assign w4564 = v2186;
assign w4565 = w4562 & w4563;
assign v2187 = ~(w4564 | w4565);
assign w4566 = v2187;
assign w4567 = w4561 & ~w4566;
assign w4568 = ~w4561 & w4566;
assign v2188 = ~(w4567 | w4568);
assign w4569 = v2188;
assign w4570 = w4560 & ~w4569;
assign w4571 = ~w4560 & w4569;
assign v2189 = ~(w4570 | w4571);
assign w4572 = v2189;
assign w4573 = w4540 & w4572;
assign v2190 = ~(w4540 | w4572);
assign w4574 = v2190;
assign v2191 = ~(w4573 | w4574);
assign w4575 = v2191;
assign w4576 = w4521 & w4575;
assign v2192 = ~(w4521 | w4575);
assign w4577 = v2192;
assign v2193 = ~(w4576 | w4577);
assign w4578 = v2193;
assign w4579 = w4488 & w4578;
assign v2194 = ~(w4488 | w4578);
assign w4580 = v2194;
assign v2195 = ~(w4579 | w4580);
assign w4581 = v2195;
assign w4582 = w4466 & w4581;
assign v2196 = ~(w4466 | w4581);
assign w4583 = v2196;
assign v2197 = ~(w4582 | w4583);
assign w4584 = v2197;
assign w4585 = ~w4441 & w4584;
assign w4586 = w4441 & ~w4584;
assign v2198 = ~(w4585 | w4586);
assign w4587 = v2198;
assign w4588 = w4440 & w4587;
assign v2199 = ~(w4440 | w4587);
assign w4589 = v2199;
assign v2200 = ~(w4588 | w4589);
assign w4590 = v2200;
assign w4591 = ~w4404 & w4590;
assign w4592 = w4404 & ~w4590;
assign v2201 = ~(w4591 | w4592);
assign w4593 = v2201;
assign v2202 = ~(w4210 | w4398);
assign w4594 = v2202;
assign w4595 = ~w4215 & w4594;
assign v2203 = ~(w4399 | w4595);
assign w4596 = v2203;
assign w4597 = w4593 & w4596;
assign v2204 = ~(w4593 | w4596);
assign w4598 = v2204;
assign v2205 = ~(w4597 | w4598);
assign w4599 = v2205;
assign v2206 = ~(w4399 | w4591);
assign w4600 = v2206;
assign w4601 = (~w4215 & w16526) | (~w4215 & w16527) | (w16526 & w16527);
assign v2207 = ~(w4585 | w4588);
assign w4602 = v2207;
assign v2208 = ~(w4435 | w4438);
assign w4603 = v2208;
assign v2209 = ~(w4427 | w4430);
assign w4604 = v2209;
assign v2210 = ~(w4461 | w4465);
assign w4605 = v2210;
assign w4606 = (~w4453 & ~w4455) | (~w4453 & w17095) | (~w4455 & w17095);
assign w4607 = pi14 & pi34;
assign w4608 = pi06 & pi42;
assign w4609 = pi13 & pi35;
assign v2211 = ~(w4608 | w4609);
assign w4610 = v2211;
assign w4611 = w4608 & w4609;
assign v2212 = ~(w4610 | w4611);
assign w4612 = v2212;
assign w4613 = w4607 & ~w4612;
assign w4614 = ~w4607 & w4612;
assign v2213 = ~(w4613 | w4614);
assign w4615 = v2213;
assign w4616 = pi07 & pi41;
assign w4617 = pi12 & pi36;
assign w4618 = pi08 & pi40;
assign v2214 = ~(w4617 | w4618);
assign w4619 = v2214;
assign w4620 = w4617 & w4618;
assign v2215 = ~(w4619 | w4620);
assign w4621 = v2215;
assign w4622 = w4616 & ~w4621;
assign w4623 = ~w4616 & w4621;
assign v2216 = ~(w4622 | w4623);
assign w4624 = v2216;
assign v2217 = ~(w4615 | w4624);
assign w4625 = v2217;
assign w4626 = w4615 & w4624;
assign v2218 = ~(w4625 | w4626);
assign w4627 = v2218;
assign w4628 = pi09 & pi39;
assign w4629 = pi11 & pi37;
assign w4630 = pi10 & pi38;
assign v2219 = ~(w4629 | w4630);
assign w4631 = v2219;
assign w4632 = pi11 & pi38;
assign w4633 = w4541 & w4632;
assign v2220 = ~(w4631 | w4633);
assign w4634 = v2220;
assign w4635 = w4628 & ~w4634;
assign w4636 = ~w4628 & w4634;
assign v2221 = ~(w4635 | w4636);
assign w4637 = v2221;
assign w4638 = w4627 & ~w4637;
assign w4639 = ~w4627 & w4637;
assign v2222 = ~(w4638 | w4639);
assign w4640 = v2222;
assign w4641 = ~w4606 & w4640;
assign w4642 = w4606 & ~w4640;
assign v2223 = ~(w4641 | w4642);
assign w4643 = v2223;
assign w4644 = pi04 & pi44;
assign w4645 = pi05 & pi43;
assign w4646 = pi15 & pi33;
assign v2224 = ~(w4645 | w4646);
assign w4647 = v2224;
assign w4648 = w4645 & w4646;
assign v2225 = ~(w4647 | w4648);
assign w4649 = v2225;
assign w4650 = w4644 & ~w4649;
assign w4651 = ~w4644 & w4649;
assign v2226 = ~(w4650 | w4651);
assign w4652 = v2226;
assign w4653 = pi20 & pi28;
assign w4654 = pi21 & pi27;
assign w4655 = pi22 & pi26;
assign v2227 = ~(w4654 | w4655);
assign w4656 = v2227;
assign w4657 = w4654 & w4655;
assign v2228 = ~(w4656 | w4657);
assign w4658 = v2228;
assign w4659 = w4653 & ~w4658;
assign w4660 = ~w4653 & w4658;
assign v2229 = ~(w4659 | w4660);
assign w4661 = v2229;
assign v2230 = ~(w4652 | w4661);
assign w4662 = v2230;
assign w4663 = w4652 & w4661;
assign v2231 = ~(w4662 | w4663);
assign w4664 = v2231;
assign w4665 = pi17 & pi31;
assign w4666 = pi18 & pi30;
assign w4667 = pi19 & pi29;
assign v2232 = ~(w4666 | w4667);
assign w4668 = v2232;
assign w4669 = w4666 & w4667;
assign v2233 = ~(w4668 | w4669);
assign w4670 = v2233;
assign w4671 = w4665 & ~w4670;
assign w4672 = ~w4665 & w4670;
assign v2234 = ~(w4671 | w4672);
assign w4673 = v2234;
assign w4674 = w4664 & ~w4673;
assign w4675 = ~w4664 & w4673;
assign v2235 = ~(w4674 | w4675);
assign w4676 = v2235;
assign v2236 = ~(w4643 | w4676);
assign w4677 = v2236;
assign w4678 = w4643 & w4676;
assign v2237 = ~(w4677 | w4678);
assign w4679 = v2237;
assign w4680 = ~w4605 & w4679;
assign w4681 = w4605 & ~w4679;
assign v2238 = ~(w4680 | w4681);
assign w4682 = v2238;
assign w4683 = ~w4604 & w4682;
assign w4684 = w4604 & ~w4682;
assign v2239 = ~(w4683 | w4684);
assign w4685 = v2239;
assign w4686 = ~w4603 & w4685;
assign w4687 = w4603 & ~w4685;
assign v2240 = ~(w4686 | w4687);
assign w4688 = v2240;
assign v2241 = ~(w4510 | w4514);
assign w4689 = v2241;
assign v2242 = ~(w4513 | w4689);
assign w4690 = v2242;
assign v2243 = ~(w4329 | w4553);
assign w4691 = v2243;
assign v2244 = ~(w4552 | w4691);
assign w4692 = v2244;
assign w4693 = w4690 & w4692;
assign v2245 = ~(w4690 | w4692);
assign w4694 = v2245;
assign v2246 = ~(w4693 | w4694);
assign w4695 = v2246;
assign v2247 = ~(w4561 | w4565);
assign w4696 = v2247;
assign v2248 = ~(w4564 | w4696);
assign w4697 = v2248;
assign v2249 = ~(w4695 | w4697);
assign w4698 = v2249;
assign w4699 = w4695 & w4697;
assign v2250 = ~(w4698 | w4699);
assign w4700 = v2250;
assign w4701 = (~w4558 & ~w4560) | (~w4558 & w16879) | (~w4560 & w16879);
assign w4702 = ~w4700 & w4701;
assign w4703 = w4700 & ~w4701;
assign v2251 = ~(w4702 | w4703);
assign w4704 = v2251;
assign v2252 = ~(w4444 | w4448);
assign w4705 = v2252;
assign v2253 = ~(w4447 | w4705);
assign w4706 = v2253;
assign v2254 = ~(w4541 | w4545);
assign w4707 = v2254;
assign v2255 = ~(w4544 | w4707);
assign w4708 = v2255;
assign w4709 = w4706 & w4708;
assign v2256 = ~(w4706 | w4708);
assign w4710 = v2256;
assign v2257 = ~(w4709 | w4710);
assign w4711 = v2257;
assign w4712 = pi02 & pi46;
assign w4713 = pi03 & pi45;
assign w4714 = pi16 & pi32;
assign v2258 = ~(w4713 | w4714);
assign w4715 = v2258;
assign w4716 = w4713 & w4714;
assign v2259 = ~(w4715 | w4716);
assign w4717 = v2259;
assign w4718 = w4712 & ~w4717;
assign w4719 = ~w4712 & w4717;
assign v2260 = ~(w4718 | w4719);
assign w4720 = v2260;
assign w4721 = ~w4711 & w4720;
assign w4722 = w4711 & ~w4720;
assign v2261 = ~(w4721 | w4722);
assign w4723 = v2261;
assign v2262 = ~(w4704 | w4723);
assign w4724 = v2262;
assign w4725 = w4704 & w4723;
assign v2263 = ~(w4724 | w4725);
assign w4726 = v2263;
assign v2264 = ~(w4573 | w4576);
assign w4727 = v2264;
assign w4728 = ~w4726 & w4727;
assign w4729 = w4726 & ~w4727;
assign v2265 = ~(w4728 | w4729);
assign w4730 = v2265;
assign v2266 = ~(w4498 | w4502);
assign w4731 = v2266;
assign v2267 = ~(w4501 | w4731);
assign w4732 = v2267;
assign v2268 = ~(w4529 | w4533);
assign w4733 = v2268;
assign v2269 = ~(w4532 | w4733);
assign w4734 = v2269;
assign w4735 = w4732 & w4734;
assign v2270 = ~(w4732 | w4734);
assign w4736 = v2270;
assign v2271 = ~(w4735 | w4736);
assign w4737 = v2271;
assign w4738 = w4373 & ~w4491;
assign v2272 = ~(w4493 | w4738);
assign w4739 = v2272;
assign w4740 = ~w4737 & w4739;
assign w4741 = w4737 & ~w4739;
assign v2273 = ~(w4740 | w4741);
assign w4742 = v2273;
assign w4743 = (~w4473 & ~w4475) | (~w4473 & w17096) | (~w4475 & w17096);
assign w4744 = (~w4507 & ~w4509) | (~w4507 & w16880) | (~w4509 & w16880);
assign v2274 = ~(w4743 | w4744);
assign w4745 = v2274;
assign w4746 = w4743 & w4744;
assign v2275 = ~(w4745 | w4746);
assign w4747 = v2275;
assign w4748 = w4742 & w4747;
assign v2276 = ~(w4742 | w4747);
assign w4749 = v2276;
assign v2277 = ~(w4748 | w4749);
assign w4750 = v2277;
assign w4751 = w4730 & w4750;
assign v2278 = ~(w4730 | w4750);
assign w4752 = v2278;
assign v2279 = ~(w4751 | w4752);
assign w4753 = v2279;
assign v2280 = ~(w4579 | w4582);
assign w4754 = v2280;
assign w4755 = (~w4526 & ~w4528) | (~w4526 & w17097) | (~w4528 & w17097);
assign w4756 = (~w4409 & ~w4411) | (~w4409 & w16734) | (~w4411 & w16734);
assign w4757 = pi00 & pi48;
assign w4758 = w4469 & w4757;
assign v2281 = ~(w4469 | w4757);
assign w4759 = v2281;
assign v2282 = ~(w4758 | w4759);
assign w4760 = v2282;
assign w4761 = pi23 & pi25;
assign w4762 = pi01 & pi47;
assign v2283 = ~(w4761 | w4762);
assign w4763 = v2283;
assign w4764 = w4761 & w4762;
assign v2284 = ~(w4763 | w4764);
assign w4765 = v2284;
assign w4766 = w4760 & w4765;
assign v2285 = ~(w4760 | w4765);
assign w4767 = v2285;
assign v2286 = ~(w4766 | w4767);
assign w4768 = v2286;
assign w4769 = ~w4756 & w4768;
assign w4770 = w4756 & ~w4768;
assign v2287 = ~(w4769 | w4770);
assign w4771 = v2287;
assign w4772 = w4755 & ~w4771;
assign w4773 = ~w4755 & w4771;
assign v2288 = ~(w4772 | w4773);
assign w4774 = v2288;
assign w4775 = (~w4419 & ~w4420) | (~w4419 & w17098) | (~w4420 & w17098);
assign w4776 = (~w4483 & ~w4485) | (~w4483 & w17099) | (~w4485 & w17099);
assign v2289 = ~(w4775 | w4776);
assign w4777 = v2289;
assign w4778 = w4775 & w4776;
assign v2290 = ~(w4777 | w4778);
assign w4779 = v2290;
assign w4780 = w4774 & w4779;
assign v2291 = ~(w4774 | w4779);
assign w4781 = v2291;
assign v2292 = ~(w4780 | w4781);
assign w4782 = v2292;
assign w4783 = ~w4754 & w4782;
assign w4784 = w4754 & ~w4782;
assign v2293 = ~(w4783 | w4784);
assign w4785 = v2293;
assign w4786 = w4753 & w4785;
assign v2294 = ~(w4753 | w4785);
assign w4787 = v2294;
assign v2295 = ~(w4786 | w4787);
assign w4788 = v2295;
assign w4789 = w4688 & w4788;
assign v2296 = ~(w4688 | w4788);
assign w4790 = v2296;
assign v2297 = ~(w4789 | w4790);
assign w4791 = v2297;
assign w4792 = w4602 & ~w4791;
assign w4793 = ~w4602 & w4791;
assign v2298 = ~(w4792 | w4793);
assign w4794 = v2298;
assign w4795 = w4601 & ~w4794;
assign w4796 = ~w4601 & w4794;
assign v2299 = ~(w4795 | w4796);
assign w4797 = v2299;
assign v2300 = ~(w4601 | w4793);
assign w4798 = v2300;
assign v2301 = ~(w4792 | w4798);
assign w4799 = v2301;
assign v2302 = ~(w4783 | w4786);
assign w4800 = v2302;
assign v2303 = ~(w4729 | w4751);
assign w4801 = v2303;
assign v2304 = ~(w4777 | w4780);
assign w4802 = v2304;
assign w4803 = pi22 & pi27;
assign w4804 = pi03 & pi46;
assign v2305 = ~(w4492 | w4804);
assign w4805 = v2305;
assign w4806 = pi03 & pi47;
assign w4807 = w4712 & w4806;
assign v2306 = ~(w4805 | w4807);
assign w4808 = v2306;
assign w4809 = w4803 & ~w4808;
assign w4810 = ~w4803 & w4808;
assign v2307 = ~(w4809 | w4810);
assign w4811 = v2307;
assign w4812 = pi19 & pi30;
assign w4813 = pi21 & pi28;
assign w4814 = pi20 & pi29;
assign v2308 = ~(w4813 | w4814);
assign w4815 = v2308;
assign w4816 = w4813 & w4814;
assign v2309 = ~(w4815 | w4816);
assign w4817 = v2309;
assign w4818 = w4812 & ~w4817;
assign w4819 = ~w4812 & w4817;
assign v2310 = ~(w4818 | w4819);
assign w4820 = v2310;
assign v2311 = ~(w4811 | w4820);
assign w4821 = v2311;
assign w4822 = w4811 & w4820;
assign v2312 = ~(w4821 | w4822);
assign w4823 = v2312;
assign w4824 = pi09 & pi40;
assign w4825 = pi12 & pi37;
assign w4826 = pi10 & pi39;
assign v2313 = ~(w4825 | w4826);
assign w4827 = v2313;
assign w4828 = w4825 & w4826;
assign v2314 = ~(w4827 | w4828);
assign w4829 = v2314;
assign w4830 = w4824 & ~w4829;
assign w4831 = ~w4824 & w4829;
assign v2315 = ~(w4830 | w4831);
assign w4832 = v2315;
assign w4833 = w4823 & ~w4832;
assign w4834 = ~w4823 & w4832;
assign v2316 = ~(w4833 | w4834);
assign w4835 = v2316;
assign w4836 = (~w4758 & ~w4760) | (~w4758 & w16735) | (~w4760 & w16735);
assign w4837 = pi00 & pi49;
assign w4838 = pi04 & pi45;
assign w4839 = pi05 & pi44;
assign v2317 = ~(w4838 | w4839);
assign w4840 = v2317;
assign w4841 = pi05 & pi45;
assign w4842 = w4644 & w4841;
assign v2318 = ~(w4840 | w4842);
assign w4843 = v2318;
assign w4844 = w4837 & ~w4843;
assign w4845 = ~w4837 & w4843;
assign v2319 = ~(w4844 | w4845);
assign w4846 = v2319;
assign v2320 = ~(w4836 | w4846);
assign w4847 = v2320;
assign w4848 = w4836 & w4846;
assign v2321 = ~(w4847 | w4848);
assign w4849 = v2321;
assign w4850 = pi16 & pi33;
assign w4851 = pi17 & pi32;
assign w4852 = pi18 & pi31;
assign v2322 = ~(w4851 | w4852);
assign w4853 = v2322;
assign w4854 = w4851 & w4852;
assign v2323 = ~(w4853 | w4854);
assign w4855 = v2323;
assign w4856 = w4850 & ~w4855;
assign w4857 = ~w4850 & w4855;
assign v2324 = ~(w4856 | w4857);
assign w4858 = v2324;
assign w4859 = w4849 & ~w4858;
assign w4860 = ~w4849 & w4858;
assign v2325 = ~(w4859 | w4860);
assign w4861 = v2325;
assign w4862 = w4835 & w4861;
assign v2326 = ~(w4835 | w4861);
assign w4863 = v2326;
assign v2327 = ~(w4862 | w4863);
assign w4864 = v2327;
assign w4865 = pi13 & pi36;
assign w4866 = pi08 & pi41;
assign w4867 = pi07 & pi42;
assign v2328 = ~(w4866 | w4867);
assign w4868 = v2328;
assign w4869 = pi08 & pi42;
assign w4870 = w4616 & w4869;
assign v2329 = ~(w4868 | w4870);
assign w4871 = v2329;
assign w4872 = w4865 & ~w4871;
assign w4873 = ~w4865 & w4871;
assign v2330 = ~(w4872 | w4873);
assign w4874 = v2330;
assign w4875 = pi24 & pi25;
assign w4876 = pi23 & pi26;
assign v2331 = ~(w4875 | w4876);
assign w4877 = v2331;
assign w4878 = w4875 & w4876;
assign v2332 = ~(w4877 | w4878);
assign w4879 = v2332;
assign w4880 = w4632 & ~w4879;
assign w4881 = ~w4632 & w4879;
assign v2333 = ~(w4880 | w4881);
assign w4882 = v2333;
assign v2334 = ~(w4874 | w4882);
assign w4883 = v2334;
assign w4884 = w4874 & w4882;
assign v2335 = ~(w4883 | w4884);
assign w4885 = v2335;
assign w4886 = pi15 & pi34;
assign w4887 = pi06 & pi43;
assign w4888 = pi14 & pi35;
assign v2336 = ~(w4887 | w4888);
assign w4889 = v2336;
assign w4890 = w4887 & w4888;
assign v2337 = ~(w4889 | w4890);
assign w4891 = v2337;
assign w4892 = w4886 & ~w4891;
assign w4893 = ~w4886 & w4891;
assign v2338 = ~(w4892 | w4893);
assign w4894 = v2338;
assign w4895 = w4885 & ~w4894;
assign w4896 = ~w4885 & w4894;
assign v2339 = ~(w4895 | w4896);
assign w4897 = v2339;
assign w4898 = w4864 & w4897;
assign v2340 = ~(w4864 | w4897);
assign w4899 = v2340;
assign v2341 = ~(w4898 | w4899);
assign w4900 = v2341;
assign w4901 = ~w4802 & w4900;
assign w4902 = w4802 & ~w4900;
assign v2342 = ~(w4901 | w4902);
assign w4903 = v2342;
assign w4904 = ~w4801 & w4903;
assign w4905 = w4801 & ~w4903;
assign v2343 = ~(w4904 | w4905);
assign w4906 = v2343;
assign w4907 = ~w4800 & w4906;
assign w4908 = w4800 & ~w4906;
assign v2344 = ~(w4907 | w4908);
assign w4909 = v2344;
assign v2345 = ~(w4665 | w4669);
assign w4910 = v2345;
assign v2346 = ~(w4668 | w4910);
assign w4911 = v2346;
assign v2347 = ~(w4607 | w4611);
assign w4912 = v2347;
assign v2348 = ~(w4610 | w4912);
assign w4913 = v2348;
assign w4914 = w4911 & w4913;
assign v2349 = ~(w4911 | w4913);
assign w4915 = v2349;
assign v2350 = ~(w4914 | w4915);
assign w4916 = v2350;
assign v2351 = ~(w4616 | w4620);
assign w4917 = v2351;
assign v2352 = ~(w4619 | w4917);
assign w4918 = v2352;
assign v2353 = ~(w4916 | w4918);
assign w4919 = v2353;
assign w4920 = w4916 & w4918;
assign v2354 = ~(w4919 | w4920);
assign w4921 = v2354;
assign w4922 = (~w4662 & ~w4664) | (~w4662 & w16881) | (~w4664 & w16881);
assign w4923 = ~w4921 & w4922;
assign w4924 = w4921 & ~w4922;
assign v2355 = ~(w4923 | w4924);
assign w4925 = v2355;
assign w4926 = (~w4769 & ~w4771) | (~w4769 & w16882) | (~w4771 & w16882);
assign w4927 = ~w4925 & w4926;
assign w4928 = w4925 & ~w4926;
assign v2356 = ~(w4927 | w4928);
assign w4929 = v2356;
assign v2357 = ~(w4641 | w4678);
assign w4930 = v2357;
assign w4931 = ~w4929 & w4930;
assign w4932 = w4929 & ~w4930;
assign v2358 = ~(w4931 | w4932);
assign w4933 = v2358;
assign v2359 = ~(w4644 | w4648);
assign w4934 = v2359;
assign v2360 = ~(w4647 | w4934);
assign w4935 = v2360;
assign v2361 = ~(w4712 | w4716);
assign w4936 = v2361;
assign v2362 = ~(w4715 | w4936);
assign w4937 = v2362;
assign w4938 = w4935 & w4937;
assign v2363 = ~(w4935 | w4937);
assign w4939 = v2363;
assign v2364 = ~(w4938 | w4939);
assign w4940 = v2364;
assign v2365 = ~(w4653 | w4657);
assign w4941 = v2365;
assign v2366 = ~(w4656 | w4941);
assign w4942 = v2366;
assign v2367 = ~(w4940 | w4942);
assign w4943 = v2367;
assign w4944 = w4940 & w4942;
assign v2368 = ~(w4943 | w4944);
assign w4945 = v2368;
assign w4946 = (~w4625 & ~w4627) | (~w4625 & w16883) | (~w4627 & w16883);
assign w4947 = ~pi48 & w4764;
assign w4948 = pi48 & w1296;
assign w4949 = pi01 & pi48;
assign v2369 = ~(pi25 | w4949);
assign w4950 = v2369;
assign v2370 = ~(w4948 | w4950);
assign w4951 = v2370;
assign v2371 = ~(w4764 | w4951);
assign w4952 = v2371;
assign v2372 = ~(w4947 | w4952);
assign w4953 = v2372;
assign w4954 = w4628 & ~w4631;
assign v2373 = ~(w4633 | w4954);
assign w4955 = v2373;
assign w4956 = w4953 & ~w4955;
assign w4957 = ~w4953 & w4955;
assign v2374 = ~(w4956 | w4957);
assign w4958 = v2374;
assign w4959 = ~w4946 & w4958;
assign w4960 = w4946 & ~w4958;
assign v2375 = ~(w4959 | w4960);
assign w4961 = v2375;
assign w4962 = w4945 & w4961;
assign v2376 = ~(w4945 | w4961);
assign w4963 = v2376;
assign v2377 = ~(w4962 | w4963);
assign w4964 = v2377;
assign w4965 = w4933 & w4964;
assign v2378 = ~(w4933 | w4964);
assign w4966 = v2378;
assign v2379 = ~(w4965 | w4966);
assign w4967 = v2379;
assign v2380 = ~(w4680 | w4683);
assign w4968 = v2380;
assign w4969 = (~w4735 & ~w4737) | (~w4735 & w17100) | (~w4737 & w17100);
assign w4970 = (~w4693 & ~w4695) | (~w4693 & w16736) | (~w4695 & w16736);
assign w4971 = (~w4709 & ~w4711) | (~w4709 & w16737) | (~w4711 & w16737);
assign v2381 = ~(w4970 | w4971);
assign w4972 = v2381;
assign w4973 = w4970 & w4971;
assign v2382 = ~(w4972 | w4973);
assign w4974 = v2382;
assign w4975 = w4969 & ~w4974;
assign w4976 = ~w4969 & w4974;
assign v2383 = ~(w4975 | w4976);
assign w4977 = v2383;
assign w4978 = (~w4703 & ~w4704) | (~w4703 & w17101) | (~w4704 & w17101);
assign w4979 = (~w4745 & ~w4747) | (~w4745 & w17102) | (~w4747 & w17102);
assign v2384 = ~(w4978 | w4979);
assign w4980 = v2384;
assign w4981 = w4978 & w4979;
assign v2385 = ~(w4980 | w4981);
assign w4982 = v2385;
assign v2386 = ~(w4977 | w4982);
assign w4983 = v2386;
assign w4984 = w4977 & w4982;
assign v2387 = ~(w4983 | w4984);
assign w4985 = v2387;
assign w4986 = ~w4968 & w4985;
assign w4987 = w4968 & ~w4985;
assign v2388 = ~(w4986 | w4987);
assign w4988 = v2388;
assign w4989 = w4967 & w4988;
assign v2389 = ~(w4967 | w4988);
assign w4990 = v2389;
assign v2390 = ~(w4989 | w4990);
assign w4991 = v2390;
assign w4992 = w4909 & w4991;
assign v2391 = ~(w4909 | w4991);
assign w4993 = v2391;
assign v2392 = ~(w4992 | w4993);
assign w4994 = v2392;
assign v2393 = ~(w4686 | w4789);
assign w4995 = v2393;
assign w4996 = ~w4994 & w4995;
assign w4997 = w4994 & ~w4995;
assign v2394 = ~(w4996 | w4997);
assign w4998 = v2394;
assign w4999 = w4799 & w4998;
assign v2395 = ~(w4799 | w4998);
assign w5000 = v2395;
assign v2396 = ~(w4999 | w5000);
assign w5001 = v2396;
assign v2397 = ~(w4792 | w4996);
assign w5002 = v2397;
assign w5003 = (w5002 & w4601) | (w5002 & w16528) | (w4601 & w16528);
assign v2398 = ~(w4997 | w5003);
assign w5004 = v2398;
assign v2399 = ~(w4907 | w4992);
assign w5005 = v2399;
assign v2400 = ~(w4986 | w4989);
assign w5006 = v2400;
assign v2401 = ~(w4932 | w4965);
assign w5007 = v2401;
assign v2402 = ~(w4980 | w4984);
assign w5008 = v2402;
assign w5009 = (~w4947 & ~w4953) | (~w4947 & w16884) | (~w4953 & w16884);
assign w5010 = pi22 & pi28;
assign w5011 = pi18 & pi32;
assign w5012 = pi23 & pi27;
assign v2403 = ~(w5011 | w5012);
assign w5013 = v2403;
assign w5014 = w5011 & w5012;
assign v2404 = ~(w5013 | w5014);
assign w5015 = v2404;
assign w5016 = w5010 & ~w5015;
assign w5017 = ~w5010 & w5015;
assign v2405 = ~(w5016 | w5017);
assign w5018 = v2405;
assign w5019 = pi16 & pi34;
assign w5020 = pi15 & pi35;
assign v2406 = ~(w4841 | w5020);
assign w5021 = v2406;
assign w5022 = w4841 & w5020;
assign v2407 = ~(w5021 | w5022);
assign w5023 = v2407;
assign w5024 = w5019 & ~w5023;
assign w5025 = ~w5019 & w5023;
assign v2408 = ~(w5024 | w5025);
assign w5026 = v2408;
assign v2409 = ~(w5018 | w5026);
assign w5027 = v2409;
assign w5028 = w5018 & w5026;
assign v2410 = ~(w5027 | w5028);
assign w5029 = v2410;
assign w5030 = w5009 & ~w5029;
assign w5031 = ~w5009 & w5029;
assign v2411 = ~(w5030 | w5031);
assign w5032 = v2411;
assign w5033 = pi04 & pi46;
assign w5034 = pi17 & pi33;
assign v2412 = ~(w5033 | w5034);
assign w5035 = v2412;
assign w5036 = w5033 & w5034;
assign v2413 = ~(w5035 | w5036);
assign w5037 = v2413;
assign w5038 = w4806 & ~w5037;
assign w5039 = ~w4806 & w5037;
assign v2414 = ~(w5038 | w5039);
assign w5040 = v2414;
assign w5041 = pi00 & pi50;
assign w5042 = pi02 & pi48;
assign v2415 = ~(w5041 | w5042);
assign w5043 = v2415;
assign w5044 = pi02 & pi50;
assign w5045 = w4757 & w5044;
assign v2416 = ~(w5043 | w5045);
assign w5046 = v2416;
assign w5047 = w4948 & ~w5046;
assign w5048 = ~w4948 & w5046;
assign v2417 = ~(w5047 | w5048);
assign w5049 = v2417;
assign v2418 = ~(w5040 | w5049);
assign w5050 = v2418;
assign w5051 = w5040 & w5049;
assign v2419 = ~(w5050 | w5051);
assign w5052 = v2419;
assign w5053 = pi19 & pi31;
assign w5054 = pi21 & pi29;
assign w5055 = pi20 & pi30;
assign v2420 = ~(w5054 | w5055);
assign w5056 = v2420;
assign w5057 = w5054 & w5055;
assign v2421 = ~(w5056 | w5057);
assign w5058 = v2421;
assign w5059 = w5053 & ~w5058;
assign w5060 = ~w5053 & w5058;
assign v2422 = ~(w5059 | w5060);
assign w5061 = v2422;
assign w5062 = w5052 & ~w5061;
assign w5063 = ~w5052 & w5061;
assign v2423 = ~(w5062 | w5063);
assign w5064 = v2423;
assign w5065 = pi06 & pi44;
assign w5066 = pi07 & pi43;
assign w5067 = pi14 & pi36;
assign v2424 = ~(w5066 | w5067);
assign w5068 = v2424;
assign w5069 = w5066 & w5067;
assign v2425 = ~(w5068 | w5069);
assign w5070 = v2425;
assign w5071 = w5065 & ~w5070;
assign w5072 = ~w5065 & w5070;
assign v2426 = ~(w5071 | w5072);
assign w5073 = v2426;
assign w5074 = pi13 & pi37;
assign w5075 = pi09 & pi41;
assign v2427 = ~(w5074 | w5075);
assign w5076 = v2427;
assign w5077 = w5074 & w5075;
assign v2428 = ~(w5076 | w5077);
assign w5078 = v2428;
assign w5079 = w4869 & ~w5078;
assign w5080 = ~w4869 & w5078;
assign v2429 = ~(w5079 | w5080);
assign w5081 = v2429;
assign v2430 = ~(w5073 | w5081);
assign w5082 = v2430;
assign w5083 = w5073 & w5081;
assign v2431 = ~(w5082 | w5083);
assign w5084 = v2431;
assign w5085 = pi12 & pi38;
assign w5086 = pi11 & pi39;
assign w5087 = pi10 & pi40;
assign v2432 = ~(w5086 | w5087);
assign w5088 = v2432;
assign w5089 = w5086 & w5087;
assign v2433 = ~(w5088 | w5089);
assign w5090 = v2433;
assign w5091 = w5085 & ~w5090;
assign w5092 = ~w5085 & w5090;
assign v2434 = ~(w5091 | w5092);
assign w5093 = v2434;
assign w5094 = w5084 & ~w5093;
assign w5095 = ~w5084 & w5093;
assign v2435 = ~(w5094 | w5095);
assign w5096 = v2435;
assign w5097 = w5064 & w5096;
assign v2436 = ~(w5064 | w5096);
assign w5098 = v2436;
assign v2437 = ~(w5097 | w5098);
assign w5099 = v2437;
assign v2438 = ~(w5032 | w5099);
assign w5100 = v2438;
assign w5101 = w5032 & w5099;
assign v2439 = ~(w5100 | w5101);
assign w5102 = v2439;
assign w5103 = ~w5008 & w5102;
assign w5104 = w5008 & ~w5102;
assign v2440 = ~(w5103 | w5104);
assign w5105 = v2440;
assign w5106 = ~w5007 & w5105;
assign w5107 = w5007 & ~w5105;
assign v2441 = ~(w5106 | w5107);
assign w5108 = v2441;
assign w5109 = ~w5006 & w5108;
assign w5110 = w5006 & ~w5108;
assign v2442 = ~(w5109 | w5110);
assign w5111 = v2442;
assign v2443 = ~(w4901 | w4904);
assign w5112 = v2443;
assign w5113 = w4837 & ~w4840;
assign v2444 = ~(w4842 | w5113);
assign w5114 = v2444;
assign w5115 = w4803 & ~w4805;
assign v2445 = ~(w4807 | w5115);
assign w5116 = v2445;
assign v2446 = ~(w5114 | w5116);
assign w5117 = v2446;
assign w5118 = w5114 & w5116;
assign v2447 = ~(w5117 | w5118);
assign w5119 = v2447;
assign v2448 = ~(w4886 | w4890);
assign w5120 = v2448;
assign v2449 = ~(w4889 | w5120);
assign w5121 = v2449;
assign v2450 = ~(w5119 | w5121);
assign w5122 = v2450;
assign w5123 = w5119 & w5121;
assign v2451 = ~(w5122 | w5123);
assign w5124 = v2451;
assign w5125 = (~w4914 & ~w4916) | (~w4914 & w16738) | (~w4916 & w16738);
assign w5126 = (~w4938 & ~w4940) | (~w4938 & w16739) | (~w4940 & w16739);
assign v2452 = ~(w5125 | w5126);
assign w5127 = v2452;
assign w5128 = w5125 & w5126;
assign v2453 = ~(w5127 | w5128);
assign w5129 = v2453;
assign w5130 = w5124 & w5129;
assign v2454 = ~(w5124 | w5129);
assign w5131 = v2454;
assign v2455 = ~(w5130 | w5131);
assign w5132 = v2455;
assign v2456 = ~(w4924 | w4928);
assign w5133 = v2456;
assign w5134 = (~w4959 & ~w4961) | (~w4959 & w17103) | (~w4961 & w17103);
assign v2457 = ~(w5133 | w5134);
assign w5135 = v2457;
assign w5136 = w5133 & w5134;
assign v2458 = ~(w5135 | w5136);
assign w5137 = v2458;
assign w5138 = w5132 & w5137;
assign v2459 = ~(w5132 | w5137);
assign w5139 = v2459;
assign v2460 = ~(w5138 | w5139);
assign w5140 = v2460;
assign w5141 = ~w5112 & w5140;
assign w5142 = w5112 & ~w5140;
assign v2461 = ~(w5141 | w5142);
assign w5143 = v2461;
assign w5144 = pi24 & pi26;
assign w5145 = pi01 & pi49;
assign v2462 = ~(w5144 | w5145);
assign w5146 = v2462;
assign w5147 = w5144 & w5145;
assign v2463 = ~(w5146 | w5147);
assign w5148 = v2463;
assign v2464 = ~(w4632 | w4878);
assign w5149 = v2464;
assign v2465 = ~(w4877 | w5149);
assign w5150 = v2465;
assign w5151 = w5148 & w5150;
assign v2466 = ~(w5148 | w5150);
assign w5152 = v2466;
assign v2467 = ~(w5151 | w5152);
assign w5153 = v2467;
assign v2468 = ~(w4824 | w4828);
assign w5154 = v2468;
assign v2469 = ~(w4827 | w5154);
assign w5155 = v2469;
assign w5156 = w5153 & w5155;
assign v2470 = ~(w5153 | w5155);
assign w5157 = v2470;
assign v2471 = ~(w5156 | w5157);
assign w5158 = v2471;
assign w5159 = (~w4821 & ~w4823) | (~w4821 & w16885) | (~w4823 & w16885);
assign w5160 = (~w4847 & ~w4849) | (~w4847 & w16886) | (~w4849 & w16886);
assign v2472 = ~(w5159 | w5160);
assign w5161 = v2472;
assign w5162 = w5159 & w5160;
assign v2473 = ~(w5161 | w5162);
assign w5163 = v2473;
assign w5164 = w5158 & w5163;
assign v2474 = ~(w5158 | w5163);
assign w5165 = v2474;
assign v2475 = ~(w5164 | w5165);
assign w5166 = v2475;
assign v2476 = ~(w4812 | w4816);
assign w5167 = v2476;
assign v2477 = ~(w4815 | w5167);
assign w5168 = v2477;
assign v2478 = ~(w4850 | w4854);
assign w5169 = v2478;
assign v2479 = ~(w4853 | w5169);
assign w5170 = v2479;
assign w5171 = w5168 & w5170;
assign v2480 = ~(w5168 | w5170);
assign w5172 = v2480;
assign v2481 = ~(w5171 | w5172);
assign w5173 = v2481;
assign w5174 = w4865 & ~w4868;
assign v2482 = ~(w4870 | w5174);
assign w5175 = v2482;
assign w5176 = ~w5173 & w5175;
assign w5177 = w5173 & ~w5175;
assign v2483 = ~(w5176 | w5177);
assign w5178 = v2483;
assign w5179 = (~w4883 & ~w4885) | (~w4883 & w16887) | (~w4885 & w16887);
assign w5180 = ~w5178 & w5179;
assign w5181 = w5178 & ~w5179;
assign v2484 = ~(w5180 | w5181);
assign w5182 = v2484;
assign w5183 = (~w4972 & ~w4974) | (~w4972 & w16888) | (~w4974 & w16888);
assign w5184 = ~w5182 & w5183;
assign w5185 = w5182 & ~w5183;
assign v2485 = ~(w5184 | w5185);
assign w5186 = v2485;
assign v2486 = ~(w4862 | w4898);
assign w5187 = v2486;
assign w5188 = ~w5186 & w5187;
assign w5189 = w5186 & ~w5187;
assign v2487 = ~(w5188 | w5189);
assign w5190 = v2487;
assign w5191 = w5166 & w5190;
assign v2488 = ~(w5166 | w5190);
assign w5192 = v2488;
assign v2489 = ~(w5191 | w5192);
assign w5193 = v2489;
assign w5194 = w5143 & w5193;
assign v2490 = ~(w5143 | w5193);
assign w5195 = v2490;
assign v2491 = ~(w5194 | w5195);
assign w5196 = v2491;
assign w5197 = w5111 & w5196;
assign v2492 = ~(w5111 | w5196);
assign w5198 = v2492;
assign v2493 = ~(w5197 | w5198);
assign w5199 = v2493;
assign w5200 = ~w5005 & w5199;
assign w5201 = w5005 & ~w5199;
assign v2494 = ~(w5200 | w5201);
assign w5202 = v2494;
assign w5203 = w5004 & w5202;
assign v2495 = ~(w5004 | w5202);
assign w5204 = v2495;
assign v2496 = ~(w5203 | w5204);
assign w5205 = v2496;
assign v2497 = ~(w4997 | w5200);
assign w5206 = v2497;
assign w5207 = (w4601 & w16530) | (w4601 & w16531) | (w16530 & w16531);
assign v2498 = ~(w5109 | w5197);
assign w5208 = v2498;
assign v2499 = ~(w5141 | w5194);
assign w5209 = v2499;
assign v2500 = ~(w5189 | w5191);
assign w5210 = v2500;
assign w5211 = (~w5135 & ~w5137) | (~w5135 & w17104) | (~w5137 & w17104);
assign w5212 = (~w5171 & ~w5173) | (~w5171 & w17105) | (~w5173 & w17105);
assign w5213 = pi00 & pi51;
assign w5214 = w5147 & w5213;
assign v2501 = ~(w5147 | w5213);
assign w5215 = v2501;
assign v2502 = ~(w5214 | w5215);
assign w5216 = v2502;
assign w5217 = pi01 & pi50;
assign w5218 = pi26 & w5217;
assign v2503 = ~(pi26 | w5217);
assign w5219 = v2503;
assign v2504 = ~(w5218 | w5219);
assign w5220 = v2504;
assign w5221 = w5216 & w5220;
assign v2505 = ~(w5216 | w5220);
assign w5222 = v2505;
assign v2506 = ~(w5221 | w5222);
assign w5223 = v2506;
assign w5224 = pi17 & pi34;
assign w5225 = pi20 & pi31;
assign w5226 = pi19 & pi32;
assign v2507 = ~(w5225 | w5226);
assign w5227 = v2507;
assign w5228 = w5225 & w5226;
assign v2508 = ~(w5227 | w5228);
assign w5229 = v2508;
assign w5230 = w5224 & ~w5229;
assign w5231 = ~w5224 & w5229;
assign v2509 = ~(w5230 | w5231);
assign w5232 = v2509;
assign w5233 = w5223 & ~w5232;
assign w5234 = ~w5223 & w5232;
assign v2510 = ~(w5233 | w5234);
assign w5235 = v2510;
assign w5236 = w5212 & ~w5235;
assign w5237 = ~w5212 & w5235;
assign v2511 = ~(w5236 | w5237);
assign w5238 = v2511;
assign w5239 = pi18 & pi33;
assign w5240 = pi05 & pi46;
assign w5241 = pi16 & pi35;
assign v2512 = ~(w5240 | w5241);
assign w5242 = v2512;
assign w5243 = w5240 & w5241;
assign v2513 = ~(w5242 | w5243);
assign w5244 = v2513;
assign w5245 = w5239 & ~w5244;
assign w5246 = ~w5239 & w5244;
assign v2514 = ~(w5245 | w5246);
assign w5247 = v2514;
assign w5248 = pi21 & pi30;
assign w5249 = pi22 & pi29;
assign w5250 = pi23 & pi28;
assign v2515 = ~(w5249 | w5250);
assign w5251 = v2515;
assign w5252 = w5249 & w5250;
assign v2516 = ~(w5251 | w5252);
assign w5253 = v2516;
assign w5254 = w5248 & ~w5253;
assign w5255 = ~w5248 & w5253;
assign v2517 = ~(w5254 | w5255);
assign w5256 = v2517;
assign v2518 = ~(w5247 | w5256);
assign w5257 = v2518;
assign w5258 = w5247 & w5256;
assign v2519 = ~(w5257 | w5258);
assign w5259 = v2519;
assign w5260 = pi15 & pi36;
assign w5261 = pi06 & pi45;
assign w5262 = pi14 & pi37;
assign v2520 = ~(w5261 | w5262);
assign w5263 = v2520;
assign w5264 = w5261 & w5262;
assign v2521 = ~(w5263 | w5264);
assign w5265 = v2521;
assign w5266 = w5260 & ~w5265;
assign w5267 = ~w5260 & w5265;
assign v2522 = ~(w5266 | w5267);
assign w5268 = v2522;
assign w5269 = w5259 & ~w5268;
assign w5270 = ~w5259 & w5268;
assign v2523 = ~(w5269 | w5270);
assign w5271 = v2523;
assign w5272 = pi07 & pi44;
assign w5273 = pi13 & pi38;
assign w5274 = pi08 & pi43;
assign v2524 = ~(w5273 | w5274);
assign w5275 = v2524;
assign w5276 = w5273 & w5274;
assign v2525 = ~(w5275 | w5276);
assign w5277 = v2525;
assign w5278 = w5272 & ~w5277;
assign w5279 = ~w5272 & w5277;
assign v2526 = ~(w5278 | w5279);
assign w5280 = v2526;
assign w5281 = pi09 & pi42;
assign w5282 = pi12 & pi39;
assign w5283 = pi10 & pi41;
assign v2527 = ~(w5282 | w5283);
assign w5284 = v2527;
assign w5285 = w5282 & w5283;
assign v2528 = ~(w5284 | w5285);
assign w5286 = v2528;
assign w5287 = w5281 & ~w5286;
assign w5288 = ~w5281 & w5286;
assign v2529 = ~(w5287 | w5288);
assign w5289 = v2529;
assign v2530 = ~(w5280 | w5289);
assign w5290 = v2530;
assign w5291 = w5280 & w5289;
assign v2531 = ~(w5290 | w5291);
assign w5292 = v2531;
assign w5293 = pi11 & pi40;
assign w5294 = pi25 & pi26;
assign w5295 = pi24 & pi27;
assign v2532 = ~(w5294 | w5295);
assign w5296 = v2532;
assign w5297 = w5294 & w5295;
assign v2533 = ~(w5296 | w5297);
assign w5298 = v2533;
assign w5299 = w5293 & ~w5298;
assign w5300 = ~w5293 & w5298;
assign v2534 = ~(w5299 | w5300);
assign w5301 = v2534;
assign w5302 = w5292 & ~w5301;
assign w5303 = ~w5292 & w5301;
assign v2535 = ~(w5302 | w5303);
assign w5304 = v2535;
assign w5305 = w5271 & w5304;
assign v2536 = ~(w5271 | w5304);
assign w5306 = v2536;
assign v2537 = ~(w5305 | w5306);
assign w5307 = v2537;
assign v2538 = ~(w5238 | w5307);
assign w5308 = v2538;
assign w5309 = w5238 & w5307;
assign v2539 = ~(w5308 | w5309);
assign w5310 = v2539;
assign w5311 = ~w5211 & w5310;
assign w5312 = w5211 & ~w5310;
assign v2540 = ~(w5311 | w5312);
assign w5313 = v2540;
assign w5314 = ~w5210 & w5313;
assign w5315 = w5210 & ~w5313;
assign v2541 = ~(w5314 | w5315);
assign w5316 = v2541;
assign w5317 = ~w5209 & w5316;
assign w5318 = w5209 & ~w5316;
assign v2542 = ~(w5317 | w5318);
assign w5319 = v2542;
assign v2543 = ~(w5103 | w5106);
assign w5320 = v2543;
assign v2544 = ~(w5050 | w5062);
assign w5321 = v2544;
assign w5322 = (~w5117 & ~w5119) | (~w5117 & w17106) | (~w5119 & w17106);
assign w5323 = (~w5151 & ~w5153) | (~w5151 & w17107) | (~w5153 & w17107);
assign v2545 = ~(w5322 | w5323);
assign w5324 = v2545;
assign w5325 = w5322 & w5323;
assign v2546 = ~(w5324 | w5325);
assign w5326 = v2546;
assign w5327 = w5321 & ~w5326;
assign w5328 = ~w5321 & w5326;
assign v2547 = ~(w5327 | w5328);
assign w5329 = v2547;
assign v2548 = ~(w5181 | w5185);
assign w5330 = v2548;
assign w5331 = (~w5161 & ~w5163) | (~w5161 & w17108) | (~w5163 & w17108);
assign v2549 = ~(w5330 | w5331);
assign w5332 = v2549;
assign w5333 = w5330 & w5331;
assign v2550 = ~(w5332 | w5333);
assign w5334 = v2550;
assign w5335 = w5329 & w5334;
assign v2551 = ~(w5329 | w5334);
assign w5336 = v2551;
assign v2552 = ~(w5335 | w5336);
assign w5337 = v2552;
assign w5338 = ~w5320 & w5337;
assign w5339 = w5320 & ~w5337;
assign v2553 = ~(w5338 | w5339);
assign w5340 = v2553;
assign v2554 = ~(w5097 | w5101);
assign w5341 = v2554;
assign w5342 = (~w5127 & ~w5129) | (~w5127 & w16889) | (~w5129 & w16889);
assign v2555 = ~(w5019 | w5022);
assign w5343 = v2555;
assign v2556 = ~(w5021 | w5343);
assign w5344 = v2556;
assign v2557 = ~(w5085 | w5089);
assign w5345 = v2557;
assign v2558 = ~(w5088 | w5345);
assign w5346 = v2558;
assign w5347 = w5344 & w5346;
assign v2559 = ~(w5344 | w5346);
assign w5348 = v2559;
assign v2560 = ~(w5347 | w5348);
assign w5349 = v2560;
assign w5350 = pi02 & pi49;
assign w5351 = pi03 & pi48;
assign w5352 = pi04 & pi47;
assign v2561 = ~(w5351 | w5352);
assign w5353 = v2561;
assign w5354 = pi04 & pi48;
assign w5355 = w4806 & w5354;
assign v2562 = ~(w5353 | w5355);
assign w5356 = v2562;
assign w5357 = w5350 & ~w5356;
assign w5358 = ~w5350 & w5356;
assign v2563 = ~(w5357 | w5358);
assign w5359 = v2563;
assign w5360 = ~w5349 & w5359;
assign w5361 = w5349 & ~w5359;
assign v2564 = ~(w5360 | w5361);
assign w5362 = v2564;
assign w5363 = (~w5027 & ~w5029) | (~w5027 & w16890) | (~w5029 & w16890);
assign w5364 = w5362 & ~w5363;
assign w5365 = ~w5362 & w5363;
assign v2565 = ~(w5364 | w5365);
assign w5366 = v2565;
assign w5367 = ~w5342 & w5366;
assign w5368 = w5342 & ~w5366;
assign v2566 = ~(w5367 | w5368);
assign w5369 = v2566;
assign w5370 = ~w5341 & w5369;
assign w5371 = w5341 & ~w5369;
assign v2567 = ~(w5370 | w5371);
assign w5372 = v2567;
assign v2568 = ~(w4869 | w5077);
assign w5373 = v2568;
assign v2569 = ~(w5076 | w5373);
assign w5374 = v2569;
assign v2570 = ~(w5065 | w5069);
assign w5375 = v2570;
assign v2571 = ~(w5068 | w5375);
assign w5376 = v2571;
assign w5377 = w5374 & w5376;
assign v2572 = ~(w5374 | w5376);
assign w5378 = v2572;
assign v2573 = ~(w5377 | w5378);
assign w5379 = v2573;
assign v2574 = ~(w5010 | w5014);
assign w5380 = v2574;
assign v2575 = ~(w5013 | w5380);
assign w5381 = v2575;
assign v2576 = ~(w5379 | w5381);
assign w5382 = v2576;
assign w5383 = w5379 & w5381;
assign v2577 = ~(w5382 | w5383);
assign w5384 = v2577;
assign v2578 = ~(w5082 | w5094);
assign w5385 = v2578;
assign w5386 = ~w5384 & w5385;
assign w5387 = w5384 & ~w5385;
assign v2579 = ~(w5386 | w5387);
assign w5388 = v2579;
assign v2580 = ~(w4806 | w5036);
assign w5389 = v2580;
assign v2581 = ~(w5035 | w5389);
assign w5390 = v2581;
assign v2582 = ~(w5053 | w5057);
assign w5391 = v2582;
assign v2583 = ~(w5056 | w5391);
assign w5392 = v2583;
assign w5393 = w5390 & w5392;
assign v2584 = ~(w5390 | w5392);
assign w5394 = v2584;
assign v2585 = ~(w5393 | w5394);
assign w5395 = v2585;
assign v2586 = ~(w4948 | w5045);
assign w5396 = v2586;
assign v2587 = ~(w5043 | w5396);
assign w5397 = v2587;
assign v2588 = ~(w5395 | w5397);
assign w5398 = v2588;
assign w5399 = w5395 & w5397;
assign v2589 = ~(w5398 | w5399);
assign w5400 = v2589;
assign w5401 = w5388 & w5400;
assign v2590 = ~(w5388 | w5400);
assign w5402 = v2590;
assign v2591 = ~(w5401 | w5402);
assign w5403 = v2591;
assign w5404 = w5372 & w5403;
assign v2592 = ~(w5372 | w5403);
assign w5405 = v2592;
assign v2593 = ~(w5404 | w5405);
assign w5406 = v2593;
assign w5407 = w5340 & w5406;
assign v2594 = ~(w5340 | w5406);
assign w5408 = v2594;
assign v2595 = ~(w5407 | w5408);
assign w5409 = v2595;
assign w5410 = w5319 & w5409;
assign v2596 = ~(w5319 | w5409);
assign w5411 = v2596;
assign v2597 = ~(w5410 | w5411);
assign w5412 = v2597;
assign w5413 = ~w5208 & w5412;
assign w5414 = w5208 & ~w5412;
assign v2598 = ~(w5413 | w5414);
assign w5415 = v2598;
assign v2599 = ~(w5207 | w5415);
assign w5416 = v2599;
assign w5417 = w5207 & w5415;
assign v2600 = ~(w5416 | w5417);
assign w5418 = v2600;
assign v2601 = ~(w5317 | w5410);
assign w5419 = v2601;
assign v2602 = ~(w5311 | w5314);
assign w5420 = v2602;
assign w5421 = (~w5377 & ~w5379) | (~w5377 & w17109) | (~w5379 & w17109);
assign w5422 = (~w5393 & ~w5395) | (~w5393 & w16740) | (~w5395 & w16740);
assign w5423 = pi19 & pi33;
assign w5424 = pi03 & pi49;
assign v2603 = ~(w5044 | w5424);
assign w5425 = v2603;
assign w5426 = pi03 & pi50;
assign w5427 = w5350 & w5426;
assign v2604 = ~(w5425 | w5427);
assign w5428 = v2604;
assign w5429 = w5423 & ~w5428;
assign w5430 = ~w5423 & w5428;
assign v2605 = ~(w5429 | w5430);
assign w5431 = v2605;
assign v2606 = ~(w5422 | w5431);
assign w5432 = v2606;
assign w5433 = w5422 & w5431;
assign v2607 = ~(w5432 | w5433);
assign w5434 = v2607;
assign w5435 = w5421 & ~w5434;
assign w5436 = ~w5421 & w5434;
assign v2608 = ~(w5435 | w5436);
assign w5437 = v2608;
assign v2609 = ~(w5364 | w5367);
assign w5438 = v2609;
assign w5439 = ~w5437 & w5438;
assign w5440 = w5437 & ~w5438;
assign v2610 = ~(w5439 | w5440);
assign w5441 = v2610;
assign v2611 = ~(w5290 | w5302);
assign w5442 = v2611;
assign w5443 = (~w5347 & ~w5349) | (~w5347 & w17110) | (~w5349 & w17110);
assign w5444 = pi25 & pi27;
assign w5445 = pi01 & pi51;
assign v2612 = ~(w5444 | w5445);
assign w5446 = v2612;
assign w5447 = w5444 & w5445;
assign v2613 = ~(w5446 | w5447);
assign w5448 = v2613;
assign w5449 = w5218 & w5448;
assign v2614 = ~(w5218 | w5448);
assign w5450 = v2614;
assign v2615 = ~(w5449 | w5450);
assign w5451 = v2615;
assign v2616 = ~(w5293 | w5297);
assign w5452 = v2616;
assign v2617 = ~(w5296 | w5452);
assign w5453 = v2617;
assign w5454 = w5451 & w5453;
assign v2618 = ~(w5451 | w5453);
assign w5455 = v2618;
assign v2619 = ~(w5454 | w5455);
assign w5456 = v2619;
assign w5457 = ~w5443 & w5456;
assign w5458 = w5443 & ~w5456;
assign v2620 = ~(w5457 | w5458);
assign w5459 = v2620;
assign w5460 = ~w5442 & w5459;
assign w5461 = w5442 & ~w5459;
assign v2621 = ~(w5460 | w5461);
assign w5462 = v2621;
assign w5463 = w5441 & w5462;
assign v2622 = ~(w5441 | w5462);
assign w5464 = v2622;
assign v2623 = ~(w5463 | w5464);
assign w5465 = v2623;
assign w5466 = ~w5420 & w5465;
assign w5467 = w5420 & ~w5465;
assign v2624 = ~(w5466 | w5467);
assign w5468 = v2624;
assign v2625 = ~(w5324 | w5328);
assign w5469 = v2625;
assign w5470 = (~w5214 & ~w5216) | (~w5214 & w16741) | (~w5216 & w16741);
assign v2626 = ~(w5281 | w5285);
assign w5471 = v2626;
assign v2627 = ~(w5284 | w5471);
assign w5472 = v2627;
assign w5473 = ~w5470 & w5472;
assign w5474 = w5470 & ~w5472;
assign v2628 = ~(w5473 | w5474);
assign w5475 = v2628;
assign w5476 = pi00 & pi52;
assign w5477 = pi17 & pi35;
assign v2629 = ~(w5354 | w5477);
assign w5478 = v2629;
assign w5479 = w5354 & w5477;
assign v2630 = ~(w5478 | w5479);
assign w5480 = v2630;
assign w5481 = w5476 & ~w5480;
assign w5482 = ~w5476 & w5480;
assign v2631 = ~(w5481 | w5482);
assign w5483 = v2631;
assign w5484 = ~w5475 & w5483;
assign w5485 = w5475 & ~w5483;
assign v2632 = ~(w5484 | w5485);
assign w5486 = v2632;
assign w5487 = (~w5233 & ~w5235) | (~w5233 & w17111) | (~w5235 & w17111);
assign w5488 = w5486 & ~w5487;
assign w5489 = ~w5486 & w5487;
assign v2633 = ~(w5488 | w5489);
assign w5490 = v2633;
assign w5491 = w5469 & ~w5490;
assign w5492 = ~w5469 & w5490;
assign v2634 = ~(w5491 | w5492);
assign w5493 = v2634;
assign v2635 = ~(w5305 | w5309);
assign w5494 = v2635;
assign v2636 = ~(w5272 | w5276);
assign w5495 = v2636;
assign v2637 = ~(w5275 | w5495);
assign w5496 = v2637;
assign v2638 = ~(w5239 | w5243);
assign w5497 = v2638;
assign v2639 = ~(w5242 | w5497);
assign w5498 = v2639;
assign w5499 = w5496 & w5498;
assign v2640 = ~(w5496 | w5498);
assign w5500 = v2640;
assign v2641 = ~(w5499 | w5500);
assign w5501 = v2641;
assign v2642 = ~(w5248 | w5252);
assign w5502 = v2642;
assign v2643 = ~(w5251 | w5502);
assign w5503 = v2643;
assign v2644 = ~(w5501 | w5503);
assign w5504 = v2644;
assign w5505 = w5501 & w5503;
assign v2645 = ~(w5504 | w5505);
assign w5506 = v2645;
assign v2646 = ~(w5224 | w5228);
assign w5507 = v2646;
assign v2647 = ~(w5227 | w5507);
assign w5508 = v2647;
assign w5509 = w5350 & ~w5353;
assign v2648 = ~(w5355 | w5509);
assign w5510 = v2648;
assign w5511 = w5508 & ~w5510;
assign w5512 = ~w5508 & w5510;
assign v2649 = ~(w5511 | w5512);
assign w5513 = v2649;
assign v2650 = ~(w5260 | w5264);
assign w5514 = v2650;
assign v2651 = ~(w5263 | w5514);
assign w5515 = v2651;
assign v2652 = ~(w5513 | w5515);
assign w5516 = v2652;
assign w5517 = w5513 & w5515;
assign v2653 = ~(w5516 | w5517);
assign w5518 = v2653;
assign v2654 = ~(w5257 | w5269);
assign w5519 = v2654;
assign w5520 = ~w5518 & w5519;
assign w5521 = w5518 & ~w5519;
assign v2655 = ~(w5520 | w5521);
assign w5522 = v2655;
assign w5523 = w5506 & w5522;
assign v2656 = ~(w5506 | w5522);
assign w5524 = v2656;
assign v2657 = ~(w5523 | w5524);
assign w5525 = v2657;
assign w5526 = ~w5494 & w5525;
assign w5527 = w5494 & ~w5525;
assign v2658 = ~(w5526 | w5527);
assign w5528 = v2658;
assign v2659 = ~(w5493 | w5528);
assign w5529 = v2659;
assign w5530 = w5493 & w5528;
assign v2660 = ~(w5529 | w5530);
assign w5531 = v2660;
assign v2661 = ~(w5468 | w5531);
assign w5532 = v2661;
assign w5533 = w5468 & w5531;
assign v2662 = ~(w5532 | w5533);
assign w5534 = v2662;
assign v2663 = ~(w5370 | w5404);
assign w5535 = v2663;
assign w5536 = (~w5332 & ~w5334) | (~w5332 & w17112) | (~w5334 & w17112);
assign v2664 = ~(w5387 | w5401);
assign w5537 = v2664;
assign w5538 = pi10 & pi42;
assign w5539 = pi12 & pi40;
assign w5540 = pi11 & pi41;
assign v2665 = ~(w5539 | w5540);
assign w5541 = v2665;
assign w5542 = pi12 & pi41;
assign w5543 = w5293 & w5542;
assign v2666 = ~(w5541 | w5543);
assign w5544 = v2666;
assign w5545 = w5538 & ~w5544;
assign w5546 = ~w5538 & w5544;
assign v2667 = ~(w5545 | w5546);
assign w5547 = v2667;
assign w5548 = pi05 & pi47;
assign w5549 = pi16 & pi36;
assign w5550 = pi06 & pi46;
assign v2668 = ~(w5549 | w5550);
assign w5551 = v2668;
assign w5552 = w5549 & w5550;
assign v2669 = ~(w5551 | w5552);
assign w5553 = v2669;
assign w5554 = w5548 & ~w5553;
assign w5555 = ~w5548 & w5553;
assign v2670 = ~(w5554 | w5555);
assign w5556 = v2670;
assign v2671 = ~(w5547 | w5556);
assign w5557 = v2671;
assign w5558 = w5547 & w5556;
assign v2672 = ~(w5557 | w5558);
assign w5559 = v2672;
assign w5560 = pi15 & pi37;
assign w5561 = pi08 & pi44;
assign w5562 = pi07 & pi45;
assign v2673 = ~(w5561 | w5562);
assign w5563 = v2673;
assign w5564 = pi08 & pi45;
assign w5565 = w5272 & w5564;
assign v2674 = ~(w5563 | w5565);
assign w5566 = v2674;
assign w5567 = w5560 & ~w5566;
assign w5568 = ~w5560 & w5566;
assign v2675 = ~(w5567 | w5568);
assign w5569 = v2675;
assign w5570 = w5559 & ~w5569;
assign w5571 = ~w5559 & w5569;
assign v2676 = ~(w5570 | w5571);
assign w5572 = v2676;
assign w5573 = pi18 & pi34;
assign w5574 = pi20 & pi32;
assign w5575 = pi21 & pi31;
assign v2677 = ~(w5574 | w5575);
assign w5576 = v2677;
assign w5577 = w5574 & w5575;
assign v2678 = ~(w5576 | w5577);
assign w5578 = v2678;
assign w5579 = w5573 & ~w5578;
assign w5580 = ~w5573 & w5578;
assign v2679 = ~(w5579 | w5580);
assign w5581 = v2679;
assign w5582 = pi22 & pi30;
assign w5583 = pi23 & pi29;
assign w5584 = pi24 & pi28;
assign v2680 = ~(w5583 | w5584);
assign w5585 = v2680;
assign w5586 = w5583 & w5584;
assign v2681 = ~(w5585 | w5586);
assign w5587 = v2681;
assign w5588 = w5582 & ~w5587;
assign w5589 = ~w5582 & w5587;
assign v2682 = ~(w5588 | w5589);
assign w5590 = v2682;
assign v2683 = ~(w5581 | w5590);
assign w5591 = v2683;
assign w5592 = w5581 & w5590;
assign v2684 = ~(w5591 | w5592);
assign w5593 = v2684;
assign w5594 = pi14 & pi38;
assign w5595 = pi09 & pi43;
assign w5596 = pi13 & pi39;
assign v2685 = ~(w5595 | w5596);
assign w5597 = v2685;
assign w5598 = w5595 & w5596;
assign v2686 = ~(w5597 | w5598);
assign w5599 = v2686;
assign w5600 = w5594 & ~w5599;
assign w5601 = ~w5594 & w5599;
assign v2687 = ~(w5600 | w5601);
assign w5602 = v2687;
assign w5603 = w5593 & ~w5602;
assign w5604 = ~w5593 & w5602;
assign v2688 = ~(w5603 | w5604);
assign w5605 = v2688;
assign w5606 = w5572 & w5605;
assign v2689 = ~(w5572 | w5605);
assign w5607 = v2689;
assign v2690 = ~(w5606 | w5607);
assign w5608 = v2690;
assign w5609 = ~w5537 & w5608;
assign w5610 = w5537 & ~w5608;
assign v2691 = ~(w5609 | w5610);
assign w5611 = v2691;
assign w5612 = ~w5536 & w5611;
assign w5613 = w5536 & ~w5611;
assign v2692 = ~(w5612 | w5613);
assign w5614 = v2692;
assign w5615 = w5535 & ~w5614;
assign w5616 = ~w5535 & w5614;
assign v2693 = ~(w5615 | w5616);
assign w5617 = v2693;
assign v2694 = ~(w5338 | w5407);
assign w5618 = v2694;
assign w5619 = ~w5617 & w5618;
assign w5620 = w5617 & ~w5618;
assign v2695 = ~(w5619 | w5620);
assign w5621 = v2695;
assign w5622 = w5534 & w5621;
assign v2696 = ~(w5534 | w5621);
assign w5623 = v2696;
assign v2697 = ~(w5622 | w5623);
assign w5624 = v2697;
assign w5625 = ~w5419 & w5624;
assign w5626 = w5419 & ~w5624;
assign v2698 = ~(w5414 | w5626);
assign w5627 = v2698;
assign w5628 = (w5627 & w5207) | (w5627 & w16532) | (w5207 & w16532);
assign w5629 = ~w5625 & w5628;
assign v2699 = ~(w5625 | w5626);
assign w5630 = v2699;
assign w5631 = w5207 & ~w5414;
assign v2700 = ~(w5413 | w5630);
assign w5632 = v2700;
assign w5633 = ~w5631 & w5632;
assign v2701 = ~(w5629 | w5633);
assign w5634 = v2701;
assign v2702 = ~(w5625 | w5628);
assign w5635 = v2702;
assign v2703 = ~(w5620 | w5622);
assign w5636 = v2703;
assign v2704 = ~(w5466 | w5533);
assign w5637 = v2704;
assign v2705 = ~(w5526 | w5530);
assign w5638 = v2705;
assign w5639 = (~w5432 & ~w5434) | (~w5432 & w16891) | (~w5434 & w16891);
assign w5640 = pi02 & pi51;
assign v2706 = ~(w5426 | w5640);
assign w5641 = v2706;
assign w5642 = pi03 & pi51;
assign w5643 = w5044 & w5642;
assign v2707 = ~(w5641 | w5643);
assign w5644 = v2707;
assign w5645 = w5447 & ~w5644;
assign w5646 = ~w5447 & w5644;
assign v2708 = ~(w5645 | w5646);
assign w5647 = v2708;
assign w5648 = pi04 & pi49;
assign w5649 = pi17 & pi36;
assign w5650 = pi18 & pi35;
assign v2709 = ~(w5649 | w5650);
assign w5651 = v2709;
assign w5652 = w5649 & w5650;
assign v2710 = ~(w5651 | w5652);
assign w5653 = v2710;
assign w5654 = w5648 & ~w5653;
assign w5655 = ~w5648 & w5653;
assign v2711 = ~(w5654 | w5655);
assign w5656 = v2711;
assign v2712 = ~(w5647 | w5656);
assign w5657 = v2712;
assign w5658 = w5647 & w5656;
assign v2713 = ~(w5657 | w5658);
assign w5659 = v2713;
assign w5660 = pi19 & pi34;
assign w5661 = pi21 & pi32;
assign w5662 = pi20 & pi33;
assign v2714 = ~(w5661 | w5662);
assign w5663 = v2714;
assign w5664 = w5661 & w5662;
assign v2715 = ~(w5663 | w5664);
assign w5665 = v2715;
assign w5666 = w5660 & ~w5665;
assign w5667 = ~w5660 & w5665;
assign v2716 = ~(w5666 | w5667);
assign w5668 = v2716;
assign w5669 = w5659 & ~w5668;
assign w5670 = ~w5659 & w5668;
assign v2717 = ~(w5669 | w5670);
assign w5671 = v2717;
assign w5672 = ~w5639 & w5671;
assign w5673 = w5639 & ~w5671;
assign v2718 = ~(w5672 | w5673);
assign w5674 = v2718;
assign w5675 = pi06 & pi47;
assign w5676 = pi07 & pi46;
assign w5677 = pi15 & pi38;
assign v2719 = ~(w5676 | w5677);
assign w5678 = v2719;
assign w5679 = w5676 & w5677;
assign v2720 = ~(w5678 | w5679);
assign w5680 = v2720;
assign w5681 = w5675 & ~w5680;
assign w5682 = ~w5675 & w5680;
assign v2721 = ~(w5681 | w5682);
assign w5683 = v2721;
assign w5684 = pi14 & pi39;
assign w5685 = pi09 & pi44;
assign v2722 = ~(w5684 | w5685);
assign w5686 = v2722;
assign w5687 = w5684 & w5685;
assign v2723 = ~(w5686 | w5687);
assign w5688 = v2723;
assign w5689 = w5564 & ~w5688;
assign w5690 = ~w5564 & w5688;
assign v2724 = ~(w5689 | w5690);
assign w5691 = v2724;
assign v2725 = ~(w5683 | w5691);
assign w5692 = v2725;
assign w5693 = w5683 & w5691;
assign v2726 = ~(w5692 | w5693);
assign w5694 = v2726;
assign w5695 = pi00 & pi53;
assign w5696 = pi05 & pi48;
assign w5697 = pi16 & pi37;
assign v2727 = ~(w5696 | w5697);
assign w5698 = v2727;
assign w5699 = w5696 & w5697;
assign v2728 = ~(w5698 | w5699);
assign w5700 = v2728;
assign w5701 = w5695 & ~w5700;
assign w5702 = ~w5695 & w5700;
assign v2729 = ~(w5701 | w5702);
assign w5703 = v2729;
assign w5704 = w5694 & ~w5703;
assign w5705 = ~w5694 & w5703;
assign v2730 = ~(w5704 | w5705);
assign w5706 = v2730;
assign v2731 = ~(w5674 | w5706);
assign w5707 = v2731;
assign w5708 = w5674 & w5706;
assign v2732 = ~(w5707 | w5708);
assign w5709 = v2732;
assign v2733 = ~(w5521 | w5523);
assign w5710 = v2733;
assign v2734 = ~(w5457 | w5460);
assign w5711 = v2734;
assign w5712 = pi13 & pi40;
assign w5713 = pi10 & pi43;
assign v2735 = ~(w5542 | w5713);
assign w5714 = v2735;
assign w5715 = w5542 & w5713;
assign v2736 = ~(w5714 | w5715);
assign w5716 = v2736;
assign w5717 = w5712 & ~w5716;
assign w5718 = ~w5712 & w5716;
assign v2737 = ~(w5717 | w5718);
assign w5719 = v2737;
assign w5720 = pi22 & pi31;
assign w5721 = pi24 & pi29;
assign w5722 = pi23 & pi30;
assign v2738 = ~(w5721 | w5722);
assign w5723 = v2738;
assign w5724 = w5721 & w5722;
assign v2739 = ~(w5723 | w5724);
assign w5725 = v2739;
assign w5726 = w5720 & ~w5725;
assign w5727 = ~w5720 & w5725;
assign v2740 = ~(w5726 | w5727);
assign w5728 = v2740;
assign v2741 = ~(w5719 | w5728);
assign w5729 = v2741;
assign w5730 = w5719 & w5728;
assign v2742 = ~(w5729 | w5730);
assign w5731 = v2742;
assign w5732 = pi11 & pi42;
assign w5733 = pi26 & pi27;
assign w5734 = pi25 & pi28;
assign v2743 = ~(w5733 | w5734);
assign w5735 = v2743;
assign w5736 = w5733 & w5734;
assign v2744 = ~(w5735 | w5736);
assign w5737 = v2744;
assign w5738 = w5732 & ~w5737;
assign w5739 = ~w5732 & w5737;
assign v2745 = ~(w5738 | w5739);
assign w5740 = v2745;
assign w5741 = w5731 & ~w5740;
assign w5742 = ~w5731 & w5740;
assign v2746 = ~(w5741 | w5742);
assign w5743 = v2746;
assign w5744 = ~w5711 & w5743;
assign w5745 = w5711 & ~w5743;
assign v2747 = ~(w5744 | w5745);
assign w5746 = v2747;
assign w5747 = ~w5710 & w5746;
assign w5748 = w5710 & ~w5746;
assign v2748 = ~(w5747 | w5748);
assign w5749 = v2748;
assign w5750 = w5709 & w5749;
assign v2749 = ~(w5709 | w5749);
assign w5751 = v2749;
assign v2750 = ~(w5750 | w5751);
assign w5752 = v2750;
assign w5753 = ~w5638 & w5752;
assign w5754 = w5638 & ~w5752;
assign v2751 = ~(w5753 | w5754);
assign w5755 = v2751;
assign w5756 = ~w5637 & w5755;
assign w5757 = w5637 & ~w5755;
assign v2752 = ~(w5756 | w5757);
assign w5758 = v2752;
assign v2753 = ~(w5476 | w5479);
assign w5759 = v2753;
assign v2754 = ~(w5478 | w5759);
assign w5760 = v2754;
assign w5761 = w5423 & ~w5425;
assign v2755 = ~(w5427 | w5761);
assign w5762 = v2755;
assign w5763 = w5760 & ~w5762;
assign w5764 = ~w5760 & w5762;
assign v2756 = ~(w5763 | w5764);
assign w5765 = v2756;
assign v2757 = ~(w5582 | w5586);
assign w5766 = v2757;
assign v2758 = ~(w5585 | w5766);
assign w5767 = v2758;
assign v2759 = ~(w5765 | w5767);
assign w5768 = v2759;
assign w5769 = w5765 & w5767;
assign v2760 = ~(w5768 | w5769);
assign w5770 = v2760;
assign w5771 = (~w5591 & ~w5593) | (~w5591 & w16892) | (~w5593 & w16892);
assign w5772 = (~w5473 & ~w5475) | (~w5473 & w16893) | (~w5475 & w16893);
assign v2761 = ~(w5771 | w5772);
assign w5773 = v2761;
assign w5774 = w5771 & w5772;
assign v2762 = ~(w5773 | w5774);
assign w5775 = v2762;
assign w5776 = w5770 & w5775;
assign v2763 = ~(w5770 | w5775);
assign w5777 = v2763;
assign v2764 = ~(w5776 | w5777);
assign w5778 = v2764;
assign v2765 = ~(w5573 | w5577);
assign w5779 = v2765;
assign v2766 = ~(w5576 | w5779);
assign w5780 = v2766;
assign v2767 = ~(w5548 | w5552);
assign w5781 = v2767;
assign v2768 = ~(w5551 | w5781);
assign w5782 = v2768;
assign w5783 = w5780 & w5782;
assign v2769 = ~(w5780 | w5782);
assign w5784 = v2769;
assign v2770 = ~(w5783 | w5784);
assign w5785 = v2770;
assign w5786 = w5560 & ~w5563;
assign v2771 = ~(w5565 | w5786);
assign w5787 = v2771;
assign w5788 = ~w5785 & w5787;
assign w5789 = w5785 & ~w5787;
assign v2772 = ~(w5788 | w5789);
assign w5790 = v2772;
assign v2773 = ~(w5557 | w5570);
assign w5791 = v2773;
assign w5792 = pi52 & w1542;
assign w5793 = pi01 & pi52;
assign v2774 = ~(pi27 | w5793);
assign w5794 = v2774;
assign v2775 = ~(w5792 | w5794);
assign w5795 = v2775;
assign w5796 = w5538 & ~w5541;
assign v2776 = ~(w5543 | w5796);
assign w5797 = v2776;
assign w5798 = w5795 & ~w5797;
assign w5799 = ~w5795 & w5797;
assign v2777 = ~(w5798 | w5799);
assign w5800 = v2777;
assign v2778 = ~(w5594 | w5598);
assign w5801 = v2778;
assign v2779 = ~(w5597 | w5801);
assign w5802 = v2779;
assign w5803 = w5800 & w5802;
assign v2780 = ~(w5800 | w5802);
assign w5804 = v2780;
assign v2781 = ~(w5803 | w5804);
assign w5805 = v2781;
assign w5806 = ~w5791 & w5805;
assign w5807 = w5791 & ~w5805;
assign v2782 = ~(w5806 | w5807);
assign w5808 = v2782;
assign v2783 = ~(w5790 | w5808);
assign w5809 = v2783;
assign w5810 = w5790 & w5808;
assign v2784 = ~(w5809 | w5810);
assign w5811 = v2784;
assign v2785 = ~(w5778 | w5811);
assign w5812 = v2785;
assign w5813 = w5778 & w5811;
assign v2786 = ~(w5812 | w5813);
assign w5814 = v2786;
assign w5815 = (~w5440 & ~w5441) | (~w5440 & w17113) | (~w5441 & w17113);
assign w5816 = ~w5814 & w5815;
assign w5817 = w5814 & ~w5815;
assign v2787 = ~(w5816 | w5817);
assign w5818 = v2787;
assign v2788 = ~(w5606 | w5609);
assign w5819 = v2788;
assign w5820 = (~w5511 & ~w5513) | (~w5511 & w17114) | (~w5513 & w17114);
assign w5821 = (~w5499 & ~w5501) | (~w5499 & w16742) | (~w5501 & w16742);
assign w5822 = (~w5449 & ~w5451) | (~w5449 & w16894) | (~w5451 & w16894);
assign v2789 = ~(w5821 | w5822);
assign w5823 = v2789;
assign w5824 = w5821 & w5822;
assign v2790 = ~(w5823 | w5824);
assign w5825 = v2790;
assign w5826 = w5820 & ~w5825;
assign w5827 = ~w5820 & w5825;
assign v2791 = ~(w5826 | w5827);
assign w5828 = v2791;
assign v2792 = ~(w5488 | w5492);
assign w5829 = v2792;
assign w5830 = ~w5828 & w5829;
assign w5831 = w5828 & ~w5829;
assign v2793 = ~(w5830 | w5831);
assign w5832 = v2793;
assign w5833 = ~w5819 & w5832;
assign w5834 = w5819 & ~w5832;
assign v2794 = ~(w5833 | w5834);
assign w5835 = v2794;
assign v2795 = ~(w5612 | w5616);
assign w5836 = v2795;
assign w5837 = ~w5835 & w5836;
assign w5838 = w5835 & ~w5836;
assign v2796 = ~(w5837 | w5838);
assign w5839 = v2796;
assign w5840 = w5818 & w5839;
assign v2797 = ~(w5818 | w5839);
assign w5841 = v2797;
assign v2798 = ~(w5840 | w5841);
assign w5842 = v2798;
assign w5843 = w5758 & w5842;
assign v2799 = ~(w5758 | w5842);
assign w5844 = v2799;
assign v2800 = ~(w5843 | w5844);
assign w5845 = v2800;
assign w5846 = ~w5636 & w5845;
assign w5847 = w5636 & ~w5845;
assign v2801 = ~(w5846 | w5847);
assign w5848 = v2801;
assign w5849 = w5635 & w5848;
assign v2802 = ~(w5635 | w5848);
assign w5850 = v2802;
assign v2803 = ~(w5849 | w5850);
assign w5851 = v2803;
assign v2804 = ~(w5756 | w5843);
assign w5852 = v2804;
assign v2805 = ~(w5750 | w5753);
assign w5853 = v2805;
assign w5854 = (~w5798 & ~w5800) | (~w5798 & w17115) | (~w5800 & w17115);
assign w5855 = (~w5783 & ~w5785) | (~w5783 & w16743) | (~w5785 & w16743);
assign w5856 = (~w5763 & ~w5765) | (~w5763 & w16744) | (~w5765 & w16744);
assign v2806 = ~(w5855 | w5856);
assign w5857 = v2806;
assign w5858 = w5855 & w5856;
assign v2807 = ~(w5857 | w5858);
assign w5859 = v2807;
assign w5860 = w5854 & ~w5859;
assign w5861 = ~w5854 & w5859;
assign v2808 = ~(w5860 | w5861);
assign w5862 = v2808;
assign w5863 = (~w5672 & ~w5674) | (~w5672 & w17116) | (~w5674 & w17116);
assign w5864 = ~w5862 & w5863;
assign w5865 = w5862 & ~w5863;
assign v2809 = ~(w5864 | w5865);
assign w5866 = v2809;
assign v2810 = ~(w5695 | w5699);
assign w5867 = v2810;
assign v2811 = ~(w5698 | w5867);
assign w5868 = v2811;
assign v2812 = ~(w5675 | w5679);
assign w5869 = v2812;
assign v2813 = ~(w5678 | w5869);
assign w5870 = v2813;
assign w5871 = w5868 & w5870;
assign v2814 = ~(w5868 | w5870);
assign w5872 = v2814;
assign v2815 = ~(w5871 | w5872);
assign w5873 = v2815;
assign v2816 = ~(w5732 | w5736);
assign w5874 = v2816;
assign v2817 = ~(w5735 | w5874);
assign w5875 = v2817;
assign v2818 = ~(w5873 | w5875);
assign w5876 = v2818;
assign w5877 = w5873 & w5875;
assign v2819 = ~(w5876 | w5877);
assign w5878 = v2819;
assign v2820 = ~(w5648 | w5652);
assign w5879 = v2820;
assign v2821 = ~(w5651 | w5879);
assign w5880 = v2821;
assign v2822 = ~(w5660 | w5664);
assign w5881 = v2822;
assign v2823 = ~(w5663 | w5881);
assign w5882 = v2823;
assign w5883 = w5880 & w5882;
assign v2824 = ~(w5880 | w5882);
assign w5884 = v2824;
assign v2825 = ~(w5883 | w5884);
assign w5885 = v2825;
assign v2826 = ~(w5720 | w5724);
assign w5886 = v2826;
assign v2827 = ~(w5723 | w5886);
assign w5887 = v2827;
assign v2828 = ~(w5885 | w5887);
assign w5888 = v2828;
assign w5889 = w5885 & w5887;
assign v2829 = ~(w5888 | w5889);
assign w5890 = v2829;
assign v2830 = ~(w5692 | w5704);
assign w5891 = v2830;
assign w5892 = ~w5890 & w5891;
assign w5893 = w5890 & ~w5891;
assign v2831 = ~(w5892 | w5893);
assign w5894 = v2831;
assign w5895 = w5878 & w5894;
assign v2832 = ~(w5878 | w5894);
assign w5896 = v2832;
assign v2833 = ~(w5895 | w5896);
assign w5897 = v2833;
assign w5898 = w5866 & w5897;
assign v2834 = ~(w5866 | w5897);
assign w5899 = v2834;
assign v2835 = ~(w5898 | w5899);
assign w5900 = v2835;
assign w5901 = ~w5853 & w5900;
assign w5902 = w5853 & ~w5900;
assign v2836 = ~(w5901 | w5902);
assign w5903 = v2836;
assign w5904 = (~w5823 & ~w5825) | (~w5823 & w16895) | (~w5825 & w16895);
assign w5905 = pi13 & pi41;
assign w5906 = pi12 & pi42;
assign w5907 = pi11 & pi43;
assign v2837 = ~(w5906 | w5907);
assign w5908 = v2837;
assign w5909 = pi12 & pi43;
assign w5910 = w5732 & w5909;
assign v2838 = ~(w5908 | w5910);
assign w5911 = v2838;
assign w5912 = w5905 & ~w5911;
assign w5913 = ~w5905 & w5911;
assign v2839 = ~(w5912 | w5913);
assign w5914 = v2839;
assign w5915 = pi20 & pi34;
assign w5916 = pi18 & pi36;
assign w5917 = pi05 & pi49;
assign v2840 = ~(w5916 | w5917);
assign w5918 = v2840;
assign w5919 = w5916 & w5917;
assign v2841 = ~(w5918 | w5919);
assign w5920 = v2841;
assign w5921 = w5915 & ~w5920;
assign w5922 = ~w5915 & w5920;
assign v2842 = ~(w5921 | w5922);
assign w5923 = v2842;
assign v2843 = ~(w5914 | w5923);
assign w5924 = v2843;
assign w5925 = w5914 & w5923;
assign v2844 = ~(w5924 | w5925);
assign w5926 = v2844;
assign w5927 = pi17 & pi37;
assign w5928 = pi06 & pi48;
assign w5929 = pi16 & pi38;
assign v2845 = ~(w5928 | w5929);
assign w5930 = v2845;
assign w5931 = w5928 & w5929;
assign v2846 = ~(w5930 | w5931);
assign w5932 = v2846;
assign w5933 = w5927 & ~w5932;
assign w5934 = ~w5927 & w5932;
assign v2847 = ~(w5933 | w5934);
assign w5935 = v2847;
assign w5936 = w5926 & ~w5935;
assign w5937 = ~w5926 & w5935;
assign v2848 = ~(w5936 | w5937);
assign w5938 = v2848;
assign w5939 = ~w5904 & w5938;
assign w5940 = w5904 & ~w5938;
assign v2849 = ~(w5939 | w5940);
assign w5941 = v2849;
assign w5942 = pi02 & pi52;
assign w5943 = pi04 & pi50;
assign v2850 = ~(w5642 | w5943);
assign w5944 = v2850;
assign w5945 = pi04 & pi51;
assign w5946 = w5426 & w5945;
assign v2851 = ~(w5944 | w5946);
assign w5947 = v2851;
assign w5948 = w5942 & ~w5947;
assign w5949 = ~w5942 & w5947;
assign v2852 = ~(w5948 | w5949);
assign w5950 = v2852;
assign w5951 = pi07 & pi47;
assign w5952 = pi15 & pi39;
assign w5953 = pi08 & pi46;
assign v2853 = ~(w5952 | w5953);
assign w5954 = v2853;
assign w5955 = w5952 & w5953;
assign v2854 = ~(w5954 | w5955);
assign w5956 = v2854;
assign w5957 = w5951 & ~w5956;
assign w5958 = ~w5951 & w5956;
assign v2855 = ~(w5957 | w5958);
assign w5959 = v2855;
assign v2856 = ~(w5950 | w5959);
assign w5960 = v2856;
assign w5961 = w5950 & w5959;
assign v2857 = ~(w5960 | w5961);
assign w5962 = v2857;
assign w5963 = pi09 & pi45;
assign w5964 = pi14 & pi40;
assign w5965 = pi10 & pi44;
assign v2858 = ~(w5964 | w5965);
assign w5966 = v2858;
assign w5967 = w5964 & w5965;
assign v2859 = ~(w5966 | w5967);
assign w5968 = v2859;
assign w5969 = w5963 & ~w5968;
assign w5970 = ~w5963 & w5968;
assign v2860 = ~(w5969 | w5970);
assign w5971 = v2860;
assign w5972 = w5962 & ~w5971;
assign w5973 = ~w5962 & w5971;
assign v2861 = ~(w5972 | w5973);
assign w5974 = v2861;
assign v2862 = ~(w5941 | w5974);
assign w5975 = v2862;
assign w5976 = w5941 & w5974;
assign v2863 = ~(w5975 | w5976);
assign w5977 = v2863;
assign v2864 = ~(w5744 | w5747);
assign w5978 = v2864;
assign v2865 = ~(w5564 | w5687);
assign w5979 = v2865;
assign v2866 = ~(w5686 | w5979);
assign w5980 = v2866;
assign w5981 = w5447 & ~w5641;
assign v2867 = ~(w5643 | w5981);
assign w5982 = v2867;
assign w5983 = w5980 & ~w5982;
assign w5984 = ~w5980 & w5982;
assign v2868 = ~(w5983 | w5984);
assign w5985 = v2868;
assign v2869 = ~(w5712 | w5715);
assign w5986 = v2869;
assign v2870 = ~(w5714 | w5986);
assign w5987 = v2870;
assign v2871 = ~(w5985 | w5987);
assign w5988 = v2871;
assign w5989 = w5985 & w5987;
assign v2872 = ~(w5988 | w5989);
assign w5990 = v2872;
assign w5991 = (~w5729 & ~w5731) | (~w5729 & w16896) | (~w5731 & w16896);
assign w5992 = (~w5657 & ~w5659) | (~w5657 & w16897) | (~w5659 & w16897);
assign v2873 = ~(w5991 | w5992);
assign w5993 = v2873;
assign w5994 = w5991 & w5992;
assign v2874 = ~(w5993 | w5994);
assign w5995 = v2874;
assign w5996 = w5990 & w5995;
assign v2875 = ~(w5990 | w5995);
assign w5997 = v2875;
assign v2876 = ~(w5996 | w5997);
assign w5998 = v2876;
assign w5999 = ~w5978 & w5998;
assign w6000 = w5978 & ~w5998;
assign v2877 = ~(w5999 | w6000);
assign w6001 = v2877;
assign v2878 = ~(w5977 | w6001);
assign w6002 = v2878;
assign w6003 = w5977 & w6001;
assign v2879 = ~(w6002 | w6003);
assign w6004 = v2879;
assign v2880 = ~(w5903 | w6004);
assign w6005 = v2880;
assign w6006 = w5903 & w6004;
assign v2881 = ~(w6005 | w6006);
assign w6007 = v2881;
assign v2882 = ~(w5806 | w5810);
assign w6008 = v2882;
assign w6009 = (~w5773 & ~w5775) | (~w5773 & w17117) | (~w5775 & w17117);
assign w6010 = pi00 & pi54;
assign w6011 = w5792 & w6010;
assign v2883 = ~(w5792 | w6010);
assign w6012 = v2883;
assign v2884 = ~(w6011 | w6012);
assign w6013 = v2884;
assign w6014 = pi26 & pi28;
assign w6015 = pi01 & pi53;
assign v2885 = ~(w6014 | w6015);
assign w6016 = v2885;
assign w6017 = w6014 & w6015;
assign v2886 = ~(w6016 | w6017);
assign w6018 = v2886;
assign w6019 = w6013 & w6018;
assign v2887 = ~(w6013 | w6018);
assign w6020 = v2887;
assign v2888 = ~(w6019 | w6020);
assign w6021 = v2888;
assign w6022 = pi19 & pi35;
assign w6023 = pi21 & pi33;
assign w6024 = pi22 & pi32;
assign v2889 = ~(w6023 | w6024);
assign w6025 = v2889;
assign w6026 = w6023 & w6024;
assign v2890 = ~(w6025 | w6026);
assign w6027 = v2890;
assign w6028 = w6022 & ~w6027;
assign w6029 = ~w6022 & w6027;
assign v2891 = ~(w6028 | w6029);
assign w6030 = v2891;
assign w6031 = pi23 & pi31;
assign w6032 = pi24 & pi30;
assign w6033 = pi25 & pi29;
assign v2892 = ~(w6032 | w6033);
assign w6034 = v2892;
assign w6035 = w6032 & w6033;
assign v2893 = ~(w6034 | w6035);
assign w6036 = v2893;
assign w6037 = w6031 & ~w6036;
assign w6038 = ~w6031 & w6036;
assign v2894 = ~(w6037 | w6038);
assign w6039 = v2894;
assign v2895 = ~(w6030 | w6039);
assign w6040 = v2895;
assign w6041 = w6030 & w6039;
assign v2896 = ~(w6040 | w6041);
assign w6042 = v2896;
assign w6043 = w6021 & w6042;
assign v2897 = ~(w6021 | w6042);
assign w6044 = v2897;
assign v2898 = ~(w6043 | w6044);
assign w6045 = v2898;
assign w6046 = ~w6009 & w6045;
assign w6047 = w6009 & ~w6045;
assign v2899 = ~(w6046 | w6047);
assign w6048 = v2899;
assign w6049 = ~w6008 & w6048;
assign w6050 = w6008 & ~w6048;
assign v2900 = ~(w6049 | w6050);
assign w6051 = v2900;
assign v2901 = ~(w5813 | w5817);
assign w6052 = v2901;
assign v2902 = ~(w5831 | w5833);
assign w6053 = v2902;
assign v2903 = ~(w6052 | w6053);
assign w6054 = v2903;
assign w6055 = w6052 & w6053;
assign v2904 = ~(w6054 | w6055);
assign w6056 = v2904;
assign v2905 = ~(w6051 | w6056);
assign w6057 = v2905;
assign w6058 = w6051 & w6056;
assign v2906 = ~(w6057 | w6058);
assign w6059 = v2906;
assign v2907 = ~(w5838 | w5840);
assign w6060 = v2907;
assign w6061 = w6059 & ~w6060;
assign w6062 = ~w6059 & w6060;
assign v2908 = ~(w6061 | w6062);
assign w6063 = v2908;
assign w6064 = w6007 & w6063;
assign v2909 = ~(w6007 | w6063);
assign w6065 = v2909;
assign v2910 = ~(w6064 | w6065);
assign w6066 = v2910;
assign w6067 = ~w5852 & w6066;
assign w6068 = w5852 & ~w6066;
assign v2911 = ~(w6067 | w6068);
assign w6069 = v2911;
assign v2912 = ~(w5625 | w5846);
assign w6070 = v2912;
assign w6071 = (w5207 & w16534) | (w5207 & w16535) | (w16534 & w16535);
assign w6072 = w6069 & w6071;
assign v2913 = ~(w6069 | w6071);
assign w6073 = v2913;
assign v2914 = ~(w6072 | w6073);
assign w6074 = v2914;
assign v2915 = ~(w6061 | w6064);
assign w6075 = v2915;
assign v2916 = ~(w6054 | w6058);
assign w6076 = v2916;
assign w6077 = (~w6011 & ~w6013) | (~w6011 & w16745) | (~w6013 & w16745);
assign v2917 = ~(w5951 | w5955);
assign w6078 = v2917;
assign v2918 = ~(w5954 | w6078);
assign w6079 = v2918;
assign w6080 = ~w6077 & w6079;
assign w6081 = w6077 & ~w6079;
assign v2919 = ~(w6080 | w6081);
assign w6082 = v2919;
assign w6083 = pi05 & pi50;
assign w6084 = pi18 & pi37;
assign w6085 = pi19 & pi36;
assign v2920 = ~(w6084 | w6085);
assign w6086 = v2920;
assign w6087 = w6084 & w6085;
assign v2921 = ~(w6086 | w6087);
assign w6088 = v2921;
assign w6089 = w6083 & ~w6088;
assign w6090 = ~w6083 & w6088;
assign v2922 = ~(w6089 | w6090);
assign w6091 = v2922;
assign w6092 = ~w6082 & w6091;
assign w6093 = w6082 & ~w6091;
assign v2923 = ~(w6092 | w6093);
assign w6094 = v2923;
assign v2924 = ~(w5963 | w5967);
assign w6095 = v2924;
assign v2925 = ~(w5966 | w6095);
assign w6096 = v2925;
assign w6097 = w5942 & ~w5944;
assign v2926 = ~(w5946 | w6097);
assign w6098 = v2926;
assign w6099 = w6096 & ~w6098;
assign w6100 = ~w6096 & w6098;
assign v2927 = ~(w6099 | w6100);
assign w6101 = v2927;
assign v2928 = ~(w5915 | w5919);
assign w6102 = v2928;
assign v2929 = ~(w5918 | w6102);
assign w6103 = v2929;
assign v2930 = ~(w6101 | w6103);
assign w6104 = v2930;
assign w6105 = w6101 & w6103;
assign v2931 = ~(w6104 | w6105);
assign w6106 = v2931;
assign v2932 = ~(w6040 | w6043);
assign w6107 = v2932;
assign w6108 = ~w6106 & w6107;
assign w6109 = w6106 & ~w6107;
assign v2933 = ~(w6108 | w6109);
assign w6110 = v2933;
assign w6111 = w6094 & w6110;
assign v2934 = ~(w6094 | w6110);
assign w6112 = v2934;
assign v2935 = ~(w6111 | w6112);
assign w6113 = v2935;
assign w6114 = pi54 & w1678;
assign w6115 = pi01 & pi54;
assign v2936 = ~(pi28 | w6115);
assign w6116 = v2936;
assign v2937 = ~(w6114 | w6116);
assign w6117 = v2937;
assign v2938 = ~(w6017 | w6117);
assign w6118 = v2938;
assign w6119 = ~pi54 & w6017;
assign v2939 = ~(w6118 | w6119);
assign w6120 = v2939;
assign w6121 = w5905 & ~w5908;
assign v2940 = ~(w5910 | w6121);
assign w6122 = v2940;
assign w6123 = w6120 & ~w6122;
assign w6124 = ~w6120 & w6122;
assign v2941 = ~(w6123 | w6124);
assign w6125 = v2941;
assign w6126 = (~w5871 & ~w5873) | (~w5871 & w16746) | (~w5873 & w16746);
assign w6127 = (~w5983 & ~w5985) | (~w5983 & w16747) | (~w5985 & w16747);
assign v2942 = ~(w6126 | w6127);
assign w6128 = v2942;
assign w6129 = w6126 & w6127;
assign v2943 = ~(w6128 | w6129);
assign w6130 = v2943;
assign v2944 = ~(w6125 | w6130);
assign w6131 = v2944;
assign w6132 = w6125 & w6130;
assign v2945 = ~(w6131 | w6132);
assign w6133 = v2945;
assign w6134 = (~w5939 & ~w5941) | (~w5939 & w17118) | (~w5941 & w17118);
assign w6135 = w6133 & ~w6134;
assign w6136 = ~w6133 & w6134;
assign v2946 = ~(w6135 | w6136);
assign w6137 = v2946;
assign w6138 = w6113 & w6137;
assign v2947 = ~(w6113 | w6137);
assign w6139 = v2947;
assign v2948 = ~(w6138 | w6139);
assign w6140 = v2948;
assign w6141 = ~w6076 & w6140;
assign w6142 = w6076 & ~w6140;
assign v2949 = ~(w6141 | w6142);
assign w6143 = v2949;
assign v2950 = ~(w6046 | w6049);
assign w6144 = v2950;
assign v2951 = ~(w6022 | w6026);
assign w6145 = v2951;
assign v2952 = ~(w6025 | w6145);
assign w6146 = v2952;
assign v2953 = ~(w6031 | w6035);
assign w6147 = v2953;
assign v2954 = ~(w6034 | w6147);
assign w6148 = v2954;
assign w6149 = w6146 & w6148;
assign v2955 = ~(w6146 | w6148);
assign w6150 = v2955;
assign v2956 = ~(w6149 | w6150);
assign w6151 = v2956;
assign v2957 = ~(w5927 | w5931);
assign w6152 = v2957;
assign v2958 = ~(w5930 | w6152);
assign w6153 = v2958;
assign v2959 = ~(w6151 | w6153);
assign w6154 = v2959;
assign w6155 = w6151 & w6153;
assign v2960 = ~(w6154 | w6155);
assign w6156 = v2960;
assign w6157 = (~w5924 & ~w5926) | (~w5924 & w17119) | (~w5926 & w17119);
assign w6158 = (~w5960 & ~w5962) | (~w5960 & w17120) | (~w5962 & w17120);
assign v2961 = ~(w6157 | w6158);
assign w6159 = v2961;
assign w6160 = w6157 & w6158;
assign v2962 = ~(w6159 | w6160);
assign w6161 = v2962;
assign w6162 = w6156 & w6161;
assign v2963 = ~(w6156 | w6161);
assign w6163 = v2963;
assign v2964 = ~(w6162 | w6163);
assign w6164 = v2964;
assign w6165 = ~w6144 & w6164;
assign w6166 = w6144 & ~w6164;
assign v2965 = ~(w6165 | w6166);
assign w6167 = v2965;
assign w6168 = (~w5857 & ~w5859) | (~w5857 & w16898) | (~w5859 & w16898);
assign w6169 = pi10 & pi45;
assign w6170 = pi13 & pi42;
assign w6171 = pi11 & pi44;
assign v2966 = ~(w6170 | w6171);
assign w6172 = v2966;
assign w6173 = pi13 & pi44;
assign w6174 = w5732 & w6173;
assign v2967 = ~(w6172 | w6174);
assign w6175 = v2967;
assign w6176 = w6169 & ~w6175;
assign w6177 = ~w6169 & w6175;
assign v2968 = ~(w6176 | w6177);
assign w6178 = v2968;
assign w6179 = pi27 & pi28;
assign w6180 = pi26 & pi29;
assign v2969 = ~(w6179 | w6180);
assign w6181 = v2969;
assign w6182 = w6179 & w6180;
assign v2970 = ~(w6181 | w6182);
assign w6183 = v2970;
assign w6184 = w5909 & ~w6183;
assign w6185 = ~w5909 & w6183;
assign v2971 = ~(w6184 | w6185);
assign w6186 = v2971;
assign v2972 = ~(w6178 | w6186);
assign w6187 = v2972;
assign w6188 = w6178 & w6186;
assign v2973 = ~(w6187 | w6188);
assign w6189 = v2973;
assign w6190 = pi16 & pi39;
assign w6191 = pi08 & pi47;
assign w6192 = pi07 & pi48;
assign v2974 = ~(w6191 | w6192);
assign w6193 = v2974;
assign w6194 = pi08 & pi48;
assign w6195 = w5951 & w6194;
assign v2975 = ~(w6193 | w6195);
assign w6196 = v2975;
assign w6197 = w6190 & ~w6196;
assign w6198 = ~w6190 & w6196;
assign v2976 = ~(w6197 | w6198);
assign w6199 = v2976;
assign w6200 = w6189 & ~w6199;
assign w6201 = ~w6189 & w6199;
assign v2977 = ~(w6200 | w6201);
assign w6202 = v2977;
assign w6203 = ~w6168 & w6202;
assign w6204 = w6168 & ~w6202;
assign v2978 = ~(w6203 | w6204);
assign w6205 = v2978;
assign w6206 = pi00 & pi55;
assign w6207 = pi02 & pi53;
assign v2979 = ~(w5945 | w6207);
assign w6208 = v2979;
assign w6209 = w5945 & w6207;
assign v2980 = ~(w6208 | w6209);
assign w6210 = v2980;
assign w6211 = w6206 & ~w6210;
assign w6212 = ~w6206 & w6210;
assign v2981 = ~(w6211 | w6212);
assign w6213 = v2981;
assign w6214 = pi20 & pi35;
assign w6215 = pi22 & pi33;
assign w6216 = pi21 & pi34;
assign v2982 = ~(w6215 | w6216);
assign w6217 = v2982;
assign w6218 = w6215 & w6216;
assign v2983 = ~(w6217 | w6218);
assign w6219 = v2983;
assign w6220 = w6214 & ~w6219;
assign w6221 = ~w6214 & w6219;
assign v2984 = ~(w6220 | w6221);
assign w6222 = v2984;
assign v2985 = ~(w6213 | w6222);
assign w6223 = v2985;
assign w6224 = w6213 & w6222;
assign v2986 = ~(w6223 | w6224);
assign w6225 = v2986;
assign w6226 = pi23 & pi32;
assign w6227 = pi25 & pi30;
assign w6228 = pi24 & pi31;
assign v2987 = ~(w6227 | w6228);
assign w6229 = v2987;
assign w6230 = w6227 & w6228;
assign v2988 = ~(w6229 | w6230);
assign w6231 = v2988;
assign w6232 = w6226 & ~w6231;
assign w6233 = ~w6226 & w6231;
assign v2989 = ~(w6232 | w6233);
assign w6234 = v2989;
assign w6235 = w6225 & ~w6234;
assign w6236 = ~w6225 & w6234;
assign v2990 = ~(w6235 | w6236);
assign w6237 = v2990;
assign w6238 = w6205 & w6237;
assign v2991 = ~(w6205 | w6237);
assign w6239 = v2991;
assign v2992 = ~(w6238 | w6239);
assign w6240 = v2992;
assign w6241 = w6167 & w6240;
assign v2993 = ~(w6167 | w6240);
assign w6242 = v2993;
assign v2994 = ~(w6241 | w6242);
assign w6243 = v2994;
assign v2995 = ~(w6143 | w6243);
assign w6244 = v2995;
assign w6245 = w6143 & w6243;
assign v2996 = ~(w6244 | w6245);
assign w6246 = v2996;
assign v2997 = ~(w5901 | w6006);
assign w6247 = v2997;
assign v2998 = ~(w5999 | w6003);
assign w6248 = v2998;
assign v2999 = ~(w5865 | w5898);
assign w6249 = v2999;
assign v3000 = ~(w5893 | w5895);
assign w6250 = v3000;
assign w6251 = (~w5883 & ~w5885) | (~w5883 & w16748) | (~w5885 & w16748);
assign w6252 = pi15 & pi40;
assign w6253 = pi14 & pi41;
assign w6254 = pi09 & pi46;
assign v3001 = ~(w6253 | w6254);
assign w6255 = v3001;
assign w6256 = w6253 & w6254;
assign v3002 = ~(w6255 | w6256);
assign w6257 = v3002;
assign w6258 = w6252 & ~w6257;
assign w6259 = ~w6252 & w6257;
assign v3003 = ~(w6258 | w6259);
assign w6260 = v3003;
assign w6261 = pi03 & pi52;
assign w6262 = pi06 & pi49;
assign w6263 = pi17 & pi38;
assign v3004 = ~(w6262 | w6263);
assign w6264 = v3004;
assign w6265 = w6262 & w6263;
assign v3005 = ~(w6264 | w6265);
assign w6266 = v3005;
assign w6267 = w6261 & ~w6266;
assign w6268 = ~w6261 & w6266;
assign v3006 = ~(w6267 | w6268);
assign w6269 = v3006;
assign v3007 = ~(w6260 | w6269);
assign w6270 = v3007;
assign w6271 = w6260 & w6269;
assign v3008 = ~(w6270 | w6271);
assign w6272 = v3008;
assign w6273 = w6251 & ~w6272;
assign w6274 = ~w6251 & w6272;
assign v3009 = ~(w6273 | w6274);
assign w6275 = v3009;
assign w6276 = (~w5993 & ~w5995) | (~w5993 & w17121) | (~w5995 & w17121);
assign w6277 = ~w6275 & w6276;
assign w6278 = w6275 & ~w6276;
assign v3010 = ~(w6277 | w6278);
assign w6279 = v3010;
assign w6280 = ~w6250 & w6279;
assign w6281 = w6250 & ~w6279;
assign v3011 = ~(w6280 | w6281);
assign w6282 = v3011;
assign w6283 = ~w6249 & w6282;
assign w6284 = w6249 & ~w6282;
assign v3012 = ~(w6283 | w6284);
assign w6285 = v3012;
assign w6286 = ~w6248 & w6285;
assign w6287 = w6248 & ~w6285;
assign v3013 = ~(w6286 | w6287);
assign w6288 = v3013;
assign w6289 = ~w6247 & w6288;
assign w6290 = w6247 & ~w6288;
assign v3014 = ~(w6289 | w6290);
assign w6291 = v3014;
assign w6292 = w6246 & w6291;
assign v3015 = ~(w6246 | w6291);
assign w6293 = v3015;
assign v3016 = ~(w6292 | w6293);
assign w6294 = v3016;
assign w6295 = ~w6075 & w6294;
assign w6296 = w6075 & ~w6294;
assign v3017 = ~(w6295 | w6296);
assign w6297 = v3017;
assign w6298 = (~w5207 & w16536) | (~w5207 & w16537) | (w16536 & w16537);
assign v3018 = ~(w6068 | w6298);
assign w6299 = v3018;
assign w6300 = w6297 & w6299;
assign v3019 = ~(w6297 | w6299);
assign w6301 = v3019;
assign v3020 = ~(w6300 | w6301);
assign w6302 = v3020;
assign v3021 = ~(w6289 | w6292);
assign w6303 = v3021;
assign v3022 = ~(w6278 | w6280);
assign w6304 = v3022;
assign v3023 = ~(w6214 | w6218);
assign w6305 = v3023;
assign v3024 = ~(w6217 | w6305);
assign w6306 = v3024;
assign v3025 = ~(w6226 | w6230);
assign w6307 = v3025;
assign v3026 = ~(w6229 | w6307);
assign w6308 = v3026;
assign w6309 = w6306 & w6308;
assign v3027 = ~(w6306 | w6308);
assign w6310 = v3027;
assign v3028 = ~(w6309 | w6310);
assign w6311 = v3028;
assign v3029 = ~(w6261 | w6265);
assign w6312 = v3029;
assign v3030 = ~(w6264 | w6312);
assign w6313 = v3030;
assign v3031 = ~(w6311 | w6313);
assign w6314 = v3031;
assign w6315 = w6311 & w6313;
assign v3032 = ~(w6314 | w6315);
assign w6316 = v3032;
assign w6317 = (~w6187 & ~w6189) | (~w6187 & w16899) | (~w6189 & w16899);
assign w6318 = pi27 & pi29;
assign w6319 = pi01 & pi55;
assign v3033 = ~(w6318 | w6319);
assign w6320 = v3033;
assign w6321 = w6318 & w6319;
assign v3034 = ~(w6320 | w6321);
assign w6322 = v3034;
assign v3035 = ~(w5909 | w6182);
assign w6323 = v3035;
assign v3036 = ~(w6181 | w6323);
assign w6324 = v3036;
assign w6325 = w6322 & w6324;
assign v3037 = ~(w6322 | w6324);
assign w6326 = v3037;
assign v3038 = ~(w6325 | w6326);
assign w6327 = v3038;
assign w6328 = w6169 & ~w6172;
assign v3039 = ~(w6174 | w6328);
assign w6329 = v3039;
assign w6330 = w6327 & ~w6329;
assign w6331 = ~w6327 & w6329;
assign v3040 = ~(w6330 | w6331);
assign w6332 = v3040;
assign w6333 = ~w6317 & w6332;
assign w6334 = w6317 & ~w6332;
assign v3041 = ~(w6333 | w6334);
assign w6335 = v3041;
assign w6336 = w6316 & w6335;
assign v3042 = ~(w6316 | w6335);
assign w6337 = v3042;
assign v3043 = ~(w6336 | w6337);
assign w6338 = v3043;
assign w6339 = ~w6304 & w6338;
assign w6340 = w6304 & ~w6338;
assign v3044 = ~(w6339 | w6340);
assign w6341 = v3044;
assign w6342 = w6190 & ~w6193;
assign v3045 = ~(w6195 | w6342);
assign w6343 = v3045;
assign w6344 = pi00 & pi56;
assign w6345 = pi02 & pi54;
assign v3046 = ~(w6344 | w6345);
assign w6346 = v3046;
assign w6347 = pi02 & pi56;
assign w6348 = w6010 & w6347;
assign v3047 = ~(w6346 | w6348);
assign w6349 = v3047;
assign w6350 = w6114 & ~w6349;
assign w6351 = ~w6114 & w6349;
assign v3048 = ~(w6350 | w6351);
assign w6352 = v3048;
assign v3049 = ~(w6343 | w6352);
assign w6353 = v3049;
assign w6354 = w6343 & w6352;
assign v3050 = ~(w6353 | w6354);
assign w6355 = v3050;
assign w6356 = pi03 & pi53;
assign w6357 = pi19 & pi37;
assign w6358 = pi04 & pi52;
assign v3051 = ~(w6357 | w6358);
assign w6359 = v3051;
assign w6360 = w6357 & w6358;
assign v3052 = ~(w6359 | w6360);
assign w6361 = v3052;
assign w6362 = w6356 & ~w6361;
assign w6363 = ~w6356 & w6361;
assign v3053 = ~(w6362 | w6363);
assign w6364 = v3053;
assign w6365 = ~w6355 & w6364;
assign w6366 = w6355 & ~w6364;
assign v3054 = ~(w6365 | w6366);
assign w6367 = v3054;
assign w6368 = pi11 & pi45;
assign w6369 = pi13 & pi43;
assign w6370 = pi12 & pi44;
assign v3055 = ~(w6369 | w6370);
assign w6371 = v3055;
assign w6372 = w5909 & w6173;
assign v3056 = ~(w6371 | w6372);
assign w6373 = v3056;
assign w6374 = w6368 & ~w6373;
assign w6375 = ~w6368 & w6373;
assign v3057 = ~(w6374 | w6375);
assign w6376 = v3057;
assign w6377 = pi06 & pi50;
assign w6378 = pi07 & pi49;
assign w6379 = pi17 & pi39;
assign v3058 = ~(w6378 | w6379);
assign w6380 = v3058;
assign w6381 = w6378 & w6379;
assign v3059 = ~(w6380 | w6381);
assign w6382 = v3059;
assign w6383 = w6377 & ~w6382;
assign w6384 = ~w6377 & w6382;
assign v3060 = ~(w6383 | w6384);
assign w6385 = v3060;
assign v3061 = ~(w6376 | w6385);
assign w6386 = v3061;
assign w6387 = w6376 & w6385;
assign v3062 = ~(w6386 | w6387);
assign w6388 = v3062;
assign w6389 = pi16 & pi40;
assign w6390 = pi15 & pi41;
assign v3063 = ~(w6194 | w6390);
assign w6391 = v3063;
assign w6392 = w6194 & w6390;
assign v3064 = ~(w6391 | w6392);
assign w6393 = v3064;
assign w6394 = w6389 & ~w6393;
assign w6395 = ~w6389 & w6393;
assign v3065 = ~(w6394 | w6395);
assign w6396 = v3065;
assign w6397 = w6388 & ~w6396;
assign w6398 = ~w6388 & w6396;
assign v3066 = ~(w6397 | w6398);
assign w6399 = v3066;
assign w6400 = pi20 & pi36;
assign w6401 = pi22 & pi34;
assign w6402 = pi23 & pi33;
assign v3067 = ~(w6401 | w6402);
assign w6403 = v3067;
assign w6404 = w6401 & w6402;
assign v3068 = ~(w6403 | w6404);
assign w6405 = v3068;
assign w6406 = w6400 & ~w6405;
assign w6407 = ~w6400 & w6405;
assign v3069 = ~(w6406 | w6407);
assign w6408 = v3069;
assign w6409 = pi24 & pi32;
assign w6410 = pi25 & pi31;
assign w6411 = pi26 & pi30;
assign v3070 = ~(w6410 | w6411);
assign w6412 = v3070;
assign w6413 = w6410 & w6411;
assign v3071 = ~(w6412 | w6413);
assign w6414 = v3071;
assign w6415 = w6409 & ~w6414;
assign w6416 = ~w6409 & w6414;
assign v3072 = ~(w6415 | w6416);
assign w6417 = v3072;
assign v3073 = ~(w6408 | w6417);
assign w6418 = v3073;
assign w6419 = w6408 & w6417;
assign v3074 = ~(w6418 | w6419);
assign w6420 = v3074;
assign w6421 = pi09 & pi47;
assign w6422 = pi14 & pi42;
assign w6423 = pi10 & pi46;
assign v3075 = ~(w6422 | w6423);
assign w6424 = v3075;
assign w6425 = w6422 & w6423;
assign v3076 = ~(w6424 | w6425);
assign w6426 = v3076;
assign w6427 = w6421 & ~w6426;
assign w6428 = ~w6421 & w6426;
assign v3077 = ~(w6427 | w6428);
assign w6429 = v3077;
assign w6430 = w6420 & ~w6429;
assign w6431 = ~w6420 & w6429;
assign v3078 = ~(w6430 | w6431);
assign w6432 = v3078;
assign w6433 = w6399 & w6432;
assign v3079 = ~(w6399 | w6432);
assign w6434 = v3079;
assign v3080 = ~(w6433 | w6434);
assign w6435 = v3080;
assign w6436 = w6367 & w6435;
assign v3081 = ~(w6367 | w6435);
assign w6437 = v3081;
assign v3082 = ~(w6436 | w6437);
assign w6438 = v3082;
assign v3083 = ~(w6341 | w6438);
assign w6439 = v3083;
assign w6440 = w6341 & w6438;
assign v3084 = ~(w6439 | w6440);
assign w6441 = v3084;
assign v3085 = ~(w6283 | w6286);
assign w6442 = v3085;
assign v3086 = ~(w6083 | w6087);
assign w6443 = v3086;
assign v3087 = ~(w6086 | w6443);
assign w6444 = v3087;
assign v3088 = ~(w6206 | w6209);
assign w6445 = v3088;
assign v3089 = ~(w6208 | w6445);
assign w6446 = v3089;
assign w6447 = w6444 & w6446;
assign v3090 = ~(w6444 | w6446);
assign w6448 = v3090;
assign v3091 = ~(w6447 | w6448);
assign w6449 = v3091;
assign v3092 = ~(w6252 | w6256);
assign w6450 = v3092;
assign v3093 = ~(w6255 | w6450);
assign w6451 = v3093;
assign v3094 = ~(w6449 | w6451);
assign w6452 = v3094;
assign w6453 = w6449 & w6451;
assign v3095 = ~(w6452 | w6453);
assign w6454 = v3095;
assign v3096 = ~(w6270 | w6274);
assign w6455 = v3096;
assign w6456 = ~w6454 & w6455;
assign w6457 = w6454 & ~w6455;
assign v3097 = ~(w6456 | w6457);
assign w6458 = v3097;
assign w6459 = (~w6128 & ~w6130) | (~w6128 & w16900) | (~w6130 & w16900);
assign w6460 = ~w6458 & w6459;
assign w6461 = w6458 & ~w6459;
assign v3098 = ~(w6460 | w6461);
assign w6462 = v3098;
assign w6463 = (~w6223 & ~w6225) | (~w6223 & w17753) | (~w6225 & w17753);
assign w6464 = (~w6149 & ~w6151) | (~w6149 & w17122) | (~w6151 & w17122);
assign w6465 = (~w6080 & ~w6082) | (~w6080 & w16901) | (~w6082 & w16901);
assign v3099 = ~(w6464 | w6465);
assign w6466 = v3099;
assign w6467 = w6464 & w6465;
assign v3100 = ~(w6466 | w6467);
assign w6468 = v3100;
assign w6469 = w6463 & ~w6468;
assign w6470 = ~w6463 & w6468;
assign v3101 = ~(w6469 | w6470);
assign w6471 = v3101;
assign w6472 = (~w6203 & ~w6205) | (~w6203 & w17123) | (~w6205 & w17123);
assign w6473 = w6471 & ~w6472;
assign w6474 = ~w6471 & w6472;
assign v3102 = ~(w6473 | w6474);
assign w6475 = v3102;
assign w6476 = w6462 & w6475;
assign v3103 = ~(w6462 | w6475);
assign w6477 = v3103;
assign v3104 = ~(w6476 | w6477);
assign w6478 = v3104;
assign w6479 = ~w6442 & w6478;
assign w6480 = w6442 & ~w6478;
assign v3105 = ~(w6479 | w6480);
assign w6481 = v3105;
assign w6482 = w6441 & w6481;
assign v3106 = ~(w6441 | w6481);
assign w6483 = v3106;
assign v3107 = ~(w6482 | w6483);
assign w6484 = v3107;
assign v3108 = ~(w6109 | w6111);
assign w6485 = v3108;
assign w6486 = (~w6099 & ~w6101) | (~w6099 & w17124) | (~w6101 & w17124);
assign w6487 = (~w6119 & ~w6120) | (~w6119 & w16902) | (~w6120 & w16902);
assign w6488 = pi21 & pi35;
assign w6489 = pi05 & pi51;
assign w6490 = pi18 & pi38;
assign v3109 = ~(w6489 | w6490);
assign w6491 = v3109;
assign w6492 = w6489 & w6490;
assign v3110 = ~(w6491 | w6492);
assign w6493 = v3110;
assign w6494 = w6488 & ~w6493;
assign w6495 = ~w6488 & w6493;
assign v3111 = ~(w6494 | w6495);
assign w6496 = v3111;
assign v3112 = ~(w6487 | w6496);
assign w6497 = v3112;
assign w6498 = w6487 & w6496;
assign v3113 = ~(w6497 | w6498);
assign w6499 = v3113;
assign w6500 = w6486 & ~w6499;
assign w6501 = ~w6486 & w6499;
assign v3114 = ~(w6500 | w6501);
assign w6502 = v3114;
assign w6503 = (~w6159 & ~w6161) | (~w6159 & w17754) | (~w6161 & w17754);
assign w6504 = ~w6502 & w6503;
assign w6505 = w6502 & ~w6503;
assign v3115 = ~(w6504 | w6505);
assign w6506 = v3115;
assign w6507 = w6485 & ~w6506;
assign w6508 = ~w6485 & w6506;
assign v3116 = ~(w6507 | w6508);
assign w6509 = v3116;
assign v3117 = ~(w6135 | w6138);
assign w6510 = v3117;
assign w6511 = ~w6509 & w6510;
assign w6512 = w6509 & ~w6510;
assign v3118 = ~(w6511 | w6512);
assign w6513 = v3118;
assign v3119 = ~(w6165 | w6241);
assign w6514 = v3119;
assign w6515 = ~w6513 & w6514;
assign w6516 = w6513 & ~w6514;
assign v3120 = ~(w6515 | w6516);
assign w6517 = v3120;
assign v3121 = ~(w6141 | w6245);
assign w6518 = v3121;
assign w6519 = w6517 & ~w6518;
assign w6520 = ~w6517 & w6518;
assign v3122 = ~(w6519 | w6520);
assign w6521 = v3122;
assign w6522 = w6484 & w6521;
assign v3123 = ~(w6484 | w6521);
assign w6523 = v3123;
assign v3124 = ~(w6522 | w6523);
assign w6524 = v3124;
assign w6525 = ~w6303 & w6524;
assign w6526 = w6303 & ~w6524;
assign v3125 = ~(w6525 | w6526);
assign w6527 = v3125;
assign v3126 = ~(w6068 | w6296);
assign w6528 = v3126;
assign w6529 = ~w6298 & w6528;
assign v3127 = ~(w6295 | w6529);
assign w6530 = v3127;
assign w6531 = w6527 & w6530;
assign v3128 = ~(w6527 | w6530);
assign w6532 = v3128;
assign v3129 = ~(w6531 | w6532);
assign w6533 = v3129;
assign v3130 = ~(w6519 | w6522);
assign w6534 = v3130;
assign v3131 = ~(w6512 | w6516);
assign w6535 = v3131;
assign w6536 = (~w6418 & ~w6420) | (~w6418 & w17755) | (~w6420 & w17755);
assign w6537 = (~w6325 & ~w6327) | (~w6325 & w17125) | (~w6327 & w17125);
assign w6538 = (~w6353 & ~w6355) | (~w6353 & w16903) | (~w6355 & w16903);
assign v3132 = ~(w6537 | w6538);
assign w6539 = v3132;
assign w6540 = w6537 & w6538;
assign v3133 = ~(w6539 | w6540);
assign w6541 = v3133;
assign w6542 = w6536 & ~w6541;
assign w6543 = ~w6536 & w6541;
assign v3134 = ~(w6542 | w6543);
assign w6544 = v3134;
assign v3135 = ~(w6433 | w6436);
assign w6545 = v3135;
assign w6546 = ~w6544 & w6545;
assign w6547 = w6544 & ~w6545;
assign v3136 = ~(w6546 | w6547);
assign w6548 = v3136;
assign w6549 = (~w6386 & ~w6388) | (~w6386 & w17756) | (~w6388 & w17756);
assign v3137 = ~(w6389 | w6392);
assign w6550 = v3137;
assign v3138 = ~(w6391 | w6550);
assign w6551 = v3138;
assign v3139 = ~(w6409 | w6413);
assign w6552 = v3139;
assign v3140 = ~(w6412 | w6552);
assign w6553 = v3140;
assign w6554 = w6551 & w6553;
assign v3141 = ~(w6551 | w6553);
assign w6555 = v3141;
assign v3142 = ~(w6554 | w6555);
assign w6556 = v3142;
assign v3143 = ~(w6377 | w6381);
assign w6557 = v3143;
assign v3144 = ~(w6380 | w6557);
assign w6558 = v3144;
assign v3145 = ~(w6556 | w6558);
assign w6559 = v3145;
assign w6560 = w6556 & w6558;
assign v3146 = ~(w6559 | w6560);
assign w6561 = v3146;
assign v3147 = ~(w6400 | w6404);
assign w6562 = v3147;
assign v3148 = ~(w6403 | w6562);
assign w6563 = v3148;
assign v3149 = ~(w6356 | w6360);
assign w6564 = v3149;
assign v3150 = ~(w6359 | w6564);
assign w6565 = v3150;
assign w6566 = w6563 & w6565;
assign v3151 = ~(w6563 | w6565);
assign w6567 = v3151;
assign v3152 = ~(w6566 | w6567);
assign w6568 = v3152;
assign v3153 = ~(w6114 | w6348);
assign w6569 = v3153;
assign v3154 = ~(w6346 | w6569);
assign w6570 = v3154;
assign v3155 = ~(w6568 | w6570);
assign w6571 = v3155;
assign w6572 = w6568 & w6570;
assign v3156 = ~(w6571 | w6572);
assign w6573 = v3156;
assign w6574 = w6561 & w6573;
assign v3157 = ~(w6561 | w6573);
assign w6575 = v3157;
assign v3158 = ~(w6574 | w6575);
assign w6576 = v3158;
assign w6577 = ~w6549 & w6576;
assign w6578 = w6549 & ~w6576;
assign v3159 = ~(w6577 | w6578);
assign w6579 = v3159;
assign w6580 = w6548 & w6579;
assign v3160 = ~(w6548 | w6579);
assign w6581 = v3160;
assign v3161 = ~(w6580 | w6581);
assign w6582 = v3161;
assign w6583 = ~w6535 & w6582;
assign w6584 = w6535 & ~w6582;
assign v3162 = ~(w6583 | w6584);
assign w6585 = v3162;
assign v3163 = ~(w6505 | w6508);
assign w6586 = v3163;
assign v3164 = ~(w6421 | w6425);
assign w6587 = v3164;
assign v3165 = ~(w6424 | w6587);
assign w6588 = v3165;
assign v3166 = ~(w6488 | w6492);
assign w6589 = v3166;
assign v3167 = ~(w6491 | w6589);
assign w6590 = v3167;
assign w6591 = w6588 & w6590;
assign v3168 = ~(w6588 | w6590);
assign w6592 = v3168;
assign v3169 = ~(w6591 | w6592);
assign w6593 = v3169;
assign w6594 = w6368 & ~w6371;
assign v3170 = ~(w6372 | w6594);
assign w6595 = v3170;
assign w6596 = ~w6593 & w6595;
assign w6597 = w6593 & ~w6595;
assign v3171 = ~(w6596 | w6597);
assign w6598 = v3171;
assign w6599 = (~w6497 & ~w6499) | (~w6497 & w17126) | (~w6499 & w17126);
assign w6600 = ~w6598 & w6599;
assign w6601 = w6598 & ~w6599;
assign v3172 = ~(w6600 | w6601);
assign w6602 = v3172;
assign w6603 = pi21 & pi36;
assign w6604 = pi23 & pi34;
assign w6605 = pi22 & pi35;
assign v3173 = ~(w6604 | w6605);
assign w6606 = v3173;
assign w6607 = pi23 & pi35;
assign w6608 = w6401 & w6607;
assign v3174 = ~(w6606 | w6608);
assign w6609 = v3174;
assign w6610 = w6603 & ~w6609;
assign w6611 = ~w6603 & w6609;
assign v3175 = ~(w6610 | w6611);
assign w6612 = v3175;
assign w6613 = pi07 & pi50;
assign w6614 = pi08 & pi49;
assign w6615 = pi16 & pi41;
assign v3176 = ~(w6614 | w6615);
assign w6616 = v3176;
assign w6617 = w6614 & w6615;
assign v3177 = ~(w6616 | w6617);
assign w6618 = v3177;
assign w6619 = w6613 & ~w6618;
assign w6620 = ~w6613 & w6618;
assign v3178 = ~(w6619 | w6620);
assign w6621 = v3178;
assign v3179 = ~(w6612 | w6621);
assign w6622 = v3179;
assign w6623 = w6612 & w6621;
assign v3180 = ~(w6622 | w6623);
assign w6624 = v3180;
assign w6625 = pi24 & pi33;
assign w6626 = pi26 & pi31;
assign w6627 = pi25 & pi32;
assign v3181 = ~(w6626 | w6627);
assign w6628 = v3181;
assign w6629 = w6626 & w6627;
assign v3182 = ~(w6628 | w6629);
assign w6630 = v3182;
assign w6631 = w6625 & ~w6630;
assign w6632 = ~w6625 & w6630;
assign v3183 = ~(w6631 | w6632);
assign w6633 = v3183;
assign w6634 = w6624 & ~w6633;
assign w6635 = ~w6624 & w6633;
assign v3184 = ~(w6634 | w6635);
assign w6636 = v3184;
assign w6637 = w6602 & w6636;
assign v3185 = ~(w6602 | w6636);
assign w6638 = v3185;
assign v3186 = ~(w6637 | w6638);
assign w6639 = v3186;
assign w6640 = ~w6586 & w6639;
assign w6641 = w6586 & ~w6639;
assign v3187 = ~(w6640 | w6641);
assign w6642 = v3187;
assign w6643 = (~w6466 & ~w6468) | (~w6466 & w17127) | (~w6468 & w17127);
assign w6644 = pi05 & pi52;
assign w6645 = pi20 & pi37;
assign w6646 = pi19 & pi38;
assign v3188 = ~(w6645 | w6646);
assign w6647 = v3188;
assign w6648 = pi20 & pi38;
assign w6649 = w6357 & w6648;
assign v3189 = ~(w6647 | w6649);
assign w6650 = v3189;
assign w6651 = w6644 & ~w6650;
assign w6652 = ~w6644 & w6650;
assign v3190 = ~(w6651 | w6652);
assign w6653 = v3190;
assign w6654 = pi03 & pi54;
assign w6655 = pi04 & pi53;
assign w6656 = pi02 & pi55;
assign v3191 = ~(w6655 | w6656);
assign w6657 = v3191;
assign w6658 = w6655 & w6656;
assign v3192 = ~(w6657 | w6658);
assign w6659 = v3192;
assign w6660 = w6654 & ~w6659;
assign w6661 = ~w6654 & w6659;
assign v3193 = ~(w6660 | w6661);
assign w6662 = v3193;
assign v3194 = ~(w6653 | w6662);
assign w6663 = v3194;
assign w6664 = w6653 & w6662;
assign v3195 = ~(w6663 | w6664);
assign w6665 = v3195;
assign w6666 = pi15 & pi42;
assign w6667 = pi10 & pi47;
assign w6668 = pi09 & pi48;
assign v3196 = ~(w6667 | w6668);
assign w6669 = v3196;
assign w6670 = pi10 & pi48;
assign w6671 = w6421 & w6670;
assign v3197 = ~(w6669 | w6671);
assign w6672 = v3197;
assign w6673 = w6666 & ~w6672;
assign w6674 = ~w6666 & w6672;
assign v3198 = ~(w6673 | w6674);
assign w6675 = v3198;
assign w6676 = w6665 & ~w6675;
assign w6677 = ~w6665 & w6675;
assign v3199 = ~(w6676 | w6677);
assign w6678 = v3199;
assign w6679 = pi14 & pi43;
assign w6680 = pi11 & pi46;
assign v3200 = ~(w6173 | w6680);
assign w6681 = v3200;
assign w6682 = pi13 & pi46;
assign w6683 = w6171 & w6682;
assign v3201 = ~(w6681 | w6683);
assign w6684 = v3201;
assign w6685 = w6679 & ~w6684;
assign w6686 = ~w6679 & w6684;
assign v3202 = ~(w6685 | w6686);
assign w6687 = v3202;
assign w6688 = pi12 & pi45;
assign w6689 = pi28 & pi29;
assign w6690 = pi27 & pi30;
assign v3203 = ~(w6689 | w6690);
assign w6691 = v3203;
assign w6692 = w6689 & w6690;
assign v3204 = ~(w6691 | w6692);
assign w6693 = v3204;
assign w6694 = w6688 & ~w6693;
assign w6695 = ~w6688 & w6693;
assign v3205 = ~(w6694 | w6695);
assign w6696 = v3205;
assign v3206 = ~(w6687 | w6696);
assign w6697 = v3206;
assign w6698 = w6687 & w6696;
assign v3207 = ~(w6697 | w6698);
assign w6699 = v3207;
assign w6700 = pi18 & pi39;
assign w6701 = pi06 & pi51;
assign w6702 = pi17 & pi40;
assign v3208 = ~(w6701 | w6702);
assign w6703 = v3208;
assign w6704 = w6701 & w6702;
assign v3209 = ~(w6703 | w6704);
assign w6705 = v3209;
assign w6706 = w6700 & ~w6705;
assign w6707 = ~w6700 & w6705;
assign v3210 = ~(w6706 | w6707);
assign w6708 = v3210;
assign w6709 = w6699 & ~w6708;
assign w6710 = ~w6699 & w6708;
assign v3211 = ~(w6709 | w6710);
assign w6711 = v3211;
assign w6712 = w6678 & w6711;
assign v3212 = ~(w6678 | w6711);
assign w6713 = v3212;
assign v3213 = ~(w6712 | w6713);
assign w6714 = v3213;
assign w6715 = ~w6643 & w6714;
assign w6716 = w6643 & ~w6714;
assign v3214 = ~(w6715 | w6716);
assign w6717 = v3214;
assign w6718 = w6642 & w6717;
assign v3215 = ~(w6642 | w6717);
assign w6719 = v3215;
assign v3216 = ~(w6718 | w6719);
assign w6720 = v3216;
assign v3217 = ~(w6585 | w6720);
assign w6721 = v3217;
assign w6722 = w6585 & w6720;
assign v3218 = ~(w6721 | w6722);
assign w6723 = v3218;
assign v3219 = ~(w6479 | w6482);
assign w6724 = v3219;
assign v3220 = ~(w6339 | w6440);
assign w6725 = v3220;
assign v3221 = ~(w6473 | w6476);
assign w6726 = v3221;
assign w6727 = (~w6447 & ~w6449) | (~w6447 & w17128) | (~w6449 & w17128);
assign w6728 = (~w6309 & ~w6311) | (~w6309 & w16749) | (~w6311 & w16749);
assign w6729 = pi00 & pi57;
assign w6730 = w6321 & w6729;
assign v3222 = ~(w6321 | w6729);
assign w6731 = v3222;
assign v3223 = ~(w6730 | w6731);
assign w6732 = v3223;
assign w6733 = pi01 & pi56;
assign w6734 = pi29 & w6733;
assign v3224 = ~(pi29 | w6733);
assign w6735 = v3224;
assign v3225 = ~(w6734 | w6735);
assign w6736 = v3225;
assign w6737 = w6732 & w6736;
assign v3226 = ~(w6732 | w6736);
assign w6738 = v3226;
assign v3227 = ~(w6737 | w6738);
assign w6739 = v3227;
assign w6740 = ~w6728 & w6739;
assign w6741 = w6728 & ~w6739;
assign v3228 = ~(w6740 | w6741);
assign w6742 = v3228;
assign w6743 = w6727 & ~w6742;
assign w6744 = ~w6727 & w6742;
assign v3229 = ~(w6743 | w6744);
assign w6745 = v3229;
assign w6746 = (~w6457 & ~w6458) | (~w6457 & w16904) | (~w6458 & w16904);
assign w6747 = (~w6333 & ~w6335) | (~w6333 & w17129) | (~w6335 & w17129);
assign v3230 = ~(w6746 | w6747);
assign w6748 = v3230;
assign w6749 = w6746 & w6747;
assign v3231 = ~(w6748 | w6749);
assign w6750 = v3231;
assign w6751 = w6745 & w6750;
assign v3232 = ~(w6745 | w6750);
assign w6752 = v3232;
assign v3233 = ~(w6751 | w6752);
assign w6753 = v3233;
assign w6754 = ~w6726 & w6753;
assign w6755 = w6726 & ~w6753;
assign v3234 = ~(w6754 | w6755);
assign w6756 = v3234;
assign w6757 = ~w6725 & w6756;
assign w6758 = w6725 & ~w6756;
assign v3235 = ~(w6757 | w6758);
assign w6759 = v3235;
assign w6760 = ~w6724 & w6759;
assign w6761 = w6724 & ~w6759;
assign v3236 = ~(w6760 | w6761);
assign w6762 = v3236;
assign w6763 = w6723 & w6762;
assign v3237 = ~(w6723 | w6762);
assign w6764 = v3237;
assign v3238 = ~(w6763 | w6764);
assign w6765 = v3238;
assign w6766 = ~w6534 & w6765;
assign w6767 = w6534 & ~w6765;
assign v3239 = ~(w6766 | w6767);
assign w6768 = v3239;
assign v3240 = ~(w6295 | w6525);
assign w6769 = v3240;
assign w6770 = (~w6298 & w16539) | (~w6298 & w16540) | (w16539 & w16540);
assign w6771 = w6768 & w6770;
assign v3241 = ~(w6768 | w6770);
assign w6772 = v3241;
assign v3242 = ~(w6771 | w6772);
assign w6773 = v3242;
assign v3243 = ~(w6760 | w6763);
assign w6774 = v3243;
assign v3244 = ~(w6583 | w6722);
assign w6775 = v3244;
assign v3245 = ~(w6547 | w6580);
assign w6776 = v3245;
assign w6777 = (~w6601 & ~w6602) | (~w6601 & w17757) | (~w6602 & w17757);
assign w6778 = (~w6554 & ~w6556) | (~w6554 & w17130) | (~w6556 & w17130);
assign w6779 = (~w6591 & ~w6593) | (~w6591 & w16750) | (~w6593 & w16750);
assign w6780 = (~w6566 & ~w6568) | (~w6566 & w16751) | (~w6568 & w16751);
assign v3246 = ~(w6779 | w6780);
assign w6781 = v3246;
assign w6782 = w6779 & w6780;
assign v3247 = ~(w6781 | w6782);
assign w6783 = v3247;
assign w6784 = w6778 & ~w6783;
assign w6785 = ~w6778 & w6783;
assign v3248 = ~(w6784 | w6785);
assign w6786 = v3248;
assign w6787 = (~w6574 & ~w6576) | (~w6574 & w17131) | (~w6576 & w17131);
assign w6788 = ~w6786 & w6787;
assign w6789 = w6786 & ~w6787;
assign v3249 = ~(w6788 | w6789);
assign w6790 = v3249;
assign w6791 = ~w6777 & w6790;
assign w6792 = w6777 & ~w6790;
assign v3250 = ~(w6791 | w6792);
assign w6793 = v3250;
assign w6794 = ~w6776 & w6793;
assign w6795 = w6776 & ~w6793;
assign v3251 = ~(w6794 | w6795);
assign w6796 = v3251;
assign v3252 = ~(w6640 | w6718);
assign w6797 = v3252;
assign w6798 = w6796 & ~w6797;
assign w6799 = ~w6796 & w6797;
assign v3253 = ~(w6798 | w6799);
assign w6800 = v3253;
assign w6801 = ~w6775 & w6800;
assign w6802 = w6775 & ~w6800;
assign v3254 = ~(w6801 | w6802);
assign w6803 = v3254;
assign v3255 = ~(w6754 | w6757);
assign w6804 = v3255;
assign v3256 = ~(w6712 | w6715);
assign w6805 = v3256;
assign w6806 = (~w6697 & ~w6699) | (~w6697 & w17758) | (~w6699 & w17758);
assign w6807 = (~w6663 & ~w6665) | (~w6663 & w16905) | (~w6665 & w16905);
assign w6808 = pi28 & pi30;
assign w6809 = pi01 & pi57;
assign v3257 = ~(w6808 | w6809);
assign w6810 = v3257;
assign w6811 = w6808 & w6809;
assign v3258 = ~(w6810 | w6811);
assign w6812 = v3258;
assign w6813 = w6734 & w6812;
assign v3259 = ~(w6734 | w6812);
assign w6814 = v3259;
assign v3260 = ~(w6813 | w6814);
assign w6815 = v3260;
assign v3261 = ~(w6688 | w6692);
assign w6816 = v3261;
assign v3262 = ~(w6691 | w6816);
assign w6817 = v3262;
assign w6818 = w6815 & w6817;
assign v3263 = ~(w6815 | w6817);
assign w6819 = v3263;
assign v3264 = ~(w6818 | w6819);
assign w6820 = v3264;
assign w6821 = ~w6807 & w6820;
assign w6822 = w6807 & ~w6820;
assign v3265 = ~(w6821 | w6822);
assign w6823 = v3265;
assign w6824 = ~w6806 & w6823;
assign w6825 = w6806 & ~w6823;
assign v3266 = ~(w6824 | w6825);
assign w6826 = v3266;
assign w6827 = ~w6805 & w6826;
assign w6828 = w6805 & ~w6826;
assign v3267 = ~(w6827 | w6828);
assign w6829 = v3267;
assign w6830 = (~w6622 & ~w6624) | (~w6622 & w17759) | (~w6624 & w17759);
assign v3268 = ~(w6625 | w6629);
assign w6831 = v3268;
assign v3269 = ~(w6628 | w6831);
assign w6832 = v3269;
assign w6833 = w6666 & ~w6669;
assign v3270 = ~(w6671 | w6833);
assign w6834 = v3270;
assign w6835 = w6832 & ~w6834;
assign w6836 = ~w6832 & w6834;
assign v3271 = ~(w6835 | w6836);
assign w6837 = v3271;
assign w6838 = w6603 & ~w6606;
assign v3272 = ~(w6608 | w6838);
assign w6839 = v3272;
assign w6840 = ~w6837 & w6839;
assign w6841 = w6837 & ~w6839;
assign v3273 = ~(w6840 | w6841);
assign w6842 = v3273;
assign v3274 = ~(w6654 | w6658);
assign w6843 = v3274;
assign v3275 = ~(w6657 | w6843);
assign w6844 = v3275;
assign w6845 = w6644 & ~w6647;
assign v3276 = ~(w6649 | w6845);
assign w6846 = v3276;
assign w6847 = w6844 & ~w6846;
assign w6848 = ~w6844 & w6846;
assign v3277 = ~(w6847 | w6848);
assign w6849 = v3277;
assign w6850 = w6679 & ~w6681;
assign v3278 = ~(w6683 | w6850);
assign w6851 = v3278;
assign w6852 = ~w6849 & w6851;
assign w6853 = w6849 & ~w6851;
assign v3279 = ~(w6852 | w6853);
assign w6854 = v3279;
assign w6855 = w6842 & w6854;
assign v3280 = ~(w6842 | w6854);
assign w6856 = v3280;
assign v3281 = ~(w6855 | w6856);
assign w6857 = v3281;
assign w6858 = ~w6830 & w6857;
assign w6859 = w6830 & ~w6857;
assign v3282 = ~(w6858 | w6859);
assign w6860 = v3282;
assign w6861 = w6829 & w6860;
assign v3283 = ~(w6829 | w6860);
assign w6862 = v3283;
assign v3284 = ~(w6861 | w6862);
assign w6863 = v3284;
assign w6864 = ~w6804 & w6863;
assign w6865 = w6804 & ~w6863;
assign v3285 = ~(w6864 | w6865);
assign w6866 = v3285;
assign w6867 = (~w6748 & ~w6750) | (~w6748 & w17132) | (~w6750 & w17132);
assign w6868 = (~w6730 & ~w6732) | (~w6730 & w17133) | (~w6732 & w17133);
assign v3286 = ~(w6613 | w6617);
assign w6869 = v3286;
assign v3287 = ~(w6616 | w6869);
assign w6870 = v3287;
assign v3288 = ~(w6700 | w6704);
assign w6871 = v3288;
assign v3289 = ~(w6703 | w6871);
assign w6872 = v3289;
assign w6873 = w6870 & w6872;
assign v3290 = ~(w6870 | w6872);
assign w6874 = v3290;
assign v3291 = ~(w6873 | w6874);
assign w6875 = v3291;
assign w6876 = w6868 & ~w6875;
assign w6877 = ~w6868 & w6875;
assign v3292 = ~(w6876 | w6877);
assign w6878 = v3292;
assign w6879 = (~w6740 & ~w6742) | (~w6740 & w16906) | (~w6742 & w16906);
assign w6880 = ~w6878 & w6879;
assign w6881 = w6878 & ~w6879;
assign v3293 = ~(w6880 | w6881);
assign w6882 = v3293;
assign w6883 = pi14 & pi44;
assign w6884 = pi13 & pi45;
assign w6885 = pi12 & pi46;
assign v3294 = ~(w6884 | w6885);
assign w6886 = v3294;
assign w6887 = w6682 & w6688;
assign v3295 = ~(w6886 | w6887);
assign w6888 = v3295;
assign w6889 = w6883 & ~w6888;
assign w6890 = ~w6883 & w6888;
assign v3296 = ~(w6889 | w6890);
assign w6891 = v3296;
assign w6892 = pi15 & pi43;
assign w6893 = pi11 & pi47;
assign v3297 = ~(w6892 | w6893);
assign w6894 = v3297;
assign w6895 = w6892 & w6893;
assign v3298 = ~(w6894 | w6895);
assign w6896 = v3298;
assign w6897 = w6670 & ~w6896;
assign w6898 = ~w6670 & w6896;
assign v3299 = ~(w6897 | w6898);
assign w6899 = v3299;
assign v3300 = ~(w6891 | w6899);
assign w6900 = v3300;
assign w6901 = w6891 & w6899;
assign v3301 = ~(w6900 | w6901);
assign w6902 = v3301;
assign w6903 = pi03 & pi55;
assign w6904 = pi19 & pi39;
assign w6905 = pi06 & pi52;
assign v3302 = ~(w6904 | w6905);
assign w6906 = v3302;
assign w6907 = w6904 & w6905;
assign v3303 = ~(w6906 | w6907);
assign w6908 = v3303;
assign w6909 = w6903 & ~w6908;
assign w6910 = ~w6903 & w6908;
assign v3304 = ~(w6909 | w6910);
assign w6911 = v3304;
assign w6912 = w6902 & ~w6911;
assign w6913 = ~w6902 & w6911;
assign v3305 = ~(w6912 | w6913);
assign w6914 = v3305;
assign v3306 = ~(w6882 | w6914);
assign w6915 = v3306;
assign w6916 = w6882 & w6914;
assign v3307 = ~(w6915 | w6916);
assign w6917 = v3307;
assign w6918 = ~w6867 & w6917;
assign w6919 = w6867 & ~w6917;
assign v3308 = ~(w6918 | w6919);
assign w6920 = v3308;
assign w6921 = (~w6539 & ~w6541) | (~w6539 & w17134) | (~w6541 & w17134);
assign w6922 = pi05 & pi53;
assign w6923 = pi21 & pi37;
assign v3309 = ~(w6648 | w6923);
assign w6924 = v3309;
assign w6925 = pi21 & pi38;
assign w6926 = w6645 & w6925;
assign v3310 = ~(w6924 | w6926);
assign w6927 = v3310;
assign w6928 = w6922 & ~w6927;
assign w6929 = ~w6922 & w6927;
assign v3311 = ~(w6928 | w6929);
assign w6930 = v3311;
assign w6931 = pi00 & pi58;
assign w6932 = pi04 & pi54;
assign v3312 = ~(w6931 | w6932);
assign w6933 = v3312;
assign w6934 = w6931 & w6932;
assign v3313 = ~(w6933 | w6934);
assign w6935 = v3313;
assign w6936 = w6347 & ~w6935;
assign w6937 = ~w6347 & w6935;
assign v3314 = ~(w6936 | w6937);
assign w6938 = v3314;
assign v3315 = ~(w6930 | w6938);
assign w6939 = v3315;
assign w6940 = w6930 & w6938;
assign v3316 = ~(w6939 | w6940);
assign w6941 = v3316;
assign w6942 = pi17 & pi41;
assign w6943 = pi09 & pi49;
assign w6944 = pi16 & pi42;
assign v3317 = ~(w6943 | w6944);
assign w6945 = v3317;
assign w6946 = w6943 & w6944;
assign v3318 = ~(w6945 | w6946);
assign w6947 = v3318;
assign w6948 = w6942 & ~w6947;
assign w6949 = ~w6942 & w6947;
assign v3319 = ~(w6948 | w6949);
assign w6950 = v3319;
assign w6951 = w6941 & ~w6950;
assign w6952 = ~w6941 & w6950;
assign v3320 = ~(w6951 | w6952);
assign w6953 = v3320;
assign w6954 = pi18 & pi40;
assign w6955 = pi07 & pi51;
assign w6956 = pi08 & pi50;
assign v3321 = ~(w6955 | w6956);
assign w6957 = v3321;
assign w6958 = pi08 & pi51;
assign w6959 = w6613 & w6958;
assign v3322 = ~(w6957 | w6959);
assign w6960 = v3322;
assign w6961 = w6954 & ~w6960;
assign w6962 = ~w6954 & w6960;
assign v3323 = ~(w6961 | w6962);
assign w6963 = v3323;
assign w6964 = pi22 & pi36;
assign w6965 = pi24 & pi34;
assign v3324 = ~(w6607 | w6965);
assign w6966 = v3324;
assign w6967 = pi24 & pi35;
assign w6968 = w6604 & w6967;
assign v3325 = ~(w6966 | w6968);
assign w6969 = v3325;
assign w6970 = w6964 & ~w6969;
assign w6971 = ~w6964 & w6969;
assign v3326 = ~(w6970 | w6971);
assign w6972 = v3326;
assign v3327 = ~(w6963 | w6972);
assign w6973 = v3327;
assign w6974 = w6963 & w6972;
assign v3328 = ~(w6973 | w6974);
assign w6975 = v3328;
assign w6976 = pi25 & pi33;
assign w6977 = pi26 & pi32;
assign w6978 = pi27 & pi31;
assign v3329 = ~(w6977 | w6978);
assign w6979 = v3329;
assign w6980 = w6977 & w6978;
assign v3330 = ~(w6979 | w6980);
assign w6981 = v3330;
assign w6982 = w6976 & ~w6981;
assign w6983 = ~w6976 & w6981;
assign v3331 = ~(w6982 | w6983);
assign w6984 = v3331;
assign w6985 = w6975 & ~w6984;
assign w6986 = ~w6975 & w6984;
assign v3332 = ~(w6985 | w6986);
assign w6987 = v3332;
assign w6988 = w6953 & w6987;
assign v3333 = ~(w6953 | w6987);
assign w6989 = v3333;
assign v3334 = ~(w6988 | w6989);
assign w6990 = v3334;
assign w6991 = ~w6921 & w6990;
assign w6992 = w6921 & ~w6990;
assign v3335 = ~(w6991 | w6992);
assign w6993 = v3335;
assign v3336 = ~(w6920 | w6993);
assign w6994 = v3336;
assign w6995 = w6920 & w6993;
assign v3337 = ~(w6994 | w6995);
assign w6996 = v3337;
assign v3338 = ~(w6866 | w6996);
assign w6997 = v3338;
assign w6998 = w6866 & w6996;
assign v3339 = ~(w6997 | w6998);
assign w6999 = v3339;
assign v3340 = ~(w6803 | w6999);
assign w7000 = v3340;
assign w7001 = w6803 & w6999;
assign v3341 = ~(w7000 | w7001);
assign w7002 = v3341;
assign w7003 = ~w6774 & w7002;
assign w7004 = w6774 & ~w7002;
assign v3342 = ~(w7003 | w7004);
assign w7005 = v3342;
assign w7006 = (w6298 & w16541) | (w6298 & w16542) | (w16541 & w16542);
assign v3343 = ~(w6767 | w7006);
assign w7007 = v3343;
assign w7008 = w7005 & w7007;
assign v3344 = ~(w7005 | w7007);
assign w7009 = v3344;
assign v3345 = ~(w7008 | w7009);
assign w7010 = v3345;
assign v3346 = ~(w6864 | w6998);
assign w7011 = v3346;
assign w7012 = (~w6918 & ~w6920) | (~w6918 & w17760) | (~w6920 & w17760);
assign w7013 = (~w6827 & ~w6829) | (~w6827 & w17761) | (~w6829 & w17761);
assign w7014 = (~w6881 & ~w6882) | (~w6881 & w17135) | (~w6882 & w17135);
assign w7015 = (~w6835 & ~w6837) | (~w6835 & w17762) | (~w6837 & w17762);
assign w7016 = (~w6873 & ~w6875) | (~w6873 & w17136) | (~w6875 & w17136);
assign w7017 = (~w6847 & ~w6849) | (~w6847 & w17137) | (~w6849 & w17137);
assign v3347 = ~(w7016 | w7017);
assign w7018 = v3347;
assign w7019 = w7016 & w7017;
assign v3348 = ~(w7018 | w7019);
assign w7020 = v3348;
assign w7021 = w7015 & ~w7020;
assign w7022 = ~w7015 & w7020;
assign v3349 = ~(w7021 | w7022);
assign w7023 = v3349;
assign w7024 = (~w6855 & ~w6857) | (~w6855 & w17138) | (~w6857 & w17138);
assign w7025 = ~w7023 & w7024;
assign w7026 = w7023 & ~w7024;
assign v3350 = ~(w7025 | w7026);
assign w7027 = v3350;
assign w7028 = ~w7014 & w7027;
assign w7029 = w7014 & ~w7027;
assign v3351 = ~(w7028 | w7029);
assign w7030 = v3351;
assign w7031 = ~w7013 & w7030;
assign w7032 = w7013 & ~w7030;
assign v3352 = ~(w7031 | w7032);
assign w7033 = v3352;
assign w7034 = ~w7012 & w7033;
assign w7035 = w7012 & ~w7033;
assign v3353 = ~(w7034 | w7035);
assign w7036 = v3353;
assign w7037 = ~w7011 & w7036;
assign w7038 = w7011 & ~w7036;
assign v3354 = ~(w7037 | w7038);
assign w7039 = v3354;
assign v3355 = ~(w6794 | w6798);
assign w7040 = v3355;
assign w7041 = (~w6939 & ~w6941) | (~w6939 & w17763) | (~w6941 & w17763);
assign w7042 = (~w6900 & ~w6902) | (~w6900 & w16907) | (~w6902 & w16907);
assign w7043 = (~w6973 & ~w6975) | (~w6973 & w16908) | (~w6975 & w16908);
assign v3356 = ~(w7042 | w7043);
assign w7044 = v3356;
assign w7045 = w7042 & w7043;
assign v3357 = ~(w7044 | w7045);
assign w7046 = v3357;
assign w7047 = w7041 & ~w7046;
assign w7048 = ~w7041 & w7046;
assign v3358 = ~(w7047 | w7048);
assign w7049 = v3358;
assign v3359 = ~(w6988 | w6991);
assign w7050 = v3359;
assign v3360 = ~(w6347 | w6934);
assign w7051 = v3360;
assign v3361 = ~(w6933 | w7051);
assign w7052 = v3361;
assign v3362 = ~(w6903 | w6907);
assign w7053 = v3362;
assign v3363 = ~(w6906 | w7053);
assign w7054 = v3363;
assign w7055 = w7052 & w7054;
assign v3364 = ~(w7052 | w7054);
assign w7056 = v3364;
assign v3365 = ~(w7055 | w7056);
assign w7057 = v3365;
assign v3366 = ~(w6942 | w6946);
assign w7058 = v3366;
assign v3367 = ~(w6945 | w7058);
assign w7059 = v3367;
assign v3368 = ~(w7057 | w7059);
assign w7060 = v3368;
assign w7061 = w7057 & w7059;
assign v3369 = ~(w7060 | w7061);
assign w7062 = v3369;
assign w7063 = w6922 & ~w6924;
assign v3370 = ~(w6926 | w7063);
assign w7064 = v3370;
assign w7065 = w6964 & ~w6966;
assign v3371 = ~(w6968 | w7065);
assign w7066 = v3371;
assign v3372 = ~(w7064 | w7066);
assign w7067 = v3372;
assign w7068 = w7064 & w7066;
assign v3373 = ~(w7067 | w7068);
assign w7069 = v3373;
assign w7070 = w6954 & ~w6957;
assign v3374 = ~(w6959 | w7070);
assign w7071 = v3374;
assign w7072 = ~w7069 & w7071;
assign w7073 = w7069 & ~w7071;
assign v3375 = ~(w7072 | w7073);
assign w7074 = v3375;
assign w7075 = pi58 & w1939;
assign w7076 = pi01 & pi58;
assign v3376 = ~(pi30 | w7076);
assign w7077 = v3376;
assign v3377 = ~(w7075 | w7077);
assign w7078 = v3377;
assign w7079 = w6883 & ~w6886;
assign v3378 = ~(w6887 | w7079);
assign w7080 = v3378;
assign w7081 = w7078 & ~w7080;
assign w7082 = ~w7078 & w7080;
assign v3379 = ~(w7081 | w7082);
assign w7083 = v3379;
assign v3380 = ~(w6670 | w6895);
assign w7084 = v3380;
assign v3381 = ~(w6894 | w7084);
assign w7085 = v3381;
assign w7086 = w7083 & w7085;
assign v3382 = ~(w7083 | w7085);
assign w7087 = v3382;
assign v3383 = ~(w7086 | w7087);
assign w7088 = v3383;
assign w7089 = w7074 & w7088;
assign v3384 = ~(w7074 | w7088);
assign w7090 = v3384;
assign v3385 = ~(w7089 | w7090);
assign w7091 = v3385;
assign w7092 = w7062 & w7091;
assign v3386 = ~(w7062 | w7091);
assign w7093 = v3386;
assign v3387 = ~(w7092 | w7093);
assign w7094 = v3387;
assign w7095 = ~w7050 & w7094;
assign w7096 = w7050 & ~w7094;
assign v3388 = ~(w7095 | w7096);
assign w7097 = v3388;
assign w7098 = w7049 & w7097;
assign v3389 = ~(w7049 | w7097);
assign w7099 = v3389;
assign v3390 = ~(w7098 | w7099);
assign w7100 = v3390;
assign w7101 = ~w7040 & w7100;
assign w7102 = w7040 & ~w7100;
assign v3391 = ~(w7101 | w7102);
assign w7103 = v3391;
assign w7104 = (~w6789 & ~w6790) | (~w6789 & w17764) | (~w6790 & w17764);
assign w7105 = (~w6821 & ~w6823) | (~w6821 & w17139) | (~w6823 & w17139);
assign w7106 = pi29 & pi30;
assign w7107 = pi28 & pi31;
assign v3392 = ~(w7106 | w7107);
assign w7108 = v3392;
assign w7109 = w7106 & w7107;
assign v3393 = ~(w7108 | w7109);
assign w7110 = v3393;
assign w7111 = w6682 & ~w7110;
assign w7112 = ~w6682 & w7110;
assign v3394 = ~(w7111 | w7112);
assign w7113 = v3394;
assign w7114 = pi11 & pi48;
assign w7115 = pi14 & pi45;
assign w7116 = pi12 & pi47;
assign v3395 = ~(w7115 | w7116);
assign w7117 = v3395;
assign w7118 = w7115 & w7116;
assign v3396 = ~(w7117 | w7118);
assign w7119 = v3396;
assign w7120 = w7114 & ~w7119;
assign w7121 = ~w7114 & w7119;
assign v3397 = ~(w7120 | w7121);
assign w7122 = v3397;
assign v3398 = ~(w7113 | w7122);
assign w7123 = v3398;
assign w7124 = w7113 & w7122;
assign v3399 = ~(w7123 | w7124);
assign w7125 = v3399;
assign w7126 = pi16 & pi43;
assign w7127 = pi17 & pi42;
assign v3400 = ~(w7126 | w7127);
assign w7128 = v3400;
assign w7129 = pi17 & pi43;
assign w7130 = w6944 & w7129;
assign v3401 = ~(w7128 | w7130);
assign w7131 = v3401;
assign w7132 = w6958 & ~w7131;
assign w7133 = ~w6958 & w7131;
assign v3402 = ~(w7132 | w7133);
assign w7134 = v3402;
assign w7135 = w7125 & ~w7134;
assign w7136 = ~w7125 & w7134;
assign v3403 = ~(w7135 | w7136);
assign w7137 = v3403;
assign v3404 = ~(w6976 | w6980);
assign w7138 = v3404;
assign v3405 = ~(w6979 | w7138);
assign w7139 = v3405;
assign w7140 = pi02 & pi57;
assign w7141 = pi03 & pi56;
assign v3406 = ~(w7140 | w7141);
assign w7142 = v3406;
assign w7143 = pi03 & pi57;
assign w7144 = w6347 & w7143;
assign v3407 = ~(w7142 | w7144);
assign w7145 = v3407;
assign w7146 = w6811 & ~w7145;
assign w7147 = ~w6811 & w7145;
assign v3408 = ~(w7146 | w7147);
assign w7148 = v3408;
assign w7149 = w7139 & ~w7148;
assign w7150 = ~w7139 & w7148;
assign v3409 = ~(w7149 | w7150);
assign w7151 = v3409;
assign w7152 = pi04 & pi55;
assign w7153 = pi05 & pi54;
assign w7154 = pi19 & pi40;
assign v3410 = ~(w7153 | w7154);
assign w7155 = v3410;
assign w7156 = w7153 & w7154;
assign v3411 = ~(w7155 | w7156);
assign w7157 = v3411;
assign w7158 = w7152 & ~w7157;
assign w7159 = ~w7152 & w7157;
assign v3412 = ~(w7158 | w7159);
assign w7160 = v3412;
assign w7161 = w7151 & ~w7160;
assign w7162 = ~w7151 & w7160;
assign v3413 = ~(w7161 | w7162);
assign w7163 = v3413;
assign w7164 = w7137 & w7163;
assign v3414 = ~(w7137 | w7163);
assign w7165 = v3414;
assign v3415 = ~(w7164 | w7165);
assign w7166 = v3415;
assign w7167 = ~w7105 & w7166;
assign w7168 = w7105 & ~w7166;
assign v3416 = ~(w7167 | w7168);
assign w7169 = v3416;
assign w7170 = ~w7104 & w7169;
assign w7171 = w7104 & ~w7169;
assign v3417 = ~(w7170 | w7171);
assign w7172 = v3417;
assign v3418 = ~(w6813 | w6818);
assign w7173 = v3418;
assign w7174 = pi06 & pi53;
assign w7175 = pi07 & pi52;
assign w7176 = pi18 & pi41;
assign v3419 = ~(w7175 | w7176);
assign w7177 = v3419;
assign w7178 = w7175 & w7176;
assign v3420 = ~(w7177 | w7178);
assign w7179 = v3420;
assign w7180 = w7174 & ~w7179;
assign w7181 = ~w7174 & w7179;
assign v3421 = ~(w7180 | w7181);
assign w7182 = v3421;
assign w7183 = pi09 & pi50;
assign w7184 = pi15 & pi44;
assign w7185 = pi10 & pi49;
assign v3422 = ~(w7184 | w7185);
assign w7186 = v3422;
assign w7187 = w7184 & w7185;
assign v3423 = ~(w7186 | w7187);
assign w7188 = v3423;
assign w7189 = w7183 & ~w7188;
assign w7190 = ~w7183 & w7188;
assign v3424 = ~(w7189 | w7190);
assign w7191 = v3424;
assign v3425 = ~(w7182 | w7191);
assign w7192 = v3425;
assign w7193 = w7182 & w7191;
assign v3426 = ~(w7192 | w7193);
assign w7194 = v3426;
assign w7195 = w7173 & ~w7194;
assign w7196 = ~w7173 & w7194;
assign v3427 = ~(w7195 | w7196);
assign w7197 = v3427;
assign w7198 = (~w6781 & ~w6783) | (~w6781 & w16909) | (~w6783 & w16909);
assign w7199 = ~w7197 & w7198;
assign w7200 = w7197 & ~w7198;
assign v3428 = ~(w7199 | w7200);
assign w7201 = v3428;
assign w7202 = pi20 & pi39;
assign w7203 = pi22 & pi37;
assign v3429 = ~(w6925 | w7203);
assign w7204 = v3429;
assign w7205 = pi22 & pi38;
assign w7206 = w6923 & w7205;
assign v3430 = ~(w7204 | w7206);
assign w7207 = v3430;
assign w7208 = w7202 & ~w7207;
assign w7209 = ~w7202 & w7207;
assign v3431 = ~(w7208 | w7209);
assign w7210 = v3431;
assign w7211 = pi23 & pi36;
assign w7212 = pi25 & pi34;
assign v3432 = ~(w6967 | w7212);
assign w7213 = v3432;
assign w7214 = pi25 & pi35;
assign w7215 = w6965 & w7214;
assign v3433 = ~(w7213 | w7215);
assign w7216 = v3433;
assign w7217 = w7211 & ~w7216;
assign w7218 = ~w7211 & w7216;
assign v3434 = ~(w7217 | w7218);
assign w7219 = v3434;
assign v3435 = ~(w7210 | w7219);
assign w7220 = v3435;
assign w7221 = w7210 & w7219;
assign v3436 = ~(w7220 | w7221);
assign w7222 = v3436;
assign w7223 = pi26 & pi33;
assign w7224 = pi27 & pi32;
assign w7225 = pi00 & pi59;
assign v3437 = ~(w7224 | w7225);
assign w7226 = v3437;
assign w7227 = w7224 & w7225;
assign v3438 = ~(w7226 | w7227);
assign w7228 = v3438;
assign w7229 = w7223 & ~w7228;
assign w7230 = ~w7223 & w7228;
assign v3439 = ~(w7229 | w7230);
assign w7231 = v3439;
assign w7232 = w7222 & ~w7231;
assign w7233 = ~w7222 & w7231;
assign v3440 = ~(w7232 | w7233);
assign w7234 = v3440;
assign w7235 = w7201 & w7234;
assign v3441 = ~(w7201 | w7234);
assign w7236 = v3441;
assign v3442 = ~(w7235 | w7236);
assign w7237 = v3442;
assign w7238 = w7172 & w7237;
assign v3443 = ~(w7172 | w7237);
assign w7239 = v3443;
assign v3444 = ~(w7238 | w7239);
assign w7240 = v3444;
assign w7241 = w7103 & w7240;
assign v3445 = ~(w7103 | w7240);
assign w7242 = v3445;
assign v3446 = ~(w7241 | w7242);
assign w7243 = v3446;
assign w7244 = w7039 & w7243;
assign v3447 = ~(w7039 | w7243);
assign w7245 = v3447;
assign v3448 = ~(w7244 | w7245);
assign w7246 = v3448;
assign v3449 = ~(w6801 | w7001);
assign w7247 = v3449;
assign w7248 = ~w7246 & w7247;
assign w7249 = w7246 & ~w7247;
assign v3450 = ~(w7248 | w7249);
assign w7250 = v3450;
assign v3451 = ~(w6767 | w7004);
assign w7251 = v3451;
assign w7252 = ~w7006 & w7251;
assign v3452 = ~(w7003 | w7252);
assign w7253 = v3452;
assign w7254 = w7250 & w7253;
assign v3453 = ~(w7250 | w7253);
assign w7255 = v3453;
assign v3454 = ~(w7254 | w7255);
assign w7256 = v3454;
assign v3455 = ~(w7037 | w7244);
assign w7257 = v3455;
assign v3456 = ~(w7101 | w7241);
assign w7258 = v3456;
assign v3457 = ~(w7170 | w7238);
assign w7259 = v3457;
assign w7260 = (~w7095 & ~w7097) | (~w7095 & w17765) | (~w7097 & w17765);
assign w7261 = (~w7149 & ~w7151) | (~w7149 & w16910) | (~w7151 & w16910);
assign w7262 = (~w7067 & ~w7069) | (~w7067 & w16752) | (~w7069 & w16752);
assign w7263 = (~w7055 & ~w7057) | (~w7055 & w16753) | (~w7057 & w16753);
assign v3458 = ~(w7262 | w7263);
assign w7264 = v3458;
assign w7265 = w7262 & w7263;
assign v3459 = ~(w7264 | w7265);
assign w7266 = v3459;
assign w7267 = w7261 & ~w7266;
assign w7268 = ~w7261 & w7266;
assign v3460 = ~(w7267 | w7268);
assign w7269 = v3460;
assign w7270 = (~w7044 & ~w7046) | (~w7044 & w17140) | (~w7046 & w17140);
assign w7271 = ~w7269 & w7270;
assign w7272 = w7269 & ~w7270;
assign v3461 = ~(w7271 | w7272);
assign w7273 = v3461;
assign w7274 = (~w7200 & ~w7201) | (~w7200 & w17141) | (~w7201 & w17141);
assign w7275 = w7273 & ~w7274;
assign w7276 = ~w7273 & w7274;
assign v3462 = ~(w7275 | w7276);
assign w7277 = v3462;
assign w7278 = ~w7260 & w7277;
assign w7279 = w7260 & ~w7277;
assign v3463 = ~(w7278 | w7279);
assign w7280 = v3463;
assign w7281 = ~w7259 & w7280;
assign w7282 = w7259 & ~w7280;
assign v3464 = ~(w7281 | w7282);
assign w7283 = v3464;
assign w7284 = ~w7258 & w7283;
assign w7285 = w7258 & ~w7283;
assign v3465 = ~(w7284 | w7285);
assign w7286 = v3465;
assign v3466 = ~(w7089 | w7092);
assign w7287 = v3466;
assign v3467 = ~(w7081 | w7086);
assign w7288 = v3467;
assign w7289 = pi00 & pi60;
assign w7290 = w7075 & w7289;
assign v3468 = ~(w7075 | w7289);
assign w7291 = v3468;
assign v3469 = ~(w7290 | w7291);
assign w7292 = v3469;
assign w7293 = pi01 & pi59;
assign w7294 = pi29 & pi31;
assign v3470 = ~(w7293 | w7294);
assign w7295 = v3470;
assign w7296 = w7293 & w7294;
assign v3471 = ~(w7295 | w7296);
assign w7297 = v3471;
assign w7298 = w7292 & w7297;
assign v3472 = ~(w7292 | w7297);
assign w7299 = v3472;
assign v3473 = ~(w7298 | w7299);
assign w7300 = v3473;
assign w7301 = pi27 & pi33;
assign w7302 = pi28 & pi32;
assign w7303 = pi23 & pi37;
assign v3474 = ~(w7302 | w7303);
assign w7304 = v3474;
assign w7305 = w7302 & w7303;
assign v3475 = ~(w7304 | w7305);
assign w7306 = v3475;
assign w7307 = w7301 & ~w7306;
assign w7308 = ~w7301 & w7306;
assign v3476 = ~(w7307 | w7308);
assign w7309 = v3476;
assign w7310 = w7300 & ~w7309;
assign w7311 = ~w7300 & w7309;
assign v3477 = ~(w7310 | w7311);
assign w7312 = v3477;
assign w7313 = w7288 & ~w7312;
assign w7314 = ~w7288 & w7312;
assign v3478 = ~(w7313 | w7314);
assign w7315 = v3478;
assign w7316 = pi14 & pi46;
assign w7317 = pi12 & pi48;
assign w7318 = pi13 & pi47;
assign v3479 = ~(w7317 | w7318);
assign w7319 = v3479;
assign w7320 = pi13 & pi48;
assign w7321 = w7116 & w7320;
assign v3480 = ~(w7319 | w7321);
assign w7322 = v3480;
assign w7323 = w7316 & ~w7322;
assign w7324 = ~w7316 & w7322;
assign v3481 = ~(w7323 | w7324);
assign w7325 = v3481;
assign w7326 = pi07 & pi53;
assign w7327 = pi08 & pi52;
assign w7328 = pi18 & pi42;
assign v3482 = ~(w7327 | w7328);
assign w7329 = v3482;
assign w7330 = w7327 & w7328;
assign v3483 = ~(w7329 | w7330);
assign w7331 = v3483;
assign w7332 = w7326 & ~w7331;
assign w7333 = ~w7326 & w7331;
assign v3484 = ~(w7332 | w7333);
assign w7334 = v3484;
assign v3485 = ~(w7325 | w7334);
assign w7335 = v3485;
assign w7336 = w7325 & w7334;
assign v3486 = ~(w7335 | w7336);
assign w7337 = v3486;
assign w7338 = pi05 & pi55;
assign w7339 = pi06 & pi54;
assign w7340 = pi19 & pi41;
assign v3487 = ~(w7339 | w7340);
assign w7341 = v3487;
assign w7342 = w7339 & w7340;
assign v3488 = ~(w7341 | w7342);
assign w7343 = v3488;
assign w7344 = w7338 & ~w7343;
assign w7345 = ~w7338 & w7343;
assign v3489 = ~(w7344 | w7345);
assign w7346 = v3489;
assign w7347 = w7337 & ~w7346;
assign w7348 = ~w7337 & w7346;
assign v3490 = ~(w7347 | w7348);
assign w7349 = v3490;
assign v3491 = ~(w7315 | w7349);
assign w7350 = v3491;
assign w7351 = w7315 & w7349;
assign v3492 = ~(w7350 | w7351);
assign w7352 = v3492;
assign w7353 = ~w7287 & w7352;
assign w7354 = w7287 & ~w7352;
assign v3493 = ~(w7353 | w7354);
assign w7355 = v3493;
assign v3494 = ~(w7026 | w7028);
assign w7356 = v3494;
assign w7357 = (~w7018 & ~w7020) | (~w7018 & w17572) | (~w7020 & w17572);
assign w7358 = pi02 & pi58;
assign w7359 = pi04 & pi56;
assign v3495 = ~(w7143 | w7359);
assign w7360 = v3495;
assign w7361 = pi04 & pi57;
assign w7362 = w7141 & w7361;
assign v3496 = ~(w7360 | w7362);
assign w7363 = v3496;
assign w7364 = w7358 & ~w7363;
assign w7365 = ~w7358 & w7363;
assign v3497 = ~(w7364 | w7365);
assign w7366 = v3497;
assign w7367 = pi20 & pi40;
assign w7368 = pi21 & pi39;
assign v3498 = ~(w7205 | w7368);
assign w7369 = v3498;
assign w7370 = pi22 & pi39;
assign w7371 = w6925 & w7370;
assign v3499 = ~(w7369 | w7371);
assign w7372 = v3499;
assign w7373 = w7367 & ~w7372;
assign w7374 = ~w7367 & w7372;
assign v3500 = ~(w7373 | w7374);
assign w7375 = v3500;
assign v3501 = ~(w7366 | w7375);
assign w7376 = v3501;
assign w7377 = w7366 & w7375;
assign v3502 = ~(w7376 | w7377);
assign w7378 = v3502;
assign w7379 = pi24 & pi36;
assign w7380 = pi26 & pi34;
assign v3503 = ~(w7214 | w7380);
assign w7381 = v3503;
assign w7382 = pi26 & pi35;
assign w7383 = w7212 & w7382;
assign v3504 = ~(w7381 | w7383);
assign w7384 = v3504;
assign w7385 = w7379 & ~w7384;
assign w7386 = ~w7379 & w7384;
assign v3505 = ~(w7385 | w7386);
assign w7387 = v3505;
assign w7388 = w7378 & ~w7387;
assign w7389 = ~w7378 & w7387;
assign v3506 = ~(w7388 | w7389);
assign w7390 = v3506;
assign w7391 = ~w7357 & w7390;
assign w7392 = w7357 & ~w7390;
assign v3507 = ~(w7391 | w7392);
assign w7393 = v3507;
assign v3508 = ~(w7114 | w7118);
assign w7394 = v3508;
assign v3509 = ~(w7117 | w7394);
assign w7395 = v3509;
assign w7396 = pi09 & pi51;
assign w7397 = pi16 & pi44;
assign v3510 = ~(w7396 | w7397);
assign w7398 = v3510;
assign w7399 = w7396 & w7397;
assign v3511 = ~(w7398 | w7399);
assign w7400 = v3511;
assign w7401 = w7129 & ~w7400;
assign w7402 = ~w7129 & w7400;
assign v3512 = ~(w7401 | w7402);
assign w7403 = v3512;
assign w7404 = w7395 & ~w7403;
assign w7405 = ~w7395 & w7403;
assign v3513 = ~(w7404 | w7405);
assign w7406 = v3513;
assign w7407 = pi10 & pi50;
assign w7408 = pi15 & pi45;
assign w7409 = pi11 & pi49;
assign v3514 = ~(w7408 | w7409);
assign w7410 = v3514;
assign w7411 = w7408 & w7409;
assign v3515 = ~(w7410 | w7411);
assign w7412 = v3515;
assign w7413 = w7407 & ~w7412;
assign w7414 = ~w7407 & w7412;
assign v3516 = ~(w7413 | w7414);
assign w7415 = v3516;
assign w7416 = w7406 & ~w7415;
assign w7417 = ~w7406 & w7415;
assign v3517 = ~(w7416 | w7417);
assign w7418 = v3517;
assign v3518 = ~(w7393 | w7418);
assign w7419 = v3518;
assign w7420 = w7393 & w7418;
assign v3519 = ~(w7419 | w7420);
assign w7421 = v3519;
assign w7422 = ~w7356 & w7421;
assign w7423 = w7356 & ~w7421;
assign v3520 = ~(w7422 | w7423);
assign w7424 = v3520;
assign v3521 = ~(w7355 | w7424);
assign w7425 = v3521;
assign w7426 = w7355 & w7424;
assign v3522 = ~(w7425 | w7426);
assign w7427 = v3522;
assign v3523 = ~(w7031 | w7034);
assign w7428 = v3523;
assign v3524 = ~(w7174 | w7178);
assign w7429 = v3524;
assign v3525 = ~(w7177 | w7429);
assign w7430 = v3525;
assign w7431 = w6958 & ~w7128;
assign v3526 = ~(w7130 | w7431);
assign w7432 = v3526;
assign w7433 = w7430 & ~w7432;
assign w7434 = ~w7430 & w7432;
assign v3527 = ~(w7433 | w7434);
assign w7435 = v3527;
assign v3528 = ~(w6682 | w7109);
assign w7436 = v3528;
assign v3529 = ~(w7108 | w7436);
assign w7437 = v3529;
assign v3530 = ~(w7435 | w7437);
assign w7438 = v3530;
assign w7439 = w7435 & w7437;
assign v3531 = ~(w7438 | w7439);
assign w7440 = v3531;
assign v3532 = ~(w7220 | w7232);
assign w7441 = v3532;
assign w7442 = ~w7440 & w7441;
assign w7443 = w7440 & ~w7441;
assign v3533 = ~(w7442 | w7443);
assign w7444 = v3533;
assign v3534 = ~(w7123 | w7135);
assign w7445 = v3534;
assign w7446 = ~w7444 & w7445;
assign w7447 = w7444 & ~w7445;
assign v3535 = ~(w7446 | w7447);
assign w7448 = v3535;
assign v3536 = ~(w7164 | w7167);
assign w7449 = v3536;
assign v3537 = ~(w7192 | w7196);
assign w7450 = v3537;
assign v3538 = ~(w7152 | w7156);
assign w7451 = v3538;
assign v3539 = ~(w7155 | w7451);
assign w7452 = v3539;
assign w7453 = w7202 & ~w7204;
assign v3540 = ~(w7206 | w7453);
assign w7454 = v3540;
assign w7455 = w7452 & ~w7454;
assign w7456 = ~w7452 & w7454;
assign v3541 = ~(w7455 | w7456);
assign w7457 = v3541;
assign w7458 = w7211 & ~w7213;
assign v3542 = ~(w7215 | w7458);
assign w7459 = v3542;
assign w7460 = ~w7457 & w7459;
assign w7461 = w7457 & ~w7459;
assign v3543 = ~(w7460 | w7461);
assign w7462 = v3543;
assign v3544 = ~(w7223 | w7227);
assign w7463 = v3544;
assign v3545 = ~(w7226 | w7463);
assign w7464 = v3545;
assign w7465 = w6811 & ~w7142;
assign v3546 = ~(w7144 | w7465);
assign w7466 = v3546;
assign w7467 = w7464 & ~w7466;
assign w7468 = ~w7464 & w7466;
assign v3547 = ~(w7467 | w7468);
assign w7469 = v3547;
assign v3548 = ~(w7183 | w7187);
assign w7470 = v3548;
assign v3549 = ~(w7186 | w7470);
assign w7471 = v3549;
assign v3550 = ~(w7469 | w7471);
assign w7472 = v3550;
assign w7473 = w7469 & w7471;
assign v3551 = ~(w7472 | w7473);
assign w7474 = v3551;
assign w7475 = w7462 & w7474;
assign v3552 = ~(w7462 | w7474);
assign w7476 = v3552;
assign v3553 = ~(w7475 | w7476);
assign w7477 = v3553;
assign w7478 = ~w7450 & w7477;
assign w7479 = w7450 & ~w7477;
assign v3554 = ~(w7478 | w7479);
assign w7480 = v3554;
assign w7481 = ~w7449 & w7480;
assign w7482 = w7449 & ~w7480;
assign v3555 = ~(w7481 | w7482);
assign w7483 = v3555;
assign w7484 = w7448 & w7483;
assign v3556 = ~(w7448 | w7483);
assign w7485 = v3556;
assign v3557 = ~(w7484 | w7485);
assign w7486 = v3557;
assign w7487 = ~w7428 & w7486;
assign w7488 = w7428 & ~w7486;
assign v3558 = ~(w7487 | w7488);
assign w7489 = v3558;
assign w7490 = w7427 & w7489;
assign v3559 = ~(w7427 | w7489);
assign w7491 = v3559;
assign v3560 = ~(w7490 | w7491);
assign w7492 = v3560;
assign w7493 = w7286 & w7492;
assign v3561 = ~(w7286 | w7492);
assign w7494 = v3561;
assign v3562 = ~(w7493 | w7494);
assign w7495 = v3562;
assign w7496 = w7257 & ~w7495;
assign w7497 = ~w7257 & w7495;
assign v3563 = ~(w7496 | w7497);
assign w7498 = v3563;
assign v3564 = ~(w7003 | w7249);
assign w7499 = v3564;
assign w7500 = (~w7006 & w16544) | (~w7006 & w16545) | (w16544 & w16545);
assign w7501 = w7498 & w7500;
assign v3565 = ~(w7498 | w7500);
assign w7502 = v3565;
assign v3566 = ~(w7501 | w7502);
assign w7503 = v3566;
assign v3567 = ~(w7284 | w7493);
assign w7504 = v3567;
assign w7505 = (~w7481 & ~w7483) | (~w7481 & w17766) | (~w7483 & w17766);
assign v3568 = ~(w7272 | w7275);
assign w7506 = v3568;
assign w7507 = (~w7264 & ~w7266) | (~w7264 & w16911) | (~w7266 & w16911);
assign w7508 = pi11 & pi50;
assign w7509 = pi14 & pi47;
assign w7510 = pi12 & pi49;
assign v3569 = ~(w7509 | w7510);
assign w7511 = v3569;
assign w7512 = w7509 & w7510;
assign v3570 = ~(w7511 | w7512);
assign w7513 = v3570;
assign w7514 = w7508 & ~w7513;
assign w7515 = ~w7508 & w7513;
assign v3571 = ~(w7514 | w7515);
assign w7516 = v3571;
assign w7517 = pi16 & pi45;
assign w7518 = pi15 & pi46;
assign w7519 = pi10 & pi51;
assign v3572 = ~(w7518 | w7519);
assign w7520 = v3572;
assign w7521 = w7518 & w7519;
assign v3573 = ~(w7520 | w7521);
assign w7522 = v3573;
assign w7523 = w7517 & ~w7522;
assign w7524 = ~w7517 & w7522;
assign v3574 = ~(w7523 | w7524);
assign w7525 = v3574;
assign v3575 = ~(w7516 | w7525);
assign w7526 = v3575;
assign w7527 = w7516 & w7525;
assign v3576 = ~(w7526 | w7527);
assign w7528 = v3576;
assign w7529 = pi30 & pi31;
assign w7530 = pi29 & pi32;
assign v3577 = ~(w7529 | w7530);
assign w7531 = v3577;
assign w7532 = w7529 & w7530;
assign v3578 = ~(w7531 | w7532);
assign w7533 = v3578;
assign w7534 = w7320 & ~w7533;
assign w7535 = ~w7320 & w7533;
assign v3579 = ~(w7534 | w7535);
assign w7536 = v3579;
assign w7537 = w7528 & ~w7536;
assign w7538 = ~w7528 & w7536;
assign v3580 = ~(w7537 | w7538);
assign w7539 = v3580;
assign w7540 = ~w7507 & w7539;
assign w7541 = w7507 & ~w7539;
assign v3581 = ~(w7540 | w7541);
assign w7542 = v3581;
assign w7543 = pi06 & pi55;
assign w7544 = pi20 & pi41;
assign w7545 = pi21 & pi40;
assign v3582 = ~(w7544 | w7545);
assign w7546 = v3582;
assign w7547 = pi21 & pi41;
assign w7548 = w7367 & w7547;
assign v3583 = ~(w7546 | w7548);
assign w7549 = v3583;
assign w7550 = w7543 & ~w7549;
assign w7551 = ~w7543 & w7549;
assign v3584 = ~(w7550 | w7551);
assign w7552 = v3584;
assign w7553 = pi00 & pi61;
assign w7554 = pi02 & pi59;
assign w7555 = pi05 & pi56;
assign v3585 = ~(w7554 | w7555);
assign w7556 = v3585;
assign w7557 = w7554 & w7555;
assign v3586 = ~(w7556 | w7557);
assign w7558 = v3586;
assign w7559 = w7553 & ~w7558;
assign w7560 = ~w7553 & w7558;
assign v3587 = ~(w7559 | w7560);
assign w7561 = v3587;
assign v3588 = ~(w7552 | w7561);
assign w7562 = v3588;
assign w7563 = w7552 & w7561;
assign v3589 = ~(w7562 | w7563);
assign w7564 = v3589;
assign w7565 = pi24 & pi37;
assign w7566 = pi25 & pi36;
assign v3590 = ~(w7565 | w7566);
assign w7567 = v3590;
assign w7568 = w7565 & w7566;
assign v3591 = ~(w7567 | w7568);
assign w7569 = v3591;
assign w7570 = w7370 & ~w7569;
assign w7571 = ~w7370 & w7569;
assign v3592 = ~(w7570 | w7571);
assign w7572 = v3592;
assign w7573 = w7564 & ~w7572;
assign w7574 = ~w7564 & w7572;
assign v3593 = ~(w7573 | w7574);
assign w7575 = v3593;
assign v3594 = ~(w7542 | w7575);
assign w7576 = v3594;
assign w7577 = w7542 & w7575;
assign v3595 = ~(w7576 | w7577);
assign w7578 = v3595;
assign w7579 = ~w7506 & w7578;
assign w7580 = w7506 & ~w7578;
assign v3596 = ~(w7579 | w7580);
assign w7581 = v3596;
assign w7582 = ~w7505 & w7581;
assign w7583 = w7505 & ~w7581;
assign v3597 = ~(w7582 | w7583);
assign w7584 = v3597;
assign v3598 = ~(w7278 | w7281);
assign w7585 = v3598;
assign v3599 = ~(w7351 | w7353);
assign w7586 = v3599;
assign w7587 = (~w7290 & ~w7292) | (~w7290 & w17142) | (~w7292 & w17142);
assign v3600 = ~(w7326 | w7330);
assign w7588 = v3600;
assign v3601 = ~(w7329 | w7588);
assign w7589 = v3601;
assign v3602 = ~(w7129 | w7399);
assign w7590 = v3602;
assign v3603 = ~(w7398 | w7590);
assign w7591 = v3603;
assign w7592 = w7589 & w7591;
assign v3604 = ~(w7589 | w7591);
assign w7593 = v3604;
assign v3605 = ~(w7592 | w7593);
assign w7594 = v3605;
assign w7595 = w7587 & ~w7594;
assign w7596 = ~w7587 & w7594;
assign v3606 = ~(w7595 | w7596);
assign w7597 = v3606;
assign v3607 = ~(w7335 | w7347);
assign w7598 = v3607;
assign w7599 = ~w7597 & w7598;
assign w7600 = w7597 & ~w7598;
assign v3608 = ~(w7599 | w7600);
assign w7601 = v3608;
assign v3609 = ~(w7310 | w7314);
assign w7602 = v3609;
assign w7603 = ~w7601 & w7602;
assign w7604 = w7601 & ~w7602;
assign v3610 = ~(w7603 | w7604);
assign w7605 = v3610;
assign v3611 = ~(w7376 | w7388);
assign w7606 = v3611;
assign v3612 = ~(w7301 | w7305);
assign w7607 = v3612;
assign v3613 = ~(w7304 | w7607);
assign w7608 = v3613;
assign w7609 = w7379 & ~w7381;
assign v3614 = ~(w7383 | w7609);
assign w7610 = v3614;
assign w7611 = w7608 & ~w7610;
assign w7612 = ~w7608 & w7610;
assign v3615 = ~(w7611 | w7612);
assign w7613 = v3615;
assign w7614 = w7367 & ~w7369;
assign v3616 = ~(w7371 | w7614);
assign w7615 = v3616;
assign w7616 = ~w7613 & w7615;
assign w7617 = w7613 & ~w7615;
assign v3617 = ~(w7616 | w7617);
assign w7618 = v3617;
assign v3618 = ~(w7338 | w7342);
assign w7619 = v3618;
assign v3619 = ~(w7341 | w7619);
assign w7620 = v3619;
assign w7621 = w7358 & ~w7360;
assign v3620 = ~(w7362 | w7621);
assign w7622 = v3620;
assign w7623 = w7620 & ~w7622;
assign w7624 = ~w7620 & w7622;
assign v3621 = ~(w7623 | w7624);
assign w7625 = v3621;
assign v3622 = ~(w7407 | w7411);
assign w7626 = v3622;
assign v3623 = ~(w7410 | w7626);
assign w7627 = v3623;
assign v3624 = ~(w7625 | w7627);
assign w7628 = v3624;
assign w7629 = w7625 & w7627;
assign v3625 = ~(w7628 | w7629);
assign w7630 = v3625;
assign w7631 = w7618 & w7630;
assign v3626 = ~(w7618 | w7630);
assign w7632 = v3626;
assign v3627 = ~(w7631 | w7632);
assign w7633 = v3627;
assign w7634 = ~w7606 & w7633;
assign w7635 = w7606 & ~w7633;
assign v3628 = ~(w7634 | w7635);
assign w7636 = v3628;
assign v3629 = ~(w7605 | w7636);
assign w7637 = v3629;
assign w7638 = w7605 & w7636;
assign v3630 = ~(w7637 | w7638);
assign w7639 = v3630;
assign w7640 = w7586 & w7639;
assign v3631 = ~(w7586 | w7639);
assign w7641 = v3631;
assign v3632 = ~(w7640 | w7641);
assign w7642 = v3632;
assign v3633 = ~(w7585 | w7642);
assign w7643 = v3633;
assign w7644 = w7585 & w7642;
assign v3634 = ~(w7643 | w7644);
assign w7645 = v3634;
assign w7646 = w7584 & w7645;
assign v3635 = ~(w7584 | w7645);
assign w7647 = v3635;
assign v3636 = ~(w7646 | w7647);
assign w7648 = v3636;
assign v3637 = ~(w7487 | w7490);
assign w7649 = v3637;
assign w7650 = (~w7422 & ~w7424) | (~w7422 & w17767) | (~w7424 & w17767);
assign w7651 = (~w7391 & ~w7393) | (~w7391 & w17768) | (~w7393 & w17768);
assign v3638 = ~(w7404 | w7416);
assign w7652 = v3638;
assign w7653 = (~w7455 & ~w7457) | (~w7455 & w17769) | (~w7457 & w17769);
assign w7654 = pi01 & pi60;
assign w7655 = ~w7296 & w17573;
assign w7656 = (w7654 & w7296) | (w7654 & w17574) | (w7296 & w17574);
assign v3639 = ~(w7655 | w7656);
assign w7657 = v3639;
assign w7658 = w7316 & ~w7319;
assign v3640 = ~(w7321 | w7658);
assign w7659 = v3640;
assign v3641 = ~(w7657 | w7659);
assign w7660 = v3641;
assign w7661 = w7657 & w7659;
assign v3642 = ~(w7660 | w7661);
assign w7662 = v3642;
assign w7663 = ~w7653 & w7662;
assign w7664 = w7653 & ~w7662;
assign v3643 = ~(w7663 | w7664);
assign w7665 = v3643;
assign w7666 = ~w7652 & w7665;
assign w7667 = w7652 & ~w7665;
assign v3644 = ~(w7666 | w7667);
assign w7668 = v3644;
assign w7669 = (~w7467 & ~w7469) | (~w7467 & w17770) | (~w7469 & w17770);
assign w7670 = (~w7433 & ~w7435) | (~w7433 & w17143) | (~w7435 & w17143);
assign w7671 = pi23 & pi38;
assign w7672 = pi03 & pi58;
assign v3645 = ~(w7361 | w7672);
assign w7673 = v3645;
assign w7674 = pi04 & pi58;
assign w7675 = w7143 & w7674;
assign v3646 = ~(w7673 | w7675);
assign w7676 = v3646;
assign w7677 = w7671 & ~w7676;
assign w7678 = ~w7671 & w7676;
assign v3647 = ~(w7677 | w7678);
assign w7679 = v3647;
assign v3648 = ~(w7670 | w7679);
assign w7680 = v3648;
assign w7681 = w7670 & w7679;
assign v3649 = ~(w7680 | w7681);
assign w7682 = v3649;
assign w7683 = ~w7669 & w7682;
assign w7684 = w7669 & ~w7682;
assign v3650 = ~(w7683 | w7684);
assign w7685 = v3650;
assign w7686 = w7668 & w7685;
assign v3651 = ~(w7668 | w7685);
assign w7687 = v3651;
assign v3652 = ~(w7686 | w7687);
assign w7688 = v3652;
assign w7689 = ~w7651 & w7688;
assign w7690 = w7651 & ~w7688;
assign v3653 = ~(w7689 | w7690);
assign w7691 = v3653;
assign v3654 = ~(w7443 | w7447);
assign w7692 = v3654;
assign w7693 = (~w7475 & ~w7477) | (~w7475 & w17771) | (~w7477 & w17771);
assign w7694 = pi19 & pi42;
assign w7695 = pi07 & pi54;
assign w7696 = pi08 & pi53;
assign v3655 = ~(w7695 | w7696);
assign w7697 = v3655;
assign w7698 = pi08 & pi54;
assign w7699 = w7326 & w7698;
assign v3656 = ~(w7697 | w7699);
assign w7700 = v3656;
assign w7701 = w7694 & ~w7700;
assign w7702 = ~w7694 & w7700;
assign v3657 = ~(w7701 | w7702);
assign w7703 = v3657;
assign w7704 = pi18 & pi43;
assign w7705 = pi09 & pi52;
assign w7706 = pi17 & pi44;
assign v3658 = ~(w7705 | w7706);
assign w7707 = v3658;
assign w7708 = w7705 & w7706;
assign v3659 = ~(w7707 | w7708);
assign w7709 = v3659;
assign w7710 = w7704 & ~w7709;
assign w7711 = ~w7704 & w7709;
assign v3660 = ~(w7710 | w7711);
assign w7712 = v3660;
assign v3661 = ~(w7703 | w7712);
assign w7713 = v3661;
assign w7714 = w7703 & w7712;
assign v3662 = ~(w7713 | w7714);
assign w7715 = v3662;
assign w7716 = pi27 & pi34;
assign w7717 = pi28 & pi33;
assign v3663 = ~(w7716 | w7717);
assign w7718 = v3663;
assign w7719 = w7716 & w7717;
assign v3664 = ~(w7718 | w7719);
assign w7720 = v3664;
assign w7721 = w7382 & ~w7720;
assign w7722 = ~w7382 & w7720;
assign v3665 = ~(w7721 | w7722);
assign w7723 = v3665;
assign w7724 = w7715 & ~w7723;
assign w7725 = ~w7715 & w7723;
assign v3666 = ~(w7724 | w7725);
assign w7726 = v3666;
assign w7727 = ~w7693 & w7726;
assign w7728 = w7693 & ~w7726;
assign v3667 = ~(w7727 | w7728);
assign w7729 = v3667;
assign w7730 = ~w7692 & w7729;
assign w7731 = w7692 & ~w7729;
assign v3668 = ~(w7730 | w7731);
assign w7732 = v3668;
assign w7733 = w7691 & w7732;
assign v3669 = ~(w7691 | w7732);
assign w7734 = v3669;
assign v3670 = ~(w7733 | w7734);
assign w7735 = v3670;
assign w7736 = ~w7650 & w7735;
assign w7737 = w7650 & ~w7735;
assign v3671 = ~(w7736 | w7737);
assign w7738 = v3671;
assign w7739 = ~w7649 & w7738;
assign w7740 = w7649 & ~w7738;
assign v3672 = ~(w7739 | w7740);
assign w7741 = v3672;
assign w7742 = w7648 & w7741;
assign v3673 = ~(w7648 | w7741);
assign w7743 = v3673;
assign v3674 = ~(w7742 | w7743);
assign w7744 = v3674;
assign w7745 = ~w7504 & w7744;
assign w7746 = w7504 & ~w7744;
assign v3675 = ~(w7745 | w7746);
assign w7747 = v3675;
assign w7748 = (w7006 & w16546) | (w7006 & w16547) | (w16546 & w16547);
assign v3676 = ~(w7496 | w7748);
assign w7749 = v3676;
assign w7750 = w7747 & w7749;
assign v3677 = ~(w7747 | w7749);
assign w7751 = v3677;
assign v3678 = ~(w7750 | w7751);
assign w7752 = v3678;
assign v3679 = ~(w7496 | w7746);
assign w7753 = v3679;
assign w7754 = (~w7006 & w16548) | (~w7006 & w16549) | (w16548 & w16549);
assign v3680 = ~(w7745 | w7754);
assign w7755 = v3680;
assign v3681 = ~(w7739 | w7742);
assign w7756 = v3681;
assign v3682 = ~(w7733 | w7736);
assign w7757 = v3682;
assign w7758 = (~w7680 & ~w7682) | (~w7680 & w17575) | (~w7682 & w17575);
assign v3683 = ~(w7704 | w7708);
assign w7759 = v3683;
assign v3684 = ~(w7707 | w7759);
assign w7760 = v3684;
assign v3685 = ~(w7517 | w7521);
assign w7761 = v3685;
assign v3686 = ~(w7520 | w7761);
assign w7762 = v3686;
assign w7763 = w7760 & w7762;
assign v3687 = ~(w7760 | w7762);
assign w7764 = v3687;
assign v3688 = ~(w7763 | w7764);
assign w7765 = v3688;
assign w7766 = pi03 & pi59;
assign w7767 = pi05 & pi57;
assign v3689 = ~(w7674 | w7767);
assign w7768 = v3689;
assign w7769 = pi05 & pi58;
assign w7770 = w7361 & w7769;
assign v3690 = ~(w7768 | w7770);
assign w7771 = v3690;
assign w7772 = w7766 & ~w7771;
assign w7773 = ~w7766 & w7771;
assign v3691 = ~(w7772 | w7773);
assign w7774 = v3691;
assign w7775 = ~w7765 & w7774;
assign w7776 = w7765 & ~w7774;
assign v3692 = ~(w7775 | w7776);
assign w7777 = v3692;
assign w7778 = (~w7713 & ~w7715) | (~w7713 & w17576) | (~w7715 & w17576);
assign w7779 = w7777 & ~w7778;
assign w7780 = ~w7777 & w7778;
assign v3693 = ~(w7779 | w7780);
assign w7781 = v3693;
assign w7782 = w7758 & ~w7781;
assign w7783 = ~w7758 & w7781;
assign v3694 = ~(w7782 | w7783);
assign w7784 = v3694;
assign w7785 = (~w7611 & ~w7613) | (~w7611 & w17772) | (~w7613 & w17772);
assign w7786 = (~w7592 & ~w7594) | (~w7592 & w17144) | (~w7594 & w17144);
assign w7787 = ~pi60 & w7296;
assign v3695 = ~(w7660 | w7787);
assign w7788 = v3695;
assign v3696 = ~(w7786 | w7788);
assign w7789 = v3696;
assign w7790 = w7786 & w7788;
assign v3697 = ~(w7789 | w7790);
assign w7791 = v3697;
assign w7792 = w7785 & ~w7791;
assign w7793 = ~w7785 & w7791;
assign v3698 = ~(w7792 | w7793);
assign w7794 = v3698;
assign w7795 = (w7542 & w17577) | (w7542 & w17578) | (w17577 & w17578);
assign w7796 = (~w7542 & w17579) | (~w7542 & w17580) | (w17579 & w17580);
assign v3699 = ~(w7795 | w7796);
assign w7797 = v3699;
assign w7798 = w7784 & w7797;
assign v3700 = ~(w7784 | w7797);
assign w7799 = v3700;
assign v3701 = ~(w7798 | w7799);
assign w7800 = v3701;
assign w7801 = ~w7757 & w7800;
assign w7802 = w7757 & ~w7800;
assign v3702 = ~(w7801 | w7802);
assign w7803 = v3702;
assign v3703 = ~(w7686 | w7689);
assign w7804 = v3703;
assign w7805 = pi19 & pi43;
assign w7806 = pi18 & pi44;
assign v3704 = ~(w7698 | w7806);
assign w7807 = v3704;
assign w7808 = w7698 & w7806;
assign v3705 = ~(w7807 | w7808);
assign w7809 = v3705;
assign w7810 = w7805 & ~w7809;
assign w7811 = ~w7805 & w7809;
assign v3706 = ~(w7810 | w7811);
assign w7812 = v3706;
assign w7813 = pi27 & pi35;
assign w7814 = pi28 & pi34;
assign w7815 = pi29 & pi33;
assign v3707 = ~(w7814 | w7815);
assign w7816 = v3707;
assign w7817 = w7814 & w7815;
assign v3708 = ~(w7816 | w7817);
assign w7818 = v3708;
assign w7819 = w7813 & ~w7818;
assign w7820 = ~w7813 & w7818;
assign v3709 = ~(w7819 | w7820);
assign w7821 = v3709;
assign v3710 = ~(w7812 | w7821);
assign w7822 = v3710;
assign w7823 = w7812 & w7821;
assign v3711 = ~(w7822 | w7823);
assign w7824 = v3711;
assign w7825 = pi22 & pi40;
assign w7826 = pi23 & pi39;
assign w7827 = pi24 & pi38;
assign v3712 = ~(w7826 | w7827);
assign w7828 = v3712;
assign w7829 = pi24 & pi39;
assign w7830 = w7671 & w7829;
assign v3713 = ~(w7828 | w7830);
assign w7831 = v3713;
assign w7832 = w7825 & ~w7831;
assign w7833 = ~w7825 & w7831;
assign v3714 = ~(w7832 | w7833);
assign w7834 = v3714;
assign w7835 = w7824 & ~w7834;
assign w7836 = ~w7824 & w7834;
assign v3715 = ~(w7835 | w7836);
assign w7837 = v3715;
assign w7838 = pi31 & w7654;
assign w7839 = pi00 & pi62;
assign w7840 = pi02 & pi60;
assign v3716 = ~(w7839 | w7840);
assign w7841 = v3716;
assign w7842 = pi02 & pi62;
assign w7843 = w7289 & w7842;
assign v3717 = ~(w7841 | w7843);
assign w7844 = v3717;
assign w7845 = w7838 & ~w7844;
assign w7846 = ~w7838 & w7844;
assign v3718 = ~(w7845 | w7846);
assign w7847 = v3718;
assign w7848 = pi25 & pi37;
assign w7849 = pi26 & pi36;
assign v3719 = ~(w7848 | w7849);
assign w7850 = v3719;
assign w7851 = w7848 & w7849;
assign v3720 = ~(w7850 | w7851);
assign w7852 = v3720;
assign w7853 = w7547 & ~w7852;
assign w7854 = ~w7547 & w7852;
assign v3721 = ~(w7853 | w7854);
assign w7855 = v3721;
assign v3722 = ~(w7847 | w7855);
assign w7856 = v3722;
assign w7857 = w7847 & w7855;
assign v3723 = ~(w7856 | w7857);
assign w7858 = v3723;
assign w7859 = pi09 & pi53;
assign w7860 = pi17 & pi45;
assign w7861 = pi10 & pi52;
assign v3724 = ~(w7860 | w7861);
assign w7862 = v3724;
assign w7863 = w7860 & w7861;
assign v3725 = ~(w7862 | w7863);
assign w7864 = v3725;
assign w7865 = w7859 & ~w7864;
assign w7866 = ~w7859 & w7864;
assign v3726 = ~(w7865 | w7866);
assign w7867 = v3726;
assign w7868 = w7858 & ~w7867;
assign w7869 = ~w7858 & w7867;
assign v3727 = ~(w7868 | w7869);
assign w7870 = v3727;
assign w7871 = pi12 & pi50;
assign w7872 = pi13 & pi49;
assign w7873 = pi14 & pi48;
assign v3728 = ~(w7872 | w7873);
assign w7874 = v3728;
assign w7875 = pi14 & pi49;
assign w7876 = w7320 & w7875;
assign v3729 = ~(w7874 | w7876);
assign w7877 = v3729;
assign w7878 = w7871 & ~w7877;
assign w7879 = ~w7871 & w7877;
assign v3730 = ~(w7878 | w7879);
assign w7880 = v3730;
assign w7881 = pi16 & pi46;
assign w7882 = pi15 & pi47;
assign w7883 = pi11 & pi51;
assign v3731 = ~(w7882 | w7883);
assign w7884 = v3731;
assign w7885 = w7882 & w7883;
assign v3732 = ~(w7884 | w7885);
assign w7886 = v3732;
assign w7887 = w7881 & ~w7886;
assign w7888 = ~w7881 & w7886;
assign v3733 = ~(w7887 | w7888);
assign w7889 = v3733;
assign v3734 = ~(w7880 | w7889);
assign w7890 = v3734;
assign w7891 = w7880 & w7889;
assign v3735 = ~(w7890 | w7891);
assign w7892 = v3735;
assign w7893 = pi20 & pi42;
assign w7894 = pi06 & pi56;
assign w7895 = pi07 & pi55;
assign v3736 = ~(w7894 | w7895);
assign w7896 = v3736;
assign w7897 = pi07 & pi56;
assign w7898 = w7543 & w7897;
assign v3737 = ~(w7896 | w7898);
assign w7899 = v3737;
assign w7900 = w7893 & ~w7899;
assign w7901 = ~w7893 & w7899;
assign v3738 = ~(w7900 | w7901);
assign w7902 = v3738;
assign w7903 = w7892 & ~w7902;
assign w7904 = ~w7892 & w7902;
assign v3739 = ~(w7903 | w7904);
assign w7905 = v3739;
assign w7906 = w7870 & w7905;
assign v3740 = ~(w7870 | w7905);
assign w7907 = v3740;
assign v3741 = ~(w7906 | w7907);
assign w7908 = v3741;
assign w7909 = w7837 & w7908;
assign v3742 = ~(w7837 | w7908);
assign w7910 = v3742;
assign v3743 = ~(w7909 | w7910);
assign w7911 = v3743;
assign w7912 = ~w7804 & w7911;
assign w7913 = w7804 & ~w7911;
assign v3744 = ~(w7912 | w7913);
assign w7914 = v3744;
assign v3745 = ~(w7637 | w7640);
assign w7915 = v3745;
assign w7916 = w7914 & w7915;
assign v3746 = ~(w7914 | w7915);
assign w7917 = v3746;
assign v3747 = ~(w7916 | w7917);
assign w7918 = v3747;
assign v3748 = ~(w7803 | w7918);
assign w7919 = v3748;
assign w7920 = w7803 & w7918;
assign v3749 = ~(w7919 | w7920);
assign w7921 = v3749;
assign v3750 = ~(w7643 | w7646);
assign w7922 = v3750;
assign w7923 = (~w7526 & ~w7528) | (~w7526 & w17581) | (~w7528 & w17581);
assign w7924 = (~w7623 & ~w7625) | (~w7623 & w17146) | (~w7625 & w17146);
assign w7925 = (~w7562 & ~w7564) | (~w7562 & w16912) | (~w7564 & w16912);
assign v3751 = ~(w7924 | w7925);
assign w7926 = v3751;
assign w7927 = w7924 & w7925;
assign v3752 = ~(w7926 | w7927);
assign w7928 = v3752;
assign w7929 = w7923 & ~w7928;
assign w7930 = ~w7923 & w7928;
assign v3753 = ~(w7929 | w7930);
assign w7931 = v3753;
assign v3754 = ~(w7553 | w7557);
assign w7932 = v3754;
assign v3755 = ~(w7556 | w7932);
assign w7933 = v3755;
assign w7934 = w7543 & ~w7546;
assign v3756 = ~(w7548 | w7934);
assign w7935 = v3756;
assign w7936 = w7933 & ~w7935;
assign w7937 = ~w7933 & w7935;
assign v3757 = ~(w7936 | w7937);
assign w7938 = v3757;
assign w7939 = w7694 & ~w7697;
assign v3758 = ~(w7699 | w7939);
assign w7940 = v3758;
assign w7941 = ~w7938 & w7940;
assign w7942 = w7938 & ~w7940;
assign v3759 = ~(w7941 | w7942);
assign w7943 = v3759;
assign v3760 = ~(w7382 | w7719);
assign w7944 = v3760;
assign v3761 = ~(w7718 | w7944);
assign w7945 = v3761;
assign w7946 = w7671 & ~w7673;
assign v3762 = ~(w7675 | w7946);
assign w7947 = v3762;
assign w7948 = w7945 & ~w7947;
assign w7949 = ~w7945 & w7947;
assign v3763 = ~(w7948 | w7949);
assign w7950 = v3763;
assign v3764 = ~(w7370 | w7568);
assign w7951 = v3764;
assign v3765 = ~(w7567 | w7951);
assign w7952 = v3765;
assign v3766 = ~(w7950 | w7952);
assign w7953 = v3766;
assign w7954 = w7950 & w7952;
assign v3767 = ~(w7953 | w7954);
assign w7955 = v3767;
assign w7956 = pi30 & pi32;
assign w7957 = pi01 & pi61;
assign v3768 = ~(w7956 | w7957);
assign w7958 = v3768;
assign w7959 = w7956 & w7957;
assign v3769 = ~(w7958 | w7959);
assign w7960 = v3769;
assign v3770 = ~(w7320 | w7532);
assign w7961 = v3770;
assign v3771 = ~(w7531 | w7961);
assign w7962 = v3771;
assign w7963 = w7960 & w7962;
assign v3772 = ~(w7960 | w7962);
assign w7964 = v3772;
assign v3773 = ~(w7963 | w7964);
assign w7965 = v3773;
assign v3774 = ~(w7508 | w7512);
assign w7966 = v3774;
assign v3775 = ~(w7511 | w7966);
assign w7967 = v3775;
assign w7968 = w7965 & w7967;
assign v3776 = ~(w7965 | w7967);
assign w7969 = v3776;
assign v3777 = ~(w7968 | w7969);
assign w7970 = v3777;
assign w7971 = w7955 & w7970;
assign v3778 = ~(w7955 | w7970);
assign w7972 = v3778;
assign v3779 = ~(w7971 | w7972);
assign w7973 = v3779;
assign v3780 = ~(w7943 | w7973);
assign w7974 = v3780;
assign w7975 = w7943 & w7973;
assign v3781 = ~(w7974 | w7975);
assign w7976 = v3781;
assign v3782 = ~(w7931 | w7976);
assign w7977 = v3782;
assign w7978 = w7931 & w7976;
assign v3783 = ~(w7977 | w7978);
assign w7979 = v3783;
assign v3784 = ~(w7727 | w7730);
assign w7980 = v3784;
assign w7981 = ~w7979 & w7980;
assign w7982 = w7979 & ~w7980;
assign v3785 = ~(w7981 | w7982);
assign w7983 = v3785;
assign v3786 = ~(w7600 | w7604);
assign w7984 = v3786;
assign w7985 = (~w7631 & ~w7633) | (~w7631 & w17773) | (~w7633 & w17773);
assign v3787 = ~(w7663 | w7666);
assign w7986 = v3787;
assign v3788 = ~(w7985 | w7986);
assign w7987 = v3788;
assign w7988 = w7985 & w7986;
assign v3789 = ~(w7987 | w7988);
assign w7989 = v3789;
assign w7990 = w7984 & ~w7989;
assign w7991 = ~w7984 & w7989;
assign v3790 = ~(w7990 | w7991);
assign w7992 = v3790;
assign w7993 = (~w7579 & ~w7581) | (~w7579 & w17774) | (~w7581 & w17774);
assign w7994 = ~w7992 & w7993;
assign w7995 = w7992 & ~w7993;
assign v3791 = ~(w7994 | w7995);
assign w7996 = v3791;
assign w7997 = w7983 & w7996;
assign v3792 = ~(w7983 | w7996);
assign w7998 = v3792;
assign v3793 = ~(w7997 | w7998);
assign w7999 = v3793;
assign w8000 = ~w7922 & w7999;
assign w8001 = w7922 & ~w7999;
assign v3794 = ~(w8000 | w8001);
assign w8002 = v3794;
assign w8003 = w7921 & w8002;
assign v3795 = ~(w7921 | w8002);
assign w8004 = v3795;
assign v3796 = ~(w8003 | w8004);
assign w8005 = v3796;
assign w8006 = ~w7756 & w8005;
assign w8007 = w7756 & ~w8005;
assign v3797 = ~(w8006 | w8007);
assign w8008 = v3797;
assign w8009 = w7755 & w8008;
assign v3798 = ~(w7755 | w8008);
assign w8010 = v3798;
assign v3799 = ~(w8009 | w8010);
assign w8011 = v3799;
assign v3800 = ~(w7745 | w8006);
assign w8012 = v3800;
assign w8013 = (~w7006 & w17775) | (~w7006 & w17776) | (w17775 & w17776);
assign v3801 = ~(w8000 | w8003);
assign w8014 = v3801;
assign v3802 = ~(w7995 | w7997);
assign w8015 = v3802;
assign v3803 = ~(w7987 | w7991);
assign w8016 = v3803;
assign v3804 = ~(w7813 | w7817);
assign w8017 = v3804;
assign v3805 = ~(w7816 | w8017);
assign w8018 = v3805;
assign v3806 = ~(w7859 | w7863);
assign w8019 = v3806;
assign v3807 = ~(w7862 | w8019);
assign w8020 = v3807;
assign w8021 = w8018 & w8020;
assign v3808 = ~(w8018 | w8020);
assign w8022 = v3808;
assign v3809 = ~(w8021 | w8022);
assign w8023 = v3809;
assign v3810 = ~(w7805 | w7808);
assign w8024 = v3810;
assign v3811 = ~(w7807 | w8024);
assign w8025 = v3811;
assign v3812 = ~(w8023 | w8025);
assign w8026 = v3812;
assign w8027 = w8023 & w8025;
assign v3813 = ~(w8026 | w8027);
assign w8028 = v3813;
assign w8029 = (~w7822 & ~w7824) | (~w7822 & w16754) | (~w7824 & w16754);
assign w8030 = ~w8028 & w8029;
assign w8031 = w8028 & ~w8029;
assign v3814 = ~(w8030 | w8031);
assign w8032 = v3814;
assign w8033 = (~w7890 & ~w7892) | (~w7890 & w17147) | (~w7892 & w17147);
assign w8034 = ~w8032 & w8033;
assign w8035 = w8032 & ~w8033;
assign v3815 = ~(w8034 | w8035);
assign w8036 = v3815;
assign w8037 = pi00 & pi63;
assign w8038 = w7959 & w8037;
assign v3816 = ~(w7959 | w8037);
assign w8039 = v3816;
assign v3817 = ~(w8038 | w8039);
assign w8040 = v3817;
assign w8041 = pi01 & pi62;
assign w8042 = pi32 & ~w8041;
assign w8043 = ~pi32 & w8041;
assign v3818 = ~(w8042 | w8043);
assign w8044 = v3818;
assign w8045 = w8040 & ~w8044;
assign w8046 = ~w8040 & w8044;
assign v3819 = ~(w8045 | w8046);
assign w8047 = v3819;
assign w8048 = pi26 & pi37;
assign w8049 = pi25 & pi38;
assign v3820 = ~(w8048 | w8049);
assign w8050 = v3820;
assign w8051 = pi26 & pi38;
assign w8052 = w7848 & w8051;
assign v3821 = ~(w8050 | w8052);
assign w8053 = v3821;
assign w8054 = w7829 & ~w8053;
assign w8055 = ~w7829 & w8053;
assign v3822 = ~(w8054 | w8055);
assign w8056 = v3822;
assign w8057 = pi27 & pi36;
assign w8058 = pi29 & pi34;
assign w8059 = pi28 & pi35;
assign v3823 = ~(w8058 | w8059);
assign w8060 = v3823;
assign w8061 = pi29 & pi35;
assign w8062 = w7814 & w8061;
assign v3824 = ~(w8060 | w8062);
assign w8063 = v3824;
assign w8064 = w8057 & ~w8063;
assign w8065 = ~w8057 & w8063;
assign v3825 = ~(w8064 | w8065);
assign w8066 = v3825;
assign v3826 = ~(w8056 | w8066);
assign w8067 = v3826;
assign w8068 = w8056 & w8066;
assign v3827 = ~(w8067 | w8068);
assign w8069 = v3827;
assign w8070 = w8047 & w8069;
assign v3828 = ~(w8047 | w8069);
assign w8071 = v3828;
assign v3829 = ~(w8070 | w8071);
assign w8072 = v3829;
assign w8073 = (~w7789 & ~w7791) | (~w7789 & w17582) | (~w7791 & w17582);
assign v3830 = ~(w7856 | w7868);
assign w8074 = v3830;
assign v3831 = ~(w8073 | w8074);
assign w8075 = v3831;
assign w8076 = w8073 & w8074;
assign v3832 = ~(w8075 | w8076);
assign w8077 = v3832;
assign v3833 = ~(w8072 | w8077);
assign w8078 = v3833;
assign w8079 = w8072 & w8077;
assign v3834 = ~(w8078 | w8079);
assign w8080 = v3834;
assign v3835 = ~(w8036 | w8080);
assign w8081 = v3835;
assign w8082 = w8036 & w8080;
assign v3836 = ~(w8081 | w8082);
assign w8083 = v3836;
assign w8084 = ~w8016 & w8083;
assign w8085 = w8016 & ~w8083;
assign v3837 = ~(w8084 | w8085);
assign w8086 = v3837;
assign w8087 = ~w8015 & w8086;
assign w8088 = w8015 & ~w8086;
assign v3838 = ~(w8087 | w8088);
assign w8089 = v3838;
assign v3839 = ~(w7978 | w7982);
assign w8090 = v3839;
assign w8091 = (~w7795 & ~w7797) | (~w7795 & w17777) | (~w7797 & w17777);
assign w8092 = pi31 & pi32;
assign w8093 = pi30 & pi33;
assign v3840 = ~(w8092 | w8093);
assign w8094 = v3840;
assign w8095 = w8092 & w8093;
assign v3841 = ~(w8094 | w8095);
assign w8096 = v3841;
assign w8097 = w7875 & ~w8096;
assign w8098 = ~w7875 & w8096;
assign v3842 = ~(w8097 | w8098);
assign w8099 = v3842;
assign w8100 = pi23 & pi40;
assign w8101 = pi06 & pi57;
assign w8102 = pi20 & pi43;
assign v3843 = ~(w8101 | w8102);
assign w8103 = v3843;
assign w8104 = w8101 & w8102;
assign v3844 = ~(w8103 | w8104);
assign w8105 = v3844;
assign w8106 = w8100 & ~w8105;
assign w8107 = ~w8100 & w8105;
assign v3845 = ~(w8106 | w8107);
assign w8108 = v3845;
assign v3846 = ~(w8099 | w8108);
assign w8109 = v3846;
assign w8110 = w8099 & w8108;
assign v3847 = ~(w8109 | w8110);
assign w8111 = v3847;
assign w8112 = pi08 & pi55;
assign w8113 = pi19 & pi44;
assign v3848 = ~(w8112 | w8113);
assign w8114 = v3848;
assign w8115 = w8112 & w8113;
assign v3849 = ~(w8114 | w8115);
assign w8116 = v3849;
assign w8117 = w7897 & ~w8116;
assign w8118 = ~w7897 & w8116;
assign v3850 = ~(w8117 | w8118);
assign w8119 = v3850;
assign w8120 = w8111 & ~w8119;
assign w8121 = ~w8111 & w8119;
assign v3851 = ~(w8120 | w8121);
assign w8122 = v3851;
assign v3852 = ~(w7881 | w7885);
assign w8123 = v3852;
assign v3853 = ~(w7884 | w8123);
assign w8124 = v3853;
assign w8125 = pi02 & pi61;
assign w8126 = pi03 & pi60;
assign w8127 = pi04 & pi59;
assign v3854 = ~(w8126 | w8127);
assign w8128 = v3854;
assign w8129 = pi04 & pi60;
assign w8130 = w7766 & w8129;
assign v3855 = ~(w8128 | w8130);
assign w8131 = v3855;
assign w8132 = w8125 & ~w8131;
assign w8133 = ~w8125 & w8131;
assign v3856 = ~(w8132 | w8133);
assign w8134 = v3856;
assign w8135 = w8124 & ~w8134;
assign w8136 = ~w8124 & w8134;
assign v3857 = ~(w8135 | w8136);
assign w8137 = v3857;
assign w8138 = pi22 & pi41;
assign w8139 = pi21 & pi42;
assign v3858 = ~(w8138 | w8139);
assign w8140 = v3858;
assign w8141 = pi22 & pi42;
assign w8142 = w7547 & w8141;
assign v3859 = ~(w8140 | w8142);
assign w8143 = v3859;
assign w8144 = w7769 & ~w8143;
assign w8145 = ~w7769 & w8143;
assign v3860 = ~(w8144 | w8145);
assign w8146 = v3860;
assign w8147 = w8137 & ~w8146;
assign w8148 = ~w8137 & w8146;
assign v3861 = ~(w8147 | w8148);
assign w8149 = v3861;
assign w8150 = w8122 & w8149;
assign v3862 = ~(w8122 | w8149);
assign w8151 = v3862;
assign v3863 = ~(w8150 | w8151);
assign w8152 = v3863;
assign w8153 = pi18 & pi45;
assign w8154 = pi17 & pi46;
assign w8155 = pi09 & pi54;
assign v3864 = ~(w8154 | w8155);
assign w8156 = v3864;
assign w8157 = w8154 & w8155;
assign v3865 = ~(w8156 | w8157);
assign w8158 = v3865;
assign w8159 = w8153 & ~w8158;
assign w8160 = ~w8153 & w8158;
assign v3866 = ~(w8159 | w8160);
assign w8161 = v3866;
assign w8162 = pi10 & pi53;
assign w8163 = pi16 & pi47;
assign w8164 = pi11 & pi52;
assign v3867 = ~(w8163 | w8164);
assign w8165 = v3867;
assign w8166 = w8163 & w8164;
assign v3868 = ~(w8165 | w8166);
assign w8167 = v3868;
assign w8168 = w8162 & ~w8167;
assign w8169 = ~w8162 & w8167;
assign v3869 = ~(w8168 | w8169);
assign w8170 = v3869;
assign v3870 = ~(w8161 | w8170);
assign w8171 = v3870;
assign w8172 = w8161 & w8170;
assign v3871 = ~(w8171 | w8172);
assign w8173 = v3871;
assign w8174 = pi15 & pi48;
assign w8175 = pi12 & pi51;
assign w8176 = pi13 & pi50;
assign v3872 = ~(w8175 | w8176);
assign w8177 = v3872;
assign w8178 = pi13 & pi51;
assign w8179 = w7871 & w8178;
assign v3873 = ~(w8177 | w8179);
assign w8180 = v3873;
assign w8181 = w8174 & ~w8180;
assign w8182 = ~w8174 & w8180;
assign v3874 = ~(w8181 | w8182);
assign w8183 = v3874;
assign w8184 = w8173 & ~w8183;
assign w8185 = ~w8173 & w8183;
assign v3875 = ~(w8184 | w8185);
assign w8186 = v3875;
assign w8187 = w8152 & w8186;
assign v3876 = ~(w8152 | w8186);
assign w8188 = v3876;
assign v3877 = ~(w8187 | w8188);
assign w8189 = v3877;
assign w8190 = ~w8091 & w8189;
assign w8191 = w8091 & ~w8189;
assign v3878 = ~(w8190 | w8191);
assign w8192 = v3878;
assign w8193 = ~w8090 & w8192;
assign w8194 = w8090 & ~w8192;
assign v3879 = ~(w8193 | w8194);
assign w8195 = v3879;
assign v3880 = ~(w8089 | w8195);
assign w8196 = v3880;
assign w8197 = w8089 & w8195;
assign v3881 = ~(w8196 | w8197);
assign w8198 = v3881;
assign v3882 = ~(w7801 | w7920);
assign w8199 = v3882;
assign v3883 = ~(w7912 | w7916);
assign w8200 = v3883;
assign v3884 = ~(w7779 | w7783);
assign w8201 = v3884;
assign w8202 = (~w7971 & ~w7973) | (~w7971 & w17148) | (~w7973 & w17148);
assign w8203 = (~w7926 & ~w7928) | (~w7926 & w17149) | (~w7928 & w17149);
assign v3885 = ~(w8202 | w8203);
assign w8204 = v3885;
assign w8205 = w8202 & w8203;
assign v3886 = ~(w8204 | w8205);
assign w8206 = v3886;
assign w8207 = w8201 & ~w8206;
assign w8208 = ~w8201 & w8206;
assign v3887 = ~(w8207 | w8208);
assign w8209 = v3887;
assign w8210 = (~w7963 & ~w7965) | (~w7963 & w17583) | (~w7965 & w17583);
assign w8211 = (~w7763 & ~w7765) | (~w7763 & w16913) | (~w7765 & w16913);
assign w8212 = (~w7948 & ~w7950) | (~w7948 & w16914) | (~w7950 & w16914);
assign v3888 = ~(w8211 | w8212);
assign w8213 = v3888;
assign w8214 = w8211 & w8212;
assign v3889 = ~(w8213 | w8214);
assign w8215 = v3889;
assign w8216 = w8210 & ~w8215;
assign w8217 = ~w8210 & w8215;
assign v3890 = ~(w8216 | w8217);
assign w8218 = v3890;
assign w8219 = (~w7906 & ~w7908) | (~w7906 & w17584) | (~w7908 & w17584);
assign w8220 = ~w8218 & w8219;
assign w8221 = w8218 & ~w8219;
assign v3891 = ~(w8220 | w8221);
assign w8222 = v3891;
assign w8223 = w7825 & ~w7828;
assign v3892 = ~(w7830 | w8223);
assign w8224 = v3892;
assign w8225 = w7893 & ~w7896;
assign v3893 = ~(w7898 | w8225);
assign w8226 = v3893;
assign v3894 = ~(w8224 | w8226);
assign w8227 = v3894;
assign w8228 = w8224 & w8226;
assign v3895 = ~(w8227 | w8228);
assign w8229 = v3895;
assign w8230 = w7871 & ~w7874;
assign v3896 = ~(w7876 | w8230);
assign w8231 = v3896;
assign w8232 = ~w8229 & w8231;
assign w8233 = w8229 & ~w8231;
assign v3897 = ~(w8232 | w8233);
assign w8234 = v3897;
assign v3898 = ~(w7547 | w7851);
assign w8235 = v3898;
assign v3899 = ~(w7850 | w8235);
assign w8236 = v3899;
assign w8237 = w7766 & ~w7768;
assign v3900 = ~(w7770 | w8237);
assign w8238 = v3900;
assign w8239 = w8236 & ~w8238;
assign w8240 = ~w8236 & w8238;
assign v3901 = ~(w8239 | w8240);
assign w8241 = v3901;
assign w8242 = w7838 & ~w7841;
assign v3902 = ~(w7843 | w8242);
assign w8243 = v3902;
assign w8244 = ~w8241 & w8243;
assign w8245 = w8241 & ~w8243;
assign v3903 = ~(w8244 | w8245);
assign w8246 = v3903;
assign w8247 = (~w7936 & ~w7938) | (~w7936 & w16915) | (~w7938 & w16915);
assign w8248 = ~w8246 & w8247;
assign w8249 = w8246 & ~w8247;
assign v3904 = ~(w8248 | w8249);
assign w8250 = v3904;
assign w8251 = w8234 & w8250;
assign v3905 = ~(w8234 | w8250);
assign w8252 = v3905;
assign v3906 = ~(w8251 | w8252);
assign w8253 = v3906;
assign w8254 = w8222 & w8253;
assign v3907 = ~(w8222 | w8253);
assign w8255 = v3907;
assign v3908 = ~(w8254 | w8255);
assign w8256 = v3908;
assign v3909 = ~(w8209 | w8256);
assign w8257 = v3909;
assign w8258 = w8209 & w8256;
assign v3910 = ~(w8257 | w8258);
assign w8259 = v3910;
assign w8260 = w8200 & ~w8259;
assign w8261 = ~w8200 & w8259;
assign v3911 = ~(w8260 | w8261);
assign w8262 = v3911;
assign w8263 = ~w8199 & w8262;
assign w8264 = w8199 & ~w8262;
assign v3912 = ~(w8263 | w8264);
assign w8265 = v3912;
assign v3913 = ~(w8198 | w8265);
assign w8266 = v3913;
assign w8267 = w8198 & w8265;
assign v3914 = ~(w8266 | w8267);
assign w8268 = v3914;
assign w8269 = w8014 & ~w8268;
assign w8270 = ~w8014 & w8268;
assign v3915 = ~(w8269 | w8270);
assign w8271 = v3915;
assign v3916 = ~(w8013 | w8271);
assign w8272 = v3916;
assign w8273 = w8013 & w8271;
assign v3917 = ~(w8272 | w8273);
assign w8274 = v3917;
assign w8275 = w7829 & ~w8050;
assign v3918 = ~(w8052 | w8275);
assign w8276 = v3918;
assign w8277 = w8174 & ~w8177;
assign v3919 = ~(w8179 | w8277);
assign w8278 = v3919;
assign v3920 = ~(w8276 | w8278);
assign w8279 = v3920;
assign w8280 = w8276 & w8278;
assign v3921 = ~(w8279 | w8280);
assign w8281 = v3921;
assign v3922 = ~(w8162 | w8166);
assign w8282 = v3922;
assign v3923 = ~(w8165 | w8282);
assign w8283 = v3923;
assign v3924 = ~(w8281 | w8283);
assign w8284 = v3924;
assign w8285 = w8281 & w8283;
assign v3925 = ~(w8284 | w8285);
assign w8286 = v3925;
assign w8287 = (~w8109 & ~w8111) | (~w8109 & w17585) | (~w8111 & w17585);
assign w8288 = ~w8286 & w8287;
assign w8289 = w8286 & ~w8287;
assign v3926 = ~(w8288 | w8289);
assign w8290 = v3926;
assign v3927 = ~(w8171 | w8184);
assign w8291 = v3927;
assign w8292 = ~w8290 & w8291;
assign w8293 = w8290 & ~w8291;
assign v3928 = ~(w8292 | w8293);
assign w8294 = v3928;
assign w8295 = (~w8204 & ~w8206) | (~w8204 & w17586) | (~w8206 & w17586);
assign w8296 = ~w8294 & w8295;
assign w8297 = w8294 & ~w8295;
assign v3929 = ~(w8296 | w8297);
assign w8298 = v3929;
assign v3930 = ~(w7875 | w8095);
assign w8299 = v3930;
assign v3931 = ~(w8094 | w8299);
assign w8300 = v3931;
assign w8301 = pi32 & pi62;
assign w8302 = pi32 & pi63;
assign w8303 = w8041 & w8302;
assign w8304 = (pi01 & w8301) | (pi01 & w16755) | (w8301 & w16755);
assign w8305 = ~w8303 & w8304;
assign w8306 = w8300 & w8305;
assign v3932 = ~(w8300 | w8305);
assign w8307 = v3932;
assign v3933 = ~(w8306 | w8307);
assign w8308 = v3933;
assign w8309 = pi11 & pi53;
assign w8310 = pi12 & pi52;
assign v3934 = ~(w8309 | w8310);
assign w8311 = v3934;
assign w8312 = pi12 & pi53;
assign w8313 = w8164 & w8312;
assign v3935 = ~(w8311 | w8313);
assign w8314 = v3935;
assign w8315 = w8178 & ~w8314;
assign w8316 = ~w8178 & w8314;
assign v3936 = ~(w8315 | w8316);
assign w8317 = v3936;
assign w8318 = pi09 & pi55;
assign w8319 = pi15 & pi49;
assign w8320 = pi10 & pi54;
assign v3937 = ~(w8319 | w8320);
assign w8321 = v3937;
assign w8322 = w8319 & w8320;
assign v3938 = ~(w8321 | w8322);
assign w8323 = v3938;
assign w8324 = w8318 & ~w8323;
assign w8325 = ~w8318 & w8323;
assign v3939 = ~(w8324 | w8325);
assign w8326 = v3939;
assign v3940 = ~(w8317 | w8326);
assign w8327 = v3940;
assign w8328 = w8317 & w8326;
assign v3941 = ~(w8327 | w8328);
assign w8329 = v3941;
assign w8330 = w8308 & w8329;
assign v3942 = ~(w8308 | w8329);
assign w8331 = v3942;
assign v3943 = ~(w8330 | w8331);
assign w8332 = v3943;
assign w8333 = (~w8213 & ~w8215) | (~w8213 & w17150) | (~w8215 & w17150);
assign v3944 = ~(w8135 | w8147);
assign w8334 = v3944;
assign v3945 = ~(w8333 | w8334);
assign w8335 = v3945;
assign w8336 = w8333 & w8334;
assign v3946 = ~(w8335 | w8336);
assign w8337 = v3946;
assign v3947 = ~(w8332 | w8337);
assign w8338 = v3947;
assign w8339 = w8332 & w8337;
assign v3948 = ~(w8338 | w8339);
assign w8340 = v3948;
assign v3949 = ~(w8298 | w8340);
assign w8341 = v3949;
assign w8342 = w8298 & w8340;
assign v3950 = ~(w8341 | w8342);
assign w8343 = v3950;
assign v3951 = ~(w8258 | w8261);
assign w8344 = v3951;
assign w8345 = w8343 & ~w8344;
assign w8346 = ~w8343 & w8344;
assign v3952 = ~(w8345 | w8346);
assign w8347 = v3952;
assign w8348 = (~w8221 & ~w8222) | (~w8221 & w17778) | (~w8222 & w17778);
assign w8349 = pi16 & pi48;
assign w8350 = pi08 & pi56;
assign v3953 = ~(w8349 | w8350);
assign w8351 = v3953;
assign w8352 = w8349 & w8350;
assign v3954 = ~(w8351 | w8352);
assign w8353 = v3954;
assign w8354 = w8051 & ~w8353;
assign w8355 = ~w8051 & w8353;
assign v3955 = ~(w8354 | w8355);
assign w8356 = v3955;
assign w8357 = pi27 & pi37;
assign w8358 = pi28 & pi36;
assign v3956 = ~(w8061 | w8358);
assign w8359 = v3956;
assign w8360 = w8061 & w8358;
assign v3957 = ~(w8359 | w8360);
assign w8361 = v3957;
assign w8362 = w8357 & ~w8361;
assign w8363 = ~w8357 & w8361;
assign v3958 = ~(w8362 | w8363);
assign w8364 = v3958;
assign v3959 = ~(w8356 | w8364);
assign w8365 = v3959;
assign w8366 = w8356 & w8364;
assign v3960 = ~(w8365 | w8366);
assign w8367 = v3960;
assign w8368 = pi14 & pi50;
assign w8369 = pi31 & pi33;
assign w8370 = pi30 & pi34;
assign v3961 = ~(w8369 | w8370);
assign w8371 = v3961;
assign w8372 = w8369 & w8370;
assign v3962 = ~(w8371 | w8372);
assign w8373 = v3962;
assign w8374 = w8368 & ~w8373;
assign w8375 = ~w8368 & w8373;
assign v3963 = ~(w8374 | w8375);
assign w8376 = v3963;
assign w8377 = w8367 & ~w8376;
assign w8378 = ~w8367 & w8376;
assign v3964 = ~(w8377 | w8378);
assign w8379 = v3964;
assign w8380 = (~w8038 & ~w8040) | (~w8038 & w17151) | (~w8040 & w17151);
assign w8381 = pi05 & pi59;
assign w8382 = pi18 & pi46;
assign w8383 = pi19 & pi45;
assign v3965 = ~(w8382 | w8383);
assign w8384 = v3965;
assign w8385 = pi19 & pi46;
assign w8386 = w8153 & w8385;
assign v3966 = ~(w8384 | w8386);
assign w8387 = v3966;
assign w8388 = w8381 & ~w8387;
assign w8389 = ~w8381 & w8387;
assign v3967 = ~(w8388 | w8389);
assign w8390 = v3967;
assign v3968 = ~(w8380 | w8390);
assign w8391 = v3968;
assign w8392 = w8380 & w8390;
assign v3969 = ~(w8391 | w8392);
assign w8393 = v3969;
assign w8394 = pi03 & pi61;
assign v3970 = ~(w8129 | w8394);
assign w8395 = v3970;
assign w8396 = pi04 & pi61;
assign w8397 = w8126 & w8396;
assign v3971 = ~(w8395 | w8397);
assign w8398 = v3971;
assign w8399 = w7842 & ~w8398;
assign w8400 = ~w7842 & w8398;
assign v3972 = ~(w8399 | w8400);
assign w8401 = v3972;
assign w8402 = w8393 & ~w8401;
assign w8403 = ~w8393 & w8401;
assign v3973 = ~(w8402 | w8403);
assign w8404 = v3973;
assign w8405 = w8379 & w8404;
assign v3974 = ~(w8379 | w8404);
assign w8406 = v3974;
assign v3975 = ~(w8405 | w8406);
assign w8407 = v3975;
assign w8408 = pi20 & pi44;
assign w8409 = pi21 & pi43;
assign v3976 = ~(w8141 | w8409);
assign w8410 = v3976;
assign w8411 = pi22 & pi43;
assign w8412 = w8139 & w8411;
assign v3977 = ~(w8410 | w8412);
assign w8413 = v3977;
assign w8414 = w8408 & ~w8413;
assign w8415 = ~w8408 & w8413;
assign v3978 = ~(w8414 | w8415);
assign w8416 = v3978;
assign w8417 = pi06 & pi58;
assign w8418 = pi17 & pi47;
assign w8419 = pi07 & pi57;
assign v3979 = ~(w8418 | w8419);
assign w8420 = v3979;
assign w8421 = w8418 & w8419;
assign v3980 = ~(w8420 | w8421);
assign w8422 = v3980;
assign w8423 = w8417 & ~w8422;
assign w8424 = ~w8417 & w8422;
assign v3981 = ~(w8423 | w8424);
assign w8425 = v3981;
assign v3982 = ~(w8416 | w8425);
assign w8426 = v3982;
assign w8427 = w8416 & w8425;
assign v3983 = ~(w8426 | w8427);
assign w8428 = v3983;
assign w8429 = pi23 & pi41;
assign w8430 = pi24 & pi40;
assign w8431 = pi25 & pi39;
assign v3984 = ~(w8430 | w8431);
assign w8432 = v3984;
assign w8433 = w8430 & w8431;
assign v3985 = ~(w8432 | w8433);
assign w8434 = v3985;
assign w8435 = w8429 & ~w8434;
assign w8436 = ~w8429 & w8434;
assign v3986 = ~(w8435 | w8436);
assign w8437 = v3986;
assign w8438 = w8428 & ~w8437;
assign w8439 = ~w8428 & w8437;
assign v3987 = ~(w8438 | w8439);
assign w8440 = v3987;
assign w8441 = w8407 & w8440;
assign v3988 = ~(w8407 | w8440);
assign w8442 = v3988;
assign v3989 = ~(w8441 | w8442);
assign w8443 = v3989;
assign w8444 = ~w8348 & w8443;
assign w8445 = w8348 & ~w8443;
assign v3990 = ~(w8444 | w8445);
assign w8446 = v3990;
assign w8447 = (~w8239 & ~w8241) | (~w8239 & w17152) | (~w8241 & w17152);
assign w8448 = (~w8227 & ~w8229) | (~w8227 & w16756) | (~w8229 & w16756);
assign w8449 = (~w8021 & ~w8023) | (~w8021 & w16757) | (~w8023 & w16757);
assign v3991 = ~(w8448 | w8449);
assign w8450 = v3991;
assign w8451 = w8448 & w8449;
assign v3992 = ~(w8450 | w8451);
assign w8452 = v3992;
assign w8453 = w8447 & ~w8452;
assign w8454 = ~w8447 & w8452;
assign v3993 = ~(w8453 | w8454);
assign w8455 = v3993;
assign w8456 = (~w8031 & ~w8032) | (~w8031 & w16916) | (~w8032 & w16916);
assign w8457 = (~w8249 & ~w8250) | (~w8249 & w16917) | (~w8250 & w16917);
assign v3994 = ~(w8456 | w8457);
assign w8458 = v3994;
assign w8459 = w8456 & w8457;
assign v3995 = ~(w8458 | w8459);
assign w8460 = v3995;
assign w8461 = w8455 & w8460;
assign v3996 = ~(w8455 | w8460);
assign w8462 = v3996;
assign v3997 = ~(w8461 | w8462);
assign w8463 = v3997;
assign w8464 = w8446 & w8463;
assign v3998 = ~(w8446 | w8463);
assign w8465 = v3998;
assign v3999 = ~(w8464 | w8465);
assign w8466 = v3999;
assign w8467 = w8347 & w8466;
assign v4000 = ~(w8347 | w8466);
assign w8468 = v4000;
assign v4001 = ~(w8467 | w8468);
assign w8469 = v4001;
assign v4002 = ~(w8087 | w8197);
assign w8470 = v4002;
assign v4003 = ~(w8190 | w8193);
assign w8471 = v4003;
assign w8472 = (~w8082 & ~w8083) | (~w8082 & w17779) | (~w8083 & w17779);
assign v4004 = ~(w8067 | w8070);
assign w8473 = v4004;
assign v4005 = ~(w8153 | w8157);
assign w8474 = v4005;
assign v4006 = ~(w8156 | w8474);
assign w8475 = v4006;
assign v4007 = ~(w8100 | w8104);
assign w8476 = v4007;
assign v4008 = ~(w8103 | w8476);
assign w8477 = v4008;
assign w8478 = w8475 & w8477;
assign v4009 = ~(w8475 | w8477);
assign w8479 = v4009;
assign v4010 = ~(w8478 | w8479);
assign w8480 = v4010;
assign w8481 = w8057 & ~w8060;
assign v4011 = ~(w8062 | w8481);
assign w8482 = v4011;
assign w8483 = ~w8480 & w8482;
assign w8484 = w8480 & ~w8482;
assign v4012 = ~(w8483 | w8484);
assign w8485 = v4012;
assign w8486 = w8125 & ~w8128;
assign v4013 = ~(w8130 | w8486);
assign w8487 = v4013;
assign w8488 = w7769 & ~w8140;
assign v4014 = ~(w8142 | w8488);
assign w8489 = v4014;
assign v4015 = ~(w8487 | w8489);
assign w8490 = v4015;
assign w8491 = w8487 & w8489;
assign v4016 = ~(w8490 | w8491);
assign w8492 = v4016;
assign v4017 = ~(w7897 | w8115);
assign w8493 = v4017;
assign v4018 = ~(w8114 | w8493);
assign w8494 = v4018;
assign v4019 = ~(w8492 | w8494);
assign w8495 = v4019;
assign w8496 = w8492 & w8494;
assign v4020 = ~(w8495 | w8496);
assign w8497 = v4020;
assign w8498 = w8485 & w8497;
assign v4021 = ~(w8485 | w8497);
assign w8499 = v4021;
assign v4022 = ~(w8498 | w8499);
assign w8500 = v4022;
assign w8501 = ~w8473 & w8500;
assign w8502 = w8473 & ~w8500;
assign v4023 = ~(w8501 | w8502);
assign w8503 = v4023;
assign v4024 = ~(w8150 | w8187);
assign w8504 = v4024;
assign w8505 = (~w8075 & ~w8077) | (~w8075 & w17780) | (~w8077 & w17780);
assign v4025 = ~(w8504 | w8505);
assign w8506 = v4025;
assign w8507 = w8504 & w8505;
assign v4026 = ~(w8506 | w8507);
assign w8508 = v4026;
assign v4027 = ~(w8503 | w8508);
assign w8509 = v4027;
assign w8510 = w8503 & w8508;
assign v4028 = ~(w8509 | w8510);
assign w8511 = v4028;
assign w8512 = ~w8472 & w8511;
assign w8513 = w8472 & ~w8511;
assign v4029 = ~(w8512 | w8513);
assign w8514 = v4029;
assign w8515 = ~w8471 & w8514;
assign w8516 = w8471 & ~w8514;
assign v4030 = ~(w8515 | w8516);
assign w8517 = v4030;
assign w8518 = ~w8470 & w8517;
assign w8519 = w8470 & ~w8517;
assign v4031 = ~(w8518 | w8519);
assign w8520 = v4031;
assign w8521 = w8469 & w8520;
assign v4032 = ~(w8469 | w8520);
assign w8522 = v4032;
assign v4033 = ~(w8521 | w8522);
assign w8523 = v4033;
assign v4034 = ~(w8263 | w8267);
assign w8524 = v4034;
assign w8525 = w8523 & ~w8524;
assign w8526 = ~w8523 & w8524;
assign v4035 = ~(w8269 | w8526);
assign w8527 = v4035;
assign w8528 = (~w7006 & w17781) | (~w7006 & w17782) | (w17781 & w17782);
assign w8529 = ~w8525 & w8528;
assign v4036 = ~(w8525 | w8526);
assign w8530 = v4036;
assign w8531 = w8013 & ~w8269;
assign v4037 = ~(w8270 | w8530);
assign w8532 = v4037;
assign w8533 = ~w8531 & w8532;
assign v4038 = ~(w8529 | w8533);
assign w8534 = v4038;
assign v4039 = ~(w8525 | w8528);
assign w8535 = v4039;
assign v4040 = ~(w8518 | w8521);
assign w8536 = v4040;
assign v4041 = ~(w8345 | w8467);
assign w8537 = v4041;
assign v4042 = ~(w8444 | w8464);
assign w8538 = v4042;
assign w8539 = (~w8297 & ~w8298) | (~w8297 & w17783) | (~w8298 & w17783);
assign w8540 = (~w8327 & ~w8329) | (~w8327 & w17587) | (~w8329 & w17587);
assign v4043 = ~(w8429 | w8433);
assign w8541 = v4043;
assign v4044 = ~(w8432 | w8541);
assign w8542 = v4044;
assign v4045 = ~(w8318 | w8322);
assign w8543 = v4045;
assign v4046 = ~(w8321 | w8543);
assign w8544 = v4046;
assign w8545 = w8542 & w8544;
assign v4047 = ~(w8542 | w8544);
assign w8546 = v4047;
assign v4048 = ~(w8545 | w8546);
assign w8547 = v4048;
assign v4049 = ~(w8417 | w8421);
assign w8548 = v4049;
assign v4050 = ~(w8420 | w8548);
assign w8549 = v4050;
assign v4051 = ~(w8547 | w8549);
assign w8550 = v4051;
assign w8551 = w8547 & w8549;
assign v4052 = ~(w8550 | w8551);
assign w8552 = v4052;
assign w8553 = w7842 & ~w8395;
assign v4053 = ~(w8397 | w8553);
assign w8554 = v4053;
assign w8555 = w8381 & ~w8384;
assign v4054 = ~(w8386 | w8555);
assign w8556 = v4054;
assign v4055 = ~(w8554 | w8556);
assign w8557 = v4055;
assign w8558 = w8554 & w8556;
assign v4056 = ~(w8557 | w8558);
assign w8559 = v4056;
assign v4057 = ~(w8051 | w8352);
assign w8560 = v4057;
assign v4058 = ~(w8351 | w8560);
assign w8561 = v4058;
assign v4059 = ~(w8559 | w8561);
assign w8562 = v4059;
assign w8563 = w8559 & w8561;
assign v4060 = ~(w8562 | w8563);
assign w8564 = v4060;
assign w8565 = w8552 & w8564;
assign v4061 = ~(w8552 | w8564);
assign w8566 = v4061;
assign v4062 = ~(w8565 | w8566);
assign w8567 = v4062;
assign w8568 = ~w8540 & w8567;
assign w8569 = w8540 & ~w8567;
assign v4063 = ~(w8568 | w8569);
assign w8570 = v4063;
assign w8571 = (~w8405 & ~w8407) | (~w8405 & w17784) | (~w8407 & w17784);
assign w8572 = (~w8335 & ~w8337) | (~w8335 & w17588) | (~w8337 & w17588);
assign v4064 = ~(w8571 | w8572);
assign w8573 = v4064;
assign w8574 = w8571 & w8572;
assign v4065 = ~(w8573 | w8574);
assign w8575 = v4065;
assign v4066 = ~(w8570 | w8575);
assign w8576 = v4066;
assign w8577 = w8570 & w8575;
assign v4067 = ~(w8576 | w8577);
assign w8578 = v4067;
assign w8579 = ~w8539 & w8578;
assign w8580 = w8539 & ~w8578;
assign v4068 = ~(w8579 | w8580);
assign w8581 = v4068;
assign w8582 = ~w8538 & w8581;
assign w8583 = w8538 & ~w8581;
assign v4069 = ~(w8582 | w8583);
assign w8584 = v4069;
assign w8585 = ~w8537 & w8584;
assign w8586 = w8537 & ~w8584;
assign v4070 = ~(w8585 | w8586);
assign w8587 = v4070;
assign v4071 = ~(w8490 | w8496);
assign w8588 = v4071;
assign w8589 = (~w8279 & ~w8281) | (~w8279 & w17785) | (~w8281 & w17785);
assign w8590 = (~w8478 & ~w8480) | (~w8478 & w17786) | (~w8480 & w17786);
assign v4072 = ~(w8589 | w8590);
assign w8591 = v4072;
assign w8592 = w8589 & w8590;
assign v4073 = ~(w8591 | w8592);
assign w8593 = v4073;
assign w8594 = w8588 & ~w8593;
assign w8595 = ~w8588 & w8593;
assign v4074 = ~(w8594 | w8595);
assign w8596 = v4074;
assign w8597 = (~w8498 & ~w8500) | (~w8498 & w17787) | (~w8500 & w17787);
assign w8598 = (~w8289 & ~w8290) | (~w8289 & w17788) | (~w8290 & w17788);
assign v4075 = ~(w8597 | w8598);
assign w8599 = v4075;
assign w8600 = w8597 & w8598;
assign v4076 = ~(w8599 | w8600);
assign w8601 = v4076;
assign v4077 = ~(w8596 | w8601);
assign w8602 = v4077;
assign w8603 = w8596 & w8601;
assign v4078 = ~(w8602 | w8603);
assign w8604 = v4078;
assign v4079 = ~(w8506 | w8510);
assign w8605 = v4079;
assign w8606 = pi29 & pi36;
assign w8607 = pi11 & pi54;
assign v4080 = ~(w8385 | w8607);
assign w8608 = v4080;
assign w8609 = w8385 & w8607;
assign v4081 = ~(w8608 | w8609);
assign w8610 = v4081;
assign w8611 = w8606 & ~w8610;
assign w8612 = ~w8606 & w8610;
assign v4082 = ~(w8611 | w8612);
assign w8613 = v4082;
assign w8614 = pi30 & pi35;
assign w8615 = pi31 & pi34;
assign w8616 = pi32 & pi33;
assign v4083 = ~(w8615 | w8616);
assign w8617 = v4083;
assign w8618 = w8615 & w8616;
assign v4084 = ~(w8617 | w8618);
assign w8619 = v4084;
assign w8620 = w8614 & ~w8619;
assign w8621 = ~w8614 & w8619;
assign v4085 = ~(w8620 | w8621);
assign w8622 = v4085;
assign v4086 = ~(w8613 | w8622);
assign w8623 = v4086;
assign w8624 = w8613 & w8622;
assign v4087 = ~(w8623 | w8624);
assign w8625 = v4087;
assign w8626 = pi17 & pi48;
assign w8627 = pi03 & pi62;
assign v4088 = ~(pi33 | w8627);
assign w8628 = v4088;
assign w8629 = pi33 & w8627;
assign v4089 = ~(w8628 | w8629);
assign w8630 = v4089;
assign w8631 = w8626 & ~w8630;
assign w8632 = ~w8626 & w8630;
assign v4090 = ~(w8631 | w8632);
assign w8633 = v4090;
assign w8634 = w8625 & ~w8633;
assign w8635 = ~w8625 & w8633;
assign v4091 = ~(w8634 | w8635);
assign w8636 = v4091;
assign w8637 = (~w8303 & ~w8300) | (~w8303 & w16758) | (~w8300 & w16758);
assign w8638 = pi08 & pi57;
assign w8639 = pi21 & pi44;
assign v4092 = ~(w8411 | w8639);
assign w8640 = v4092;
assign w8641 = pi22 & pi44;
assign w8642 = w8409 & w8641;
assign v4093 = ~(w8640 | w8642);
assign w8643 = v4093;
assign w8644 = w8638 & ~w8643;
assign w8645 = ~w8638 & w8643;
assign v4094 = ~(w8644 | w8645);
assign w8646 = v4094;
assign v4095 = ~(w8637 | w8646);
assign w8647 = v4095;
assign w8648 = w8637 & w8646;
assign v4096 = ~(w8647 | w8648);
assign w8649 = v4096;
assign w8650 = pi05 & pi60;
assign w8651 = pi06 & pi59;
assign w8652 = pi07 & pi58;
assign v4097 = ~(w8651 | w8652);
assign w8653 = v4097;
assign w8654 = pi07 & pi59;
assign w8655 = w8417 & w8654;
assign v4098 = ~(w8653 | w8655);
assign w8656 = v4098;
assign w8657 = w8650 & ~w8656;
assign w8658 = ~w8650 & w8656;
assign v4099 = ~(w8657 | w8658);
assign w8659 = v4099;
assign w8660 = w8649 & ~w8659;
assign w8661 = ~w8649 & w8659;
assign v4100 = ~(w8660 | w8661);
assign w8662 = v4100;
assign w8663 = w8636 & w8662;
assign v4101 = ~(w8636 | w8662);
assign w8664 = v4101;
assign v4102 = ~(w8663 | w8664);
assign w8665 = v4102;
assign w8666 = pi23 & pi42;
assign w8667 = pi25 & pi40;
assign w8668 = pi24 & pi41;
assign v4103 = ~(w8667 | w8668);
assign w8669 = v4103;
assign w8670 = pi25 & pi41;
assign w8671 = w8430 & w8670;
assign v4104 = ~(w8669 | w8671);
assign w8672 = v4104;
assign w8673 = w8666 & ~w8672;
assign w8674 = ~w8666 & w8672;
assign v4105 = ~(w8673 | w8674);
assign w8675 = v4105;
assign w8676 = pi09 & pi56;
assign w8677 = pi10 & pi55;
assign w8678 = pi20 & pi45;
assign v4106 = ~(w8677 | w8678);
assign w8679 = v4106;
assign w8680 = w8677 & w8678;
assign v4107 = ~(w8679 | w8680);
assign w8681 = v4107;
assign w8682 = w8676 & ~w8681;
assign w8683 = ~w8676 & w8681;
assign v4108 = ~(w8682 | w8683);
assign w8684 = v4108;
assign v4109 = ~(w8675 | w8684);
assign w8685 = v4109;
assign w8686 = w8675 & w8684;
assign v4110 = ~(w8685 | w8686);
assign w8687 = v4110;
assign w8688 = pi26 & pi39;
assign w8689 = pi28 & pi37;
assign w8690 = pi27 & pi38;
assign v4111 = ~(w8689 | w8690);
assign w8691 = v4111;
assign w8692 = pi28 & pi38;
assign w8693 = w8357 & w8692;
assign v4112 = ~(w8691 | w8693);
assign w8694 = v4112;
assign w8695 = w8688 & ~w8694;
assign w8696 = ~w8688 & w8694;
assign v4113 = ~(w8695 | w8696);
assign w8697 = v4113;
assign w8698 = w8687 & ~w8697;
assign w8699 = ~w8687 & w8697;
assign v4114 = ~(w8698 | w8699);
assign w8700 = v4114;
assign w8701 = w8665 & w8700;
assign v4115 = ~(w8665 | w8700);
assign w8702 = v4115;
assign v4116 = ~(w8701 | w8702);
assign w8703 = v4116;
assign w8704 = ~w8605 & w8703;
assign w8705 = w8605 & ~w8703;
assign v4117 = ~(w8704 | w8705);
assign w8706 = v4117;
assign w8707 = w8604 & w8706;
assign v4118 = ~(w8604 | w8706);
assign w8708 = v4118;
assign v4119 = ~(w8707 | w8708);
assign w8709 = v4119;
assign v4120 = ~(w8512 | w8515);
assign w8710 = v4120;
assign w8711 = pi02 & pi63;
assign v4121 = ~(w8396 | w8711);
assign w8712 = v4121;
assign w8713 = w8396 & w8711;
assign v4122 = ~(w8712 | w8713);
assign w8714 = v4122;
assign v4123 = ~(w8368 | w8372);
assign w8715 = v4123;
assign v4124 = ~(w8371 | w8715);
assign w8716 = v4124;
assign w8717 = w8714 & w8716;
assign v4125 = ~(w8714 | w8716);
assign w8718 = v4125;
assign v4126 = ~(w8717 | w8718);
assign w8719 = v4126;
assign w8720 = pi16 & pi49;
assign w8721 = pi15 & pi50;
assign w8722 = pi14 & pi51;
assign v4127 = ~(w8721 | w8722);
assign w8723 = v4127;
assign w8724 = pi15 & pi51;
assign w8725 = w8368 & w8724;
assign v4128 = ~(w8723 | w8725);
assign w8726 = v4128;
assign w8727 = w8720 & ~w8726;
assign w8728 = ~w8720 & w8726;
assign v4129 = ~(w8727 | w8728);
assign w8729 = v4129;
assign w8730 = pi13 & pi52;
assign w8731 = pi18 & pi47;
assign v4130 = ~(w8730 | w8731);
assign w8732 = v4130;
assign w8733 = w8730 & w8731;
assign v4131 = ~(w8732 | w8733);
assign w8734 = v4131;
assign w8735 = w8312 & ~w8734;
assign w8736 = ~w8312 & w8734;
assign v4132 = ~(w8735 | w8736);
assign w8737 = v4132;
assign v4133 = ~(w8729 | w8737);
assign w8738 = v4133;
assign w8739 = w8729 & w8737;
assign v4134 = ~(w8738 | w8739);
assign w8740 = v4134;
assign w8741 = w8719 & w8740;
assign v4135 = ~(w8719 | w8740);
assign w8742 = v4135;
assign v4136 = ~(w8741 | w8742);
assign w8743 = v4136;
assign w8744 = (~w8450 & ~w8452) | (~w8450 & w16918) | (~w8452 & w16918);
assign v4137 = ~(w8391 | w8402);
assign w8745 = v4137;
assign v4138 = ~(w8744 | w8745);
assign w8746 = v4138;
assign w8747 = w8744 & w8745;
assign v4139 = ~(w8746 | w8747);
assign w8748 = v4139;
assign v4140 = ~(w8743 | w8748);
assign w8749 = v4140;
assign w8750 = w8743 & w8748;
assign v4141 = ~(w8749 | w8750);
assign w8751 = v4141;
assign v4142 = ~(w8357 | w8360);
assign w8752 = v4142;
assign v4143 = ~(w8359 | w8752);
assign w8753 = v4143;
assign w8754 = w8408 & ~w8410;
assign v4144 = ~(w8412 | w8754);
assign w8755 = v4144;
assign w8756 = w8753 & ~w8755;
assign w8757 = ~w8753 & w8755;
assign v4145 = ~(w8756 | w8757);
assign w8758 = v4145;
assign w8759 = w8178 & ~w8311;
assign v4146 = ~(w8313 | w8759);
assign w8760 = v4146;
assign w8761 = ~w8758 & w8760;
assign w8762 = w8758 & ~w8760;
assign v4147 = ~(w8761 | w8762);
assign w8763 = v4147;
assign w8764 = (~w8365 & ~w8367) | (~w8365 & w16919) | (~w8367 & w16919);
assign w8765 = ~w8763 & w8764;
assign w8766 = w8763 & ~w8764;
assign v4148 = ~(w8765 | w8766);
assign w8767 = v4148;
assign w8768 = (~w8426 & ~w8428) | (~w8426 & w17589) | (~w8428 & w17589);
assign w8769 = ~w8767 & w8768;
assign w8770 = w8767 & ~w8768;
assign v4149 = ~(w8769 | w8770);
assign w8771 = v4149;
assign w8772 = (~w8458 & ~w8460) | (~w8458 & w17153) | (~w8460 & w17153);
assign w8773 = ~w8771 & w8772;
assign w8774 = w8771 & ~w8772;
assign v4150 = ~(w8773 | w8774);
assign w8775 = v4150;
assign w8776 = w8751 & w8775;
assign v4151 = ~(w8751 | w8775);
assign w8777 = v4151;
assign v4152 = ~(w8776 | w8777);
assign w8778 = v4152;
assign w8779 = ~w8710 & w8778;
assign w8780 = w8710 & ~w8778;
assign v4153 = ~(w8779 | w8780);
assign w8781 = v4153;
assign w8782 = w8709 & w8781;
assign v4154 = ~(w8709 | w8781);
assign w8783 = v4154;
assign v4155 = ~(w8782 | w8783);
assign w8784 = v4155;
assign w8785 = w8587 & w8784;
assign v4156 = ~(w8587 | w8784);
assign w8786 = v4156;
assign v4157 = ~(w8785 | w8786);
assign w8787 = v4157;
assign w8788 = ~w8536 & w8787;
assign w8789 = w8536 & ~w8787;
assign v4158 = ~(w8788 | w8789);
assign w8790 = v4158;
assign w8791 = w8535 & w8790;
assign v4159 = ~(w8535 | w8790);
assign w8792 = v4159;
assign v4160 = ~(w8791 | w8792);
assign w8793 = v4160;
assign v4161 = ~(w8525 | w8788);
assign w8794 = v4161;
assign w8795 = (~w7006 & w17789) | (~w7006 & w17790) | (w17789 & w17790);
assign v4162 = ~(w8585 | w8785);
assign w8796 = v4162;
assign w8797 = (~w8573 & ~w8575) | (~w8573 & w17791) | (~w8575 & w17791);
assign w8798 = pi03 & pi63;
assign w8799 = pi05 & pi61;
assign w8800 = pi04 & pi62;
assign v4163 = ~(w8799 | w8800);
assign w8801 = v4163;
assign w8802 = pi05 & pi62;
assign w8803 = w8396 & w8802;
assign v4164 = ~(w8801 | w8803);
assign w8804 = v4164;
assign w8805 = w8798 & ~w8804;
assign w8806 = ~w8798 & w8804;
assign v4165 = ~(w8805 | w8806);
assign w8807 = v4165;
assign w8808 = pi27 & pi39;
assign w8809 = pi29 & pi37;
assign v4166 = ~(w8692 | w8809);
assign w8810 = v4166;
assign w8811 = pi29 & pi38;
assign w8812 = w8689 & w8811;
assign v4167 = ~(w8810 | w8812);
assign w8813 = v4167;
assign w8814 = w8808 & ~w8813;
assign w8815 = ~w8808 & w8813;
assign v4168 = ~(w8814 | w8815);
assign w8816 = v4168;
assign v4169 = ~(w8807 | w8816);
assign w8817 = v4169;
assign w8818 = w8807 & w8816;
assign v4170 = ~(w8817 | w8818);
assign w8819 = v4170;
assign w8820 = pi11 & pi55;
assign w8821 = pi19 & pi47;
assign w8822 = pi12 & pi54;
assign v4171 = ~(w8821 | w8822);
assign w8823 = v4171;
assign w8824 = w8821 & w8822;
assign v4172 = ~(w8823 | w8824);
assign w8825 = v4172;
assign w8826 = w8820 & ~w8825;
assign w8827 = ~w8820 & w8825;
assign v4173 = ~(w8826 | w8827);
assign w8828 = v4173;
assign w8829 = w8819 & ~w8828;
assign w8830 = ~w8819 & w8828;
assign v4174 = ~(w8829 | w8830);
assign w8831 = v4174;
assign w8832 = pi20 & pi46;
assign w8833 = pi21 & pi45;
assign v4175 = ~(w8641 | w8833);
assign w8834 = v4175;
assign w8835 = pi22 & pi45;
assign w8836 = w8639 & w8835;
assign v4176 = ~(w8834 | w8836);
assign w8837 = v4176;
assign w8838 = w8832 & ~w8837;
assign w8839 = ~w8832 & w8837;
assign v4177 = ~(w8838 | w8839);
assign w8840 = v4177;
assign w8841 = pi23 & pi43;
assign w8842 = pi09 & pi57;
assign w8843 = pi24 & pi42;
assign v4178 = ~(w8842 | w8843);
assign w8844 = v4178;
assign w8845 = w8842 & w8843;
assign v4179 = ~(w8844 | w8845);
assign w8846 = v4179;
assign w8847 = w8841 & ~w8846;
assign w8848 = ~w8841 & w8846;
assign v4180 = ~(w8847 | w8848);
assign w8849 = v4180;
assign v4181 = ~(w8840 | w8849);
assign w8850 = v4181;
assign w8851 = w8840 & w8849;
assign v4182 = ~(w8850 | w8851);
assign w8852 = v4182;
assign w8853 = pi10 & pi56;
assign w8854 = pi26 & pi40;
assign v4183 = ~(w8670 | w8854);
assign w8855 = v4183;
assign w8856 = pi26 & pi41;
assign w8857 = w8667 & w8856;
assign v4184 = ~(w8855 | w8857);
assign w8858 = v4184;
assign w8859 = w8853 & ~w8858;
assign w8860 = ~w8853 & w8858;
assign v4185 = ~(w8859 | w8860);
assign w8861 = v4185;
assign w8862 = w8852 & ~w8861;
assign w8863 = ~w8852 & w8861;
assign v4186 = ~(w8862 | w8863);
assign w8864 = v4186;
assign w8865 = pi14 & pi52;
assign w8866 = pi31 & pi35;
assign w8867 = pi30 & pi36;
assign v4187 = ~(w8866 | w8867);
assign w8868 = v4187;
assign w8869 = w8866 & w8867;
assign v4188 = ~(w8868 | w8869);
assign w8870 = v4188;
assign w8871 = w8865 & ~w8870;
assign w8872 = ~w8865 & w8870;
assign v4189 = ~(w8871 | w8872);
assign w8873 = v4189;
assign w8874 = pi18 & pi48;
assign w8875 = pi13 & pi53;
assign v4190 = ~(w8724 | w8875);
assign w8876 = v4190;
assign w8877 = w8724 & w8875;
assign v4191 = ~(w8876 | w8877);
assign w8878 = v4191;
assign w8879 = w8874 & ~w8878;
assign w8880 = ~w8874 & w8878;
assign v4192 = ~(w8879 | w8880);
assign w8881 = v4192;
assign v4193 = ~(w8873 | w8881);
assign w8882 = v4193;
assign w8883 = w8873 & w8881;
assign v4194 = ~(w8882 | w8883);
assign w8884 = v4194;
assign w8885 = pi32 & pi34;
assign w8886 = pi17 & pi49;
assign w8887 = pi16 & pi50;
assign v4195 = ~(w8886 | w8887);
assign w8888 = v4195;
assign w8889 = pi17 & pi50;
assign w8890 = w8720 & w8889;
assign v4196 = ~(w8888 | w8890);
assign w8891 = v4196;
assign w8892 = w8885 & ~w8891;
assign w8893 = ~w8885 & w8891;
assign v4197 = ~(w8892 | w8893);
assign w8894 = v4197;
assign w8895 = w8884 & ~w8894;
assign w8896 = ~w8884 & w8894;
assign v4198 = ~(w8895 | w8896);
assign w8897 = v4198;
assign w8898 = w8864 & w8897;
assign v4199 = ~(w8864 | w8897);
assign w8899 = v4199;
assign v4200 = ~(w8898 | w8899);
assign w8900 = v4200;
assign w8901 = w8831 & w8900;
assign v4201 = ~(w8831 | w8900);
assign w8902 = v4201;
assign v4202 = ~(w8901 | w8902);
assign w8903 = v4202;
assign w8904 = ~w8797 & w8903;
assign w8905 = w8797 & ~w8903;
assign v4203 = ~(w8904 | w8905);
assign w8906 = v4203;
assign v4204 = ~(w8756 | w8762);
assign w8907 = v4204;
assign w8908 = (~w8545 & ~w8547) | (~w8545 & w17792) | (~w8547 & w17792);
assign w8909 = (~w8557 & ~w8559) | (~w8557 & w17793) | (~w8559 & w17793);
assign v4205 = ~(w8908 | w8909);
assign w8910 = v4205;
assign w8911 = w8908 & w8909;
assign v4206 = ~(w8910 | w8911);
assign w8912 = v4206;
assign w8913 = w8907 & ~w8912;
assign w8914 = ~w8907 & w8912;
assign v4207 = ~(w8913 | w8914);
assign w8915 = v4207;
assign w8916 = (~w8565 & ~w8567) | (~w8565 & w17154) | (~w8567 & w17154);
assign w8917 = (~w8766 & ~w8767) | (~w8766 & w17155) | (~w8767 & w17155);
assign v4208 = ~(w8916 | w8917);
assign w8918 = v4208;
assign w8919 = w8916 & w8917;
assign v4209 = ~(w8918 | w8919);
assign w8920 = v4209;
assign v4210 = ~(w8915 | w8920);
assign w8921 = v4210;
assign w8922 = w8915 & w8920;
assign v4211 = ~(w8921 | w8922);
assign w8923 = v4211;
assign w8924 = w8906 & w8923;
assign v4212 = ~(w8906 | w8923);
assign w8925 = v4212;
assign v4213 = ~(w8924 | w8925);
assign w8926 = v4213;
assign v4214 = ~(w8579 | w8582);
assign w8927 = v4214;
assign v4215 = ~(w8704 | w8707);
assign w8928 = v4215;
assign v4216 = ~(w8927 | w8928);
assign w8929 = v4216;
assign w8930 = w8927 & w8928;
assign v4217 = ~(w8929 | w8930);
assign w8931 = v4217;
assign w8932 = w8926 & w8931;
assign v4218 = ~(w8926 | w8931);
assign w8933 = v4218;
assign v4219 = ~(w8932 | w8933);
assign w8934 = v4219;
assign v4220 = ~(w8779 | w8782);
assign w8935 = v4220;
assign v4221 = ~(w8599 | w8603);
assign w8936 = v4221;
assign v4222 = ~(w8591 | w8595);
assign w8937 = v4222;
assign w8938 = (~w8713 & ~w8716) | (~w8713 & w17156) | (~w8716 & w17156);
assign w8939 = w8688 & ~w8691;
assign v4223 = ~(w8693 | w8939);
assign w8940 = v4223;
assign v4224 = ~(w8938 | w8940);
assign w8941 = v4224;
assign w8942 = w8938 & w8940;
assign v4225 = ~(w8941 | w8942);
assign w8943 = v4225;
assign w8944 = pi06 & pi60;
assign w8945 = pi08 & pi58;
assign v4226 = ~(w8654 | w8945);
assign w8946 = v4226;
assign w8947 = pi08 & pi59;
assign w8948 = w8652 & w8947;
assign v4227 = ~(w8946 | w8948);
assign w8949 = v4227;
assign w8950 = w8944 & ~w8949;
assign w8951 = ~w8944 & w8949;
assign v4228 = ~(w8950 | w8951);
assign w8952 = v4228;
assign w8953 = ~w8943 & w8952;
assign w8954 = w8943 & ~w8952;
assign v4229 = ~(w8953 | w8954);
assign w8955 = v4229;
assign v4230 = ~(w8738 | w8741);
assign w8956 = v4230;
assign w8957 = w8955 & ~w8956;
assign w8958 = ~w8955 & w8956;
assign v4231 = ~(w8957 | w8958);
assign w8959 = v4231;
assign w8960 = w8937 & ~w8959;
assign w8961 = ~w8937 & w8959;
assign v4232 = ~(w8960 | w8961);
assign w8962 = v4232;
assign v4233 = ~(w8614 | w8618);
assign w8963 = v4233;
assign v4234 = ~(w8617 | w8963);
assign w8964 = v4234;
assign v4235 = ~(w8626 | w8629);
assign w8965 = v4235;
assign v4236 = ~(w8628 | w8965);
assign w8966 = v4236;
assign w8967 = w8964 & w8966;
assign v4237 = ~(w8964 | w8966);
assign w8968 = v4237;
assign v4238 = ~(w8967 | w8968);
assign w8969 = v4238;
assign w8970 = w8720 & ~w8723;
assign v4239 = ~(w8725 | w8970);
assign w8971 = v4239;
assign w8972 = ~w8969 & w8971;
assign w8973 = w8969 & ~w8971;
assign v4240 = ~(w8972 | w8973);
assign w8974 = v4240;
assign w8975 = w8638 & ~w8640;
assign v4241 = ~(w8642 | w8975);
assign w8976 = v4241;
assign w8977 = w8650 & ~w8653;
assign v4242 = ~(w8655 | w8977);
assign w8978 = v4242;
assign v4243 = ~(w8976 | w8978);
assign w8979 = v4243;
assign w8980 = w8976 & w8978;
assign v4244 = ~(w8979 | w8980);
assign w8981 = v4244;
assign v4245 = ~(w8606 | w8609);
assign w8982 = v4245;
assign v4246 = ~(w8608 | w8982);
assign w8983 = v4246;
assign v4247 = ~(w8981 | w8983);
assign w8984 = v4247;
assign w8985 = w8981 & w8983;
assign v4248 = ~(w8984 | w8985);
assign w8986 = v4248;
assign w8987 = (~w8623 & ~w8625) | (~w8623 & w16920) | (~w8625 & w16920);
assign w8988 = ~w8986 & w8987;
assign w8989 = w8986 & ~w8987;
assign v4249 = ~(w8988 | w8989);
assign w8990 = v4249;
assign w8991 = w8974 & w8990;
assign v4250 = ~(w8974 | w8990);
assign w8992 = v4250;
assign v4251 = ~(w8991 | w8992);
assign w8993 = v4251;
assign w8994 = w8962 & w8993;
assign v4252 = ~(w8962 | w8993);
assign w8995 = v4252;
assign v4253 = ~(w8994 | w8995);
assign w8996 = v4253;
assign w8997 = ~w8936 & w8996;
assign w8998 = w8936 & ~w8996;
assign v4254 = ~(w8997 | w8998);
assign w8999 = v4254;
assign w9000 = (~w8774 & ~w8775) | (~w8774 & w17590) | (~w8775 & w17590);
assign v4255 = ~(w8676 | w8680);
assign w9001 = v4255;
assign v4256 = ~(w8679 | w9001);
assign w9002 = v4256;
assign v4257 = ~(w8312 | w8733);
assign w9003 = v4257;
assign v4258 = ~(w8732 | w9003);
assign w9004 = v4258;
assign w9005 = w9002 & w9004;
assign v4259 = ~(w9002 | w9004);
assign w9006 = v4259;
assign v4260 = ~(w9005 | w9006);
assign w9007 = v4260;
assign w9008 = w8666 & ~w8669;
assign v4261 = ~(w8671 | w9008);
assign w9009 = v4261;
assign w9010 = ~w9007 & w9009;
assign w9011 = w9007 & ~w9009;
assign v4262 = ~(w9010 | w9011);
assign w9012 = v4262;
assign w9013 = (~w8647 & ~w8649) | (~w8647 & w16921) | (~w8649 & w16921);
assign w9014 = ~w9012 & w9013;
assign w9015 = w9012 & ~w9013;
assign v4263 = ~(w9014 | w9015);
assign w9016 = v4263;
assign w9017 = (~w8685 & ~w8687) | (~w8685 & w17591) | (~w8687 & w17591);
assign w9018 = ~w9016 & w9017;
assign w9019 = w9016 & ~w9017;
assign v4264 = ~(w9018 | w9019);
assign w9020 = v4264;
assign w9021 = (~w8663 & ~w8665) | (~w8663 & w17592) | (~w8665 & w17592);
assign w9022 = (~w8746 & ~w8748) | (~w8746 & w17157) | (~w8748 & w17157);
assign v4265 = ~(w9021 | w9022);
assign w9023 = v4265;
assign w9024 = w9021 & w9022;
assign v4266 = ~(w9023 | w9024);
assign w9025 = v4266;
assign w9026 = w9020 & w9025;
assign v4267 = ~(w9020 | w9025);
assign w9027 = v4267;
assign v4268 = ~(w9026 | w9027);
assign w9028 = v4268;
assign w9029 = ~w9000 & w9028;
assign w9030 = w9000 & ~w9028;
assign v4269 = ~(w9029 | w9030);
assign w9031 = v4269;
assign v4270 = ~(w8999 | w9031);
assign w9032 = v4270;
assign w9033 = w8999 & w9031;
assign v4271 = ~(w9032 | w9033);
assign w9034 = v4271;
assign w9035 = ~w8935 & w9034;
assign w9036 = w8935 & ~w9034;
assign v4272 = ~(w9035 | w9036);
assign w9037 = v4272;
assign w9038 = w8934 & w9037;
assign v4273 = ~(w8934 | w9037);
assign w9039 = v4273;
assign v4274 = ~(w9038 | w9039);
assign w9040 = v4274;
assign w9041 = ~w8796 & w9040;
assign w9042 = w8796 & ~w9040;
assign v4275 = ~(w9041 | w9042);
assign w9043 = v4275;
assign w9044 = w8795 & ~w9043;
assign w9045 = ~w8795 & w9043;
assign v4276 = ~(w9044 | w9045);
assign w9046 = v4276;
assign v4277 = ~(w9035 | w9038);
assign w9047 = v4277;
assign v4278 = ~(w8929 | w8932);
assign w9048 = v4278;
assign v4279 = ~(w8994 | w8997);
assign w9049 = v4279;
assign w9050 = (~w8918 & ~w8920) | (~w8918 & w17593) | (~w8920 & w17593);
assign v4280 = ~(w8817 | w8829);
assign w9051 = v4280;
assign w9052 = (~w8850 & ~w8852) | (~w8850 & w17594) | (~w8852 & w17594);
assign w9053 = (~w8941 & ~w8943) | (~w8941 & w17595) | (~w8943 & w17595);
assign v4281 = ~(w9052 | w9053);
assign w9054 = v4281;
assign w9055 = w9052 & w9053;
assign v4282 = ~(w9054 | w9055);
assign w9056 = v4282;
assign w9057 = w9051 & ~w9056;
assign w9058 = ~w9051 & w9056;
assign v4283 = ~(w9057 | w9058);
assign w9059 = v4283;
assign w9060 = w8798 & ~w8801;
assign v4284 = ~(w8803 | w9060);
assign w9061 = v4284;
assign w9062 = w8944 & ~w8946;
assign v4285 = ~(w8948 | w9062);
assign w9063 = v4285;
assign v4286 = ~(w9061 | w9063);
assign w9064 = v4286;
assign w9065 = w9061 & w9063;
assign v4287 = ~(w9064 | w9065);
assign w9066 = v4287;
assign w9067 = w8808 & ~w8810;
assign v4288 = ~(w8812 | w9067);
assign w9068 = v4288;
assign w9069 = ~w9066 & w9068;
assign w9070 = w9066 & ~w9068;
assign v4289 = ~(w9069 | w9070);
assign w9071 = v4289;
assign v4290 = ~(w8841 | w8845);
assign w9072 = v4290;
assign v4291 = ~(w8844 | w9072);
assign w9073 = v4291;
assign w9074 = w8853 & ~w8855;
assign v4292 = ~(w8857 | w9074);
assign w9075 = v4292;
assign w9076 = w9073 & ~w9075;
assign w9077 = ~w9073 & w9075;
assign v4293 = ~(w9076 | w9077);
assign w9078 = v4293;
assign w9079 = w8832 & ~w8834;
assign v4294 = ~(w8836 | w9079);
assign w9080 = v4294;
assign w9081 = ~w9078 & w9080;
assign w9082 = w9078 & ~w9080;
assign v4295 = ~(w9081 | w9082);
assign w9083 = v4295;
assign w9084 = pi06 & pi61;
assign w9085 = w8885 & ~w8888;
assign w9086 = (w9084 & w9085) | (w9084 & w16759) | (w9085 & w16759);
assign w9087 = ~w9085 & w16760;
assign v4296 = ~(w9086 | w9087);
assign w9088 = v4296;
assign v4297 = ~(w8865 | w8869);
assign w9089 = v4297;
assign v4298 = ~(w8868 | w9089);
assign w9090 = v4298;
assign v4299 = ~(w9088 | w9090);
assign w9091 = v4299;
assign w9092 = w9088 & w9090;
assign v4300 = ~(w9091 | w9092);
assign w9093 = v4300;
assign w9094 = w9083 & w9093;
assign v4301 = ~(w9083 | w9093);
assign w9095 = v4301;
assign v4302 = ~(w9094 | w9095);
assign w9096 = v4302;
assign w9097 = w9071 & w9096;
assign v4303 = ~(w9071 | w9096);
assign w9098 = v4303;
assign v4304 = ~(w9097 | w9098);
assign w9099 = v4304;
assign w9100 = w9059 & w9099;
assign v4305 = ~(w9059 | w9099);
assign w9101 = v4305;
assign v4306 = ~(w9100 | w9101);
assign w9102 = v4306;
assign w9103 = ~w9050 & w9102;
assign w9104 = w9050 & ~w9102;
assign v4307 = ~(w9103 | w9104);
assign w9105 = v4307;
assign w9106 = ~w9049 & w9105;
assign w9107 = w9049 & ~w9105;
assign v4308 = ~(w9106 | w9107);
assign w9108 = v4308;
assign v4309 = ~(w8910 | w8914);
assign w9109 = v4309;
assign v4310 = ~(w8874 | w8877);
assign w9110 = v4310;
assign v4311 = ~(w8876 | w9110);
assign w9111 = v4311;
assign v4312 = ~(w8820 | w8824);
assign w9112 = v4312;
assign v4313 = ~(w8823 | w9112);
assign w9113 = v4313;
assign w9114 = w9111 & w9113;
assign v4314 = ~(w9111 | w9113);
assign w9115 = v4314;
assign v4315 = ~(w9114 | w9115);
assign w9116 = v4315;
assign w9117 = pi10 & pi57;
assign w9118 = pi11 & pi56;
assign w9119 = pi20 & pi47;
assign v4316 = ~(w9118 | w9119);
assign w9120 = v4316;
assign w9121 = w9118 & w9119;
assign v4317 = ~(w9120 | w9121);
assign w9122 = v4317;
assign w9123 = w9117 & ~w9122;
assign w9124 = ~w9117 & w9122;
assign v4318 = ~(w9123 | w9124);
assign w9125 = v4318;
assign w9126 = ~w9116 & w9125;
assign w9127 = w9116 & ~w9125;
assign v4319 = ~(w9126 | w9127);
assign w9128 = v4319;
assign v4320 = ~(w8882 | w8895);
assign w9129 = v4320;
assign w9130 = w9128 & ~w9129;
assign w9131 = ~w9128 & w9129;
assign v4321 = ~(w9130 | w9131);
assign w9132 = v4321;
assign w9133 = w9109 & ~w9132;
assign w9134 = ~w9109 & w9132;
assign v4322 = ~(w9133 | w9134);
assign w9135 = v4322;
assign v4323 = ~(w8898 | w8901);
assign w9136 = v4323;
assign v4324 = ~(w8957 | w8961);
assign w9137 = v4324;
assign v4325 = ~(w9136 | w9137);
assign w9138 = v4325;
assign w9139 = w9136 & w9137;
assign v4326 = ~(w9138 | w9139);
assign w9140 = v4326;
assign w9141 = w9135 & w9140;
assign v4327 = ~(w9135 | w9140);
assign w9142 = v4327;
assign v4328 = ~(w9141 | w9142);
assign w9143 = v4328;
assign w9144 = w9108 & w9143;
assign v4329 = ~(w9108 | w9143);
assign w9145 = v4329;
assign v4330 = ~(w9144 | w9145);
assign w9146 = v4330;
assign w9147 = ~w9048 & w9146;
assign w9148 = w9048 & ~w9146;
assign v4331 = ~(w9147 | w9148);
assign w9149 = v4331;
assign w9150 = pi19 & pi48;
assign w9151 = pi14 & pi53;
assign v4332 = ~(w8889 | w9151);
assign w9152 = v4332;
assign w9153 = w8889 & w9151;
assign v4333 = ~(w9152 | w9153);
assign w9154 = v4333;
assign w9155 = w9150 & ~w9154;
assign w9156 = ~w9150 & w9154;
assign v4334 = ~(w9155 | w9156);
assign w9157 = v4334;
assign w9158 = pi25 & pi42;
assign w9159 = pi21 & pi46;
assign v4335 = ~(w8856 | w9159);
assign w9160 = v4335;
assign w9161 = w8856 & w9159;
assign v4336 = ~(w9160 | w9161);
assign w9162 = v4336;
assign w9163 = w9158 & ~w9162;
assign w9164 = ~w9158 & w9162;
assign v4337 = ~(w9163 | w9164);
assign w9165 = v4337;
assign v4338 = ~(w9157 | w9165);
assign w9166 = v4338;
assign w9167 = w9157 & w9165;
assign v4339 = ~(w9166 | w9167);
assign w9168 = v4339;
assign w9169 = pi04 & pi63;
assign w9170 = pi27 & pi40;
assign w9171 = pi28 & pi39;
assign v4340 = ~(w9170 | w9171);
assign w9172 = v4340;
assign w9173 = w9170 & w9171;
assign v4341 = ~(w9172 | w9173);
assign w9174 = v4341;
assign w9175 = w9169 & ~w9174;
assign w9176 = ~w9169 & w9174;
assign v4342 = ~(w9175 | w9176);
assign w9177 = v4342;
assign w9178 = w9168 & ~w9177;
assign w9179 = ~w9168 & w9177;
assign v4343 = ~(w9178 | w9179);
assign w9180 = v4343;
assign w9181 = pi18 & pi49;
assign w9182 = pi62 & w3094;
assign v4344 = ~(pi34 | w8802);
assign w9183 = v4344;
assign v4345 = ~(w9182 | w9183);
assign w9184 = v4345;
assign w9185 = w9181 & ~w9184;
assign w9186 = ~w9181 & w9184;
assign v4346 = ~(w9185 | w9186);
assign w9187 = v4346;
assign w9188 = pi31 & pi36;
assign w9189 = pi33 & pi34;
assign w9190 = pi32 & pi35;
assign v4347 = ~(w9189 | w9190);
assign w9191 = v4347;
assign w9192 = pi33 & pi35;
assign w9193 = w8885 & w9192;
assign v4348 = ~(w9191 | w9193);
assign w9194 = v4348;
assign w9195 = w9188 & ~w9194;
assign w9196 = ~w9188 & w9194;
assign v4349 = ~(w9195 | w9196);
assign w9197 = v4349;
assign v4350 = ~(w9187 | w9197);
assign w9198 = v4350;
assign w9199 = w9187 & w9197;
assign v4351 = ~(w9198 | w9199);
assign w9200 = v4351;
assign w9201 = pi12 & pi55;
assign w9202 = pi13 & pi54;
assign v4352 = ~(w9201 | w9202);
assign w9203 = v4352;
assign w9204 = pi13 & pi55;
assign w9205 = w8822 & w9204;
assign v4353 = ~(w9203 | w9205);
assign w9206 = v4353;
assign w9207 = w8811 & ~w9206;
assign w9208 = ~w8811 & w9206;
assign v4354 = ~(w9207 | w9208);
assign w9209 = v4354;
assign w9210 = w9200 & ~w9209;
assign w9211 = ~w9200 & w9209;
assign v4355 = ~(w9210 | w9211);
assign w9212 = v4355;
assign w9213 = pi07 & pi60;
assign w9214 = pi09 & pi58;
assign v4356 = ~(w8947 | w9214);
assign w9215 = v4356;
assign w9216 = pi09 & pi59;
assign w9217 = w8945 & w9216;
assign v4357 = ~(w9215 | w9217);
assign w9218 = v4357;
assign w9219 = w9213 & ~w9218;
assign w9220 = ~w9213 & w9218;
assign v4358 = ~(w9219 | w9220);
assign w9221 = v4358;
assign w9222 = pi23 & pi44;
assign w9223 = pi24 & pi43;
assign v4359 = ~(w9222 | w9223);
assign w9224 = v4359;
assign w9225 = pi24 & pi44;
assign w9226 = w8841 & w9225;
assign v4360 = ~(w9224 | w9226);
assign w9227 = v4360;
assign w9228 = w8835 & ~w9227;
assign w9229 = ~w8835 & w9227;
assign v4361 = ~(w9228 | w9229);
assign w9230 = v4361;
assign v4362 = ~(w9221 | w9230);
assign w9231 = v4362;
assign w9232 = w9221 & w9230;
assign v4363 = ~(w9231 | w9232);
assign w9233 = v4363;
assign w9234 = pi15 & pi52;
assign w9235 = pi16 & pi51;
assign w9236 = pi30 & pi37;
assign v4364 = ~(w9235 | w9236);
assign w9237 = v4364;
assign w9238 = w9235 & w9236;
assign v4365 = ~(w9237 | w9238);
assign w9239 = v4365;
assign w9240 = w9234 & ~w9239;
assign w9241 = ~w9234 & w9239;
assign v4366 = ~(w9240 | w9241);
assign w9242 = v4366;
assign w9243 = w9233 & ~w9242;
assign w9244 = ~w9233 & w9242;
assign v4367 = ~(w9243 | w9244);
assign w9245 = v4367;
assign w9246 = w9212 & w9245;
assign v4368 = ~(w9212 | w9245);
assign w9247 = v4368;
assign v4369 = ~(w9246 | w9247);
assign w9248 = v4369;
assign w9249 = w9180 & w9248;
assign v4370 = ~(w9180 | w9248);
assign w9250 = v4370;
assign v4371 = ~(w9249 | w9250);
assign w9251 = v4371;
assign w9252 = (w9025 & w17794) | (w9025 & w17795) | (w17794 & w17795);
assign w9253 = (~w9025 & w17796) | (~w9025 & w17797) | (w17796 & w17797);
assign v4372 = ~(w9252 | w9253);
assign w9254 = v4372;
assign w9255 = (~w8967 & ~w8969) | (~w8967 & w17798) | (~w8969 & w17798);
assign w9256 = (~w8979 & ~w8981) | (~w8979 & w17158) | (~w8981 & w17158);
assign w9257 = (~w9005 & ~w9007) | (~w9005 & w17159) | (~w9007 & w17159);
assign v4373 = ~(w9256 | w9257);
assign w9258 = v4373;
assign w9259 = w9256 & w9257;
assign v4374 = ~(w9258 | w9259);
assign w9260 = v4374;
assign w9261 = w9255 & ~w9260;
assign w9262 = ~w9255 & w9260;
assign v4375 = ~(w9261 | w9262);
assign w9263 = v4375;
assign w9264 = (~w8989 & ~w8990) | (~w8989 & w17160) | (~w8990 & w17160);
assign w9265 = (~w9015 & ~w9016) | (~w9015 & w17161) | (~w9016 & w17161);
assign v4376 = ~(w9264 | w9265);
assign w9266 = v4376;
assign w9267 = w9264 & w9265;
assign v4377 = ~(w9266 | w9267);
assign w9268 = v4377;
assign w9269 = w9263 & w9268;
assign v4378 = ~(w9263 | w9268);
assign w9270 = v4378;
assign v4379 = ~(w9269 | w9270);
assign w9271 = v4379;
assign w9272 = w9254 & w9271;
assign v4380 = ~(w9254 | w9271);
assign w9273 = v4380;
assign v4381 = ~(w9272 | w9273);
assign w9274 = v4381;
assign w9275 = (~w9029 & ~w9031) | (~w9029 & w17799) | (~w9031 & w17799);
assign v4382 = ~(w8904 | w8924);
assign w9276 = v4382;
assign v4383 = ~(w9275 | w9276);
assign w9277 = v4383;
assign w9278 = w9275 & w9276;
assign v4384 = ~(w9277 | w9278);
assign w9279 = v4384;
assign v4385 = ~(w9274 | w9279);
assign w9280 = v4385;
assign w9281 = w9274 & w9279;
assign v4386 = ~(w9280 | w9281);
assign w9282 = v4386;
assign w9283 = w9149 & w9282;
assign v4387 = ~(w9149 | w9282);
assign w9284 = v4387;
assign v4388 = ~(w9283 | w9284);
assign w9285 = v4388;
assign w9286 = ~w9047 & w9285;
assign w9287 = w9047 & ~w9285;
assign v4389 = ~(w9286 | w9287);
assign w9288 = v4389;
assign w9289 = (w7754 & w17800) | (w7754 & w17801) | (w17800 & w17801);
assign w9290 = w9288 & w9289;
assign v4390 = ~(w9288 | w9289);
assign w9291 = v4390;
assign v4391 = ~(w9290 | w9291);
assign w9292 = v4391;
assign v4392 = ~(w9106 | w9144);
assign w9293 = v4392;
assign v4393 = ~(w9252 | w9272);
assign w9294 = v4393;
assign v4394 = ~(w9138 | w9141);
assign w9295 = v4394;
assign v4395 = ~(w9130 | w9134);
assign w9296 = v4395;
assign w9297 = (~w9094 & ~w9096) | (~w9094 & w17802) | (~w9096 & w17802);
assign w9298 = (~w9054 & ~w9056) | (~w9054 & w17803) | (~w9056 & w17803);
assign v4396 = ~(w9297 | w9298);
assign w9299 = v4396;
assign w9300 = w9297 & w9298;
assign v4397 = ~(w9299 | w9300);
assign w9301 = v4397;
assign w9302 = w9296 & ~w9301;
assign w9303 = ~w9296 & w9301;
assign v4398 = ~(w9302 | w9303);
assign w9304 = v4398;
assign w9305 = pi10 & pi58;
assign w9306 = pi11 & pi57;
assign v4399 = ~(w9305 | w9306);
assign w9307 = v4399;
assign w9308 = pi11 & pi58;
assign w9309 = w9117 & w9308;
assign v4400 = ~(w9307 | w9309);
assign w9310 = v4400;
assign w9311 = w9216 & ~w9310;
assign w9312 = ~w9216 & w9310;
assign v4401 = ~(w9311 | w9312);
assign w9313 = v4401;
assign w9314 = pi27 & pi41;
assign w9315 = pi28 & pi40;
assign w9316 = pi29 & pi39;
assign v4402 = ~(w9315 | w9316);
assign w9317 = v4402;
assign w9318 = w9315 & w9316;
assign v4403 = ~(w9317 | w9318);
assign w9319 = v4403;
assign w9320 = w9314 & ~w9319;
assign w9321 = ~w9314 & w9319;
assign v4404 = ~(w9320 | w9321);
assign w9322 = v4404;
assign v4405 = ~(w9313 | w9322);
assign w9323 = v4405;
assign w9324 = w9313 & w9322;
assign v4406 = ~(w9323 | w9324);
assign w9325 = v4406;
assign w9326 = pi21 & pi47;
assign w9327 = pi05 & pi63;
assign w9328 = pi06 & pi62;
assign v4407 = ~(w9327 | w9328);
assign w9329 = v4407;
assign w9330 = pi06 & pi63;
assign w9331 = w8802 & w9330;
assign v4408 = ~(w9329 | w9331);
assign w9332 = v4408;
assign w9333 = w9326 & ~w9332;
assign w9334 = ~w9326 & w9332;
assign v4409 = ~(w9333 | w9334);
assign w9335 = v4409;
assign w9336 = w9325 & ~w9335;
assign w9337 = ~w9325 & w9335;
assign v4410 = ~(w9336 | w9337);
assign w9338 = v4410;
assign w9339 = pi18 & pi50;
assign w9340 = pi19 & pi49;
assign v4411 = ~(w9339 | w9340);
assign w9341 = v4411;
assign w9342 = pi19 & pi50;
assign w9343 = w9181 & w9342;
assign v4412 = ~(w9341 | w9343);
assign w9344 = v4412;
assign w9345 = w9192 & ~w9344;
assign w9346 = ~w9192 & w9344;
assign v4413 = ~(w9345 | w9346);
assign w9347 = v4413;
assign w9348 = pi30 & pi38;
assign w9349 = pi32 & pi36;
assign w9350 = pi31 & pi37;
assign v4414 = ~(w9349 | w9350);
assign w9351 = v4414;
assign w9352 = w9349 & w9350;
assign v4415 = ~(w9351 | w9352);
assign w9353 = v4415;
assign w9354 = w9348 & ~w9353;
assign w9355 = ~w9348 & w9353;
assign v4416 = ~(w9354 | w9355);
assign w9356 = v4416;
assign v4417 = ~(w9347 | w9356);
assign w9357 = v4417;
assign w9358 = w9347 & w9356;
assign v4418 = ~(w9357 | w9358);
assign w9359 = v4418;
assign w9360 = pi12 & pi56;
assign w9361 = pi17 & pi51;
assign v4419 = ~(w9204 | w9361);
assign w9362 = v4419;
assign w9363 = w9204 & w9361;
assign v4420 = ~(w9362 | w9363);
assign w9364 = v4420;
assign w9365 = w9360 & ~w9364;
assign w9366 = ~w9360 & w9364;
assign v4421 = ~(w9365 | w9366);
assign w9367 = v4421;
assign w9368 = w9359 & ~w9367;
assign w9369 = ~w9359 & w9367;
assign v4422 = ~(w9368 | w9369);
assign w9370 = v4422;
assign w9371 = pi14 & pi54;
assign w9372 = pi16 & pi52;
assign w9373 = pi15 & pi53;
assign v4423 = ~(w9372 | w9373);
assign w9374 = v4423;
assign w9375 = pi16 & pi53;
assign w9376 = w9234 & w9375;
assign v4424 = ~(w9374 | w9376);
assign w9377 = v4424;
assign w9378 = w9371 & ~w9377;
assign w9379 = ~w9371 & w9377;
assign v4425 = ~(w9378 | w9379);
assign w9380 = v4425;
assign w9381 = pi20 & pi48;
assign w9382 = pi22 & pi46;
assign w9383 = pi23 & pi45;
assign v4426 = ~(w9382 | w9383);
assign w9384 = v4426;
assign w9385 = pi23 & pi46;
assign w9386 = w8835 & w9385;
assign v4427 = ~(w9384 | w9386);
assign w9387 = v4427;
assign w9388 = w9381 & ~w9387;
assign w9389 = ~w9381 & w9387;
assign v4428 = ~(w9388 | w9389);
assign w9390 = v4428;
assign v4429 = ~(w9380 | w9390);
assign w9391 = v4429;
assign w9392 = w9380 & w9390;
assign v4430 = ~(w9391 | w9392);
assign w9393 = v4430;
assign w9394 = pi25 & pi43;
assign w9395 = pi26 & pi42;
assign v4431 = ~(w9394 | w9395);
assign w9396 = v4431;
assign w9397 = pi26 & pi43;
assign w9398 = w9158 & w9397;
assign v4432 = ~(w9396 | w9398);
assign w9399 = v4432;
assign w9400 = w9225 & ~w9399;
assign w9401 = ~w9225 & w9399;
assign v4433 = ~(w9400 | w9401);
assign w9402 = v4433;
assign w9403 = w9393 & ~w9402;
assign w9404 = ~w9393 & w9402;
assign v4434 = ~(w9403 | w9404);
assign w9405 = v4434;
assign w9406 = w9370 & w9405;
assign v4435 = ~(w9370 | w9405);
assign w9407 = v4435;
assign v4436 = ~(w9406 | w9407);
assign w9408 = v4436;
assign w9409 = w9338 & w9408;
assign v4437 = ~(w9338 | w9408);
assign w9410 = v4437;
assign v4438 = ~(w9409 | w9410);
assign w9411 = v4438;
assign w9412 = w9304 & w9411;
assign v4439 = ~(w9304 | w9411);
assign w9413 = v4439;
assign v4440 = ~(w9412 | w9413);
assign w9414 = v4440;
assign w9415 = ~w9295 & w9414;
assign w9416 = w9295 & ~w9414;
assign v4441 = ~(w9415 | w9416);
assign w9417 = v4441;
assign w9418 = ~w9294 & w9417;
assign w9419 = w9294 & ~w9417;
assign v4442 = ~(w9418 | w9419);
assign w9420 = v4442;
assign w9421 = ~w9293 & w9420;
assign w9422 = w9293 & ~w9420;
assign v4443 = ~(w9421 | w9422);
assign w9423 = v4443;
assign v4444 = ~(w9277 | w9281);
assign w9424 = v4444;
assign w9425 = (~w9266 & ~w9268) | (~w9266 & w17599) | (~w9268 & w17599);
assign v4445 = ~(w9158 | w9161);
assign w9426 = v4445;
assign v4446 = ~(w9160 | w9426);
assign w9427 = v4446;
assign v4447 = ~(w9150 | w9153);
assign w9428 = v4447;
assign v4448 = ~(w9152 | w9428);
assign w9429 = v4448;
assign w9430 = w9427 & w9429;
assign v4449 = ~(w9427 | w9429);
assign w9431 = v4449;
assign v4450 = ~(w9430 | w9431);
assign w9432 = v4450;
assign w9433 = w8811 & ~w9203;
assign v4451 = ~(w9205 | w9433);
assign w9434 = v4451;
assign w9435 = ~w9432 & w9434;
assign w9436 = w9432 & ~w9434;
assign v4452 = ~(w9435 | w9436);
assign w9437 = v4452;
assign w9438 = (~w9166 & ~w9168) | (~w9166 & w17600) | (~w9168 & w17600);
assign w9439 = (~w9198 & ~w9200) | (~w9198 & w17601) | (~w9200 & w17601);
assign v4453 = ~(w9438 | w9439);
assign w9440 = v4453;
assign w9441 = w9438 & w9439;
assign v4454 = ~(w9440 | w9441);
assign w9442 = v4454;
assign w9443 = w9437 & w9442;
assign v4455 = ~(w9437 | w9442);
assign w9444 = v4455;
assign v4456 = ~(w9443 | w9444);
assign w9445 = v4456;
assign w9446 = (~w9258 & ~w9260) | (~w9258 & w17602) | (~w9260 & w17602);
assign v4457 = ~(w9117 | w9121);
assign w9447 = v4457;
assign v4458 = ~(w9120 | w9447);
assign w9448 = v4458;
assign w9449 = w8835 & ~w9224;
assign v4459 = ~(w9226 | w9449);
assign w9450 = v4459;
assign w9451 = w9448 & ~w9450;
assign w9452 = ~w9448 & w9450;
assign v4460 = ~(w9451 | w9452);
assign w9453 = v4460;
assign w9454 = w9213 & ~w9215;
assign v4461 = ~(w9217 | w9454);
assign w9455 = v4461;
assign w9456 = ~w9453 & w9455;
assign w9457 = w9453 & ~w9455;
assign v4462 = ~(w9456 | w9457);
assign w9458 = v4462;
assign v4463 = ~(w9169 | w9173);
assign w9459 = v4463;
assign v4464 = ~(w9172 | w9459);
assign w9460 = v4464;
assign w9461 = w9188 & ~w9191;
assign v4465 = ~(w9193 | w9461);
assign w9462 = v4465;
assign w9463 = w9460 & ~w9462;
assign w9464 = ~w9460 & w9462;
assign v4466 = ~(w9463 | w9464);
assign w9465 = v4466;
assign v4467 = ~(w9234 | w9238);
assign w9466 = v4467;
assign v4468 = ~(w9237 | w9466);
assign w9467 = v4468;
assign v4469 = ~(w9465 | w9467);
assign w9468 = v4469;
assign w9469 = w9465 & w9467;
assign v4470 = ~(w9468 | w9469);
assign w9470 = v4470;
assign w9471 = w9458 & w9470;
assign v4471 = ~(w9458 | w9470);
assign w9472 = v4471;
assign v4472 = ~(w9471 | w9472);
assign w9473 = v4472;
assign w9474 = ~w9446 & w9473;
assign w9475 = w9446 & ~w9473;
assign v4473 = ~(w9474 | w9475);
assign w9476 = v4473;
assign w9477 = w9445 & w9476;
assign v4474 = ~(w9445 | w9476);
assign w9478 = v4474;
assign v4475 = ~(w9477 | w9478);
assign w9479 = v4475;
assign w9480 = ~w9425 & w9479;
assign w9481 = w9425 & ~w9479;
assign v4476 = ~(w9480 | w9481);
assign w9482 = v4476;
assign v4477 = ~(w9100 | w9103);
assign w9483 = v4477;
assign v4478 = ~(w9246 | w9249);
assign w9484 = v4478;
assign w9485 = (~w9231 & ~w9233) | (~w9231 & w16922) | (~w9233 & w16922);
assign w9486 = (~w9114 & ~w9116) | (~w9114 & w16761) | (~w9116 & w16761);
assign w9487 = (~w9076 & ~w9078) | (~w9076 & w16762) | (~w9078 & w16762);
assign v4479 = ~(w9486 | w9487);
assign w9488 = v4479;
assign w9489 = w9486 & w9487;
assign v4480 = ~(w9488 | w9489);
assign w9490 = v4480;
assign w9491 = w9485 & ~w9490;
assign w9492 = ~w9485 & w9490;
assign v4481 = ~(w9491 | w9492);
assign w9493 = v4481;
assign w9494 = (~w9064 & ~w9066) | (~w9064 & w17162) | (~w9066 & w17162);
assign w9495 = (~w9086 & ~w9088) | (~w9086 & w16923) | (~w9088 & w16923);
assign w9496 = pi08 & pi60;
assign w9497 = pi07 & pi61;
assign v4482 = ~(w9496 | w9497);
assign w9498 = v4482;
assign w9499 = pi08 & pi61;
assign w9500 = w9213 & w9499;
assign v4483 = ~(w9498 | w9500);
assign w9501 = v4483;
assign w9502 = w9181 & ~w9183;
assign v4484 = ~(w9182 | w9502);
assign w9503 = v4484;
assign w9504 = w9501 & ~w9503;
assign w9505 = ~w9501 & w9503;
assign v4485 = ~(w9504 | w9505);
assign w9506 = v4485;
assign w9507 = ~w9495 & w9506;
assign w9508 = w9495 & ~w9506;
assign v4486 = ~(w9507 | w9508);
assign w9509 = v4486;
assign w9510 = w9494 & ~w9509;
assign w9511 = ~w9494 & w9509;
assign v4487 = ~(w9510 | w9511);
assign w9512 = v4487;
assign w9513 = w9493 & w9512;
assign v4488 = ~(w9493 | w9512);
assign w9514 = v4488;
assign v4489 = ~(w9513 | w9514);
assign w9515 = v4489;
assign w9516 = ~w9484 & w9515;
assign w9517 = w9484 & ~w9515;
assign v4490 = ~(w9516 | w9517);
assign w9518 = v4490;
assign w9519 = ~w9483 & w9518;
assign w9520 = w9483 & ~w9518;
assign v4491 = ~(w9519 | w9520);
assign w9521 = v4491;
assign v4492 = ~(w9482 | w9521);
assign w9522 = v4492;
assign w9523 = w9482 & w9521;
assign v4493 = ~(w9522 | w9523);
assign w9524 = v4493;
assign w9525 = ~w9424 & w9524;
assign w9526 = w9424 & ~w9524;
assign v4494 = ~(w9525 | w9526);
assign w9527 = v4494;
assign w9528 = w9423 & w9527;
assign v4495 = ~(w9423 | w9527);
assign w9529 = v4495;
assign v4496 = ~(w9528 | w9529);
assign w9530 = v4496;
assign v4497 = ~(w9147 | w9283);
assign w9531 = v4497;
assign w9532 = ~w9530 & w9531;
assign w9533 = w9530 & ~w9531;
assign v4498 = ~(w9532 | w9533);
assign w9534 = v4498;
assign v4499 = ~(w9042 | w9287);
assign w9535 = v4499;
assign w9536 = (~w7754 & w17804) | (~w7754 & w17805) | (w17804 & w17805);
assign w9537 = w9534 & w9536;
assign v4500 = ~(w9534 | w9536);
assign w9538 = v4500;
assign v4501 = ~(w9537 | w9538);
assign w9539 = v4501;
assign v4502 = ~(w9525 | w9528);
assign w9540 = v4502;
assign v4503 = ~(w9418 | w9421);
assign w9541 = v4503;
assign v4504 = ~(w9477 | w9480);
assign w9542 = v4504;
assign v4505 = ~(w9406 | w9409);
assign w9543 = v4505;
assign v4506 = ~(w9471 | w9474);
assign w9544 = v4506;
assign v4507 = ~(w9360 | w9363);
assign w9545 = v4507;
assign v4508 = ~(w9362 | w9545);
assign w9546 = v4508;
assign w9547 = w9225 & ~w9396;
assign v4509 = ~(w9398 | w9547);
assign w9548 = v4509;
assign w9549 = w9546 & ~w9548;
assign w9550 = ~w9546 & w9548;
assign v4510 = ~(w9549 | w9550);
assign w9551 = v4510;
assign v4511 = ~(w9314 | w9318);
assign w9552 = v4511;
assign v4512 = ~(w9317 | w9552);
assign w9553 = v4512;
assign v4513 = ~(w9551 | w9553);
assign w9554 = v4513;
assign w9555 = w9551 & w9553;
assign v4514 = ~(w9554 | w9555);
assign w9556 = v4514;
assign w9557 = (~w9463 & ~w9465) | (~w9463 & w16763) | (~w9465 & w16763);
assign w9558 = (~w9430 & ~w9432) | (~w9430 & w16764) | (~w9432 & w16764);
assign v4515 = ~(w9557 | w9558);
assign w9559 = v4515;
assign w9560 = w9557 & w9558;
assign v4516 = ~(w9559 | w9560);
assign w9561 = v4516;
assign w9562 = w9556 & w9561;
assign v4517 = ~(w9556 | w9561);
assign w9563 = v4517;
assign v4518 = ~(w9562 | w9563);
assign w9564 = v4518;
assign w9565 = ~w9544 & w9564;
assign w9566 = w9544 & ~w9564;
assign v4519 = ~(w9565 | w9566);
assign w9567 = v4519;
assign w9568 = ~w9543 & w9567;
assign w9569 = w9543 & ~w9567;
assign v4520 = ~(w9568 | w9569);
assign w9570 = v4520;
assign w9571 = ~w9542 & w9570;
assign w9572 = w9542 & ~w9570;
assign v4521 = ~(w9571 | w9572);
assign w9573 = v4521;
assign v4522 = ~(w9299 | w9303);
assign w9574 = v4522;
assign w9575 = (~w9507 & ~w9509) | (~w9507 & w17163) | (~w9509 & w17163);
assign w9576 = (~w9357 & ~w9359) | (~w9357 & w16924) | (~w9359 & w16924);
assign w9577 = (~w9391 & ~w9393) | (~w9391 & w16925) | (~w9393 & w16925);
assign v4523 = ~(w9576 | w9577);
assign w9578 = v4523;
assign w9579 = w9576 & w9577;
assign v4524 = ~(w9578 | w9579);
assign w9580 = v4524;
assign w9581 = w9575 & ~w9580;
assign w9582 = ~w9575 & w9580;
assign v4525 = ~(w9581 | w9582);
assign w9583 = v4525;
assign w9584 = w9216 & ~w9307;
assign v4526 = ~(w9309 | w9584);
assign w9585 = v4526;
assign w9586 = w9326 & ~w9329;
assign v4527 = ~(w9331 | w9586);
assign w9587 = v4527;
assign v4528 = ~(w9585 | w9587);
assign w9588 = v4528;
assign w9589 = w9585 & w9587;
assign v4529 = ~(w9588 | w9589);
assign w9590 = v4529;
assign w9591 = w9381 & ~w9384;
assign v4530 = ~(w9386 | w9591);
assign w9592 = v4530;
assign w9593 = ~w9590 & w9592;
assign w9594 = w9590 & ~w9592;
assign v4531 = ~(w9593 | w9594);
assign w9595 = v4531;
assign v4532 = ~(w9348 | w9352);
assign w9596 = v4532;
assign v4533 = ~(w9351 | w9596);
assign w9597 = v4533;
assign w9598 = w9192 & ~w9341;
assign v4534 = ~(w9343 | w9598);
assign w9599 = v4534;
assign w9600 = w9597 & ~w9599;
assign w9601 = ~w9597 & w9599;
assign v4535 = ~(w9600 | w9601);
assign w9602 = v4535;
assign w9603 = w9371 & ~w9374;
assign v4536 = ~(w9376 | w9603);
assign w9604 = v4536;
assign w9605 = ~w9602 & w9604;
assign w9606 = w9602 & ~w9604;
assign v4537 = ~(w9605 | w9606);
assign w9607 = v4537;
assign w9608 = (~w9323 & ~w9325) | (~w9323 & w16926) | (~w9325 & w16926);
assign w9609 = ~w9607 & w9608;
assign w9610 = w9607 & ~w9608;
assign v4538 = ~(w9609 | w9610);
assign w9611 = v4538;
assign w9612 = w9595 & w9611;
assign v4539 = ~(w9595 | w9611);
assign w9613 = v4539;
assign v4540 = ~(w9612 | w9613);
assign w9614 = v4540;
assign w9615 = w9583 & w9614;
assign v4541 = ~(w9583 | w9614);
assign w9616 = v4541;
assign v4542 = ~(w9615 | w9616);
assign w9617 = v4542;
assign w9618 = w9574 & ~w9617;
assign w9619 = ~w9574 & w9617;
assign v4543 = ~(w9618 | w9619);
assign w9620 = v4543;
assign w9621 = w9573 & w9620;
assign v4544 = ~(w9573 | w9620);
assign w9622 = v4544;
assign v4545 = ~(w9621 | w9622);
assign w9623 = v4545;
assign w9624 = ~w9541 & w9623;
assign w9625 = w9541 & ~w9623;
assign v4546 = ~(w9624 | w9625);
assign w9626 = v4546;
assign w9627 = (~w9488 & ~w9490) | (~w9488 & w16927) | (~w9490 & w16927);
assign w9628 = pi09 & pi60;
assign w9629 = pi10 & pi59;
assign v4547 = ~(w9628 | w9629);
assign w9630 = v4547;
assign w9631 = pi10 & pi60;
assign w9632 = w9216 & w9631;
assign v4548 = ~(w9630 | w9632);
assign w9633 = v4548;
assign w9634 = w9499 & ~w9633;
assign w9635 = ~w9499 & w9633;
assign v4549 = ~(w9634 | w9635);
assign w9636 = v4549;
assign w9637 = pi24 & pi45;
assign w9638 = pi25 & pi44;
assign v4550 = ~(w9637 | w9638);
assign w9639 = v4550;
assign w9640 = pi25 & pi45;
assign w9641 = w9225 & w9640;
assign v4551 = ~(w9639 | w9641);
assign w9642 = v4551;
assign w9643 = w9385 & ~w9642;
assign w9644 = ~w9385 & w9642;
assign v4552 = ~(w9643 | w9644);
assign w9645 = v4552;
assign v4553 = ~(w9636 | w9645);
assign w9646 = v4553;
assign w9647 = w9636 & w9645;
assign v4554 = ~(w9646 | w9647);
assign w9648 = v4554;
assign w9649 = pi27 & pi42;
assign v4555 = ~(w9397 | w9649);
assign w9650 = v4555;
assign w9651 = pi27 & pi43;
assign w9652 = w9395 & w9651;
assign v4556 = ~(w9650 | w9652);
assign w9653 = v4556;
assign w9654 = w9330 & ~w9653;
assign w9655 = ~w9330 & w9653;
assign v4557 = ~(w9654 | w9655);
assign w9656 = v4557;
assign w9657 = w9648 & ~w9656;
assign w9658 = ~w9648 & w9656;
assign v4558 = ~(w9657 | w9658);
assign w9659 = v4558;
assign w9660 = ~w9627 & w9659;
assign w9661 = w9627 & ~w9659;
assign v4559 = ~(w9660 | w9661);
assign w9662 = v4559;
assign w9663 = (~w9500 & w9503) | (~w9500 & w16765) | (w9503 & w16765);
assign w9664 = pi13 & pi56;
assign w9665 = pi12 & pi57;
assign v4560 = ~(w9664 | w9665);
assign w9666 = v4560;
assign w9667 = pi13 & pi57;
assign w9668 = w9360 & w9667;
assign v4561 = ~(w9666 | w9668);
assign w9669 = v4561;
assign w9670 = w9308 & ~w9669;
assign w9671 = ~w9308 & w9669;
assign v4562 = ~(w9670 | w9671);
assign w9672 = v4562;
assign v4563 = ~(w9663 | w9672);
assign w9673 = v4563;
assign w9674 = w9663 & w9672;
assign v4564 = ~(w9673 | w9674);
assign w9675 = v4564;
assign w9676 = pi14 & pi55;
assign w9677 = pi21 & pi48;
assign w9678 = pi22 & pi47;
assign v4565 = ~(w9677 | w9678);
assign w9679 = v4565;
assign w9680 = pi22 & pi48;
assign w9681 = w9326 & w9680;
assign v4566 = ~(w9679 | w9681);
assign w9682 = v4566;
assign w9683 = w9676 & ~w9682;
assign w9684 = ~w9676 & w9682;
assign v4567 = ~(w9683 | w9684);
assign w9685 = v4567;
assign w9686 = w9675 & ~w9685;
assign w9687 = ~w9675 & w9685;
assign v4568 = ~(w9686 | w9687);
assign w9688 = v4568;
assign w9689 = w9662 & w9688;
assign v4569 = ~(w9662 | w9688);
assign w9690 = v4569;
assign v4570 = ~(w9689 | w9690);
assign w9691 = v4570;
assign v4571 = ~(w9513 | w9516);
assign w9692 = v4571;
assign w9693 = (~w9440 & ~w9442) | (~w9440 & w17806) | (~w9442 & w17806);
assign w9694 = (~w9451 & ~w9453) | (~w9451 & w17164) | (~w9453 & w17164);
assign w9695 = pi18 & pi51;
assign w9696 = pi17 & pi52;
assign v4572 = ~(w9695 | w9696);
assign w9697 = v4572;
assign w9698 = pi18 & pi52;
assign w9699 = w9361 & w9698;
assign v4573 = ~(w9697 | w9699);
assign w9700 = v4573;
assign w9701 = w9342 & ~w9700;
assign w9702 = ~w9342 & w9700;
assign v4574 = ~(w9701 | w9702);
assign w9703 = v4574;
assign w9704 = pi28 & pi41;
assign w9705 = pi29 & pi40;
assign w9706 = pi30 & pi39;
assign v4575 = ~(w9705 | w9706);
assign w9707 = v4575;
assign w9708 = w9705 & w9706;
assign v4576 = ~(w9707 | w9708);
assign w9709 = v4576;
assign w9710 = w9704 & ~w9709;
assign w9711 = ~w9704 & w9709;
assign v4577 = ~(w9710 | w9711);
assign w9712 = v4577;
assign v4578 = ~(w9703 | w9712);
assign w9713 = v4578;
assign w9714 = w9703 & w9712;
assign v4579 = ~(w9713 | w9714);
assign w9715 = v4579;
assign w9716 = w9694 & ~w9715;
assign w9717 = ~w9694 & w9715;
assign v4580 = ~(w9716 | w9717);
assign w9718 = v4580;
assign w9719 = pi07 & pi62;
assign w9720 = ~pi34 & pi35;
assign w9721 = w9719 & ~w9720;
assign w9722 = ~w9719 & w9720;
assign v4581 = ~(w9721 | w9722);
assign w9723 = v4581;
assign w9724 = pi31 & pi38;
assign w9725 = pi32 & pi37;
assign w9726 = pi33 & pi36;
assign v4582 = ~(w9725 | w9726);
assign w9727 = v4582;
assign w9728 = w9725 & w9726;
assign v4583 = ~(w9727 | w9728);
assign w9729 = v4583;
assign w9730 = w9724 & ~w9729;
assign w9731 = ~w9724 & w9729;
assign v4584 = ~(w9730 | w9731);
assign w9732 = v4584;
assign v4585 = ~(w9723 | w9732);
assign w9733 = v4585;
assign w9734 = w9723 & w9732;
assign v4586 = ~(w9733 | w9734);
assign w9735 = v4586;
assign w9736 = pi15 & pi54;
assign w9737 = pi20 & pi49;
assign v4587 = ~(w9375 | w9737);
assign w9738 = v4587;
assign w9739 = w9375 & w9737;
assign v4588 = ~(w9738 | w9739);
assign w9740 = v4588;
assign w9741 = w9736 & ~w9740;
assign w9742 = ~w9736 & w9740;
assign v4589 = ~(w9741 | w9742);
assign w9743 = v4589;
assign w9744 = w9735 & ~w9743;
assign w9745 = ~w9735 & w9743;
assign v4590 = ~(w9744 | w9745);
assign w9746 = v4590;
assign v4591 = ~(w9718 | w9746);
assign w9747 = v4591;
assign w9748 = w9718 & w9746;
assign v4592 = ~(w9747 | w9748);
assign w9749 = v4592;
assign w9750 = w9693 & w9749;
assign v4593 = ~(w9693 | w9749);
assign w9751 = v4593;
assign v4594 = ~(w9750 | w9751);
assign w9752 = v4594;
assign v4595 = ~(w9692 | w9752);
assign w9753 = v4595;
assign w9754 = w9692 & w9752;
assign v4596 = ~(w9753 | w9754);
assign w9755 = v4596;
assign w9756 = w9691 & w9755;
assign v4597 = ~(w9691 | w9755);
assign w9757 = v4597;
assign v4598 = ~(w9756 | w9757);
assign w9758 = v4598;
assign w9759 = (~w9519 & ~w9521) | (~w9519 & w17807) | (~w9521 & w17807);
assign v4599 = ~(w9412 | w9415);
assign w9760 = v4599;
assign v4600 = ~(w9759 | w9760);
assign w9761 = v4600;
assign w9762 = w9759 & w9760;
assign v4601 = ~(w9761 | w9762);
assign w9763 = v4601;
assign w9764 = w9758 & w9763;
assign v4602 = ~(w9758 | w9763);
assign w9765 = v4602;
assign v4603 = ~(w9764 | w9765);
assign w9766 = v4603;
assign w9767 = w9626 & w9766;
assign v4604 = ~(w9626 | w9766);
assign w9768 = v4604;
assign v4605 = ~(w9767 | w9768);
assign w9769 = v4605;
assign w9770 = ~w9540 & w9769;
assign w9771 = w9540 & ~w9769;
assign v4606 = ~(w9770 | w9771);
assign w9772 = v4606;
assign v4607 = ~(w9286 | w9533);
assign w9773 = v4607;
assign w9774 = (w8795 & w16560) | (w8795 & w16561) | (w16560 & w16561);
assign w9775 = w9772 & w9774;
assign v4608 = ~(w9772 | w9774);
assign w9776 = v4608;
assign v4609 = ~(w9775 | w9776);
assign w9777 = v4609;
assign v4610 = ~(w9624 | w9767);
assign w9778 = v4610;
assign w9779 = (~w9571 & ~w9573) | (~w9571 & w17808) | (~w9573 & w17808);
assign v4611 = ~(w9704 | w9708);
assign w9780 = v4611;
assign v4612 = ~(w9707 | w9780);
assign w9781 = v4612;
assign w9782 = w9330 & ~w9650;
assign v4613 = ~(w9652 | w9782);
assign w9783 = v4613;
assign w9784 = w9781 & ~w9783;
assign w9785 = ~w9781 & w9783;
assign v4614 = ~(w9784 | w9785);
assign w9786 = v4614;
assign w9787 = w9385 & ~w9639;
assign v4615 = ~(w9641 | w9787);
assign w9788 = v4615;
assign w9789 = ~w9786 & w9788;
assign w9790 = w9786 & ~w9788;
assign v4616 = ~(w9789 | w9790);
assign w9791 = v4616;
assign w9792 = pi08 & pi62;
assign v4617 = ~(pi34 | w9719);
assign w9793 = v4617;
assign w9794 = pi35 & ~w9793;
assign w9795 = w9792 & w9794;
assign v4618 = ~(w9792 | w9794);
assign w9796 = v4618;
assign v4619 = ~(w9795 | w9796);
assign w9797 = v4619;
assign v4620 = ~(w9724 | w9728);
assign w9798 = v4620;
assign v4621 = ~(w9727 | w9798);
assign w9799 = v4621;
assign w9800 = ~w9797 & w9799;
assign w9801 = w9797 & ~w9799;
assign v4622 = ~(w9800 | w9801);
assign w9802 = v4622;
assign w9803 = ~w9791 & w9802;
assign w9804 = w9791 & ~w9802;
assign v4623 = ~(w9803 | w9804);
assign w9805 = v4623;
assign v4624 = ~(w9713 | w9717);
assign w9806 = v4624;
assign w9807 = ~w9805 & w9806;
assign w9808 = w9805 & ~w9806;
assign v4625 = ~(w9807 | w9808);
assign w9809 = v4625;
assign w9810 = (~w9733 & ~w9735) | (~w9733 & w17452) | (~w9735 & w17452);
assign w9811 = (~w9646 & ~w9648) | (~w9646 & w16928) | (~w9648 & w16928);
assign w9812 = (~w9673 & ~w9675) | (~w9673 & w16929) | (~w9675 & w16929);
assign v4626 = ~(w9811 | w9812);
assign w9813 = v4626;
assign w9814 = w9811 & w9812;
assign v4627 = ~(w9813 | w9814);
assign w9815 = v4627;
assign w9816 = w9810 & ~w9815;
assign w9817 = ~w9810 & w9815;
assign v4628 = ~(w9816 | w9817);
assign w9818 = v4628;
assign v4629 = ~(w9747 | w9750);
assign w9819 = v4629;
assign w9820 = w9818 & w9819;
assign v4630 = ~(w9818 | w9819);
assign w9821 = v4630;
assign v4631 = ~(w9820 | w9821);
assign w9822 = v4631;
assign v4632 = ~(w9809 | w9822);
assign w9823 = v4632;
assign w9824 = w9809 & w9822;
assign v4633 = ~(w9823 | w9824);
assign w9825 = v4633;
assign w9826 = ~w9779 & w9825;
assign w9827 = w9779 & ~w9825;
assign v4634 = ~(w9826 | w9827);
assign w9828 = v4634;
assign w9829 = (~w9565 & ~w9567) | (~w9565 & w17809) | (~w9567 & w17809);
assign w9830 = pi09 & pi61;
assign w9831 = pi11 & pi59;
assign v4635 = ~(w9631 | w9831);
assign w9832 = v4635;
assign w9833 = pi11 & pi60;
assign w9834 = w9629 & w9833;
assign v4636 = ~(w9832 | w9834);
assign w9835 = v4636;
assign w9836 = w9830 & ~w9835;
assign w9837 = ~w9830 & w9835;
assign v4637 = ~(w9836 | w9837);
assign w9838 = v4637;
assign w9839 = pi17 & pi53;
assign w9840 = pi16 & pi54;
assign v4638 = ~(w9839 | w9840);
assign w9841 = v4638;
assign w9842 = pi17 & pi54;
assign w9843 = w9375 & w9842;
assign v4639 = ~(w9841 | w9843);
assign w9844 = v4639;
assign w9845 = w9698 & ~w9844;
assign w9846 = ~w9698 & w9844;
assign v4640 = ~(w9845 | w9846);
assign w9847 = v4640;
assign v4641 = ~(w9838 | w9847);
assign w9848 = v4641;
assign w9849 = w9838 & w9847;
assign v4642 = ~(w9848 | w9849);
assign w9850 = v4642;
assign w9851 = pi12 & pi58;
assign w9852 = pi24 & pi46;
assign v4643 = ~(w9667 | w9852);
assign w9853 = v4643;
assign w9854 = w9667 & w9852;
assign v4644 = ~(w9853 | w9854);
assign w9855 = v4644;
assign w9856 = w9851 & ~w9855;
assign w9857 = ~w9851 & w9855;
assign v4645 = ~(w9856 | w9857);
assign w9858 = v4645;
assign w9859 = w9850 & ~w9858;
assign w9860 = ~w9850 & w9858;
assign v4646 = ~(w9859 | w9860);
assign w9861 = v4646;
assign v4647 = ~(w9736 | w9739);
assign w9862 = v4647;
assign v4648 = ~(w9738 | w9862);
assign w9863 = v4648;
assign w9864 = w9342 & ~w9697;
assign v4649 = ~(w9699 | w9864);
assign w9865 = v4649;
assign w9866 = w9863 & ~w9865;
assign w9867 = ~w9863 & w9865;
assign v4650 = ~(w9866 | w9867);
assign w9868 = v4650;
assign w9869 = pi32 & pi38;
assign w9870 = pi33 & pi37;
assign w9871 = pi34 & pi36;
assign v4651 = ~(w9870 | w9871);
assign w9872 = v4651;
assign w9873 = w9870 & w9871;
assign v4652 = ~(w9872 | w9873);
assign w9874 = v4652;
assign w9875 = w9869 & ~w9874;
assign w9876 = ~w9869 & w9874;
assign v4653 = ~(w9875 | w9876);
assign w9877 = v4653;
assign w9878 = ~w9868 & w9877;
assign w9879 = w9868 & ~w9877;
assign v4654 = ~(w9878 | w9879);
assign w9880 = v4654;
assign w9881 = (~w9559 & ~w9561) | (~w9559 & w16930) | (~w9561 & w16930);
assign w9882 = w9880 & ~w9881;
assign w9883 = ~w9880 & w9881;
assign v4655 = ~(w9882 | w9883);
assign w9884 = v4655;
assign w9885 = w9861 & w9884;
assign v4656 = ~(w9861 | w9884);
assign w9886 = v4656;
assign v4657 = ~(w9885 | w9886);
assign w9887 = v4657;
assign w9888 = ~w9829 & w9887;
assign w9889 = w9829 & ~w9887;
assign v4658 = ~(w9888 | w9889);
assign w9890 = v4658;
assign w9891 = (~w9610 & ~w9611) | (~w9610 & w17165) | (~w9611 & w17165);
assign w9892 = (~w9600 & ~w9602) | (~w9600 & w17166) | (~w9602 & w17166);
assign w9893 = pi28 & pi42;
assign w9894 = pi23 & pi47;
assign w9895 = pi07 & pi63;
assign v4659 = ~(w9894 | w9895);
assign w9896 = v4659;
assign w9897 = w9894 & w9895;
assign v4660 = ~(w9896 | w9897);
assign w9898 = v4660;
assign w9899 = w9893 & ~w9898;
assign w9900 = ~w9893 & w9898;
assign v4661 = ~(w9899 | w9900);
assign w9901 = v4661;
assign w9902 = pi29 & pi41;
assign w9903 = pi30 & pi40;
assign w9904 = pi31 & pi39;
assign v4662 = ~(w9903 | w9904);
assign w9905 = v4662;
assign w9906 = w9903 & w9904;
assign v4663 = ~(w9905 | w9906);
assign w9907 = v4663;
assign w9908 = w9902 & ~w9907;
assign w9909 = ~w9902 & w9907;
assign v4664 = ~(w9908 | w9909);
assign w9910 = v4664;
assign v4665 = ~(w9901 | w9910);
assign w9911 = v4665;
assign w9912 = w9901 & w9910;
assign v4666 = ~(w9911 | w9912);
assign w9913 = v4666;
assign w9914 = w9892 & ~w9913;
assign w9915 = ~w9892 & w9913;
assign v4667 = ~(w9914 | w9915);
assign w9916 = v4667;
assign w9917 = pi14 & pi56;
assign w9918 = pi15 & pi55;
assign v4668 = ~(w9917 | w9918);
assign w9919 = v4668;
assign w9920 = pi15 & pi56;
assign w9921 = w9676 & w9920;
assign v4669 = ~(w9919 | w9921);
assign w9922 = v4669;
assign w9923 = w9680 & ~w9922;
assign w9924 = ~w9680 & w9922;
assign v4670 = ~(w9923 | w9924);
assign w9925 = v4670;
assign w9926 = pi26 & pi44;
assign v4671 = ~(w9651 | w9926);
assign w9927 = v4671;
assign w9928 = pi27 & pi44;
assign w9929 = w9397 & w9928;
assign v4672 = ~(w9927 | w9929);
assign w9930 = v4672;
assign w9931 = w9640 & ~w9930;
assign w9932 = ~w9640 & w9930;
assign v4673 = ~(w9931 | w9932);
assign w9933 = v4673;
assign v4674 = ~(w9925 | w9933);
assign w9934 = v4674;
assign w9935 = w9925 & w9933;
assign v4675 = ~(w9934 | w9935);
assign w9936 = v4675;
assign w9937 = pi21 & pi49;
assign w9938 = pi19 & pi51;
assign w9939 = pi20 & pi50;
assign v4676 = ~(w9938 | w9939);
assign w9940 = v4676;
assign w9941 = pi20 & pi51;
assign w9942 = w9342 & w9941;
assign v4677 = ~(w9940 | w9942);
assign w9943 = v4677;
assign w9944 = w9937 & ~w9943;
assign w9945 = ~w9937 & w9943;
assign v4678 = ~(w9944 | w9945);
assign w9946 = v4678;
assign w9947 = w9936 & ~w9946;
assign w9948 = ~w9936 & w9946;
assign v4679 = ~(w9947 | w9948);
assign w9949 = v4679;
assign v4680 = ~(w9916 | w9949);
assign w9950 = v4680;
assign w9951 = w9916 & w9949;
assign v4681 = ~(w9950 | w9951);
assign w9952 = v4681;
assign w9953 = w9891 & w9952;
assign v4682 = ~(w9891 | w9952);
assign w9954 = v4682;
assign v4683 = ~(w9953 | w9954);
assign w9955 = v4683;
assign w9956 = w9890 & ~w9955;
assign w9957 = ~w9890 & w9955;
assign v4684 = ~(w9956 | w9957);
assign w9958 = v4684;
assign w9959 = w9828 & w9958;
assign v4685 = ~(w9828 | w9958);
assign w9960 = v4685;
assign v4686 = ~(w9959 | w9960);
assign w9961 = v4686;
assign v4687 = ~(w9753 | w9756);
assign w9962 = v4687;
assign v4688 = ~(w9615 | w9619);
assign w9963 = v4688;
assign w9964 = (~w9660 & ~w9662) | (~w9660 & w17167) | (~w9662 & w17167);
assign w9965 = (~w9578 & ~w9580) | (~w9578 & w17168) | (~w9580 & w17168);
assign w9966 = w9499 & ~w9630;
assign v4689 = ~(w9632 | w9966);
assign w9967 = v4689;
assign w9968 = w9308 & ~w9666;
assign v4690 = ~(w9668 | w9968);
assign w9969 = v4690;
assign v4691 = ~(w9967 | w9969);
assign w9970 = v4691;
assign w9971 = w9967 & w9969;
assign v4692 = ~(w9970 | w9971);
assign w9972 = v4692;
assign w9973 = w9676 & ~w9679;
assign v4693 = ~(w9681 | w9973);
assign w9974 = v4693;
assign w9975 = ~w9972 & w9974;
assign w9976 = w9972 & ~w9974;
assign v4694 = ~(w9975 | w9976);
assign w9977 = v4694;
assign w9978 = (~w9588 & ~w9590) | (~w9588 & w16766) | (~w9590 & w16766);
assign w9979 = (~w9549 & ~w9551) | (~w9549 & w16767) | (~w9551 & w16767);
assign v4695 = ~(w9978 | w9979);
assign w9980 = v4695;
assign w9981 = w9978 & w9979;
assign v4696 = ~(w9980 | w9981);
assign w9982 = v4696;
assign w9983 = w9977 & w9982;
assign v4697 = ~(w9977 | w9982);
assign w9984 = v4697;
assign v4698 = ~(w9983 | w9984);
assign w9985 = v4698;
assign w9986 = ~w9965 & w9985;
assign w9987 = w9965 & ~w9985;
assign v4699 = ~(w9986 | w9987);
assign w9988 = v4699;
assign w9989 = ~w9964 & w9988;
assign w9990 = w9964 & ~w9988;
assign v4700 = ~(w9989 | w9990);
assign w9991 = v4700;
assign w9992 = ~w9963 & w9991;
assign w9993 = w9963 & ~w9991;
assign v4701 = ~(w9992 | w9993);
assign w9994 = v4701;
assign w9995 = w9962 & ~w9994;
assign w9996 = ~w9962 & w9994;
assign v4702 = ~(w9995 | w9996);
assign w9997 = v4702;
assign v4703 = ~(w9761 | w9764);
assign w9998 = v4703;
assign w9999 = w9997 & ~w9998;
assign w10000 = ~w9997 & w9998;
assign v4704 = ~(w9999 | w10000);
assign w10001 = v4704;
assign w10002 = w9961 & w10001;
assign v4705 = ~(w9961 | w10001);
assign w10003 = v4705;
assign v4706 = ~(w10002 | w10003);
assign w10004 = v4706;
assign w10005 = ~w9778 & w10004;
assign w10006 = w9778 & ~w10004;
assign v4707 = ~(w10005 | w10006);
assign w10007 = v4707;
assign w10008 = (~w7754 & w17605) | (~w7754 & w17606) | (w17605 & w17606);
assign w10009 = (w7754 & w17810) | (w7754 & w17811) | (w17810 & w17811);
assign w10010 = w10007 & w10009;
assign v4708 = ~(w10007 | w10009);
assign w10011 = v4708;
assign v4709 = ~(w10010 | w10011);
assign w10012 = v4709;
assign v4710 = ~(w9771 | w10006);
assign w10013 = v4710;
assign w10014 = (~w7754 & w17812) | (~w7754 & w17813) | (w17812 & w17813);
assign v4711 = ~(w9999 | w10002);
assign w10015 = v4711;
assign v4712 = ~(w9888 | w9956);
assign w10016 = v4712;
assign w10017 = (~w9784 & ~w9786) | (~w9784 & w17169) | (~w9786 & w17169);
assign w10018 = (~w9866 & ~w9868) | (~w9866 & w16768) | (~w9868 & w16768);
assign v4713 = ~(w9795 | w9799);
assign w10019 = v4713;
assign v4714 = ~(w9796 | w10019);
assign w10020 = v4714;
assign w10021 = ~w10018 & w10020;
assign w10022 = w10018 & ~w10020;
assign v4715 = ~(w10021 | w10022);
assign w10023 = v4715;
assign w10024 = w10017 & ~w10023;
assign w10025 = ~w10017 & w10023;
assign v4716 = ~(w10024 | w10025);
assign w10026 = v4716;
assign w10027 = (~w9804 & ~w9805) | (~w9804 & w17170) | (~w9805 & w17170);
assign w10028 = ~w10026 & w10027;
assign w10029 = w10026 & ~w10027;
assign v4717 = ~(w10028 | w10029);
assign w10030 = v4717;
assign w10031 = (~w9882 & ~w9884) | (~w9882 & w17171) | (~w9884 & w17171);
assign w10032 = ~w10030 & w10031;
assign w10033 = w10030 & ~w10031;
assign v4718 = ~(w10032 | w10033);
assign w10034 = v4718;
assign v4719 = ~(w9820 | w9824);
assign w10035 = v4719;
assign w10036 = ~w10034 & w10035;
assign w10037 = w10034 & ~w10035;
assign v4720 = ~(w10036 | w10037);
assign w10038 = v4720;
assign w10039 = w10016 & ~w10038;
assign w10040 = ~w10016 & w10038;
assign v4721 = ~(w10039 | w10040);
assign w10041 = v4721;
assign v4722 = ~(w9826 | w9959);
assign w10042 = v4722;
assign w10043 = ~w10041 & w10042;
assign w10044 = w10041 & ~w10042;
assign v4723 = ~(w10043 | w10044);
assign w10045 = v4723;
assign v4724 = ~(w9992 | w9996);
assign w10046 = v4724;
assign w10047 = (~w9934 & ~w9936) | (~w9934 & w17455) | (~w9936 & w17455);
assign w10048 = (~w9848 & ~w9850) | (~w9848 & w16931) | (~w9850 & w16931);
assign w10049 = (~w9970 & ~w9972) | (~w9970 & w17172) | (~w9972 & w17172);
assign v4725 = ~(w10048 | w10049);
assign w10050 = v4725;
assign w10051 = w10048 & w10049;
assign v4726 = ~(w10050 | w10051);
assign w10052 = v4726;
assign w10053 = w10047 & ~w10052;
assign w10054 = ~w10047 & w10052;
assign v4727 = ~(w10053 | w10054);
assign w10055 = v4727;
assign v4728 = ~(w9950 | w9953);
assign w10056 = v4728;
assign w10057 = w10055 & w10056;
assign v4729 = ~(w10055 | w10056);
assign w10058 = v4729;
assign v4730 = ~(w10057 | w10058);
assign w10059 = v4730;
assign v4731 = ~(w9911 | w9915);
assign w10060 = v4731;
assign v4732 = ~(w9851 | w9854);
assign w10061 = v4732;
assign v4733 = ~(w9853 | w10061);
assign w10062 = v4733;
assign w10063 = w9830 & ~w9832;
assign v4734 = ~(w9834 | w10063);
assign w10064 = v4734;
assign w10065 = w10062 & ~w10064;
assign w10066 = ~w10062 & w10064;
assign v4735 = ~(w10065 | w10066);
assign w10067 = v4735;
assign w10068 = w9640 & ~w9927;
assign v4736 = ~(w9929 | w10068);
assign w10069 = v4736;
assign w10070 = ~w10067 & w10069;
assign w10071 = w10067 & ~w10069;
assign v4737 = ~(w10070 | w10071);
assign w10072 = v4737;
assign v4738 = ~(w9902 | w9906);
assign w10073 = v4738;
assign v4739 = ~(w9905 | w10073);
assign w10074 = v4739;
assign w10075 = w9680 & ~w9919;
assign v4740 = ~(w9921 | w10075);
assign w10076 = v4740;
assign w10077 = w10074 & ~w10076;
assign w10078 = ~w10074 & w10076;
assign v4741 = ~(w10077 | w10078);
assign w10079 = v4741;
assign v4742 = ~(w9893 | w9897);
assign w10080 = v4742;
assign v4743 = ~(w9896 | w10080);
assign w10081 = v4743;
assign v4744 = ~(w10079 | w10081);
assign w10082 = v4744;
assign w10083 = w10079 & w10081;
assign v4745 = ~(w10082 | w10083);
assign w10084 = v4745;
assign w10085 = w10072 & w10084;
assign v4746 = ~(w10072 | w10084);
assign w10086 = v4746;
assign v4747 = ~(w10085 | w10086);
assign w10087 = v4747;
assign w10088 = ~w10060 & w10087;
assign w10089 = w10060 & ~w10087;
assign v4748 = ~(w10088 | w10089);
assign w10090 = v4748;
assign w10091 = w10059 & w10090;
assign v4749 = ~(w10059 | w10090);
assign w10092 = v4749;
assign v4750 = ~(w10091 | w10092);
assign w10093 = v4750;
assign w10094 = ~w10046 & w10093;
assign w10095 = w10046 & ~w10093;
assign v4751 = ~(w10094 | w10095);
assign w10096 = v4751;
assign v4752 = ~(w9986 | w9989);
assign w10097 = v4752;
assign w10098 = pi22 & pi49;
assign w10099 = pi62 & w4081;
assign w10100 = pi09 & pi62;
assign v4753 = ~(pi36 | w10100);
assign w10101 = v4753;
assign v4754 = ~(w10099 | w10101);
assign w10102 = v4754;
assign w10103 = w10098 & ~w10102;
assign w10104 = ~w10098 & w10102;
assign v4755 = ~(w10103 | w10104);
assign w10105 = v4755;
assign w10106 = pi21 & pi50;
assign w10107 = pi19 & pi52;
assign v4756 = ~(w9941 | w10107);
assign w10108 = v4756;
assign w10109 = pi20 & pi52;
assign w10110 = w9938 & w10109;
assign v4757 = ~(w10108 | w10110);
assign w10111 = v4757;
assign w10112 = w10106 & ~w10111;
assign w10113 = ~w10106 & w10111;
assign v4758 = ~(w10112 | w10113);
assign w10114 = v4758;
assign v4759 = ~(w10105 | w10114);
assign w10115 = v4759;
assign w10116 = w10105 & w10114;
assign v4760 = ~(w10115 | w10116);
assign w10117 = v4760;
assign w10118 = pi33 & pi38;
assign w10119 = pi34 & pi37;
assign w10120 = pi35 & pi36;
assign v4761 = ~(w10119 | w10120);
assign w10121 = v4761;
assign w10122 = w10119 & w10120;
assign v4762 = ~(w10121 | w10122);
assign w10123 = v4762;
assign w10124 = w10118 & ~w10123;
assign w10125 = ~w10118 & w10123;
assign v4763 = ~(w10124 | w10125);
assign w10126 = v4763;
assign w10127 = w10117 & ~w10126;
assign w10128 = ~w10117 & w10126;
assign v4764 = ~(w10127 | w10128);
assign w10129 = v4764;
assign v4765 = ~(w9869 | w9873);
assign w10130 = v4765;
assign v4766 = ~(w9872 | w10130);
assign w10131 = v4766;
assign w10132 = w9698 & ~w9841;
assign v4767 = ~(w9843 | w10132);
assign w10133 = v4767;
assign w10134 = w10131 & ~w10133;
assign w10135 = ~w10131 & w10133;
assign v4768 = ~(w10134 | w10135);
assign w10136 = v4768;
assign w10137 = pi08 & pi63;
assign w10138 = pi10 & pi61;
assign v4769 = ~(w10137 | w10138);
assign w10139 = v4769;
assign w10140 = w10137 & w10138;
assign v4770 = ~(w10139 | w10140);
assign w10141 = v4770;
assign w10142 = w9833 & ~w10141;
assign w10143 = ~w9833 & w10141;
assign v4771 = ~(w10142 | w10143);
assign w10144 = v4771;
assign w10145 = ~w10136 & w10144;
assign w10146 = w10136 & ~w10144;
assign v4772 = ~(w10145 | w10146);
assign w10147 = v4772;
assign w10148 = (~w9980 & ~w9982) | (~w9980 & w16932) | (~w9982 & w16932);
assign w10149 = w10147 & ~w10148;
assign w10150 = ~w10147 & w10148;
assign v4773 = ~(w10149 | w10150);
assign w10151 = v4773;
assign w10152 = w10129 & w10151;
assign v4774 = ~(w10129 | w10151);
assign w10153 = v4774;
assign v4775 = ~(w10152 | w10153);
assign w10154 = v4775;
assign w10155 = ~w10097 & w10154;
assign w10156 = w10097 & ~w10154;
assign v4776 = ~(w10155 | w10156);
assign w10157 = v4776;
assign w10158 = (~w9813 & ~w9815) | (~w9813 & w17173) | (~w9815 & w17173);
assign w10159 = pi28 & pi43;
assign w10160 = pi29 & pi42;
assign v4777 = ~(w10159 | w10160);
assign w10161 = v4777;
assign w10162 = pi29 & pi43;
assign w10163 = w9893 & w10162;
assign v4778 = ~(w10161 | w10163);
assign w10164 = v4778;
assign w10165 = w9928 & ~w10164;
assign w10166 = ~w9928 & w10164;
assign v4779 = ~(w10165 | w10166);
assign w10167 = v4779;
assign w10168 = pi30 & pi41;
assign w10169 = pi31 & pi40;
assign w10170 = pi32 & pi39;
assign v4780 = ~(w10169 | w10170);
assign w10171 = v4780;
assign w10172 = w10169 & w10170;
assign v4781 = ~(w10171 | w10172);
assign w10173 = v4781;
assign w10174 = w10168 & ~w10173;
assign w10175 = ~w10168 & w10173;
assign v4782 = ~(w10174 | w10175);
assign w10176 = v4782;
assign v4783 = ~(w10167 | w10176);
assign w10177 = v4783;
assign w10178 = w10167 & w10176;
assign v4784 = ~(w10177 | w10178);
assign w10179 = v4784;
assign w10180 = pi23 & pi48;
assign w10181 = pi18 & pi53;
assign v4785 = ~(w9842 | w10181);
assign w10182 = v4785;
assign w10183 = pi18 & pi54;
assign w10184 = w9839 & w10183;
assign v4786 = ~(w10182 | w10184);
assign w10185 = v4786;
assign w10186 = w10180 & ~w10185;
assign w10187 = ~w10180 & w10185;
assign v4787 = ~(w10186 | w10187);
assign w10188 = v4787;
assign w10189 = w10179 & ~w10188;
assign w10190 = ~w10179 & w10188;
assign v4788 = ~(w10189 | w10190);
assign w10191 = v4788;
assign w10192 = pi13 & pi58;
assign w10193 = pi12 & pi59;
assign v4789 = ~(w10192 | w10193);
assign w10194 = v4789;
assign w10195 = pi13 & pi59;
assign w10196 = w9851 & w10195;
assign v4790 = ~(w10194 | w10196);
assign w10197 = v4790;
assign w10198 = w9937 & ~w9940;
assign v4791 = ~(w9942 | w10198);
assign w10199 = v4791;
assign w10200 = w10197 & ~w10199;
assign w10201 = ~w10197 & w10199;
assign v4792 = ~(w10200 | w10201);
assign w10202 = v4792;
assign w10203 = pi14 & pi57;
assign w10204 = pi16 & pi55;
assign v4793 = ~(w9920 | w10204);
assign w10205 = v4793;
assign w10206 = pi16 & pi56;
assign w10207 = w9918 & w10206;
assign v4794 = ~(w10205 | w10207);
assign w10208 = v4794;
assign w10209 = w10203 & ~w10208;
assign w10210 = ~w10203 & w10208;
assign v4795 = ~(w10209 | w10210);
assign w10211 = v4795;
assign w10212 = pi24 & pi47;
assign w10213 = pi25 & pi46;
assign w10214 = pi26 & pi45;
assign v4796 = ~(w10213 | w10214);
assign w10215 = v4796;
assign w10216 = pi26 & pi46;
assign w10217 = w9640 & w10216;
assign v4797 = ~(w10215 | w10217);
assign w10218 = v4797;
assign w10219 = w10212 & ~w10218;
assign w10220 = ~w10212 & w10218;
assign v4798 = ~(w10219 | w10220);
assign w10221 = v4798;
assign v4799 = ~(w10211 | w10221);
assign w10222 = v4799;
assign w10223 = w10211 & w10221;
assign v4800 = ~(w10222 | w10223);
assign w10224 = v4800;
assign w10225 = w10202 & w10224;
assign v4801 = ~(w10202 | w10224);
assign w10226 = v4801;
assign v4802 = ~(w10225 | w10226);
assign w10227 = v4802;
assign w10228 = w10191 & w10227;
assign v4803 = ~(w10191 | w10227);
assign w10229 = v4803;
assign v4804 = ~(w10228 | w10229);
assign w10230 = v4804;
assign w10231 = ~w10158 & w10230;
assign w10232 = w10158 & ~w10230;
assign v4805 = ~(w10231 | w10232);
assign w10233 = v4805;
assign w10234 = w10157 & w10233;
assign v4806 = ~(w10157 | w10233);
assign w10235 = v4806;
assign v4807 = ~(w10234 | w10235);
assign w10236 = v4807;
assign w10237 = w10096 & w10236;
assign v4808 = ~(w10096 | w10236);
assign w10238 = v4808;
assign v4809 = ~(w10237 | w10238);
assign w10239 = v4809;
assign v4810 = ~(w10045 | w10239);
assign w10240 = v4810;
assign w10241 = w10045 & w10239;
assign v4811 = ~(w10240 | w10241);
assign w10242 = v4811;
assign w10243 = w10015 & ~w10242;
assign w10244 = ~w10015 & w10242;
assign v4812 = ~(w10243 | w10244);
assign w10245 = v4812;
assign w10246 = w10014 & w10245;
assign v4813 = ~(w10014 | w10245);
assign w10247 = v4813;
assign v4814 = ~(w10246 | w10247);
assign w10248 = v4814;
assign v4815 = ~(w10005 | w10244);
assign w10249 = v4815;
assign w10250 = (w7754 & w17814) | (w7754 & w17815) | (w17814 & w17815);
assign w10251 = (~w10155 & ~w10157) | (~w10155 & w17456) | (~w10157 & w17456);
assign w10252 = (~w10085 & ~w10087) | (~w10085 & w17174) | (~w10087 & w17174);
assign w10253 = (~w10077 & ~w10079) | (~w10077 & w17175) | (~w10079 & w17175);
assign w10254 = (~w10134 & ~w10136) | (~w10134 & w16769) | (~w10136 & w16769);
assign w10255 = pi31 & pi41;
assign w10256 = pi30 & pi42;
assign v4816 = ~(w10255 | w10256);
assign w10257 = v4816;
assign w10258 = pi31 & pi42;
assign w10259 = w10168 & w10258;
assign v4817 = ~(w10257 | w10259);
assign w10260 = v4817;
assign w10261 = w10162 & ~w10260;
assign w10262 = ~w10162 & w10260;
assign v4818 = ~(w10261 | w10262);
assign w10263 = v4818;
assign v4819 = ~(w10254 | w10263);
assign w10264 = v4819;
assign w10265 = w10254 & w10263;
assign v4820 = ~(w10264 | w10265);
assign w10266 = v4820;
assign w10267 = w10253 & ~w10266;
assign w10268 = ~w10253 & w10266;
assign v4821 = ~(w10267 | w10268);
assign w10269 = v4821;
assign w10270 = ~w10252 & w10269;
assign w10271 = w10252 & ~w10269;
assign v4822 = ~(w10270 | w10271);
assign w10272 = v4822;
assign w10273 = (~w10149 & ~w10151) | (~w10149 & w17176) | (~w10151 & w17176);
assign w10274 = ~w10272 & w10273;
assign w10275 = w10272 & ~w10273;
assign v4823 = ~(w10274 | w10275);
assign w10276 = v4823;
assign w10277 = (~w10057 & ~w10059) | (~w10057 & w17457) | (~w10059 & w17457);
assign w10278 = ~w10276 & w10277;
assign w10279 = w10276 & ~w10277;
assign v4824 = ~(w10278 | w10279);
assign w10280 = v4824;
assign w10281 = w10251 & ~w10280;
assign w10282 = ~w10251 & w10280;
assign v4825 = ~(w10281 | w10282);
assign w10283 = v4825;
assign v4826 = ~(w10094 | w10237);
assign w10284 = v4826;
assign w10285 = ~w10283 & w10284;
assign w10286 = w10283 & ~w10284;
assign v4827 = ~(w10285 | w10286);
assign w10287 = v4827;
assign v4828 = ~(w10037 | w10040);
assign w10288 = v4828;
assign w10289 = (~w10115 & ~w10117) | (~w10115 & w17458) | (~w10117 & w17458);
assign w10290 = (~w10177 & ~w10179) | (~w10177 & w16933) | (~w10179 & w16933);
assign w10291 = (~w10065 & ~w10067) | (~w10065 & w17177) | (~w10067 & w17177);
assign v4829 = ~(w10290 | w10291);
assign w10292 = v4829;
assign w10293 = w10290 & w10291;
assign v4830 = ~(w10292 | w10293);
assign w10294 = v4830;
assign w10295 = w10289 & ~w10294;
assign w10296 = ~w10289 & w10294;
assign v4831 = ~(w10295 | w10296);
assign w10297 = v4831;
assign v4832 = ~(w10228 | w10231);
assign w10298 = v4832;
assign w10299 = ~w10297 & w10298;
assign w10300 = w10297 & ~w10298;
assign v4833 = ~(w10299 | w10300);
assign w10301 = v4833;
assign w10302 = (~w10222 & ~w10224) | (~w10222 & w17459) | (~w10224 & w17459);
assign w10303 = w9928 & ~w10161;
assign v4834 = ~(w10163 | w10303);
assign w10304 = v4834;
assign w10305 = w10180 & ~w10182;
assign v4835 = ~(w10184 | w10305);
assign w10306 = v4835;
assign v4836 = ~(w10304 | w10306);
assign w10307 = v4836;
assign w10308 = w10304 & w10306;
assign v4837 = ~(w10307 | w10308);
assign w10309 = v4837;
assign v4838 = ~(w10168 | w10172);
assign w10310 = v4838;
assign v4839 = ~(w10171 | w10310);
assign w10311 = v4839;
assign v4840 = ~(w10309 | w10311);
assign w10312 = v4840;
assign w10313 = w10309 & w10311;
assign v4841 = ~(w10312 | w10313);
assign w10314 = v4841;
assign w10315 = w10098 & ~w10101;
assign v4842 = ~(w10099 | w10315);
assign w10316 = v4842;
assign v4843 = ~(w10118 | w10122);
assign w10317 = v4843;
assign v4844 = ~(w10121 | w10317);
assign w10318 = v4844;
assign w10319 = ~w10316 & w10318;
assign w10320 = w10316 & ~w10318;
assign v4845 = ~(w10319 | w10320);
assign w10321 = v4845;
assign w10322 = w10106 & ~w10108;
assign v4846 = ~(w10110 | w10322);
assign w10323 = v4846;
assign w10324 = ~w10321 & w10323;
assign w10325 = w10321 & ~w10323;
assign v4847 = ~(w10324 | w10325);
assign w10326 = v4847;
assign w10327 = w10314 & w10326;
assign v4848 = ~(w10314 | w10326);
assign w10328 = v4848;
assign v4849 = ~(w10327 | w10328);
assign w10329 = v4849;
assign w10330 = ~w10302 & w10329;
assign w10331 = w10302 & ~w10329;
assign v4850 = ~(w10330 | w10331);
assign w10332 = v4850;
assign w10333 = w10301 & w10332;
assign v4851 = ~(w10301 | w10332);
assign w10334 = v4851;
assign v4852 = ~(w10333 | w10334);
assign w10335 = v4852;
assign w10336 = ~w10288 & w10335;
assign w10337 = w10288 & ~w10335;
assign v4853 = ~(w10336 | w10337);
assign w10338 = v4853;
assign w10339 = (~w10050 & ~w10052) | (~w10050 & w17178) | (~w10052 & w17178);
assign w10340 = (~w10196 & w10199) | (~w10196 & w17179) | (w10199 & w17179);
assign w10341 = pi12 & pi60;
assign w10342 = pi25 & pi47;
assign w10343 = pi24 & pi48;
assign v4854 = ~(w10342 | w10343);
assign w10344 = v4854;
assign w10345 = pi25 & pi48;
assign w10346 = w10212 & w10345;
assign v4855 = ~(w10344 | w10346);
assign w10347 = v4855;
assign w10348 = w10341 & ~w10347;
assign w10349 = ~w10341 & w10347;
assign v4856 = ~(w10348 | w10349);
assign w10350 = v4856;
assign v4857 = ~(w10340 | w10350);
assign w10351 = v4857;
assign w10352 = w10340 & w10350;
assign v4858 = ~(w10351 | w10352);
assign w10353 = v4858;
assign w10354 = pi09 & pi63;
assign w10355 = pi10 & pi62;
assign w10356 = pi11 & pi61;
assign v4859 = ~(w10355 | w10356);
assign w10357 = v4859;
assign w10358 = pi11 & pi62;
assign w10359 = w10138 & w10358;
assign v4860 = ~(w10357 | w10359);
assign w10360 = v4860;
assign w10361 = w10354 & ~w10360;
assign w10362 = ~w10354 & w10360;
assign v4861 = ~(w10361 | w10362);
assign w10363 = v4861;
assign w10364 = w10353 & ~w10363;
assign w10365 = ~w10353 & w10363;
assign v4862 = ~(w10364 | w10365);
assign w10366 = v4862;
assign w10367 = pi35 & pi37;
assign w10368 = pi21 & pi51;
assign w10369 = pi22 & pi50;
assign v4863 = ~(w10368 | w10369);
assign w10370 = v4863;
assign w10371 = pi22 & pi51;
assign w10372 = w10106 & w10371;
assign v4864 = ~(w10370 | w10372);
assign w10373 = v4864;
assign w10374 = w10367 & ~w10373;
assign w10375 = ~w10367 & w10373;
assign v4865 = ~(w10374 | w10375);
assign w10376 = v4865;
assign w10377 = pi32 & pi40;
assign w10378 = pi23 & pi49;
assign v4866 = ~(w10206 | w10378);
assign w10379 = v4866;
assign w10380 = w10206 & w10378;
assign v4867 = ~(w10379 | w10380);
assign w10381 = v4867;
assign w10382 = w10377 & ~w10381;
assign w10383 = ~w10377 & w10381;
assign v4868 = ~(w10382 | w10383);
assign w10384 = v4868;
assign v4869 = ~(w10376 | w10384);
assign w10385 = v4869;
assign w10386 = w10376 & w10384;
assign v4870 = ~(w10385 | w10386);
assign w10387 = v4870;
assign w10388 = pi17 & pi55;
assign v4871 = ~(w10109 | w10183);
assign w10389 = v4871;
assign w10390 = w10109 & w10183;
assign v4872 = ~(w10389 | w10390);
assign w10391 = v4872;
assign w10392 = w10388 & ~w10391;
assign w10393 = ~w10388 & w10391;
assign v4873 = ~(w10392 | w10393);
assign w10394 = v4873;
assign w10395 = w10387 & ~w10394;
assign w10396 = ~w10387 & w10394;
assign v4874 = ~(w10395 | w10396);
assign w10397 = v4874;
assign w10398 = w10366 & w10397;
assign v4875 = ~(w10366 | w10397);
assign w10399 = v4875;
assign v4876 = ~(w10398 | w10399);
assign w10400 = v4876;
assign w10401 = ~w10339 & w10400;
assign w10402 = w10339 & ~w10400;
assign v4877 = ~(w10401 | w10402);
assign w10403 = v4877;
assign v4878 = ~(w10029 | w10033);
assign w10404 = v4878;
assign w10405 = w10203 & ~w10205;
assign v4879 = ~(w10207 | w10405);
assign w10406 = v4879;
assign w10407 = w10212 & ~w10215;
assign v4880 = ~(w10217 | w10407);
assign w10408 = v4880;
assign v4881 = ~(w10406 | w10408);
assign w10409 = v4881;
assign w10410 = w10406 & w10408;
assign v4882 = ~(w10409 | w10410);
assign w10411 = v4882;
assign v4883 = ~(w9833 | w10140);
assign w10412 = v4883;
assign v4884 = ~(w10139 | w10412);
assign w10413 = v4884;
assign v4885 = ~(w10411 | w10413);
assign w10414 = v4885;
assign w10415 = w10411 & w10413;
assign v4886 = ~(w10414 | w10415);
assign w10416 = v4886;
assign w10417 = (~w10021 & ~w10023) | (~w10021 & w16934) | (~w10023 & w16934);
assign w10418 = ~w10416 & w10417;
assign w10419 = w10416 & ~w10417;
assign v4887 = ~(w10418 | w10419);
assign w10420 = v4887;
assign w10421 = pi14 & pi58;
assign w10422 = pi15 & pi57;
assign v4888 = ~(w10421 | w10422);
assign w10423 = v4888;
assign w10424 = pi15 & pi58;
assign w10425 = w10203 & w10424;
assign v4889 = ~(w10423 | w10425);
assign w10426 = v4889;
assign w10427 = w10195 & ~w10426;
assign w10428 = ~w10195 & w10426;
assign v4890 = ~(w10427 | w10428);
assign w10429 = v4890;
assign w10430 = pi27 & pi45;
assign w10431 = pi28 & pi44;
assign v4891 = ~(w10430 | w10431);
assign w10432 = v4891;
assign w10433 = pi28 & pi45;
assign w10434 = w9928 & w10433;
assign v4892 = ~(w10432 | w10434);
assign w10435 = v4892;
assign w10436 = w10216 & ~w10435;
assign w10437 = ~w10216 & w10435;
assign v4893 = ~(w10436 | w10437);
assign w10438 = v4893;
assign v4894 = ~(w10429 | w10438);
assign w10439 = v4894;
assign w10440 = w10429 & w10438;
assign v4895 = ~(w10439 | w10440);
assign w10441 = v4895;
assign w10442 = pi19 & pi53;
assign w10443 = pi34 & pi38;
assign w10444 = pi33 & pi39;
assign v4896 = ~(w10443 | w10444);
assign w10445 = v4896;
assign w10446 = pi34 & pi39;
assign w10447 = w10118 & w10446;
assign v4897 = ~(w10445 | w10447);
assign w10448 = v4897;
assign w10449 = w10442 & ~w10448;
assign w10450 = ~w10442 & w10448;
assign v4898 = ~(w10449 | w10450);
assign w10451 = v4898;
assign w10452 = w10441 & ~w10451;
assign w10453 = ~w10441 & w10451;
assign v4899 = ~(w10452 | w10453);
assign w10454 = v4899;
assign v4900 = ~(w10420 | w10454);
assign w10455 = v4900;
assign w10456 = w10420 & w10454;
assign v4901 = ~(w10455 | w10456);
assign w10457 = v4901;
assign w10458 = ~w10404 & w10457;
assign w10459 = w10404 & ~w10457;
assign v4902 = ~(w10458 | w10459);
assign w10460 = v4902;
assign v4903 = ~(w10403 | w10460);
assign w10461 = v4903;
assign w10462 = w10403 & w10460;
assign v4904 = ~(w10461 | w10462);
assign w10463 = v4904;
assign v4905 = ~(w10338 | w10463);
assign w10464 = v4905;
assign w10465 = w10338 & w10463;
assign v4906 = ~(w10464 | w10465);
assign w10466 = v4906;
assign v4907 = ~(w10287 | w10466);
assign w10467 = v4907;
assign w10468 = w10287 & w10466;
assign v4908 = ~(w10467 | w10468);
assign w10469 = v4908;
assign v4909 = ~(w10044 | w10241);
assign w10470 = v4909;
assign w10471 = ~w10469 & w10470;
assign w10472 = w10469 & ~w10470;
assign v4910 = ~(w10471 | w10472);
assign w10473 = v4910;
assign w10474 = w10250 & ~w10473;
assign w10475 = ~w10250 & w10473;
assign v4911 = ~(w10474 | w10475);
assign w10476 = v4911;
assign v4912 = ~(w10286 | w10468);
assign w10477 = v4912;
assign v4913 = ~(w10336 | w10465);
assign w10478 = v4913;
assign w10479 = (~w10458 & ~w10460) | (~w10458 & w17460) | (~w10460 & w17460);
assign w10480 = (~w10300 & ~w10301) | (~w10300 & w17461) | (~w10301 & w17461);
assign w10481 = (~w10419 & ~w10420) | (~w10419 & w17180) | (~w10420 & w17180);
assign v4914 = ~(w10307 | w10313);
assign w10482 = v4914;
assign w10483 = (~w10409 & ~w10411) | (~w10409 & w17181) | (~w10411 & w17181);
assign w10484 = pi33 & pi40;
assign w10485 = pi32 & pi41;
assign v4915 = ~(w10484 | w10485);
assign w10486 = v4915;
assign w10487 = pi33 & pi41;
assign w10488 = w10377 & w10487;
assign v4916 = ~(w10486 | w10488);
assign w10489 = v4916;
assign w10490 = w10258 & ~w10489;
assign w10491 = ~w10258 & w10489;
assign v4917 = ~(w10490 | w10491);
assign w10492 = v4917;
assign v4918 = ~(w10483 | w10492);
assign w10493 = v4918;
assign w10494 = w10483 & w10492;
assign v4919 = ~(w10493 | w10494);
assign w10495 = v4919;
assign w10496 = w10482 & ~w10495;
assign w10497 = ~w10482 & w10495;
assign v4920 = ~(w10496 | w10497);
assign w10498 = v4920;
assign w10499 = (~w10327 & ~w10329) | (~w10327 & w17182) | (~w10329 & w17182);
assign w10500 = ~w10498 & w10499;
assign w10501 = w10498 & ~w10499;
assign v4921 = ~(w10500 | w10501);
assign w10502 = v4921;
assign w10503 = ~w10481 & w10502;
assign w10504 = w10481 & ~w10502;
assign v4922 = ~(w10503 | w10504);
assign w10505 = v4922;
assign w10506 = ~w10480 & w10505;
assign w10507 = w10480 & ~w10505;
assign v4923 = ~(w10506 | w10507);
assign w10508 = v4923;
assign w10509 = ~w10479 & w10508;
assign w10510 = w10479 & ~w10508;
assign v4924 = ~(w10509 | w10510);
assign w10511 = v4924;
assign w10512 = ~w10478 & w10511;
assign w10513 = w10478 & ~w10511;
assign v4925 = ~(w10512 | w10513);
assign w10514 = v4925;
assign w10515 = (~w10439 & ~w10441) | (~w10439 & w17816) | (~w10441 & w17816);
assign w10516 = (~w10351 & ~w10353) | (~w10351 & w17462) | (~w10353 & w17462);
assign w10517 = (~w10319 & ~w10321) | (~w10319 & w17609) | (~w10321 & w17609);
assign v4926 = ~(w10516 | w10517);
assign w10518 = v4926;
assign w10519 = w10516 & w10517;
assign v4927 = ~(w10518 | w10519);
assign w10520 = v4927;
assign w10521 = w10515 & ~w10520;
assign w10522 = ~w10515 & w10520;
assign v4928 = ~(w10521 | w10522);
assign w10523 = v4928;
assign v4929 = ~(w10398 | w10401);
assign w10524 = v4929;
assign w10525 = ~w10523 & w10524;
assign w10526 = w10523 & ~w10524;
assign v4930 = ~(w10525 | w10526);
assign w10527 = v4930;
assign w10528 = (~w10385 & ~w10387) | (~w10385 & w17817) | (~w10387 & w17817);
assign w10529 = pi13 & pi60;
assign w10530 = w10367 & ~w10370;
assign w10531 = (w10529 & w10530) | (w10529 & w17463) | (w10530 & w17463);
assign w10532 = ~w10530 & w17464;
assign v4931 = ~(w10531 | w10532);
assign w10533 = v4931;
assign w10534 = w10442 & ~w10445;
assign v4932 = ~(w10447 | w10534);
assign w10535 = v4932;
assign w10536 = ~w10533 & w10535;
assign w10537 = w10533 & ~w10535;
assign v4933 = ~(w10536 | w10537);
assign w10538 = v4933;
assign w10539 = w10354 & ~w10357;
assign v4934 = ~(w10359 | w10539);
assign w10540 = v4934;
assign w10541 = w10341 & ~w10344;
assign v4935 = ~(w10346 | w10541);
assign w10542 = v4935;
assign v4936 = ~(w10540 | w10542);
assign w10543 = v4936;
assign w10544 = w10540 & w10542;
assign v4937 = ~(w10543 | w10544);
assign w10545 = v4937;
assign v4938 = ~(w10388 | w10390);
assign w10546 = v4938;
assign v4939 = ~(w10389 | w10546);
assign w10547 = v4939;
assign v4940 = ~(w10545 | w10547);
assign w10548 = v4940;
assign w10549 = w10545 & w10547;
assign v4941 = ~(w10548 | w10549);
assign w10550 = v4941;
assign w10551 = w10538 & w10550;
assign v4942 = ~(w10538 | w10550);
assign w10552 = v4942;
assign v4943 = ~(w10551 | w10552);
assign w10553 = v4943;
assign w10554 = ~w10528 & w10553;
assign w10555 = w10528 & ~w10553;
assign v4944 = ~(w10554 | w10555);
assign w10556 = v4944;
assign w10557 = w10527 & w10556;
assign v4945 = ~(w10527 | w10556);
assign w10558 = v4945;
assign v4946 = ~(w10557 | w10558);
assign w10559 = v4946;
assign w10560 = (w10559 & w10282) | (w10559 & w17610) | (w10282 & w17610);
assign w10561 = ~w10282 & w17611;
assign v4947 = ~(w10560 | w10561);
assign w10562 = v4947;
assign w10563 = (~w10292 & ~w10294) | (~w10292 & w17183) | (~w10294 & w17183);
assign v4948 = ~(w10377 | w10380);
assign w10564 = v4948;
assign v4949 = ~(w10379 | w10564);
assign w10565 = v4949;
assign w10566 = pi17 & pi56;
assign w10567 = pi26 & pi47;
assign w10568 = pi27 & pi46;
assign v4950 = ~(w10567 | w10568);
assign w10569 = v4950;
assign w10570 = pi27 & pi47;
assign w10571 = w10216 & w10570;
assign v4951 = ~(w10569 | w10571);
assign w10572 = v4951;
assign w10573 = w10566 & ~w10572;
assign w10574 = ~w10566 & w10572;
assign v4952 = ~(w10573 | w10574);
assign w10575 = v4952;
assign w10576 = w10565 & ~w10575;
assign w10577 = ~w10565 & w10575;
assign v4953 = ~(w10576 | w10577);
assign w10578 = v4953;
assign w10579 = pi14 & pi59;
assign w10580 = pi16 & pi57;
assign v4954 = ~(w10424 | w10580);
assign w10581 = v4954;
assign w10582 = pi16 & pi58;
assign w10583 = w10422 & w10582;
assign v4955 = ~(w10581 | w10583);
assign w10584 = v4955;
assign w10585 = w10579 & ~w10584;
assign w10586 = ~w10579 & w10584;
assign v4956 = ~(w10585 | w10586);
assign w10587 = v4956;
assign w10588 = w10578 & ~w10587;
assign w10589 = ~w10578 & w10587;
assign v4957 = ~(w10588 | w10589);
assign w10590 = v4957;
assign w10591 = pi23 & pi50;
assign w10592 = pi62 & w4629;
assign v4958 = ~(pi37 | w10358);
assign w10593 = v4958;
assign v4959 = ~(w10592 | w10593);
assign w10594 = v4959;
assign w10595 = w10591 & ~w10594;
assign w10596 = ~w10591 & w10594;
assign v4960 = ~(w10595 | w10596);
assign w10597 = v4960;
assign w10598 = pi18 & pi55;
assign w10599 = pi24 & pi49;
assign w10600 = pi19 & pi54;
assign v4961 = ~(w10599 | w10600);
assign w10601 = v4961;
assign w10602 = w10599 & w10600;
assign v4962 = ~(w10601 | w10602);
assign w10603 = v4962;
assign w10604 = w10598 & ~w10603;
assign w10605 = ~w10598 & w10603;
assign v4963 = ~(w10604 | w10605);
assign w10606 = v4963;
assign v4964 = ~(w10597 | w10606);
assign w10607 = v4964;
assign w10608 = w10597 & w10606;
assign v4965 = ~(w10607 | w10608);
assign w10609 = v4965;
assign w10610 = pi20 & pi53;
assign w10611 = pi21 & pi52;
assign v4966 = ~(w10610 | w10611);
assign w10612 = v4966;
assign w10613 = pi21 & pi53;
assign w10614 = w10109 & w10613;
assign v4967 = ~(w10612 | w10614);
assign w10615 = v4967;
assign w10616 = w10371 & ~w10615;
assign w10617 = ~w10371 & w10615;
assign v4968 = ~(w10616 | w10617);
assign w10618 = v4968;
assign w10619 = w10609 & ~w10618;
assign w10620 = ~w10609 & w10618;
assign v4969 = ~(w10619 | w10620);
assign w10621 = v4969;
assign w10622 = w10590 & w10621;
assign v4970 = ~(w10590 | w10621);
assign w10623 = v4970;
assign v4971 = ~(w10622 | w10623);
assign w10624 = v4971;
assign w10625 = w10563 & ~w10624;
assign w10626 = ~w10563 & w10624;
assign v4972 = ~(w10625 | w10626);
assign w10627 = v4972;
assign v4973 = ~(w10270 | w10275);
assign w10628 = v4973;
assign w10629 = w10195 & ~w10423;
assign v4974 = ~(w10425 | w10629);
assign w10630 = v4974;
assign w10631 = w10216 & ~w10432;
assign v4975 = ~(w10434 | w10631);
assign w10632 = v4975;
assign v4976 = ~(w10630 | w10632);
assign w10633 = v4976;
assign w10634 = w10630 & w10632;
assign v4977 = ~(w10633 | w10634);
assign w10635 = v4977;
assign w10636 = w10162 & ~w10257;
assign v4978 = ~(w10259 | w10636);
assign w10637 = v4978;
assign w10638 = ~w10635 & w10637;
assign w10639 = w10635 & ~w10637;
assign v4979 = ~(w10638 | w10639);
assign w10640 = v4979;
assign w10641 = (~w10264 & ~w10266) | (~w10264 & w16935) | (~w10266 & w16935);
assign w10642 = ~w10640 & w10641;
assign w10643 = w10640 & ~w10641;
assign v4980 = ~(w10642 | w10643);
assign w10644 = v4980;
assign w10645 = pi29 & pi44;
assign w10646 = pi30 & pi43;
assign v4981 = ~(w10645 | w10646);
assign w10647 = v4981;
assign w10648 = pi30 & pi44;
assign w10649 = w10162 & w10648;
assign v4982 = ~(w10647 | w10649);
assign w10650 = v4982;
assign w10651 = w10433 & ~w10650;
assign w10652 = ~w10433 & w10650;
assign v4983 = ~(w10651 | w10652);
assign w10653 = v4983;
assign w10654 = pi10 & pi63;
assign w10655 = pi12 & pi61;
assign v4984 = ~(w10654 | w10655);
assign w10656 = v4984;
assign w10657 = w10654 & w10655;
assign v4985 = ~(w10656 | w10657);
assign w10658 = v4985;
assign w10659 = w10345 & ~w10658;
assign w10660 = ~w10345 & w10658;
assign v4986 = ~(w10659 | w10660);
assign w10661 = v4986;
assign v4987 = ~(w10653 | w10661);
assign w10662 = v4987;
assign w10663 = w10653 & w10661;
assign v4988 = ~(w10662 | w10663);
assign w10664 = v4988;
assign w10665 = pi36 & pi37;
assign w10666 = pi35 & pi38;
assign v4989 = ~(w10665 | w10666);
assign w10667 = v4989;
assign w10668 = pi36 & pi38;
assign w10669 = w10367 & w10668;
assign v4990 = ~(w10667 | w10669);
assign w10670 = v4990;
assign w10671 = w10446 & ~w10670;
assign w10672 = ~w10446 & w10670;
assign v4991 = ~(w10671 | w10672);
assign w10673 = v4991;
assign w10674 = w10664 & ~w10673;
assign w10675 = ~w10664 & w10673;
assign v4992 = ~(w10674 | w10675);
assign w10676 = v4992;
assign v4993 = ~(w10644 | w10676);
assign w10677 = v4993;
assign w10678 = w10644 & w10676;
assign v4994 = ~(w10677 | w10678);
assign w10679 = v4994;
assign w10680 = ~w10628 & w10679;
assign w10681 = w10628 & ~w10679;
assign v4995 = ~(w10680 | w10681);
assign w10682 = v4995;
assign v4996 = ~(w10627 | w10682);
assign w10683 = v4996;
assign w10684 = w10627 & w10682;
assign v4997 = ~(w10683 | w10684);
assign w10685 = v4997;
assign v4998 = ~(w10562 | w10685);
assign w10686 = v4998;
assign w10687 = w10562 & w10685;
assign v4999 = ~(w10686 | w10687);
assign w10688 = v4999;
assign v5000 = ~(w10514 | w10688);
assign w10689 = v5000;
assign w10690 = w10514 & w10688;
assign v5001 = ~(w10689 | w10690);
assign w10691 = v5001;
assign w10692 = w10477 & ~w10691;
assign w10693 = ~w10477 & w10691;
assign v5002 = ~(w10692 | w10693);
assign w10694 = v5002;
assign w10695 = (w7754 & w17818) | (w7754 & w17819) | (w17818 & w17819);
assign w10696 = w10694 & w10695;
assign v5003 = ~(w10694 | w10695);
assign w10697 = v5003;
assign v5004 = ~(w10696 | w10697);
assign w10698 = v5004;
assign v5005 = ~(w10512 | w10690);
assign w10699 = v5005;
assign w10700 = (~w10560 & ~w10562) | (~w10560 & w17820) | (~w10562 & w17820);
assign w10701 = (~w10680 & ~w10682) | (~w10680 & w17467) | (~w10682 & w17467);
assign w10702 = (~w10526 & ~w10527) | (~w10526 & w17468) | (~w10527 & w17468);
assign w10703 = (~w10576 & ~w10578) | (~w10576 & w17614) | (~w10578 & w17614);
assign w10704 = (~w10543 & ~w10545) | (~w10543 & w17469) | (~w10545 & w17469);
assign w10705 = (~w10531 & ~w10533) | (~w10531 & w17615) | (~w10533 & w17615);
assign v5006 = ~(w10704 | w10705);
assign w10706 = v5006;
assign w10707 = w10704 & w10705;
assign v5007 = ~(w10706 | w10707);
assign w10708 = v5007;
assign w10709 = w10703 & ~w10708;
assign w10710 = ~w10703 & w10708;
assign v5008 = ~(w10709 | w10710);
assign w10711 = v5008;
assign w10712 = (~w10551 & ~w10553) | (~w10551 & w17616) | (~w10553 & w17616);
assign w10713 = (~w10518 & ~w10520) | (~w10518 & w17617) | (~w10520 & w17617);
assign v5009 = ~(w10712 | w10713);
assign w10714 = v5009;
assign w10715 = w10712 & w10713;
assign v5010 = ~(w10714 | w10715);
assign w10716 = v5010;
assign w10717 = w10711 & w10716;
assign v5011 = ~(w10711 | w10716);
assign w10718 = v5011;
assign v5012 = ~(w10717 | w10718);
assign w10719 = v5012;
assign w10720 = ~w10702 & w10719;
assign w10721 = w10702 & ~w10719;
assign v5013 = ~(w10720 | w10721);
assign w10722 = v5013;
assign w10723 = ~w10701 & w10722;
assign w10724 = w10701 & ~w10722;
assign v5014 = ~(w10723 | w10724);
assign w10725 = v5014;
assign w10726 = ~w10700 & w10725;
assign w10727 = w10700 & ~w10725;
assign v5015 = ~(w10726 | w10727);
assign w10728 = v5015;
assign v5016 = ~(w10493 | w10497);
assign w10729 = v5016;
assign w10730 = w10258 & ~w10486;
assign v5017 = ~(w10488 | w10730);
assign w10731 = v5017;
assign w10732 = w10446 & ~w10667;
assign v5018 = ~(w10669 | w10732);
assign w10733 = v5018;
assign v5019 = ~(w10731 | w10733);
assign w10734 = v5019;
assign w10735 = w10731 & w10733;
assign v5020 = ~(w10734 | w10735);
assign w10736 = v5020;
assign w10737 = pi14 & pi60;
assign w10738 = pi15 & pi59;
assign v5021 = ~(w10582 | w10738);
assign w10739 = v5021;
assign w10740 = pi16 & pi59;
assign w10741 = w10424 & w10740;
assign v5022 = ~(w10739 | w10741);
assign w10742 = v5022;
assign w10743 = w10737 & ~w10742;
assign w10744 = ~w10737 & w10742;
assign v5023 = ~(w10743 | w10744);
assign w10745 = v5023;
assign w10746 = ~w10736 & w10745;
assign w10747 = w10736 & ~w10745;
assign v5024 = ~(w10746 | w10747);
assign w10748 = v5024;
assign v5025 = ~(w10607 | w10619);
assign w10749 = v5025;
assign w10750 = w10748 & ~w10749;
assign w10751 = ~w10748 & w10749;
assign v5026 = ~(w10750 | w10751);
assign w10752 = v5026;
assign w10753 = w10729 & ~w10752;
assign w10754 = ~w10729 & w10752;
assign v5027 = ~(w10753 | w10754);
assign w10755 = v5027;
assign v5028 = ~(w10622 | w10626);
assign w10756 = v5028;
assign w10757 = (~w10643 & ~w10644) | (~w10643 & w17184) | (~w10644 & w17184);
assign v5029 = ~(w10756 | w10757);
assign w10758 = v5029;
assign w10759 = w10756 & w10757;
assign v5030 = ~(w10758 | w10759);
assign w10760 = v5030;
assign w10761 = w10755 & w10760;
assign v5031 = ~(w10755 | w10760);
assign w10762 = v5031;
assign v5032 = ~(w10761 | w10762);
assign w10763 = v5032;
assign w10764 = (w10763 & w10509) | (w10763 & w17618) | (w10509 & w17618);
assign w10765 = ~w10509 & w17619;
assign v5033 = ~(w10764 | w10765);
assign w10766 = v5033;
assign w10767 = w10566 & ~w10569;
assign v5034 = ~(w10571 | w10767);
assign w10768 = v5034;
assign w10769 = w10433 & ~w10647;
assign v5035 = ~(w10649 | w10769);
assign w10770 = v5035;
assign v5036 = ~(w10768 | w10770);
assign w10771 = v5036;
assign w10772 = w10768 & w10770;
assign v5037 = ~(w10771 | w10772);
assign w10773 = v5037;
assign w10774 = w10579 & ~w10581;
assign v5038 = ~(w10583 | w10774);
assign w10775 = v5038;
assign w10776 = ~w10773 & w10775;
assign w10777 = w10773 & ~w10775;
assign v5039 = ~(w10776 | w10777);
assign w10778 = v5039;
assign v5040 = ~(w10598 | w10602);
assign w10779 = v5040;
assign v5041 = ~(w10601 | w10779);
assign w10780 = v5041;
assign w10781 = w10371 & ~w10612;
assign v5042 = ~(w10614 | w10781);
assign w10782 = v5042;
assign w10783 = w10780 & ~w10782;
assign w10784 = ~w10780 & w10782;
assign v5043 = ~(w10783 | w10784);
assign w10785 = v5043;
assign v5044 = ~(w10345 | w10657);
assign w10786 = v5044;
assign v5045 = ~(w10656 | w10786);
assign w10787 = v5045;
assign v5046 = ~(w10785 | w10787);
assign w10788 = v5046;
assign w10789 = w10785 & w10787;
assign v5047 = ~(w10788 | w10789);
assign w10790 = v5047;
assign w10791 = (~w10662 & ~w10664) | (~w10662 & w17470) | (~w10664 & w17470);
assign w10792 = ~w10790 & w10791;
assign w10793 = w10790 & ~w10791;
assign v5048 = ~(w10792 | w10793);
assign w10794 = v5048;
assign w10795 = w10778 & w10794;
assign v5049 = ~(w10778 | w10794);
assign w10796 = v5049;
assign v5050 = ~(w10795 | w10796);
assign w10797 = v5050;
assign w10798 = (w10797 & w10503) | (w10797 & w17471) | (w10503 & w17471);
assign w10799 = ~w10503 & w17472;
assign v5051 = ~(w10798 | w10799);
assign w10800 = v5051;
assign v5052 = ~(w10633 | w10639);
assign w10801 = v5052;
assign w10802 = pi13 & pi61;
assign w10803 = pi12 & pi62;
assign v5053 = ~(w10802 | w10803);
assign w10804 = v5053;
assign w10805 = pi13 & pi62;
assign w10806 = w10655 & w10805;
assign v5054 = ~(w10804 | w10806);
assign w10807 = v5054;
assign w10808 = w10591 & ~w10593;
assign v5055 = ~(w10592 | w10808);
assign w10809 = v5055;
assign w10810 = w10807 & ~w10809;
assign w10811 = ~w10807 & w10809;
assign v5056 = ~(w10810 | w10811);
assign w10812 = v5056;
assign w10813 = pi29 & pi45;
assign w10814 = pi17 & pi57;
assign v5057 = ~(w10648 | w10814);
assign w10815 = v5057;
assign w10816 = w10648 & w10814;
assign v5058 = ~(w10815 | w10816);
assign w10817 = v5058;
assign w10818 = w10813 & ~w10817;
assign w10819 = ~w10813 & w10817;
assign v5059 = ~(w10818 | w10819);
assign w10820 = v5059;
assign w10821 = w10812 & ~w10820;
assign w10822 = ~w10812 & w10820;
assign v5060 = ~(w10821 | w10822);
assign w10823 = v5060;
assign w10824 = w10801 & ~w10823;
assign w10825 = ~w10801 & w10823;
assign v5061 = ~(w10824 | w10825);
assign w10826 = v5061;
assign w10827 = pi11 & pi63;
assign w10828 = pi31 & pi43;
assign w10829 = pi32 & pi42;
assign v5062 = ~(w10828 | w10829);
assign w10830 = v5062;
assign w10831 = pi32 & pi43;
assign w10832 = w10258 & w10831;
assign v5063 = ~(w10830 | w10832);
assign w10833 = v5063;
assign w10834 = w10827 & ~w10833;
assign w10835 = ~w10827 & w10833;
assign v5064 = ~(w10834 | w10835);
assign w10836 = v5064;
assign w10837 = pi18 & pi56;
assign w10838 = pi25 & pi49;
assign v5065 = ~(w10837 | w10838);
assign w10839 = v5065;
assign w10840 = w10837 & w10838;
assign v5066 = ~(w10839 | w10840);
assign w10841 = v5066;
assign w10842 = w10487 & ~w10841;
assign w10843 = ~w10487 & w10841;
assign v5067 = ~(w10842 | w10843);
assign w10844 = v5067;
assign v5068 = ~(w10836 | w10844);
assign w10845 = v5068;
assign w10846 = w10836 & w10844;
assign v5069 = ~(w10845 | w10846);
assign w10847 = v5069;
assign w10848 = pi26 & pi48;
assign w10849 = pi28 & pi46;
assign v5070 = ~(w10570 | w10849);
assign w10850 = v5070;
assign w10851 = pi28 & pi47;
assign w10852 = w10568 & w10851;
assign v5071 = ~(w10850 | w10852);
assign w10853 = v5071;
assign w10854 = w10848 & ~w10853;
assign w10855 = ~w10848 & w10853;
assign v5072 = ~(w10854 | w10855);
assign w10856 = v5072;
assign w10857 = w10847 & ~w10856;
assign w10858 = ~w10847 & w10856;
assign v5073 = ~(w10857 | w10858);
assign w10859 = v5073;
assign w10860 = pi20 & pi54;
assign w10861 = pi35 & pi39;
assign w10862 = pi34 & pi40;
assign v5074 = ~(w10861 | w10862);
assign w10863 = v5074;
assign w10864 = pi35 & pi40;
assign w10865 = w10446 & w10864;
assign v5075 = ~(w10863 | w10865);
assign w10866 = v5075;
assign w10867 = w10860 & ~w10866;
assign w10868 = ~w10860 & w10866;
assign v5076 = ~(w10867 | w10868);
assign w10869 = v5076;
assign w10870 = pi22 & pi52;
assign w10871 = pi19 & pi55;
assign v5077 = ~(w10613 | w10871);
assign w10872 = v5077;
assign w10873 = w10613 & w10871;
assign v5078 = ~(w10872 | w10873);
assign w10874 = v5078;
assign w10875 = w10870 & ~w10874;
assign w10876 = ~w10870 & w10874;
assign v5079 = ~(w10875 | w10876);
assign w10877 = v5079;
assign v5080 = ~(w10869 | w10877);
assign w10878 = v5080;
assign w10879 = w10869 & w10877;
assign v5081 = ~(w10878 | w10879);
assign w10880 = v5081;
assign w10881 = pi23 & pi51;
assign w10882 = pi24 & pi50;
assign v5082 = ~(w10881 | w10882);
assign w10883 = v5082;
assign w10884 = pi24 & pi51;
assign w10885 = w10591 & w10884;
assign v5083 = ~(w10883 | w10885);
assign w10886 = v5083;
assign w10887 = w10668 & ~w10886;
assign w10888 = ~w10668 & w10886;
assign v5084 = ~(w10887 | w10888);
assign w10889 = v5084;
assign w10890 = w10880 & ~w10889;
assign w10891 = ~w10880 & w10889;
assign v5085 = ~(w10890 | w10891);
assign w10892 = v5085;
assign w10893 = w10859 & w10892;
assign v5086 = ~(w10859 | w10892);
assign w10894 = v5086;
assign v5087 = ~(w10893 | w10894);
assign w10895 = v5087;
assign v5088 = ~(w10826 | w10895);
assign w10896 = v5088;
assign w10897 = w10826 & w10895;
assign v5089 = ~(w10896 | w10897);
assign w10898 = v5089;
assign v5090 = ~(w10800 | w10898);
assign w10899 = v5090;
assign w10900 = w10800 & w10898;
assign v5091 = ~(w10899 | w10900);
assign w10901 = v5091;
assign w10902 = w10766 & w10901;
assign v5092 = ~(w10766 | w10901);
assign w10903 = v5092;
assign v5093 = ~(w10902 | w10903);
assign w10904 = v5093;
assign w10905 = w10728 & w10904;
assign v5094 = ~(w10728 | w10904);
assign w10906 = v5094;
assign v5095 = ~(w10905 | w10906);
assign w10907 = v5095;
assign w10908 = w10699 & ~w10907;
assign w10909 = ~w10699 & w10907;
assign v5096 = ~(w10908 | w10909);
assign w10910 = v5096;
assign v5097 = ~(w10471 | w10692);
assign w10911 = v5097;
assign w10912 = (~w8795 & w17620) | (~w8795 & w17621) | (w17620 & w17621);
assign w10913 = w10910 & w10912;
assign v5098 = ~(w10910 | w10912);
assign w10914 = v5098;
assign v5099 = ~(w10913 | w10914);
assign w10915 = v5099;
assign v5100 = ~(w10726 | w10905);
assign w10916 = v5100;
assign w10917 = (~w10771 & ~w10773) | (~w10771 & w17185) | (~w10773 & w17185);
assign w10918 = (~w10734 & ~w10736) | (~w10734 & w16770) | (~w10736 & w16770);
assign w10919 = (~w10783 & ~w10785) | (~w10783 & w16771) | (~w10785 & w16771);
assign v5101 = ~(w10918 | w10919);
assign w10920 = v5101;
assign w10921 = w10918 & w10919;
assign v5102 = ~(w10920 | w10921);
assign w10922 = v5102;
assign w10923 = w10917 & ~w10922;
assign w10924 = ~w10917 & w10922;
assign v5103 = ~(w10923 | w10924);
assign w10925 = v5103;
assign w10926 = (~w10893 & ~w10895) | (~w10893 & w17821) | (~w10895 & w17821);
assign w10927 = ~w10925 & w10926;
assign w10928 = w10925 & ~w10926;
assign v5104 = ~(w10927 | w10928);
assign w10929 = v5104;
assign v5105 = ~(w10821 | w10825);
assign w10930 = v5105;
assign w10931 = w10668 & ~w10883;
assign v5106 = ~(w10885 | w10931);
assign w10932 = v5106;
assign w10933 = w10860 & ~w10863;
assign v5107 = ~(w10865 | w10933);
assign w10934 = v5107;
assign v5108 = ~(w10932 | w10934);
assign w10935 = v5108;
assign w10936 = w10932 & w10934;
assign v5109 = ~(w10935 | w10936);
assign w10937 = v5109;
assign v5110 = ~(w10870 | w10873);
assign w10938 = v5110;
assign v5111 = ~(w10872 | w10938);
assign w10939 = v5111;
assign v5112 = ~(w10937 | w10939);
assign w10940 = v5112;
assign w10941 = w10937 & w10939;
assign v5113 = ~(w10940 | w10941);
assign w10942 = v5113;
assign w10943 = (~w10806 & w10809) | (~w10806 & w17186) | (w10809 & w17186);
assign v5114 = ~(w10487 | w10840);
assign w10944 = v5114;
assign v5115 = ~(w10839 | w10944);
assign w10945 = v5115;
assign w10946 = w10827 & ~w10830;
assign v5116 = ~(w10832 | w10946);
assign w10947 = v5116;
assign w10948 = w10945 & ~w10947;
assign w10949 = ~w10945 & w10947;
assign v5117 = ~(w10948 | w10949);
assign w10950 = v5117;
assign w10951 = w10943 & ~w10950;
assign w10952 = ~w10943 & w10950;
assign v5118 = ~(w10951 | w10952);
assign w10953 = v5118;
assign w10954 = w10942 & w10953;
assign v5119 = ~(w10942 | w10953);
assign w10955 = v5119;
assign v5120 = ~(w10954 | w10955);
assign w10956 = v5120;
assign w10957 = ~w10930 & w10956;
assign w10958 = w10930 & ~w10956;
assign v5121 = ~(w10957 | w10958);
assign w10959 = v5121;
assign w10960 = w10929 & w10959;
assign v5122 = ~(w10929 | w10959);
assign w10961 = v5122;
assign v5123 = ~(w10960 | w10961);
assign w10962 = v5123;
assign w10963 = (w10962 & w10723) | (w10962 & w17622) | (w10723 & w17622);
assign w10964 = ~w10723 & w17623;
assign v5124 = ~(w10963 | w10964);
assign w10965 = v5124;
assign w10966 = (~w10714 & ~w10716) | (~w10714 & w17822) | (~w10716 & w17822);
assign v5125 = ~(w10813 | w10816);
assign w10967 = v5125;
assign v5126 = ~(w10815 | w10967);
assign w10968 = v5126;
assign w10969 = w10848 & ~w10850;
assign v5127 = ~(w10852 | w10969);
assign w10970 = v5127;
assign w10971 = w10968 & ~w10970;
assign w10972 = ~w10968 & w10970;
assign v5128 = ~(w10971 | w10972);
assign w10973 = v5128;
assign w10974 = w10737 & ~w10739;
assign v5129 = ~(w10741 | w10974);
assign w10975 = v5129;
assign w10976 = ~w10973 & w10975;
assign w10977 = w10973 & ~w10975;
assign v5130 = ~(w10976 | w10977);
assign w10978 = v5130;
assign w10979 = (~w10878 & ~w10880) | (~w10878 & w16936) | (~w10880 & w16936);
assign w10980 = (~w10845 & ~w10847) | (~w10845 & w16937) | (~w10847 & w16937);
assign v5131 = ~(w10979 | w10980);
assign w10981 = v5131;
assign w10982 = w10979 & w10980;
assign v5132 = ~(w10981 | w10982);
assign w10983 = v5132;
assign w10984 = w10978 & w10983;
assign v5133 = ~(w10978 | w10983);
assign w10985 = v5133;
assign v5134 = ~(w10984 | w10985);
assign w10986 = v5134;
assign w10987 = ~w10966 & w10986;
assign w10988 = w10966 & ~w10986;
assign v5135 = ~(w10987 | w10988);
assign w10989 = v5135;
assign w10990 = (~w10706 & ~w10708) | (~w10706 & w17624) | (~w10708 & w17624);
assign w10991 = pi23 & pi52;
assign w10992 = pi36 & pi39;
assign v5136 = ~(w10864 | w10992);
assign w10993 = v5136;
assign w10994 = w10864 & w10992;
assign v5137 = ~(w10993 | w10994);
assign w10995 = v5137;
assign w10996 = w10991 & ~w10995;
assign w10997 = ~w10991 & w10995;
assign v5138 = ~(w10996 | w10997);
assign w10998 = v5138;
assign w10999 = pi30 & pi45;
assign w11000 = pi12 & pi63;
assign w11001 = pi19 & pi56;
assign v5139 = ~(w11000 | w11001);
assign w11002 = v5139;
assign w11003 = w11000 & w11001;
assign v5140 = ~(w11002 | w11003);
assign w11004 = v5140;
assign w11005 = w10999 & ~w11004;
assign w11006 = ~w10999 & w11004;
assign v5141 = ~(w11005 | w11006);
assign w11007 = v5141;
assign v5142 = ~(w10998 | w11007);
assign w11008 = v5142;
assign w11009 = w10998 & w11007;
assign v5143 = ~(w11008 | w11009);
assign w11010 = v5143;
assign w11011 = ~pi37 & pi38;
assign w11012 = w10805 & ~w11011;
assign w11013 = ~w10805 & w11011;
assign v5144 = ~(w11012 | w11013);
assign w11014 = v5144;
assign w11015 = w11010 & ~w11014;
assign w11016 = ~w11010 & w11014;
assign v5145 = ~(w11015 | w11016);
assign w11017 = v5145;
assign w11018 = ~w10990 & w11017;
assign w11019 = w10990 & ~w11017;
assign v5146 = ~(w11018 | w11019);
assign w11020 = v5146;
assign w11021 = pi14 & pi61;
assign w11022 = pi15 & pi60;
assign v5147 = ~(w10740 | w11022);
assign w11023 = v5147;
assign w11024 = pi16 & pi60;
assign w11025 = w10738 & w11024;
assign v5148 = ~(w11023 | w11025);
assign w11026 = v5148;
assign w11027 = w11021 & ~w11026;
assign w11028 = ~w11021 & w11026;
assign v5149 = ~(w11027 | w11028);
assign w11029 = v5149;
assign w11030 = pi17 & pi58;
assign w11031 = pi26 & pi49;
assign w11032 = pi18 & pi57;
assign v5150 = ~(w11031 | w11032);
assign w11033 = v5150;
assign w11034 = w11031 & w11032;
assign v5151 = ~(w11033 | w11034);
assign w11035 = v5151;
assign w11036 = w11030 & ~w11035;
assign w11037 = ~w11030 & w11035;
assign v5152 = ~(w11036 | w11037);
assign w11038 = v5152;
assign v5153 = ~(w11029 | w11038);
assign w11039 = v5153;
assign w11040 = w11029 & w11038;
assign v5154 = ~(w11039 | w11040);
assign w11041 = v5154;
assign w11042 = pi27 & pi48;
assign w11043 = pi29 & pi46;
assign v5155 = ~(w10851 | w11043);
assign w11044 = v5155;
assign w11045 = pi29 & pi47;
assign w11046 = w10849 & w11045;
assign v5156 = ~(w11044 | w11046);
assign w11047 = v5156;
assign w11048 = w11042 & ~w11047;
assign w11049 = ~w11042 & w11047;
assign v5157 = ~(w11048 | w11049);
assign w11050 = v5157;
assign w11051 = w11041 & ~w11050;
assign w11052 = ~w11041 & w11050;
assign v5158 = ~(w11051 | w11052);
assign w11053 = v5158;
assign w11054 = w11020 & w11053;
assign v5159 = ~(w11020 | w11053);
assign w11055 = v5159;
assign v5160 = ~(w11054 | w11055);
assign w11056 = v5160;
assign w11057 = w10989 & w11056;
assign v5161 = ~(w10989 | w11056);
assign w11058 = v5161;
assign v5162 = ~(w11057 | w11058);
assign w11059 = v5162;
assign v5163 = ~(w10965 | w11059);
assign w11060 = v5163;
assign w11061 = w10965 & w11059;
assign v5164 = ~(w11060 | w11061);
assign w11062 = v5164;
assign w11063 = (~w10798 & ~w10800) | (~w10798 & w17625) | (~w10800 & w17625);
assign w11064 = (~w10758 & ~w10760) | (~w10758 & w17474) | (~w10760 & w17474);
assign v5165 = ~(w10750 | w10754);
assign w11065 = v5165;
assign w11066 = (~w10793 & ~w10794) | (~w10793 & w17626) | (~w10794 & w17626);
assign w11067 = pi31 & pi44;
assign w11068 = pi33 & pi42;
assign v5166 = ~(w10831 | w11068);
assign w11069 = v5166;
assign w11070 = pi33 & pi43;
assign w11071 = w10829 & w11070;
assign v5167 = ~(w11069 | w11071);
assign w11072 = v5167;
assign w11073 = w11067 & ~w11072;
assign w11074 = ~w11067 & w11072;
assign v5168 = ~(w11073 | w11074);
assign w11075 = v5168;
assign w11076 = pi34 & pi41;
assign w11077 = pi20 & pi55;
assign w11078 = pi25 & pi50;
assign v5169 = ~(w11077 | w11078);
assign w11079 = v5169;
assign w11080 = w11077 & w11078;
assign v5170 = ~(w11079 | w11080);
assign w11081 = v5170;
assign w11082 = w11076 & ~w11081;
assign w11083 = ~w11076 & w11081;
assign v5171 = ~(w11082 | w11083);
assign w11084 = v5171;
assign v5172 = ~(w11075 | w11084);
assign w11085 = v5172;
assign w11086 = w11075 & w11084;
assign v5173 = ~(w11085 | w11086);
assign w11087 = v5173;
assign w11088 = pi21 & pi54;
assign w11089 = pi22 & pi53;
assign v5174 = ~(w10884 | w11089);
assign w11090 = v5174;
assign w11091 = w10884 & w11089;
assign v5175 = ~(w11090 | w11091);
assign w11092 = v5175;
assign w11093 = w11088 & ~w11092;
assign w11094 = ~w11088 & w11092;
assign v5176 = ~(w11093 | w11094);
assign w11095 = v5176;
assign w11096 = w11087 & ~w11095;
assign w11097 = ~w11087 & w11095;
assign v5177 = ~(w11096 | w11097);
assign w11098 = v5177;
assign w11099 = ~w11066 & w11098;
assign w11100 = w11066 & ~w11098;
assign v5178 = ~(w11099 | w11100);
assign w11101 = v5178;
assign w11102 = ~w11065 & w11101;
assign w11103 = w11065 & ~w11101;
assign v5179 = ~(w11102 | w11103);
assign w11104 = v5179;
assign w11105 = ~w11064 & w11104;
assign w11106 = w11064 & ~w11104;
assign v5180 = ~(w11105 | w11106);
assign w11107 = v5180;
assign w11108 = w11063 & ~w11107;
assign w11109 = ~w11063 & w11107;
assign v5181 = ~(w11108 | w11109);
assign w11110 = v5181;
assign w11111 = (~w10764 & ~w10766) | (~w10764 & w17823) | (~w10766 & w17823);
assign w11112 = ~w11110 & w11111;
assign w11113 = w11110 & ~w11111;
assign v5182 = ~(w11112 | w11113);
assign w11114 = v5182;
assign w11115 = w11062 & w11114;
assign v5183 = ~(w11062 | w11114);
assign w11116 = v5183;
assign v5184 = ~(w11115 | w11116);
assign w11117 = v5184;
assign w11118 = ~w10916 & w11117;
assign w11119 = w10916 & ~w11117;
assign v5185 = ~(w11118 | w11119);
assign w11120 = v5185;
assign v5186 = ~(w10693 | w10909);
assign w11121 = v5186;
assign w11122 = (w8795 & w17475) | (w8795 & w17476) | (w17475 & w17476);
assign w11123 = w11120 & w11122;
assign v5187 = ~(w11120 | w11122);
assign w11124 = v5187;
assign v5188 = ~(w11123 | w11124);
assign w11125 = v5188;
assign v5189 = ~(w11113 | w11115);
assign w11126 = v5189;
assign w11127 = (~w10963 & ~w10965) | (~w10963 & w17824) | (~w10965 & w17824);
assign v5190 = ~(w10987 | w11057);
assign w11128 = v5190;
assign v5191 = ~(w10928 | w10960);
assign w11129 = v5191;
assign v5192 = ~(w10954 | w10957);
assign w11130 = v5192;
assign w11131 = (~w10981 & ~w10983) | (~w10981 & w17187) | (~w10983 & w17187);
assign w11132 = pi13 & pi63;
assign w11133 = pi31 & pi45;
assign w11134 = pi32 & pi44;
assign v5193 = ~(w11133 | w11134);
assign w11135 = v5193;
assign w11136 = pi32 & pi45;
assign w11137 = w11067 & w11136;
assign v5194 = ~(w11135 | w11137);
assign w11138 = v5194;
assign w11139 = w11132 & ~w11138;
assign w11140 = ~w11132 & w11138;
assign v5195 = ~(w11139 | w11140);
assign w11141 = v5195;
assign w11142 = pi19 & pi57;
assign w11143 = pi23 & pi53;
assign v5196 = ~(w11142 | w11143);
assign w11144 = v5196;
assign w11145 = w11142 & w11143;
assign v5197 = ~(w11144 | w11145);
assign w11146 = v5197;
assign w11147 = w11070 & ~w11146;
assign w11148 = ~w11070 & w11146;
assign v5198 = ~(w11147 | w11148);
assign w11149 = v5198;
assign v5199 = ~(w11141 | w11149);
assign w11150 = v5199;
assign w11151 = w11141 & w11149;
assign v5200 = ~(w11150 | w11151);
assign w11152 = v5200;
assign w11153 = pi20 & pi56;
assign w11154 = pi21 & pi55;
assign w11155 = pi22 & pi54;
assign v5201 = ~(w11154 | w11155);
assign w11156 = v5201;
assign w11157 = pi22 & pi55;
assign w11158 = w11088 & w11157;
assign v5202 = ~(w11156 | w11158);
assign w11159 = v5202;
assign w11160 = w11153 & ~w11159;
assign w11161 = ~w11153 & w11159;
assign v5203 = ~(w11160 | w11161);
assign w11162 = v5203;
assign w11163 = w11152 & ~w11162;
assign w11164 = ~w11152 & w11162;
assign v5204 = ~(w11163 | w11164);
assign w11165 = v5204;
assign w11166 = ~w11131 & w11165;
assign w11167 = w11131 & ~w11165;
assign v5205 = ~(w11166 | w11167);
assign w11168 = v5205;
assign w11169 = ~w11130 & w11168;
assign w11170 = w11130 & ~w11168;
assign v5206 = ~(w11169 | w11170);
assign w11171 = v5206;
assign w11172 = ~w11129 & w11171;
assign w11173 = w11129 & ~w11171;
assign v5207 = ~(w11172 | w11173);
assign w11174 = v5207;
assign w11175 = ~w11128 & w11174;
assign w11176 = w11128 & ~w11174;
assign v5208 = ~(w11175 | w11176);
assign w11177 = v5208;
assign w11178 = ~w11127 & w11177;
assign w11179 = w11127 & ~w11177;
assign v5209 = ~(w11178 | w11179);
assign w11180 = v5209;
assign v5210 = ~(w10935 | w10941);
assign w11181 = v5210;
assign w11182 = (~w10948 & ~w10950) | (~w10948 & w17188) | (~w10950 & w17188);
assign w11183 = (~w10971 & ~w10973) | (~w10971 & w17189) | (~w10973 & w17189);
assign v5211 = ~(w11182 | w11183);
assign w11184 = v5211;
assign w11185 = w11182 & w11183;
assign v5212 = ~(w11184 | w11185);
assign w11186 = v5212;
assign w11187 = w11181 & ~w11186;
assign w11188 = ~w11181 & w11186;
assign v5213 = ~(w11187 | w11188);
assign w11189 = v5213;
assign w11190 = (~w11018 & ~w11020) | (~w11018 & w17825) | (~w11020 & w17825);
assign w11191 = ~w11189 & w11190;
assign w11192 = w11189 & ~w11190;
assign v5214 = ~(w11191 | w11192);
assign w11193 = v5214;
assign v5215 = ~(w11076 | w11080);
assign w11194 = v5215;
assign v5216 = ~(w11079 | w11194);
assign w11195 = v5216;
assign w11196 = w11042 & ~w11044;
assign v5217 = ~(w11046 | w11196);
assign w11197 = v5217;
assign w11198 = w11195 & ~w11197;
assign w11199 = ~w11195 & w11197;
assign v5218 = ~(w11198 | w11199);
assign w11200 = v5218;
assign v5219 = ~(w10999 | w11003);
assign w11201 = v5219;
assign v5220 = ~(w11002 | w11201);
assign w11202 = v5220;
assign v5221 = ~(w11200 | w11202);
assign w11203 = v5221;
assign w11204 = w11200 & w11202;
assign v5222 = ~(w11203 | w11204);
assign w11205 = v5222;
assign v5223 = ~(w11085 | w11096);
assign w11206 = v5223;
assign w11207 = pi14 & pi62;
assign v5224 = ~(pi37 | w10805);
assign w11208 = v5224;
assign w11209 = pi38 & ~w11208;
assign v5225 = ~(w11207 | w11209);
assign w11210 = v5225;
assign w11211 = w11207 & w11209;
assign v5226 = ~(w11210 | w11211);
assign w11212 = v5226;
assign v5227 = ~(w10991 | w10994);
assign w11213 = v5227;
assign v5228 = ~(w10993 | w11213);
assign w11214 = v5228;
assign w11215 = ~w11212 & w11214;
assign w11216 = w11212 & ~w11214;
assign v5229 = ~(w11215 | w11216);
assign w11217 = v5229;
assign v5230 = ~(w11206 | w11217);
assign w11218 = v5230;
assign w11219 = w11206 & w11217;
assign v5231 = ~(w11218 | w11219);
assign w11220 = v5231;
assign v5232 = ~(w11205 | w11220);
assign w11221 = v5232;
assign w11222 = w11205 & w11220;
assign v5233 = ~(w11221 | w11222);
assign w11223 = v5233;
assign v5234 = ~(w11193 | w11223);
assign w11224 = v5234;
assign w11225 = w11193 & w11223;
assign v5235 = ~(w11224 | w11225);
assign w11226 = v5235;
assign w11227 = (~w11105 & ~w11107) | (~w11105 & w17627) | (~w11107 & w17627);
assign w11228 = w11226 & ~w11227;
assign w11229 = ~w11226 & w11227;
assign v5236 = ~(w11228 | w11229);
assign w11230 = v5236;
assign v5237 = ~(w11099 | w11102);
assign w11231 = v5237;
assign v5238 = ~(w11030 | w11034);
assign w11232 = v5238;
assign v5239 = ~(w11033 | w11232);
assign w11233 = v5239;
assign w11234 = w11021 & ~w11023;
assign v5240 = ~(w11025 | w11234);
assign w11235 = v5240;
assign w11236 = w11233 & ~w11235;
assign w11237 = ~w11233 & w11235;
assign v5241 = ~(w11236 | w11237);
assign w11238 = v5241;
assign w11239 = w11067 & ~w11069;
assign v5242 = ~(w11071 | w11239);
assign w11240 = v5242;
assign w11241 = ~w11238 & w11240;
assign w11242 = w11238 & ~w11240;
assign v5243 = ~(w11241 | w11242);
assign w11243 = v5243;
assign w11244 = (~w11039 & ~w11041) | (~w11039 & w16938) | (~w11041 & w16938);
assign w11245 = (~w11008 & ~w11010) | (~w11008 & w16939) | (~w11010 & w16939);
assign v5244 = ~(w11244 | w11245);
assign w11246 = v5244;
assign w11247 = w11244 & w11245;
assign v5245 = ~(w11246 | w11247);
assign w11248 = v5245;
assign w11249 = w11243 & w11248;
assign v5246 = ~(w11243 | w11248);
assign w11250 = v5246;
assign v5247 = ~(w11249 | w11250);
assign w11251 = v5247;
assign w11252 = ~w11231 & w11251;
assign w11253 = w11231 & ~w11251;
assign v5248 = ~(w11252 | w11253);
assign w11254 = v5248;
assign w11255 = (~w10920 & ~w10922) | (~w10920 & w16940) | (~w10922 & w16940);
assign w11256 = pi28 & pi48;
assign w11257 = pi30 & pi46;
assign v5249 = ~(w11045 | w11257);
assign w11258 = v5249;
assign w11259 = pi30 & pi47;
assign w11260 = w11043 & w11259;
assign v5250 = ~(w11258 | w11260);
assign w11261 = v5250;
assign w11262 = w11256 & ~w11261;
assign w11263 = ~w11256 & w11261;
assign v5251 = ~(w11262 | w11263);
assign w11264 = v5251;
assign w11265 = pi34 & pi42;
assign w11266 = pi36 & pi40;
assign w11267 = pi35 & pi41;
assign v5252 = ~(w11266 | w11267);
assign w11268 = v5252;
assign w11269 = pi36 & pi41;
assign w11270 = w10864 & w11269;
assign v5253 = ~(w11268 | w11270);
assign w11271 = v5253;
assign w11272 = w11265 & ~w11271;
assign w11273 = ~w11265 & w11271;
assign v5254 = ~(w11272 | w11273);
assign w11274 = v5254;
assign v5255 = ~(w11264 | w11274);
assign w11275 = v5255;
assign w11276 = w11264 & w11274;
assign v5256 = ~(w11275 | w11276);
assign w11277 = v5256;
assign w11278 = pi37 & pi39;
assign w11279 = pi25 & pi51;
assign w11280 = pi24 & pi52;
assign v5257 = ~(w11279 | w11280);
assign w11281 = v5257;
assign w11282 = pi25 & pi52;
assign w11283 = w10884 & w11282;
assign v5258 = ~(w11281 | w11283);
assign w11284 = v5258;
assign w11285 = w11278 & ~w11284;
assign w11286 = ~w11278 & w11284;
assign v5259 = ~(w11285 | w11286);
assign w11287 = v5259;
assign w11288 = w11277 & ~w11287;
assign w11289 = ~w11277 & w11287;
assign v5260 = ~(w11288 | w11289);
assign w11290 = v5260;
assign w11291 = ~w11255 & w11290;
assign w11292 = w11255 & ~w11290;
assign v5261 = ~(w11291 | w11292);
assign w11293 = v5261;
assign v5262 = ~(w11088 | w11091);
assign w11294 = v5262;
assign v5263 = ~(w11090 | w11294);
assign w11295 = v5263;
assign w11296 = pi15 & pi61;
assign w11297 = pi17 & pi59;
assign v5264 = ~(w11024 | w11297);
assign w11298 = v5264;
assign w11299 = pi17 & pi60;
assign w11300 = w10740 & w11299;
assign v5265 = ~(w11298 | w11300);
assign w11301 = v5265;
assign w11302 = w11296 & ~w11301;
assign w11303 = ~w11296 & w11301;
assign v5266 = ~(w11302 | w11303);
assign w11304 = v5266;
assign w11305 = w11295 & ~w11304;
assign w11306 = ~w11295 & w11304;
assign v5267 = ~(w11305 | w11306);
assign w11307 = v5267;
assign w11308 = pi18 & pi58;
assign w11309 = pi26 & pi50;
assign w11310 = pi27 & pi49;
assign v5268 = ~(w11309 | w11310);
assign w11311 = v5268;
assign w11312 = pi27 & pi50;
assign w11313 = w11031 & w11312;
assign v5269 = ~(w11311 | w11313);
assign w11314 = v5269;
assign w11315 = w11308 & ~w11314;
assign w11316 = ~w11308 & w11314;
assign v5270 = ~(w11315 | w11316);
assign w11317 = v5270;
assign w11318 = w11307 & ~w11317;
assign w11319 = ~w11307 & w11317;
assign v5271 = ~(w11318 | w11319);
assign w11320 = v5271;
assign w11321 = w11293 & w11320;
assign v5272 = ~(w11293 | w11320);
assign w11322 = v5272;
assign v5273 = ~(w11321 | w11322);
assign w11323 = v5273;
assign w11324 = w11254 & w11323;
assign v5274 = ~(w11254 | w11323);
assign w11325 = v5274;
assign v5275 = ~(w11324 | w11325);
assign w11326 = v5275;
assign w11327 = w11230 & w11326;
assign v5276 = ~(w11230 | w11326);
assign w11328 = v5276;
assign v5277 = ~(w11327 | w11328);
assign w11329 = v5277;
assign w11330 = w11180 & w11329;
assign v5278 = ~(w11180 | w11329);
assign w11331 = v5278;
assign v5279 = ~(w11330 | w11331);
assign w11332 = v5279;
assign w11333 = ~w11126 & w11332;
assign w11334 = w11126 & ~w11332;
assign v5280 = ~(w11333 | w11334);
assign w11335 = v5280;
assign w11336 = (w7754 & w17826) | (w7754 & w17827) | (w17826 & w17827);
assign w11337 = w11335 & w11336;
assign v5281 = ~(w11335 | w11336);
assign w11338 = v5281;
assign v5282 = ~(w11337 | w11338);
assign w11339 = v5282;
assign v5283 = ~(w11178 | w11330);
assign w11340 = v5283;
assign w11341 = (~w11228 & ~w11230) | (~w11228 & w17828) | (~w11230 & w17828);
assign v5284 = ~(w11252 | w11324);
assign w11342 = v5284;
assign v5285 = ~(w11192 | w11225);
assign w11343 = v5285;
assign v5286 = ~(w11218 | w11222);
assign w11344 = v5286;
assign w11345 = (~w11246 & ~w11248) | (~w11246 & w17190) | (~w11248 & w17190);
assign w11346 = pi24 & pi53;
assign w11347 = pi23 & pi54;
assign v5287 = ~(w11346 | w11347);
assign w11348 = v5287;
assign w11349 = pi24 & pi54;
assign w11350 = w11143 & w11349;
assign v5288 = ~(w11348 | w11350);
assign w11351 = v5288;
assign w11352 = w11282 & ~w11351;
assign w11353 = ~w11282 & w11351;
assign v5289 = ~(w11352 | w11353);
assign w11354 = v5289;
assign w11355 = pi34 & pi43;
assign w11356 = pi26 & pi51;
assign v5290 = ~(w11157 | w11356);
assign w11357 = v5290;
assign w11358 = w11157 & w11356;
assign v5291 = ~(w11357 | w11358);
assign w11359 = v5291;
assign w11360 = w11355 & ~w11359;
assign w11361 = ~w11355 & w11359;
assign v5292 = ~(w11360 | w11361);
assign w11362 = v5292;
assign v5293 = ~(w11354 | w11362);
assign w11363 = v5293;
assign w11364 = w11354 & w11362;
assign v5294 = ~(w11363 | w11364);
assign w11365 = v5294;
assign w11366 = pi16 & pi61;
assign w11367 = pi33 & pi44;
assign v5295 = ~(w11136 | w11367);
assign w11368 = v5295;
assign w11369 = pi33 & pi45;
assign w11370 = w11134 & w11369;
assign v5296 = ~(w11368 | w11370);
assign w11371 = v5296;
assign w11372 = w11366 & ~w11371;
assign w11373 = ~w11366 & w11371;
assign v5297 = ~(w11372 | w11373);
assign w11374 = v5297;
assign w11375 = w11365 & ~w11374;
assign w11376 = ~w11365 & w11374;
assign v5298 = ~(w11375 | w11376);
assign w11377 = v5298;
assign w11378 = ~w11345 & w11377;
assign w11379 = w11345 & ~w11377;
assign v5299 = ~(w11378 | w11379);
assign w11380 = v5299;
assign w11381 = ~w11344 & w11380;
assign w11382 = w11344 & ~w11380;
assign v5300 = ~(w11381 | w11382);
assign w11383 = v5300;
assign w11384 = ~w11343 & w11383;
assign w11385 = w11343 & ~w11383;
assign v5301 = ~(w11384 | w11385);
assign w11386 = v5301;
assign w11387 = ~w11342 & w11386;
assign w11388 = w11342 & ~w11386;
assign v5302 = ~(w11387 | w11388);
assign w11389 = v5302;
assign w11390 = ~w11341 & w11389;
assign w11391 = w11341 & ~w11389;
assign v5303 = ~(w11390 | w11391);
assign w11392 = v5303;
assign v5304 = ~(w11172 | w11175);
assign w11393 = v5304;
assign w11394 = (~w11198 & ~w11200) | (~w11198 & w17191) | (~w11200 & w17191);
assign w11395 = (~w11236 & ~w11238) | (~w11236 & w16772) | (~w11238 & w16772);
assign w11396 = pi18 & pi59;
assign v5305 = ~(w11299 | w11396);
assign w11397 = v5305;
assign w11398 = pi18 & pi60;
assign w11399 = w11297 & w11398;
assign v5306 = ~(w11397 | w11399);
assign w11400 = v5306;
assign w11401 = w11278 & ~w11281;
assign v5307 = ~(w11283 | w11401);
assign w11402 = v5307;
assign w11403 = w11400 & ~w11402;
assign w11404 = ~w11400 & w11402;
assign v5308 = ~(w11403 | w11404);
assign w11405 = v5308;
assign w11406 = ~w11395 & w11405;
assign w11407 = w11395 & ~w11405;
assign v5309 = ~(w11406 | w11407);
assign w11408 = v5309;
assign w11409 = w11394 & ~w11408;
assign w11410 = ~w11394 & w11408;
assign v5310 = ~(w11409 | w11410);
assign w11411 = v5310;
assign w11412 = (~w11291 & ~w11293) | (~w11291 & w17192) | (~w11293 & w17192);
assign w11413 = ~w11411 & w11412;
assign w11414 = w11411 & ~w11412;
assign v5311 = ~(w11413 | w11414);
assign w11415 = v5311;
assign w11416 = w11153 & ~w11156;
assign v5312 = ~(w11158 | w11416);
assign w11417 = v5312;
assign w11418 = w11256 & ~w11258;
assign v5313 = ~(w11260 | w11418);
assign w11419 = v5313;
assign v5314 = ~(w11417 | w11419);
assign w11420 = v5314;
assign w11421 = w11417 & w11419;
assign v5315 = ~(w11420 | w11421);
assign w11422 = v5315;
assign w11423 = w11132 & ~w11135;
assign v5316 = ~(w11137 | w11423);
assign w11424 = v5316;
assign w11425 = ~w11422 & w11424;
assign w11426 = w11422 & ~w11424;
assign v5317 = ~(w11425 | w11426);
assign w11427 = v5317;
assign w11428 = w11296 & ~w11298;
assign v5318 = ~(w11300 | w11428);
assign w11429 = v5318;
assign w11430 = w11308 & ~w11311;
assign v5319 = ~(w11313 | w11430);
assign w11431 = v5319;
assign v5320 = ~(w11429 | w11431);
assign w11432 = v5320;
assign w11433 = w11429 & w11431;
assign v5321 = ~(w11432 | w11433);
assign w11434 = v5321;
assign v5322 = ~(w11070 | w11145);
assign w11435 = v5322;
assign v5323 = ~(w11144 | w11435);
assign w11436 = v5323;
assign v5324 = ~(w11434 | w11436);
assign w11437 = v5324;
assign w11438 = w11434 & w11436;
assign v5325 = ~(w11437 | w11438);
assign w11439 = v5325;
assign w11440 = (~w11150 & ~w11152) | (~w11150 & w17829) | (~w11152 & w17829);
assign w11441 = ~w11439 & w11440;
assign w11442 = w11439 & ~w11440;
assign v5326 = ~(w11441 | w11442);
assign w11443 = v5326;
assign w11444 = w11427 & w11443;
assign v5327 = ~(w11427 | w11443);
assign w11445 = v5327;
assign v5328 = ~(w11444 | w11445);
assign w11446 = v5328;
assign w11447 = w11415 & w11446;
assign v5329 = ~(w11415 | w11446);
assign w11448 = v5329;
assign v5330 = ~(w11447 | w11448);
assign w11449 = v5330;
assign w11450 = ~w11393 & w11449;
assign w11451 = w11393 & ~w11449;
assign v5331 = ~(w11450 | w11451);
assign w11452 = v5331;
assign w11453 = (~w11275 & ~w11277) | (~w11275 & w17830) | (~w11277 & w17830);
assign w11454 = (~w11305 & ~w11307) | (~w11305 & w16941) | (~w11307 & w16941);
assign v5332 = ~(w11211 | w11214);
assign w11455 = v5332;
assign v5333 = ~(w11210 | w11455);
assign w11456 = v5333;
assign w11457 = ~w11454 & w11456;
assign w11458 = w11454 & ~w11456;
assign v5334 = ~(w11457 | w11458);
assign w11459 = v5334;
assign w11460 = w11453 & ~w11459;
assign w11461 = ~w11453 & w11459;
assign v5335 = ~(w11460 | w11461);
assign w11462 = v5335;
assign v5336 = ~(w11166 | w11169);
assign w11463 = v5336;
assign w11464 = ~w11462 & w11463;
assign w11465 = w11462 & ~w11463;
assign v5337 = ~(w11464 | w11465);
assign w11466 = v5337;
assign v5338 = ~(w11184 | w11188);
assign w11467 = v5338;
assign w11468 = pi35 & pi42;
assign w11469 = pi37 & pi40;
assign v5339 = ~(w11269 | w11469);
assign w11470 = v5339;
assign w11471 = pi37 & pi41;
assign w11472 = w11266 & w11471;
assign v5340 = ~(w11470 | w11472);
assign w11473 = v5340;
assign w11474 = w11468 & ~w11473;
assign w11475 = ~w11468 & w11473;
assign v5341 = ~(w11474 | w11475);
assign w11476 = v5341;
assign w11477 = pi14 & pi63;
assign w11478 = pi31 & pi46;
assign v5342 = ~(w11477 | w11478);
assign w11479 = v5342;
assign w11480 = w11477 & w11478;
assign v5343 = ~(w11479 | w11480);
assign w11481 = v5343;
assign w11482 = w11259 & ~w11481;
assign w11483 = ~w11259 & w11481;
assign v5344 = ~(w11482 | w11483);
assign w11484 = v5344;
assign v5345 = ~(w11476 | w11484);
assign w11485 = v5345;
assign w11486 = w11476 & w11484;
assign v5346 = ~(w11485 | w11486);
assign w11487 = v5346;
assign w11488 = pi15 & pi62;
assign w11489 = ~pi38 & pi39;
assign w11490 = w11488 & ~w11489;
assign w11491 = ~w11488 & w11489;
assign v5347 = ~(w11490 | w11491);
assign w11492 = v5347;
assign w11493 = w11487 & ~w11492;
assign w11494 = ~w11487 & w11492;
assign v5348 = ~(w11493 | w11494);
assign w11495 = v5348;
assign w11496 = ~w11467 & w11495;
assign w11497 = w11467 & ~w11495;
assign v5349 = ~(w11496 | w11497);
assign w11498 = v5349;
assign w11499 = pi19 & pi58;
assign w11500 = pi20 & pi57;
assign w11501 = pi21 & pi56;
assign v5350 = ~(w11500 | w11501);
assign w11502 = v5350;
assign w11503 = pi21 & pi57;
assign w11504 = w11153 & w11503;
assign v5351 = ~(w11502 | w11504);
assign w11505 = v5351;
assign w11506 = w11499 & ~w11505;
assign w11507 = ~w11499 & w11505;
assign v5352 = ~(w11506 | w11507);
assign w11508 = v5352;
assign w11509 = w11265 & ~w11268;
assign v5353 = ~(w11270 | w11509);
assign w11510 = v5353;
assign v5354 = ~(w11508 | w11510);
assign w11511 = v5354;
assign w11512 = w11508 & w11510;
assign v5355 = ~(w11511 | w11512);
assign w11513 = v5355;
assign w11514 = pi28 & pi49;
assign w11515 = pi29 & pi48;
assign v5356 = ~(w11514 | w11515);
assign w11516 = v5356;
assign w11517 = pi29 & pi49;
assign w11518 = w11256 & w11517;
assign v5357 = ~(w11516 | w11518);
assign w11519 = v5357;
assign w11520 = w11312 & ~w11519;
assign w11521 = ~w11312 & w11519;
assign v5358 = ~(w11520 | w11521);
assign w11522 = v5358;
assign w11523 = w11513 & ~w11522;
assign w11524 = ~w11513 & w11522;
assign v5359 = ~(w11523 | w11524);
assign w11525 = v5359;
assign w11526 = w11498 & w11525;
assign v5360 = ~(w11498 | w11525);
assign w11527 = v5360;
assign v5361 = ~(w11526 | w11527);
assign w11528 = v5361;
assign w11529 = w11466 & w11528;
assign v5362 = ~(w11466 | w11528);
assign w11530 = v5362;
assign v5363 = ~(w11529 | w11530);
assign w11531 = v5363;
assign w11532 = w11452 & w11531;
assign v5364 = ~(w11452 | w11531);
assign w11533 = v5364;
assign v5365 = ~(w11532 | w11533);
assign w11534 = v5365;
assign w11535 = w11392 & w11534;
assign v5366 = ~(w11392 | w11534);
assign w11536 = v5366;
assign v5367 = ~(w11535 | w11536);
assign w11537 = v5367;
assign w11538 = ~w11340 & w11537;
assign w11539 = w11340 & ~w11537;
assign v5368 = ~(w11538 | w11539);
assign w11540 = v5368;
assign v5369 = ~(w11119 | w11334);
assign w11541 = v5369;
assign w11542 = (~w7754 & w17831) | (~w7754 & w17832) | (w17831 & w17832);
assign w11543 = w11540 & w11542;
assign v5370 = ~(w11540 | w11542);
assign w11544 = v5370;
assign v5371 = ~(w11543 | w11544);
assign w11545 = v5371;
assign v5372 = ~(w11333 | w11538);
assign w11546 = v5372;
assign w11547 = (w8795 & w17628) | (w8795 & w17629) | (w17628 & w17629);
assign v5373 = ~(w11390 | w11535);
assign w11548 = v5373;
assign v5374 = ~(w11465 | w11529);
assign w11549 = v5374;
assign v5375 = ~(w11414 | w11447);
assign w11550 = v5375;
assign w11551 = (~w11457 & ~w11459) | (~w11457 & w17193) | (~w11459 & w17193);
assign w11552 = pi27 & pi51;
assign w11553 = pi28 & pi50;
assign v5376 = ~(w11517 | w11553);
assign w11554 = v5376;
assign w11555 = pi29 & pi50;
assign w11556 = w11514 & w11555;
assign v5377 = ~(w11554 | w11556);
assign w11557 = v5377;
assign w11558 = w11552 & ~w11557;
assign w11559 = ~w11552 & w11557;
assign v5378 = ~(w11558 | w11559);
assign w11560 = v5378;
assign w11561 = pi19 & pi59;
assign v5379 = ~(w11503 | w11561);
assign w11562 = v5379;
assign w11563 = w11503 & w11561;
assign v5380 = ~(w11562 | w11563);
assign w11564 = v5380;
assign w11565 = w11398 & ~w11564;
assign w11566 = ~w11398 & w11564;
assign v5381 = ~(w11565 | w11566);
assign w11567 = v5381;
assign v5382 = ~(w11560 | w11567);
assign w11568 = v5382;
assign w11569 = w11560 & w11567;
assign v5383 = ~(w11568 | w11569);
assign w11570 = v5383;
assign w11571 = pi15 & pi63;
assign w11572 = pi16 & pi62;
assign w11573 = pi17 & pi61;
assign v5384 = ~(w11572 | w11573);
assign w11574 = v5384;
assign w11575 = pi17 & pi62;
assign w11576 = w11366 & w11575;
assign v5385 = ~(w11574 | w11576);
assign w11577 = v5385;
assign w11578 = w11571 & ~w11577;
assign w11579 = ~w11571 & w11577;
assign v5386 = ~(w11578 | w11579);
assign w11580 = v5386;
assign w11581 = w11570 & ~w11580;
assign w11582 = ~w11570 & w11580;
assign v5387 = ~(w11581 | w11582);
assign w11583 = v5387;
assign w11584 = pi32 & pi46;
assign w11585 = pi34 & pi44;
assign v5388 = ~(w11369 | w11585);
assign w11586 = v5388;
assign w11587 = pi34 & pi45;
assign w11588 = w11367 & w11587;
assign v5389 = ~(w11586 | w11588);
assign w11589 = v5389;
assign w11590 = w11584 & ~w11589;
assign w11591 = ~w11584 & w11589;
assign v5390 = ~(w11590 | w11591);
assign w11592 = v5390;
assign w11593 = pi20 & pi58;
assign w11594 = pi31 & pi47;
assign w11595 = pi30 & pi48;
assign v5391 = ~(w11594 | w11595);
assign w11596 = v5391;
assign w11597 = pi31 & pi48;
assign w11598 = w11259 & w11597;
assign v5392 = ~(w11596 | w11598);
assign w11599 = v5392;
assign w11600 = w11593 & ~w11599;
assign w11601 = ~w11593 & w11599;
assign v5393 = ~(w11600 | w11601);
assign w11602 = v5393;
assign v5394 = ~(w11592 | w11602);
assign w11603 = v5394;
assign w11604 = w11592 & w11602;
assign v5395 = ~(w11603 | w11604);
assign w11605 = v5395;
assign w11606 = pi25 & pi53;
assign w11607 = pi22 & pi56;
assign v5396 = ~(w11349 | w11607);
assign w11608 = v5396;
assign w11609 = w11349 & w11607;
assign v5397 = ~(w11608 | w11609);
assign w11610 = v5397;
assign w11611 = w11606 & ~w11610;
assign w11612 = ~w11606 & w11610;
assign v5398 = ~(w11611 | w11612);
assign w11613 = v5398;
assign w11614 = w11605 & ~w11613;
assign w11615 = ~w11605 & w11613;
assign v5399 = ~(w11614 | w11615);
assign w11616 = v5399;
assign w11617 = w11583 & w11616;
assign v5400 = ~(w11583 | w11616);
assign w11618 = v5400;
assign v5401 = ~(w11617 | w11618);
assign w11619 = v5401;
assign w11620 = ~w11551 & w11619;
assign w11621 = w11551 & ~w11619;
assign v5402 = ~(w11620 | w11621);
assign w11622 = v5402;
assign w11623 = ~w11550 & w11622;
assign w11624 = w11550 & ~w11622;
assign v5403 = ~(w11623 | w11624);
assign w11625 = v5403;
assign w11626 = w11549 & ~w11625;
assign w11627 = ~w11549 & w11625;
assign v5404 = ~(w11626 | w11627);
assign w11628 = v5404;
assign v5405 = ~(w11450 | w11532);
assign w11629 = v5405;
assign w11630 = ~w11628 & w11629;
assign w11631 = w11628 & ~w11629;
assign v5406 = ~(w11630 | w11631);
assign w11632 = v5406;
assign v5407 = ~(w11384 | w11387);
assign w11633 = v5407;
assign w11634 = (~w11363 & ~w11365) | (~w11363 & w17833) | (~w11365 & w17833);
assign w11635 = (~w11511 & ~w11513) | (~w11511 & w16942) | (~w11513 & w16942);
assign w11636 = (~w11485 & ~w11487) | (~w11485 & w16943) | (~w11487 & w16943);
assign v5408 = ~(w11635 | w11636);
assign w11637 = v5408;
assign w11638 = w11635 & w11636;
assign v5409 = ~(w11637 | w11638);
assign w11639 = v5409;
assign w11640 = w11634 & ~w11639;
assign w11641 = ~w11634 & w11639;
assign v5410 = ~(w11640 | w11641);
assign w11642 = v5410;
assign v5411 = ~(w11442 | w11444);
assign w11643 = v5411;
assign w11644 = ~w11642 & w11643;
assign w11645 = w11642 & ~w11643;
assign v5412 = ~(w11644 | w11645);
assign w11646 = v5412;
assign v5413 = ~(pi38 | w11488);
assign w11647 = v5413;
assign w11648 = pi39 & ~w11647;
assign w11649 = w11468 & ~w11470;
assign v5414 = ~(w11472 | w11649);
assign w11650 = v5414;
assign w11651 = w11648 & ~w11650;
assign w11652 = ~w11648 & w11650;
assign v5415 = ~(w11651 | w11652);
assign w11653 = v5415;
assign w11654 = w11282 & ~w11348;
assign v5416 = ~(w11350 | w11654);
assign w11655 = v5416;
assign w11656 = ~w11653 & w11655;
assign w11657 = w11653 & ~w11655;
assign v5417 = ~(w11656 | w11657);
assign w11658 = v5417;
assign v5418 = ~(w11259 | w11480);
assign w11659 = v5418;
assign v5419 = ~(w11479 | w11659);
assign w11660 = v5419;
assign w11661 = w11312 & ~w11516;
assign v5420 = ~(w11518 | w11661);
assign w11662 = v5420;
assign w11663 = w11660 & ~w11662;
assign w11664 = ~w11660 & w11662;
assign v5421 = ~(w11663 | w11664);
assign w11665 = v5421;
assign w11666 = w11366 & ~w11368;
assign v5422 = ~(w11370 | w11666);
assign w11667 = v5422;
assign w11668 = ~w11665 & w11667;
assign w11669 = w11665 & ~w11667;
assign v5423 = ~(w11668 | w11669);
assign w11670 = v5423;
assign w11671 = (~w11432 & ~w11434) | (~w11432 & w17194) | (~w11434 & w17194);
assign w11672 = ~w11670 & w11671;
assign w11673 = w11670 & ~w11671;
assign v5424 = ~(w11672 | w11673);
assign w11674 = v5424;
assign w11675 = w11658 & w11674;
assign v5425 = ~(w11658 | w11674);
assign w11676 = v5425;
assign v5426 = ~(w11675 | w11676);
assign w11677 = v5426;
assign w11678 = w11646 & w11677;
assign v5427 = ~(w11646 | w11677);
assign w11679 = v5427;
assign v5428 = ~(w11678 | w11679);
assign w11680 = v5428;
assign w11681 = ~w11633 & w11680;
assign w11682 = w11633 & ~w11680;
assign v5429 = ~(w11681 | w11682);
assign w11683 = v5429;
assign w11684 = (~w11420 & ~w11422) | (~w11420 & w16773) | (~w11422 & w16773);
assign w11685 = pi23 & pi55;
assign w11686 = pi35 & pi43;
assign w11687 = pi36 & pi42;
assign v5430 = ~(w11686 | w11687);
assign w11688 = v5430;
assign w11689 = pi36 & pi43;
assign w11690 = w11468 & w11689;
assign v5431 = ~(w11688 | w11690);
assign w11691 = v5431;
assign w11692 = w11685 & ~w11691;
assign w11693 = ~w11685 & w11691;
assign v5432 = ~(w11692 | w11693);
assign w11694 = v5432;
assign w11695 = pi38 & pi40;
assign w11696 = pi26 & pi52;
assign v5433 = ~(w11695 | w11696);
assign w11697 = v5433;
assign w11698 = w11695 & w11696;
assign v5434 = ~(w11697 | w11698);
assign w11699 = v5434;
assign w11700 = w11471 & ~w11699;
assign w11701 = ~w11471 & w11699;
assign v5435 = ~(w11700 | w11701);
assign w11702 = v5435;
assign v5436 = ~(w11694 | w11702);
assign w11703 = v5436;
assign w11704 = w11694 & w11702;
assign v5437 = ~(w11703 | w11704);
assign w11705 = v5437;
assign w11706 = w11684 & ~w11705;
assign w11707 = ~w11684 & w11705;
assign v5438 = ~(w11706 | w11707);
assign w11708 = v5438;
assign w11709 = (~w11399 & w11402) | (~w11399 & w16944) | (w11402 & w16944);
assign v5439 = ~(w11355 | w11358);
assign w11710 = v5439;
assign v5440 = ~(w11357 | w11710);
assign w11711 = v5440;
assign w11712 = w11499 & ~w11502;
assign v5441 = ~(w11504 | w11712);
assign w11713 = v5441;
assign w11714 = w11711 & ~w11713;
assign w11715 = ~w11711 & w11713;
assign v5442 = ~(w11714 | w11715);
assign w11716 = v5442;
assign w11717 = w11709 & ~w11716;
assign w11718 = ~w11709 & w11716;
assign v5443 = ~(w11717 | w11718);
assign w11719 = v5443;
assign w11720 = (~w11406 & ~w11408) | (~w11406 & w16945) | (~w11408 & w16945);
assign w11721 = ~w11719 & w11720;
assign w11722 = w11719 & ~w11720;
assign v5444 = ~(w11721 | w11722);
assign w11723 = v5444;
assign w11724 = w11708 & w11723;
assign v5445 = ~(w11708 | w11723);
assign w11725 = v5445;
assign v5446 = ~(w11724 | w11725);
assign w11726 = v5446;
assign v5447 = ~(w11378 | w11381);
assign w11727 = v5447;
assign v5448 = ~(w11496 | w11526);
assign w11728 = v5448;
assign v5449 = ~(w11727 | w11728);
assign w11729 = v5449;
assign w11730 = w11727 & w11728;
assign v5450 = ~(w11729 | w11730);
assign w11731 = v5450;
assign w11732 = w11726 & w11731;
assign v5451 = ~(w11726 | w11731);
assign w11733 = v5451;
assign v5452 = ~(w11732 | w11733);
assign w11734 = v5452;
assign w11735 = w11683 & w11734;
assign v5453 = ~(w11683 | w11734);
assign w11736 = v5453;
assign v5454 = ~(w11735 | w11736);
assign w11737 = v5454;
assign w11738 = w11632 & w11737;
assign v5455 = ~(w11632 | w11737);
assign w11739 = v5455;
assign v5456 = ~(w11738 | w11739);
assign w11740 = v5456;
assign w11741 = ~w11548 & w11740;
assign w11742 = w11548 & ~w11740;
assign v5457 = ~(w11741 | w11742);
assign w11743 = v5457;
assign w11744 = w11547 & ~w11743;
assign w11745 = ~w11547 & w11743;
assign v5458 = ~(w11744 | w11745);
assign w11746 = v5458;
assign v5459 = ~(w11631 | w11738);
assign w11747 = v5459;
assign v5460 = ~(w11729 | w11732);
assign w11748 = v5460;
assign v5461 = ~(w11617 | w11620);
assign w11749 = v5461;
assign v5462 = ~(w11398 | w11563);
assign w11750 = v5462;
assign v5463 = ~(w11562 | w11750);
assign w11751 = v5463;
assign w11752 = w11552 & ~w11554;
assign v5464 = ~(w11556 | w11752);
assign w11753 = v5464;
assign w11754 = w11751 & ~w11753;
assign w11755 = ~w11751 & w11753;
assign v5465 = ~(w11754 | w11755);
assign w11756 = v5465;
assign v5466 = ~(w11606 | w11609);
assign w11757 = v5466;
assign v5467 = ~(w11608 | w11757);
assign w11758 = v5467;
assign v5468 = ~(w11756 | w11758);
assign w11759 = v5468;
assign w11760 = w11756 & w11758;
assign v5469 = ~(w11759 | w11760);
assign w11761 = v5469;
assign v5470 = ~(w11703 | w11707);
assign w11762 = v5470;
assign w11763 = ~w11761 & w11762;
assign w11764 = w11761 & ~w11762;
assign v5471 = ~(w11763 | w11764);
assign w11765 = v5471;
assign w11766 = (~w11714 & ~w11716) | (~w11714 & w16946) | (~w11716 & w16946);
assign w11767 = pi16 & pi63;
assign w11768 = pi35 & pi44;
assign v5472 = ~(w11587 | w11768);
assign w11769 = v5472;
assign w11770 = pi35 & pi45;
assign w11771 = w11585 & w11770;
assign v5473 = ~(w11769 | w11771);
assign w11772 = v5473;
assign w11773 = w11767 & ~w11772;
assign w11774 = ~w11767 & w11772;
assign v5474 = ~(w11773 | w11774);
assign w11775 = v5474;
assign w11776 = pi23 & pi56;
assign w11777 = pi27 & pi52;
assign v5475 = ~(w11776 | w11777);
assign w11778 = v5475;
assign w11779 = w11776 & w11777;
assign v5476 = ~(w11778 | w11779);
assign w11780 = v5476;
assign w11781 = w11689 & ~w11780;
assign w11782 = ~w11689 & w11780;
assign v5477 = ~(w11781 | w11782);
assign w11783 = v5477;
assign v5478 = ~(w11775 | w11783);
assign w11784 = v5478;
assign w11785 = w11775 & w11783;
assign v5479 = ~(w11784 | w11785);
assign w11786 = v5479;
assign w11787 = w11766 & ~w11786;
assign w11788 = ~w11766 & w11786;
assign v5480 = ~(w11787 | w11788);
assign w11789 = v5480;
assign w11790 = w11765 & w11789;
assign v5481 = ~(w11765 | w11789);
assign w11791 = v5481;
assign v5482 = ~(w11790 | w11791);
assign w11792 = v5482;
assign w11793 = ~w11749 & w11792;
assign w11794 = w11749 & ~w11792;
assign v5483 = ~(w11793 | w11794);
assign w11795 = v5483;
assign v5484 = ~(w11603 | w11614);
assign w11796 = v5484;
assign w11797 = pi18 & pi61;
assign v5485 = ~(w11471 | w11698);
assign w11798 = v5485;
assign w11799 = ~w11798 & w17195;
assign w11800 = (~w11797 & w11798) | (~w11797 & w17196) | (w11798 & w17196);
assign v5486 = ~(w11799 | w11800);
assign w11801 = v5486;
assign w11802 = w11685 & ~w11688;
assign v5487 = ~(w11690 | w11802);
assign w11803 = v5487;
assign w11804 = ~w11801 & w11803;
assign w11805 = w11801 & ~w11803;
assign v5488 = ~(w11804 | w11805);
assign w11806 = v5488;
assign w11807 = w11571 & ~w11574;
assign v5489 = ~(w11576 | w11807);
assign w11808 = v5489;
assign w11809 = w11593 & ~w11596;
assign v5490 = ~(w11598 | w11809);
assign w11810 = v5490;
assign v5491 = ~(w11808 | w11810);
assign w11811 = v5491;
assign w11812 = w11808 & w11810;
assign v5492 = ~(w11811 | w11812);
assign w11813 = v5492;
assign w11814 = w11584 & ~w11586;
assign v5493 = ~(w11588 | w11814);
assign w11815 = v5493;
assign w11816 = ~w11813 & w11815;
assign w11817 = w11813 & ~w11815;
assign v5494 = ~(w11816 | w11817);
assign w11818 = v5494;
assign w11819 = w11806 & w11818;
assign v5495 = ~(w11806 | w11818);
assign w11820 = v5495;
assign v5496 = ~(w11819 | w11820);
assign w11821 = v5496;
assign w11822 = ~w11796 & w11821;
assign w11823 = w11796 & ~w11821;
assign v5497 = ~(w11822 | w11823);
assign w11824 = v5497;
assign w11825 = w11795 & w11824;
assign v5498 = ~(w11795 | w11824);
assign w11826 = v5498;
assign v5499 = ~(w11825 | w11826);
assign w11827 = v5499;
assign w11828 = ~w11748 & w11827;
assign w11829 = w11748 & ~w11827;
assign v5500 = ~(w11828 | w11829);
assign w11830 = v5500;
assign v5501 = ~(w11623 | w11627);
assign w11831 = v5501;
assign w11832 = ~w11830 & w11831;
assign w11833 = w11830 & ~w11831;
assign v5502 = ~(w11832 | w11833);
assign w11834 = v5502;
assign v5503 = ~(w11645 | w11678);
assign w11835 = v5503;
assign w11836 = (~w11673 & ~w11674) | (~w11673 & w17197) | (~w11674 & w17197);
assign w11837 = pi24 & pi55;
assign w11838 = pi26 & pi53;
assign w11839 = pi25 & pi54;
assign v5504 = ~(w11838 | w11839);
assign w11840 = v5504;
assign w11841 = pi26 & pi54;
assign w11842 = w11606 & w11841;
assign v5505 = ~(w11840 | w11842);
assign w11843 = v5505;
assign w11844 = w11837 & ~w11843;
assign w11845 = ~w11837 & w11843;
assign v5506 = ~(w11844 | w11845);
assign w11846 = v5506;
assign w11847 = pi37 & pi42;
assign w11848 = pi39 & pi40;
assign w11849 = pi38 & pi41;
assign v5507 = ~(w11848 | w11849);
assign w11850 = v5507;
assign w11851 = pi39 & pi41;
assign w11852 = w11695 & w11851;
assign v5508 = ~(w11850 | w11852);
assign w11853 = v5508;
assign w11854 = w11847 & ~w11853;
assign w11855 = ~w11847 & w11853;
assign v5509 = ~(w11854 | w11855);
assign w11856 = v5509;
assign v5510 = ~(w11846 | w11856);
assign w11857 = v5510;
assign w11858 = w11846 & w11856;
assign v5511 = ~(w11857 | w11858);
assign w11859 = v5511;
assign w11860 = pi28 & pi51;
assign v5512 = ~(pi40 | w11575);
assign w11861 = v5512;
assign w11862 = pi62 & w6702;
assign v5513 = ~(w11861 | w11862);
assign w11863 = v5513;
assign w11864 = w11860 & ~w11863;
assign w11865 = ~w11860 & w11863;
assign v5514 = ~(w11864 | w11865);
assign w11866 = v5514;
assign w11867 = w11859 & ~w11866;
assign w11868 = ~w11859 & w11866;
assign v5515 = ~(w11867 | w11868);
assign w11869 = v5515;
assign w11870 = pi19 & pi60;
assign w11871 = pi20 & pi59;
assign w11872 = pi21 & pi58;
assign v5516 = ~(w11871 | w11872);
assign w11873 = v5516;
assign w11874 = pi21 & pi59;
assign w11875 = w11593 & w11874;
assign v5517 = ~(w11873 | w11875);
assign w11876 = v5517;
assign w11877 = w11870 & ~w11876;
assign w11878 = ~w11870 & w11876;
assign v5518 = ~(w11877 | w11878);
assign w11879 = v5518;
assign w11880 = pi22 & pi57;
assign w11881 = pi30 & pi49;
assign v5519 = ~(w11555 | w11881);
assign w11882 = v5519;
assign w11883 = pi30 & pi50;
assign w11884 = w11517 & w11883;
assign v5520 = ~(w11882 | w11884);
assign w11885 = v5520;
assign w11886 = w11880 & ~w11885;
assign w11887 = ~w11880 & w11885;
assign v5521 = ~(w11886 | w11887);
assign w11888 = v5521;
assign v5522 = ~(w11879 | w11888);
assign w11889 = v5522;
assign w11890 = w11879 & w11888;
assign v5523 = ~(w11889 | w11890);
assign w11891 = v5523;
assign w11892 = pi33 & pi46;
assign w11893 = pi32 & pi47;
assign v5524 = ~(w11892 | w11893);
assign w11894 = v5524;
assign w11895 = pi33 & pi47;
assign w11896 = w11584 & w11895;
assign v5525 = ~(w11894 | w11896);
assign w11897 = v5525;
assign w11898 = w11597 & ~w11897;
assign w11899 = ~w11597 & w11897;
assign v5526 = ~(w11898 | w11899);
assign w11900 = v5526;
assign w11901 = w11891 & ~w11900;
assign w11902 = ~w11891 & w11900;
assign v5527 = ~(w11901 | w11902);
assign w11903 = v5527;
assign w11904 = w11869 & w11903;
assign v5528 = ~(w11869 | w11903);
assign w11905 = v5528;
assign v5529 = ~(w11904 | w11905);
assign w11906 = v5529;
assign w11907 = ~w11836 & w11906;
assign w11908 = w11836 & ~w11906;
assign v5530 = ~(w11907 | w11908);
assign w11909 = v5530;
assign w11910 = ~w11835 & w11909;
assign w11911 = w11835 & ~w11909;
assign v5531 = ~(w11910 | w11911);
assign w11912 = v5531;
assign w11913 = (~w11568 & ~w11570) | (~w11568 & w17198) | (~w11570 & w17198);
assign w11914 = (~w11663 & ~w11665) | (~w11663 & w16947) | (~w11665 & w16947);
assign w11915 = (~w11651 & ~w11653) | (~w11651 & w16948) | (~w11653 & w16948);
assign v5532 = ~(w11914 | w11915);
assign w11916 = v5532;
assign w11917 = w11914 & w11915;
assign v5533 = ~(w11916 | w11917);
assign w11918 = v5533;
assign w11919 = w11913 & ~w11918;
assign w11920 = ~w11913 & w11918;
assign v5534 = ~(w11919 | w11920);
assign w11921 = v5534;
assign w11922 = (~w11637 & ~w11639) | (~w11637 & w17199) | (~w11639 & w17199);
assign w11923 = ~w11921 & w11922;
assign w11924 = w11921 & ~w11922;
assign v5535 = ~(w11923 | w11924);
assign w11925 = v5535;
assign w11926 = (~w11722 & ~w11723) | (~w11722 & w17200) | (~w11723 & w17200);
assign w11927 = w11925 & ~w11926;
assign w11928 = ~w11925 & w11926;
assign v5536 = ~(w11927 | w11928);
assign w11929 = v5536;
assign w11930 = w11912 & w11929;
assign v5537 = ~(w11912 | w11929);
assign w11931 = v5537;
assign v5538 = ~(w11930 | w11931);
assign w11932 = v5538;
assign v5539 = ~(w11681 | w11735);
assign w11933 = v5539;
assign w11934 = w11932 & ~w11933;
assign w11935 = ~w11932 & w11933;
assign v5540 = ~(w11934 | w11935);
assign w11936 = v5540;
assign w11937 = w11834 & w11936;
assign v5541 = ~(w11834 | w11936);
assign w11938 = v5541;
assign v5542 = ~(w11937 | w11938);
assign w11939 = v5542;
assign w11940 = ~w11747 & w11939;
assign w11941 = w11747 & ~w11939;
assign v5543 = ~(w11940 | w11941);
assign w11942 = v5543;
assign w11943 = (w7754 & w17834) | (w7754 & w17835) | (w17834 & w17835);
assign w11944 = w11942 & w11943;
assign v5544 = ~(w11942 | w11943);
assign w11945 = v5544;
assign v5545 = ~(w11944 | w11945);
assign w11946 = v5545;
assign v5546 = ~(w11742 | w11941);
assign w11947 = v5546;
assign w11948 = (~w7754 & w17836) | (~w7754 & w17837) | (w17836 & w17837);
assign v5547 = ~(w11934 | w11937);
assign w11949 = v5547;
assign v5548 = ~(w11828 | w11833);
assign w11950 = v5548;
assign w11951 = (~w11793 & ~w11795) | (~w11793 & w17838) | (~w11795 & w17838);
assign w11952 = pi19 & pi61;
assign w11953 = pi18 & pi62;
assign v5549 = ~(w11952 | w11953);
assign w11954 = v5549;
assign w11955 = pi19 & pi62;
assign w11956 = w11797 & w11955;
assign v5550 = ~(w11954 | w11956);
assign w11957 = v5550;
assign v5551 = ~(w11860 | w11862);
assign w11958 = v5551;
assign v5552 = ~(w11861 | w11958);
assign w11959 = v5552;
assign w11960 = w11957 & w11959;
assign v5553 = ~(w11957 | w11959);
assign w11961 = v5553;
assign v5554 = ~(w11960 | w11961);
assign w11962 = v5554;
assign w11963 = pi34 & pi46;
assign w11964 = pi36 & pi44;
assign v5555 = ~(w11770 | w11964);
assign w11965 = v5555;
assign w11966 = pi36 & pi45;
assign w11967 = w11768 & w11966;
assign v5556 = ~(w11965 | w11967);
assign w11968 = v5556;
assign w11969 = w11963 & ~w11968;
assign w11970 = ~w11963 & w11968;
assign v5557 = ~(w11969 | w11970);
assign w11971 = v5557;
assign w11972 = pi17 & pi63;
assign w11973 = pi29 & pi51;
assign v5558 = ~(w11972 | w11973);
assign w11974 = v5558;
assign w11975 = w11972 & w11973;
assign v5559 = ~(w11974 | w11975);
assign w11976 = v5559;
assign w11977 = w11895 & ~w11976;
assign w11978 = ~w11895 & w11976;
assign v5560 = ~(w11977 | w11978);
assign w11979 = v5560;
assign v5561 = ~(w11971 | w11979);
assign w11980 = v5561;
assign w11981 = w11971 & w11979;
assign v5562 = ~(w11980 | w11981);
assign w11982 = v5562;
assign w11983 = w11962 & w11982;
assign v5563 = ~(w11962 | w11982);
assign w11984 = v5563;
assign v5564 = ~(w11983 | w11984);
assign w11985 = v5564;
assign w11986 = pi20 & pi60;
assign w11987 = pi22 & pi58;
assign v5565 = ~(w11874 | w11987);
assign w11988 = v5565;
assign w11989 = pi22 & pi59;
assign w11990 = w11872 & w11989;
assign v5566 = ~(w11988 | w11990);
assign w11991 = v5566;
assign w11992 = w11986 & ~w11991;
assign w11993 = ~w11986 & w11991;
assign v5567 = ~(w11992 | w11993);
assign w11994 = v5567;
assign w11995 = w11847 & ~w11850;
assign v5568 = ~(w11852 | w11995);
assign w11996 = v5568;
assign v5569 = ~(w11994 | w11996);
assign w11997 = v5569;
assign w11998 = w11994 & w11996;
assign v5570 = ~(w11997 | w11998);
assign w11999 = v5570;
assign w12000 = pi31 & pi49;
assign w12001 = pi32 & pi48;
assign v5571 = ~(w12000 | w12001);
assign w12002 = v5571;
assign w12003 = pi32 & pi49;
assign w12004 = w11597 & w12003;
assign v5572 = ~(w12002 | w12004);
assign w12005 = v5572;
assign w12006 = w11883 & ~w12005;
assign w12007 = ~w11883 & w12005;
assign v5573 = ~(w12006 | w12007);
assign w12008 = v5573;
assign w12009 = ~w11999 & w12008;
assign w12010 = w11999 & ~w12008;
assign v5574 = ~(w12009 | w12010);
assign w12011 = v5574;
assign w12012 = pi25 & pi55;
assign w12013 = pi38 & pi42;
assign w12014 = pi37 & pi43;
assign v5575 = ~(w12013 | w12014);
assign w12015 = v5575;
assign w12016 = pi38 & pi43;
assign w12017 = w11847 & w12016;
assign v5576 = ~(w12015 | w12017);
assign w12018 = v5576;
assign w12019 = w12012 & ~w12018;
assign w12020 = ~w12012 & w12018;
assign v5577 = ~(w12019 | w12020);
assign w12021 = v5577;
assign w12022 = pi23 & pi57;
assign w12023 = pi24 & pi56;
assign v5578 = ~(w11841 | w12023);
assign w12024 = v5578;
assign w12025 = w11841 & w12023;
assign v5579 = ~(w12024 | w12025);
assign w12026 = v5579;
assign w12027 = w12022 & ~w12026;
assign w12028 = ~w12022 & w12026;
assign v5580 = ~(w12027 | w12028);
assign w12029 = v5580;
assign v5581 = ~(w12021 | w12029);
assign w12030 = v5581;
assign w12031 = w12021 & w12029;
assign v5582 = ~(w12030 | w12031);
assign w12032 = v5582;
assign w12033 = pi28 & pi52;
assign w12034 = pi27 & pi53;
assign v5583 = ~(w12033 | w12034);
assign w12035 = v5583;
assign w12036 = pi28 & pi53;
assign w12037 = w11777 & w12036;
assign v5584 = ~(w12035 | w12037);
assign w12038 = v5584;
assign w12039 = w11851 & ~w12038;
assign w12040 = ~w11851 & w12038;
assign v5585 = ~(w12039 | w12040);
assign w12041 = v5585;
assign w12042 = w12032 & ~w12041;
assign w12043 = ~w12032 & w12041;
assign v5586 = ~(w12042 | w12043);
assign w12044 = v5586;
assign w12045 = w12011 & w12044;
assign v5587 = ~(w12011 | w12044);
assign w12046 = v5587;
assign v5588 = ~(w12045 | w12046);
assign w12047 = v5588;
assign w12048 = w11985 & w12047;
assign v5589 = ~(w11985 | w12047);
assign w12049 = v5589;
assign v5590 = ~(w12048 | w12049);
assign w12050 = v5590;
assign w12051 = (w12050 & w11927) | (w12050 & w17839) | (w11927 & w17839);
assign w12052 = ~w11927 & w17840;
assign v5591 = ~(w12051 | w12052);
assign w12053 = v5591;
assign w12054 = ~w11951 & w12053;
assign w12055 = w11951 & ~w12053;
assign v5592 = ~(w12054 | w12055);
assign w12056 = v5592;
assign w12057 = ~w11950 & w12056;
assign w12058 = w11950 & ~w12056;
assign v5593 = ~(w12057 | w12058);
assign w12059 = v5593;
assign v5594 = ~(w11910 | w11930);
assign w12060 = v5594;
assign v5595 = ~(w11904 | w11907);
assign w12061 = v5595;
assign w12062 = w11767 & ~w11769;
assign v5596 = ~(w11771 | w12062);
assign w12063 = v5596;
assign w12064 = w11837 & ~w11840;
assign v5597 = ~(w11842 | w12064);
assign w12065 = v5597;
assign v5598 = ~(w12063 | w12065);
assign w12066 = v5598;
assign w12067 = w12063 & w12065;
assign v5599 = ~(w12066 | w12067);
assign w12068 = v5599;
assign v5600 = ~(w11689 | w11779);
assign w12069 = v5600;
assign v5601 = ~(w11778 | w12069);
assign w12070 = v5601;
assign v5602 = ~(w12068 | w12070);
assign w12071 = v5602;
assign w12072 = w12068 & w12070;
assign v5603 = ~(w12071 | w12072);
assign w12073 = v5603;
assign v5604 = ~(w11784 | w11788);
assign w12074 = v5604;
assign w12075 = ~w12073 & w12074;
assign w12076 = w12073 & ~w12074;
assign v5605 = ~(w12075 | w12076);
assign w12077 = v5605;
assign w12078 = (~w11916 & ~w11918) | (~w11916 & w17201) | (~w11918 & w17201);
assign w12079 = ~w12077 & w12078;
assign w12080 = w12077 & ~w12078;
assign v5606 = ~(w12079 | w12080);
assign w12081 = v5606;
assign w12082 = ~w12061 & w12081;
assign w12083 = w12061 & ~w12081;
assign v5607 = ~(w12082 | w12083);
assign w12084 = v5607;
assign w12085 = w11870 & ~w11873;
assign v5608 = ~(w11875 | w12085);
assign w12086 = v5608;
assign w12087 = w11880 & ~w11882;
assign v5609 = ~(w11884 | w12087);
assign w12088 = v5609;
assign v5610 = ~(w12086 | w12088);
assign w12089 = v5610;
assign w12090 = w12086 & w12088;
assign v5611 = ~(w12089 | w12090);
assign w12091 = v5611;
assign w12092 = w11597 & ~w11894;
assign v5612 = ~(w11896 | w12092);
assign w12093 = v5612;
assign w12094 = ~w12091 & w12093;
assign w12095 = w12091 & ~w12093;
assign v5613 = ~(w12094 | w12095);
assign w12096 = v5613;
assign w12097 = (~w11857 & ~w11859) | (~w11857 & w17202) | (~w11859 & w17202);
assign w12098 = (~w11889 & ~w11891) | (~w11889 & w17203) | (~w11891 & w17203);
assign v5614 = ~(w12097 | w12098);
assign w12099 = v5614;
assign w12100 = w12097 & w12098;
assign v5615 = ~(w12099 | w12100);
assign w12101 = v5615;
assign w12102 = w12096 & w12101;
assign v5616 = ~(w12096 | w12101);
assign w12103 = v5616;
assign v5617 = ~(w12102 | w12103);
assign w12104 = v5617;
assign w12105 = w12084 & w12104;
assign v5618 = ~(w12084 | w12104);
assign w12106 = v5618;
assign v5619 = ~(w12105 | w12106);
assign w12107 = v5619;
assign v5620 = ~(w11799 | w11805);
assign w12108 = v5620;
assign w12109 = (~w11754 & ~w11756) | (~w11754 & w17204) | (~w11756 & w17204);
assign w12110 = (~w11811 & ~w11813) | (~w11811 & w17205) | (~w11813 & w17205);
assign v5621 = ~(w12109 | w12110);
assign w12111 = v5621;
assign w12112 = w12109 & w12110;
assign v5622 = ~(w12111 | w12112);
assign w12113 = v5622;
assign w12114 = w12108 & ~w12113;
assign w12115 = ~w12108 & w12113;
assign v5623 = ~(w12114 | w12115);
assign w12116 = v5623;
assign w12117 = (~w11764 & ~w11765) | (~w11764 & w16949) | (~w11765 & w16949);
assign w12118 = (~w11819 & ~w11821) | (~w11819 & w17206) | (~w11821 & w17206);
assign v5624 = ~(w12117 | w12118);
assign w12119 = v5624;
assign w12120 = w12117 & w12118;
assign v5625 = ~(w12119 | w12120);
assign w12121 = v5625;
assign v5626 = ~(w12116 | w12121);
assign w12122 = v5626;
assign w12123 = w12116 & w12121;
assign v5627 = ~(w12122 | w12123);
assign w12124 = v5627;
assign w12125 = w12107 & w12124;
assign v5628 = ~(w12107 | w12124);
assign w12126 = v5628;
assign v5629 = ~(w12125 | w12126);
assign w12127 = v5629;
assign w12128 = ~w12060 & w12127;
assign w12129 = w12060 & ~w12127;
assign v5630 = ~(w12128 | w12129);
assign w12130 = v5630;
assign w12131 = w12059 & w12130;
assign v5631 = ~(w12059 | w12130);
assign w12132 = v5631;
assign v5632 = ~(w12131 | w12132);
assign w12133 = v5632;
assign w12134 = ~w11949 & w12133;
assign w12135 = w11949 & ~w12133;
assign v5633 = ~(w12134 | w12135);
assign w12136 = v5633;
assign w12137 = w11948 & w12136;
assign v5634 = ~(w11948 | w12136);
assign w12138 = v5634;
assign v5635 = ~(w12137 | w12138);
assign w12139 = v5635;
assign v5636 = ~(w11940 | w12134);
assign w12140 = v5636;
assign w12141 = (w8795 & w17630) | (w8795 & w17631) | (w17630 & w17631);
assign v5637 = ~(w12057 | w12131);
assign w12142 = v5637;
assign v5638 = ~(w12051 | w12054);
assign w12143 = v5638;
assign v5639 = ~(w12066 | w12072);
assign w12144 = v5639;
assign v5640 = ~(w12089 | w12095);
assign w12145 = v5640;
assign w12146 = pi27 & pi54;
assign w12147 = pi39 & pi42;
assign v5641 = ~(w12016 | w12147);
assign w12148 = v5641;
assign w12149 = pi39 & pi43;
assign w12150 = w12013 & w12149;
assign v5642 = ~(w12148 | w12150);
assign w12151 = v5642;
assign w12152 = w12146 & ~w12151;
assign w12153 = ~w12146 & w12151;
assign v5643 = ~(w12152 | w12153);
assign w12154 = v5643;
assign v5644 = ~(w12145 | w12154);
assign w12155 = v5644;
assign w12156 = w12145 & w12154;
assign v5645 = ~(w12155 | w12156);
assign w12157 = v5645;
assign w12158 = w12144 & ~w12157;
assign w12159 = ~w12144 & w12157;
assign v5646 = ~(w12158 | w12159);
assign w12160 = v5646;
assign w12161 = (~w12076 & ~w12077) | (~w12076 & w17207) | (~w12077 & w17207);
assign v5647 = ~(w12099 | w12102);
assign w12162 = v5647;
assign v5648 = ~(w12161 | w12162);
assign w12163 = v5648;
assign w12164 = w12161 & w12162;
assign v5649 = ~(w12163 | w12164);
assign w12165 = v5649;
assign w12166 = w12160 & w12165;
assign v5650 = ~(w12160 | w12165);
assign w12167 = v5650;
assign v5651 = ~(w12166 | w12167);
assign w12168 = v5651;
assign w12169 = ~w12143 & w12168;
assign w12170 = w12143 & ~w12168;
assign v5652 = ~(w12169 | w12170);
assign w12171 = v5652;
assign w12172 = w12012 & ~w12015;
assign v5653 = ~(w12017 | w12172);
assign w12173 = v5653;
assign w12174 = w11851 & ~w12035;
assign v5654 = ~(w12037 | w12174);
assign w12175 = v5654;
assign v5655 = ~(w12173 | w12175);
assign w12176 = v5655;
assign w12177 = w12173 & w12175;
assign v5656 = ~(w12176 | w12177);
assign w12178 = v5656;
assign v5657 = ~(w12022 | w12025);
assign w12179 = v5657;
assign v5658 = ~(w12024 | w12179);
assign w12180 = v5658;
assign v5659 = ~(w12178 | w12180);
assign w12181 = v5659;
assign w12182 = w12178 & w12180;
assign v5660 = ~(w12181 | w12182);
assign w12183 = v5660;
assign w12184 = (~w12030 & ~w12032) | (~w12030 & w17841) | (~w12032 & w17841);
assign w12185 = (~w11997 & ~w11999) | (~w11997 & w17842) | (~w11999 & w17842);
assign v5661 = ~(w12184 | w12185);
assign w12186 = v5661;
assign w12187 = w12184 & w12185;
assign v5662 = ~(w12186 | w12187);
assign w12188 = v5662;
assign w12189 = w12183 & w12188;
assign v5663 = ~(w12183 | w12188);
assign w12190 = v5663;
assign v5664 = ~(w12189 | w12190);
assign w12191 = v5664;
assign v5665 = ~(w11956 | w11960);
assign w12192 = v5665;
assign w12193 = w11963 & ~w11965;
assign v5666 = ~(w11967 | w12193);
assign w12194 = v5666;
assign v5667 = ~(w12192 | w12194);
assign w12195 = v5667;
assign w12196 = w12192 & w12194;
assign v5668 = ~(w12195 | w12196);
assign w12197 = v5668;
assign w12198 = pi30 & pi51;
assign w12199 = pi31 & pi50;
assign v5669 = ~(w12003 | w12199);
assign w12200 = v5669;
assign w12201 = pi32 & pi50;
assign w12202 = w12000 & w12201;
assign v5670 = ~(w12200 | w12202);
assign w12203 = v5670;
assign w12204 = w12198 & ~w12203;
assign w12205 = ~w12198 & w12203;
assign v5671 = ~(w12204 | w12205);
assign w12206 = v5671;
assign w12207 = ~w12197 & w12206;
assign w12208 = w12197 & ~w12206;
assign v5672 = ~(w12207 | w12208);
assign w12209 = v5672;
assign v5673 = ~(w11895 | w11975);
assign w12210 = v5673;
assign v5674 = ~(w11974 | w12210);
assign w12211 = v5674;
assign w12212 = w11883 & ~w12002;
assign v5675 = ~(w12004 | w12212);
assign w12213 = v5675;
assign w12214 = w12211 & ~w12213;
assign w12215 = ~w12211 & w12213;
assign v5676 = ~(w12214 | w12215);
assign w12216 = v5676;
assign w12217 = w11986 & ~w11988;
assign v5677 = ~(w11990 | w12217);
assign w12218 = v5677;
assign w12219 = ~w12216 & w12218;
assign w12220 = w12216 & ~w12218;
assign v5678 = ~(w12219 | w12220);
assign w12221 = v5678;
assign w12222 = (~w11980 & ~w11982) | (~w11980 & w17843) | (~w11982 & w17843);
assign w12223 = ~w12221 & w12222;
assign w12224 = w12221 & ~w12222;
assign v5679 = ~(w12223 | w12224);
assign w12225 = v5679;
assign w12226 = w12209 & w12225;
assign v5680 = ~(w12209 | w12225);
assign w12227 = v5680;
assign v5681 = ~(w12226 | w12227);
assign w12228 = v5681;
assign v5682 = ~(w12045 | w12048);
assign w12229 = v5682;
assign w12230 = w12228 & ~w12229;
assign w12231 = ~w12228 & w12229;
assign v5683 = ~(w12230 | w12231);
assign w12232 = v5683;
assign w12233 = w12191 & w12232;
assign v5684 = ~(w12191 | w12232);
assign w12234 = v5684;
assign v5685 = ~(w12233 | w12234);
assign w12235 = v5685;
assign w12236 = w12171 & w12235;
assign v5686 = ~(w12171 | w12235);
assign w12237 = v5686;
assign v5687 = ~(w12236 | w12237);
assign w12238 = v5687;
assign v5688 = ~(w12125 | w12128);
assign w12239 = v5688;
assign w12240 = (~w12082 & ~w12084) | (~w12082 & w17844) | (~w12084 & w17844);
assign w12241 = (~w12119 & ~w12121) | (~w12119 & w17208) | (~w12121 & w17208);
assign w12242 = (~w12111 & ~w12113) | (~w12111 & w17845) | (~w12113 & w17845);
assign w12243 = ~pi40 & pi41;
assign w12244 = w11955 & ~w12243;
assign w12245 = ~w11955 & w12243;
assign v5689 = ~(w12244 | w12245);
assign w12246 = v5689;
assign w12247 = pi25 & pi56;
assign w12248 = pi23 & pi58;
assign v5690 = ~(w12247 | w12248);
assign w12249 = v5690;
assign w12250 = w12247 & w12248;
assign v5691 = ~(w12249 | w12250);
assign w12251 = v5691;
assign w12252 = w11989 & ~w12251;
assign w12253 = ~w11989 & w12251;
assign v5692 = ~(w12252 | w12253);
assign w12254 = v5692;
assign v5693 = ~(w12246 | w12254);
assign w12255 = v5693;
assign w12256 = w12246 & w12254;
assign v5694 = ~(w12255 | w12256);
assign w12257 = v5694;
assign w12258 = pi24 & pi57;
assign w12259 = pi33 & pi48;
assign w12260 = pi34 & pi47;
assign v5695 = ~(w12259 | w12260);
assign w12261 = v5695;
assign w12262 = pi34 & pi48;
assign w12263 = w11895 & w12262;
assign v5696 = ~(w12261 | w12263);
assign w12264 = v5696;
assign w12265 = w12258 & ~w12264;
assign w12266 = ~w12258 & w12264;
assign v5697 = ~(w12265 | w12266);
assign w12267 = v5697;
assign w12268 = w12257 & ~w12267;
assign w12269 = ~w12257 & w12267;
assign v5698 = ~(w12268 | w12269);
assign w12270 = v5698;
assign w12271 = ~w12242 & w12270;
assign w12272 = w12242 & ~w12270;
assign v5699 = ~(w12271 | w12272);
assign w12273 = v5699;
assign w12274 = pi18 & pi63;
assign w12275 = pi20 & pi61;
assign w12276 = pi21 & pi60;
assign v5700 = ~(w12275 | w12276);
assign w12277 = v5700;
assign w12278 = pi21 & pi61;
assign w12279 = w11986 & w12278;
assign v5701 = ~(w12277 | w12279);
assign w12280 = v5701;
assign w12281 = w12274 & ~w12280;
assign w12282 = ~w12274 & w12280;
assign v5702 = ~(w12281 | w12282);
assign w12283 = v5702;
assign w12284 = pi35 & pi46;
assign w12285 = pi37 & pi44;
assign v5703 = ~(w11966 | w12285);
assign w12286 = v5703;
assign w12287 = pi37 & pi45;
assign w12288 = w11964 & w12287;
assign v5704 = ~(w12286 | w12288);
assign w12289 = v5704;
assign w12290 = w12284 & ~w12289;
assign w12291 = ~w12284 & w12289;
assign v5705 = ~(w12290 | w12291);
assign w12292 = v5705;
assign v5706 = ~(w12283 | w12292);
assign w12293 = v5706;
assign w12294 = w12283 & w12292;
assign v5707 = ~(w12293 | w12294);
assign w12295 = v5707;
assign w12296 = pi26 & pi55;
assign w12297 = pi29 & pi52;
assign v5708 = ~(w12036 | w12297);
assign w12298 = v5708;
assign w12299 = pi29 & pi53;
assign w12300 = w12033 & w12299;
assign v5709 = ~(w12298 | w12300);
assign w12301 = v5709;
assign w12302 = w12296 & ~w12301;
assign w12303 = ~w12296 & w12301;
assign v5710 = ~(w12302 | w12303);
assign w12304 = v5710;
assign w12305 = w12295 & ~w12304;
assign w12306 = ~w12295 & w12304;
assign v5711 = ~(w12305 | w12306);
assign w12307 = v5711;
assign v5712 = ~(w12273 | w12307);
assign w12308 = v5712;
assign w12309 = w12273 & w12307;
assign v5713 = ~(w12308 | w12309);
assign w12310 = v5713;
assign w12311 = ~w12241 & w12310;
assign w12312 = w12241 & ~w12310;
assign v5714 = ~(w12311 | w12312);
assign w12313 = v5714;
assign w12314 = ~w12240 & w12313;
assign w12315 = w12240 & ~w12313;
assign v5715 = ~(w12314 | w12315);
assign w12316 = v5715;
assign w12317 = ~w12239 & w12316;
assign w12318 = w12239 & ~w12316;
assign v5716 = ~(w12317 | w12318);
assign w12319 = v5716;
assign w12320 = w12238 & w12319;
assign v5717 = ~(w12238 | w12319);
assign w12321 = v5717;
assign v5718 = ~(w12320 | w12321);
assign w12322 = v5718;
assign w12323 = w12142 & ~w12322;
assign w12324 = ~w12142 & w12322;
assign v5719 = ~(w12323 | w12324);
assign w12325 = v5719;
assign w12326 = w12141 & ~w12325;
assign w12327 = ~w12141 & w12325;
assign v5720 = ~(w12326 | w12327);
assign w12328 = v5720;
assign w12329 = (~w7754 & w17846) | (~w7754 & w17847) | (w17846 & w17847);
assign v5721 = ~(w12317 | w12320);
assign w12330 = v5721;
assign w12331 = (~w12311 & ~w12313) | (~w12311 & w17848) | (~w12313 & w17848);
assign v5722 = ~(w12176 | w12182);
assign w12332 = v5722;
assign v5723 = ~(w12214 | w12220);
assign w12333 = v5723;
assign w12334 = pi28 & pi54;
assign w12335 = pi27 & pi55;
assign w12336 = pi25 & pi57;
assign v5724 = ~(w12335 | w12336);
assign w12337 = v5724;
assign w12338 = w12335 & w12336;
assign v5725 = ~(w12337 | w12338);
assign w12339 = v5725;
assign w12340 = w12334 & ~w12339;
assign w12341 = ~w12334 & w12339;
assign v5726 = ~(w12340 | w12341);
assign w12342 = v5726;
assign v5727 = ~(w12333 | w12342);
assign w12343 = v5727;
assign w12344 = w12333 & w12342;
assign v5728 = ~(w12343 | w12344);
assign w12345 = v5728;
assign w12346 = w12332 & ~w12345;
assign w12347 = ~w12332 & w12345;
assign v5729 = ~(w12346 | w12347);
assign w12348 = v5729;
assign v5730 = ~(w12224 | w12226);
assign w12349 = v5730;
assign v5731 = ~(w12186 | w12189);
assign w12350 = v5731;
assign v5732 = ~(w12349 | w12350);
assign w12351 = v5732;
assign w12352 = w12349 & w12350;
assign v5733 = ~(w12351 | w12352);
assign w12353 = v5733;
assign w12354 = w12348 & w12353;
assign v5734 = ~(w12348 | w12353);
assign w12355 = v5734;
assign v5735 = ~(w12354 | w12355);
assign w12356 = v5735;
assign w12357 = ~w12331 & w12356;
assign w12358 = w12331 & ~w12356;
assign v5736 = ~(w12357 | w12358);
assign w12359 = v5736;
assign v5737 = ~(w12271 | w12309);
assign w12360 = v5737;
assign w12361 = w12198 & ~w12200;
assign v5738 = ~(w12202 | w12361);
assign w12362 = v5738;
assign w12363 = w12258 & ~w12261;
assign v5739 = ~(w12263 | w12363);
assign w12364 = v5739;
assign v5740 = ~(w12362 | w12364);
assign w12365 = v5740;
assign w12366 = w12362 & w12364;
assign v5741 = ~(w12365 | w12366);
assign w12367 = v5741;
assign w12368 = w12296 & ~w12298;
assign v5742 = ~(w12300 | w12368);
assign w12369 = v5742;
assign w12370 = ~w12367 & w12369;
assign w12371 = w12367 & ~w12369;
assign v5743 = ~(w12370 | w12371);
assign w12372 = v5743;
assign v5744 = ~(w11989 | w12250);
assign w12373 = v5744;
assign v5745 = ~(w12249 | w12373);
assign w12374 = v5745;
assign w12375 = w12274 & ~w12277;
assign v5746 = ~(w12279 | w12375);
assign w12376 = v5746;
assign w12377 = w12374 & ~w12376;
assign w12378 = ~w12374 & w12376;
assign v5747 = ~(w12377 | w12378);
assign w12379 = v5747;
assign w12380 = w12284 & ~w12286;
assign v5748 = ~(w12288 | w12380);
assign w12381 = v5748;
assign w12382 = ~w12379 & w12381;
assign w12383 = w12379 & ~w12381;
assign v5749 = ~(w12382 | w12383);
assign w12384 = v5749;
assign v5750 = ~(w12293 | w12305);
assign w12385 = v5750;
assign w12386 = ~w12384 & w12385;
assign w12387 = w12384 & ~w12385;
assign v5751 = ~(w12386 | w12387);
assign w12388 = v5751;
assign w12389 = w12372 & w12388;
assign v5752 = ~(w12372 | w12388);
assign w12390 = v5752;
assign v5753 = ~(w12389 | w12390);
assign w12391 = v5753;
assign w12392 = ~w12360 & w12391;
assign w12393 = w12360 & ~w12391;
assign v5754 = ~(w12392 | w12393);
assign w12394 = v5754;
assign v5755 = ~(w12195 | w12208);
assign w12395 = v5755;
assign v5756 = ~(w12255 | w12268);
assign w12396 = v5756;
assign v5757 = ~(w12395 | w12396);
assign w12397 = v5757;
assign w12398 = w12395 & w12396;
assign v5758 = ~(w12397 | w12398);
assign w12399 = v5758;
assign w12400 = pi19 & pi63;
assign v5759 = ~(pi40 | w11955);
assign w12401 = v5759;
assign w12402 = pi41 & ~w12401;
assign v5760 = ~(w12400 | w12402);
assign w12403 = v5760;
assign w12404 = w12400 & w12402;
assign v5761 = ~(w12403 | w12404);
assign w12405 = v5761;
assign w12406 = w12146 & ~w12148;
assign v5762 = ~(w12150 | w12406);
assign w12407 = v5762;
assign w12408 = w12405 & ~w12407;
assign w12409 = ~w12405 & w12407;
assign v5763 = ~(w12408 | w12409);
assign w12410 = v5763;
assign w12411 = w12399 & w12410;
assign v5764 = ~(w12399 | w12410);
assign w12412 = v5764;
assign v5765 = ~(w12411 | w12412);
assign w12413 = v5765;
assign w12414 = w12394 & w12413;
assign v5766 = ~(w12394 | w12413);
assign w12415 = v5766;
assign v5767 = ~(w12414 | w12415);
assign w12416 = v5767;
assign w12417 = w12359 & w12416;
assign v5768 = ~(w12359 | w12416);
assign w12418 = v5768;
assign v5769 = ~(w12417 | w12418);
assign w12419 = v5769;
assign v5770 = ~(w12169 | w12236);
assign w12420 = v5770;
assign v5771 = ~(w12230 | w12233);
assign w12421 = v5771;
assign v5772 = ~(w12163 | w12166);
assign w12422 = v5772;
assign v5773 = ~(w12155 | w12159);
assign w12423 = v5773;
assign w12424 = pi33 & pi49;
assign v5774 = ~(w12262 | w12424);
assign w12425 = v5774;
assign w12426 = pi34 & pi49;
assign w12427 = w12259 & w12426;
assign v5775 = ~(w12425 | w12427);
assign w12428 = v5775;
assign w12429 = w12201 & ~w12428;
assign w12430 = ~w12201 & w12428;
assign v5776 = ~(w12429 | w12430);
assign w12431 = v5776;
assign w12432 = pi20 & pi62;
assign w12433 = pi31 & pi51;
assign v5777 = ~(w12278 | w12433);
assign w12434 = v5777;
assign w12435 = w12278 & w12433;
assign v5778 = ~(w12434 | w12435);
assign w12436 = v5778;
assign w12437 = w12432 & ~w12436;
assign w12438 = ~w12432 & w12436;
assign v5779 = ~(w12437 | w12438);
assign w12439 = v5779;
assign v5780 = ~(w12431 | w12439);
assign w12440 = v5780;
assign w12441 = w12431 & w12439;
assign v5781 = ~(w12440 | w12441);
assign w12442 = v5781;
assign w12443 = pi22 & pi60;
assign w12444 = pi24 & pi58;
assign w12445 = pi23 & pi59;
assign v5782 = ~(w12444 | w12445);
assign w12446 = v5782;
assign w12447 = pi24 & pi59;
assign w12448 = w12248 & w12447;
assign v5783 = ~(w12446 | w12448);
assign w12449 = v5783;
assign w12450 = w12443 & ~w12449;
assign w12451 = ~w12443 & w12449;
assign v5784 = ~(w12450 | w12451);
assign w12452 = v5784;
assign w12453 = w12442 & ~w12452;
assign w12454 = ~w12442 & w12452;
assign v5785 = ~(w12453 | w12454);
assign w12455 = v5785;
assign w12456 = ~w12423 & w12455;
assign w12457 = w12423 & ~w12455;
assign v5786 = ~(w12456 | w12457);
assign w12458 = v5786;
assign w12459 = pi40 & pi42;
assign w12460 = pi30 & pi52;
assign v5787 = ~(w12299 | w12460);
assign w12461 = v5787;
assign w12462 = pi30 & pi53;
assign w12463 = w12297 & w12462;
assign v5788 = ~(w12461 | w12463);
assign w12464 = v5788;
assign w12465 = w12459 & ~w12464;
assign w12466 = ~w12459 & w12464;
assign v5789 = ~(w12465 | w12466);
assign w12467 = v5789;
assign w12468 = pi26 & pi56;
assign w12469 = pi38 & pi44;
assign v5790 = ~(w12149 | w12469);
assign w12470 = v5790;
assign w12471 = pi39 & pi44;
assign w12472 = w12016 & w12471;
assign v5791 = ~(w12470 | w12472);
assign w12473 = v5791;
assign w12474 = w12468 & ~w12473;
assign w12475 = ~w12468 & w12473;
assign v5792 = ~(w12474 | w12475);
assign w12476 = v5792;
assign v5793 = ~(w12467 | w12476);
assign w12477 = v5793;
assign w12478 = w12467 & w12476;
assign v5794 = ~(w12477 | w12478);
assign w12479 = v5794;
assign w12480 = pi35 & pi47;
assign w12481 = pi36 & pi46;
assign v5795 = ~(w12287 | w12481);
assign w12482 = v5795;
assign w12483 = pi37 & pi46;
assign w12484 = w11966 & w12483;
assign v5796 = ~(w12482 | w12484);
assign w12485 = v5796;
assign w12486 = w12480 & ~w12485;
assign w12487 = ~w12480 & w12485;
assign v5797 = ~(w12486 | w12487);
assign w12488 = v5797;
assign w12489 = w12479 & ~w12488;
assign w12490 = ~w12479 & w12488;
assign v5798 = ~(w12489 | w12490);
assign w12491 = v5798;
assign v5799 = ~(w12458 | w12491);
assign w12492 = v5799;
assign w12493 = w12458 & w12491;
assign v5800 = ~(w12492 | w12493);
assign w12494 = v5800;
assign w12495 = ~w12422 & w12494;
assign w12496 = w12422 & ~w12494;
assign v5801 = ~(w12495 | w12496);
assign w12497 = v5801;
assign w12498 = ~w12421 & w12497;
assign w12499 = w12421 & ~w12497;
assign v5802 = ~(w12498 | w12499);
assign w12500 = v5802;
assign w12501 = ~w12420 & w12500;
assign w12502 = w12420 & ~w12500;
assign v5803 = ~(w12501 | w12502);
assign w12503 = v5803;
assign w12504 = w12419 & w12503;
assign v5804 = ~(w12419 | w12503);
assign w12505 = v5804;
assign v5805 = ~(w12504 | w12505);
assign w12506 = v5805;
assign w12507 = ~w12330 & w12506;
assign w12508 = w12330 & ~w12506;
assign v5806 = ~(w12507 | w12508);
assign w12509 = v5806;
assign w12510 = (~w10008 & w17849) | (~w10008 & w17850) | (w17849 & w17850);
assign w12511 = (w10008 & w17851) | (w10008 & w17852) | (w17851 & w17852);
assign v5807 = ~(w12510 | w12511);
assign w12512 = v5807;
assign v5808 = ~(w12501 | w12504);
assign w12513 = v5808;
assign v5809 = ~(w12357 | w12417);
assign w12514 = v5809;
assign v5810 = ~(w12392 | w12414);
assign w12515 = v5810;
assign v5811 = ~(w12351 | w12354);
assign w12516 = v5811;
assign v5812 = ~(w12343 | w12347);
assign w12517 = v5812;
assign w12518 = pi29 & pi54;
assign w12519 = pi40 & pi43;
assign v5813 = ~(w12471 | w12519);
assign w12520 = v5813;
assign w12521 = pi40 & pi44;
assign w12522 = w12149 & w12521;
assign v5814 = ~(w12520 | w12522);
assign w12523 = v5814;
assign w12524 = w12518 & ~w12523;
assign w12525 = ~w12518 & w12523;
assign v5815 = ~(w12524 | w12525);
assign w12526 = v5815;
assign w12527 = pi21 & pi62;
assign w12528 = ~pi41 & pi42;
assign w12529 = w12527 & ~w12528;
assign w12530 = ~w12527 & w12528;
assign v5816 = ~(w12529 | w12530);
assign w12531 = v5816;
assign v5817 = ~(w12526 | w12531);
assign w12532 = v5817;
assign w12533 = w12526 & w12531;
assign v5818 = ~(w12532 | w12533);
assign w12534 = v5818;
assign w12535 = pi33 & pi50;
assign w12536 = pi35 & pi48;
assign v5819 = ~(w12426 | w12536);
assign w12537 = v5819;
assign w12538 = pi35 & pi49;
assign w12539 = w12262 & w12538;
assign v5820 = ~(w12537 | w12539);
assign w12540 = v5820;
assign w12541 = w12535 & ~w12540;
assign w12542 = ~w12535 & w12540;
assign v5821 = ~(w12541 | w12542);
assign w12543 = v5821;
assign w12544 = w12534 & ~w12543;
assign w12545 = ~w12534 & w12543;
assign v5822 = ~(w12544 | w12545);
assign w12546 = v5822;
assign w12547 = ~w12517 & w12546;
assign w12548 = w12517 & ~w12546;
assign v5823 = ~(w12547 | w12548);
assign w12549 = v5823;
assign w12550 = pi36 & pi47;
assign w12551 = pi38 & pi45;
assign v5824 = ~(w12483 | w12551);
assign w12552 = v5824;
assign w12553 = pi38 & pi46;
assign w12554 = w12287 & w12553;
assign v5825 = ~(w12552 | w12554);
assign w12555 = v5825;
assign w12556 = w12550 & ~w12555;
assign w12557 = ~w12550 & w12555;
assign v5826 = ~(w12556 | w12557);
assign w12558 = v5826;
assign w12559 = pi25 & pi58;
assign w12560 = pi26 & pi57;
assign w12561 = pi32 & pi51;
assign v5827 = ~(w12560 | w12561);
assign w12562 = v5827;
assign w12563 = w12560 & w12561;
assign v5828 = ~(w12562 | w12563);
assign w12564 = v5828;
assign w12565 = w12559 & ~w12564;
assign w12566 = ~w12559 & w12564;
assign v5829 = ~(w12565 | w12566);
assign w12567 = v5829;
assign v5830 = ~(w12558 | w12567);
assign w12568 = v5830;
assign w12569 = w12558 & w12567;
assign v5831 = ~(w12568 | w12569);
assign w12570 = v5831;
assign w12571 = pi27 & pi56;
assign w12572 = pi20 & pi63;
assign w12573 = pi22 & pi61;
assign v5832 = ~(w12572 | w12573);
assign w12574 = v5832;
assign w12575 = w12572 & w12573;
assign v5833 = ~(w12574 | w12575);
assign w12576 = v5833;
assign w12577 = w12571 & ~w12576;
assign w12578 = ~w12571 & w12576;
assign v5834 = ~(w12577 | w12578);
assign w12579 = v5834;
assign w12580 = w12570 & ~w12579;
assign w12581 = ~w12570 & w12579;
assign v5835 = ~(w12580 | w12581);
assign w12582 = v5835;
assign v5836 = ~(w12549 | w12582);
assign w12583 = v5836;
assign w12584 = w12549 & w12582;
assign v5837 = ~(w12583 | w12584);
assign w12585 = v5837;
assign w12586 = ~w12516 & w12585;
assign w12587 = w12516 & ~w12585;
assign v5838 = ~(w12586 | w12587);
assign w12588 = v5838;
assign w12589 = ~w12515 & w12588;
assign w12590 = w12515 & ~w12588;
assign v5839 = ~(w12589 | w12590);
assign w12591 = v5839;
assign w12592 = ~w12514 & w12591;
assign w12593 = w12514 & ~w12591;
assign v5840 = ~(w12592 | w12593);
assign w12594 = v5840;
assign w12595 = w12443 & ~w12446;
assign v5841 = ~(w12448 | w12595);
assign w12596 = v5841;
assign w12597 = w12480 & ~w12482;
assign v5842 = ~(w12484 | w12597);
assign w12598 = v5842;
assign v5843 = ~(w12596 | w12598);
assign w12599 = v5843;
assign w12600 = w12596 & w12598;
assign v5844 = ~(w12599 | w12600);
assign w12601 = v5844;
assign w12602 = w12468 & ~w12470;
assign v5845 = ~(w12472 | w12602);
assign w12603 = v5845;
assign w12604 = ~w12601 & w12603;
assign w12605 = w12601 & ~w12603;
assign v5846 = ~(w12604 | w12605);
assign w12606 = v5846;
assign v5847 = ~(w12432 | w12435);
assign w12607 = v5847;
assign v5848 = ~(w12434 | w12607);
assign w12608 = v5848;
assign w12609 = w12201 & ~w12425;
assign v5849 = ~(w12427 | w12609);
assign w12610 = v5849;
assign w12611 = w12608 & ~w12610;
assign w12612 = ~w12608 & w12610;
assign v5850 = ~(w12611 | w12612);
assign w12613 = v5850;
assign v5851 = ~(w12334 | w12338);
assign w12614 = v5851;
assign v5852 = ~(w12337 | w12614);
assign w12615 = v5852;
assign v5853 = ~(w12613 | w12615);
assign w12616 = v5853;
assign w12617 = w12613 & w12615;
assign v5854 = ~(w12616 | w12617);
assign w12618 = v5854;
assign v5855 = ~(w12477 | w12489);
assign w12619 = v5855;
assign w12620 = ~w12618 & w12619;
assign w12621 = w12618 & ~w12619;
assign v5856 = ~(w12620 | w12621);
assign w12622 = v5856;
assign w12623 = w12606 & w12622;
assign v5857 = ~(w12606 | w12622);
assign w12624 = v5857;
assign v5858 = ~(w12623 | w12624);
assign w12625 = v5858;
assign v5859 = ~(w12456 | w12493);
assign w12626 = v5859;
assign v5860 = ~(w12387 | w12389);
assign w12627 = v5860;
assign v5861 = ~(w12626 | w12627);
assign w12628 = v5861;
assign w12629 = w12626 & w12627;
assign v5862 = ~(w12628 | w12629);
assign w12630 = v5862;
assign w12631 = w12625 & w12630;
assign v5863 = ~(w12625 | w12630);
assign w12632 = v5863;
assign v5864 = ~(w12631 | w12632);
assign w12633 = v5864;
assign v5865 = ~(w12495 | w12498);
assign w12634 = v5865;
assign v5866 = ~(w12440 | w12453);
assign w12635 = v5866;
assign v5867 = ~(w12365 | w12371);
assign w12636 = v5867;
assign v5868 = ~(w12377 | w12383);
assign w12637 = v5868;
assign v5869 = ~(w12636 | w12637);
assign w12638 = v5869;
assign w12639 = w12636 & w12637;
assign v5870 = ~(w12638 | w12639);
assign w12640 = v5870;
assign w12641 = w12635 & ~w12640;
assign w12642 = ~w12635 & w12640;
assign v5871 = ~(w12641 | w12642);
assign w12643 = v5871;
assign w12644 = pi23 & pi60;
assign v5872 = ~(w12447 | w12644);
assign w12645 = v5872;
assign w12646 = pi24 & pi60;
assign w12647 = w12445 & w12646;
assign v5873 = ~(w12645 | w12647);
assign w12648 = v5873;
assign w12649 = w12459 & ~w12461;
assign v5874 = ~(w12463 | w12649);
assign w12650 = v5874;
assign w12651 = w12648 & ~w12650;
assign w12652 = ~w12648 & w12650;
assign v5875 = ~(w12651 | w12652);
assign w12653 = v5875;
assign w12654 = pi31 & pi52;
assign w12655 = pi28 & pi55;
assign v5876 = ~(w12462 | w12655);
assign w12656 = v5876;
assign w12657 = w12462 & w12655;
assign v5877 = ~(w12656 | w12657);
assign w12658 = v5877;
assign w12659 = w12654 & ~w12658;
assign w12660 = ~w12654 & w12658;
assign v5878 = ~(w12659 | w12660);
assign w12661 = v5878;
assign w12662 = w12653 & ~w12661;
assign w12663 = ~w12653 & w12661;
assign v5879 = ~(w12662 | w12663);
assign w12664 = v5879;
assign v5880 = ~(w12404 | w12408);
assign w12665 = v5880;
assign w12666 = ~w12664 & w12665;
assign w12667 = w12664 & ~w12665;
assign v5881 = ~(w12666 | w12667);
assign w12668 = v5881;
assign v5882 = ~(w12397 | w12411);
assign w12669 = v5882;
assign w12670 = ~w12668 & w12669;
assign w12671 = w12668 & ~w12669;
assign v5883 = ~(w12670 | w12671);
assign w12672 = v5883;
assign w12673 = w12643 & w12672;
assign v5884 = ~(w12643 | w12672);
assign w12674 = v5884;
assign v5885 = ~(w12673 | w12674);
assign w12675 = v5885;
assign w12676 = ~w12634 & w12675;
assign w12677 = w12634 & ~w12675;
assign v5886 = ~(w12676 | w12677);
assign w12678 = v5886;
assign w12679 = w12633 & w12678;
assign v5887 = ~(w12633 | w12678);
assign w12680 = v5887;
assign v5888 = ~(w12679 | w12680);
assign w12681 = v5888;
assign v5889 = ~(w12594 | w12681);
assign w12682 = v5889;
assign w12683 = w12594 & w12681;
assign v5890 = ~(w12682 | w12683);
assign w12684 = v5890;
assign w12685 = ~w12513 & w12684;
assign w12686 = w12513 & ~w12684;
assign v5891 = ~(w12685 | w12686);
assign w12687 = v5891;
assign v5892 = ~(w12323 | w12508);
assign w12688 = v5892;
assign w12689 = (~w8795 & w17632) | (~w8795 & w17633) | (w17632 & w17633);
assign w12690 = w12687 & w12689;
assign v5893 = ~(w12687 | w12689);
assign w12691 = v5893;
assign v5894 = ~(w12690 | w12691);
assign w12692 = v5894;
assign v5895 = ~(w12507 | w12685);
assign w12693 = v5895;
assign v5896 = ~(w12592 | w12683);
assign w12694 = v5896;
assign v5897 = ~(w12676 | w12679);
assign w12695 = v5897;
assign v5898 = ~(w12638 | w12642);
assign w12696 = v5898;
assign w12697 = (~w12647 & w12650) | (~w12647 & w16774) | (w12650 & w16774);
assign v5899 = ~(w12571 | w12575);
assign w12698 = v5899;
assign v5900 = ~(w12574 | w12698);
assign w12699 = v5900;
assign w12700 = ~w12697 & w12699;
assign w12701 = w12697 & ~w12699;
assign v5901 = ~(w12700 | w12701);
assign w12702 = v5901;
assign w12703 = pi26 & pi58;
assign w12704 = pi31 & pi53;
assign w12705 = pi32 & pi52;
assign v5902 = ~(w12704 | w12705);
assign w12706 = v5902;
assign w12707 = pi32 & pi53;
assign w12708 = w12654 & w12707;
assign v5903 = ~(w12706 | w12708);
assign w12709 = v5903;
assign w12710 = w12703 & ~w12709;
assign w12711 = ~w12703 & w12709;
assign v5904 = ~(w12710 | w12711);
assign w12712 = v5904;
assign w12713 = ~w12702 & w12712;
assign w12714 = w12702 & ~w12712;
assign v5905 = ~(w12713 | w12714);
assign w12715 = v5905;
assign v5906 = ~(w12662 | w12667);
assign w12716 = v5906;
assign w12717 = w12715 & ~w12716;
assign w12718 = ~w12715 & w12716;
assign v5907 = ~(w12717 | w12718);
assign w12719 = v5907;
assign w12720 = w12696 & ~w12719;
assign w12721 = ~w12696 & w12719;
assign v5908 = ~(w12720 | w12721);
assign w12722 = v5908;
assign v5909 = ~(w12671 | w12673);
assign w12723 = v5909;
assign w12724 = ~w12722 & w12723;
assign w12725 = w12722 & ~w12723;
assign v5910 = ~(w12724 | w12725);
assign w12726 = v5910;
assign w12727 = w12535 & ~w12537;
assign v5911 = ~(w12539 | w12727);
assign w12728 = v5911;
assign w12729 = w12550 & ~w12552;
assign v5912 = ~(w12554 | w12729);
assign w12730 = v5912;
assign v5913 = ~(w12728 | w12730);
assign w12731 = v5913;
assign w12732 = w12728 & w12730;
assign v5914 = ~(w12731 | w12732);
assign w12733 = v5914;
assign v5915 = ~(w12559 | w12563);
assign w12734 = v5915;
assign v5916 = ~(w12562 | w12734);
assign w12735 = v5916;
assign v5917 = ~(w12733 | w12735);
assign w12736 = v5917;
assign w12737 = w12733 & w12735;
assign v5918 = ~(w12736 | w12737);
assign w12738 = v5918;
assign w12739 = (~w12599 & ~w12601) | (~w12599 & w16775) | (~w12601 & w16775);
assign w12740 = (~w12611 & ~w12613) | (~w12611 & w16776) | (~w12613 & w16776);
assign v5919 = ~(w12739 | w12740);
assign w12741 = v5919;
assign w12742 = w12739 & w12740;
assign v5920 = ~(w12741 | w12742);
assign w12743 = v5920;
assign w12744 = w12738 & w12743;
assign v5921 = ~(w12738 | w12743);
assign w12745 = v5921;
assign v5922 = ~(w12744 | w12745);
assign w12746 = v5922;
assign w12747 = pi21 & pi63;
assign w12748 = pi22 & pi62;
assign w12749 = pi23 & pi61;
assign v5923 = ~(w12748 | w12749);
assign w12750 = v5923;
assign w12751 = pi23 & pi62;
assign w12752 = w12573 & w12751;
assign v5924 = ~(w12750 | w12752);
assign w12753 = v5924;
assign w12754 = w12747 & ~w12753;
assign w12755 = ~w12747 & w12753;
assign v5925 = ~(w12754 | w12755);
assign w12756 = v5925;
assign w12757 = pi33 & pi51;
assign w12758 = pi25 & pi59;
assign v5926 = ~(w12646 | w12758);
assign w12759 = v5926;
assign w12760 = pi25 & pi60;
assign w12761 = w12447 & w12760;
assign v5927 = ~(w12759 | w12761);
assign w12762 = v5927;
assign w12763 = w12757 & ~w12762;
assign w12764 = ~w12757 & w12762;
assign v5928 = ~(w12763 | w12764);
assign w12765 = v5928;
assign v5929 = ~(w12756 | w12765);
assign w12766 = v5929;
assign w12767 = w12756 & w12765;
assign v5930 = ~(w12766 | w12767);
assign w12768 = v5930;
assign w12769 = pi34 & pi50;
assign w12770 = pi36 & pi48;
assign v5931 = ~(w12538 | w12770);
assign w12771 = v5931;
assign w12772 = pi36 & pi49;
assign w12773 = w12536 & w12772;
assign v5932 = ~(w12771 | w12773);
assign w12774 = v5932;
assign w12775 = w12769 & ~w12774;
assign w12776 = ~w12769 & w12774;
assign v5933 = ~(w12775 | w12776);
assign w12777 = v5933;
assign w12778 = w12768 & ~w12777;
assign w12779 = ~w12768 & w12777;
assign v5934 = ~(w12778 | w12779);
assign w12780 = v5934;
assign w12781 = pi39 & pi45;
assign w12782 = pi41 & pi43;
assign v5935 = ~(w12521 | w12782);
assign w12783 = v5935;
assign w12784 = pi41 & pi44;
assign w12785 = w12519 & w12784;
assign v5936 = ~(w12783 | w12785);
assign w12786 = v5936;
assign w12787 = w12781 & ~w12786;
assign w12788 = ~w12781 & w12786;
assign v5937 = ~(w12787 | w12788);
assign w12789 = v5937;
assign w12790 = pi28 & pi56;
assign w12791 = pi29 & pi55;
assign v5938 = ~(w12553 | w12791);
assign w12792 = v5938;
assign w12793 = w12553 & w12791;
assign v5939 = ~(w12792 | w12793);
assign w12794 = v5939;
assign w12795 = w12790 & ~w12794;
assign w12796 = ~w12790 & w12794;
assign v5940 = ~(w12795 | w12796);
assign w12797 = v5940;
assign v5941 = ~(w12789 | w12797);
assign w12798 = v5941;
assign w12799 = w12789 & w12797;
assign v5942 = ~(w12798 | w12799);
assign w12800 = v5942;
assign w12801 = pi37 & pi47;
assign w12802 = pi27 & pi57;
assign w12803 = pi30 & pi54;
assign v5943 = ~(w12802 | w12803);
assign w12804 = v5943;
assign w12805 = w12802 & w12803;
assign v5944 = ~(w12804 | w12805);
assign w12806 = v5944;
assign w12807 = w12801 & ~w12806;
assign w12808 = ~w12801 & w12806;
assign v5945 = ~(w12807 | w12808);
assign w12809 = v5945;
assign w12810 = w12800 & ~w12809;
assign w12811 = ~w12800 & w12809;
assign v5946 = ~(w12810 | w12811);
assign w12812 = v5946;
assign w12813 = w12780 & w12812;
assign v5947 = ~(w12780 | w12812);
assign w12814 = v5947;
assign v5948 = ~(w12813 | w12814);
assign w12815 = v5948;
assign w12816 = w12746 & w12815;
assign v5949 = ~(w12746 | w12815);
assign w12817 = v5949;
assign v5950 = ~(w12816 | w12817);
assign w12818 = v5950;
assign w12819 = w12726 & w12818;
assign v5951 = ~(w12726 | w12818);
assign w12820 = v5951;
assign v5952 = ~(w12819 | w12820);
assign w12821 = v5952;
assign w12822 = ~w12695 & w12821;
assign w12823 = w12695 & ~w12821;
assign v5953 = ~(w12822 | w12823);
assign w12824 = v5953;
assign v5954 = ~(pi41 | w12527);
assign w12825 = v5954;
assign w12826 = pi42 & ~w12825;
assign w12827 = w12518 & ~w12520;
assign v5955 = ~(w12522 | w12827);
assign w12828 = v5955;
assign w12829 = w12826 & ~w12828;
assign w12830 = ~w12826 & w12828;
assign v5956 = ~(w12829 | w12830);
assign w12831 = v5956;
assign v5957 = ~(w12654 | w12657);
assign w12832 = v5957;
assign v5958 = ~(w12656 | w12832);
assign w12833 = v5958;
assign v5959 = ~(w12831 | w12833);
assign w12834 = v5959;
assign w12835 = w12831 & w12833;
assign v5960 = ~(w12834 | w12835);
assign w12836 = v5960;
assign w12837 = (~w12568 & ~w12570) | (~w12568 & w16950) | (~w12570 & w16950);
assign w12838 = (~w12532 & ~w12534) | (~w12532 & w16951) | (~w12534 & w16951);
assign v5961 = ~(w12837 | w12838);
assign w12839 = v5961;
assign w12840 = w12837 & w12838;
assign v5962 = ~(w12839 | w12840);
assign w12841 = v5962;
assign w12842 = w12836 & w12841;
assign v5963 = ~(w12836 | w12841);
assign w12843 = v5963;
assign v5964 = ~(w12842 | w12843);
assign w12844 = v5964;
assign v5965 = ~(w12547 | w12584);
assign w12845 = v5965;
assign v5966 = ~(w12621 | w12623);
assign w12846 = v5966;
assign v5967 = ~(w12845 | w12846);
assign w12847 = v5967;
assign w12848 = w12845 & w12846;
assign v5968 = ~(w12847 | w12848);
assign w12849 = v5968;
assign w12850 = w12844 & w12849;
assign v5969 = ~(w12844 | w12849);
assign w12851 = v5969;
assign v5970 = ~(w12850 | w12851);
assign w12852 = v5970;
assign v5971 = ~(w12586 | w12589);
assign w12853 = v5971;
assign v5972 = ~(w12628 | w12631);
assign w12854 = v5972;
assign v5973 = ~(w12853 | w12854);
assign w12855 = v5973;
assign w12856 = w12853 & w12854;
assign v5974 = ~(w12855 | w12856);
assign w12857 = v5974;
assign w12858 = w12852 & w12857;
assign v5975 = ~(w12852 | w12857);
assign w12859 = v5975;
assign v5976 = ~(w12858 | w12859);
assign w12860 = v5976;
assign w12861 = w12824 & w12860;
assign v5977 = ~(w12824 | w12860);
assign w12862 = v5977;
assign v5978 = ~(w12861 | w12862);
assign w12863 = v5978;
assign w12864 = w12694 & ~w12863;
assign w12865 = ~w12694 & w12863;
assign v5979 = ~(w12864 | w12865);
assign w12866 = v5979;
assign w12867 = (~w10008 & w17853) | (~w10008 & w17854) | (w17853 & w17854);
assign w12868 = (w10008 & w17855) | (w10008 & w17856) | (w17855 & w17856);
assign v5980 = ~(w12867 | w12868);
assign w12869 = v5980;
assign w12870 = (w8795 & w17634) | (w8795 & w17635) | (w17634 & w17635);
assign v5981 = ~(w12822 | w12861);
assign w12871 = v5981;
assign v5982 = ~(w12847 | w12850);
assign w12872 = v5982;
assign w12873 = (~w12700 & ~w12702) | (~w12700 & w16952) | (~w12702 & w16952);
assign w12874 = (~w12731 & ~w12733) | (~w12731 & w16777) | (~w12733 & w16777);
assign w12875 = (~w12829 & ~w12831) | (~w12829 & w16778) | (~w12831 & w16778);
assign v5983 = ~(w12874 | w12875);
assign w12876 = v5983;
assign w12877 = w12874 & w12875;
assign v5984 = ~(w12876 | w12877);
assign w12878 = v5984;
assign w12879 = w12873 & ~w12878;
assign w12880 = ~w12873 & w12878;
assign v5985 = ~(w12879 | w12880);
assign w12881 = v5985;
assign v5986 = ~(w12717 | w12721);
assign w12882 = v5986;
assign w12883 = ~w12881 & w12882;
assign w12884 = w12881 & ~w12882;
assign v5987 = ~(w12883 | w12884);
assign w12885 = v5987;
assign v5988 = ~(w12813 | w12816);
assign w12886 = v5988;
assign w12887 = w12885 & ~w12886;
assign w12888 = ~w12885 & w12886;
assign v5989 = ~(w12887 | w12888);
assign w12889 = v5989;
assign w12890 = ~w12872 & w12889;
assign w12891 = w12872 & ~w12889;
assign v5990 = ~(w12890 | w12891);
assign w12892 = v5990;
assign v5991 = ~(w12725 | w12819);
assign w12893 = v5991;
assign w12894 = w12892 & ~w12893;
assign w12895 = ~w12892 & w12893;
assign v5992 = ~(w12894 | w12895);
assign w12896 = v5992;
assign v5993 = ~(w12855 | w12858);
assign w12897 = v5993;
assign w12898 = w12747 & ~w12750;
assign v5994 = ~(w12752 | w12898);
assign w12899 = v5994;
assign w12900 = w12769 & ~w12771;
assign v5995 = ~(w12773 | w12900);
assign w12901 = v5995;
assign v5996 = ~(w12899 | w12901);
assign w12902 = v5996;
assign w12903 = w12899 & w12901;
assign v5997 = ~(w12902 | w12903);
assign w12904 = v5997;
assign w12905 = w12757 & ~w12759;
assign v5998 = ~(w12761 | w12905);
assign w12906 = v5998;
assign w12907 = ~w12904 & w12906;
assign w12908 = w12904 & ~w12906;
assign v5999 = ~(w12907 | w12908);
assign w12909 = v5999;
assign w12910 = (~w12798 & ~w12800) | (~w12798 & w16953) | (~w12800 & w16953);
assign w12911 = (~w12766 & ~w12768) | (~w12766 & w16954) | (~w12768 & w16954);
assign v6000 = ~(w12910 | w12911);
assign w12912 = v6000;
assign w12913 = w12910 & w12911;
assign v6001 = ~(w12912 | w12913);
assign w12914 = v6001;
assign w12915 = w12909 & w12914;
assign v6002 = ~(w12909 | w12914);
assign w12916 = v6002;
assign v6003 = ~(w12915 | w12916);
assign w12917 = v6003;
assign w12918 = (~w12741 & ~w12743) | (~w12741 & w16955) | (~w12743 & w16955);
assign w12919 = pi24 & pi61;
assign w12920 = w12781 & ~w12783;
assign w12921 = (w12919 & w12920) | (w12919 & w16779) | (w12920 & w16779);
assign w12922 = ~w12920 & w16780;
assign v6004 = ~(w12921 | w12922);
assign w12923 = v6004;
assign v6005 = ~(w12790 | w12793);
assign w12924 = v6005;
assign v6006 = ~(w12792 | w12924);
assign w12925 = v6006;
assign v6007 = ~(w12923 | w12925);
assign w12926 = v6007;
assign w12927 = w12923 & w12925;
assign v6008 = ~(w12926 | w12927);
assign w12928 = v6008;
assign v6009 = ~(w12801 | w12805);
assign w12929 = v6009;
assign v6010 = ~(w12804 | w12929);
assign w12930 = v6010;
assign w12931 = w12703 & ~w12706;
assign v6011 = ~(w12708 | w12931);
assign w12932 = v6011;
assign w12933 = w12930 & ~w12932;
assign w12934 = ~w12930 & w12932;
assign v6012 = ~(w12933 | w12934);
assign w12935 = v6012;
assign w12936 = pi26 & pi59;
assign w12937 = pi27 & pi58;
assign v6013 = ~(w12936 | w12937);
assign w12938 = v6013;
assign w12939 = pi27 & pi59;
assign w12940 = w12703 & w12939;
assign v6014 = ~(w12938 | w12940);
assign w12941 = v6014;
assign w12942 = w12760 & ~w12941;
assign w12943 = ~w12760 & w12941;
assign v6015 = ~(w12942 | w12943);
assign w12944 = v6015;
assign w12945 = ~w12935 & w12944;
assign w12946 = w12935 & ~w12944;
assign v6016 = ~(w12945 | w12946);
assign w12947 = v6016;
assign v6017 = ~(w12928 | w12947);
assign w12948 = v6017;
assign w12949 = w12928 & w12947;
assign v6018 = ~(w12948 | w12949);
assign w12950 = v6018;
assign w12951 = w12918 & ~w12950;
assign w12952 = ~w12918 & w12950;
assign v6019 = ~(w12951 | w12952);
assign w12953 = v6019;
assign w12954 = w12917 & w12953;
assign v6020 = ~(w12917 | w12953);
assign w12955 = v6020;
assign v6021 = ~(w12954 | w12955);
assign w12956 = v6021;
assign w12957 = (~w12839 & ~w12841) | (~w12839 & w17209) | (~w12841 & w17209);
assign w12958 = pi33 & pi52;
assign w12959 = pi34 & pi51;
assign v6022 = ~(w12958 | w12959);
assign w12960 = v6022;
assign w12961 = pi34 & pi52;
assign w12962 = w12757 & w12961;
assign v6023 = ~(w12960 | w12962);
assign w12963 = v6023;
assign w12964 = w12707 & ~w12963;
assign w12965 = ~w12707 & w12963;
assign v6024 = ~(w12964 | w12965);
assign w12966 = v6024;
assign w12967 = pi35 & pi50;
assign w12968 = pi28 & pi57;
assign w12969 = pi22 & pi63;
assign v6025 = ~(w12968 | w12969);
assign w12970 = v6025;
assign w12971 = w12968 & w12969;
assign v6026 = ~(w12970 | w12971);
assign w12972 = v6026;
assign w12973 = w12967 & ~w12972;
assign w12974 = ~w12967 & w12972;
assign v6027 = ~(w12973 | w12974);
assign w12975 = v6027;
assign v6028 = ~(w12966 | w12975);
assign w12976 = v6028;
assign w12977 = w12966 & w12975;
assign v6029 = ~(w12976 | w12977);
assign w12978 = v6029;
assign w12979 = pi39 & pi46;
assign w12980 = pi40 & pi45;
assign v6030 = ~(w12784 | w12980);
assign w12981 = v6030;
assign w12982 = pi41 & pi45;
assign w12983 = w12521 & w12982;
assign v6031 = ~(w12981 | w12983);
assign w12984 = v6031;
assign w12985 = w12979 & ~w12984;
assign w12986 = ~w12979 & w12984;
assign v6032 = ~(w12985 | w12986);
assign w12987 = v6032;
assign w12988 = w12978 & ~w12987;
assign w12989 = ~w12978 & w12987;
assign v6033 = ~(w12988 | w12989);
assign w12990 = v6033;
assign w12991 = pi37 & pi48;
assign w12992 = pi38 & pi47;
assign v6034 = ~(w12991 | w12992);
assign w12993 = v6034;
assign w12994 = pi38 & pi48;
assign w12995 = w12801 & w12994;
assign v6035 = ~(w12993 | w12995);
assign w12996 = v6035;
assign w12997 = w12772 & ~w12996;
assign w12998 = ~w12772 & w12996;
assign v6036 = ~(w12997 | w12998);
assign w12999 = v6036;
assign w13000 = ~pi42 & pi43;
assign w13001 = w12751 & ~w13000;
assign w13002 = ~w12751 & w13000;
assign v6037 = ~(w13001 | w13002);
assign w13003 = v6037;
assign v6038 = ~(w12999 | w13003);
assign w13004 = v6038;
assign w13005 = w12999 & w13003;
assign v6039 = ~(w13004 | w13005);
assign w13006 = v6039;
assign w13007 = pi29 & pi56;
assign w13008 = pi30 & pi55;
assign w13009 = pi31 & pi54;
assign v6040 = ~(w13008 | w13009);
assign w13010 = v6040;
assign w13011 = pi31 & pi55;
assign w13012 = w12803 & w13011;
assign v6041 = ~(w13010 | w13012);
assign w13013 = v6041;
assign w13014 = w13007 & ~w13013;
assign w13015 = ~w13007 & w13013;
assign v6042 = ~(w13014 | w13015);
assign w13016 = v6042;
assign w13017 = w13006 & ~w13016;
assign w13018 = ~w13006 & w13016;
assign v6043 = ~(w13017 | w13018);
assign w13019 = v6043;
assign w13020 = w12990 & w13019;
assign v6044 = ~(w12990 | w13019);
assign w13021 = v6044;
assign v6045 = ~(w13020 | w13021);
assign w13022 = v6045;
assign w13023 = ~w12957 & w13022;
assign w13024 = w12957 & ~w13022;
assign v6046 = ~(w13023 | w13024);
assign w13025 = v6046;
assign v6047 = ~(w12956 | w13025);
assign w13026 = v6047;
assign w13027 = w12956 & w13025;
assign v6048 = ~(w13026 | w13027);
assign w13028 = v6048;
assign w13029 = ~w12897 & w13028;
assign w13030 = w12897 & ~w13028;
assign v6049 = ~(w13029 | w13030);
assign w13031 = v6049;
assign w13032 = w12896 & w13031;
assign v6050 = ~(w12896 | w13031);
assign w13033 = v6050;
assign v6051 = ~(w13032 | w13033);
assign w13034 = v6051;
assign w13035 = ~w12871 & w13034;
assign w13036 = w12871 & ~w13034;
assign v6052 = ~(w13035 | w13036);
assign w13037 = v6052;
assign w13038 = w12870 & w13037;
assign v6053 = ~(w12870 | w13037);
assign w13039 = v6053;
assign v6054 = ~(w13038 | w13039);
assign w13040 = v6054;
assign v6055 = ~(w12864 | w13036);
assign w13041 = v6055;
assign w13042 = (~w8795 & w17636) | (~w8795 & w17637) | (w17636 & w17637);
assign v6056 = ~(w13029 | w13032);
assign w13043 = v6056;
assign w13044 = (~w12902 & ~w12904) | (~w12902 & w17210) | (~w12904 & w17210);
assign w13045 = (~w12921 & ~w12923) | (~w12921 & w16956) | (~w12923 & w16956);
assign w13046 = pi25 & pi61;
assign w13047 = pi24 & pi62;
assign v6057 = ~(w13046 | w13047);
assign w13048 = v6057;
assign w13049 = pi25 & pi62;
assign w13050 = w12919 & w13049;
assign v6058 = ~(w13048 | w13050);
assign w13051 = v6058;
assign w13052 = (pi43 & w12751) | (pi43 & w16957) | (w12751 & w16957);
assign w13053 = w13051 & w13052;
assign v6059 = ~(w13051 | w13052);
assign w13054 = v6059;
assign v6060 = ~(w13053 | w13054);
assign w13055 = v6060;
assign w13056 = ~w13045 & w13055;
assign w13057 = w13045 & ~w13055;
assign v6061 = ~(w13056 | w13057);
assign w13058 = v6061;
assign w13059 = w13044 & ~w13058;
assign w13060 = ~w13044 & w13058;
assign v6062 = ~(w13059 | w13060);
assign w13061 = v6062;
assign w13062 = (w13061 & w12952) | (w13061 & w17211) | (w12952 & w17211);
assign w13063 = ~w12952 & w17212;
assign v6063 = ~(w13062 | w13063);
assign w13064 = v6063;
assign v6064 = ~(w13020 | w13023);
assign w13065 = v6064;
assign w13066 = w13064 & ~w13065;
assign w13067 = ~w13064 & w13065;
assign v6065 = ~(w13066 | w13067);
assign w13068 = v6065;
assign v6066 = ~(w12954 | w13027);
assign w13069 = v6066;
assign v6067 = ~(w12884 | w12887);
assign w13070 = v6067;
assign v6068 = ~(w13069 | w13070);
assign w13071 = v6068;
assign w13072 = w13069 & w13070;
assign v6069 = ~(w13071 | w13072);
assign w13073 = v6069;
assign w13074 = w13068 & w13073;
assign v6070 = ~(w13068 | w13073);
assign w13075 = v6070;
assign v6071 = ~(w13074 | w13075);
assign w13076 = v6071;
assign v6072 = ~(w12890 | w12894);
assign w13077 = v6072;
assign w13078 = (~w12912 & ~w12914) | (~w12912 & w17213) | (~w12914 & w17213);
assign w13079 = pi23 & pi63;
assign w13080 = pi36 & pi50;
assign w13081 = pi37 & pi49;
assign v6073 = ~(w13080 | w13081);
assign w13082 = v6073;
assign w13083 = pi37 & pi50;
assign w13084 = w12772 & w13083;
assign v6074 = ~(w13082 | w13084);
assign w13085 = v6074;
assign w13086 = w13079 & ~w13085;
assign w13087 = ~w13079 & w13085;
assign v6075 = ~(w13086 | w13087);
assign w13088 = v6075;
assign w13089 = pi33 & pi53;
assign w13090 = pi35 & pi51;
assign v6076 = ~(w12961 | w13090);
assign w13091 = v6076;
assign w13092 = pi35 & pi52;
assign w13093 = w12959 & w13092;
assign v6077 = ~(w13091 | w13093);
assign w13094 = v6077;
assign w13095 = w13089 & ~w13094;
assign w13096 = ~w13089 & w13094;
assign v6078 = ~(w13095 | w13096);
assign w13097 = v6078;
assign v6079 = ~(w13088 | w13097);
assign w13098 = v6079;
assign w13099 = w13088 & w13097;
assign v6080 = ~(w13098 | w13099);
assign w13100 = v6080;
assign w13101 = pi29 & pi57;
assign v6081 = ~(w13011 | w13101);
assign w13102 = v6081;
assign w13103 = w13011 & w13101;
assign v6082 = ~(w13102 | w13103);
assign w13104 = v6082;
assign w13105 = w12994 & ~w13104;
assign w13106 = ~w12994 & w13104;
assign v6083 = ~(w13105 | w13106);
assign w13107 = v6083;
assign w13108 = w13100 & ~w13107;
assign w13109 = ~w13100 & w13107;
assign v6084 = ~(w13108 | w13109);
assign w13110 = v6084;
assign w13111 = pi26 & pi60;
assign w13112 = pi28 & pi58;
assign v6085 = ~(w12939 | w13112);
assign w13113 = v6085;
assign w13114 = pi28 & pi59;
assign w13115 = w12937 & w13114;
assign v6086 = ~(w13113 | w13115);
assign w13116 = v6086;
assign w13117 = w13111 & ~w13116;
assign w13118 = ~w13111 & w13116;
assign v6087 = ~(w13117 | w13118);
assign w13119 = v6087;
assign w13120 = pi42 & pi44;
assign w13121 = pi32 & pi54;
assign v6088 = ~(w13120 | w13121);
assign w13122 = v6088;
assign w13123 = w13120 & w13121;
assign v6089 = ~(w13122 | w13123);
assign w13124 = v6089;
assign w13125 = w12982 & ~w13124;
assign w13126 = ~w12982 & w13124;
assign v6090 = ~(w13125 | w13126);
assign w13127 = v6090;
assign v6091 = ~(w13119 | w13127);
assign w13128 = v6091;
assign w13129 = w13119 & w13127;
assign v6092 = ~(w13128 | w13129);
assign w13130 = v6092;
assign w13131 = pi30 & pi56;
assign w13132 = pi40 & pi46;
assign w13133 = pi39 & pi47;
assign v6093 = ~(w13132 | w13133);
assign w13134 = v6093;
assign w13135 = pi40 & pi47;
assign w13136 = w12979 & w13135;
assign v6094 = ~(w13134 | w13136);
assign w13137 = v6094;
assign w13138 = w13131 & ~w13137;
assign w13139 = ~w13131 & w13137;
assign v6095 = ~(w13138 | w13139);
assign w13140 = v6095;
assign w13141 = w13130 & ~w13140;
assign w13142 = ~w13130 & w13140;
assign v6096 = ~(w13141 | w13142);
assign w13143 = v6096;
assign w13144 = w13110 & w13143;
assign v6097 = ~(w13110 | w13143);
assign w13145 = v6097;
assign v6098 = ~(w13144 | w13145);
assign w13146 = v6098;
assign w13147 = ~w13078 & w13146;
assign w13148 = w13078 & ~w13146;
assign v6099 = ~(w13147 | w13148);
assign w13149 = v6099;
assign v6100 = ~(w13004 | w13017);
assign w13150 = v6100;
assign w13151 = (~w12933 & ~w12935) | (~w12933 & w17214) | (~w12935 & w17214);
assign w13152 = (~w12976 & ~w12978) | (~w12976 & w16958) | (~w12978 & w16958);
assign v6101 = ~(w13151 | w13152);
assign w13153 = v6101;
assign w13154 = w13151 & w13152;
assign v6102 = ~(w13153 | w13154);
assign w13155 = v6102;
assign w13156 = w13150 & ~w13155;
assign w13157 = ~w13150 & w13155;
assign v6103 = ~(w13156 | w13157);
assign w13158 = v6103;
assign w13159 = (~w12876 & ~w12878) | (~w12876 & w16959) | (~w12878 & w16959);
assign w13160 = w12979 & ~w12981;
assign v6104 = ~(w12983 | w13160);
assign w13161 = v6104;
assign w13162 = w13007 & ~w13010;
assign v6105 = ~(w13012 | w13162);
assign w13163 = v6105;
assign v6106 = ~(w13161 | w13163);
assign w13164 = v6106;
assign w13165 = w13161 & w13163;
assign v6107 = ~(w13164 | w13165);
assign w13166 = v6107;
assign w13167 = w12772 & ~w12993;
assign v6108 = ~(w12995 | w13167);
assign w13168 = v6108;
assign w13169 = ~w13166 & w13168;
assign w13170 = w13166 & ~w13168;
assign v6109 = ~(w13169 | w13170);
assign w13171 = v6109;
assign w13172 = w12760 & ~w12938;
assign v6110 = ~(w12940 | w13172);
assign w13173 = v6110;
assign w13174 = w12707 & ~w12960;
assign v6111 = ~(w12962 | w13174);
assign w13175 = v6111;
assign v6112 = ~(w13173 | w13175);
assign w13176 = v6112;
assign w13177 = w13173 & w13175;
assign v6113 = ~(w13176 | w13177);
assign w13178 = v6113;
assign v6114 = ~(w12967 | w12971);
assign w13179 = v6114;
assign v6115 = ~(w12970 | w13179);
assign w13180 = v6115;
assign v6116 = ~(w13178 | w13180);
assign w13181 = v6116;
assign w13182 = w13178 & w13180;
assign v6117 = ~(w13181 | w13182);
assign w13183 = v6117;
assign w13184 = w13171 & w13183;
assign v6118 = ~(w13171 | w13183);
assign w13185 = v6118;
assign v6119 = ~(w13184 | w13185);
assign w13186 = v6119;
assign w13187 = ~w13159 & w13186;
assign w13188 = w13159 & ~w13186;
assign v6120 = ~(w13187 | w13188);
assign w13189 = v6120;
assign w13190 = w13158 & w13189;
assign v6121 = ~(w13158 | w13189);
assign w13191 = v6121;
assign v6122 = ~(w13190 | w13191);
assign w13192 = v6122;
assign w13193 = w13149 & w13192;
assign v6123 = ~(w13149 | w13192);
assign w13194 = v6123;
assign v6124 = ~(w13193 | w13194);
assign w13195 = v6124;
assign w13196 = ~w13077 & w13195;
assign w13197 = w13077 & ~w13195;
assign v6125 = ~(w13196 | w13197);
assign w13198 = v6125;
assign w13199 = w13076 & w13198;
assign v6126 = ~(w13076 | w13198);
assign w13200 = v6126;
assign v6127 = ~(w13199 | w13200);
assign w13201 = v6127;
assign w13202 = ~w13043 & w13201;
assign w13203 = w13043 & ~w13201;
assign v6128 = ~(w13202 | w13203);
assign w13204 = v6128;
assign w13205 = w13042 & w13204;
assign v6129 = ~(w13042 | w13204);
assign w13206 = v6129;
assign v6130 = ~(w13205 | w13206);
assign w13207 = v6130;
assign v6131 = ~(w13035 | w13202);
assign w13208 = v6131;
assign v6132 = ~(w13196 | w13199);
assign w13209 = v6132;
assign v6133 = ~(w13144 | w13147);
assign w13210 = v6133;
assign v6134 = ~(w13128 | w13141);
assign w13211 = v6134;
assign w13212 = (~w13164 & ~w13166) | (~w13164 & w17215) | (~w13166 & w17215);
assign w13213 = (~w13098 & ~w13100) | (~w13098 & w16960) | (~w13100 & w16960);
assign v6135 = ~(w13212 | w13213);
assign w13214 = v6135;
assign w13215 = w13212 & w13213;
assign v6136 = ~(w13214 | w13215);
assign w13216 = v6136;
assign w13217 = w13211 & ~w13216;
assign w13218 = ~w13211 & w13216;
assign v6137 = ~(w13217 | w13218);
assign w13219 = v6137;
assign w13220 = ~w13210 & w13219;
assign w13221 = w13210 & ~w13219;
assign v6138 = ~(w13220 | w13221);
assign w13222 = v6138;
assign v6139 = ~(w13062 | w13066);
assign w13223 = v6139;
assign w13224 = ~w13222 & w13223;
assign w13225 = w13222 & ~w13223;
assign v6140 = ~(w13224 | w13225);
assign w13226 = v6140;
assign v6141 = ~(w13071 | w13074);
assign w13227 = v6141;
assign w13228 = ~w13226 & w13227;
assign w13229 = w13226 & ~w13227;
assign v6142 = ~(w13228 | w13229);
assign w13230 = v6142;
assign v6143 = ~(w13190 | w13193);
assign w13231 = v6143;
assign w13232 = (~w13176 & ~w13178) | (~w13176 & w17216) | (~w13178 & w17216);
assign w13233 = ~pi43 & pi44;
assign w13234 = w13049 & ~w13233;
assign w13235 = ~w13049 & w13233;
assign v6144 = ~(w13234 | w13235);
assign w13236 = v6144;
assign w13237 = pi31 & pi56;
assign w13238 = pi33 & pi54;
assign v6145 = ~(w13237 | w13238);
assign w13239 = v6145;
assign w13240 = w13237 & w13238;
assign v6146 = ~(w13239 | w13240);
assign w13241 = v6146;
assign w13242 = w13135 & ~w13241;
assign w13243 = ~w13135 & w13241;
assign v6147 = ~(w13242 | w13243);
assign w13244 = v6147;
assign v6148 = ~(w13236 | w13244);
assign w13245 = v6148;
assign w13246 = w13236 & w13244;
assign v6149 = ~(w13245 | w13246);
assign w13247 = v6149;
assign w13248 = w13232 & ~w13247;
assign w13249 = ~w13232 & w13247;
assign v6150 = ~(w13248 | w13249);
assign w13250 = v6150;
assign w13251 = pi24 & pi63;
assign w13252 = pi26 & pi61;
assign w13253 = pi27 & pi60;
assign v6151 = ~(w13252 | w13253);
assign w13254 = v6151;
assign w13255 = pi27 & pi61;
assign w13256 = w13111 & w13255;
assign v6152 = ~(w13254 | w13256);
assign w13257 = v6152;
assign w13258 = w13251 & ~w13257;
assign w13259 = ~w13251 & w13257;
assign v6153 = ~(w13258 | w13259);
assign w13260 = v6153;
assign w13261 = pi38 & pi49;
assign w13262 = pi39 & pi48;
assign v6154 = ~(w13261 | w13262);
assign w13263 = v6154;
assign w13264 = pi39 & pi49;
assign w13265 = w12994 & w13264;
assign v6155 = ~(w13263 | w13265);
assign w13266 = v6155;
assign w13267 = w13083 & ~w13266;
assign w13268 = ~w13083 & w13266;
assign v6156 = ~(w13267 | w13268);
assign w13269 = v6156;
assign v6157 = ~(w13260 | w13269);
assign w13270 = v6157;
assign w13271 = w13260 & w13269;
assign v6158 = ~(w13270 | w13271);
assign w13272 = v6158;
assign w13273 = pi32 & pi55;
assign w13274 = pi41 & pi46;
assign w13275 = pi42 & pi45;
assign v6159 = ~(w13274 | w13275);
assign w13276 = v6159;
assign w13277 = pi42 & pi46;
assign w13278 = w12982 & w13277;
assign v6160 = ~(w13276 | w13278);
assign w13279 = v6160;
assign w13280 = w13273 & ~w13279;
assign w13281 = ~w13273 & w13279;
assign v6161 = ~(w13280 | w13281);
assign w13282 = v6161;
assign w13283 = w13272 & ~w13282;
assign w13284 = ~w13272 & w13282;
assign v6162 = ~(w13283 | w13284);
assign w13285 = v6162;
assign v6163 = ~(w13250 | w13285);
assign w13286 = v6163;
assign w13287 = w13250 & w13285;
assign v6164 = ~(w13286 | w13287);
assign w13288 = v6164;
assign w13289 = (~w13050 & ~w13051) | (~w13050 & w16961) | (~w13051 & w16961);
assign w13290 = pi30 & pi57;
assign w13291 = pi34 & pi53;
assign v6165 = ~(w13290 | w13291);
assign w13292 = v6165;
assign w13293 = w13290 & w13291;
assign v6166 = ~(w13292 | w13293);
assign w13294 = v6166;
assign w13295 = w13114 & ~w13294;
assign w13296 = ~w13114 & w13294;
assign v6167 = ~(w13295 | w13296);
assign w13297 = v6167;
assign v6168 = ~(w13289 | w13297);
assign w13298 = v6168;
assign w13299 = w13289 & w13297;
assign v6169 = ~(w13298 | w13299);
assign w13300 = v6169;
assign w13301 = pi29 & pi58;
assign w13302 = pi36 & pi51;
assign v6170 = ~(w13301 | w13302);
assign w13303 = v6170;
assign w13304 = w13301 & w13302;
assign v6171 = ~(w13303 | w13304);
assign w13305 = v6171;
assign w13306 = w13092 & ~w13305;
assign w13307 = ~w13092 & w13305;
assign v6172 = ~(w13306 | w13307);
assign w13308 = v6172;
assign w13309 = w13300 & ~w13308;
assign w13310 = ~w13300 & w13308;
assign v6173 = ~(w13309 | w13310);
assign w13311 = v6173;
assign w13312 = w13288 & w13311;
assign v6174 = ~(w13288 | w13311);
assign w13313 = v6174;
assign v6175 = ~(w13312 | w13313);
assign w13314 = v6175;
assign w13315 = ~w13231 & w13314;
assign w13316 = w13231 & ~w13314;
assign v6176 = ~(w13315 | w13316);
assign w13317 = v6176;
assign w13318 = (~w13056 & ~w13058) | (~w13056 & w17217) | (~w13058 & w17217);
assign v6177 = ~(w12982 | w13123);
assign w13319 = v6177;
assign v6178 = ~(w13122 | w13319);
assign w13320 = v6178;
assign w13321 = w13131 & ~w13134;
assign v6179 = ~(w13136 | w13321);
assign w13322 = v6179;
assign w13323 = w13320 & ~w13322;
assign w13324 = ~w13320 & w13322;
assign v6180 = ~(w13323 | w13324);
assign w13325 = v6180;
assign v6181 = ~(w12994 | w13103);
assign w13326 = v6181;
assign v6182 = ~(w13102 | w13326);
assign w13327 = v6182;
assign v6183 = ~(w13325 | w13327);
assign w13328 = v6183;
assign w13329 = w13325 & w13327;
assign v6184 = ~(w13328 | w13329);
assign w13330 = v6184;
assign w13331 = w13089 & ~w13091;
assign v6185 = ~(w13093 | w13331);
assign w13332 = v6185;
assign w13333 = w13111 & ~w13113;
assign v6186 = ~(w13115 | w13333);
assign w13334 = v6186;
assign v6187 = ~(w13332 | w13334);
assign w13335 = v6187;
assign w13336 = w13332 & w13334;
assign v6188 = ~(w13335 | w13336);
assign w13337 = v6188;
assign w13338 = w13079 & ~w13082;
assign v6189 = ~(w13084 | w13338);
assign w13339 = v6189;
assign w13340 = ~w13337 & w13339;
assign w13341 = w13337 & ~w13339;
assign v6190 = ~(w13340 | w13341);
assign w13342 = v6190;
assign w13343 = w13330 & w13342;
assign v6191 = ~(w13330 | w13342);
assign w13344 = v6191;
assign v6192 = ~(w13343 | w13344);
assign w13345 = v6192;
assign w13346 = ~w13318 & w13345;
assign w13347 = w13318 & ~w13345;
assign v6193 = ~(w13346 | w13347);
assign w13348 = v6193;
assign v6194 = ~(w13184 | w13187);
assign w13349 = v6194;
assign w13350 = (~w13153 & ~w13155) | (~w13153 & w17218) | (~w13155 & w17218);
assign v6195 = ~(w13349 | w13350);
assign w13351 = v6195;
assign w13352 = w13349 & w13350;
assign v6196 = ~(w13351 | w13352);
assign w13353 = v6196;
assign w13354 = w13348 & w13353;
assign v6197 = ~(w13348 | w13353);
assign w13355 = v6197;
assign v6198 = ~(w13354 | w13355);
assign w13356 = v6198;
assign w13357 = w13317 & w13356;
assign v6199 = ~(w13317 | w13356);
assign w13358 = v6199;
assign v6200 = ~(w13357 | w13358);
assign w13359 = v6200;
assign v6201 = ~(w13230 | w13359);
assign w13360 = v6201;
assign w13361 = w13230 & w13359;
assign v6202 = ~(w13360 | w13361);
assign w13362 = v6202;
assign w13363 = w13209 & ~w13362;
assign w13364 = ~w13209 & w13362;
assign v6203 = ~(w13363 | w13364);
assign w13365 = v6203;
assign w13366 = (~w10008 & w17857) | (~w10008 & w17858) | (w17857 & w17858);
assign w13367 = (w10008 & w17859) | (w10008 & w17860) | (w17859 & w17860);
assign v6204 = ~(w13366 | w13367);
assign w13368 = v6204;
assign v6205 = ~(w13229 | w13361);
assign w13369 = v6205;
assign v6206 = ~(w13315 | w13357);
assign w13370 = v6206;
assign w13371 = (~w13351 & ~w13353) | (~w13351 & w17219) | (~w13353 & w17219);
assign v6207 = ~(w13270 | w13283);
assign w13372 = v6207;
assign w13373 = (~w13335 & ~w13337) | (~w13335 & w17220) | (~w13337 & w17220);
assign w13374 = (~w13298 & ~w13300) | (~w13298 & w16962) | (~w13300 & w16962);
assign v6208 = ~(w13373 | w13374);
assign w13375 = v6208;
assign w13376 = w13373 & w13374;
assign v6209 = ~(w13375 | w13376);
assign w13377 = v6209;
assign w13378 = w13372 & ~w13377;
assign w13379 = ~w13372 & w13377;
assign v6210 = ~(w13378 | w13379);
assign w13380 = v6210;
assign v6211 = ~(w13287 | w13312);
assign w13381 = v6211;
assign w13382 = ~w13380 & w13381;
assign w13383 = w13380 & ~w13381;
assign v6212 = ~(w13382 | w13383);
assign w13384 = v6212;
assign w13385 = ~w13371 & w13384;
assign w13386 = w13371 & ~w13384;
assign v6213 = ~(w13385 | w13386);
assign w13387 = v6213;
assign w13388 = ~w13370 & w13387;
assign w13389 = w13370 & ~w13387;
assign v6214 = ~(w13388 | w13389);
assign w13390 = v6214;
assign v6215 = ~(w13114 | w13293);
assign w13391 = v6215;
assign v6216 = ~(w13292 | w13391);
assign w13392 = v6216;
assign w13393 = w13251 & ~w13254;
assign v6217 = ~(w13256 | w13393);
assign w13394 = v6217;
assign w13395 = w13392 & ~w13394;
assign w13396 = ~w13392 & w13394;
assign v6218 = ~(w13395 | w13396);
assign w13397 = v6218;
assign w13398 = w13083 & ~w13263;
assign v6219 = ~(w13265 | w13398);
assign w13399 = v6219;
assign w13400 = ~w13397 & w13399;
assign w13401 = w13397 & ~w13399;
assign v6220 = ~(w13400 | w13401);
assign w13402 = v6220;
assign v6221 = ~(w13135 | w13240);
assign w13403 = v6221;
assign v6222 = ~(w13239 | w13403);
assign w13404 = v6222;
assign v6223 = ~(w13092 | w13304);
assign w13405 = v6223;
assign v6224 = ~(w13303 | w13405);
assign w13406 = v6224;
assign w13407 = w13404 & w13406;
assign v6225 = ~(w13404 | w13406);
assign w13408 = v6225;
assign v6226 = ~(w13407 | w13408);
assign w13409 = v6226;
assign w13410 = pi43 & pi45;
assign w13411 = pi33 & pi55;
assign w13412 = pi34 & pi54;
assign v6227 = ~(w13411 | w13412);
assign w13413 = v6227;
assign w13414 = pi34 & pi55;
assign w13415 = w13238 & w13414;
assign v6228 = ~(w13413 | w13415);
assign w13416 = v6228;
assign w13417 = w13410 & ~w13416;
assign w13418 = ~w13410 & w13416;
assign v6229 = ~(w13417 | w13418);
assign w13419 = v6229;
assign w13420 = ~w13409 & w13419;
assign w13421 = w13409 & ~w13419;
assign v6230 = ~(w13420 | w13421);
assign w13422 = v6230;
assign v6231 = ~(w13245 | w13249);
assign w13423 = v6231;
assign w13424 = w13422 & ~w13423;
assign w13425 = ~w13422 & w13423;
assign v6232 = ~(w13424 | w13425);
assign w13426 = v6232;
assign w13427 = w13402 & w13426;
assign v6233 = ~(w13402 | w13426);
assign w13428 = v6233;
assign v6234 = ~(w13427 | w13428);
assign w13429 = v6234;
assign w13430 = (~w13343 & ~w13345) | (~w13343 & w17221) | (~w13345 & w17221);
assign w13431 = (~w13214 & ~w13216) | (~w13214 & w17222) | (~w13216 & w17222);
assign v6235 = ~(w13430 | w13431);
assign w13432 = v6235;
assign w13433 = w13430 & w13431;
assign v6236 = ~(w13432 | w13433);
assign w13434 = v6236;
assign w13435 = w13429 & w13434;
assign v6237 = ~(w13429 | w13434);
assign w13436 = v6237;
assign v6238 = ~(w13435 | w13436);
assign w13437 = v6238;
assign v6239 = ~(w13220 | w13225);
assign w13438 = v6239;
assign w13439 = pi26 & pi62;
assign w13440 = pi28 & pi60;
assign v6240 = ~(w13255 | w13440);
assign w13441 = v6240;
assign w13442 = pi28 & pi61;
assign w13443 = w13253 & w13442;
assign v6241 = ~(w13441 | w13443);
assign w13444 = v6241;
assign w13445 = w13439 & ~w13444;
assign w13446 = ~w13439 & w13444;
assign v6242 = ~(w13445 | w13446);
assign w13447 = v6242;
assign w13448 = pi31 & pi57;
assign w13449 = pi41 & pi47;
assign v6243 = ~(w13277 | w13449);
assign w13450 = v6243;
assign w13451 = pi42 & pi47;
assign w13452 = w13274 & w13451;
assign v6244 = ~(w13450 | w13452);
assign w13453 = v6244;
assign w13454 = w13448 & ~w13453;
assign w13455 = ~w13448 & w13453;
assign v6245 = ~(w13454 | w13455);
assign w13456 = v6245;
assign v6246 = ~(w13447 | w13456);
assign w13457 = v6246;
assign w13458 = w13447 & w13456;
assign v6247 = ~(w13457 | w13458);
assign w13459 = v6247;
assign w13460 = pi35 & pi53;
assign w13461 = pi37 & pi51;
assign w13462 = pi36 & pi52;
assign v6248 = ~(w13461 | w13462);
assign w13463 = v6248;
assign w13464 = pi37 & pi52;
assign w13465 = w13302 & w13464;
assign v6249 = ~(w13463 | w13465);
assign w13466 = v6249;
assign w13467 = w13460 & ~w13466;
assign w13468 = ~w13460 & w13466;
assign v6250 = ~(w13467 | w13468);
assign w13469 = v6250;
assign w13470 = w13459 & ~w13469;
assign w13471 = ~w13459 & w13469;
assign v6251 = ~(w13470 | w13471);
assign w13472 = v6251;
assign w13473 = (~w13323 & ~w13325) | (~w13323 & w17223) | (~w13325 & w17223);
assign w13474 = pi29 & pi59;
assign w13475 = pi38 & pi50;
assign v6252 = ~(w13264 | w13475);
assign w13476 = v6252;
assign w13477 = pi39 & pi50;
assign w13478 = w13261 & w13477;
assign v6253 = ~(w13476 | w13478);
assign w13479 = v6253;
assign w13480 = w13474 & ~w13479;
assign w13481 = ~w13474 & w13479;
assign v6254 = ~(w13480 | w13481);
assign w13482 = v6254;
assign w13483 = pi40 & pi48;
assign w13484 = pi30 & pi58;
assign w13485 = pi32 & pi56;
assign v6255 = ~(w13484 | w13485);
assign w13486 = v6255;
assign w13487 = w13484 & w13485;
assign v6256 = ~(w13486 | w13487);
assign w13488 = v6256;
assign w13489 = w13483 & ~w13488;
assign w13490 = ~w13483 & w13488;
assign v6257 = ~(w13489 | w13490);
assign w13491 = v6257;
assign v6258 = ~(w13482 | w13491);
assign w13492 = v6258;
assign w13493 = w13482 & w13491;
assign v6259 = ~(w13492 | w13493);
assign w13494 = v6259;
assign w13495 = w13473 & ~w13494;
assign w13496 = ~w13473 & w13494;
assign v6260 = ~(w13495 | w13496);
assign w13497 = v6260;
assign w13498 = pi25 & pi63;
assign v6261 = ~(pi43 | w13049);
assign w13499 = v6261;
assign w13500 = pi44 & ~w13499;
assign w13501 = w13498 & w13500;
assign v6262 = ~(w13498 | w13500);
assign w13502 = v6262;
assign v6263 = ~(w13501 | w13502);
assign w13503 = v6263;
assign w13504 = w13273 & ~w13276;
assign v6264 = ~(w13278 | w13504);
assign w13505 = v6264;
assign w13506 = ~w13503 & w13505;
assign w13507 = w13503 & ~w13505;
assign v6265 = ~(w13506 | w13507);
assign w13508 = v6265;
assign w13509 = w13497 & w13508;
assign v6266 = ~(w13497 | w13508);
assign w13510 = v6266;
assign v6267 = ~(w13509 | w13510);
assign w13511 = v6267;
assign w13512 = w13472 & w13511;
assign v6268 = ~(w13472 | w13511);
assign w13513 = v6268;
assign v6269 = ~(w13512 | w13513);
assign w13514 = v6269;
assign w13515 = ~w13438 & w13514;
assign w13516 = w13438 & ~w13514;
assign v6270 = ~(w13515 | w13516);
assign w13517 = v6270;
assign w13518 = w13437 & w13517;
assign v6271 = ~(w13437 | w13517);
assign w13519 = v6271;
assign v6272 = ~(w13518 | w13519);
assign w13520 = v6272;
assign v6273 = ~(w13390 | w13520);
assign w13521 = v6273;
assign w13522 = w13390 & w13520;
assign v6274 = ~(w13521 | w13522);
assign w13523 = v6274;
assign w13524 = w13369 & ~w13523;
assign w13525 = ~w13369 & w13523;
assign v6275 = ~(w13524 | w13525);
assign w13526 = v6275;
assign w13527 = (w11122 & w17638) | (w11122 & w17639) | (w17638 & w17639);
assign w13528 = (~w11122 & w17640) | (~w11122 & w17641) | (w17640 & w17641);
assign v6276 = ~(w13527 | w13528);
assign w13529 = v6276;
assign v6277 = ~(w13388 | w13522);
assign w13530 = v6277;
assign v6278 = ~(w13407 | w13421);
assign w13531 = v6278;
assign w13532 = (~w13395 & ~w13397) | (~w13395 & w17224) | (~w13397 & w17224);
assign v6279 = ~(w13501 | w13507);
assign w13533 = v6279;
assign v6280 = ~(w13532 | w13533);
assign w13534 = v6280;
assign w13535 = w13532 & w13533;
assign v6281 = ~(w13534 | w13535);
assign w13536 = v6281;
assign w13537 = w13531 & ~w13536;
assign w13538 = ~w13531 & w13536;
assign v6282 = ~(w13537 | w13538);
assign w13539 = v6282;
assign w13540 = (~w13375 & ~w13377) | (~w13375 & w17225) | (~w13377 & w17225);
assign w13541 = ~w13539 & w13540;
assign w13542 = w13539 & ~w13540;
assign v6283 = ~(w13541 | w13542);
assign w13543 = v6283;
assign v6284 = ~(w13424 | w13427);
assign w13544 = v6284;
assign w13545 = w13543 & ~w13544;
assign w13546 = ~w13543 & w13544;
assign v6285 = ~(w13545 | w13546);
assign w13547 = v6285;
assign v6286 = ~(w13383 | w13385);
assign w13548 = v6286;
assign w13549 = w13439 & ~w13441;
assign v6287 = ~(w13443 | w13549);
assign w13550 = v6287;
assign w13551 = w13460 & ~w13463;
assign v6288 = ~(w13465 | w13551);
assign w13552 = v6288;
assign v6289 = ~(w13550 | w13552);
assign w13553 = v6289;
assign w13554 = w13550 & w13552;
assign v6290 = ~(w13553 | w13554);
assign w13555 = v6290;
assign v6291 = ~(w13483 | w13487);
assign w13556 = v6291;
assign v6292 = ~(w13486 | w13556);
assign w13557 = v6292;
assign v6293 = ~(w13555 | w13557);
assign w13558 = v6293;
assign w13559 = w13555 & w13557;
assign v6294 = ~(w13558 | w13559);
assign w13560 = v6294;
assign w13561 = pi29 & pi60;
assign v6295 = ~(w13442 | w13561);
assign w13562 = v6295;
assign w13563 = pi29 & pi61;
assign w13564 = w13440 & w13563;
assign v6296 = ~(w13562 | w13564);
assign w13565 = v6296;
assign w13566 = w13410 & ~w13413;
assign v6297 = ~(w13415 | w13566);
assign w13567 = v6297;
assign w13568 = w13565 & ~w13567;
assign w13569 = ~w13565 & w13567;
assign v6298 = ~(w13568 | w13569);
assign w13570 = v6298;
assign w13571 = pi43 & pi46;
assign v6299 = ~(w13451 | w13571);
assign w13572 = v6299;
assign w13573 = pi43 & pi47;
assign w13574 = w13277 & w13573;
assign v6300 = ~(w13572 | w13574);
assign w13575 = v6300;
assign w13576 = w13414 & ~w13575;
assign w13577 = ~w13414 & w13575;
assign v6301 = ~(w13576 | w13577);
assign w13578 = v6301;
assign w13579 = pi27 & pi62;
assign w13580 = ~pi44 & pi45;
assign w13581 = w13579 & ~w13580;
assign w13582 = ~w13579 & w13580;
assign v6302 = ~(w13581 | w13582);
assign w13583 = v6302;
assign v6303 = ~(w13578 | w13583);
assign w13584 = v6303;
assign w13585 = w13578 & w13583;
assign v6304 = ~(w13584 | w13585);
assign w13586 = v6304;
assign w13587 = w13570 & w13586;
assign v6305 = ~(w13570 | w13586);
assign w13588 = v6305;
assign v6306 = ~(w13587 | w13588);
assign w13589 = v6306;
assign v6307 = ~(w13560 | w13589);
assign w13590 = v6307;
assign w13591 = w13560 & w13589;
assign v6308 = ~(w13590 | w13591);
assign w13592 = v6308;
assign w13593 = pi36 & pi53;
assign w13594 = pi38 & pi51;
assign v6309 = ~(w13464 | w13594);
assign w13595 = v6309;
assign w13596 = pi38 & pi52;
assign w13597 = w13461 & w13596;
assign v6310 = ~(w13595 | w13597);
assign w13598 = v6310;
assign w13599 = w13593 & ~w13598;
assign w13600 = ~w13593 & w13598;
assign v6311 = ~(w13599 | w13600);
assign w13601 = v6311;
assign w13602 = pi41 & pi48;
assign w13603 = pi33 & pi56;
assign w13604 = pi35 & pi54;
assign v6312 = ~(w13603 | w13604);
assign w13605 = v6312;
assign w13606 = w13603 & w13604;
assign v6313 = ~(w13605 | w13606);
assign w13607 = v6313;
assign w13608 = w13602 & ~w13607;
assign w13609 = ~w13602 & w13607;
assign v6314 = ~(w13608 | w13609);
assign w13610 = v6314;
assign v6315 = ~(w13601 | w13610);
assign w13611 = v6315;
assign w13612 = w13601 & w13610;
assign v6316 = ~(w13611 | w13612);
assign w13613 = v6316;
assign w13614 = pi30 & pi59;
assign w13615 = pi32 & pi57;
assign w13616 = pi31 & pi58;
assign v6317 = ~(w13615 | w13616);
assign w13617 = v6317;
assign w13618 = pi32 & pi58;
assign w13619 = w13448 & w13618;
assign v6318 = ~(w13617 | w13619);
assign w13620 = v6318;
assign w13621 = w13614 & ~w13620;
assign w13622 = ~w13614 & w13620;
assign v6319 = ~(w13621 | w13622);
assign w13623 = v6319;
assign w13624 = w13613 & ~w13623;
assign w13625 = ~w13613 & w13623;
assign v6320 = ~(w13624 | w13625);
assign w13626 = v6320;
assign w13627 = w13592 & w13626;
assign v6321 = ~(w13592 | w13626);
assign w13628 = v6321;
assign v6322 = ~(w13627 | w13628);
assign w13629 = v6322;
assign w13630 = ~w13548 & w13629;
assign w13631 = w13548 & ~w13629;
assign v6323 = ~(w13630 | w13631);
assign w13632 = v6323;
assign w13633 = w13547 & w13632;
assign v6324 = ~(w13547 | w13632);
assign w13634 = v6324;
assign v6325 = ~(w13633 | w13634);
assign w13635 = v6325;
assign v6326 = ~(w13432 | w13435);
assign w13636 = v6326;
assign v6327 = ~(w13509 | w13512);
assign w13637 = v6327;
assign w13638 = w13448 & ~w13450;
assign v6328 = ~(w13452 | w13638);
assign w13639 = v6328;
assign w13640 = w13474 & ~w13476;
assign v6329 = ~(w13478 | w13640);
assign w13641 = v6329;
assign v6330 = ~(w13639 | w13641);
assign w13642 = v6330;
assign w13643 = w13639 & w13641;
assign v6331 = ~(w13642 | w13643);
assign w13644 = v6331;
assign w13645 = pi26 & pi63;
assign w13646 = pi40 & pi49;
assign v6332 = ~(w13477 | w13646);
assign w13647 = v6332;
assign w13648 = pi40 & pi50;
assign w13649 = w13264 & w13648;
assign v6333 = ~(w13647 | w13649);
assign w13650 = v6333;
assign w13651 = w13645 & ~w13650;
assign w13652 = ~w13645 & w13650;
assign v6334 = ~(w13651 | w13652);
assign w13653 = v6334;
assign w13654 = ~w13644 & w13653;
assign w13655 = w13644 & ~w13653;
assign v6335 = ~(w13654 | w13655);
assign w13656 = v6335;
assign v6336 = ~(w13492 | w13496);
assign w13657 = v6336;
assign v6337 = ~(w13457 | w13470);
assign w13658 = v6337;
assign v6338 = ~(w13657 | w13658);
assign w13659 = v6338;
assign w13660 = w13657 & w13658;
assign v6339 = ~(w13659 | w13660);
assign w13661 = v6339;
assign v6340 = ~(w13656 | w13661);
assign w13662 = v6340;
assign w13663 = w13656 & w13661;
assign v6341 = ~(w13662 | w13663);
assign w13664 = v6341;
assign w13665 = ~w13637 & w13664;
assign w13666 = w13637 & ~w13664;
assign v6342 = ~(w13665 | w13666);
assign w13667 = v6342;
assign w13668 = ~w13636 & w13667;
assign w13669 = w13636 & ~w13667;
assign v6343 = ~(w13668 | w13669);
assign w13670 = v6343;
assign v6344 = ~(w13515 | w13518);
assign w13671 = v6344;
assign w13672 = w13670 & ~w13671;
assign w13673 = ~w13670 & w13671;
assign v6345 = ~(w13672 | w13673);
assign w13674 = v6345;
assign w13675 = w13635 & w13674;
assign v6346 = ~(w13635 | w13674);
assign w13676 = v6346;
assign v6347 = ~(w13675 | w13676);
assign w13677 = v6347;
assign w13678 = ~w13530 & w13677;
assign w13679 = w13530 & ~w13677;
assign v6348 = ~(w13678 | w13679);
assign w13680 = v6348;
assign v6349 = ~(w13363 | w13524);
assign w13681 = v6349;
assign w13682 = (~w11122 & w17642) | (~w11122 & w17643) | (w17642 & w17643);
assign w13683 = (w11122 & w17644) | (w11122 & w17645) | (w17644 & w17645);
assign v6350 = ~(w13682 | w13683);
assign w13684 = v6350;
assign v6351 = ~(w13525 | w13678);
assign w13685 = v6351;
assign v6352 = ~(w13672 | w13675);
assign w13686 = v6352;
assign v6353 = ~(w13542 | w13545);
assign w13687 = v6353;
assign v6354 = ~(w13591 | w13627);
assign w13688 = v6354;
assign v6355 = ~(pi44 | w13579);
assign w13689 = v6355;
assign w13690 = pi45 & ~w13689;
assign w13691 = w13414 & ~w13572;
assign v6356 = ~(w13574 | w13691);
assign w13692 = v6356;
assign w13693 = w13690 & ~w13692;
assign w13694 = ~w13690 & w13692;
assign v6357 = ~(w13693 | w13694);
assign w13695 = v6357;
assign v6358 = ~(w13602 | w13606);
assign w13696 = v6358;
assign v6359 = ~(w13605 | w13696);
assign w13697 = v6359;
assign v6360 = ~(w13695 | w13697);
assign w13698 = v6360;
assign w13699 = w13695 & w13697;
assign v6361 = ~(w13698 | w13699);
assign w13700 = v6361;
assign v6362 = ~(w13584 | w13587);
assign w13701 = v6362;
assign v6363 = ~(w13611 | w13624);
assign w13702 = v6363;
assign v6364 = ~(w13701 | w13702);
assign w13703 = v6364;
assign w13704 = w13701 & w13702;
assign v6365 = ~(w13703 | w13704);
assign w13705 = v6365;
assign w13706 = w13700 & w13705;
assign v6366 = ~(w13700 | w13705);
assign w13707 = v6366;
assign v6367 = ~(w13706 | w13707);
assign w13708 = v6367;
assign w13709 = ~w13688 & w13708;
assign w13710 = w13688 & ~w13708;
assign v6368 = ~(w13709 | w13710);
assign w13711 = v6368;
assign w13712 = w13687 & ~w13711;
assign w13713 = ~w13687 & w13711;
assign v6369 = ~(w13712 | w13713);
assign w13714 = v6369;
assign v6370 = ~(w13630 | w13633);
assign w13715 = v6370;
assign w13716 = ~w13714 & w13715;
assign w13717 = w13714 & ~w13715;
assign v6371 = ~(w13716 | w13717);
assign w13718 = v6371;
assign v6372 = ~(w13665 | w13668);
assign w13719 = v6372;
assign w13720 = w13614 & ~w13617;
assign v6373 = ~(w13619 | w13720);
assign w13721 = v6373;
assign w13722 = w13593 & ~w13595;
assign v6374 = ~(w13597 | w13722);
assign w13723 = v6374;
assign v6375 = ~(w13721 | w13723);
assign w13724 = v6375;
assign w13725 = w13721 & w13723;
assign v6376 = ~(w13724 | w13725);
assign w13726 = v6376;
assign w13727 = w13645 & ~w13647;
assign v6377 = ~(w13649 | w13727);
assign w13728 = v6377;
assign w13729 = ~w13726 & w13728;
assign w13730 = w13726 & ~w13728;
assign v6378 = ~(w13729 | w13730);
assign w13731 = v6378;
assign v6379 = ~(w13534 | w13538);
assign w13732 = v6379;
assign w13733 = ~w13731 & w13732;
assign w13734 = w13731 & ~w13732;
assign v6380 = ~(w13733 | w13734);
assign w13735 = v6380;
assign w13736 = pi35 & pi55;
assign w13737 = pi33 & pi57;
assign w13738 = pi34 & pi56;
assign v6381 = ~(w13737 | w13738);
assign w13739 = v6381;
assign w13740 = pi34 & pi57;
assign w13741 = w13603 & w13740;
assign v6382 = ~(w13739 | w13741);
assign w13742 = v6382;
assign w13743 = w13736 & ~w13742;
assign w13744 = ~w13736 & w13742;
assign v6383 = ~(w13743 | w13744);
assign w13745 = v6383;
assign w13746 = pi36 & pi54;
assign w13747 = pi37 & pi53;
assign v6384 = ~(w13596 | w13747);
assign w13748 = v6384;
assign w13749 = pi38 & pi53;
assign w13750 = w13464 & w13749;
assign v6385 = ~(w13748 | w13750);
assign w13751 = v6385;
assign w13752 = w13746 & ~w13751;
assign w13753 = ~w13746 & w13751;
assign v6386 = ~(w13752 | w13753);
assign w13754 = v6386;
assign v6387 = ~(w13745 | w13754);
assign w13755 = v6387;
assign w13756 = w13745 & w13754;
assign v6388 = ~(w13755 | w13756);
assign w13757 = v6388;
assign w13758 = pi42 & pi48;
assign w13759 = pi44 & pi46;
assign v6389 = ~(w13573 | w13759);
assign w13760 = v6389;
assign w13761 = pi44 & pi47;
assign w13762 = w13571 & w13761;
assign v6390 = ~(w13760 | w13762);
assign w13763 = v6390;
assign w13764 = w13758 & ~w13763;
assign w13765 = ~w13758 & w13763;
assign v6391 = ~(w13764 | w13765);
assign w13766 = v6391;
assign w13767 = w13757 & ~w13766;
assign w13768 = ~w13757 & w13766;
assign v6392 = ~(w13767 | w13768);
assign w13769 = v6392;
assign w13770 = w13735 & w13769;
assign v6393 = ~(w13735 | w13769);
assign w13771 = v6393;
assign v6394 = ~(w13770 | w13771);
assign w13772 = v6394;
assign w13773 = ~w13719 & w13772;
assign w13774 = w13719 & ~w13772;
assign v6395 = ~(w13773 | w13774);
assign w13775 = v6395;
assign v6396 = ~(w13659 | w13663);
assign w13776 = v6396;
assign v6397 = ~(w13642 | w13655);
assign w13777 = v6397;
assign w13778 = (~w13553 & ~w13555) | (~w13553 & w17226) | (~w13555 & w17226);
assign w13779 = pi39 & pi51;
assign w13780 = pi41 & pi49;
assign v6398 = ~(w13648 | w13780);
assign w13781 = v6398;
assign w13782 = pi41 & pi50;
assign w13783 = w13646 & w13782;
assign v6399 = ~(w13781 | w13783);
assign w13784 = v6399;
assign w13785 = w13779 & ~w13784;
assign w13786 = ~w13779 & w13784;
assign v6400 = ~(w13785 | w13786);
assign w13787 = v6400;
assign v6401 = ~(w13778 | w13787);
assign w13788 = v6401;
assign w13789 = w13778 & w13787;
assign v6402 = ~(w13788 | w13789);
assign w13790 = v6402;
assign w13791 = w13777 & ~w13790;
assign w13792 = ~w13777 & w13790;
assign v6403 = ~(w13791 | w13792);
assign w13793 = v6403;
assign v6404 = ~(w13564 | w13568);
assign w13794 = v6404;
assign w13795 = pi30 & pi60;
assign w13796 = pi31 & pi59;
assign v6405 = ~(w13618 | w13796);
assign w13797 = v6405;
assign w13798 = pi32 & pi59;
assign w13799 = w13616 & w13798;
assign v6406 = ~(w13797 | w13799);
assign w13800 = v6406;
assign w13801 = w13795 & ~w13800;
assign w13802 = ~w13795 & w13800;
assign v6407 = ~(w13801 | w13802);
assign w13803 = v6407;
assign v6408 = ~(w13794 | w13803);
assign w13804 = v6408;
assign w13805 = w13794 & w13803;
assign v6409 = ~(w13804 | w13805);
assign w13806 = v6409;
assign w13807 = pi27 & pi63;
assign w13808 = pi28 & pi62;
assign v6410 = ~(w13563 | w13808);
assign w13809 = v6410;
assign w13810 = pi29 & pi62;
assign w13811 = w13442 & w13810;
assign v6411 = ~(w13809 | w13811);
assign w13812 = v6411;
assign w13813 = w13807 & ~w13812;
assign w13814 = ~w13807 & w13812;
assign v6412 = ~(w13813 | w13814);
assign w13815 = v6412;
assign w13816 = w13806 & ~w13815;
assign w13817 = ~w13806 & w13815;
assign v6413 = ~(w13816 | w13817);
assign w13818 = v6413;
assign w13819 = w13793 & w13818;
assign v6414 = ~(w13793 | w13818);
assign w13820 = v6414;
assign v6415 = ~(w13819 | w13820);
assign w13821 = v6415;
assign w13822 = ~w13776 & w13821;
assign w13823 = w13776 & ~w13821;
assign v6416 = ~(w13822 | w13823);
assign w13824 = v6416;
assign w13825 = w13775 & w13824;
assign v6417 = ~(w13775 | w13824);
assign w13826 = v6417;
assign v6418 = ~(w13825 | w13826);
assign w13827 = v6418;
assign v6419 = ~(w13718 | w13827);
assign w13828 = v6419;
assign w13829 = w13718 & w13827;
assign v6420 = ~(w13828 | w13829);
assign w13830 = v6420;
assign w13831 = ~w13686 & w13830;
assign w13832 = w13686 & ~w13830;
assign v6421 = ~(w13831 | w13832);
assign w13833 = v6421;
assign w13834 = (~w10008 & w17861) | (~w10008 & w17862) | (w17861 & w17862);
assign w13835 = (w10008 & w17863) | (w10008 & w17864) | (w17863 & w17864);
assign v6422 = ~(w13834 | w13835);
assign w13836 = v6422;
assign v6423 = ~(w13717 | w13829);
assign w13837 = v6423;
assign w13838 = w13746 & ~w13748;
assign v6424 = ~(w13750 | w13838);
assign w13839 = v6424;
assign w13840 = w13807 & ~w13809;
assign v6425 = ~(w13811 | w13840);
assign w13841 = v6425;
assign v6426 = ~(w13839 | w13841);
assign w13842 = v6426;
assign w13843 = w13839 & w13841;
assign v6427 = ~(w13842 | w13843);
assign w13844 = v6427;
assign w13845 = w13795 & ~w13797;
assign v6428 = ~(w13799 | w13845);
assign w13846 = v6428;
assign w13847 = ~w13844 & w13846;
assign w13848 = w13844 & ~w13846;
assign v6429 = ~(w13847 | w13848);
assign w13849 = v6429;
assign v6430 = ~(w13788 | w13792);
assign w13850 = v6430;
assign w13851 = ~w13849 & w13850;
assign w13852 = w13849 & ~w13850;
assign v6431 = ~(w13851 | w13852);
assign w13853 = v6431;
assign w13854 = pi28 & pi63;
assign w13855 = pi40 & pi51;
assign v6432 = ~(w13782 | w13855);
assign w13856 = v6432;
assign w13857 = pi41 & pi51;
assign w13858 = w13648 & w13857;
assign v6433 = ~(w13856 | w13858);
assign w13859 = v6433;
assign w13860 = w13854 & ~w13859;
assign w13861 = ~w13854 & w13859;
assign v6434 = ~(w13860 | w13861);
assign w13862 = v6434;
assign w13863 = pi35 & pi56;
assign w13864 = pi43 & pi48;
assign v6435 = ~(w13761 | w13864);
assign w13865 = v6435;
assign w13866 = pi44 & pi48;
assign w13867 = w13573 & w13866;
assign v6436 = ~(w13865 | w13867);
assign w13868 = v6436;
assign w13869 = w13863 & ~w13868;
assign w13870 = ~w13863 & w13868;
assign v6437 = ~(w13869 | w13870);
assign w13871 = v6437;
assign v6438 = ~(w13862 | w13871);
assign w13872 = v6438;
assign w13873 = w13862 & w13871;
assign v6439 = ~(w13872 | w13873);
assign w13874 = v6439;
assign w13875 = ~pi45 & pi46;
assign w13876 = w13810 & ~w13875;
assign w13877 = ~w13810 & w13875;
assign v6440 = ~(w13876 | w13877);
assign w13878 = v6440;
assign w13879 = w13874 & ~w13878;
assign w13880 = ~w13874 & w13878;
assign v6441 = ~(w13879 | w13880);
assign w13881 = v6441;
assign v6442 = ~(w13853 | w13881);
assign w13882 = v6442;
assign w13883 = w13853 & w13881;
assign v6443 = ~(w13882 | w13883);
assign w13884 = v6443;
assign v6444 = ~(w13709 | w13713);
assign w13885 = v6444;
assign w13886 = ~w13884 & w13885;
assign w13887 = w13884 & ~w13885;
assign v6445 = ~(w13886 | w13887);
assign w13888 = v6445;
assign v6446 = ~(w13724 | w13730);
assign w13889 = v6446;
assign v6447 = ~(w13693 | w13699);
assign w13890 = v6447;
assign w13891 = pi42 & pi49;
assign w13892 = pi36 & pi55;
assign v6448 = ~(w13740 | w13892);
assign w13893 = v6448;
assign w13894 = w13740 & w13892;
assign v6449 = ~(w13893 | w13894);
assign w13895 = v6449;
assign w13896 = w13891 & ~w13895;
assign w13897 = ~w13891 & w13895;
assign v6450 = ~(w13896 | w13897);
assign w13898 = v6450;
assign v6451 = ~(w13890 | w13898);
assign w13899 = v6451;
assign w13900 = w13890 & w13898;
assign v6452 = ~(w13899 | w13900);
assign w13901 = v6452;
assign w13902 = w13889 & ~w13901;
assign w13903 = ~w13889 & w13901;
assign v6453 = ~(w13902 | w13903);
assign w13904 = v6453;
assign v6454 = ~(w13703 | w13706);
assign w13905 = v6454;
assign w13906 = pi37 & pi54;
assign w13907 = pi39 & pi52;
assign v6455 = ~(w13749 | w13907);
assign w13908 = v6455;
assign w13909 = pi39 & pi53;
assign w13910 = w13596 & w13909;
assign v6456 = ~(w13908 | w13910);
assign w13911 = v6456;
assign w13912 = w13906 & ~w13911;
assign w13913 = ~w13906 & w13911;
assign v6457 = ~(w13912 | w13913);
assign w13914 = v6457;
assign w13915 = w13779 & ~w13781;
assign v6458 = ~(w13783 | w13915);
assign w13916 = v6458;
assign v6459 = ~(w13914 | w13916);
assign w13917 = v6459;
assign w13918 = w13914 & w13916;
assign v6460 = ~(w13917 | w13918);
assign w13919 = v6460;
assign w13920 = pi31 & pi60;
assign w13921 = pi33 & pi58;
assign v6461 = ~(w13798 | w13921);
assign w13922 = v6461;
assign w13923 = pi33 & pi59;
assign w13924 = w13618 & w13923;
assign v6462 = ~(w13922 | w13924);
assign w13925 = v6462;
assign w13926 = w13920 & ~w13925;
assign w13927 = ~w13920 & w13925;
assign v6463 = ~(w13926 | w13927);
assign w13928 = v6463;
assign w13929 = w13919 & ~w13928;
assign w13930 = ~w13919 & w13928;
assign v6464 = ~(w13929 | w13930);
assign w13931 = v6464;
assign w13932 = ~w13905 & w13931;
assign w13933 = w13905 & ~w13931;
assign v6465 = ~(w13932 | w13933);
assign w13934 = v6465;
assign w13935 = w13904 & w13934;
assign v6466 = ~(w13904 | w13934);
assign w13936 = v6466;
assign v6467 = ~(w13935 | w13936);
assign w13937 = v6467;
assign w13938 = w13888 & w13937;
assign v6468 = ~(w13888 | w13937);
assign w13939 = v6468;
assign v6469 = ~(w13938 | w13939);
assign w13940 = v6469;
assign v6470 = ~(w13773 | w13825);
assign w13941 = v6470;
assign v6471 = ~(w13819 | w13822);
assign w13942 = v6471;
assign v6472 = ~(w13734 | w13770);
assign w13943 = v6472;
assign w13944 = pi30 & pi61;
assign w13945 = w13758 & ~w13760;
assign v6473 = ~(w13762 | w13945);
assign w13946 = v6473;
assign w13947 = w13944 & ~w13946;
assign w13948 = ~w13944 & w13946;
assign v6474 = ~(w13947 | w13948);
assign w13949 = v6474;
assign w13950 = w13736 & ~w13739;
assign v6475 = ~(w13741 | w13950);
assign w13951 = v6475;
assign w13952 = ~w13949 & w13951;
assign w13953 = w13949 & ~w13951;
assign v6476 = ~(w13952 | w13953);
assign w13954 = v6476;
assign v6477 = ~(w13804 | w13816);
assign w13955 = v6477;
assign v6478 = ~(w13755 | w13767);
assign w13956 = v6478;
assign v6479 = ~(w13955 | w13956);
assign w13957 = v6479;
assign w13958 = w13955 & w13956;
assign v6480 = ~(w13957 | w13958);
assign w13959 = v6480;
assign w13960 = w13954 & w13959;
assign v6481 = ~(w13954 | w13959);
assign w13961 = v6481;
assign v6482 = ~(w13960 | w13961);
assign w13962 = v6482;
assign w13963 = ~w13943 & w13962;
assign w13964 = w13943 & ~w13962;
assign v6483 = ~(w13963 | w13964);
assign w13965 = v6483;
assign w13966 = ~w13942 & w13965;
assign w13967 = w13942 & ~w13965;
assign v6484 = ~(w13966 | w13967);
assign w13968 = v6484;
assign w13969 = ~w13941 & w13968;
assign w13970 = w13941 & ~w13968;
assign v6485 = ~(w13969 | w13970);
assign w13971 = v6485;
assign w13972 = w13940 & w13971;
assign v6486 = ~(w13940 | w13971);
assign w13973 = v6486;
assign v6487 = ~(w13972 | w13973);
assign w13974 = v6487;
assign w13975 = ~w13837 & w13974;
assign w13976 = w13837 & ~w13974;
assign v6488 = ~(w13975 | w13976);
assign w13977 = v6488;
assign w13978 = (~w8795 & w17646) | (~w8795 & w17647) | (w17646 & w17647);
assign w13979 = (w11122 & w17648) | (w11122 & w17649) | (w17648 & w17649);
assign w13980 = (~w11122 & w17650) | (~w11122 & w17651) | (w17650 & w17651);
assign v6489 = ~(w13979 | w13980);
assign w13981 = v6489;
assign v6490 = ~(w13832 | w13976);
assign w13982 = v6490;
assign v6491 = ~(w13963 | w13966);
assign w13983 = v6491;
assign v6492 = ~(w13932 | w13935);
assign w13984 = v6492;
assign v6493 = ~(w13957 | w13960);
assign w13985 = v6493;
assign v6494 = ~(w13947 | w13953);
assign w13986 = v6494;
assign w13987 = pi31 & pi61;
assign w13988 = pi30 & pi62;
assign v6495 = ~(w13987 | w13988);
assign w13989 = v6495;
assign w13990 = pi31 & pi62;
assign w13991 = w13944 & w13990;
assign v6496 = ~(w13989 | w13991);
assign w13992 = v6496;
assign v6497 = ~(pi45 | w13810);
assign w13993 = v6497;
assign w13994 = pi46 & ~w13993;
assign w13995 = w13992 & w13994;
assign v6498 = ~(w13992 | w13994);
assign w13996 = v6498;
assign v6499 = ~(w13995 | w13996);
assign w13997 = v6499;
assign w13998 = pi40 & pi52;
assign v6500 = ~(w13857 | w13998);
assign w13999 = v6500;
assign w14000 = pi41 & pi52;
assign w14001 = w13855 & w14000;
assign v6501 = ~(w13999 | w14001);
assign w14002 = v6501;
assign w14003 = w13909 & ~w14002;
assign w14004 = ~w13909 & w14002;
assign v6502 = ~(w14003 | w14004);
assign w14005 = v6502;
assign w14006 = w13997 & ~w14005;
assign w14007 = ~w13997 & w14005;
assign v6503 = ~(w14006 | w14007);
assign w14008 = v6503;
assign w14009 = w13986 & ~w14008;
assign w14010 = ~w13986 & w14008;
assign v6504 = ~(w14009 | w14010);
assign w14011 = v6504;
assign w14012 = pi43 & pi49;
assign w14013 = pi45 & pi47;
assign v6505 = ~(w13866 | w14013);
assign w14014 = v6505;
assign w14015 = pi45 & pi48;
assign w14016 = w13761 & w14015;
assign v6506 = ~(w14014 | w14016);
assign w14017 = v6506;
assign w14018 = w14012 & ~w14017;
assign w14019 = ~w14012 & w14017;
assign v6507 = ~(w14018 | w14019);
assign w14020 = v6507;
assign w14021 = pi34 & pi58;
assign w14022 = pi35 & pi57;
assign w14023 = pi42 & pi50;
assign v6508 = ~(w14022 | w14023);
assign w14024 = v6508;
assign w14025 = w14022 & w14023;
assign v6509 = ~(w14024 | w14025);
assign w14026 = v6509;
assign w14027 = w14021 & ~w14026;
assign w14028 = ~w14021 & w14026;
assign v6510 = ~(w14027 | w14028);
assign w14029 = v6510;
assign v6511 = ~(w14020 | w14029);
assign w14030 = v6511;
assign w14031 = w14020 & w14029;
assign v6512 = ~(w14030 | w14031);
assign w14032 = v6512;
assign w14033 = pi36 & pi56;
assign w14034 = pi29 & pi63;
assign v6513 = ~(w13923 | w14034);
assign w14035 = v6513;
assign w14036 = w13923 & w14034;
assign v6514 = ~(w14035 | w14036);
assign w14037 = v6514;
assign w14038 = w14033 & ~w14037;
assign w14039 = ~w14033 & w14037;
assign v6515 = ~(w14038 | w14039);
assign w14040 = v6515;
assign w14041 = w14032 & ~w14040;
assign w14042 = ~w14032 & w14040;
assign v6516 = ~(w14041 | w14042);
assign w14043 = v6516;
assign v6517 = ~(w14011 | w14043);
assign w14044 = v6517;
assign w14045 = w14011 & w14043;
assign v6518 = ~(w14044 | w14045);
assign w14046 = v6518;
assign w14047 = ~w13985 & w14046;
assign w14048 = w13985 & ~w14046;
assign v6519 = ~(w14047 | w14048);
assign w14049 = v6519;
assign w14050 = ~w13984 & w14049;
assign w14051 = w13984 & ~w14049;
assign v6520 = ~(w14050 | w14051);
assign w14052 = v6520;
assign w14053 = ~w13983 & w14052;
assign w14054 = w13983 & ~w14052;
assign v6521 = ~(w14053 | w14054);
assign w14055 = v6521;
assign v6522 = ~(w13887 | w13938);
assign w14056 = v6522;
assign v6523 = ~(w13872 | w13879);
assign w14057 = v6523;
assign v6524 = ~(w13917 | w13929);
assign w14058 = v6524;
assign v6525 = ~(w13842 | w13848);
assign w14059 = v6525;
assign v6526 = ~(w14058 | w14059);
assign w14060 = v6526;
assign w14061 = w14058 & w14059;
assign v6527 = ~(w14060 | w14061);
assign w14062 = v6527;
assign w14063 = w14057 & ~w14062;
assign w14064 = ~w14057 & w14062;
assign v6528 = ~(w14063 | w14064);
assign w14065 = v6528;
assign v6529 = ~(w13852 | w13883);
assign w14066 = v6529;
assign v6530 = ~(w13899 | w13903);
assign w14067 = v6530;
assign w14068 = w13920 & ~w13922;
assign v6531 = ~(w13924 | w14068);
assign w14069 = v6531;
assign w14070 = w13906 & ~w13908;
assign v6532 = ~(w13910 | w14070);
assign w14071 = v6532;
assign v6533 = ~(w14069 | w14071);
assign w14072 = v6533;
assign w14073 = w14069 & w14071;
assign v6534 = ~(w14072 | w14073);
assign w14074 = v6534;
assign w14075 = w13854 & ~w13856;
assign v6535 = ~(w13858 | w14075);
assign w14076 = v6535;
assign w14077 = ~w14074 & w14076;
assign w14078 = w14074 & ~w14076;
assign v6536 = ~(w14077 | w14078);
assign w14079 = v6536;
assign v6537 = ~(w13891 | w13894);
assign w14080 = v6537;
assign v6538 = ~(w13893 | w14080);
assign w14081 = v6538;
assign w14082 = w13863 & ~w13865;
assign v6539 = ~(w13867 | w14082);
assign w14083 = v6539;
assign w14084 = w14081 & ~w14083;
assign w14085 = ~w14081 & w14083;
assign v6540 = ~(w14084 | w14085);
assign w14086 = v6540;
assign w14087 = pi32 & pi60;
assign w14088 = pi37 & pi55;
assign w14089 = pi38 & pi54;
assign v6541 = ~(w14088 | w14089);
assign w14090 = v6541;
assign w14091 = pi38 & pi55;
assign w14092 = w13906 & w14091;
assign v6542 = ~(w14090 | w14092);
assign w14093 = v6542;
assign w14094 = w14087 & ~w14093;
assign w14095 = ~w14087 & w14093;
assign v6543 = ~(w14094 | w14095);
assign w14096 = v6543;
assign w14097 = ~w14086 & w14096;
assign w14098 = w14086 & ~w14096;
assign v6544 = ~(w14097 | w14098);
assign w14099 = v6544;
assign v6545 = ~(w14079 | w14099);
assign w14100 = v6545;
assign w14101 = w14079 & w14099;
assign v6546 = ~(w14100 | w14101);
assign w14102 = v6546;
assign w14103 = ~w14067 & w14102;
assign w14104 = w14067 & ~w14102;
assign v6547 = ~(w14103 | w14104);
assign w14105 = v6547;
assign w14106 = ~w14066 & w14105;
assign w14107 = w14066 & ~w14105;
assign v6548 = ~(w14106 | w14107);
assign w14108 = v6548;
assign w14109 = w14065 & w14108;
assign v6549 = ~(w14065 | w14108);
assign w14110 = v6549;
assign v6550 = ~(w14109 | w14110);
assign w14111 = v6550;
assign w14112 = ~w14056 & w14111;
assign w14113 = w14056 & ~w14111;
assign v6551 = ~(w14112 | w14113);
assign w14114 = v6551;
assign w14115 = w14055 & w14114;
assign v6552 = ~(w14055 | w14114);
assign w14116 = v6552;
assign v6553 = ~(w14115 | w14116);
assign w14117 = v6553;
assign v6554 = ~(w13969 | w13972);
assign w14118 = v6554;
assign w14119 = w14117 & ~w14118;
assign w14120 = ~w14117 & w14118;
assign v6555 = ~(w14119 | w14120);
assign w14121 = v6555;
assign w14122 = (w12329 & w17493) | (w12329 & w17494) | (w17493 & w17494);
assign w14123 = (~w12329 & w17495) | (~w12329 & w17496) | (w17495 & w17496);
assign v6556 = ~(w14122 | w14123);
assign w14124 = v6556;
assign v6557 = ~(w13975 | w14119);
assign w14125 = v6557;
assign v6558 = ~(w14112 | w14115);
assign w14126 = v6558;
assign v6559 = ~(w14050 | w14053);
assign w14127 = v6559;
assign v6560 = ~(w14030 | w14041);
assign w14128 = v6560;
assign v6561 = ~(w14084 | w14098);
assign w14129 = v6561;
assign v6562 = ~(w14072 | w14078);
assign w14130 = v6562;
assign v6563 = ~(w14129 | w14130);
assign w14131 = v6563;
assign w14132 = w14129 & w14130;
assign v6564 = ~(w14131 | w14132);
assign w14133 = v6564;
assign w14134 = w14128 & ~w14133;
assign w14135 = ~w14128 & w14133;
assign v6565 = ~(w14134 | w14135);
assign w14136 = v6565;
assign v6566 = ~(w14101 | w14103);
assign w14137 = v6566;
assign w14138 = ~w14136 & w14137;
assign w14139 = w14136 & ~w14137;
assign v6567 = ~(w14138 | w14139);
assign w14140 = v6567;
assign v6568 = ~(w14006 | w14010);
assign w14141 = v6568;
assign v6569 = ~(w14021 | w14025);
assign w14142 = v6569;
assign v6570 = ~(w14024 | w14142);
assign w14143 = v6570;
assign w14144 = w14012 & ~w14014;
assign v6571 = ~(w14016 | w14144);
assign w14145 = v6571;
assign w14146 = w14143 & ~w14145;
assign w14147 = ~w14143 & w14145;
assign v6572 = ~(w14146 | w14147);
assign w14148 = v6572;
assign w14149 = w13909 & ~w13999;
assign v6573 = ~(w14001 | w14149);
assign w14150 = v6573;
assign w14151 = ~w14148 & w14150;
assign w14152 = w14148 & ~w14150;
assign v6574 = ~(w14151 | w14152);
assign w14153 = v6574;
assign v6575 = ~(w13991 | w13995);
assign w14154 = v6575;
assign v6576 = ~(w14033 | w14036);
assign w14155 = v6576;
assign v6577 = ~(w14035 | w14155);
assign w14156 = v6577;
assign w14157 = w14087 & ~w14090;
assign v6578 = ~(w14092 | w14157);
assign w14158 = v6578;
assign w14159 = w14156 & ~w14158;
assign w14160 = ~w14156 & w14158;
assign v6579 = ~(w14159 | w14160);
assign w14161 = v6579;
assign w14162 = w14154 & ~w14161;
assign w14163 = ~w14154 & w14161;
assign v6580 = ~(w14162 | w14163);
assign w14164 = v6580;
assign w14165 = w14153 & w14164;
assign v6581 = ~(w14153 | w14164);
assign w14166 = v6581;
assign v6582 = ~(w14165 | w14166);
assign w14167 = v6582;
assign w14168 = ~w14141 & w14167;
assign w14169 = w14141 & ~w14167;
assign v6583 = ~(w14168 | w14169);
assign w14170 = v6583;
assign w14171 = w14140 & w14170;
assign v6584 = ~(w14140 | w14170);
assign w14172 = v6584;
assign v6585 = ~(w14171 | w14172);
assign w14173 = v6585;
assign w14174 = ~w14127 & w14173;
assign w14175 = w14127 & ~w14173;
assign v6586 = ~(w14174 | w14175);
assign w14176 = v6586;
assign v6587 = ~(w14106 | w14109);
assign w14177 = v6587;
assign v6588 = ~(w14045 | w14047);
assign w14178 = v6588;
assign v6589 = ~(w14060 | w14064);
assign w14179 = v6589;
assign w14180 = pi30 & pi63;
assign w14181 = pi32 & pi61;
assign w14182 = pi33 & pi60;
assign v6590 = ~(w14181 | w14182);
assign w14183 = v6590;
assign w14184 = pi33 & pi61;
assign w14185 = w14087 & w14184;
assign v6591 = ~(w14183 | w14185);
assign w14186 = v6591;
assign w14187 = w14180 & ~w14186;
assign w14188 = ~w14180 & w14186;
assign v6592 = ~(w14187 | w14188);
assign w14189 = v6592;
assign w14190 = pi35 & pi58;
assign w14191 = pi36 & pi57;
assign w14192 = pi39 & pi54;
assign v6593 = ~(w14191 | w14192);
assign w14193 = v6593;
assign w14194 = w14191 & w14192;
assign v6594 = ~(w14193 | w14194);
assign w14195 = v6594;
assign w14196 = w14190 & ~w14195;
assign w14197 = ~w14190 & w14195;
assign v6595 = ~(w14196 | w14197);
assign w14198 = v6595;
assign v6596 = ~(w14189 | w14198);
assign w14199 = v6596;
assign w14200 = w14189 & w14198;
assign v6597 = ~(w14199 | w14200);
assign w14201 = v6597;
assign w14202 = pi34 & pi59;
assign w14203 = pi40 & pi53;
assign v6598 = ~(w14000 | w14203);
assign w14204 = v6598;
assign w14205 = pi41 & pi53;
assign w14206 = w13998 & w14205;
assign v6599 = ~(w14204 | w14206);
assign w14207 = v6599;
assign w14208 = w14202 & ~w14207;
assign w14209 = ~w14202 & w14207;
assign v6600 = ~(w14208 | w14209);
assign w14210 = v6600;
assign w14211 = w14201 & ~w14210;
assign w14212 = ~w14201 & w14210;
assign v6601 = ~(w14211 | w14212);
assign w14213 = v6601;
assign w14214 = pi42 & pi51;
assign w14215 = pi44 & pi49;
assign w14216 = pi43 & pi50;
assign v6602 = ~(w14215 | w14216);
assign w14217 = v6602;
assign w14218 = pi44 & pi50;
assign w14219 = w14012 & w14218;
assign v6603 = ~(w14217 | w14219);
assign w14220 = v6603;
assign w14221 = w14214 & ~w14220;
assign w14222 = ~w14214 & w14220;
assign v6604 = ~(w14221 | w14222);
assign w14223 = v6604;
assign w14224 = pi37 & pi56;
assign v6605 = ~(w14015 | w14091);
assign w14225 = v6605;
assign w14226 = w14015 & w14091;
assign v6606 = ~(w14225 | w14226);
assign w14227 = v6606;
assign w14228 = w14224 & ~w14227;
assign w14229 = ~w14224 & w14227;
assign v6607 = ~(w14228 | w14229);
assign w14230 = v6607;
assign v6608 = ~(w14223 | w14230);
assign w14231 = v6608;
assign w14232 = w14223 & w14230;
assign v6609 = ~(w14231 | w14232);
assign w14233 = v6609;
assign w14234 = ~pi46 & pi47;
assign w14235 = w13990 & ~w14234;
assign w14236 = ~w13990 & w14234;
assign v6610 = ~(w14235 | w14236);
assign w14237 = v6610;
assign w14238 = w14233 & ~w14237;
assign w14239 = ~w14233 & w14237;
assign v6611 = ~(w14238 | w14239);
assign w14240 = v6611;
assign w14241 = w14213 & w14240;
assign v6612 = ~(w14213 | w14240);
assign w14242 = v6612;
assign v6613 = ~(w14241 | w14242);
assign w14243 = v6613;
assign w14244 = ~w14179 & w14243;
assign w14245 = w14179 & ~w14243;
assign v6614 = ~(w14244 | w14245);
assign w14246 = v6614;
assign w14247 = ~w14178 & w14246;
assign w14248 = w14178 & ~w14246;
assign v6615 = ~(w14247 | w14248);
assign w14249 = v6615;
assign w14250 = w14177 & ~w14249;
assign w14251 = ~w14177 & w14249;
assign v6616 = ~(w14250 | w14251);
assign w14252 = v6616;
assign w14253 = w14176 & w14252;
assign v6617 = ~(w14176 | w14252);
assign w14254 = v6617;
assign v6618 = ~(w14253 | w14254);
assign w14255 = v6618;
assign w14256 = ~w14126 & w14255;
assign w14257 = w14126 & ~w14255;
assign v6619 = ~(w14256 | w14257);
assign w14258 = v6619;
assign w14259 = (w11122 & w17652) | (w11122 & w17653) | (w17652 & w17653);
assign w14260 = (~w11122 & w17654) | (~w11122 & w17655) | (w17654 & w17655);
assign v6620 = ~(w14259 | w14260);
assign w14261 = v6620;
assign v6621 = ~(w14247 | w14251);
assign w14262 = v6621;
assign v6622 = ~(w14241 | w14244);
assign w14263 = v6622;
assign v6623 = ~(w14199 | w14211);
assign w14264 = v6623;
assign v6624 = ~(w14159 | w14163);
assign w14265 = v6624;
assign v6625 = ~(w14146 | w14152);
assign w14266 = v6625;
assign v6626 = ~(w14265 | w14266);
assign w14267 = v6626;
assign w14268 = w14265 & w14266;
assign v6627 = ~(w14267 | w14268);
assign w14269 = v6627;
assign w14270 = w14264 & ~w14269;
assign w14271 = ~w14264 & w14269;
assign v6628 = ~(w14270 | w14271);
assign w14272 = v6628;
assign v6629 = ~(w14165 | w14168);
assign w14273 = v6629;
assign w14274 = ~w14272 & w14273;
assign w14275 = w14272 & ~w14273;
assign v6630 = ~(w14274 | w14275);
assign w14276 = v6630;
assign w14277 = ~w14263 & w14276;
assign w14278 = w14263 & ~w14276;
assign v6631 = ~(w14277 | w14278);
assign w14279 = v6631;
assign w14280 = ~w14262 & w14279;
assign w14281 = w14262 & ~w14279;
assign v6632 = ~(w14280 | w14281);
assign w14282 = v6632;
assign v6633 = ~(w14139 | w14171);
assign w14283 = v6633;
assign v6634 = ~(w14231 | w14238);
assign w14284 = v6634;
assign w14285 = pi31 & pi63;
assign v6635 = ~(pi46 | w13990);
assign w14286 = v6635;
assign w14287 = pi47 & ~w14286;
assign w14288 = w14285 & w14287;
assign v6636 = ~(w14285 | w14287);
assign w14289 = v6636;
assign v6637 = ~(w14288 | w14289);
assign w14290 = v6637;
assign v6638 = ~(w14224 | w14226);
assign w14291 = v6638;
assign v6639 = ~(w14225 | w14291);
assign w14292 = v6639;
assign w14293 = w14290 & w14292;
assign v6640 = ~(w14290 | w14292);
assign w14294 = v6640;
assign v6641 = ~(w14293 | w14294);
assign w14295 = v6641;
assign w14296 = w14284 & ~w14295;
assign w14297 = ~w14284 & w14295;
assign v6642 = ~(w14296 | w14297);
assign w14298 = v6642;
assign v6643 = ~(w14190 | w14194);
assign w14299 = v6643;
assign v6644 = ~(w14193 | w14299);
assign w14300 = v6644;
assign w14301 = w14180 & ~w14183;
assign v6645 = ~(w14185 | w14301);
assign w14302 = v6645;
assign w14303 = w14300 & ~w14302;
assign w14304 = ~w14300 & w14302;
assign v6646 = ~(w14303 | w14304);
assign w14305 = v6646;
assign w14306 = w14202 & ~w14204;
assign v6647 = ~(w14206 | w14306);
assign w14307 = v6647;
assign w14308 = ~w14305 & w14307;
assign w14309 = w14305 & ~w14307;
assign v6648 = ~(w14308 | w14309);
assign w14310 = v6648;
assign w14311 = w14298 & w14310;
assign v6649 = ~(w14298 | w14310);
assign w14312 = v6649;
assign v6650 = ~(w14311 | w14312);
assign w14313 = v6650;
assign w14314 = ~w14283 & w14313;
assign w14315 = w14283 & ~w14313;
assign v6651 = ~(w14314 | w14315);
assign w14316 = v6651;
assign v6652 = ~(w14131 | w14135);
assign w14317 = v6652;
assign w14318 = pi36 & pi58;
assign w14319 = pi43 & pi51;
assign v6653 = ~(w14218 | w14319);
assign w14320 = v6653;
assign w14321 = pi44 & pi51;
assign w14322 = w14216 & w14321;
assign v6654 = ~(w14320 | w14322);
assign w14323 = v6654;
assign w14324 = w14318 & ~w14323;
assign w14325 = ~w14318 & w14323;
assign v6655 = ~(w14324 | w14325);
assign w14326 = v6655;
assign w14327 = pi40 & pi54;
assign w14328 = pi42 & pi52;
assign v6656 = ~(w14205 | w14328);
assign w14329 = v6656;
assign w14330 = pi42 & pi53;
assign w14331 = w14000 & w14330;
assign v6657 = ~(w14329 | w14331);
assign w14332 = v6657;
assign w14333 = w14327 & ~w14332;
assign w14334 = ~w14327 & w14332;
assign v6658 = ~(w14333 | w14334);
assign w14335 = v6658;
assign v6659 = ~(w14326 | w14335);
assign w14336 = v6659;
assign w14337 = w14326 & w14335;
assign v6660 = ~(w14336 | w14337);
assign w14338 = v6660;
assign w14339 = pi45 & pi49;
assign w14340 = pi38 & pi56;
assign w14341 = pi46 & pi48;
assign v6661 = ~(w14340 | w14341);
assign w14342 = v6661;
assign w14343 = w14340 & w14341;
assign v6662 = ~(w14342 | w14343);
assign w14344 = v6662;
assign w14345 = w14339 & ~w14344;
assign w14346 = ~w14339 & w14344;
assign v6663 = ~(w14345 | w14346);
assign w14347 = v6663;
assign w14348 = w14338 & ~w14347;
assign w14349 = ~w14338 & w14347;
assign v6664 = ~(w14348 | w14349);
assign w14350 = v6664;
assign w14351 = ~w14317 & w14350;
assign w14352 = w14317 & ~w14350;
assign v6665 = ~(w14351 | w14352);
assign w14353 = v6665;
assign w14354 = w14214 & ~w14217;
assign v6666 = ~(w14219 | w14354);
assign w14355 = v6666;
assign w14356 = pi35 & pi59;
assign v6667 = ~(w14184 | w14356);
assign w14357 = v6667;
assign w14358 = w14184 & w14356;
assign v6668 = ~(w14357 | w14358);
assign w14359 = v6668;
assign w14360 = w8301 & ~w14359;
assign w14361 = ~w8301 & w14359;
assign v6669 = ~(w14360 | w14361);
assign w14362 = v6669;
assign v6670 = ~(w14355 | w14362);
assign w14363 = v6670;
assign w14364 = w14355 & w14362;
assign v6671 = ~(w14363 | w14364);
assign w14365 = v6671;
assign w14366 = pi37 & pi57;
assign w14367 = pi34 & pi60;
assign w14368 = pi39 & pi55;
assign v6672 = ~(w14367 | w14368);
assign w14369 = v6672;
assign w14370 = w14367 & w14368;
assign v6673 = ~(w14369 | w14370);
assign w14371 = v6673;
assign w14372 = w14366 & ~w14371;
assign w14373 = ~w14366 & w14371;
assign v6674 = ~(w14372 | w14373);
assign w14374 = v6674;
assign w14375 = w14365 & ~w14374;
assign w14376 = ~w14365 & w14374;
assign v6675 = ~(w14375 | w14376);
assign w14377 = v6675;
assign w14378 = w14353 & w14377;
assign v6676 = ~(w14353 | w14377);
assign w14379 = v6676;
assign v6677 = ~(w14378 | w14379);
assign w14380 = v6677;
assign w14381 = w14316 & w14380;
assign v6678 = ~(w14316 | w14380);
assign w14382 = v6678;
assign v6679 = ~(w14381 | w14382);
assign w14383 = v6679;
assign v6680 = ~(w14282 | w14383);
assign w14384 = v6680;
assign w14385 = w14282 & w14383;
assign v6681 = ~(w14384 | w14385);
assign w14386 = v6681;
assign v6682 = ~(w14174 | w14253);
assign w14387 = v6682;
assign w14388 = ~w14386 & w14387;
assign w14389 = w14386 & ~w14387;
assign v6683 = ~(w14388 | w14389);
assign w14390 = v6683;
assign w14391 = (~w12329 & w17497) | (~w12329 & w17498) | (w17497 & w17498);
assign w14392 = (w12329 & w17499) | (w12329 & w17500) | (w17499 & w17500);
assign v6684 = ~(w14391 | w14392);
assign w14393 = v6684;
assign v6685 = ~(w14314 | w14381);
assign w14394 = v6685;
assign v6686 = ~(w14351 | w14378);
assign w14395 = v6686;
assign v6687 = ~(w14303 | w14309);
assign w14396 = v6687;
assign w14397 = pi36 & pi59;
assign w14398 = pi35 & pi60;
assign v6688 = ~(w14397 | w14398);
assign w14399 = v6688;
assign w14400 = pi36 & pi60;
assign w14401 = w14356 & w14400;
assign v6689 = ~(w14399 | w14401);
assign w14402 = v6689;
assign v6690 = ~(w14339 | w14343);
assign w14403 = v6690;
assign v6691 = ~(w14342 | w14403);
assign w14404 = v6691;
assign w14405 = w14402 & w14404;
assign v6692 = ~(w14402 | w14404);
assign w14406 = v6692;
assign v6693 = ~(w14405 | w14406);
assign w14407 = v6693;
assign v6694 = ~(w14288 | w14293);
assign w14408 = v6694;
assign w14409 = w14407 & ~w14408;
assign w14410 = ~w14407 & w14408;
assign v6695 = ~(w14409 | w14410);
assign w14411 = v6695;
assign w14412 = w14396 & ~w14411;
assign w14413 = ~w14396 & w14411;
assign v6696 = ~(w14412 | w14413);
assign w14414 = v6696;
assign v6697 = ~(w14297 | w14311);
assign w14415 = v6697;
assign w14416 = ~w14414 & w14415;
assign w14417 = w14414 & ~w14415;
assign v6698 = ~(w14416 | w14417);
assign w14418 = v6698;
assign w14419 = ~w14395 & w14418;
assign w14420 = w14395 & ~w14418;
assign v6699 = ~(w14419 | w14420);
assign w14421 = v6699;
assign w14422 = ~w14394 & w14421;
assign w14423 = w14394 & ~w14421;
assign v6700 = ~(w14422 | w14423);
assign w14424 = v6700;
assign v6701 = ~(w14267 | w14271);
assign w14425 = v6701;
assign w14426 = pi39 & pi56;
assign w14427 = pi46 & pi49;
assign w14428 = pi45 & pi50;
assign v6702 = ~(w14427 | w14428);
assign w14429 = v6702;
assign w14430 = pi46 & pi50;
assign w14431 = w14339 & w14430;
assign v6703 = ~(w14429 | w14431);
assign w14432 = v6703;
assign w14433 = w14426 & ~w14432;
assign w14434 = ~w14426 & w14432;
assign v6704 = ~(w14433 | w14434);
assign w14435 = v6704;
assign w14436 = pi33 & pi62;
assign w14437 = ~pi47 & pi48;
assign w14438 = w14436 & ~w14437;
assign w14439 = ~w14436 & w14437;
assign v6705 = ~(w14438 | w14439);
assign w14440 = v6705;
assign v6706 = ~(w14435 | w14440);
assign w14441 = v6706;
assign w14442 = w14435 & w14440;
assign v6707 = ~(w14441 | w14442);
assign w14443 = v6707;
assign w14444 = pi43 & pi52;
assign v6708 = ~(w14321 | w14444);
assign w14445 = v6708;
assign w14446 = pi44 & pi52;
assign w14447 = w14319 & w14446;
assign v6709 = ~(w14445 | w14447);
assign w14448 = v6709;
assign w14449 = w14330 & ~w14448;
assign w14450 = ~w14330 & w14448;
assign v6710 = ~(w14449 | w14450);
assign w14451 = v6710;
assign w14452 = w14443 & ~w14451;
assign w14453 = ~w14443 & w14451;
assign v6711 = ~(w14452 | w14453);
assign w14454 = v6711;
assign w14455 = ~w14425 & w14454;
assign w14456 = w14425 & ~w14454;
assign v6712 = ~(w14455 | w14456);
assign w14457 = v6712;
assign w14458 = w14318 & ~w14320;
assign v6713 = ~(w14322 | w14458);
assign w14459 = v6713;
assign w14460 = pi37 & pi58;
assign w14461 = pi40 & pi55;
assign w14462 = pi38 & pi57;
assign v6714 = ~(w14461 | w14462);
assign w14463 = v6714;
assign w14464 = w14461 & w14462;
assign v6715 = ~(w14463 | w14464);
assign w14465 = v6715;
assign w14466 = w14460 & ~w14465;
assign w14467 = ~w14460 & w14465;
assign v6716 = ~(w14466 | w14467);
assign w14468 = v6716;
assign v6717 = ~(w14459 | w14468);
assign w14469 = v6717;
assign w14470 = w14459 & w14468;
assign v6718 = ~(w14469 | w14470);
assign w14471 = v6718;
assign w14472 = pi41 & pi54;
assign w14473 = pi34 & pi61;
assign v6719 = ~(w8302 | w14473);
assign w14474 = v6719;
assign w14475 = w8302 & w14473;
assign v6720 = ~(w14474 | w14475);
assign w14476 = v6720;
assign w14477 = w14472 & ~w14476;
assign w14478 = ~w14472 & w14476;
assign v6721 = ~(w14477 | w14478);
assign w14479 = v6721;
assign w14480 = w14471 & ~w14479;
assign w14481 = ~w14471 & w14479;
assign v6722 = ~(w14480 | w14481);
assign w14482 = v6722;
assign v6723 = ~(w14457 | w14482);
assign w14483 = v6723;
assign w14484 = w14457 & w14482;
assign v6724 = ~(w14483 | w14484);
assign w14485 = v6724;
assign v6725 = ~(w14275 | w14277);
assign w14486 = v6725;
assign v6726 = ~(w8301 | w14358);
assign w14487 = v6726;
assign v6727 = ~(w14357 | w14487);
assign w14488 = v6727;
assign v6728 = ~(w14366 | w14370);
assign w14489 = v6728;
assign v6729 = ~(w14369 | w14489);
assign w14490 = v6729;
assign w14491 = w14488 & w14490;
assign v6730 = ~(w14488 | w14490);
assign w14492 = v6730;
assign v6731 = ~(w14491 | w14492);
assign w14493 = v6731;
assign w14494 = w14327 & ~w14329;
assign v6732 = ~(w14331 | w14494);
assign w14495 = v6732;
assign w14496 = ~w14493 & w14495;
assign w14497 = w14493 & ~w14495;
assign v6733 = ~(w14496 | w14497);
assign w14498 = v6733;
assign v6734 = ~(w14336 | w14348);
assign w14499 = v6734;
assign v6735 = ~(w14363 | w14375);
assign w14500 = v6735;
assign v6736 = ~(w14499 | w14500);
assign w14501 = v6736;
assign w14502 = w14499 & w14500;
assign v6737 = ~(w14501 | w14502);
assign w14503 = v6737;
assign w14504 = w14498 & w14503;
assign v6738 = ~(w14498 | w14503);
assign w14505 = v6738;
assign v6739 = ~(w14504 | w14505);
assign w14506 = v6739;
assign w14507 = ~w14486 & w14506;
assign w14508 = w14486 & ~w14506;
assign v6740 = ~(w14507 | w14508);
assign w14509 = v6740;
assign w14510 = w14485 & w14509;
assign v6741 = ~(w14485 | w14509);
assign w14511 = v6741;
assign v6742 = ~(w14510 | w14511);
assign w14512 = v6742;
assign v6743 = ~(w14424 | w14512);
assign w14513 = v6743;
assign w14514 = w14424 & w14512;
assign v6744 = ~(w14513 | w14514);
assign w14515 = v6744;
assign v6745 = ~(w14280 | w14385);
assign w14516 = v6745;
assign w14517 = w14515 & ~w14516;
assign w14518 = ~w14515 & w14516;
assign v6746 = ~(w14517 | w14518);
assign w14519 = v6746;
assign v6747 = ~(w14257 | w14388);
assign w14520 = v6747;
assign w14521 = (w12329 & w17501) | (w12329 & w17502) | (w17501 & w17502);
assign w14522 = (~w12329 & w17503) | (~w12329 & w17504) | (w17503 & w17504);
assign v6748 = ~(w14521 | w14522);
assign w14523 = v6748;
assign v6749 = ~(w14389 | w14517);
assign w14524 = v6749;
assign v6750 = ~(w14422 | w14514);
assign w14525 = v6750;
assign v6751 = ~(w14417 | w14419);
assign w14526 = v6751;
assign v6752 = ~(pi47 | w14436);
assign w14527 = v6752;
assign w14528 = pi48 & ~w14527;
assign w14529 = w14426 & ~w14429;
assign v6753 = ~(w14431 | w14529);
assign w14530 = v6753;
assign w14531 = w14528 & ~w14530;
assign w14532 = ~w14528 & w14530;
assign v6754 = ~(w14531 | w14532);
assign w14533 = v6754;
assign w14534 = w14330 & ~w14445;
assign v6755 = ~(w14447 | w14534);
assign w14535 = v6755;
assign w14536 = ~w14533 & w14535;
assign w14537 = w14533 & ~w14535;
assign v6756 = ~(w14536 | w14537);
assign w14538 = v6756;
assign v6757 = ~(w14469 | w14480);
assign w14539 = v6757;
assign v6758 = ~(w14441 | w14452);
assign w14540 = v6758;
assign v6759 = ~(w14539 | w14540);
assign w14541 = v6759;
assign w14542 = w14539 & w14540;
assign v6760 = ~(w14541 | w14542);
assign w14543 = v6760;
assign w14544 = w14538 & w14543;
assign v6761 = ~(w14538 | w14543);
assign w14545 = v6761;
assign v6762 = ~(w14544 | w14545);
assign w14546 = v6762;
assign w14547 = ~w14526 & w14546;
assign w14548 = w14526 & ~w14546;
assign v6763 = ~(w14547 | w14548);
assign w14549 = v6763;
assign v6764 = ~(w14491 | w14497);
assign w14550 = v6764;
assign w14551 = pi33 & pi63;
assign w14552 = pi35 & pi61;
assign w14553 = pi34 & pi62;
assign v6765 = ~(w14552 | w14553);
assign w14554 = v6765;
assign w14555 = pi35 & pi62;
assign w14556 = w14473 & w14555;
assign v6766 = ~(w14554 | w14556);
assign w14557 = v6766;
assign w14558 = w14551 & ~w14557;
assign w14559 = ~w14551 & w14557;
assign v6767 = ~(w14558 | w14559);
assign w14560 = v6767;
assign w14561 = pi41 & pi55;
assign w14562 = pi42 & pi54;
assign w14563 = pi43 & pi53;
assign v6768 = ~(w14562 | w14563);
assign w14564 = v6768;
assign w14565 = pi43 & pi54;
assign w14566 = w14330 & w14565;
assign v6769 = ~(w14564 | w14566);
assign w14567 = v6769;
assign w14568 = w14561 & ~w14567;
assign w14569 = ~w14561 & w14567;
assign v6770 = ~(w14568 | w14569);
assign w14570 = v6770;
assign v6771 = ~(w14560 | w14570);
assign w14571 = v6771;
assign w14572 = w14560 & w14570;
assign v6772 = ~(w14571 | w14572);
assign w14573 = v6772;
assign w14574 = w14550 & ~w14573;
assign w14575 = ~w14550 & w14573;
assign v6773 = ~(w14574 | w14575);
assign w14576 = v6773;
assign v6774 = ~(w14401 | w14405);
assign w14577 = v6774;
assign v6775 = ~(w14472 | w14475);
assign w14578 = v6775;
assign v6776 = ~(w14474 | w14578);
assign w14579 = v6776;
assign v6777 = ~(w14460 | w14464);
assign w14580 = v6777;
assign v6778 = ~(w14463 | w14580);
assign w14581 = v6778;
assign w14582 = w14579 & w14581;
assign v6779 = ~(w14579 | w14581);
assign w14583 = v6779;
assign v6780 = ~(w14582 | w14583);
assign w14584 = v6780;
assign w14585 = w14577 & ~w14584;
assign w14586 = ~w14577 & w14584;
assign v6781 = ~(w14585 | w14586);
assign w14587 = v6781;
assign v6782 = ~(w14409 | w14413);
assign w14588 = v6782;
assign w14589 = ~w14587 & w14588;
assign w14590 = w14587 & ~w14588;
assign v6783 = ~(w14589 | w14590);
assign w14591 = v6783;
assign w14592 = w14576 & w14591;
assign v6784 = ~(w14576 | w14591);
assign w14593 = v6784;
assign v6785 = ~(w14592 | w14593);
assign w14594 = v6785;
assign w14595 = w14549 & w14594;
assign v6786 = ~(w14549 | w14594);
assign w14596 = v6786;
assign v6787 = ~(w14595 | w14596);
assign w14597 = v6787;
assign v6788 = ~(w14507 | w14510);
assign w14598 = v6788;
assign v6789 = ~(w14455 | w14484);
assign w14599 = v6789;
assign v6790 = ~(w14501 | w14504);
assign w14600 = v6790;
assign w14601 = pi39 & pi57;
assign w14602 = pi38 & pi58;
assign v6791 = ~(w14601 | w14602);
assign w14603 = v6791;
assign w14604 = pi39 & pi58;
assign w14605 = w14462 & w14604;
assign v6792 = ~(w14603 | w14605);
assign w14606 = v6792;
assign w14607 = w14446 & ~w14606;
assign w14608 = ~w14446 & w14606;
assign v6793 = ~(w14607 | w14608);
assign w14609 = v6793;
assign w14610 = pi37 & pi59;
assign w14611 = pi40 & pi56;
assign v6794 = ~(w14610 | w14611);
assign w14612 = v6794;
assign w14613 = w14610 & w14611;
assign v6795 = ~(w14612 | w14613);
assign w14614 = v6795;
assign w14615 = w14400 & ~w14614;
assign w14616 = ~w14400 & w14614;
assign v6796 = ~(w14615 | w14616);
assign w14617 = v6796;
assign v6797 = ~(w14609 | w14617);
assign w14618 = v6797;
assign w14619 = w14609 & w14617;
assign v6798 = ~(w14618 | w14619);
assign w14620 = v6798;
assign w14621 = pi45 & pi51;
assign w14622 = pi47 & pi49;
assign v6799 = ~(w14430 | w14622);
assign w14623 = v6799;
assign w14624 = pi47 & pi50;
assign w14625 = w14427 & w14624;
assign v6800 = ~(w14623 | w14625);
assign w14626 = v6800;
assign w14627 = w14621 & ~w14626;
assign w14628 = ~w14621 & w14626;
assign v6801 = ~(w14627 | w14628);
assign w14629 = v6801;
assign w14630 = w14620 & ~w14629;
assign w14631 = ~w14620 & w14629;
assign v6802 = ~(w14630 | w14631);
assign w14632 = v6802;
assign w14633 = ~w14600 & w14632;
assign w14634 = w14600 & ~w14632;
assign v6803 = ~(w14633 | w14634);
assign w14635 = v6803;
assign w14636 = ~w14599 & w14635;
assign w14637 = w14599 & ~w14635;
assign v6804 = ~(w14636 | w14637);
assign w14638 = v6804;
assign w14639 = ~w14598 & w14638;
assign w14640 = w14598 & ~w14638;
assign v6805 = ~(w14639 | w14640);
assign w14641 = v6805;
assign w14642 = w14597 & w14641;
assign v6806 = ~(w14597 | w14641);
assign w14643 = v6806;
assign v6807 = ~(w14642 | w14643);
assign w14644 = v6807;
assign w14645 = ~w14525 & w14644;
assign w14646 = w14525 & ~w14644;
assign v6808 = ~(w14645 | w14646);
assign w14647 = v6808;
assign w14648 = (w11122 & w17656) | (w11122 & w17657) | (w17656 & w17657);
assign w14649 = (~w11122 & w17658) | (~w11122 & w17659) | (w17658 & w17659);
assign v6809 = ~(w14648 | w14649);
assign w14650 = v6809;
assign v6810 = ~(w14639 | w14642);
assign w14651 = v6810;
assign v6811 = ~(w14633 | w14636);
assign w14652 = v6811;
assign w14653 = pi36 & pi61;
assign w14654 = w14621 & ~w14623;
assign w14655 = (w14653 & w14654) | (w14653 & w16781) | (w14654 & w16781);
assign w14656 = ~w14654 & w16782;
assign v6812 = ~(w14655 | w14656);
assign w14657 = v6812;
assign w14658 = w14446 & ~w14603;
assign v6813 = ~(w14605 | w14658);
assign w14659 = v6813;
assign w14660 = ~w14657 & w14659;
assign w14661 = w14657 & ~w14659;
assign v6814 = ~(w14660 | w14661);
assign w14662 = v6814;
assign v6815 = ~(w14618 | w14630);
assign w14663 = v6815;
assign v6816 = ~(w14582 | w14586);
assign w14664 = v6816;
assign v6817 = ~(w14663 | w14664);
assign w14665 = v6817;
assign w14666 = w14663 & w14664;
assign v6818 = ~(w14665 | w14666);
assign w14667 = v6818;
assign w14668 = w14662 & w14667;
assign v6819 = ~(w14662 | w14667);
assign w14669 = v6819;
assign v6820 = ~(w14668 | w14669);
assign w14670 = v6820;
assign w14671 = (~w14531 & ~w14533) | (~w14531 & w16783) | (~w14533 & w16783);
assign w14672 = pi40 & pi57;
assign w14673 = pi46 & pi51;
assign v6821 = ~(w14624 | w14673);
assign w14674 = v6821;
assign w14675 = pi47 & pi51;
assign w14676 = w14430 & w14675;
assign v6822 = ~(w14674 | w14676);
assign w14677 = v6822;
assign w14678 = w14672 & ~w14677;
assign w14679 = ~w14672 & w14677;
assign v6823 = ~(w14678 | w14679);
assign w14680 = v6823;
assign w14681 = ~pi48 & pi49;
assign w14682 = w14555 & ~w14681;
assign w14683 = ~w14555 & w14681;
assign v6824 = ~(w14682 | w14683);
assign w14684 = v6824;
assign v6825 = ~(w14680 | w14684);
assign w14685 = v6825;
assign w14686 = w14680 & w14684;
assign v6826 = ~(w14685 | w14686);
assign w14687 = v6826;
assign w14688 = w14671 & ~w14687;
assign w14689 = ~w14671 & w14687;
assign v6827 = ~(w14688 | w14689);
assign w14690 = v6827;
assign v6828 = ~(w14400 | w14613);
assign w14691 = v6828;
assign v6829 = ~(w14612 | w14691);
assign w14692 = v6829;
assign w14693 = w14551 & ~w14554;
assign v6830 = ~(w14556 | w14693);
assign w14694 = v6830;
assign w14695 = w14692 & ~w14694;
assign w14696 = ~w14692 & w14694;
assign v6831 = ~(w14695 | w14696);
assign w14697 = v6831;
assign w14698 = w14561 & ~w14564;
assign v6832 = ~(w14566 | w14698);
assign w14699 = v6832;
assign w14700 = ~w14697 & w14699;
assign w14701 = w14697 & ~w14699;
assign v6833 = ~(w14700 | w14701);
assign w14702 = v6833;
assign v6834 = ~(w14571 | w14575);
assign w14703 = v6834;
assign w14704 = ~w14702 & w14703;
assign w14705 = w14702 & ~w14703;
assign v6835 = ~(w14704 | w14705);
assign w14706 = v6835;
assign w14707 = w14690 & w14706;
assign v6836 = ~(w14690 | w14706);
assign w14708 = v6836;
assign v6837 = ~(w14707 | w14708);
assign w14709 = v6837;
assign w14710 = w14670 & w14709;
assign v6838 = ~(w14670 | w14709);
assign w14711 = v6838;
assign v6839 = ~(w14710 | w14711);
assign w14712 = v6839;
assign w14713 = w14652 & ~w14712;
assign w14714 = ~w14652 & w14712;
assign v6840 = ~(w14713 | w14714);
assign w14715 = v6840;
assign v6841 = ~(w14547 | w14595);
assign w14716 = v6841;
assign v6842 = ~(w14590 | w14592);
assign w14717 = v6842;
assign v6843 = ~(w14541 | w14544);
assign w14718 = v6843;
assign w14719 = pi37 & pi60;
assign w14720 = pi38 & pi59;
assign v6844 = ~(w14604 | w14720);
assign w14721 = v6844;
assign w14722 = pi39 & pi59;
assign w14723 = w14602 & w14722;
assign v6845 = ~(w14721 | w14723);
assign w14724 = v6845;
assign w14725 = w14719 & ~w14724;
assign w14726 = ~w14719 & w14724;
assign v6846 = ~(w14725 | w14726);
assign w14727 = v6846;
assign w14728 = pi41 & pi56;
assign w14729 = pi34 & pi63;
assign w14730 = pi42 & pi55;
assign v6847 = ~(w14729 | w14730);
assign w14731 = v6847;
assign w14732 = w14729 & w14730;
assign v6848 = ~(w14731 | w14732);
assign w14733 = v6848;
assign w14734 = w14728 & ~w14733;
assign w14735 = ~w14728 & w14733;
assign v6849 = ~(w14734 | w14735);
assign w14736 = v6849;
assign v6850 = ~(w14727 | w14736);
assign w14737 = v6850;
assign w14738 = w14727 & w14736;
assign v6851 = ~(w14737 | w14738);
assign w14739 = v6851;
assign w14740 = pi45 & pi52;
assign w14741 = pi44 & pi53;
assign v6852 = ~(w14740 | w14741);
assign w14742 = v6852;
assign w14743 = pi45 & pi53;
assign w14744 = w14446 & w14743;
assign v6853 = ~(w14742 | w14744);
assign w14745 = v6853;
assign w14746 = w14565 & ~w14745;
assign w14747 = ~w14565 & w14745;
assign v6854 = ~(w14746 | w14747);
assign w14748 = v6854;
assign w14749 = w14739 & ~w14748;
assign w14750 = ~w14739 & w14748;
assign v6855 = ~(w14749 | w14750);
assign w14751 = v6855;
assign w14752 = ~w14718 & w14751;
assign w14753 = w14718 & ~w14751;
assign v6856 = ~(w14752 | w14753);
assign w14754 = v6856;
assign w14755 = ~w14717 & w14754;
assign w14756 = w14717 & ~w14754;
assign v6857 = ~(w14755 | w14756);
assign w14757 = v6857;
assign w14758 = ~w14716 & w14757;
assign w14759 = w14716 & ~w14757;
assign v6858 = ~(w14758 | w14759);
assign w14760 = v6858;
assign w14761 = w14715 & w14760;
assign v6859 = ~(w14715 | w14760);
assign w14762 = v6859;
assign v6860 = ~(w14761 | w14762);
assign w14763 = v6860;
assign w14764 = ~w14651 & w14763;
assign w14765 = w14651 & ~w14763;
assign v6861 = ~(w14764 | w14765);
assign w14766 = v6861;
assign w14767 = (~w12329 & w17505) | (~w12329 & w17506) | (w17505 & w17506);
assign w14768 = (w12329 & w17507) | (w12329 & w17508) | (w17507 & w17508);
assign v6862 = ~(w14767 | w14768);
assign w14769 = v6862;
assign v6863 = ~(w14758 | w14761);
assign w14770 = v6863;
assign v6864 = ~(w14710 | w14714);
assign w14771 = v6864;
assign v6865 = ~(w14705 | w14707);
assign w14772 = v6865;
assign w14773 = pi44 & pi54;
assign w14774 = pi43 & pi55;
assign v6866 = ~(w14773 | w14774);
assign w14775 = v6866;
assign w14776 = pi44 & pi55;
assign w14777 = w14565 & w14776;
assign v6867 = ~(w14775 | w14777);
assign w14778 = v6867;
assign w14779 = pi35 & pi63;
assign w14780 = ~w14778 & w14779;
assign w14781 = w14778 & ~w14779;
assign v6868 = ~(w14780 | w14781);
assign w14782 = v6868;
assign w14783 = w14672 & ~w14674;
assign v6869 = ~(w14676 | w14783);
assign w14784 = v6869;
assign v6870 = ~(w14782 | w14784);
assign w14785 = v6870;
assign w14786 = w14782 & w14784;
assign v6871 = ~(w14785 | w14786);
assign w14787 = v6871;
assign w14788 = pi38 & pi60;
assign w14789 = pi42 & pi56;
assign w14790 = pi41 & pi57;
assign v6872 = ~(w14789 | w14790);
assign w14791 = v6872;
assign w14792 = pi42 & pi57;
assign w14793 = w14728 & w14792;
assign v6873 = ~(w14791 | w14793);
assign w14794 = v6873;
assign w14795 = w14788 & ~w14794;
assign w14796 = ~w14788 & w14794;
assign v6874 = ~(w14795 | w14796);
assign w14797 = v6874;
assign w14798 = ~w14787 & w14797;
assign w14799 = w14787 & ~w14797;
assign v6875 = ~(w14798 | w14799);
assign w14800 = v6875;
assign v6876 = ~(w14665 | w14668);
assign w14801 = v6876;
assign w14802 = w14800 & ~w14801;
assign w14803 = ~w14800 & w14801;
assign v6877 = ~(w14802 | w14803);
assign w14804 = v6877;
assign w14805 = ~w14772 & w14804;
assign w14806 = w14772 & ~w14804;
assign v6878 = ~(w14805 | w14806);
assign w14807 = v6878;
assign w14808 = ~w14771 & w14807;
assign w14809 = w14771 & ~w14807;
assign v6879 = ~(w14808 | w14809);
assign w14810 = v6879;
assign v6880 = ~(w14752 | w14755);
assign w14811 = v6880;
assign w14812 = (~w14737 & ~w14739) | (~w14737 & w16963) | (~w14739 & w16963);
assign w14813 = (~w14695 & ~w14697) | (~w14695 & w16784) | (~w14697 & w16784);
assign w14814 = (~w14655 & ~w14657) | (~w14655 & w16964) | (~w14657 & w16964);
assign v6881 = ~(w14813 | w14814);
assign w14815 = v6881;
assign w14816 = w14813 & w14814;
assign v6882 = ~(w14815 | w14816);
assign w14817 = v6882;
assign w14818 = w14812 & ~w14817;
assign w14819 = ~w14812 & w14817;
assign v6883 = ~(w14818 | w14819);
assign w14820 = v6883;
assign v6884 = ~(w14728 | w14732);
assign w14821 = v6884;
assign v6885 = ~(w14731 | w14821);
assign w14822 = v6885;
assign w14823 = w14719 & ~w14721;
assign v6886 = ~(w14723 | w14823);
assign w14824 = v6886;
assign w14825 = w14822 & ~w14824;
assign w14826 = ~w14822 & w14824;
assign v6887 = ~(w14825 | w14826);
assign w14827 = v6887;
assign w14828 = w14565 & ~w14742;
assign v6888 = ~(w14744 | w14828);
assign w14829 = v6888;
assign w14830 = ~w14827 & w14829;
assign w14831 = w14827 & ~w14829;
assign v6889 = ~(w14830 | w14831);
assign w14832 = v6889;
assign v6890 = ~(w14685 | w14689);
assign w14833 = v6890;
assign w14834 = ~w14832 & w14833;
assign w14835 = w14832 & ~w14833;
assign v6891 = ~(w14834 | w14835);
assign w14836 = v6891;
assign w14837 = pi36 & pi62;
assign w14838 = pi37 & pi61;
assign v6892 = ~(w14837 | w14838);
assign w14839 = v6892;
assign w14840 = pi37 & pi62;
assign w14841 = w14653 & w14840;
assign v6893 = ~(w14839 | w14841);
assign w14842 = v6893;
assign w14843 = (pi49 & w14555) | (pi49 & w16965) | (w14555 & w16965);
assign w14844 = w14842 & w14843;
assign v6894 = ~(w14842 | w14843);
assign w14845 = v6894;
assign v6895 = ~(w14844 | w14845);
assign w14846 = v6895;
assign w14847 = pi46 & pi52;
assign w14848 = pi48 & pi50;
assign v6896 = ~(w14675 | w14848);
assign w14849 = v6896;
assign w14850 = pi48 & pi51;
assign w14851 = w14624 & w14850;
assign v6897 = ~(w14849 | w14851);
assign w14852 = v6897;
assign w14853 = w14847 & ~w14852;
assign w14854 = ~w14847 & w14852;
assign v6898 = ~(w14853 | w14854);
assign w14855 = v6898;
assign w14856 = pi40 & pi58;
assign v6899 = ~(w14722 | w14856);
assign w14857 = v6899;
assign w14858 = pi40 & pi59;
assign w14859 = w14604 & w14858;
assign v6900 = ~(w14857 | w14859);
assign w14860 = v6900;
assign w14861 = w14743 & ~w14860;
assign w14862 = ~w14743 & w14860;
assign v6901 = ~(w14861 | w14862);
assign w14863 = v6901;
assign v6902 = ~(w14855 | w14863);
assign w14864 = v6902;
assign w14865 = w14855 & w14863;
assign v6903 = ~(w14864 | w14865);
assign w14866 = v6903;
assign w14867 = w14846 & w14866;
assign v6904 = ~(w14846 | w14866);
assign w14868 = v6904;
assign v6905 = ~(w14867 | w14868);
assign w14869 = v6905;
assign v6906 = ~(w14836 | w14869);
assign w14870 = v6906;
assign w14871 = w14836 & w14869;
assign v6907 = ~(w14870 | w14871);
assign w14872 = v6907;
assign v6908 = ~(w14820 | w14872);
assign w14873 = v6908;
assign w14874 = w14820 & w14872;
assign v6909 = ~(w14873 | w14874);
assign w14875 = v6909;
assign w14876 = w14811 & ~w14875;
assign w14877 = ~w14811 & w14875;
assign v6910 = ~(w14876 | w14877);
assign w14878 = v6910;
assign w14879 = w14810 & w14878;
assign v6911 = ~(w14810 | w14878);
assign w14880 = v6911;
assign v6912 = ~(w14879 | w14880);
assign w14881 = v6912;
assign w14882 = w14770 & ~w14881;
assign w14883 = ~w14770 & w14881;
assign v6913 = ~(w14882 | w14883);
assign w14884 = v6913;
assign v6914 = ~(w14646 | w14765);
assign w14885 = v6914;
assign w14886 = (w12329 & w17509) | (w12329 & w17510) | (w17509 & w17510);
assign w14887 = (~w12329 & w17511) | (~w12329 & w17512) | (w17511 & w17512);
assign v6915 = ~(w14886 | w14887);
assign w14888 = v6915;
assign v6916 = ~(w14808 | w14879);
assign w14889 = v6916;
assign v6917 = ~(w14802 | w14805);
assign w14890 = v6917;
assign w14891 = (~w14785 & ~w14787) | (~w14785 & w16966) | (~w14787 & w16966);
assign w14892 = (~w14825 & ~w14827) | (~w14825 & w16785) | (~w14827 & w16785);
assign w14893 = ~pi49 & pi50;
assign w14894 = w14840 & ~w14893;
assign w14895 = ~w14840 & w14893;
assign v6918 = ~(w14894 | w14895);
assign w14896 = v6918;
assign v6919 = ~(w14892 | w14896);
assign w14897 = v6919;
assign w14898 = w14892 & w14896;
assign v6920 = ~(w14897 | w14898);
assign w14899 = v6920;
assign w14900 = w14891 & ~w14899;
assign w14901 = ~w14891 & w14899;
assign v6921 = ~(w14900 | w14901);
assign w14902 = v6921;
assign w14903 = (~w14841 & ~w14842) | (~w14841 & w16967) | (~w14842 & w16967);
assign w14904 = w14788 & ~w14791;
assign v6922 = ~(w14793 | w14904);
assign w14905 = v6922;
assign v6923 = ~(w14903 | w14905);
assign w14906 = v6923;
assign w14907 = w14903 & w14905;
assign v6924 = ~(w14906 | w14907);
assign w14908 = v6924;
assign w14909 = pi36 & pi63;
assign w14910 = pi39 & pi60;
assign w14911 = pi38 & pi61;
assign v6925 = ~(w14910 | w14911);
assign w14912 = v6925;
assign w14913 = pi39 & pi61;
assign w14914 = w14788 & w14913;
assign v6926 = ~(w14912 | w14914);
assign w14915 = v6926;
assign w14916 = w14909 & ~w14915;
assign w14917 = ~w14909 & w14915;
assign v6927 = ~(w14916 | w14917);
assign w14918 = v6927;
assign w14919 = ~w14908 & w14918;
assign w14920 = w14908 & ~w14918;
assign v6928 = ~(w14919 | w14920);
assign w14921 = v6928;
assign w14922 = w14743 & ~w14857;
assign v6929 = ~(w14859 | w14922);
assign w14923 = v6929;
assign w14924 = w14847 & ~w14849;
assign v6930 = ~(w14851 | w14924);
assign w14925 = v6930;
assign v6931 = ~(w14923 | w14925);
assign w14926 = v6931;
assign w14927 = w14923 & w14925;
assign v6932 = ~(w14926 | w14927);
assign w14928 = v6932;
assign w14929 = ~w14775 & w14779;
assign v6933 = ~(w14777 | w14929);
assign w14930 = v6933;
assign w14931 = ~w14928 & w14930;
assign w14932 = w14928 & ~w14930;
assign v6934 = ~(w14931 | w14932);
assign w14933 = v6934;
assign w14934 = (~w14864 & ~w14866) | (~w14864 & w16968) | (~w14866 & w16968);
assign w14935 = ~w14933 & w14934;
assign w14936 = w14933 & ~w14934;
assign v6935 = ~(w14935 | w14936);
assign w14937 = v6935;
assign w14938 = w14921 & w14937;
assign v6936 = ~(w14921 | w14937);
assign w14939 = v6936;
assign v6937 = ~(w14938 | w14939);
assign w14940 = v6937;
assign v6938 = ~(w14902 | w14940);
assign w14941 = v6938;
assign w14942 = w14902 & w14940;
assign v6939 = ~(w14941 | w14942);
assign w14943 = v6939;
assign w14944 = ~w14890 & w14943;
assign w14945 = w14890 & ~w14943;
assign v6940 = ~(w14944 | w14945);
assign w14946 = v6940;
assign w14947 = (~w14835 & ~w14836) | (~w14835 & w16969) | (~w14836 & w16969);
assign w14948 = (~w14815 & ~w14817) | (~w14815 & w16970) | (~w14817 & w16970);
assign w14949 = pi45 & pi54;
assign w14950 = pi47 & pi52;
assign w14951 = pi46 & pi53;
assign v6941 = ~(w14950 | w14951);
assign w14952 = v6941;
assign w14953 = pi47 & pi53;
assign w14954 = w14847 & w14953;
assign v6942 = ~(w14952 | w14954);
assign w14955 = v6942;
assign w14956 = w14949 & ~w14955;
assign w14957 = ~w14949 & w14955;
assign v6943 = ~(w14956 | w14957);
assign w14958 = v6943;
assign w14959 = pi41 & pi58;
assign v6944 = ~(w14776 | w14959);
assign w14960 = v6944;
assign w14961 = w14776 & w14959;
assign v6945 = ~(w14960 | w14961);
assign w14962 = v6945;
assign w14963 = w14858 & ~w14962;
assign w14964 = ~w14858 & w14962;
assign v6946 = ~(w14963 | w14964);
assign w14965 = v6946;
assign v6947 = ~(w14958 | w14965);
assign w14966 = v6947;
assign w14967 = w14958 & w14965;
assign v6948 = ~(w14966 | w14967);
assign w14968 = v6948;
assign w14969 = pi43 & pi56;
assign v6949 = ~(w14792 | w14969);
assign w14970 = v6949;
assign w14971 = pi43 & pi57;
assign w14972 = w14789 & w14971;
assign v6950 = ~(w14970 | w14972);
assign w14973 = v6950;
assign w14974 = w14850 & ~w14973;
assign w14975 = ~w14850 & w14973;
assign v6951 = ~(w14974 | w14975);
assign w14976 = v6951;
assign w14977 = w14968 & ~w14976;
assign w14978 = ~w14968 & w14976;
assign v6952 = ~(w14977 | w14978);
assign w14979 = v6952;
assign w14980 = ~w14948 & w14979;
assign w14981 = w14948 & ~w14979;
assign v6953 = ~(w14980 | w14981);
assign w14982 = v6953;
assign w14983 = w14947 & ~w14982;
assign w14984 = ~w14947 & w14982;
assign v6954 = ~(w14983 | w14984);
assign w14985 = v6954;
assign v6955 = ~(w14874 | w14877);
assign w14986 = v6955;
assign w14987 = w14985 & ~w14986;
assign w14988 = ~w14985 & w14986;
assign v6956 = ~(w14987 | w14988);
assign w14989 = v6956;
assign w14990 = w14946 & w14989;
assign v6957 = ~(w14946 | w14989);
assign w14991 = v6957;
assign v6958 = ~(w14990 | w14991);
assign w14992 = v6958;
assign w14993 = ~w14889 & w14992;
assign w14994 = w14889 & ~w14992;
assign v6959 = ~(w14993 | w14994);
assign w14995 = v6959;
assign v6960 = ~(w14764 | w14883);
assign w14996 = v6960;
assign w14997 = (w11122 & w17660) | (w11122 & w17661) | (w17660 & w17661);
assign w14998 = (~w11122 & w17662) | (~w11122 & w17663) | (w17662 & w17663);
assign v6961 = ~(w14997 | w14998);
assign w14999 = v6961;
assign v6962 = ~(w14987 | w14990);
assign w15000 = v6962;
assign w15001 = (~w14906 & ~w14908) | (~w14906 & w17237) | (~w14908 & w17237);
assign w15002 = (~w14926 & ~w14928) | (~w14926 & w16786) | (~w14928 & w16786);
assign w15003 = pi49 & pi51;
assign w15004 = pi48 & pi52;
assign v6963 = ~(w15003 | w15004);
assign w15005 = v6963;
assign w15006 = pi49 & pi52;
assign w15007 = w14850 & w15006;
assign v6964 = ~(w15005 | w15007);
assign w15008 = v6964;
assign w15009 = w14953 & ~w15008;
assign w15010 = ~w14953 & w15008;
assign v6965 = ~(w15009 | w15010);
assign w15011 = v6965;
assign v6966 = ~(w15002 | w15011);
assign w15012 = v6966;
assign w15013 = w15002 & w15011;
assign v6967 = ~(w15012 | w15013);
assign w15014 = v6967;
assign w15015 = w15001 & ~w15014;
assign w15016 = ~w15001 & w15014;
assign v6968 = ~(w15015 | w15016);
assign w15017 = v6968;
assign w15018 = ~w14984 & w17238;
assign w15019 = (w15017 & w14984) | (w15017 & w17239) | (w14984 & w17239);
assign v6969 = ~(w15018 | w15019);
assign w15020 = v6969;
assign w15021 = w14909 & ~w14912;
assign v6970 = ~(w14914 | w15021);
assign w15022 = v6970;
assign w15023 = w14949 & ~w14952;
assign v6971 = ~(w14954 | w15023);
assign w15024 = v6971;
assign v6972 = ~(w15022 | w15024);
assign w15025 = v6972;
assign w15026 = w15022 & w15024;
assign v6973 = ~(w15025 | w15026);
assign w15027 = v6973;
assign v6974 = ~(w14858 | w14961);
assign w15028 = v6974;
assign v6975 = ~(w14960 | w15028);
assign w15029 = v6975;
assign v6976 = ~(w15027 | w15029);
assign w15030 = v6976;
assign w15031 = w15027 & w15029;
assign v6977 = ~(w15030 | w15031);
assign w15032 = v6977;
assign v6978 = ~(w14966 | w14977);
assign w15033 = v6978;
assign w15034 = ~w15032 & w15033;
assign w15035 = w15032 & ~w15033;
assign v6979 = ~(w15034 | w15035);
assign w15036 = v6979;
assign w15037 = pi37 & pi63;
assign v6980 = ~(pi49 | w14840);
assign w15038 = v6980;
assign w15039 = pi50 & ~w15038;
assign w15040 = w15037 & w15039;
assign v6981 = ~(w15037 | w15039);
assign w15041 = v6981;
assign v6982 = ~(w15040 | w15041);
assign w15042 = v6982;
assign w15043 = w14850 & ~w14970;
assign v6983 = ~(w14972 | w15043);
assign w15044 = v6983;
assign w15045 = ~w15042 & w15044;
assign w15046 = w15042 & ~w15044;
assign v6984 = ~(w15045 | w15046);
assign w15047 = v6984;
assign w15048 = w15036 & w15047;
assign v6985 = ~(w15036 | w15047);
assign w15049 = v6985;
assign v6986 = ~(w15048 | w15049);
assign w15050 = v6986;
assign w15051 = w15020 & w15050;
assign v6987 = ~(w15020 | w15050);
assign w15052 = v6987;
assign v6988 = ~(w15051 | w15052);
assign w15053 = v6988;
assign v6989 = ~(w14942 | w14944);
assign w15054 = v6989;
assign w15055 = (~w14936 & ~w14937) | (~w14936 & w17240) | (~w14937 & w17240);
assign w15056 = (~w14897 & ~w14899) | (~w14897 & w16971) | (~w14899 & w16971);
assign w15057 = pi45 & pi55;
assign w15058 = pi44 & pi56;
assign v6990 = ~(w15057 | w15058);
assign w15059 = v6990;
assign w15060 = pi45 & pi56;
assign w15061 = w14776 & w15060;
assign v6991 = ~(w15059 | w15061);
assign w15062 = v6991;
assign w15063 = w14971 & ~w15062;
assign w15064 = ~w14971 & w15062;
assign v6992 = ~(w15063 | w15064);
assign w15065 = v6992;
assign w15066 = pi38 & pi62;
assign w15067 = pi40 & pi60;
assign v6993 = ~(w14913 | w15067);
assign w15068 = v6993;
assign w15069 = pi40 & pi61;
assign w15070 = w14910 & w15069;
assign v6994 = ~(w15068 | w15070);
assign w15071 = v6994;
assign w15072 = w15066 & ~w15071;
assign w15073 = ~w15066 & w15071;
assign v6995 = ~(w15072 | w15073);
assign w15074 = v6995;
assign v6996 = ~(w15065 | w15074);
assign w15075 = v6996;
assign w15076 = w15065 & w15074;
assign v6997 = ~(w15075 | w15076);
assign w15077 = v6997;
assign w15078 = pi46 & pi54;
assign w15079 = pi42 & pi58;
assign w15080 = pi41 & pi59;
assign v6998 = ~(w15079 | w15080);
assign w15081 = v6998;
assign w15082 = pi42 & pi59;
assign w15083 = w14959 & w15082;
assign v6999 = ~(w15081 | w15083);
assign w15084 = v6999;
assign w15085 = w15078 & ~w15084;
assign w15086 = ~w15078 & w15084;
assign v7000 = ~(w15085 | w15086);
assign w15087 = v7000;
assign w15088 = w15077 & ~w15087;
assign w15089 = ~w15077 & w15087;
assign v7001 = ~(w15088 | w15089);
assign w15090 = v7001;
assign w15091 = ~w15056 & w15090;
assign w15092 = w15056 & ~w15090;
assign v7002 = ~(w15091 | w15092);
assign w15093 = v7002;
assign w15094 = ~w15055 & w15093;
assign w15095 = w15055 & ~w15093;
assign v7003 = ~(w15094 | w15095);
assign w15096 = v7003;
assign w15097 = ~w15054 & w15096;
assign w15098 = w15054 & ~w15096;
assign v7004 = ~(w15097 | w15098);
assign w15099 = v7004;
assign w15100 = w15053 & w15099;
assign v7005 = ~(w15053 | w15099);
assign w15101 = v7005;
assign v7006 = ~(w15100 | w15101);
assign w15102 = v7006;
assign w15103 = ~w15000 & w15102;
assign w15104 = w15000 & ~w15102;
assign v7007 = ~(w15103 | w15104);
assign w15105 = v7007;
assign w15106 = (~w12329 & w17513) | (~w12329 & w17514) | (w17513 & w17514);
assign w15107 = (w12329 & w17515) | (w12329 & w17516) | (w17515 & w17516);
assign v7008 = ~(w15106 | w15107);
assign w15108 = v7008;
assign v7009 = ~(w14994 | w15104);
assign w15109 = v7009;
assign v7010 = ~(w15097 | w15100);
assign w15110 = v7010;
assign v7011 = ~(w15019 | w15051);
assign w15111 = v7011;
assign w15112 = (~w15012 & ~w15014) | (~w15012 & w16972) | (~w15014 & w16972);
assign w15113 = pi38 & pi63;
assign w15114 = pi47 & pi54;
assign w15115 = pi46 & pi55;
assign v7012 = ~(w15114 | w15115);
assign w15116 = v7012;
assign w15117 = pi47 & pi55;
assign w15118 = w15078 & w15117;
assign v7013 = ~(w15116 | w15118);
assign w15119 = v7013;
assign w15120 = w15113 & ~w15119;
assign w15121 = ~w15113 & w15119;
assign v7014 = ~(w15120 | w15121);
assign w15122 = v7014;
assign w15123 = pi43 & pi58;
assign v7015 = ~(w15060 | w15123);
assign w15124 = v7015;
assign w15125 = w15060 & w15123;
assign v7016 = ~(w15124 | w15125);
assign w15126 = v7016;
assign w15127 = w15082 & ~w15126;
assign w15128 = ~w15082 & w15126;
assign v7017 = ~(w15127 | w15128);
assign w15129 = v7017;
assign v7018 = ~(w15122 | w15129);
assign w15130 = v7018;
assign w15131 = w15122 & w15129;
assign v7019 = ~(w15130 | w15131);
assign w15132 = v7019;
assign w15133 = pi48 & pi53;
assign w15134 = pi44 & pi57;
assign v7020 = ~(w15006 | w15134);
assign w15135 = v7020;
assign w15136 = w15006 & w15134;
assign v7021 = ~(w15135 | w15136);
assign w15137 = v7021;
assign w15138 = w15133 & ~w15137;
assign w15139 = ~w15133 & w15137;
assign v7022 = ~(w15138 | w15139);
assign w15140 = v7022;
assign w15141 = w15132 & ~w15140;
assign w15142 = ~w15132 & w15140;
assign v7023 = ~(w15141 | w15142);
assign w15143 = v7023;
assign w15144 = ~w15112 & w15143;
assign w15145 = w15112 & ~w15143;
assign v7024 = ~(w15144 | w15145);
assign w15146 = v7024;
assign v7025 = ~(w15040 | w15046);
assign w15147 = v7025;
assign w15148 = pi41 & pi60;
assign v7026 = ~(w15069 | w15148);
assign w15149 = v7026;
assign w15150 = pi41 & pi61;
assign w15151 = w15067 & w15150;
assign v7027 = ~(w15149 | w15151);
assign w15152 = v7027;
assign w15153 = w14953 & ~w15005;
assign v7028 = ~(w15007 | w15153);
assign w15154 = v7028;
assign w15155 = w15152 & ~w15154;
assign w15156 = ~w15152 & w15154;
assign v7029 = ~(w15155 | w15156);
assign w15157 = v7029;
assign w15158 = pi39 & pi62;
assign w15159 = ~pi50 & pi51;
assign w15160 = w15158 & ~w15159;
assign w15161 = ~w15158 & w15159;
assign v7030 = ~(w15160 | w15161);
assign w15162 = v7030;
assign w15163 = w15157 & ~w15162;
assign w15164 = ~w15157 & w15162;
assign v7031 = ~(w15163 | w15164);
assign w15165 = v7031;
assign w15166 = ~w15147 & w15165;
assign w15167 = w15147 & ~w15165;
assign v7032 = ~(w15166 | w15167);
assign w15168 = v7032;
assign w15169 = w15146 & w15168;
assign v7033 = ~(w15146 | w15168);
assign w15170 = v7033;
assign v7034 = ~(w15169 | w15170);
assign w15171 = v7034;
assign w15172 = ~w15111 & w15171;
assign w15173 = w15111 & ~w15171;
assign v7035 = ~(w15172 | w15173);
assign w15174 = v7035;
assign w15175 = w15066 & ~w15068;
assign v7036 = ~(w15070 | w15175);
assign w15176 = v7036;
assign w15177 = w15078 & ~w15081;
assign v7037 = ~(w15083 | w15177);
assign w15178 = v7037;
assign v7038 = ~(w15176 | w15178);
assign w15179 = v7038;
assign w15180 = w15176 & w15178;
assign v7039 = ~(w15179 | w15180);
assign w15181 = v7039;
assign w15182 = w14971 & ~w15059;
assign v7040 = ~(w15061 | w15182);
assign w15183 = v7040;
assign w15184 = ~w15181 & w15183;
assign w15185 = w15181 & ~w15183;
assign v7041 = ~(w15184 | w15185);
assign w15186 = v7041;
assign v7042 = ~(w15075 | w15088);
assign w15187 = v7042;
assign v7043 = ~(w15025 | w15031);
assign w15188 = v7043;
assign v7044 = ~(w15187 | w15188);
assign w15189 = v7044;
assign w15190 = w15187 & w15188;
assign v7045 = ~(w15189 | w15190);
assign w15191 = v7045;
assign w15192 = w15186 & w15191;
assign v7046 = ~(w15186 | w15191);
assign w15193 = v7046;
assign v7047 = ~(w15192 | w15193);
assign w15194 = v7047;
assign w15195 = (~w15091 & ~w15093) | (~w15091 & w17245) | (~w15093 & w17245);
assign v7048 = ~(w15035 | w15048);
assign w15196 = v7048;
assign v7049 = ~(w15195 | w15196);
assign w15197 = v7049;
assign w15198 = w15195 & w15196;
assign v7050 = ~(w15197 | w15198);
assign w15199 = v7050;
assign w15200 = w15194 & w15199;
assign v7051 = ~(w15194 | w15199);
assign w15201 = v7051;
assign v7052 = ~(w15200 | w15201);
assign w15202 = v7052;
assign w15203 = w15174 & w15202;
assign v7053 = ~(w15174 | w15202);
assign w15204 = v7053;
assign v7054 = ~(w15203 | w15204);
assign w15205 = v7054;
assign w15206 = ~w15110 & w15205;
assign w15207 = w15110 & ~w15205;
assign v7055 = ~(w15206 | w15207);
assign w15208 = v7055;
assign w15209 = (w12329 & w17517) | (w12329 & w17518) | (w17517 & w17518);
assign w15210 = (~w12329 & w17519) | (~w12329 & w17520) | (w17519 & w17520);
assign v7056 = ~(w15209 | w15210);
assign w15211 = v7056;
assign v7057 = ~(w15103 | w15206);
assign w15212 = v7057;
assign w15213 = (~w10008 & w17521) | (~w10008 & w17522) | (w17521 & w17522);
assign v7058 = ~(w15172 | w15203);
assign w15214 = v7058;
assign v7059 = ~(w15197 | w15200);
assign w15215 = v7059;
assign w15216 = (~w15151 & w15154) | (~w15151 & w17248) | (w15154 & w17248);
assign v7060 = ~(w15082 | w15125);
assign w15217 = v7060;
assign v7061 = ~(w15124 | w15217);
assign w15218 = v7061;
assign w15219 = ~w15216 & w15218;
assign w15220 = w15216 & ~w15218;
assign v7062 = ~(w15219 | w15220);
assign w15221 = v7062;
assign w15222 = pi39 & pi63;
assign w15223 = pi42 & pi60;
assign v7063 = ~(w15150 | w15223);
assign w15224 = v7063;
assign w15225 = pi42 & pi61;
assign w15226 = w15148 & w15225;
assign v7064 = ~(w15224 | w15226);
assign w15227 = v7064;
assign w15228 = w15222 & ~w15227;
assign w15229 = ~w15222 & w15227;
assign v7065 = ~(w15228 | w15229);
assign w15230 = v7065;
assign w15231 = ~w15221 & w15230;
assign w15232 = w15221 & ~w15230;
assign v7066 = ~(w15231 | w15232);
assign w15233 = v7066;
assign w15234 = (~w15163 & ~w15165) | (~w15163 & w17249) | (~w15165 & w17249);
assign w15235 = w15233 & ~w15234;
assign w15236 = ~w15233 & w15234;
assign v7067 = ~(w15235 | w15236);
assign w15237 = v7067;
assign w15238 = pi40 & pi62;
assign w15239 = pi44 & pi58;
assign w15240 = pi43 & pi59;
assign v7068 = ~(w15239 | w15240);
assign w15241 = v7068;
assign w15242 = pi44 & pi59;
assign w15243 = w15123 & w15242;
assign v7069 = ~(w15241 | w15243);
assign w15244 = v7069;
assign w15245 = w15238 & ~w15244;
assign w15246 = ~w15238 & w15244;
assign v7070 = ~(w15245 | w15246);
assign w15247 = v7070;
assign w15248 = pi45 & pi57;
assign w15249 = pi46 & pi56;
assign v7071 = ~(w15117 | w15249);
assign w15250 = v7071;
assign w15251 = pi47 & pi56;
assign w15252 = w15115 & w15251;
assign v7072 = ~(w15250 | w15252);
assign w15253 = v7072;
assign w15254 = w15248 & ~w15253;
assign w15255 = ~w15248 & w15253;
assign v7073 = ~(w15254 | w15255);
assign w15256 = v7073;
assign v7074 = ~(w15247 | w15256);
assign w15257 = v7074;
assign w15258 = w15247 & w15256;
assign v7075 = ~(w15257 | w15258);
assign w15259 = v7075;
assign w15260 = pi48 & pi54;
assign w15261 = pi49 & pi53;
assign w15262 = pi50 & pi52;
assign v7076 = ~(w15261 | w15262);
assign w15263 = v7076;
assign w15264 = pi50 & pi53;
assign w15265 = w15006 & w15264;
assign v7077 = ~(w15263 | w15265);
assign w15266 = v7077;
assign w15267 = w15260 & ~w15266;
assign w15268 = ~w15260 & w15266;
assign v7078 = ~(w15267 | w15268);
assign w15269 = v7078;
assign w15270 = w15259 & ~w15269;
assign w15271 = ~w15259 & w15269;
assign v7079 = ~(w15270 | w15271);
assign w15272 = v7079;
assign w15273 = w15237 & w15272;
assign v7080 = ~(w15237 | w15272);
assign w15274 = v7080;
assign v7081 = ~(w15273 | w15274);
assign w15275 = v7081;
assign w15276 = ~w15215 & w15275;
assign w15277 = w15215 & ~w15275;
assign v7082 = ~(w15276 | w15277);
assign w15278 = v7082;
assign v7083 = ~(pi50 | w15158);
assign w15279 = v7083;
assign w15280 = pi51 & ~w15279;
assign v7084 = ~(w15133 | w15136);
assign w15281 = v7084;
assign v7085 = ~(w15135 | w15281);
assign w15282 = v7085;
assign w15283 = w15280 & w15282;
assign v7086 = ~(w15280 | w15282);
assign w15284 = v7086;
assign v7087 = ~(w15283 | w15284);
assign w15285 = v7087;
assign w15286 = w15113 & ~w15116;
assign v7088 = ~(w15118 | w15286);
assign w15287 = v7088;
assign w15288 = ~w15285 & w15287;
assign w15289 = w15285 & ~w15287;
assign v7089 = ~(w15288 | w15289);
assign w15290 = v7089;
assign v7090 = ~(w15179 | w15185);
assign w15291 = v7090;
assign w15292 = ~w15290 & w15291;
assign w15293 = w15290 & ~w15291;
assign v7091 = ~(w15292 | w15293);
assign w15294 = v7091;
assign v7092 = ~(w15130 | w15141);
assign w15295 = v7092;
assign w15296 = ~w15294 & w15295;
assign w15297 = w15294 & ~w15295;
assign v7093 = ~(w15296 | w15297);
assign w15298 = v7093;
assign w15299 = (~w15144 & ~w15146) | (~w15144 & w17250) | (~w15146 & w17250);
assign v7094 = ~(w15189 | w15192);
assign w15300 = v7094;
assign v7095 = ~(w15299 | w15300);
assign w15301 = v7095;
assign w15302 = w15299 & w15300;
assign v7096 = ~(w15301 | w15302);
assign w15303 = v7096;
assign w15304 = w15298 & w15303;
assign v7097 = ~(w15298 | w15303);
assign w15305 = v7097;
assign v7098 = ~(w15304 | w15305);
assign w15306 = v7098;
assign w15307 = w15278 & w15306;
assign v7099 = ~(w15278 | w15306);
assign w15308 = v7099;
assign v7100 = ~(w15307 | w15308);
assign w15309 = v7100;
assign w15310 = w15214 & ~w15309;
assign w15311 = ~w15214 & w15309;
assign v7101 = ~(w15310 | w15311);
assign w15312 = v7101;
assign w15313 = (~w10008 & w17865) | (~w10008 & w17866) | (w17865 & w17866);
assign w15314 = (w10008 & w17867) | (w10008 & w17868) | (w17867 & w17868);
assign v7102 = ~(w15313 | w15314);
assign w15315 = v7102;
assign v7103 = ~(w15257 | w15270);
assign w15316 = v7103;
assign v7104 = ~(w15219 | w15232);
assign w15317 = v7104;
assign v7105 = ~(w15283 | w15289);
assign w15318 = v7105;
assign v7106 = ~(w15317 | w15318);
assign w15319 = v7106;
assign w15320 = w15317 & w15318;
assign v7107 = ~(w15319 | w15320);
assign w15321 = v7107;
assign w15322 = w15316 & ~w15321;
assign w15323 = ~w15316 & w15321;
assign v7108 = ~(w15322 | w15323);
assign w15324 = v7108;
assign v7109 = ~(w15235 | w15273);
assign w15325 = v7109;
assign v7110 = ~(w15293 | w15297);
assign w15326 = v7110;
assign v7111 = ~(w15325 | w15326);
assign w15327 = v7111;
assign w15328 = w15325 & w15326;
assign v7112 = ~(w15327 | w15328);
assign w15329 = v7112;
assign w15330 = w15324 & w15329;
assign v7113 = ~(w15324 | w15329);
assign w15331 = v7113;
assign v7114 = ~(w15330 | w15331);
assign w15332 = v7114;
assign v7115 = ~(w15301 | w15304);
assign w15333 = v7115;
assign w15334 = pi40 & pi63;
assign w15335 = w15260 & ~w15263;
assign v7116 = ~(w15265 | w15335);
assign w15336 = v7116;
assign w15337 = w15334 & ~w15336;
assign w15338 = ~w15334 & w15336;
assign v7117 = ~(w15337 | w15338);
assign w15339 = v7117;
assign w15340 = w15248 & ~w15250;
assign v7118 = ~(w15252 | w15340);
assign w15341 = v7118;
assign w15342 = ~w15339 & w15341;
assign w15343 = w15339 & ~w15341;
assign v7119 = ~(w15342 | w15343);
assign w15344 = v7119;
assign w15345 = w15222 & ~w15224;
assign v7120 = ~(w15226 | w15345);
assign w15346 = v7120;
assign w15347 = w15238 & ~w15241;
assign v7121 = ~(w15243 | w15347);
assign w15348 = v7121;
assign v7122 = ~(w15346 | w15348);
assign w15349 = v7122;
assign w15350 = w15346 & w15348;
assign v7123 = ~(w15349 | w15350);
assign w15351 = v7123;
assign w15352 = pi45 & pi58;
assign v7124 = ~(w15242 | w15352);
assign w15353 = v7124;
assign w15354 = pi45 & pi59;
assign w15355 = w15239 & w15354;
assign v7125 = ~(w15353 | w15355);
assign w15356 = v7125;
assign w15357 = w15225 & ~w15356;
assign w15358 = ~w15225 & w15356;
assign v7126 = ~(w15357 | w15358);
assign w15359 = v7126;
assign w15360 = ~w15351 & w15359;
assign w15361 = w15351 & ~w15359;
assign v7127 = ~(w15360 | w15361);
assign w15362 = v7127;
assign v7128 = ~(w15344 | w15362);
assign w15363 = v7128;
assign w15364 = w15344 & w15362;
assign v7129 = ~(w15363 | w15364);
assign w15365 = v7129;
assign w15366 = pi43 & pi60;
assign w15367 = pi46 & pi57;
assign v7130 = ~(w15251 | w15367);
assign w15368 = v7130;
assign w15369 = pi47 & pi57;
assign w15370 = w15249 & w15369;
assign v7131 = ~(w15368 | w15370);
assign w15371 = v7131;
assign w15372 = w15366 & ~w15371;
assign w15373 = ~w15366 & w15371;
assign v7132 = ~(w15372 | w15373);
assign w15374 = v7132;
assign w15375 = pi48 & pi55;
assign w15376 = pi49 & pi54;
assign v7133 = ~(w15264 | w15376);
assign w15377 = v7133;
assign w15378 = pi50 & pi54;
assign w15379 = w15261 & w15378;
assign v7134 = ~(w15377 | w15379);
assign w15380 = v7134;
assign w15381 = w15375 & ~w15380;
assign w15382 = ~w15375 & w15380;
assign v7135 = ~(w15381 | w15382);
assign w15383 = v7135;
assign v7136 = ~(w15374 | w15383);
assign w15384 = v7136;
assign w15385 = w15374 & w15383;
assign v7137 = ~(w15384 | w15385);
assign w15386 = v7137;
assign w15387 = pi41 & pi62;
assign w15388 = ~pi51 & pi52;
assign w15389 = w15387 & ~w15388;
assign w15390 = ~w15387 & w15388;
assign v7138 = ~(w15389 | w15390);
assign w15391 = v7138;
assign w15392 = w15386 & ~w15391;
assign w15393 = ~w15386 & w15391;
assign v7139 = ~(w15392 | w15393);
assign w15394 = v7139;
assign w15395 = w15365 & w15394;
assign v7140 = ~(w15365 | w15394);
assign w15396 = v7140;
assign v7141 = ~(w15395 | w15396);
assign w15397 = v7141;
assign w15398 = ~w15333 & w15397;
assign w15399 = w15333 & ~w15397;
assign v7142 = ~(w15398 | w15399);
assign w15400 = v7142;
assign w15401 = w15332 & w15400;
assign v7143 = ~(w15332 | w15400);
assign w15402 = v7143;
assign v7144 = ~(w15401 | w15402);
assign w15403 = v7144;
assign v7145 = ~(w15276 | w15307);
assign w15404 = v7145;
assign w15405 = w15403 & ~w15404;
assign w15406 = ~w15403 & w15404;
assign v7146 = ~(w15405 | w15406);
assign w15407 = v7146;
assign w15408 = (~w13978 & w17375) | (~w13978 & w17376) | (w17375 & w17376);
assign w15409 = (w13978 & w17377) | (w13978 & w17378) | (w17377 & w17378);
assign v7147 = ~(w15408 | w15409);
assign w15410 = v7147;
assign v7148 = ~(w15310 | w15406);
assign w15411 = v7148;
assign v7149 = ~(w15398 | w15401);
assign w15412 = v7149;
assign v7150 = ~(w15327 | w15330);
assign w15413 = v7150;
assign w15414 = w15366 & ~w15368;
assign v7151 = ~(w15370 | w15414);
assign w15415 = v7151;
assign w15416 = w15375 & ~w15377;
assign v7152 = ~(w15379 | w15416);
assign w15417 = v7152;
assign v7153 = ~(w15415 | w15417);
assign w15418 = v7153;
assign w15419 = w15415 & w15417;
assign v7154 = ~(w15418 | w15419);
assign w15420 = v7154;
assign w15421 = w15225 & ~w15353;
assign v7155 = ~(w15355 | w15421);
assign w15422 = v7155;
assign w15423 = ~w15420 & w15422;
assign w15424 = w15420 & ~w15422;
assign v7156 = ~(w15423 | w15424);
assign w15425 = v7156;
assign v7157 = ~(w15384 | w15392);
assign w15426 = v7157;
assign w15427 = ~w15425 & w15426;
assign w15428 = w15425 & ~w15426;
assign v7158 = ~(w15427 | w15428);
assign w15429 = v7158;
assign w15430 = pi46 & pi58;
assign w15431 = pi48 & pi56;
assign v7159 = ~(w15369 | w15431);
assign w15432 = v7159;
assign w15433 = pi48 & pi57;
assign w15434 = w15251 & w15433;
assign v7160 = ~(w15432 | w15434);
assign w15435 = v7160;
assign w15436 = w15430 & ~w15435;
assign w15437 = ~w15430 & w15435;
assign v7161 = ~(w15436 | w15437);
assign w15438 = v7161;
assign w15439 = pi44 & pi60;
assign w15440 = pi43 & pi61;
assign v7162 = ~(w15354 | w15440);
assign w15441 = v7162;
assign w15442 = w15354 & w15440;
assign v7163 = ~(w15441 | w15442);
assign w15443 = v7163;
assign w15444 = w15439 & ~w15443;
assign w15445 = ~w15439 & w15443;
assign v7164 = ~(w15444 | w15445);
assign w15446 = v7164;
assign v7165 = ~(w15438 | w15446);
assign w15447 = v7165;
assign w15448 = w15438 & w15446;
assign v7166 = ~(w15447 | w15448);
assign w15449 = v7166;
assign w15450 = pi49 & pi55;
assign w15451 = pi51 & pi53;
assign v7167 = ~(w15378 | w15451);
assign w15452 = v7167;
assign w15453 = pi51 & pi54;
assign w15454 = w15264 & w15453;
assign v7168 = ~(w15452 | w15454);
assign w15455 = v7168;
assign w15456 = w15450 & ~w15455;
assign w15457 = ~w15450 & w15455;
assign v7169 = ~(w15456 | w15457);
assign w15458 = v7169;
assign w15459 = w15449 & ~w15458;
assign w15460 = ~w15449 & w15458;
assign v7170 = ~(w15459 | w15460);
assign w15461 = v7170;
assign w15462 = w15429 & w15461;
assign v7171 = ~(w15429 | w15461);
assign w15463 = v7171;
assign v7172 = ~(w15462 | w15463);
assign w15464 = v7172;
assign w15465 = ~w15413 & w15464;
assign w15466 = w15413 & ~w15464;
assign v7173 = ~(w15465 | w15466);
assign w15467 = v7173;
assign v7174 = ~(w15337 | w15343);
assign w15468 = v7174;
assign w15469 = pi41 & pi63;
assign w15470 = pi42 & pi62;
assign v7175 = ~(w15469 | w15470);
assign w15471 = v7175;
assign w15472 = pi42 & pi63;
assign w15473 = w15387 & w15472;
assign v7176 = ~(w15471 | w15473);
assign w15474 = v7176;
assign v7177 = ~(pi51 | w15387);
assign w15475 = v7177;
assign w15476 = pi52 & ~w15475;
assign w15477 = w15474 & w15476;
assign v7178 = ~(w15474 | w15476);
assign w15478 = v7178;
assign v7179 = ~(w15477 | w15478);
assign w15479 = v7179;
assign w15480 = ~w15468 & w15479;
assign w15481 = w15468 & ~w15479;
assign v7180 = ~(w15480 | w15481);
assign w15482 = v7180;
assign v7181 = ~(w15349 | w15361);
assign w15483 = v7181;
assign w15484 = ~w15482 & w15483;
assign w15485 = w15482 & ~w15483;
assign v7182 = ~(w15484 | w15485);
assign w15486 = v7182;
assign v7183 = ~(w15364 | w15395);
assign w15487 = v7183;
assign v7184 = ~(w15319 | w15323);
assign w15488 = v7184;
assign v7185 = ~(w15487 | w15488);
assign w15489 = v7185;
assign w15490 = w15487 & w15488;
assign v7186 = ~(w15489 | w15490);
assign w15491 = v7186;
assign w15492 = w15486 & w15491;
assign v7187 = ~(w15486 | w15491);
assign w15493 = v7187;
assign v7188 = ~(w15492 | w15493);
assign w15494 = v7188;
assign w15495 = w15467 & w15494;
assign v7189 = ~(w15467 | w15494);
assign w15496 = v7189;
assign v7190 = ~(w15495 | w15496);
assign w15497 = v7190;
assign w15498 = ~w15412 & w15497;
assign w15499 = w15412 & ~w15497;
assign v7191 = ~(w15498 | w15499);
assign w15500 = v7191;
assign w15501 = (w13978 & w17379) | (w13978 & w17380) | (w17379 & w17380);
assign w15502 = (~w13978 & w17381) | (~w13978 & w17382) | (w17381 & w17382);
assign v7192 = ~(w15501 | w15502);
assign w15503 = v7192;
assign w15504 = w15430 & ~w15432;
assign v7193 = ~(w15434 | w15504);
assign w15505 = v7193;
assign w15506 = w15450 & ~w15452;
assign v7194 = ~(w15454 | w15506);
assign w15507 = v7194;
assign v7195 = ~(w15505 | w15507);
assign w15508 = v7195;
assign w15509 = w15505 & w15507;
assign v7196 = ~(w15508 | w15509);
assign w15510 = v7196;
assign v7197 = ~(w15439 | w15442);
assign w15511 = v7197;
assign v7198 = ~(w15441 | w15511);
assign w15512 = v7198;
assign v7199 = ~(w15510 | w15512);
assign w15513 = v7199;
assign w15514 = w15510 & w15512;
assign v7200 = ~(w15513 | w15514);
assign w15515 = v7200;
assign v7201 = ~(w15447 | w15459);
assign w15516 = v7201;
assign w15517 = ~w15515 & w15516;
assign w15518 = w15515 & ~w15516;
assign v7202 = ~(w15517 | w15518);
assign w15519 = v7202;
assign v7203 = ~(w15480 | w15485);
assign w15520 = v7203;
assign w15521 = ~w15519 & w15520;
assign w15522 = w15519 & ~w15520;
assign v7204 = ~(w15521 | w15522);
assign w15523 = v7204;
assign v7205 = ~(w15489 | w15492);
assign w15524 = v7205;
assign w15525 = ~w15523 & w15524;
assign w15526 = w15523 & ~w15524;
assign v7206 = ~(w15525 | w15526);
assign w15527 = v7206;
assign v7207 = ~(w15428 | w15462);
assign w15528 = v7207;
assign v7208 = ~(w15418 | w15424);
assign w15529 = v7208;
assign w15530 = pi49 & pi56;
assign w15531 = pi50 & pi55;
assign v7209 = ~(w15453 | w15531);
assign w15532 = v7209;
assign w15533 = pi51 & pi55;
assign w15534 = w15378 & w15533;
assign v7210 = ~(w15532 | w15534);
assign w15535 = v7210;
assign w15536 = w15530 & ~w15535;
assign w15537 = ~w15530 & w15535;
assign v7211 = ~(w15536 | w15537);
assign w15538 = v7211;
assign w15539 = pi43 & pi62;
assign w15540 = ~pi52 & pi53;
assign w15541 = w15539 & ~w15540;
assign w15542 = ~w15539 & w15540;
assign v7212 = ~(w15541 | w15542);
assign w15543 = v7212;
assign v7213 = ~(w15538 | w15543);
assign w15544 = v7213;
assign w15545 = w15538 & w15543;
assign v7214 = ~(w15544 | w15545);
assign w15546 = v7214;
assign w15547 = w15529 & ~w15546;
assign w15548 = ~w15529 & w15546;
assign v7215 = ~(w15547 | w15548);
assign w15549 = v7215;
assign v7216 = ~(w15473 | w15477);
assign w15550 = v7216;
assign w15551 = pi44 & pi61;
assign w15552 = pi45 & pi60;
assign v7217 = ~(w15551 | w15552);
assign w15553 = v7217;
assign w15554 = pi45 & pi61;
assign w15555 = w15439 & w15554;
assign v7218 = ~(w15553 | w15555);
assign w15556 = v7218;
assign w15557 = w15472 & ~w15556;
assign w15558 = ~w15472 & w15556;
assign v7219 = ~(w15557 | w15558);
assign w15559 = v7219;
assign v7220 = ~(w15550 | w15559);
assign w15560 = v7220;
assign w15561 = w15550 & w15559;
assign v7221 = ~(w15560 | w15561);
assign w15562 = v7221;
assign w15563 = pi46 & pi59;
assign w15564 = pi47 & pi58;
assign v7222 = ~(w15433 | w15564);
assign w15565 = v7222;
assign w15566 = pi48 & pi58;
assign w15567 = w15369 & w15566;
assign v7223 = ~(w15565 | w15567);
assign w15568 = v7223;
assign w15569 = w15563 & ~w15568;
assign w15570 = ~w15563 & w15568;
assign v7224 = ~(w15569 | w15570);
assign w15571 = v7224;
assign w15572 = w15562 & ~w15571;
assign w15573 = ~w15562 & w15571;
assign v7225 = ~(w15572 | w15573);
assign w15574 = v7225;
assign w15575 = w15549 & w15574;
assign v7226 = ~(w15549 | w15574);
assign w15576 = v7226;
assign v7227 = ~(w15575 | w15576);
assign w15577 = v7227;
assign w15578 = ~w15528 & w15577;
assign w15579 = w15528 & ~w15577;
assign v7228 = ~(w15578 | w15579);
assign w15580 = v7228;
assign w15581 = w15527 & w15580;
assign v7229 = ~(w15527 | w15580);
assign w15582 = v7229;
assign v7230 = ~(w15581 | w15582);
assign w15583 = v7230;
assign v7231 = ~(w15465 | w15495);
assign w15584 = v7231;
assign w15585 = ~w15583 & w15584;
assign w15586 = w15583 & ~w15584;
assign v7232 = ~(w15585 | w15586);
assign w15587 = v7232;
assign v7233 = ~(w15405 | w15498);
assign w15588 = v7233;
assign w15589 = (~w12329 & w17523) | (~w12329 & w17524) | (w17523 & w17524);
assign w15590 = (w12329 & w17525) | (w12329 & w17526) | (w17525 & w17526);
assign v7234 = ~(w15589 | w15590);
assign w15591 = v7234;
assign v7235 = ~(w15526 | w15581);
assign w15592 = v7235;
assign w15593 = pi43 & pi63;
assign v7236 = ~(pi52 | w15539);
assign w15594 = v7236;
assign w15595 = pi53 & ~w15594;
assign w15596 = w15593 & w15595;
assign v7237 = ~(w15593 | w15595);
assign w15597 = v7237;
assign v7238 = ~(w15596 | w15597);
assign w15598 = v7238;
assign w15599 = w15530 & ~w15532;
assign v7239 = ~(w15534 | w15599);
assign w15600 = v7239;
assign w15601 = ~w15598 & w15600;
assign w15602 = w15598 & ~w15600;
assign v7240 = ~(w15601 | w15602);
assign w15603 = v7240;
assign v7241 = ~(w15560 | w15572);
assign w15604 = v7241;
assign w15605 = ~w15603 & w15604;
assign w15606 = w15603 & ~w15604;
assign v7242 = ~(w15605 | w15606);
assign w15607 = v7242;
assign v7243 = ~(w15544 | w15548);
assign w15608 = v7243;
assign w15609 = ~w15607 & w15608;
assign w15610 = w15607 & ~w15608;
assign v7244 = ~(w15609 | w15610);
assign w15611 = v7244;
assign v7245 = ~(w15575 | w15578);
assign w15612 = v7245;
assign w15613 = ~w15611 & w15612;
assign w15614 = w15611 & ~w15612;
assign v7246 = ~(w15613 | w15614);
assign w15615 = v7246;
assign v7247 = ~(w15518 | w15522);
assign w15616 = v7247;
assign v7248 = ~(w15508 | w15514);
assign w15617 = v7248;
assign w15618 = pi47 & pi59;
assign w15619 = pi49 & pi57;
assign v7249 = ~(w15566 | w15619);
assign w15620 = v7249;
assign w15621 = pi49 & pi58;
assign w15622 = w15433 & w15621;
assign v7250 = ~(w15620 | w15622);
assign w15623 = v7250;
assign w15624 = w15618 & ~w15623;
assign w15625 = ~w15618 & w15623;
assign v7251 = ~(w15624 | w15625);
assign w15626 = v7251;
assign w15627 = pi50 & pi56;
assign w15628 = pi52 & pi54;
assign v7252 = ~(w15533 | w15628);
assign w15629 = v7252;
assign w15630 = pi52 & pi55;
assign w15631 = w15453 & w15630;
assign v7253 = ~(w15629 | w15631);
assign w15632 = v7253;
assign w15633 = w15627 & ~w15632;
assign w15634 = ~w15627 & w15632;
assign v7254 = ~(w15633 | w15634);
assign w15635 = v7254;
assign v7255 = ~(w15626 | w15635);
assign w15636 = v7255;
assign w15637 = w15626 & w15635;
assign v7256 = ~(w15636 | w15637);
assign w15638 = v7256;
assign w15639 = w15617 & ~w15638;
assign w15640 = ~w15617 & w15638;
assign v7257 = ~(w15639 | w15640);
assign w15641 = v7257;
assign w15642 = w15472 & ~w15553;
assign v7258 = ~(w15555 | w15642);
assign w15643 = v7258;
assign w15644 = w15563 & ~w15565;
assign v7259 = ~(w15567 | w15644);
assign w15645 = v7259;
assign v7260 = ~(w15643 | w15645);
assign w15646 = v7260;
assign w15647 = w15643 & w15645;
assign v7261 = ~(w15646 | w15647);
assign w15648 = v7261;
assign w15649 = pi44 & pi62;
assign w15650 = pi46 & pi60;
assign v7262 = ~(w15554 | w15650);
assign w15651 = v7262;
assign w15652 = pi46 & pi61;
assign w15653 = w15552 & w15652;
assign v7263 = ~(w15651 | w15653);
assign w15654 = v7263;
assign w15655 = w15649 & ~w15654;
assign w15656 = ~w15649 & w15654;
assign v7264 = ~(w15655 | w15656);
assign w15657 = v7264;
assign w15658 = ~w15648 & w15657;
assign w15659 = w15648 & ~w15657;
assign v7265 = ~(w15658 | w15659);
assign w15660 = v7265;
assign v7266 = ~(w15641 | w15660);
assign w15661 = v7266;
assign w15662 = w15641 & w15660;
assign v7267 = ~(w15661 | w15662);
assign w15663 = v7267;
assign w15664 = w15616 & w15663;
assign v7268 = ~(w15616 | w15663);
assign w15665 = v7268;
assign v7269 = ~(w15664 | w15665);
assign w15666 = v7269;
assign w15667 = w15615 & ~w15666;
assign w15668 = ~w15615 & w15666;
assign v7270 = ~(w15667 | w15668);
assign w15669 = v7270;
assign w15670 = ~w15592 & w15669;
assign w15671 = w15592 & ~w15669;
assign v7271 = ~(w15670 | w15671);
assign w15672 = v7271;
assign w15673 = (~w13978 & w17383) | (~w13978 & w17384) | (w17383 & w17384);
assign w15674 = (w13978 & w17385) | (w13978 & w17386) | (w17385 & w17386);
assign v7272 = ~(w15673 | w15674);
assign w15675 = v7272;
assign v7273 = ~(w15585 | w15671);
assign w15676 = v7273;
assign v7274 = ~(w15614 | w15667);
assign w15677 = v7274;
assign v7275 = ~(w15606 | w15610);
assign w15678 = v7275;
assign w15679 = w15618 & ~w15620;
assign v7276 = ~(w15622 | w15679);
assign w15680 = v7276;
assign w15681 = w15649 & ~w15651;
assign v7277 = ~(w15653 | w15681);
assign w15682 = v7277;
assign v7278 = ~(w15680 | w15682);
assign w15683 = v7278;
assign w15684 = w15680 & w15682;
assign v7279 = ~(w15683 | w15684);
assign w15685 = v7279;
assign w15686 = pi48 & pi59;
assign w15687 = pi44 & pi63;
assign v7280 = ~(w15621 | w15687);
assign w15688 = v7280;
assign w15689 = w15621 & w15687;
assign v7281 = ~(w15688 | w15689);
assign w15690 = v7281;
assign w15691 = w15686 & ~w15690;
assign w15692 = ~w15686 & w15690;
assign v7282 = ~(w15691 | w15692);
assign w15693 = v7282;
assign w15694 = ~w15685 & w15693;
assign w15695 = w15685 & ~w15693;
assign v7283 = ~(w15694 | w15695);
assign w15696 = v7283;
assign w15697 = pi47 & pi60;
assign v7284 = ~(w15652 | w15697);
assign w15698 = v7284;
assign w15699 = pi47 & pi61;
assign w15700 = w15650 & w15699;
assign v7285 = ~(w15698 | w15700);
assign w15701 = v7285;
assign w15702 = w15627 & ~w15629;
assign v7286 = ~(w15631 | w15702);
assign w15703 = v7286;
assign w15704 = w15701 & ~w15703;
assign w15705 = ~w15701 & w15703;
assign v7287 = ~(w15704 | w15705);
assign w15706 = v7287;
assign w15707 = pi50 & pi57;
assign w15708 = pi51 & pi56;
assign v7288 = ~(w15630 | w15708);
assign w15709 = v7288;
assign w15710 = pi52 & pi56;
assign w15711 = w15533 & w15710;
assign v7289 = ~(w15709 | w15711);
assign w15712 = v7289;
assign w15713 = w15707 & ~w15712;
assign w15714 = ~w15707 & w15712;
assign v7290 = ~(w15713 | w15714);
assign w15715 = v7290;
assign w15716 = pi45 & pi62;
assign w15717 = ~pi53 & pi54;
assign w15718 = w15716 & ~w15717;
assign w15719 = ~w15716 & w15717;
assign v7291 = ~(w15718 | w15719);
assign w15720 = v7291;
assign v7292 = ~(w15715 | w15720);
assign w15721 = v7292;
assign w15722 = w15715 & w15720;
assign v7293 = ~(w15721 | w15722);
assign w15723 = v7293;
assign w15724 = w15706 & w15723;
assign v7294 = ~(w15706 | w15723);
assign w15725 = v7294;
assign v7295 = ~(w15724 | w15725);
assign w15726 = v7295;
assign w15727 = w15696 & w15726;
assign v7296 = ~(w15696 | w15726);
assign w15728 = v7296;
assign v7297 = ~(w15727 | w15728);
assign w15729 = v7297;
assign w15730 = w15678 & ~w15729;
assign w15731 = ~w15678 & w15729;
assign v7298 = ~(w15730 | w15731);
assign w15732 = v7298;
assign v7299 = ~(w15636 | w15640);
assign w15733 = v7299;
assign v7300 = ~(w15646 | w15659);
assign w15734 = v7300;
assign v7301 = ~(w15596 | w15602);
assign w15735 = v7301;
assign v7302 = ~(w15734 | w15735);
assign w15736 = v7302;
assign w15737 = w15734 & w15735;
assign v7303 = ~(w15736 | w15737);
assign w15738 = v7303;
assign w15739 = w15733 & ~w15738;
assign w15740 = ~w15733 & w15738;
assign v7304 = ~(w15739 | w15740);
assign w15741 = v7304;
assign v7305 = ~(w15661 | w15664);
assign w15742 = v7305;
assign w15743 = w15741 & w15742;
assign v7306 = ~(w15741 | w15742);
assign w15744 = v7306;
assign v7307 = ~(w15743 | w15744);
assign w15745 = v7307;
assign w15746 = w15732 & w15745;
assign v7308 = ~(w15732 | w15745);
assign w15747 = v7308;
assign v7309 = ~(w15746 | w15747);
assign w15748 = v7309;
assign w15749 = w15677 & ~w15748;
assign w15750 = ~w15677 & w15748;
assign v7310 = ~(w15749 | w15750);
assign w15751 = v7310;
assign w15752 = (w13978 & w17387) | (w13978 & w17388) | (w17387 & w17388);
assign w15753 = (~w13978 & w17389) | (~w13978 & w17390) | (w17389 & w17390);
assign v7311 = ~(w15752 | w15753);
assign w15754 = v7311;
assign v7312 = ~(w15670 | w15750);
assign w15755 = v7312;
assign v7313 = ~(w15743 | w15746);
assign w15756 = v7313;
assign v7314 = ~(pi53 | w15716);
assign w15757 = v7314;
assign w15758 = pi54 & ~w15757;
assign w15759 = w15707 & ~w15709;
assign v7315 = ~(w15711 | w15759);
assign w15760 = v7315;
assign w15761 = w15758 & ~w15760;
assign w15762 = ~w15758 & w15760;
assign v7316 = ~(w15761 | w15762);
assign w15763 = v7316;
assign v7317 = ~(w15686 | w15689);
assign w15764 = v7317;
assign v7318 = ~(w15688 | w15764);
assign w15765 = v7318;
assign v7319 = ~(w15763 | w15765);
assign w15766 = v7319;
assign w15767 = w15763 & w15765;
assign v7320 = ~(w15766 | w15767);
assign w15768 = v7320;
assign v7321 = ~(w15736 | w15740);
assign w15769 = v7321;
assign w15770 = ~w15768 & w15769;
assign w15771 = w15768 & ~w15769;
assign v7322 = ~(w15770 | w15771);
assign w15772 = v7322;
assign v7323 = ~(w15700 | w15704);
assign w15773 = v7323;
assign w15774 = pi45 & pi63;
assign w15775 = pi46 & pi62;
assign v7324 = ~(w15699 | w15775);
assign w15776 = v7324;
assign w15777 = pi47 & pi62;
assign w15778 = w15652 & w15777;
assign v7325 = ~(w15776 | w15778);
assign w15779 = v7325;
assign w15780 = w15774 & ~w15779;
assign w15781 = ~w15774 & w15779;
assign v7326 = ~(w15780 | w15781);
assign w15782 = v7326;
assign v7327 = ~(w15773 | w15782);
assign w15783 = v7327;
assign w15784 = w15773 & w15782;
assign v7328 = ~(w15783 | w15784);
assign w15785 = v7328;
assign w15786 = pi48 & pi60;
assign w15787 = pi49 & pi59;
assign w15788 = pi50 & pi58;
assign v7329 = ~(w15787 | w15788);
assign w15789 = v7329;
assign w15790 = pi50 & pi59;
assign w15791 = w15621 & w15790;
assign v7330 = ~(w15789 | w15791);
assign w15792 = v7330;
assign w15793 = w15786 & ~w15792;
assign w15794 = ~w15786 & w15792;
assign v7331 = ~(w15793 | w15794);
assign w15795 = v7331;
assign w15796 = w15785 & ~w15795;
assign w15797 = ~w15785 & w15795;
assign v7332 = ~(w15796 | w15797);
assign w15798 = v7332;
assign w15799 = w15772 & w15798;
assign v7333 = ~(w15772 | w15798);
assign w15800 = v7333;
assign v7334 = ~(w15799 | w15800);
assign w15801 = v7334;
assign v7335 = ~(w15727 | w15731);
assign w15802 = v7335;
assign v7336 = ~(w15721 | w15724);
assign w15803 = v7336;
assign v7337 = ~(w15683 | w15695);
assign w15804 = v7337;
assign w15805 = pi51 & pi57;
assign w15806 = pi53 & pi55;
assign v7338 = ~(w15710 | w15806);
assign w15807 = v7338;
assign w15808 = pi53 & pi56;
assign w15809 = w15630 & w15808;
assign v7339 = ~(w15807 | w15809);
assign w15810 = v7339;
assign w15811 = w15805 & ~w15810;
assign w15812 = ~w15805 & w15810;
assign v7340 = ~(w15811 | w15812);
assign w15813 = v7340;
assign v7341 = ~(w15804 | w15813);
assign w15814 = v7341;
assign w15815 = w15804 & w15813;
assign v7342 = ~(w15814 | w15815);
assign w15816 = v7342;
assign w15817 = ~w15803 & w15816;
assign w15818 = w15803 & ~w15816;
assign v7343 = ~(w15817 | w15818);
assign w15819 = v7343;
assign w15820 = ~w15802 & w15819;
assign w15821 = w15802 & ~w15819;
assign v7344 = ~(w15820 | w15821);
assign w15822 = v7344;
assign w15823 = w15801 & w15822;
assign v7345 = ~(w15801 | w15822);
assign w15824 = v7345;
assign v7346 = ~(w15823 | w15824);
assign w15825 = v7346;
assign w15826 = w15756 & ~w15825;
assign w15827 = ~w15756 & w15825;
assign v7347 = ~(w15826 | w15827);
assign w15828 = v7347;
assign w15829 = (~w12329 & w17527) | (~w12329 & w17528) | (w17527 & w17528);
assign w15830 = (w12329 & w17529) | (w12329 & w17530) | (w17529 & w17530);
assign v7348 = ~(w15829 | w15830);
assign w15831 = v7348;
assign v7349 = ~(w15820 | w15823);
assign w15832 = v7349;
assign v7350 = ~(w15783 | w15796);
assign w15833 = v7350;
assign v7351 = ~(w15761 | w15767);
assign w15834 = v7351;
assign w15835 = ~pi54 & pi55;
assign w15836 = w15777 & ~w15835;
assign w15837 = ~w15777 & w15835;
assign v7352 = ~(w15836 | w15837);
assign w15838 = v7352;
assign v7353 = ~(w15834 | w15838);
assign w15839 = v7353;
assign w15840 = w15834 & w15838;
assign v7354 = ~(w15839 | w15840);
assign w15841 = v7354;
assign w15842 = w15833 & ~w15841;
assign w15843 = ~w15833 & w15841;
assign v7355 = ~(w15842 | w15843);
assign w15844 = v7355;
assign v7356 = ~(w15771 | w15799);
assign w15845 = v7356;
assign w15846 = ~w15844 & w15845;
assign w15847 = w15844 & ~w15845;
assign v7357 = ~(w15846 | w15847);
assign w15848 = v7357;
assign w15849 = pi46 & pi63;
assign w15850 = w15805 & ~w15807;
assign v7358 = ~(w15809 | w15850);
assign w15851 = v7358;
assign w15852 = w15849 & ~w15851;
assign w15853 = ~w15849 & w15851;
assign v7359 = ~(w15852 | w15853);
assign w15854 = v7359;
assign w15855 = w15786 & ~w15789;
assign v7360 = ~(w15791 | w15855);
assign w15856 = v7360;
assign w15857 = ~w15854 & w15856;
assign w15858 = w15854 & ~w15856;
assign v7361 = ~(w15857 | w15858);
assign w15859 = v7361;
assign v7362 = ~(w15814 | w15817);
assign w15860 = v7362;
assign w15861 = ~w15859 & w15860;
assign w15862 = w15859 & ~w15860;
assign v7363 = ~(w15861 | w15862);
assign w15863 = v7363;
assign w15864 = pi48 & pi61;
assign w15865 = pi49 & pi60;
assign v7364 = ~(w15790 | w15865);
assign w15866 = v7364;
assign w15867 = pi50 & pi60;
assign w15868 = w15787 & w15867;
assign v7365 = ~(w15866 | w15868);
assign w15869 = v7365;
assign w15870 = w15864 & ~w15869;
assign w15871 = ~w15864 & w15869;
assign v7366 = ~(w15870 | w15871);
assign w15872 = v7366;
assign w15873 = w15774 & ~w15776;
assign v7367 = ~(w15778 | w15873);
assign w15874 = v7367;
assign v7368 = ~(w15872 | w15874);
assign w15875 = v7368;
assign w15876 = w15872 & w15874;
assign v7369 = ~(w15875 | w15876);
assign w15877 = v7369;
assign w15878 = pi51 & pi58;
assign w15879 = pi52 & pi57;
assign v7370 = ~(w15808 | w15879);
assign w15880 = v7370;
assign w15881 = pi53 & pi57;
assign w15882 = w15710 & w15881;
assign v7371 = ~(w15880 | w15882);
assign w15883 = v7371;
assign w15884 = w15878 & ~w15883;
assign w15885 = ~w15878 & w15883;
assign v7372 = ~(w15884 | w15885);
assign w15886 = v7372;
assign w15887 = w15877 & ~w15886;
assign w15888 = ~w15877 & w15886;
assign v7373 = ~(w15887 | w15888);
assign w15889 = v7373;
assign w15890 = w15863 & w15889;
assign v7374 = ~(w15863 | w15889);
assign w15891 = v7374;
assign v7375 = ~(w15890 | w15891);
assign w15892 = v7375;
assign w15893 = w15848 & w15892;
assign v7376 = ~(w15848 | w15892);
assign w15894 = v7376;
assign v7377 = ~(w15893 | w15894);
assign w15895 = v7377;
assign w15896 = ~w15832 & w15895;
assign w15897 = w15832 & ~w15895;
assign v7378 = ~(w15896 | w15897);
assign w15898 = v7378;
assign w15899 = (~w13978 & w17391) | (~w13978 & w17392) | (w17391 & w17392);
assign w15900 = (w13978 & w17393) | (w13978 & w17394) | (w17393 & w17394);
assign v7379 = ~(w15899 | w15900);
assign w15901 = v7379;
assign v7380 = ~(w15826 | w15897);
assign w15902 = v7380;
assign v7381 = ~(w15847 | w15893);
assign w15903 = v7381;
assign v7382 = ~(w15839 | w15843);
assign w15904 = v7382;
assign w15905 = w15864 & ~w15866;
assign v7383 = ~(w15868 | w15905);
assign w15906 = v7383;
assign w15907 = w15878 & ~w15880;
assign v7384 = ~(w15882 | w15907);
assign w15908 = v7384;
assign v7385 = ~(w15906 | w15908);
assign w15909 = v7385;
assign w15910 = w15906 & w15908;
assign v7386 = ~(w15909 | w15910);
assign w15911 = v7386;
assign w15912 = pi49 & pi61;
assign w15913 = pi51 & pi59;
assign v7387 = ~(w15867 | w15913);
assign w15914 = v7387;
assign w15915 = pi51 & pi60;
assign w15916 = w15790 & w15915;
assign v7388 = ~(w15914 | w15916);
assign w15917 = v7388;
assign w15918 = w15912 & ~w15917;
assign w15919 = ~w15912 & w15917;
assign v7389 = ~(w15918 | w15919);
assign w15920 = v7389;
assign w15921 = ~w15911 & w15920;
assign w15922 = w15911 & ~w15920;
assign v7390 = ~(w15921 | w15922);
assign w15923 = v7390;
assign v7391 = ~(w15875 | w15887);
assign w15924 = v7391;
assign w15925 = w15923 & ~w15924;
assign w15926 = ~w15923 & w15924;
assign v7392 = ~(w15925 | w15926);
assign w15927 = v7392;
assign w15928 = w15904 & ~w15927;
assign w15929 = ~w15904 & w15927;
assign v7393 = ~(w15928 | w15929);
assign w15930 = v7393;
assign w15931 = pi47 & pi63;
assign w15932 = pi48 & pi62;
assign v7394 = ~(w15931 | w15932);
assign w15933 = v7394;
assign w15934 = pi48 & pi63;
assign w15935 = w15777 & w15934;
assign v7395 = ~(w15933 | w15935);
assign w15936 = v7395;
assign v7396 = ~(pi54 | w15777);
assign w15937 = v7396;
assign w15938 = pi55 & ~w15937;
assign w15939 = w15936 & w15938;
assign v7397 = ~(w15936 | w15938);
assign w15940 = v7397;
assign v7398 = ~(w15939 | w15940);
assign w15941 = v7398;
assign w15942 = pi52 & pi58;
assign w15943 = pi54 & pi56;
assign v7399 = ~(w15881 | w15943);
assign w15944 = v7399;
assign w15945 = pi54 & pi57;
assign w15946 = w15808 & w15945;
assign v7400 = ~(w15944 | w15946);
assign w15947 = v7400;
assign w15948 = w15942 & ~w15947;
assign w15949 = ~w15942 & w15947;
assign v7401 = ~(w15948 | w15949);
assign w15950 = v7401;
assign w15951 = ~w15941 & w15950;
assign w15952 = w15941 & ~w15950;
assign v7402 = ~(w15951 | w15952);
assign w15953 = v7402;
assign v7403 = ~(w15852 | w15858);
assign w15954 = v7403;
assign w15955 = ~w15953 & w15954;
assign w15956 = w15953 & ~w15954;
assign v7404 = ~(w15955 | w15956);
assign w15957 = v7404;
assign v7405 = ~(w15862 | w15890);
assign w15958 = v7405;
assign w15959 = w15957 & ~w15958;
assign w15960 = ~w15957 & w15958;
assign v7406 = ~(w15959 | w15960);
assign w15961 = v7406;
assign w15962 = w15930 & w15961;
assign v7407 = ~(w15930 | w15961);
assign w15963 = v7407;
assign v7408 = ~(w15962 | w15963);
assign w15964 = v7408;
assign w15965 = ~w15903 & w15964;
assign w15966 = w15903 & ~w15964;
assign v7409 = ~(w15965 | w15966);
assign w15967 = v7409;
assign w15968 = (w13978 & w17395) | (w13978 & w17396) | (w17395 & w17396);
assign w15969 = (~w13978 & w17397) | (~w13978 & w17398) | (w17397 & w17398);
assign v7410 = ~(w15968 | w15969);
assign w15970 = v7410;
assign v7411 = ~(w15896 | w15965);
assign w15971 = v7411;
assign v7412 = ~(w15959 | w15962);
assign w15972 = v7412;
assign v7413 = ~(w15935 | w15939);
assign w15973 = v7413;
assign w15974 = w15912 & ~w15914;
assign v7414 = ~(w15916 | w15974);
assign w15975 = v7414;
assign w15976 = w15942 & ~w15944;
assign v7415 = ~(w15946 | w15976);
assign w15977 = v7415;
assign v7416 = ~(w15975 | w15977);
assign w15978 = v7416;
assign w15979 = w15975 & w15977;
assign v7417 = ~(w15978 | w15979);
assign w15980 = v7417;
assign w15981 = w15973 & ~w15980;
assign w15982 = ~w15973 & w15980;
assign v7418 = ~(w15981 | w15982);
assign w15983 = v7418;
assign v7419 = ~(w15909 | w15922);
assign w15984 = v7419;
assign w15985 = ~w15983 & w15984;
assign w15986 = w15983 & ~w15984;
assign v7420 = ~(w15985 | w15986);
assign w15987 = v7420;
assign v7421 = ~(w15952 | w15956);
assign w15988 = v7421;
assign w15989 = ~w15987 & w15988;
assign w15990 = w15987 & ~w15988;
assign v7422 = ~(w15989 | w15990);
assign w15991 = v7422;
assign v7423 = ~(w15925 | w15929);
assign w15992 = v7423;
assign w15993 = pi50 & pi61;
assign v7424 = ~(w15915 | w15993);
assign w15994 = v7424;
assign w15995 = pi51 & pi61;
assign w15996 = w15867 & w15995;
assign v7425 = ~(w15994 | w15996);
assign w15997 = v7425;
assign w15998 = w15934 & ~w15997;
assign w15999 = ~w15934 & w15997;
assign v7426 = ~(w15998 | w15999);
assign w16000 = v7426;
assign w16001 = pi49 & pi62;
assign w16002 = ~pi55 & pi56;
assign w16003 = w16001 & ~w16002;
assign w16004 = ~w16001 & w16002;
assign v7427 = ~(w16003 | w16004);
assign w16005 = v7427;
assign v7428 = ~(w16000 | w16005);
assign w16006 = v7428;
assign w16007 = w16000 & w16005;
assign v7429 = ~(w16006 | w16007);
assign w16008 = v7429;
assign w16009 = pi52 & pi59;
assign w16010 = pi53 & pi58;
assign v7430 = ~(w15945 | w16010);
assign w16011 = v7430;
assign w16012 = pi54 & pi58;
assign w16013 = w15881 & w16012;
assign v7431 = ~(w16011 | w16013);
assign w16014 = v7431;
assign w16015 = w16009 & ~w16014;
assign w16016 = ~w16009 & w16014;
assign v7432 = ~(w16015 | w16016);
assign w16017 = v7432;
assign w16018 = w16008 & ~w16017;
assign w16019 = ~w16008 & w16017;
assign v7433 = ~(w16018 | w16019);
assign w16020 = v7433;
assign w16021 = ~w15992 & w16020;
assign w16022 = w15992 & ~w16020;
assign v7434 = ~(w16021 | w16022);
assign w16023 = v7434;
assign w16024 = w15991 & w16023;
assign v7435 = ~(w15991 | w16023);
assign w16025 = v7435;
assign v7436 = ~(w16024 | w16025);
assign w16026 = v7436;
assign w16027 = ~w15972 & w16026;
assign w16028 = w15972 & ~w16026;
assign v7437 = ~(w16027 | w16028);
assign w16029 = v7437;
assign w16030 = (~w11122 & w17664) | (~w11122 & w17665) | (w17664 & w17665);
assign w16031 = (w11122 & w17666) | (w11122 & w17667) | (w17666 & w17667);
assign v7438 = ~(w16030 | w16031);
assign w16032 = v7438;
assign v7439 = ~(w16021 | w16024);
assign w16033 = v7439;
assign v7440 = ~(w15986 | w15990);
assign w16034 = v7440;
assign w16035 = pi49 & pi63;
assign w16036 = pi52 & pi60;
assign v7441 = ~(w15995 | w16036);
assign w16037 = v7441;
assign w16038 = pi52 & pi61;
assign w16039 = w15915 & w16038;
assign v7442 = ~(w16037 | w16039);
assign w16040 = v7442;
assign w16041 = w16035 & ~w16040;
assign w16042 = ~w16035 & w16040;
assign v7443 = ~(w16041 | w16042);
assign w16043 = v7443;
assign w16044 = w15934 & ~w15994;
assign v7444 = ~(w15996 | w16044);
assign w16045 = v7444;
assign v7445 = ~(w16043 | w16045);
assign w16046 = v7445;
assign w16047 = w16043 & w16045;
assign v7446 = ~(w16046 | w16047);
assign w16048 = v7446;
assign w16049 = pi53 & pi59;
assign w16050 = pi55 & pi57;
assign v7447 = ~(w16012 | w16050);
assign w16051 = v7447;
assign w16052 = pi55 & pi58;
assign w16053 = w15945 & w16052;
assign v7448 = ~(w16051 | w16053);
assign w16054 = v7448;
assign w16055 = w16049 & ~w16054;
assign w16056 = ~w16049 & w16054;
assign v7449 = ~(w16055 | w16056);
assign w16057 = v7449;
assign w16058 = w16048 & ~w16057;
assign w16059 = ~w16048 & w16057;
assign v7450 = ~(w16058 | w16059);
assign w16060 = v7450;
assign w16061 = ~w16034 & w16060;
assign w16062 = w16034 & ~w16060;
assign v7451 = ~(w16061 | w16062);
assign w16063 = v7451;
assign w16064 = pi50 & pi62;
assign v7452 = ~(pi55 | w16001);
assign w16065 = v7452;
assign w16066 = pi56 & ~w16065;
assign w16067 = w16064 & w16066;
assign v7453 = ~(w16064 | w16066);
assign w16068 = v7453;
assign v7454 = ~(w16067 | w16068);
assign w16069 = v7454;
assign w16070 = w16009 & ~w16011;
assign v7455 = ~(w16013 | w16070);
assign w16071 = v7455;
assign w16072 = w16069 & ~w16071;
assign w16073 = ~w16069 & w16071;
assign v7456 = ~(w16072 | w16073);
assign w16074 = v7456;
assign v7457 = ~(w15978 | w15982);
assign w16075 = v7457;
assign v7458 = ~(w16006 | w16018);
assign w16076 = v7458;
assign v7459 = ~(w16075 | w16076);
assign w16077 = v7459;
assign w16078 = w16075 & w16076;
assign v7460 = ~(w16077 | w16078);
assign w16079 = v7460;
assign w16080 = w16074 & w16079;
assign v7461 = ~(w16074 | w16079);
assign w16081 = v7461;
assign v7462 = ~(w16080 | w16081);
assign w16082 = v7462;
assign w16083 = w16063 & w16082;
assign v7463 = ~(w16063 | w16082);
assign w16084 = v7463;
assign v7464 = ~(w16083 | w16084);
assign w16085 = v7464;
assign w16086 = ~w16033 & w16085;
assign w16087 = w16033 & ~w16085;
assign v7465 = ~(w16028 | w16087);
assign w16088 = v7465;
assign w16089 = (w11122 & w17668) | (w11122 & w17669) | (w17668 & w17669);
assign v7466 = ~(w16086 | w16087);
assign w16090 = v7466;
assign v7467 = ~(w16027 | w16090);
assign w16091 = v7467;
assign w16092 = (w13978 & w17401) | (w13978 & w17402) | (w17401 & w17402);
assign v7468 = ~(w16089 | w16092);
assign w16093 = v7468;
assign v7469 = ~(w16061 | w16083);
assign w16094 = v7469;
assign v7470 = ~(w16046 | w16058);
assign w16095 = v7470;
assign w16096 = pi53 & pi60;
assign v7471 = ~(w16038 | w16096);
assign w16097 = v7471;
assign w16098 = pi53 & pi61;
assign w16099 = w16036 & w16098;
assign v7472 = ~(w16097 | w16099);
assign w16100 = v7472;
assign w16101 = w16049 & ~w16051;
assign v7473 = ~(w16053 | w16101);
assign w16102 = v7473;
assign w16103 = w16100 & ~w16102;
assign w16104 = ~w16100 & w16102;
assign v7474 = ~(w16103 | w16104);
assign w16105 = v7474;
assign v7475 = ~(w16067 | w16072);
assign w16106 = v7475;
assign w16107 = w16105 & ~w16106;
assign w16108 = ~w16105 & w16106;
assign v7476 = ~(w16107 | w16108);
assign w16109 = v7476;
assign w16110 = w16095 & ~w16109;
assign w16111 = ~w16095 & w16109;
assign v7477 = ~(w16110 | w16111);
assign w16112 = v7477;
assign v7478 = ~(w16077 | w16080);
assign w16113 = v7478;
assign w16114 = pi50 & pi63;
assign w16115 = pi54 & pi59;
assign v7479 = ~(w16052 | w16115);
assign w16116 = v7479;
assign w16117 = pi55 & pi59;
assign w16118 = w16012 & w16117;
assign v7480 = ~(w16116 | w16118);
assign w16119 = v7480;
assign w16120 = w16114 & ~w16119;
assign w16121 = ~w16114 & w16119;
assign v7481 = ~(w16120 | w16121);
assign w16122 = v7481;
assign w16123 = w16035 & ~w16037;
assign v7482 = ~(w16039 | w16123);
assign w16124 = v7482;
assign v7483 = ~(w16122 | w16124);
assign w16125 = v7483;
assign w16126 = w16122 & w16124;
assign v7484 = ~(w16125 | w16126);
assign w16127 = v7484;
assign w16128 = pi51 & pi62;
assign w16129 = ~pi56 & pi57;
assign w16130 = w16128 & ~w16129;
assign w16131 = ~w16128 & w16129;
assign v7485 = ~(w16130 | w16131);
assign w16132 = v7485;
assign w16133 = w16127 & ~w16132;
assign w16134 = ~w16127 & w16132;
assign v7486 = ~(w16133 | w16134);
assign w16135 = v7486;
assign w16136 = ~w16113 & w16135;
assign w16137 = w16113 & ~w16135;
assign v7487 = ~(w16136 | w16137);
assign w16138 = v7487;
assign v7488 = ~(w16112 | w16138);
assign w16139 = v7488;
assign w16140 = w16112 & w16138;
assign v7489 = ~(w16139 | w16140);
assign w16141 = v7489;
assign w16142 = w16094 & ~w16141;
assign w16143 = ~w16094 & w16141;
assign v7490 = ~(w16142 | w16143);
assign w16144 = v7490;
assign w16145 = (w13978 & w17403) | (w13978 & w17404) | (w17403 & w17404);
assign w16146 = (~w13978 & w17405) | (~w13978 & w17406) | (w17405 & w17406);
assign v7491 = ~(w16145 | w16146);
assign w16147 = v7491;
assign v7492 = ~(w16086 | w16143);
assign w16148 = v7492;
assign v7493 = ~(w16136 | w16140);
assign w16149 = v7493;
assign v7494 = ~(w16099 | w16103);
assign w16150 = v7494;
assign v7495 = ~(pi56 | w16128);
assign w16151 = v7495;
assign w16152 = pi57 & ~w16151;
assign w16153 = w16114 & ~w16116;
assign v7496 = ~(w16118 | w16153);
assign w16154 = v7496;
assign w16155 = w16152 & ~w16154;
assign w16156 = ~w16152 & w16154;
assign v7497 = ~(w16155 | w16156);
assign w16157 = v7497;
assign w16158 = w16150 & ~w16157;
assign w16159 = ~w16150 & w16157;
assign v7498 = ~(w16158 | w16159);
assign w16160 = v7498;
assign v7499 = ~(w16107 | w16111);
assign w16161 = v7499;
assign w16162 = ~w16160 & w16161;
assign w16163 = w16160 & ~w16161;
assign v7500 = ~(w16162 | w16163);
assign w16164 = v7500;
assign v7501 = ~(w16125 | w16133);
assign w16165 = v7501;
assign w16166 = pi54 & pi60;
assign w16167 = pi56 & pi58;
assign v7502 = ~(w16117 | w16167);
assign w16168 = v7502;
assign w16169 = pi56 & pi59;
assign w16170 = w16052 & w16169;
assign v7503 = ~(w16168 | w16170);
assign w16171 = v7503;
assign w16172 = w16166 & ~w16171;
assign w16173 = ~w16166 & w16171;
assign v7504 = ~(w16172 | w16173);
assign w16174 = v7504;
assign w16175 = pi51 & pi63;
assign w16176 = pi52 & pi62;
assign v7505 = ~(w16098 | w16176);
assign w16177 = v7505;
assign w16178 = pi53 & pi62;
assign w16179 = w16038 & w16178;
assign v7506 = ~(w16177 | w16179);
assign w16180 = v7506;
assign w16181 = w16175 & ~w16180;
assign w16182 = ~w16175 & w16180;
assign v7507 = ~(w16181 | w16182);
assign w16183 = v7507;
assign v7508 = ~(w16174 | w16183);
assign w16184 = v7508;
assign w16185 = w16174 & w16183;
assign v7509 = ~(w16184 | w16185);
assign w16186 = v7509;
assign w16187 = w16165 & ~w16186;
assign w16188 = ~w16165 & w16186;
assign v7510 = ~(w16187 | w16188);
assign w16189 = v7510;
assign w16190 = w16164 & w16189;
assign v7511 = ~(w16164 | w16189);
assign w16191 = v7511;
assign v7512 = ~(w16190 | w16191);
assign w16192 = v7512;
assign w16193 = w16149 & ~w16192;
assign w16194 = ~w16149 & w16192;
assign v7513 = ~(w16193 | w16194);
assign w16195 = v7513;
assign w16196 = (~w12329 & w17531) | (~w12329 & w17532) | (w17531 & w17532);
assign w16197 = (w12329 & w17533) | (w12329 & w17534) | (w17533 & w17534);
assign v7514 = ~(w16196 | w16197);
assign w16198 = v7514;
assign v7515 = ~(w16163 | w16190);
assign w16199 = v7515;
assign v7516 = ~(w16155 | w16159);
assign w16200 = v7516;
assign w16201 = pi54 & pi61;
assign w16202 = pi55 & pi60;
assign v7517 = ~(w16169 | w16202);
assign w16203 = v7517;
assign w16204 = pi56 & pi60;
assign w16205 = w16117 & w16204;
assign v7518 = ~(w16203 | w16205);
assign w16206 = v7518;
assign w16207 = w16201 & ~w16206;
assign w16208 = ~w16201 & w16206;
assign v7519 = ~(w16207 | w16208);
assign w16209 = v7519;
assign w16210 = ~pi57 & pi58;
assign w16211 = w16178 & ~w16210;
assign w16212 = ~w16178 & w16210;
assign v7520 = ~(w16211 | w16212);
assign w16213 = v7520;
assign v7521 = ~(w16209 | w16213);
assign w16214 = v7521;
assign w16215 = w16209 & w16213;
assign v7522 = ~(w16214 | w16215);
assign w16216 = v7522;
assign w16217 = w16200 & ~w16216;
assign w16218 = ~w16200 & w16216;
assign v7523 = ~(w16217 | w16218);
assign w16219 = v7523;
assign w16220 = pi52 & pi63;
assign w16221 = w16166 & ~w16168;
assign v7524 = ~(w16170 | w16221);
assign w16222 = v7524;
assign w16223 = w16220 & ~w16222;
assign w16224 = ~w16220 & w16222;
assign v7525 = ~(w16223 | w16224);
assign w16225 = v7525;
assign w16226 = w16175 & ~w16177;
assign v7526 = ~(w16179 | w16226);
assign w16227 = v7526;
assign w16228 = ~w16225 & w16227;
assign w16229 = w16225 & ~w16227;
assign v7527 = ~(w16228 | w16229);
assign w16230 = v7527;
assign v7528 = ~(w16184 | w16188);
assign w16231 = v7528;
assign w16232 = ~w16230 & w16231;
assign w16233 = w16230 & ~w16231;
assign v7529 = ~(w16232 | w16233);
assign w16234 = v7529;
assign w16235 = w16219 & w16234;
assign v7530 = ~(w16219 | w16234);
assign w16236 = v7530;
assign v7531 = ~(w16235 | w16236);
assign w16237 = v7531;
assign w16238 = ~w16199 & w16237;
assign w16239 = w16199 & ~w16237;
assign v7532 = ~(w16238 | w16239);
assign w16240 = v7532;
assign w16241 = (~w13978 & w17407) | (~w13978 & w17408) | (w17407 & w17408);
assign w16242 = (w13978 & w17409) | (w13978 & w17410) | (w17409 & w17410);
assign v7533 = ~(w16241 | w16242);
assign w16243 = v7533;
assign v7534 = ~(w16193 | w16239);
assign w16244 = v7534;
assign w16245 = pi54 & pi62;
assign w16246 = pi53 & pi63;
assign v7535 = ~(w16245 | w16246);
assign w16247 = v7535;
assign w16248 = pi54 & pi63;
assign w16249 = w16178 & w16248;
assign v7536 = ~(w16247 | w16249);
assign w16250 = v7536;
assign v7537 = ~(pi57 | w16178);
assign w16251 = v7537;
assign w16252 = pi58 & ~w16251;
assign w16253 = w16250 & w16252;
assign v7538 = ~(w16250 | w16252);
assign w16254 = v7538;
assign v7539 = ~(w16253 | w16254);
assign w16255 = v7539;
assign w16256 = pi55 & pi61;
assign w16257 = pi57 & pi59;
assign v7540 = ~(w16204 | w16257);
assign w16258 = v7540;
assign w16259 = pi57 & pi60;
assign w16260 = w16169 & w16259;
assign v7541 = ~(w16258 | w16260);
assign w16261 = v7541;
assign w16262 = w16256 & ~w16261;
assign w16263 = ~w16256 & w16261;
assign v7542 = ~(w16262 | w16263);
assign w16264 = v7542;
assign w16265 = w16201 & ~w16203;
assign v7543 = ~(w16205 | w16265);
assign w16266 = v7543;
assign v7544 = ~(w16264 | w16266);
assign w16267 = v7544;
assign w16268 = w16264 & w16266;
assign v7545 = ~(w16267 | w16268);
assign w16269 = v7545;
assign w16270 = w16255 & w16269;
assign v7546 = ~(w16255 | w16269);
assign w16271 = v7546;
assign v7547 = ~(w16270 | w16271);
assign w16272 = v7547;
assign v7548 = ~(w16214 | w16218);
assign w16273 = v7548;
assign v7549 = ~(w16223 | w16229);
assign w16274 = v7549;
assign v7550 = ~(w16273 | w16274);
assign w16275 = v7550;
assign w16276 = w16273 & w16274;
assign v7551 = ~(w16275 | w16276);
assign w16277 = v7551;
assign w16278 = w16272 & w16277;
assign v7552 = ~(w16272 | w16277);
assign w16279 = v7552;
assign v7553 = ~(w16278 | w16279);
assign w16280 = v7553;
assign v7554 = ~(w16233 | w16235);
assign w16281 = v7554;
assign w16282 = w16280 & ~w16281;
assign w16283 = ~w16280 & w16281;
assign v7555 = ~(w16282 | w16283);
assign w16284 = v7555;
assign w16285 = (w13978 & w17411) | (w13978 & w17412) | (w17411 & w17412);
assign w16286 = (~w13978 & w17413) | (~w13978 & w17414) | (w17413 & w17414);
assign v7556 = ~(w16285 | w16286);
assign w16287 = v7556;
assign v7557 = ~(w16238 | w16282);
assign w16288 = v7557;
assign v7558 = ~(w16275 | w16278);
assign w16289 = v7558;
assign v7559 = ~(w16249 | w16253);
assign w16290 = v7559;
assign w16291 = w16256 & ~w16258;
assign v7560 = ~(w16260 | w16291);
assign w16292 = v7560;
assign v7561 = ~(w16290 | w16292);
assign w16293 = v7561;
assign w16294 = w16290 & w16292;
assign v7562 = ~(w16293 | w16294);
assign w16295 = v7562;
assign w16296 = pi56 & pi61;
assign v7563 = ~(w16259 | w16296);
assign w16297 = v7563;
assign w16298 = pi57 & pi61;
assign w16299 = w16204 & w16298;
assign v7564 = ~(w16297 | w16299);
assign w16300 = v7564;
assign w16301 = w16248 & ~w16300;
assign w16302 = ~w16248 & w16300;
assign v7565 = ~(w16301 | w16302);
assign w16303 = v7565;
assign w16304 = ~w16295 & w16303;
assign w16305 = w16295 & ~w16303;
assign v7566 = ~(w16304 | w16305);
assign w16306 = v7566;
assign v7567 = ~(w16267 | w16270);
assign w16307 = v7567;
assign w16308 = pi55 & pi62;
assign w16309 = ~pi58 & pi59;
assign w16310 = w16308 & ~w16309;
assign w16311 = ~w16308 & w16309;
assign v7568 = ~(w16310 | w16311);
assign w16312 = v7568;
assign v7569 = ~(w16307 | w16312);
assign w16313 = v7569;
assign w16314 = w16307 & w16312;
assign v7570 = ~(w16313 | w16314);
assign w16315 = v7570;
assign w16316 = w16306 & w16315;
assign v7571 = ~(w16306 | w16315);
assign w16317 = v7571;
assign v7572 = ~(w16316 | w16317);
assign w16318 = v7572;
assign w16319 = w16289 & ~w16318;
assign w16320 = ~w16289 & w16318;
assign v7573 = ~(w16319 | w16320);
assign w16321 = v7573;
assign w16322 = (w11122 & w17670) | (w11122 & w17671) | (w17670 & w17671);
assign w16323 = (~w11122 & w17672) | (~w11122 & w17673) | (w17672 & w17673);
assign v7574 = ~(w16322 | w16323);
assign w16324 = v7574;
assign w16325 = pi55 & pi63;
assign v7575 = ~(pi58 | w16308);
assign w16326 = v7575;
assign w16327 = pi59 & ~w16326;
assign w16328 = w16325 & w16327;
assign v7576 = ~(w16325 | w16327);
assign w16329 = v7576;
assign v7577 = ~(w16328 | w16329);
assign w16330 = v7577;
assign w16331 = w16248 & ~w16297;
assign v7578 = ~(w16299 | w16331);
assign w16332 = v7578;
assign w16333 = ~w16330 & w16332;
assign w16334 = w16330 & ~w16332;
assign v7579 = ~(w16333 | w16334);
assign w16335 = v7579;
assign v7580 = ~(w16293 | w16305);
assign w16336 = v7580;
assign w16337 = pi56 & pi62;
assign w16338 = pi58 & pi60;
assign v7581 = ~(w16298 | w16338);
assign w16339 = v7581;
assign w16340 = pi58 & pi61;
assign w16341 = w16259 & w16340;
assign v7582 = ~(w16339 | w16341);
assign w16342 = v7582;
assign w16343 = w16337 & ~w16342;
assign w16344 = ~w16337 & w16342;
assign v7583 = ~(w16343 | w16344);
assign w16345 = v7583;
assign v7584 = ~(w16336 | w16345);
assign w16346 = v7584;
assign w16347 = w16336 & w16345;
assign v7585 = ~(w16346 | w16347);
assign w16348 = v7585;
assign v7586 = ~(w16335 | w16348);
assign w16349 = v7586;
assign w16350 = w16335 & w16348;
assign v7587 = ~(w16349 | w16350);
assign w16351 = v7587;
assign v7588 = ~(w16313 | w16316);
assign w16352 = v7588;
assign w16353 = ~w16351 & w16352;
assign w16354 = w16351 & ~w16352;
assign v7589 = ~(w16353 | w16354);
assign w16355 = v7589;
assign w16356 = (w15213 & w17325) | (w15213 & w17326) | (w17325 & w17326);
assign w16357 = (~w15213 & w17327) | (~w15213 & w17328) | (w17327 & w17328);
assign v7590 = ~(w16356 | w16357);
assign w16358 = v7590;
assign v7591 = ~(w16328 | w16334);
assign w16359 = v7591;
assign w16360 = pi56 & pi63;
assign v7592 = ~(w16340 | w16360);
assign w16361 = v7592;
assign w16362 = w16340 & w16360;
assign v7593 = ~(w16361 | w16362);
assign w16363 = v7593;
assign w16364 = w16337 & ~w16339;
assign v7594 = ~(w16341 | w16364);
assign w16365 = v7594;
assign w16366 = w16363 & ~w16365;
assign w16367 = ~w16363 & w16365;
assign v7595 = ~(w16366 | w16367);
assign w16368 = v7595;
assign w16369 = pi57 & pi62;
assign w16370 = ~pi59 & pi60;
assign w16371 = w16369 & ~w16370;
assign w16372 = ~w16369 & w16370;
assign v7596 = ~(w16371 | w16372);
assign w16373 = v7596;
assign w16374 = w16368 & ~w16373;
assign w16375 = ~w16368 & w16373;
assign v7597 = ~(w16374 | w16375);
assign w16376 = v7597;
assign w16377 = w16359 & ~w16376;
assign w16378 = ~w16359 & w16376;
assign v7598 = ~(w16377 | w16378);
assign w16379 = v7598;
assign v7599 = ~(w16346 | w16350);
assign w16380 = v7599;
assign w16381 = w16379 & ~w16380;
assign w16382 = ~w16379 & w16380;
assign v7600 = ~(w16381 | w16382);
assign w16383 = v7600;
assign v7601 = ~(w16319 | w16353);
assign w16384 = v7601;
assign w16385 = (~w15213 & w17329) | (~w15213 & w17330) | (w17329 & w17330);
assign w16386 = (w15213 & w17331) | (w15213 & w17332) | (w17331 & w17332);
assign v7602 = ~(w16385 | w16386);
assign w16387 = v7602;
assign v7603 = ~(w16354 | w16381);
assign w16388 = v7603;
assign v7604 = ~(w16374 | w16378);
assign w16389 = v7604;
assign v7605 = ~(w16362 | w16366);
assign w16390 = v7605;
assign v7606 = ~(pi59 | w16369);
assign w16391 = v7606;
assign w16392 = pi60 & ~w16391;
assign w16393 = ~w16390 & w16392;
assign w16394 = w16390 & ~w16392;
assign v7607 = ~(w16393 | w16394);
assign w16395 = v7607;
assign w16396 = pi57 & pi63;
assign w16397 = pi59 & pi61;
assign w16398 = pi58 & pi62;
assign v7608 = ~(w16397 | w16398);
assign w16399 = v7608;
assign w16400 = pi59 & pi62;
assign w16401 = w16340 & w16400;
assign v7609 = ~(w16399 | w16401);
assign w16402 = v7609;
assign w16403 = w16396 & ~w16402;
assign w16404 = ~w16396 & w16402;
assign v7610 = ~(w16403 | w16404);
assign w16405 = v7610;
assign w16406 = w16395 & ~w16405;
assign w16407 = ~w16395 & w16405;
assign v7611 = ~(w16406 | w16407);
assign w16408 = v7611;
assign w16409 = ~w16389 & w16408;
assign w16410 = w16389 & ~w16408;
assign v7612 = ~(w16409 | w16410);
assign w16411 = v7612;
assign w16412 = (~w13978 & w17416) | (~w13978 & w17417) | (w17416 & w17417);
assign w16413 = (w13978 & w17418) | (w13978 & w17419) | (w17418 & w17419);
assign v7613 = ~(w16412 | w16413);
assign w16414 = v7613;
assign w16415 = pi58 & pi63;
assign w16416 = w16396 & ~w16399;
assign v7614 = ~(w16401 | w16416);
assign w16417 = v7614;
assign w16418 = ~w16415 & w16417;
assign w16419 = w16415 & ~w16417;
assign v7615 = ~(w16418 | w16419);
assign w16420 = v7615;
assign w16421 = ~pi60 & pi61;
assign w16422 = w16400 & ~w16421;
assign w16423 = ~w16400 & w16421;
assign v7616 = ~(w16422 | w16423);
assign w16424 = v7616;
assign w16425 = ~w16420 & w16424;
assign w16426 = w16420 & ~w16424;
assign v7617 = ~(w16425 | w16426);
assign w16427 = v7617;
assign v7618 = ~(w16393 | w16406);
assign w16428 = v7618;
assign w16429 = ~w16427 & w16428;
assign w16430 = w16427 & ~w16428;
assign v7619 = ~(w16429 | w16430);
assign w16431 = v7619;
assign w16432 = (w15213 & w17333) | (w15213 & w17334) | (w17333 & w17334);
assign w16433 = (~w15213 & w17335) | (~w15213 & w17336) | (w17335 & w17336);
assign v7620 = ~(w16432 | w16433);
assign w16434 = v7620;
assign v7621 = ~(w16410 | w16429);
assign w16435 = v7621;
assign v7622 = ~(w16419 | w16426);
assign w16436 = v7622;
assign w16437 = pi59 & pi63;
assign w16438 = pi60 & pi62;
assign v7623 = ~(w16437 | w16438);
assign w16439 = v7623;
assign w16440 = pi60 & pi63;
assign w16441 = w16400 & w16440;
assign v7624 = ~(w16439 | w16441);
assign w16442 = v7624;
assign v7625 = ~(pi60 | w16400);
assign w16443 = v7625;
assign w16444 = pi61 & ~w16443;
assign w16445 = w16442 & w16444;
assign v7626 = ~(w16442 | w16444);
assign w16446 = v7626;
assign v7627 = ~(w16445 | w16446);
assign w16447 = v7627;
assign w16448 = w16436 & ~w16447;
assign w16449 = ~w16436 & w16447;
assign v7628 = ~(w16448 | w16449);
assign w16450 = v7628;
assign w16451 = (w10008 & w17869) | (w10008 & w17870) | (w17869 & w17870);
assign w16452 = (~w10008 & w17871) | (~w10008 & w17872) | (w17871 & w17872);
assign v7629 = ~(w16451 | w16452);
assign w16453 = v7629;
assign v7630 = ~(w16430 | w16449);
assign w16454 = v7630;
assign v7631 = ~(w16441 | w16445);
assign w16455 = v7631;
assign w16456 = ~pi61 & pi62;
assign w16457 = ~w16440 & w16456;
assign w16458 = w16440 & ~w16456;
assign v7632 = ~(w16457 | w16458);
assign w16459 = v7632;
assign w16460 = w16455 & w16459;
assign v7633 = ~(w16455 | w16459);
assign w16461 = v7633;
assign v7634 = ~(w16460 | w16461);
assign w16462 = v7634;
assign w16463 = (~w10008 & w17873) | (~w10008 & w17874) | (w17873 & w17874);
assign w16464 = (w10008 & w17875) | (w10008 & w17876) | (w17875 & w17876);
assign v7635 = ~(w16463 | w16464);
assign w16465 = v7635;
assign w16466 = pi61 & pi63;
assign w16467 = pi62 & w16466;
assign w16468 = pi62 & w16459;
assign v7636 = ~(w16466 | w16468);
assign w16469 = v7636;
assign v7637 = ~(w16467 | w16469);
assign w16470 = v7637;
assign w16471 = (~w10008 & w17877) | (~w10008 & w17878) | (w17877 & w17878);
assign w16472 = (w10008 & w17879) | (w10008 & w17880) | (w17879 & w17880);
assign v7638 = ~(w16471 | w16472);
assign w16473 = v7638;
assign v7639 = ~(w16460 | w16469);
assign w16474 = v7639;
assign w16475 = ~pi62 & pi63;
assign w16476 = (~w10008 & w17881) | (~w10008 & w17882) | (w17881 & w17882);
assign w16477 = pi63 & ~w16456;
assign w16478 = (w10008 & w17883) | (w10008 & w17884) | (w17883 & w17884);
assign v7640 = ~(w16476 | w16478);
assign w16479 = v7640;
assign w16480 = (w10008 & w17885) | (w10008 & w17886) | (w17885 & w17886);
assign w16481 = pi63 & ~w16480;
assign v7641 = ~(w26 | w23);
assign w16482 = v7641;
assign v7642 = ~(w2 | w6);
assign w16483 = v7642;
assign w16484 = w26 & w23;
assign w16485 = w36 & ~w50;
assign w16486 = w110 & ~w107;
assign v7643 = ~(w119 | w121);
assign w16487 = v7643;
assign v7644 = ~(w162 | w158);
assign w16488 = v7644;
assign v7645 = ~(w235 | w226);
assign w16489 = v7645;
assign w16490 = w206 & ~w196;
assign v7646 = ~(w257 | w271);
assign w16491 = v7646;
assign v7647 = ~(w392 | w387);
assign w16492 = v7647;
assign w16493 = ~w511 & w16682;
assign w16494 = w518 & ~w510;
assign v7648 = ~(w589 | w581);
assign w16495 = v7648;
assign w16496 = ~w740 & w902;
assign w16497 = (w816 & ~w898) | (w816 & w16803) | (~w898 & w16803);
assign v7649 = ~(w1093 | w1084);
assign w16498 = v7649;
assign w16499 = ~w1283 & w17337;
assign w16500 = w1505 & ~w1393;
assign w16501 = w1505 & ~w16499;
assign w16502 = w1391 & ~w1502;
assign v7650 = ~(w1863 | w1737);
assign w16503 = v7650;
assign w16504 = w1860 & w1993;
assign w16505 = w2259 & ~w1993;
assign w16506 = w2259 & ~w16504;
assign w16507 = w2122 & ~w2257;
assign w16508 = w2402 & w2257;
assign w16509 = w2402 & ~w16507;
assign w16510 = (~w2543 & w16508) | (~w2543 & w16683) | (w16508 & w16683);
assign w16511 = (~w2543 & w16509) | (~w2543 & w16683) | (w16509 & w16683);
assign w16512 = w2688 & w2997;
assign w16513 = w3160 & ~w16512;
assign v7651 = ~(w2995 | w16513);
assign w16514 = v7651;
assign w16515 = (~w2995 & ~w3160) | (~w2995 & w16684) | (~w3160 & w16684);
assign w16516 = ~w3321 & w16804;
assign v7652 = ~(w3500 | w3491);
assign w16517 = v7652;
assign w16518 = ~w3665 & w3491;
assign w16519 = (~w3665 & w3500) | (~w3665 & w16518) | (w3500 & w16518);
assign w16520 = ~w4023 & w4029;
assign v7653 = ~(w4021 | w4029);
assign w16521 = v7653;
assign v7654 = ~(w4021 | w16520);
assign w16522 = v7654;
assign v7655 = ~(w4209 | w16521);
assign w16523 = v7655;
assign w16524 = (~w4209 & w16520) | (~w4209 & w16685) | (w16520 & w16685);
assign w16525 = ~w4594 & w4600;
assign v7656 = ~(w4592 | w4600);
assign w16526 = v7656;
assign v7657 = ~(w4592 | w16525);
assign w16527 = v7657;
assign w16528 = w4793 & w5002;
assign w16529 = w5206 & ~w5002;
assign v7658 = ~(w5201 | w16529);
assign w16530 = v7658;
assign w16531 = (~w5201 & w16528) | (~w5201 & w16686) | (w16528 & w16686);
assign w16532 = w5413 & w5627;
assign w16533 = w6070 & ~w5627;
assign v7659 = ~(w5847 | w16533);
assign w16534 = v7659;
assign w16535 = (~w5847 & w16532) | (~w5847 & w16687) | (w16532 & w16687);
assign v7660 = ~(w6067 | w16534);
assign w16536 = v7660;
assign v7661 = ~(w6067 | w16535);
assign w16537 = v7661;
assign w16538 = ~w6525 & w16688;
assign v7662 = ~(w6526 | w6769);
assign w16539 = v7662;
assign v7663 = ~(w6526 | w16538);
assign w16540 = v7663;
assign v7664 = ~(w6766 | w16539);
assign w16541 = v7664;
assign v7665 = ~(w6766 | w16540);
assign w16542 = v7665;
assign w16543 = ~w7251 & w7499;
assign v7666 = ~(w7248 | w7499);
assign w16544 = v7666;
assign v7667 = ~(w7248 | w16543);
assign w16545 = v7667;
assign v7668 = ~(w7497 | w16544);
assign w16546 = v7668;
assign w16547 = (~w7497 & w16543) | (~w7497 & w16689) | (w16543 & w16689);
assign w16548 = w7753 & ~w16546;
assign w16549 = w7753 & ~w16547;
assign v7669 = ~(w8012 | w8007);
assign w16550 = v7669;
assign w16551 = ~w8270 & w8007;
assign w16552 = (~w8270 & w8012) | (~w8270 & w16551) | (w8012 & w16551);
assign w16553 = ~w8526 & w16690;
assign w16554 = w8527 & ~w16552;
assign w16555 = w8794 & ~w16553;
assign v7670 = ~(w8789 | w16555);
assign w16556 = v7670;
assign w16557 = (~w8789 & w16554) | (~w8789 & w16691) | (w16554 & w16691);
assign w16558 = w9041 & w9535;
assign w16559 = w9773 & ~w9535;
assign v7671 = ~(w9532 | w16559);
assign w16560 = v7671;
assign w16561 = (~w9532 & w16558) | (~w9532 & w16692) | (w16558 & w16692);
assign w16562 = (~w9770 & w16559) | (~w9770 & w17535) | (w16559 & w17535);
assign v7672 = ~(w9770 | w16561);
assign w16563 = v7672;
assign v7673 = ~(w10243 | w10249);
assign w16564 = v7673;
assign w16565 = (~w10243 & w10013) | (~w10243 & w16564) | (w10013 & w16564);
assign v7674 = ~(w10472 | w16564);
assign w16566 = v7674;
assign v7675 = ~(w10472 | w16565);
assign w16567 = v7675;
assign w16568 = w10911 & ~w16566;
assign w16569 = w10911 & ~w16567;
assign w16570 = (w11121 & w16567) | (w11121 & w17420) | (w16567 & w17420);
assign w16571 = (~w10908 & w16568) | (~w10908 & w17536) | (w16568 & w17536);
assign v7676 = ~(w10908 | w16570);
assign w16572 = v7676;
assign w16573 = w11118 & w11541;
assign w16574 = w11546 & ~w11541;
assign v7677 = ~(w11539 | w16574);
assign w16575 = v7677;
assign w16576 = (~w11539 & w16573) | (~w11539 & w16693) | (w16573 & w16693);
assign v7678 = ~(w11741 | w16575);
assign w16577 = v7678;
assign v7679 = ~(w11741 | w16576);
assign w16578 = v7679;
assign w16579 = w11947 & ~w16577;
assign w16580 = w11947 & ~w16578;
assign w16581 = w12140 & ~w16580;
assign w16582 = (~w12135 & w16579) | (~w12135 & w17338) | (w16579 & w17338);
assign v7680 = ~(w12135 | w16581);
assign w16583 = v7680;
assign v7681 = ~(w12324 | w16582);
assign w16584 = v7681;
assign w16585 = (~w16580 & w17421) | (~w16580 & w17422) | (w17421 & w17422);
assign w16586 = ~w12688 & w12693;
assign v7682 = ~(w12686 | w12693);
assign w16587 = v7682;
assign v7683 = ~(w12686 | w16586);
assign w16588 = v7683;
assign v7684 = ~(w12865 | w16587);
assign w16589 = v7684;
assign w16590 = (~w12865 & w16586) | (~w12865 & w16694) | (w16586 & w16694);
assign w16591 = w13041 & ~w16589;
assign w16592 = w13041 & ~w16590;
assign w16593 = w13208 & ~w16592;
assign w16594 = (~w13203 & w16591) | (~w13203 & w17273) | (w16591 & w17273);
assign v7685 = ~(w13203 | w16593);
assign w16595 = v7685;
assign v7686 = ~(w13364 | w16594);
assign w16596 = v7686;
assign w16597 = (~w16592 & w17340) | (~w16592 & w17341) | (w17340 & w17341);
assign w16598 = (w13681 & w16594) | (w13681 & w17342) | (w16594 & w17342);
assign w16599 = w13681 & ~w16597;
assign w16600 = (w16594 & w17537) | (w16594 & w17538) | (w17537 & w17538);
assign w16601 = (~w16597 & w17674) | (~w16597 & w17537) | (w17674 & w17537);
assign v7687 = ~(w13831 | w16600);
assign w16602 = v7687;
assign w16603 = (w16597 & w17675) | (w16597 & w17676) | (w17675 & w17676);
assign w16604 = ~w13982 & w14125;
assign v7688 = ~(w14120 | w14125);
assign w16605 = v7688;
assign v7689 = ~(w14120 | w16604);
assign w16606 = v7689;
assign w16607 = (~w14256 & w14125) | (~w14256 & w16695) | (w14125 & w16695);
assign w16608 = (~w14256 & w16604) | (~w14256 & w16695) | (w16604 & w16695);
assign w16609 = w14520 & ~w16607;
assign w16610 = (~w16604 & w17019) | (~w16604 & w17020) | (w17019 & w17020);
assign w16611 = w14524 & ~w16610;
assign w16612 = (~w14518 & w16609) | (~w14518 & w17275) | (w16609 & w17275);
assign v7690 = ~(w14518 | w16611);
assign w16613 = v7690;
assign v7691 = ~(w14645 | w16612);
assign w16614 = v7691;
assign w16615 = (~w16610 & w17343) | (~w16610 & w17344) | (w17343 & w17344);
assign w16616 = (w14885 & w16612) | (w14885 & w17345) | (w16612 & w17345);
assign w16617 = w14885 & ~w16615;
assign w16618 = (~w16612 & w17425) | (~w16612 & w17426) | (w17425 & w17426);
assign v7692 = ~(w14882 | w16618);
assign w16619 = v7692;
assign w16620 = (~w16615 & w17540) | (~w16615 & w17541) | (w17540 & w17541);
assign v7693 = ~(w14993 | w16619);
assign w16621 = v7693;
assign v7694 = ~(w14993 | w16620);
assign w16622 = v7694;
assign w16623 = (~w16618 & w17677) | (~w16618 & w17678) | (w17677 & w17678);
assign w16624 = (w15109 & w16620) | (w15109 & w17542) | (w16620 & w17542);
assign w16625 = w15212 & ~w16623;
assign w16626 = w15212 & ~w16624;
assign v7695 = ~(w15207 | w16625);
assign w16627 = v7695;
assign v7696 = ~(w15207 | w16626);
assign w16628 = v7696;
assign w16629 = w15311 & w15411;
assign w16630 = w15588 & ~w15411;
assign v7697 = ~(w15499 | w16630);
assign w16631 = v7697;
assign w16632 = (~w15499 & w16629) | (~w15499 & w16696) | (w16629 & w16696);
assign w16633 = (~w15586 & w16630) | (~w15586 & w16805) | (w16630 & w16805);
assign v7698 = ~(w15586 | w16632);
assign w16634 = v7698;
assign w16635 = (~w16630 & w16806) | (~w16630 & w17021) | (w16806 & w17021);
assign w16636 = (w15676 & w16632) | (w15676 & w16806) | (w16632 & w16806);
assign w16637 = (~w16632 & w17022) | (~w16632 & w17023) | (w17022 & w17023);
assign w16638 = (~w15749 & w16635) | (~w15749 & w17277) | (w16635 & w17277);
assign v7699 = ~(w15749 | w16637);
assign w16639 = v7699;
assign w16640 = (~w16635 & w17278) | (~w16635 & w17346) | (w17278 & w17346);
assign w16641 = (~w15827 & w16637) | (~w15827 & w17278) | (w16637 & w17278);
assign w16642 = w15902 & ~w16640;
assign w16643 = (~w16637 & w17347) | (~w16637 & w17348) | (w17347 & w17348);
assign w16644 = (w16637 & w17428) | (w16637 & w17429) | (w17428 & w17429);
assign w16645 = (~w16640 & w17543) | (~w16640 & w17544) | (w17543 & w17544);
assign v7700 = ~(w15966 | w16644);
assign w16646 = v7700;
assign w16647 = (w16640 & w17679) | (w16640 & w17680) | (w17679 & w17680);
assign w16648 = (w16637 & w17681) | (w16637 & w17682) | (w17681 & w17682);
assign w16649 = w16088 & ~w16647;
assign w16650 = w16088 & ~w16648;
assign w16651 = w16148 & ~w16649;
assign w16652 = w16148 & ~w16650;
assign v7701 = ~(w16142 | w16651);
assign w16653 = v7701;
assign v7702 = ~(w16142 | w16652);
assign w16654 = v7702;
assign v7703 = ~(w16194 | w16653);
assign w16655 = v7703;
assign v7704 = ~(w16194 | w16654);
assign w16656 = v7704;
assign w16657 = w16244 & ~w16655;
assign w16658 = w16244 & ~w16656;
assign w16659 = w16288 & ~w16657;
assign w16660 = w16288 & ~w16658;
assign v7705 = ~(w16283 | w16659);
assign w16661 = v7705;
assign v7706 = ~(w16283 | w16660);
assign w16662 = v7706;
assign w16663 = w16320 & w16384;
assign w16664 = w16388 & ~w16384;
assign w16665 = w16388 & ~w16663;
assign v7707 = ~(w16382 | w16664);
assign w16666 = v7707;
assign v7708 = ~(w16382 | w16665);
assign w16667 = v7708;
assign v7709 = ~(w16409 | w16666);
assign w16668 = v7709;
assign v7710 = ~(w16409 | w16667);
assign w16669 = v7710;
assign w16670 = w16435 & ~w16668;
assign w16671 = w16435 & ~w16669;
assign w16672 = w16454 & ~w16670;
assign w16673 = w16454 & ~w16671;
assign v7711 = ~(w16448 | w16672);
assign w16674 = v7711;
assign v7712 = ~(w16448 | w16673);
assign w16675 = v7712;
assign v7713 = ~(w16461 | w16674);
assign w16676 = v7713;
assign v7714 = ~(w16461 | w16675);
assign w16677 = v7714;
assign v7715 = ~(w16460 | w16676);
assign w16678 = v7715;
assign v7716 = ~(w16460 | w16677);
assign w16679 = v7716;
assign w16680 = w16474 & ~w16676;
assign w16681 = w16474 & ~w16677;
assign w16682 = ~w449 & w448;
assign v7717 = ~(w2690 | w2543);
assign w16683 = v7717;
assign w16684 = w2997 & ~w2995;
assign w16685 = w4021 & ~w4209;
assign v7718 = ~(w5206 | w5201);
assign w16686 = v7718;
assign v7719 = ~(w6070 | w5847);
assign w16687 = v7719;
assign v7720 = ~(w6295 | w6528);
assign w16688 = v7720;
assign w16689 = w7248 & ~w7497;
assign v7721 = ~(w8269 | w16551);
assign w16690 = v7721;
assign v7722 = ~(w8794 | w8789);
assign w16691 = v7722;
assign v7723 = ~(w9773 | w9532);
assign w16692 = v7723;
assign v7724 = ~(w11546 | w11539);
assign w16693 = v7724;
assign w16694 = w12686 & ~w12865;
assign w16695 = w14120 & ~w14256;
assign v7725 = ~(w15588 | w15499);
assign w16696 = v7725;
assign w16697 = w327 & ~w316;
assign v7726 = ~(w376 | w372);
assign w16698 = v7726;
assign w16699 = w395 & ~w416;
assign w16700 = w437 & ~w426;
assign w16701 = w470 & ~w459;
assign w16702 = w570 & ~w559;
assign w16703 = ~w656 & w581;
assign v7727 = ~(w656 | w16495);
assign w16704 = v7727;
assign w16705 = w645 & ~w631;
assign v7728 = ~(w802 | w798);
assign w16706 = v7728;
assign v7729 = ~(w972 | w968);
assign w16707 = v7729;
assign w16708 = w998 & ~w1017;
assign w16709 = w1045 & ~w1034;
assign v7730 = ~(w1131 | w1123);
assign w16710 = v7730;
assign w16711 = w1192 & ~w1197;
assign v7731 = ~(w1306 | w1302);
assign w16712 = v7731;
assign w16713 = w1334 & ~w1323;
assign v7732 = ~(w1404 | w1406);
assign w16714 = v7732;
assign v7733 = ~(w1444 | w1440);
assign w16715 = v7733;
assign v7734 = ~(w1687 | w1683);
assign w16716 = v7734;
assign w16717 = w2055 & ~w2044;
assign v7735 = ~(w2135 | w2131);
assign w16718 = v7735;
assign w16719 = w2190 & ~w2179;
assign v7736 = ~(w2436 | w2432);
assign w16720 = v7736;
assign v7737 = ~(w2451 | w2447);
assign w16721 = v7737;
assign v7738 = ~(w3011 | w3013);
assign w16722 = v7738;
assign w16723 = w3166 & ~w3171;
assign v7739 = ~(w3295 | w3291);
assign w16724 = v7739;
assign v7740 = ~(w3309 | w3307);
assign w16725 = v7740;
assign v7741 = ~(w3233 | w3236);
assign w16726 = v7741;
assign w16727 = w3329 & ~w3364;
assign w16728 = w3377 & w3550;
assign v7742 = ~(w3377 | w3550);
assign w16729 = v7742;
assign v7743 = ~(w3360 | w3345);
assign w16730 = v7743;
assign v7744 = ~(w3632 | w3628);
assign w16731 = v7744;
assign w16732 = w3972 & ~w3961;
assign v7745 = ~(w3858 | w3854);
assign w16733 = v7745;
assign v7746 = ~(w4413 | w4409);
assign w16734 = v7746;
assign v7747 = ~(w4765 | w4758);
assign w16735 = v7747;
assign v7748 = ~(w4697 | w4693);
assign w16736 = v7748;
assign w16737 = w4720 & ~w4709;
assign v7749 = ~(w4918 | w4914);
assign w16738 = v7749;
assign v7750 = ~(w4942 | w4938);
assign w16739 = v7750;
assign v7751 = ~(w5397 | w5393);
assign w16740 = v7751;
assign v7752 = ~(w5220 | w5214);
assign w16741 = v7752;
assign v7753 = ~(w5503 | w5499);
assign w16742 = v7753;
assign w16743 = w5787 & ~w5783;
assign v7754 = ~(w5767 | w5763);
assign w16744 = v7754;
assign v7755 = ~(w6018 | w6011);
assign w16745 = v7755;
assign v7756 = ~(w5875 | w5871);
assign w16746 = v7756;
assign v7757 = ~(w5987 | w5983);
assign w16747 = v7757;
assign v7758 = ~(w5887 | w5883);
assign w16748 = v7758;
assign v7759 = ~(w6313 | w6309);
assign w16749 = v7759;
assign w16750 = w6595 & ~w6591;
assign v7760 = ~(w6570 | w6566);
assign w16751 = v7760;
assign w16752 = w7071 & ~w7067;
assign v7761 = ~(w7059 | w7055);
assign w16753 = v7761;
assign w16754 = w7834 & ~w7822;
assign w16755 = pi63 & pi01;
assign w16756 = w8231 & ~w8227;
assign v7762 = ~(w8025 | w8021);
assign w16757 = v7762;
assign v7763 = ~(w8305 | w8303);
assign w16758 = v7763;
assign w16759 = w8890 & w9084;
assign v7764 = ~(w8890 | w9084);
assign w16760 = v7764;
assign w16761 = w9125 & ~w9114;
assign w16762 = w9080 & ~w9076;
assign v7765 = ~(w9467 | w9463);
assign w16763 = v7765;
assign w16764 = w9434 & ~w9430;
assign v7766 = ~(w9501 | w9500);
assign w16765 = v7766;
assign w16766 = w9592 & ~w9588;
assign v7767 = ~(w9553 | w9549);
assign w16767 = v7767;
assign w16768 = w9877 & ~w9866;
assign w16769 = w10144 & ~w10134;
assign w16770 = w10745 & ~w10734;
assign v7768 = ~(w10787 | w10783);
assign w16771 = v7768;
assign w16772 = w11240 & ~w11236;
assign w16773 = w11424 & ~w11420;
assign v7769 = ~(w12648 | w12647);
assign w16774 = v7769;
assign w16775 = w12603 & ~w12599;
assign v7770 = ~(w12615 | w12611);
assign w16776 = v7770;
assign v7771 = ~(w12735 | w12731);
assign w16777 = v7771;
assign v7772 = ~(w12833 | w12829);
assign w16778 = v7772;
assign w16779 = w12785 & w12919;
assign v7773 = ~(w12785 | w12919);
assign w16780 = v7773;
assign w16781 = w14625 & w14653;
assign v7774 = ~(w14625 | w14653);
assign w16782 = v7774;
assign w16783 = w14535 & ~w14531;
assign w16784 = w14699 & ~w14695;
assign w16785 = w14829 & ~w14825;
assign w16786 = w14930 & ~w14926;
assign v7775 = ~(w16320 | w16662);
assign w16787 = v7775;
assign v7776 = ~(w16320 | w16661);
assign w16788 = v7776;
assign w16789 = (w16384 & w16663) | (w16384 & w16662) | (w16663 & w16662);
assign w16790 = (w16384 & w16663) | (w16384 & w16661) | (w16663 & w16661);
assign w16791 = (w16668 & w16669) | (w16668 & ~w16662) | (w16669 & ~w16662);
assign w16792 = (w16668 & w16669) | (w16668 & ~w16661) | (w16669 & ~w16661);
assign w16793 = (w16670 & w16671) | (w16670 & w16662) | (w16671 & w16662);
assign w16794 = (w16670 & w16671) | (w16670 & w16661) | (w16671 & w16661);
assign w16795 = ~w16430 & w16450;
assign w16796 = w16430 & ~w16450;
assign w16797 = (w16674 & w16675) | (w16674 & w16662) | (w16675 & w16662);
assign w16798 = (w16674 & w16675) | (w16674 & w16661) | (w16675 & w16661);
assign w16799 = (w16678 & w16679) | (w16678 & w16662) | (w16679 & w16662);
assign w16800 = (w16678 & w16679) | (w16678 & w16661) | (w16679 & w16661);
assign w16801 = (w16680 & w16681) | (w16680 & w16662) | (w16681 & w16662);
assign w16802 = (w16680 & w16681) | (w16680 & w16661) | (w16681 & w16661);
assign w16803 = w821 & w816;
assign w16804 = ~w3158 & w3157;
assign w16805 = w15499 & ~w15586;
assign w16806 = w15586 & w15676;
assign w16807 = w294 & ~w286;
assign w16808 = w360 & ~w357;
assign v7777 = ~(w490 | w501);
assign w16809 = v7777;
assign w16810 = (w16493 & w583) | (w16493 & ~w387) | (w583 & ~w387);
assign w16811 = (w16493 & w583) | (w16493 & w16492) | (w583 & w16492);
assign v7778 = ~(w529 | w525);
assign w16812 = v7778;
assign v7779 = ~(w532 | w535);
assign w16813 = v7779;
assign v7780 = ~(w593 | w598);
assign w16814 = v7780;
assign v7781 = ~(w603 | w606);
assign w16815 = v7781;
assign w16816 = w678 & ~w667;
assign v7782 = ~(w691 | w683);
assign w16817 = v7782;
assign v7783 = ~(w681 | w695);
assign w16818 = v7783;
assign w16819 = w786 & ~w775;
assign w16820 = w888 & ~w885;
assign w16821 = (w16497 & ~w899) | (w16497 & w902) | (~w899 & w902);
assign w16822 = (w16497 & ~w899) | (w16497 & w16496) | (~w899 & w16496);
assign w16823 = w953 & ~w942;
assign w16824 = w1172 & ~w1161;
assign w16825 = ~pi13 & w1215;
assign w16826 = pi13 & ~w1215;
assign v7784 = ~(w1108 | w1111);
assign w16827 = v7784;
assign v7785 = ~(w1337 | w1341);
assign w16828 = v7785;
assign w16829 = w1377 & ~w1366;
assign w16830 = w1458 & ~w1461;
assign w16831 = w1532 & ~w1521;
assign v7786 = ~(w1550 | w1546);
assign w16832 = v7786;
assign w16833 = w1720 & ~w1709;
assign w16834 = (~w1642 & w1643) | (~w1642 & w17024) | (w1643 & w17024);
assign v7787 = ~(w1757 | w1749);
assign w16835 = v7787;
assign w16836 = w1844 & ~w1833;
assign w16837 = w1746 & ~w1761;
assign v7788 = ~(w2077 | w2073);
assign w16838 = v7788;
assign v7789 = ~(w2092 | w2088);
assign w16839 = v7789;
assign v7790 = ~(w2193 | w2159);
assign w16840 = v7790;
assign w16841 = w2197 & ~w2200;
assign w16842 = w2213 & ~w2234;
assign v7791 = ~(w2303 | w2299);
assign w16843 = v7791;
assign v7792 = ~(w2306 | w2321);
assign w16844 = v7792;
assign w16845 = w2377 & ~w2366;
assign w16846 = w2267 & ~w2278;
assign v7793 = ~(w2539 | w2424);
assign w16847 = v7793;
assign v7794 = ~(w2536 | w2461);
assign w16848 = v7794;
assign w16849 = w2530 & ~w2519;
assign v7795 = ~(w2439 | w2455);
assign w16850 = v7795;
assign v7796 = ~(w2533 | w2498);
assign w16851 = v7796;
assign w16852 = w2418 & w2677;
assign v7797 = ~(w2418 | w2677);
assign w16853 = v7797;
assign w16854 = w2551 & ~w2554;
assign v7798 = ~(w2613 | w2606);
assign w16855 = v7798;
assign v7799 = ~(w2817 | w2809);
assign w16856 = v7799;
assign v7800 = ~(w2860 | w2856);
assign w16857 = v7800;
assign w16858 = w2972 & ~w2961;
assign w16859 = w2914 & ~w2904;
assign v7801 = ~(w3063 | w3059);
assign w16860 = v7801;
assign v7802 = ~(w3033 | w3029);
assign w16861 = v7802;
assign w16862 = w3100 & ~w3089;
assign w16863 = w3141 & ~w3130;
assign w16864 = w3210 & ~w3199;
assign w16865 = w3272 & ~w3261;
assign v7803 = ~(w3357 | w3353);
assign w16866 = v7803;
assign w16867 = w3592 & ~w3614;
assign v7804 = ~(w3601 | w3594);
assign w16868 = v7804;
assign v7805 = ~(w3585 | w3551);
assign w16869 = v7805;
assign w16870 = w3778 & ~w3789;
assign w16871 = w3748 & ~w3772;
assign w16872 = w3761 & ~w3766;
assign w16873 = w3944 & ~w3933;
assign w16874 = w3910 & ~w3899;
assign w16875 = w4032 & ~w4035;
assign w16876 = w4307 & ~w4296;
assign v7806 = ~(w4379 | w4375);
assign w16877 = v7806;
assign w16878 = w4334 & ~w4322;
assign w16879 = w4569 & ~w4558;
assign w16880 = w4518 & ~w4507;
assign w16881 = w4673 & ~w4662;
assign w16882 = w4755 & ~w4769;
assign w16883 = w4637 & ~w4625;
assign w16884 = w4955 & ~w4947;
assign w16885 = w4832 & ~w4821;
assign w16886 = w4858 & ~w4847;
assign w16887 = w4894 & ~w4883;
assign w16888 = w4969 & ~w4972;
assign v7807 = ~(w5124 | w5127);
assign w16889 = v7807;
assign w16890 = w5009 & ~w5027;
assign w16891 = w5421 & ~w5432;
assign w16892 = w5602 & ~w5591;
assign w16893 = w5483 & ~w5473;
assign v7808 = ~(w5453 | w5449);
assign w16894 = v7808;
assign w16895 = w5820 & ~w5823;
assign w16896 = w5740 & ~w5729;
assign w16897 = w5668 & ~w5657;
assign w16898 = w5854 & ~w5857;
assign w16899 = w6199 & ~w6187;
assign v7809 = ~(w6125 | w6128);
assign w16900 = v7809;
assign w16901 = w6091 & ~w6080;
assign w16902 = w6122 & ~w6119;
assign w16903 = w6364 & ~w6353;
assign w16904 = w6459 & ~w6457;
assign w16905 = w6675 & ~w6663;
assign w16906 = w6727 & ~w6740;
assign w16907 = w6911 & ~w6900;
assign w16908 = w6984 & ~w6973;
assign w16909 = w6778 & ~w6781;
assign w16910 = w7160 & ~w7149;
assign w16911 = w7261 & ~w7264;
assign w16912 = w7572 & ~w7562;
assign w16913 = w7774 & ~w7763;
assign v7810 = ~(w7952 | w7948);
assign w16914 = v7810;
assign w16915 = w7940 & ~w7936;
assign w16916 = w8033 & ~w8031;
assign v7811 = ~(w8234 | w8249);
assign w16917 = v7811;
assign w16918 = w8447 & ~w8450;
assign w16919 = w8376 & ~w8365;
assign w16920 = w8633 & ~w8623;
assign w16921 = w8659 & ~w8647;
assign w16922 = w9242 & ~w9231;
assign v7812 = ~(w9090 | w9086);
assign w16923 = v7812;
assign w16924 = w9367 & ~w9357;
assign w16925 = w9402 & ~w9391;
assign w16926 = w9335 & ~w9323;
assign w16927 = w9485 & ~w9488;
assign w16928 = w9656 & ~w9646;
assign w16929 = w9685 & ~w9673;
assign v7813 = ~(w9556 | w9559);
assign w16930 = v7813;
assign w16931 = w9858 & ~w9848;
assign v7814 = ~(w9977 | w9980);
assign w16932 = v7814;
assign w16933 = w10188 & ~w10177;
assign w16934 = w10017 & ~w10021;
assign w16935 = w10253 & ~w10264;
assign w16936 = w10889 & ~w10878;
assign w16937 = w10856 & ~w10845;
assign w16938 = w11050 & ~w11039;
assign w16939 = w11014 & ~w11008;
assign w16940 = w10917 & ~w10920;
assign w16941 = w11317 & ~w11305;
assign w16942 = w11522 & ~w11511;
assign w16943 = w11492 & ~w11485;
assign v7815 = ~(w11400 | w11399);
assign w16944 = v7815;
assign w16945 = w11394 & ~w11406;
assign w16946 = w11709 & ~w11714;
assign w16947 = w11667 & ~w11663;
assign w16948 = w11655 & ~w11651;
assign v7816 = ~(w11789 | w11764);
assign w16949 = v7816;
assign w16950 = w12579 & ~w12568;
assign w16951 = w12543 & ~w12532;
assign w16952 = w12712 & ~w12700;
assign w16953 = w12809 & ~w12798;
assign w16954 = w12777 & ~w12766;
assign v7817 = ~(w12738 | w12741);
assign w16955 = v7817;
assign v7818 = ~(w12925 | w12921);
assign w16956 = v7818;
assign w16957 = pi42 & pi43;
assign w16958 = w12987 & ~w12976;
assign w16959 = w12873 & ~w12876;
assign w16960 = w13107 & ~w13098;
assign v7819 = ~(w13052 | w13050);
assign w16961 = v7819;
assign w16962 = w13308 & ~w13298;
assign w16963 = w14748 & ~w14737;
assign w16964 = w14659 & ~w14655;
assign w16965 = pi48 & pi49;
assign w16966 = w14797 & ~w14785;
assign v7820 = ~(w14843 | w14841);
assign w16967 = v7820;
assign v7821 = ~(w14846 | w14864);
assign w16968 = v7821;
assign v7822 = ~(w14869 | w14835);
assign w16969 = v7822;
assign w16970 = w14812 & ~w14815;
assign w16971 = w14891 & ~w14897;
assign w16972 = w15001 & ~w15012;
assign v7823 = ~(w15311 | w16628);
assign w16973 = v7823;
assign v7824 = ~(w15311 | w16627);
assign w16974 = v7824;
assign w16975 = (w15411 & w16629) | (w15411 & w16628) | (w16629 & w16628);
assign w16976 = (w15411 & w16629) | (w15411 & w16627) | (w16629 & w16627);
assign w16977 = (w16633 & w16634) | (w16633 & ~w16628) | (w16634 & ~w16628);
assign w16978 = (w16633 & w16634) | (w16633 & ~w16627) | (w16634 & ~w16627);
assign w16979 = (w16636 & w16635) | (w16636 & w16628) | (w16635 & w16628);
assign w16980 = (w16636 & w16635) | (w16636 & w16627) | (w16635 & w16627);
assign w16981 = (w16641 & w16640) | (w16641 & ~w16628) | (w16640 & ~w16628);
assign w16982 = (w16641 & w16640) | (w16641 & ~w16627) | (w16640 & ~w16627);
assign w16983 = (w16643 & w16642) | (w16643 & w16628) | (w16642 & w16628);
assign w16984 = (w16643 & w16642) | (w16643 & w16627) | (w16642 & w16627);
assign w16985 = (w16646 & w16645) | (w16646 & w16628) | (w16645 & w16628);
assign w16986 = (w16646 & w16645) | (w16646 & w16627) | (w16645 & w16627);
assign w16987 = (w16650 & w16649) | (w16650 & w16628) | (w16649 & w16628);
assign w16988 = (w16650 & w16649) | (w16650 & w16627) | (w16649 & w16627);
assign w16989 = (w16656 & w16655) | (w16656 & ~w16628) | (w16655 & ~w16628);
assign w16990 = (w16656 & w16655) | (w16656 & ~w16627) | (w16655 & ~w16627);
assign w16991 = (w16658 & w16657) | (w16658 & w16628) | (w16657 & w16628);
assign w16992 = (w16658 & w16657) | (w16658 & w16627) | (w16657 & w16627);
assign w16993 = (w16662 & w16661) | (w16662 & w16628) | (w16661 & w16628);
assign w16994 = (w16662 & w16661) | (w16662 & w16627) | (w16661 & w16627);
assign v7825 = ~(w16319 | w16788);
assign w16995 = v7825;
assign v7826 = ~(w16319 | w16787);
assign w16996 = v7826;
assign v7827 = ~(w16354 | w16790);
assign w16997 = v7827;
assign v7828 = ~(w16354 | w16789);
assign w16998 = v7828;
assign v7829 = ~(w16410 | w16792);
assign w16999 = v7829;
assign v7830 = ~(w16410 | w16791);
assign w17000 = v7830;
assign w17001 = w16795 & ~w16794;
assign w17002 = w16795 & ~w16793;
assign w17003 = (~w16450 & w16796) | (~w16450 & w16794) | (w16796 & w16794);
assign w17004 = (~w16450 & w16796) | (~w16450 & w16793) | (w16796 & w16793);
assign w17005 = ~w16462 & w16798;
assign w17006 = ~w16462 & w16797;
assign w17007 = w16462 & ~w16798;
assign w17008 = w16462 & ~w16797;
assign w17009 = ~w16470 & w16800;
assign w17010 = ~w16470 & w16799;
assign w17011 = w16470 & ~w16800;
assign w17012 = w16470 & ~w16799;
assign w17013 = ~w16475 & w16802;
assign w17014 = ~w16475 & w16801;
assign w17015 = w16477 & ~w16802;
assign w17016 = w16477 & ~w16801;
assign v7831 = ~(pi62 | w16802);
assign w17017 = v7831;
assign v7832 = ~(pi62 | w16801);
assign w17018 = v7832;
assign w17019 = w14520 & w14256;
assign w17020 = w14520 & ~w16695;
assign w17021 = w15676 & ~w16805;
assign w17022 = w15755 & ~w15676;
assign w17023 = w15755 & ~w16806;
assign w17024 = w1644 & ~w1642;
assign v7833 = ~(w611 | w649);
assign w17025 = v7833;
assign v7834 = ~(w700 | w728);
assign w17026 = v7834;
assign v7835 = ~(w755 | w833);
assign w17027 = v7835;
assign w17028 = w755 & w833;
assign v7836 = ~(w789 | w806);
assign w17029 = v7836;
assign v7837 = ~(w881 | w875);
assign w17030 = v7837;
assign v7838 = ~(w830 | w826);
assign w17031 = v7838;
assign w17032 = (~w956 & w920) | (~w956 & w17279) | (w920 & w17279);
assign w17033 = w909 & ~w914;
assign v7839 = ~(w1069 | w1072);
assign w17034 = v7839;
assign v7840 = ~(w1066 | w1062);
assign w17035 = v7840;
assign w17036 = w1121 & ~w1144;
assign w17037 = w1120 & ~w1176;
assign v7841 = ~(w1105 | w1101);
assign w17038 = v7841;
assign v7842 = ~(w1239 | w1274);
assign w17039 = v7842;
assign w17040 = w1207 & ~w1205;
assign w17041 = (~w1435 & w1448) | (~w1435 & w17280) | (w1448 & w17280);
assign w17042 = (~w1502 & w16502) | (~w1502 & w16501) | (w16502 & w16501);
assign w17043 = (~w1502 & w16502) | (~w1502 & w16500) | (w16502 & w16500);
assign w17044 = (~w1605 & w1577) | (~w1605 & w17281) | (w1577 & w17281);
assign v7843 = ~(w1573 | w1569);
assign w17045 = v7843;
assign w17046 = w1639 & ~w1628;
assign w17047 = w1660 & ~w1671;
assign v7844 = ~(w1782 | w1803);
assign w17048 = v7844;
assign v7845 = ~(w1850 | w1848);
assign w17049 = v7845;
assign w17050 = w1892 & ~w1881;
assign v7846 = ~(w2061 | w2060);
assign w17051 = v7846;
assign w17052 = w2102 & ~w2105;
assign v7847 = ~(w2098 | w2096);
assign w17053 = v7847;
assign v7848 = ~(w2101 | w2113);
assign w17054 = v7848;
assign v7849 = ~(w2117 | w2065);
assign w17055 = v7849;
assign v7850 = ~(w2196 | w2208);
assign w17056 = v7850;
assign w17057 = w2154 & ~w2143;
assign w17058 = w2340 & ~w2331;
assign v7851 = ~(w2317 | w2313);
assign w17059 = v7851;
assign v7852 = ~(w2380 | w2345);
assign w17060 = v7852;
assign v7853 = ~(w2283 | w2286);
assign w17061 = v7853;
assign w17062 = w2407 & ~w2410;
assign w17063 = w2494 & ~w2483;
assign w17064 = w2667 & ~w2663;
assign w17065 = w2562 & w2797;
assign v7854 = ~(w2562 | w2797);
assign w17066 = v7854;
assign v7855 = ~(w2646 | w2678);
assign w17067 = v7855;
assign v7856 = ~(w2655 | w2651);
assign w17068 = v7856;
assign w17069 = w2775 & ~w2764;
assign w17070 = w2754 & ~w2743;
assign v7857 = ~(w2787 | w2783);
assign w17071 = v7857;
assign v7858 = ~(w2757 | w2723);
assign w17072 = v7858;
assign w17073 = w2875 & ~w2886;
assign w17074 = w3006 & ~w3019;
assign v7859 = ~(w3036 | w3039);
assign w17075 = v7859;
assign v7860 = ~(w3298 | w3301);
assign w17076 = v7860;
assign v7861 = ~(w3230 | w3226);
assign w17077 = v7861;
assign w17078 = w3405 & ~w3394;
assign v7862 = ~(w3478 | w3444);
assign w17079 = v7862;
assign w17080 = w3417 & ~w3436;
assign w17081 = w3648 & ~w3644;
assign v7863 = ~(w3654 | w3622);
assign w17082 = v7863;
assign w17083 = w3547 & ~w3536;
assign w17084 = w3806 & ~w3828;
assign v7864 = ~(w3818 | w3810);
assign w17085 = v7864;
assign v7865 = ~(w3987 | w3983);
assign w17086 = v7865;
assign v7866 = ~(w3997 | w4008);
assign w17087 = v7866;
assign v7867 = ~(w4053 | w4049);
assign w17088 = v7867;
assign v7868 = ~(w4064 | w4043);
assign w17089 = v7868;
assign v7869 = ~(w4056 | w4059);
assign w17090 = v7869;
assign v7870 = ~(w4148 | w4144);
assign w17091 = v7870;
assign v7871 = ~(w4242 | w4257);
assign w17092 = v7871;
assign v7872 = ~(w4251 | w4247);
assign w17093 = v7872;
assign v7873 = ~(w4365 | w4361);
assign w17094 = v7873;
assign w17095 = w4442 & ~w4453;
assign w17096 = w4477 & ~w4473;
assign w17097 = w4537 & ~w4526;
assign w17098 = w4421 & ~w4419;
assign v7874 = ~(w4480 | w4483);
assign w17099 = v7874;
assign w17100 = w4739 & ~w4735;
assign v7875 = ~(w4723 | w4703);
assign w17101 = v7875;
assign v7876 = ~(w4742 | w4745);
assign w17102 = v7876;
assign v7877 = ~(w4945 | w4959);
assign w17103 = v7877;
assign v7878 = ~(w5132 | w5135);
assign w17104 = v7878;
assign w17105 = w5175 & ~w5171;
assign v7879 = ~(w5121 | w5117);
assign w17106 = v7879;
assign v7880 = ~(w5155 | w5151);
assign w17107 = v7880;
assign v7881 = ~(w5158 | w5161);
assign w17108 = v7881;
assign v7882 = ~(w5381 | w5377);
assign w17109 = v7882;
assign w17110 = w5359 & ~w5347;
assign w17111 = w5212 & ~w5233;
assign v7883 = ~(w5329 | w5332);
assign w17112 = v7883;
assign v7884 = ~(w5462 | w5440);
assign w17113 = v7884;
assign v7885 = ~(w5515 | w5511);
assign w17114 = v7885;
assign v7886 = ~(w5802 | w5798);
assign w17115 = v7886;
assign v7887 = ~(w5706 | w5672);
assign w17116 = v7887;
assign v7888 = ~(w5770 | w5773);
assign w17117 = v7888;
assign v7889 = ~(w5974 | w5939);
assign w17118 = v7889;
assign w17119 = w5935 & ~w5924;
assign w17120 = w5971 & ~w5960;
assign v7890 = ~(w5990 | w5993);
assign w17121 = v7890;
assign v7891 = ~(w6153 | w6149);
assign w17122 = v7891;
assign v7892 = ~(w6237 | w6203);
assign w17123 = v7892;
assign v7893 = ~(w6103 | w6099);
assign w17124 = v7893;
assign w17125 = w6329 & ~w6325;
assign w17126 = w6486 & ~w6497;
assign w17127 = w6463 & ~w6466;
assign v7894 = ~(w6451 | w6447);
assign w17128 = v7894;
assign v7895 = ~(w6316 | w6333);
assign w17129 = v7895;
assign v7896 = ~(w6558 | w6554);
assign w17130 = v7896;
assign w17131 = w6549 & ~w6574;
assign w17132 = (~w6745 & w6746) | (~w6745 & w17683) | (w6746 & w17683);
assign v7897 = ~(w6736 | w6730);
assign w17133 = v7897;
assign w17134 = w6536 & ~w6539;
assign w17135 = (~w6914 & w6879) | (~w6914 & w17684) | (w6879 & w17684);
assign w17136 = w6868 & ~w6873;
assign w17137 = w6851 & ~w6847;
assign w17138 = w6830 & ~w6855;
assign w17139 = w6806 & ~w6821;
assign w17140 = w7041 & ~w7044;
assign w17141 = (~w7234 & w7198) | (~w7234 & w17685) | (w7198 & w17685);
assign v7898 = ~(w7297 | w7290);
assign w17142 = v7898;
assign v7899 = ~(w7437 | w7433);
assign w17143 = v7899;
assign w17144 = w7587 & ~w7592;
assign w17145 = (~w7575 & w7507) | (~w7575 & w17546) | (w7507 & w17546);
assign v7900 = ~(w7627 | w7623);
assign w17146 = v7900;
assign w17147 = w7902 & ~w7890;
assign v7901 = ~(w7943 | w7971);
assign w17148 = v7901;
assign w17149 = w7923 & ~w7926;
assign w17150 = w8210 & ~w8213;
assign w17151 = w8044 & ~w8038;
assign w17152 = w8243 & ~w8239;
assign v7902 = ~(w8455 | w8458);
assign w17153 = v7902;
assign w17154 = w8540 & ~w8565;
assign w17155 = w8768 & ~w8766;
assign v7903 = ~(w8714 | w8713);
assign w17156 = v7903;
assign w17157 = (~w8743 & w8744) | (~w8743 & w17547) | (w8744 & w17547);
assign v7904 = ~(w8983 | w8979);
assign w17158 = v7904;
assign w17159 = w9009 & ~w9005;
assign v7905 = ~(w8974 | w8989);
assign w17160 = v7905;
assign w17161 = w9017 & ~w9015;
assign w17162 = w9068 & ~w9064;
assign w17163 = w9494 & ~w9507;
assign w17164 = w9455 & ~w9451;
assign v7906 = ~(w9595 | w9610);
assign w17165 = v7906;
assign w17166 = w9604 & ~w9600;
assign w17167 = (~w9688 & w9627) | (~w9688 & w17430) | (w9627 & w17430);
assign w17168 = w9575 & ~w9578;
assign w17169 = w9788 & ~w9784;
assign w17170 = w9806 & ~w9804;
assign w17171 = (~w9861 & w9881) | (~w9861 & w17431) | (w9881 & w17431);
assign w17172 = w9974 & ~w9970;
assign w17173 = w9810 & ~w9813;
assign w17174 = w10060 & ~w10085;
assign v7907 = ~(w10081 | w10077);
assign w17175 = v7907;
assign w17176 = (~w10129 & w10148) | (~w10129 & w17432) | (w10148 & w17432);
assign w17177 = w10069 & ~w10065;
assign w17178 = w10047 & ~w10050;
assign v7908 = ~(w10197 | w10196);
assign w17179 = v7908;
assign w17180 = (~w10454 & w10417) | (~w10454 & w17433) | (w10417 & w17433);
assign v7909 = ~(w10413 | w10409);
assign w17181 = v7909;
assign w17182 = w10302 & ~w10327;
assign w17183 = w10289 & ~w10292;
assign w17184 = (~w10676 & w10641) | (~w10676 & w17434) | (w10641 & w17434);
assign w17185 = w10775 & ~w10771;
assign v7910 = ~(w10807 | w10806);
assign w17186 = v7910;
assign v7911 = ~(w10978 | w10981);
assign w17187 = v7911;
assign w17188 = w10943 & ~w10948;
assign w17189 = w10975 & ~w10971;
assign v7912 = ~(w11243 | w11246);
assign w17190 = v7912;
assign v7913 = ~(w11202 | w11198);
assign w17191 = v7913;
assign w17192 = (~w11320 & w11255) | (~w11320 & w17686) | (w11255 & w17686);
assign w17193 = w11453 & ~w11457;
assign v7914 = ~(w11436 | w11432);
assign w17194 = v7914;
assign w17195 = ~w11697 & w11797;
assign w17196 = w11697 & ~w11797;
assign v7915 = ~(w11658 | w11673);
assign w17197 = v7915;
assign w17198 = w11580 & ~w11568;
assign w17199 = w11634 & ~w11637;
assign w17200 = (~w11708 & w11720) | (~w11708 & w17687) | (w11720 & w17687);
assign w17201 = w11913 & ~w11916;
assign w17202 = w11866 & ~w11857;
assign w17203 = w11900 & ~w11889;
assign v7916 = ~(w11758 | w11754);
assign w17204 = v7916;
assign w17205 = w11815 & ~w11811;
assign w17206 = w11796 & ~w11819;
assign w17207 = w12078 & ~w12076;
assign w17208 = (~w12116 & w12117) | (~w12116 & w17688) | (w12117 & w17688);
assign v7917 = ~(w12836 | w12839);
assign w17209 = v7917;
assign w17210 = w12906 & ~w12902;
assign w17211 = w12949 & w13061;
assign v7918 = ~(w12949 | w13061);
assign w17212 = v7918;
assign v7919 = ~(w12909 | w12912);
assign w17213 = v7919;
assign w17214 = w12944 & ~w12933;
assign w17215 = w13168 & ~w13164;
assign v7920 = ~(w13180 | w13176);
assign w17216 = v7920;
assign w17217 = w13044 & ~w13056;
assign w17218 = w13150 & ~w13153;
assign v7921 = ~(w13348 | w13351);
assign w17219 = v7921;
assign w17220 = w13339 & ~w13335;
assign w17221 = w13318 & ~w13343;
assign w17222 = w13211 & ~w13214;
assign v7922 = ~(w13327 | w13323);
assign w17223 = v7922;
assign w17224 = w13399 & ~w13395;
assign w17225 = w13372 & ~w13375;
assign v7923 = ~(w13557 | w13553);
assign w17226 = v7923;
assign w17227 = w13982 & ~w16603;
assign w17228 = (w13982 & w16600) | (w13982 & w17689) | (w16600 & w17689);
assign w17229 = (w16607 & w16608) | (w16607 & w16603) | (w16608 & w16603);
assign w17230 = (~w16600 & w17690) | (~w16600 & w17691) | (w17690 & w17691);
assign w17231 = (w16610 & w16609) | (w16610 & ~w16603) | (w16609 & ~w16603);
assign w17232 = (w16600 & w17692) | (w16600 & w17693) | (w17692 & w17693);
assign w17233 = (w16615 & w16614) | (w16615 & w16603) | (w16614 & w16603);
assign w17234 = (~w16600 & w17694) | (~w16600 & w17695) | (w17694 & w17695);
assign w17235 = (w16617 & w16616) | (w16617 & ~w16603) | (w16616 & ~w16603);
assign w17236 = (w16600 & w17696) | (w16600 & w17697) | (w17696 & w17697);
assign w17237 = w14918 & ~w14906;
assign v7924 = ~(w14980 | w15017);
assign w17238 = v7924;
assign w17239 = w14980 & w15017;
assign v7925 = ~(w14921 | w14936);
assign w17240 = v7925;
assign w17241 = (w16622 & w16621) | (w16622 & w16603) | (w16621 & w16603);
assign w17242 = (~w16600 & w17698) | (~w16600 & w17699) | (w17698 & w17699);
assign w17243 = (w16624 & w16623) | (w16624 & ~w16603) | (w16623 & ~w16603);
assign w17244 = (w16600 & w17700) | (w16600 & w17701) | (w17700 & w17701);
assign w17245 = w15055 & ~w15091;
assign w17246 = (w16628 & w16627) | (w16628 & ~w16603) | (w16627 & ~w16603);
assign w17247 = (w16628 & w16627) | (w16628 & ~w16602) | (w16627 & ~w16602);
assign v7926 = ~(w15152 | w15151);
assign w17248 = v7926;
assign w17249 = w15147 & ~w15163;
assign v7927 = ~(w15168 | w15144);
assign w17250 = v7927;
assign v7928 = ~(w15310 | w16974);
assign w17251 = v7928;
assign v7929 = ~(w15310 | w16973);
assign w17252 = v7929;
assign v7930 = ~(w15405 | w16976);
assign w17253 = v7930;
assign v7931 = ~(w15405 | w16975);
assign w17254 = v7931;
assign v7932 = ~(w15585 | w16978);
assign w17255 = v7932;
assign v7933 = ~(w15585 | w16977);
assign w17256 = v7933;
assign v7934 = ~(w15670 | w16980);
assign w17257 = v7934;
assign v7935 = ~(w15670 | w16979);
assign w17258 = v7935;
assign v7936 = ~(w15826 | w16982);
assign w17259 = v7936;
assign v7937 = ~(w15826 | w16981);
assign w17260 = v7937;
assign v7938 = ~(w15896 | w16984);
assign w17261 = v7938;
assign v7939 = ~(w15896 | w16983);
assign w17262 = v7939;
assign w17263 = ~w16028 & w16986;
assign w17264 = ~w16028 & w16985;
assign v7940 = ~(w16086 | w16988);
assign w17265 = v7940;
assign v7941 = ~(w16086 | w16987);
assign w17266 = v7941;
assign v7942 = ~(w16193 | w16990);
assign w17267 = v7942;
assign v7943 = ~(w16193 | w16989);
assign w17268 = v7943;
assign v7944 = ~(w16238 | w16992);
assign w17269 = v7944;
assign v7945 = ~(w16238 | w16991);
assign w17270 = v7945;
assign w17271 = (w16666 & w16667) | (w16666 & w16994) | (w16667 & w16994);
assign w17272 = (w16666 & w16667) | (w16666 & w16993) | (w16667 & w16993);
assign v7946 = ~(w13208 | w13203);
assign w17273 = v7946;
assign w17274 = w13203 & ~w13364;
assign v7947 = ~(w14524 | w14518);
assign w17275 = v7947;
assign w17276 = w14518 & ~w14645;
assign v7948 = ~(w15755 | w15749);
assign w17277 = v7948;
assign w17278 = w15749 & ~w15827;
assign v7949 = ~(w919 | w956);
assign w17279 = v7949;
assign v7950 = ~(w1447 | w1435);
assign w17280 = v7950;
assign v7951 = ~(w1576 | w1605);
assign w17281 = v7951;
assign w17282 = w866 & ~w855;
assign w17283 = w961 & ~w976;
assign v7952 = ~(w1054 | w1078);
assign w17284 = v7952;
assign w17285 = w997 & ~w1049;
assign v7953 = ~(w1223 | w1234);
assign w17286 = v7953;
assign w17287 = w1270 & ~w1259;
assign v7954 = ~(w1346 | w1381);
assign w17288 = v7954;
assign w17289 = w1535 & ~w17041;
assign w17290 = w1535 & w1450;
assign w17291 = ~w1535 & w17041;
assign v7955 = ~(w1535 | w1450);
assign w17292 = v7955;
assign w17293 = w1488 & ~w1477;
assign v7956 = ~(w1676 | w1724);
assign w17294 = v7956;
assign v7957 = ~(w1650 | w1653);
assign w17295 = v7957;
assign w17296 = w12688 & ~w16585;
assign w17297 = (w16590 & w16589) | (w16590 & w16585) | (w16589 & w16585);
assign w17298 = (w16592 & w16591) | (w16592 & ~w16585) | (w16591 & ~w16585);
assign w17299 = (w16597 & w16596) | (w16597 & w16585) | (w16596 & w16585);
assign w17300 = (~w16582 & w17440) | (~w16582 & w17441) | (w17440 & w17441);
assign w17301 = (w16599 & w16598) | (w16599 & ~w16585) | (w16598 & ~w16585);
assign w17302 = (w16582 & w17442) | (w16582 & w17443) | (w17442 & w17443);
assign w17303 = (w16603 & w16602) | (w16603 & w16585) | (w16602 & w16585);
assign w17304 = (w16603 & w16602) | (w16603 & w16584) | (w16602 & w16584);
assign v7958 = ~(w13975 | w17228);
assign w17305 = v7958;
assign v7959 = ~(w13975 | w17227);
assign w17306 = v7959;
assign v7960 = ~(w14257 | w17230);
assign w17307 = v7960;
assign v7961 = ~(w14257 | w17229);
assign w17308 = v7961;
assign v7962 = ~(w14389 | w17232);
assign w17309 = v7962;
assign v7963 = ~(w14389 | w17231);
assign w17310 = v7963;
assign v7964 = ~(w14646 | w17234);
assign w17311 = v7964;
assign v7965 = ~(w14646 | w17233);
assign w17312 = v7965;
assign v7966 = ~(w14764 | w17236);
assign w17313 = v7966;
assign v7967 = ~(w14764 | w17235);
assign w17314 = v7967;
assign v7968 = ~(w14994 | w17242);
assign w17315 = v7968;
assign v7969 = ~(w14994 | w17241);
assign w17316 = v7969;
assign v7970 = ~(w15103 | w17244);
assign w17317 = v7970;
assign v7971 = ~(w15103 | w17243);
assign w17318 = v7971;
assign w17319 = (~w16602 & w17702) | (~w16602 & w17703) | (w17702 & w17703);
assign w17320 = (w16632 & w16631) | (w16632 & w17246) | (w16631 & w17246);
assign w17321 = (~w16602 & w17704) | (~w16602 & w17705) | (w17704 & w17705);
assign w17322 = (w16638 & w16639) | (w16638 & w17246) | (w16639 & w17246);
assign w17323 = (~w16602 & w17706) | (~w16602 & w17707) | (w17706 & w17707);
assign w17324 = (w16654 & w16653) | (w16654 & w17246) | (w16653 & w17246);
assign w17325 = w16355 & w16996;
assign w17326 = w16355 & w16995;
assign v7972 = ~(w16355 | w16996);
assign w17327 = v7972;
assign v7973 = ~(w16355 | w16995);
assign w17328 = v7973;
assign w17329 = w16383 & w16998;
assign w17330 = w16383 & w16997;
assign v7974 = ~(w16383 | w16998);
assign w17331 = v7974;
assign v7975 = ~(w16383 | w16997);
assign w17332 = v7975;
assign w17333 = w16431 & w17000;
assign w17334 = w16431 & w16999;
assign v7976 = ~(w16431 | w17000);
assign w17335 = v7976;
assign v7977 = ~(w16431 | w16999);
assign w17336 = v7977;
assign w17337 = ~w1186 & w1185;
assign v7978 = ~(w12140 | w12135);
assign w17338 = v7978;
assign w17339 = w11949 & w17708;
assign w17340 = w13203 & ~w13364;
assign w17341 = (~w13364 & w17274) | (~w13364 & w13208) | (w17274 & w13208);
assign w17342 = w13364 & w13681;
assign w17343 = w17276 & ~w14645;
assign w17344 = (~w14645 & w17276) | (~w14645 & w14524) | (w17276 & w14524);
assign w17345 = w14645 & w14885;
assign v7979 = ~(w15827 | w17277);
assign w17346 = v7979;
assign w17347 = w15902 & w15827;
assign w17348 = w15902 & ~w17278;
assign v7980 = ~(w11118 | w16571);
assign w17349 = v7980;
assign w17350 = (~w11118 & w16570) | (~w11118 & w17548) | (w16570 & w17548);
assign w17351 = (w11541 & w16573) | (w11541 & w16571) | (w16573 & w16571);
assign w17352 = (~w16570 & w17549) | (~w16570 & w17550) | (w17549 & w17550);
assign w17353 = (w16578 & w16577) | (w16578 & ~w16571) | (w16577 & ~w16571);
assign w17354 = (w16570 & w17551) | (w16570 & w17552) | (w17551 & w17552);
assign w17355 = (w16580 & w16579) | (w16580 & w16571) | (w16579 & w16571);
assign w17356 = (~w16570 & w17553) | (~w16570 & w17554) | (w17553 & w17554);
assign w17357 = (w16585 & w16584) | (w16585 & ~w16571) | (w16584 & ~w16571);
assign w17358 = (w16585 & w16584) | (w16585 & ~w16572) | (w16584 & ~w16572);
assign w17359 = (~w16582 & w17709) | (~w16582 & w17710) | (w17709 & w17710);
assign v7981 = ~(w12507 | w17296);
assign w17360 = v7981;
assign w17361 = (w16582 & w17711) | (w16582 & w17712) | (w17711 & w17712);
assign v7982 = ~(w12864 | w17297);
assign w17362 = v7982;
assign w17363 = (~w16582 & w17713) | (~w16582 & w17714) | (w17713 & w17714);
assign v7983 = ~(w13035 | w17298);
assign w17364 = v7983;
assign v7984 = ~(w13363 | w17299);
assign w17365 = v7984;
assign v7985 = ~(w13525 | w17301);
assign w17366 = v7985;
assign w17367 = (~w16584 & w17444) | (~w16584 & w17445) | (w17444 & w17445);
assign w17368 = (~w16602 & w17715) | (~w16602 & w17444) | (w17715 & w17444);
assign w17369 = (~w16584 & w17446) | (~w16584 & w17447) | (w17446 & w17447);
assign w17370 = (~w16602 & w17716) | (~w16602 & w17446) | (w17716 & w17446);
assign w17371 = (~w16584 & w17448) | (~w16584 & w17449) | (w17448 & w17449);
assign w17372 = (~w16602 & w17717) | (~w16602 & w17448) | (w17717 & w17448);
assign w17373 = (~w16584 & w17450) | (~w16584 & w17451) | (w17450 & w17451);
assign w17374 = (~w16602 & w17718) | (~w16602 & w17450) | (w17718 & w17450);
assign w17375 = w15407 & w17252;
assign w17376 = w15407 & w17251;
assign v7986 = ~(w15407 | w17252);
assign w17377 = v7986;
assign v7987 = ~(w15407 | w17251);
assign w17378 = v7987;
assign w17379 = w15500 & w17254;
assign w17380 = w15500 & w17253;
assign v7988 = ~(w15500 | w17254);
assign w17381 = v7988;
assign v7989 = ~(w15500 | w17253);
assign w17382 = v7989;
assign w17383 = w15672 & w17256;
assign w17384 = w15672 & w17255;
assign v7990 = ~(w15672 | w17256);
assign w17385 = v7990;
assign v7991 = ~(w15672 | w17255);
assign w17386 = v7991;
assign w17387 = w15751 & w17258;
assign w17388 = w15751 & w17257;
assign v7992 = ~(w15751 | w17258);
assign w17389 = v7992;
assign v7993 = ~(w15751 | w17257);
assign w17390 = v7993;
assign w17391 = w15898 & w17260;
assign w17392 = w15898 & w17259;
assign v7994 = ~(w15898 | w17260);
assign w17393 = v7994;
assign v7995 = ~(w15898 | w17259);
assign w17394 = v7995;
assign w17395 = w15967 & w17262;
assign w17396 = w15967 & w17261;
assign v7996 = ~(w15967 | w17262);
assign w17397 = v7996;
assign v7997 = ~(w15967 | w17261);
assign w17398 = v7997;
assign w17399 = (w16986 & w16985) | (w16986 & ~w17304) | (w16985 & ~w17304);
assign w17400 = (w16988 & w16987) | (w16988 & ~w17304) | (w16987 & ~w17304);
assign w17401 = w16091 & ~w17264;
assign w17402 = w16091 & ~w17263;
assign w17403 = w16144 & w17266;
assign w17404 = w16144 & w17265;
assign v7998 = ~(w16144 | w17266);
assign w17405 = v7998;
assign v7999 = ~(w16144 | w17265);
assign w17406 = v7999;
assign w17407 = w16240 & w17268;
assign w17408 = w16240 & w17267;
assign v8000 = ~(w16240 | w17268);
assign w17409 = v8000;
assign v8001 = ~(w16240 | w17267);
assign w17410 = v8001;
assign w17411 = w16284 & w17270;
assign w17412 = w16284 & w17269;
assign v8002 = ~(w16284 | w17270);
assign w17413 = v8002;
assign v8003 = ~(w16284 | w17269);
assign w17414 = v8003;
assign w17415 = (w16994 & w16993) | (w16994 & ~w17304) | (w16993 & ~w17304);
assign w17416 = ~w16411 & w17272;
assign w17417 = ~w16411 & w17271;
assign w17418 = w16411 & ~w17272;
assign w17419 = w16411 & ~w17271;
assign w17420 = ~w10911 & w11121;
assign w17421 = w17339 & ~w12324;
assign w17422 = (~w12324 & w17339) | (~w12324 & w12140) | (w17339 & w12140);
assign w17423 = w13685 & ~w13681;
assign w17424 = (w13685 & ~w13681) | (w13685 & w17719) | (~w13681 & w17719);
assign w17425 = w14996 & ~w14885;
assign w17426 = w14996 & ~w17345;
assign w17427 = ~w15902 & w15971;
assign w17428 = w15971 & ~w17348;
assign w17429 = w15971 & ~w17347;
assign v8004 = ~(w9659 | w9688);
assign w17430 = v8004;
assign v8005 = ~(w9880 | w9861);
assign w17431 = v8005;
assign v8006 = ~(w10147 | w10129);
assign w17432 = v8006;
assign v8007 = ~(w10416 | w10454);
assign w17433 = v8007;
assign v8008 = ~(w10640 | w10676);
assign w17434 = v8008;
assign w17435 = w12324 & w12688;
assign w17436 = w16589 & w16590;
assign w17437 = (w16590 & w16589) | (w16590 & ~w12324) | (w16589 & ~w12324);
assign w17438 = w16591 | w16592;
assign w17439 = (w16592 & w16591) | (w16592 & w12324) | (w16591 & w12324);
assign w17440 = w16596 & w16597;
assign w17441 = (w16597 & w16596) | (w16597 & ~w12324) | (w16596 & ~w12324);
assign w17442 = w16598 | w16599;
assign w17443 = (w16599 & w16598) | (w16599 & w12324) | (w16598 & w12324);
assign v8009 = ~(w13832 | w16603);
assign w17444 = v8009;
assign w17445 = (~w13832 & w16600) | (~w13832 & w17720) | (w16600 & w17720);
assign w17446 = (w16605 & w16606) | (w16605 & ~w16603) | (w16606 & ~w16603);
assign w17447 = (w16600 & w17721) | (w16600 & w17722) | (w17721 & w17722);
assign w17448 = (w16612 & w16613) | (w16612 & ~w16603) | (w16613 & ~w16603);
assign w17449 = (w16600 & w17723) | (w16600 & w17724) | (w17723 & w17724);
assign w17450 = (w16620 & w16619) | (w16620 & ~w16603) | (w16619 & ~w16603);
assign w17451 = (w16600 & w17725) | (w16600 & w17726) | (w17725 & w17726);
assign w17452 = w9743 & ~w9733;
assign w17453 = (w10013 & w16561) | (w10013 & w17555) | (w16561 & w17555);
assign w17454 = (~w16559 & w17555) | (~w16559 & w17727) | (w17555 & w17727);
assign w17455 = w9946 & ~w9934;
assign w17456 = (~w10233 & w10097) | (~w10233 & w17556) | (w10097 & w17556);
assign w17457 = (~w10090 & ~w10056) | (~w10090 & w17557) | (~w10056 & w17557);
assign w17458 = w10126 & ~w10115;
assign v8010 = ~(w10202 | w10222);
assign w17459 = v8010;
assign w17460 = (~w10403 & w10404) | (~w10403 & w17558) | (w10404 & w17558);
assign w17461 = (~w10332 & w10298) | (~w10332 & w17559) | (w10298 & w17559);
assign w17462 = w10363 & ~w10351;
assign w17463 = w10372 & w10529;
assign v8011 = ~(w10372 | w10529);
assign w17464 = v8011;
assign w17465 = (~w16561 & w17560) | (~w16561 & w17561) | (w17560 & w17561);
assign w17466 = (w16566 & w16567) | (w16566 & w16562) | (w16567 & w16562);
assign w17467 = (~w10627 & w10628) | (~w10627 & w17562) | (w10628 & w17562);
assign w17468 = (~w10556 & w10524) | (~w10556 & w17563) | (w10524 & w17563);
assign v8012 = ~(w10547 | w10543);
assign w17469 = v8012;
assign w17470 = w10673 & ~w10662;
assign w17471 = w10501 & w10797;
assign v8013 = ~(w10501 | w10797);
assign w17472 = v8013;
assign w17473 = (w16568 & w16569) | (w16568 & ~w16562) | (w16569 & ~w16562);
assign v8014 = ~(w10755 | w10758);
assign w17474 = v8014;
assign w17475 = (w16572 & w16571) | (w16572 & ~w16563) | (w16571 & ~w16563);
assign w17476 = (w16572 & w16571) | (w16572 & ~w16562) | (w16571 & ~w16562);
assign v8015 = ~(w11119 | w17350);
assign w17477 = v8015;
assign v8016 = ~(w11119 | w17349);
assign w17478 = v8016;
assign v8017 = ~(w11333 | w17352);
assign w17479 = v8017;
assign v8018 = ~(w11333 | w17351);
assign w17480 = v8018;
assign v8019 = ~(w11742 | w17354);
assign w17481 = v8019;
assign v8020 = ~(w11742 | w17353);
assign w17482 = v8020;
assign v8021 = ~(w11940 | w17356);
assign w17483 = v8021;
assign v8022 = ~(w11940 | w17355);
assign w17484 = v8022;
assign v8023 = ~(w12323 | w17358);
assign w17485 = v8023;
assign w17486 = (~w16584 & w17564) | (~w16584 & w17565) | (w17564 & w17565);
assign w17487 = (w16587 & w16588) | (w16587 & ~w17358) | (w16588 & ~w17358);
assign w17488 = (~w16584 & w17566) | (~w16584 & w17567) | (w17566 & w17567);
assign w17489 = (w16594 & w16595) | (w16594 & ~w17358) | (w16595 & ~w17358);
assign w17490 = (~w16584 & w17568) | (~w16584 & w17569) | (w17568 & w17569);
assign w17491 = (w16601 & w16600) | (w16601 & ~w17358) | (w16600 & ~w17358);
assign w17492 = (~w16584 & w17570) | (~w16584 & w17571) | (w17570 & w17571);
assign w17493 = w14121 & w17306;
assign w17494 = w14121 & w17305;
assign v8024 = ~(w14121 | w17306);
assign w17495 = v8024;
assign v8025 = ~(w14121 | w17305);
assign w17496 = v8025;
assign w17497 = w14390 & w17308;
assign w17498 = w14390 & w17307;
assign v8026 = ~(w14390 | w17308);
assign w17499 = v8026;
assign v8027 = ~(w14390 | w17307);
assign w17500 = v8027;
assign w17501 = w14519 & w17310;
assign w17502 = w14519 & w17309;
assign v8028 = ~(w14519 | w17310);
assign w17503 = v8028;
assign v8029 = ~(w14519 | w17309);
assign w17504 = v8029;
assign w17505 = w14766 & w17312;
assign w17506 = w14766 & w17311;
assign v8030 = ~(w14766 | w17312);
assign w17507 = v8030;
assign v8031 = ~(w14766 | w17311);
assign w17508 = v8031;
assign w17509 = w14884 & w17314;
assign w17510 = w14884 & w17313;
assign v8032 = ~(w14884 | w17314);
assign w17511 = v8032;
assign v8033 = ~(w14884 | w17313);
assign w17512 = v8033;
assign w17513 = w15105 & w17316;
assign w17514 = w15105 & w17315;
assign v8034 = ~(w15105 | w17316);
assign w17515 = v8034;
assign v8035 = ~(w15105 | w17315);
assign w17516 = v8035;
assign w17517 = w15208 & w17318;
assign w17518 = w15208 & w17317;
assign v8036 = ~(w15208 | w17318);
assign w17519 = v8036;
assign v8037 = ~(w15208 | w17317);
assign w17520 = v8037;
assign w17521 = (w17247 & w17246) | (w17247 & ~w17358) | (w17246 & ~w17358);
assign w17522 = (w17247 & w17246) | (w17247 & ~w17357) | (w17246 & ~w17357);
assign w17523 = w15587 & w17320;
assign w17524 = w15587 & w17319;
assign v8038 = ~(w15587 | w17320);
assign w17525 = v8038;
assign v8039 = ~(w15587 | w17319);
assign w17526 = v8039;
assign w17527 = ~w15828 & w17322;
assign w17528 = ~w15828 & w17321;
assign w17529 = w15828 & ~w17322;
assign w17530 = w15828 & ~w17321;
assign w17531 = ~w16195 & w17324;
assign w17532 = ~w16195 & w17323;
assign w17533 = w16195 & ~w17324;
assign w17534 = w16195 & ~w17323;
assign w17535 = w9532 & ~w9770;
assign v8040 = ~(w11121 | w10908);
assign w17536 = v8040;
assign v8041 = ~(w13679 | w17423);
assign w17537 = v8041;
assign v8042 = ~(w13679 | w17424);
assign w17538 = v8042;
assign w17539 = w13679 & ~w13831;
assign v8043 = ~(w14882 | w14996);
assign w17540 = v8043;
assign v8044 = ~(w14882 | w17425);
assign w17541 = v8044;
assign w17542 = w14993 & w15109;
assign v8045 = ~(w15966 | w15971);
assign w17543 = v8045;
assign v8046 = ~(w15966 | w17427);
assign w17544 = v8046;
assign w17545 = w15966 & ~w16027;
assign v8047 = ~(w7539 | w7575);
assign w17546 = v8047;
assign w17547 = w8745 & ~w8743;
assign w17548 = w10908 & ~w11118;
assign w17549 = w16573 & w11541;
assign w17550 = (w11541 & w16573) | (w11541 & ~w10908) | (w16573 & ~w10908);
assign w17551 = w16577 | w16578;
assign w17552 = (w16578 & w16577) | (w16578 & w10908) | (w16577 & w10908);
assign w17553 = w16579 & w16580;
assign w17554 = (w16580 & w16579) | (w16580 & ~w10908) | (w16579 & ~w10908);
assign w17555 = w9770 & w10013;
assign v8048 = ~(w10154 | w10233);
assign w17556 = v8048;
assign v8049 = ~(w10055 | w10090);
assign w17557 = v8049;
assign v8050 = ~(w10457 | w10403);
assign w17558 = v8050;
assign v8051 = ~(w10297 | w10332);
assign w17559 = v8051;
assign w17560 = w16567 & w16566;
assign w17561 = (w16566 & w16567) | (w16566 & ~w9770) | (w16567 & ~w9770);
assign v8052 = ~(w10679 | w10627);
assign w17562 = v8052;
assign v8053 = ~(w10523 | w10556);
assign w17563 = v8053;
assign w17564 = ~w12323 & w16571;
assign v8054 = ~(w12323 | w16585);
assign w17565 = v8054;
assign w17566 = (w16587 & w16588) | (w16587 & w16571) | (w16588 & w16571);
assign w17567 = (w16587 & w16588) | (w16587 & ~w16585) | (w16588 & ~w16585);
assign w17568 = (w16594 & w16595) | (w16594 & w16571) | (w16595 & w16571);
assign w17569 = (w16594 & w16595) | (w16594 & ~w16585) | (w16595 & ~w16585);
assign w17570 = (w16600 & w16601) | (w16600 & w16571) | (w16601 & w16571);
assign w17571 = (w16600 & w16601) | (w16600 & ~w16585) | (w16601 & ~w16585);
assign w17572 = w7015 & ~w7018;
assign w17573 = pi31 & ~w7654;
assign w17574 = ~pi31 & w7654;
assign w17575 = w7669 & ~w7680;
assign w17576 = w7723 & ~w7713;
assign w17577 = w7794 & ~w17145;
assign w17578 = w7794 & w7540;
assign w17579 = ~w7794 & w17145;
assign v8055 = ~(w7794 | w7540);
assign w17580 = v8055;
assign w17581 = w7536 & ~w7526;
assign w17582 = w7785 & ~w7789;
assign v8056 = ~(w7967 | w7963);
assign w17583 = v8056;
assign v8057 = ~(w7837 | w7906);
assign w17584 = v8057;
assign w17585 = w8119 & ~w8109;
assign w17586 = w8201 & ~w8204;
assign v8058 = ~(w8308 | w8327);
assign w17587 = v8058;
assign w17588 = (~w8332 & w8333) | (~w8332 & w17728) | (w8333 & w17728);
assign w17589 = w8437 & ~w8426;
assign v8059 = ~(w8751 | w8774);
assign w17590 = v8059;
assign w17591 = w8697 & ~w8685;
assign v8060 = ~(w8700 | w8663);
assign w17592 = v8060;
assign v8061 = ~(w8915 | w8918);
assign w17593 = v8061;
assign w17594 = w8861 & ~w8850;
assign w17595 = w8952 & ~w8941;
assign w17596 = (~w9020 & w9022) | (~w9020 & w17729) | (w9022 & w17729);
assign v8062 = ~(w9041 | w16557);
assign w17597 = v8062;
assign w17598 = (~w9041 & w16555) | (~w9041 & w17730) | (w16555 & w17730);
assign v8063 = ~(w9263 | w9266);
assign w17599 = v8063;
assign w17600 = w9177 & ~w9166;
assign w17601 = w9209 & ~w9198;
assign w17602 = w9255 & ~w9258;
assign w17603 = (w9535 & w16558) | (w9535 & w16557) | (w16558 & w16557);
assign w17604 = (~w16555 & w17731) | (~w16555 & w17732) | (w17731 & w17732);
assign w17605 = (w16562 & w16563) | (w16562 & ~w16557) | (w16563 & ~w16557);
assign w17606 = (w16562 & w16563) | (w16562 & ~w16556) | (w16563 & ~w16556);
assign w17607 = (w17454 & w17453) | (w17454 & w16557) | (w17453 & w16557);
assign w17608 = (w17454 & w17453) | (w17454 & w16556) | (w17453 & w16556);
assign w17609 = w10323 & ~w10319;
assign w17610 = w10279 & w10559;
assign v8064 = ~(w10279 | w10559);
assign w17611 = v8064;
assign w17612 = (w17466 & w17465) | (w17466 & ~w16557) | (w17465 & ~w16557);
assign w17613 = (w17466 & w17465) | (w17466 & ~w16556) | (w17465 & ~w16556);
assign w17614 = w10587 & ~w10576;
assign w17615 = w10535 & ~w10531;
assign w17616 = w10528 & ~w10551;
assign w17617 = w10515 & ~w10518;
assign w17618 = w10506 & w10763;
assign v8065 = ~(w10506 | w10763);
assign w17619 = v8065;
assign v8066 = ~(w10693 | w17473);
assign w17620 = v8066;
assign w17621 = (w16563 & w17733) | (w16563 & w17734) | (w17733 & w17734);
assign w17622 = w10720 & w10962;
assign v8067 = ~(w10720 | w10962);
assign w17623 = v8067;
assign w17624 = w10703 & ~w10706;
assign w17625 = (~w10503 & w17735) | (~w10503 & w17736) | (w17735 & w17736);
assign v8068 = ~(w10778 | w10793);
assign w17626 = v8068;
assign w17627 = w11063 & ~w11105;
assign w17628 = (w16572 & w17737) | (w16572 & w17738) | (w17737 & w17738);
assign w17629 = (w16576 & w16575) | (w16576 & w17475) | (w16575 & w17475);
assign w17630 = (w16582 & w16583) | (w16582 & w17476) | (w16583 & w17476);
assign w17631 = (w16582 & w16583) | (w16582 & w17475) | (w16583 & w17475);
assign w17632 = (w17360 & w17359) | (w17360 & ~w17476) | (w17359 & ~w17476);
assign w17633 = (w17360 & w17359) | (w17360 & ~w17475) | (w17359 & ~w17475);
assign w17634 = (w17362 & w17361) | (w17362 & w17476) | (w17361 & w17476);
assign w17635 = (w17362 & w17361) | (w17362 & w17475) | (w17361 & w17475);
assign w17636 = (w17364 & w17363) | (w17364 & ~w17476) | (w17363 & ~w17476);
assign w17637 = (w17364 & w17363) | (w17364 & ~w17475) | (w17363 & ~w17475);
assign w17638 = w13526 & w17365;
assign w17639 = ~w17300 & w17739;
assign v8069 = ~(w13526 | w17365);
assign w17640 = v8069;
assign w17641 = (~w13526 & w17300) | (~w13526 & w17740) | (w17300 & w17740);
assign w17642 = w13680 & w17366;
assign w17643 = ~w17302 & w17741;
assign v8070 = ~(w13680 | w17366);
assign w17644 = v8070;
assign w17645 = (~w13680 & w17302) | (~w13680 & w17742) | (w17302 & w17742);
assign w17646 = (w17304 & w17303) | (w17304 & ~w17476) | (w17303 & ~w17476);
assign w17647 = (w17304 & w17303) | (w17304 & ~w17475) | (w17303 & ~w17475);
assign w17648 = w13977 & w17368;
assign w17649 = w13977 & w17367;
assign v8071 = ~(w13977 | w17368);
assign w17650 = v8071;
assign v8072 = ~(w13977 | w17367);
assign w17651 = v8072;
assign w17652 = ~w14258 & w17370;
assign w17653 = ~w14258 & w17369;
assign w17654 = w14258 & ~w17370;
assign w17655 = w14258 & ~w17369;
assign w17656 = ~w14647 & w17372;
assign w17657 = ~w14647 & w17371;
assign w17658 = w14647 & ~w17372;
assign w17659 = w14647 & ~w17371;
assign w17660 = w14995 & w17374;
assign w17661 = w14995 & w17373;
assign v8073 = ~(w14995 | w17374);
assign w17662 = v8073;
assign v8074 = ~(w14995 | w17373);
assign w17663 = v8074;
assign w17664 = (w17303 & w17743) | (w17303 & w17744) | (w17743 & w17744);
assign w17665 = (w17304 & w17743) | (w17304 & w17744) | (w17743 & w17744);
assign w17666 = (~w17303 & w17745) | (~w17303 & w17746) | (w17745 & w17746);
assign w17667 = w16029 & w17399;
assign w17668 = (~w17303 & w17747) | (~w17303 & w17748) | (w17747 & w17748);
assign w17669 = ~w16086 & w17400;
assign w17670 = (~w17303 & w17749) | (~w17303 & w17750) | (w17749 & w17750);
assign w17671 = (~w17304 & w17749) | (~w17304 & w17750) | (w17749 & w17750);
assign w17672 = (w17303 & w17751) | (w17303 & w17752) | (w17751 & w17752);
assign w17673 = w16321 & ~w17415;
assign v8075 = ~(w13679 | w13685);
assign w17674 = v8075;
assign w17675 = (~w13831 & w17539) | (~w13831 & w13685) | (w17539 & w13685);
assign w17676 = (~w13831 & w17539) | (~w13831 & w17423) | (w17539 & w17423);
assign w17677 = w17542 & w15109;
assign w17678 = (w15109 & w17542) | (w15109 & ~w14882) | (w17542 & ~w14882);
assign v8076 = ~(w16027 | w17543);
assign w17679 = v8076;
assign v8077 = ~(w16027 | w17544);
assign w17680 = v8077;
assign w17681 = (~w16027 & w17545) | (~w16027 & w17429) | (w17545 & w17429);
assign w17682 = (~w16027 & w17545) | (~w16027 & w17428) | (w17545 & w17428);
assign w17683 = w6747 & ~w6745;
assign v8078 = ~(w6878 | w6914);
assign w17684 = v8078;
assign v8079 = ~(w7197 | w7234);
assign w17685 = v8079;
assign v8080 = ~(w11290 | w11320);
assign w17686 = v8080;
assign v8081 = ~(w11719 | w11708);
assign w17687 = v8081;
assign w17688 = w12118 & ~w12116;
assign w17689 = w13831 & w13982;
assign w17690 = w16608 & w16607;
assign w17691 = (w16607 & w16608) | (w16607 & ~w13831) | (w16608 & ~w13831);
assign w17692 = w16609 | w16610;
assign w17693 = (w16610 & w16609) | (w16610 & w13831) | (w16609 & w13831);
assign w17694 = w16614 & w16615;
assign w17695 = (w16615 & w16614) | (w16615 & ~w13831) | (w16614 & ~w13831);
assign w17696 = w16616 | w16617;
assign w17697 = (w16617 & w16616) | (w16617 & w13831) | (w16616 & w13831);
assign w17698 = w16621 & w16622;
assign w17699 = (w16622 & w16621) | (w16622 & ~w13831) | (w16621 & ~w13831);
assign w17700 = w16623 | w16624;
assign w17701 = (w16624 & w16623) | (w16624 & w13831) | (w16623 & w13831);
assign w17702 = (w16632 & w16631) | (w16632 & w16628) | (w16631 & w16628);
assign w17703 = (w16632 & w16631) | (w16632 & w16627) | (w16631 & w16627);
assign w17704 = (w16638 & w16639) | (w16638 & w16628) | (w16639 & w16628);
assign w17705 = (w16638 & w16639) | (w16638 & w16627) | (w16639 & w16627);
assign w17706 = (w16654 & w16653) | (w16654 & w16628) | (w16653 & w16628);
assign w17707 = (w16654 & w16653) | (w16654 & w16627) | (w16653 & w16627);
assign v8082 = ~(w12133 | w12324);
assign w17708 = v8082;
assign v8083 = ~(w12507 | w12688);
assign w17709 = v8083;
assign v8084 = ~(w12507 | w17435);
assign w17710 = v8084;
assign v8085 = ~(w12864 | w17437);
assign w17711 = v8085;
assign v8086 = ~(w12864 | w17436);
assign w17712 = v8086;
assign v8087 = ~(w13035 | w17439);
assign w17713 = v8087;
assign v8088 = ~(w13035 | w17438);
assign w17714 = v8088;
assign v8089 = ~(w13832 | w16585);
assign w17715 = v8089;
assign w17716 = (w16605 & w16606) | (w16605 & ~w16585) | (w16606 & ~w16585);
assign w17717 = (w16612 & w16613) | (w16612 & ~w16585) | (w16613 & ~w16585);
assign w17718 = (w16620 & w16619) | (w16620 & ~w16585) | (w16619 & ~w16585);
assign w17719 = ~w13364 & w13685;
assign w17720 = w13831 & ~w13832;
assign w17721 = w16606 | w16605;
assign w17722 = (w16605 & w16606) | (w16605 & w13831) | (w16606 & w13831);
assign w17723 = w16613 | w16612;
assign w17724 = (w16612 & w16613) | (w16612 & w13831) | (w16613 & w13831);
assign w17725 = w16619 | w16620;
assign w17726 = (w16620 & w16619) | (w16620 & w13831) | (w16619 & w13831);
assign w17727 = w10013 & ~w17535;
assign w17728 = w8334 & ~w8332;
assign w17729 = w9021 & ~w9020;
assign w17730 = w8789 & ~w9041;
assign w17731 = w16558 & w9535;
assign w17732 = (w9535 & w16558) | (w9535 & ~w8789) | (w16558 & ~w8789);
assign v8090 = ~(w10693 | w16568);
assign w17733 = v8090;
assign v8091 = ~(w10693 | w16569);
assign w17734 = v8091;
assign v8092 = ~(w10898 | w10797);
assign w17735 = v8092;
assign v8093 = ~(w10898 | w17471);
assign w17736 = v8093;
assign w17737 = (w16576 & w16575) | (w16576 & ~w16562) | (w16575 & ~w16562);
assign w17738 = (w16576 & w16575) | (w16576 & w16571) | (w16575 & w16571);
assign w17739 = ~w13363 & w13526;
assign w17740 = w13363 & ~w13526;
assign w17741 = ~w13525 & w13680;
assign w17742 = w13525 & ~w13680;
assign v8094 = ~(w16029 | w16986);
assign w17743 = v8094;
assign v8095 = ~(w16029 | w16985);
assign w17744 = v8095;
assign w17745 = w16029 & w16986;
assign w17746 = w16029 & w16985;
assign w17747 = ~w16086 & w16988;
assign w17748 = ~w16086 & w16987;
assign w17749 = ~w16321 & w16994;
assign w17750 = ~w16321 & w16993;
assign w17751 = w16321 & ~w16994;
assign w17752 = w16321 & ~w16993;
assign w17753 = w6234 & ~w6223;
assign v8096 = ~(w6156 | w6159);
assign w17754 = v8096;
assign w17755 = w6429 & ~w6418;
assign w17756 = w6396 & ~w6386;
assign v8097 = ~(w6636 | w6601);
assign w17757 = v8097;
assign w17758 = w6708 & ~w6697;
assign w17759 = w6633 & ~w6622;
assign v8098 = ~(w6993 | w6918);
assign w17760 = v8098;
assign v8099 = ~(w6860 | w6827);
assign w17761 = v8099;
assign w17762 = w6839 & ~w6835;
assign w17763 = w6950 & ~w6939;
assign w17764 = w6777 & ~w6789;
assign v8100 = ~(w7049 | w7095);
assign w17765 = v8100;
assign v8101 = ~(w7448 | w7481);
assign w17766 = v8101;
assign v8102 = ~(w7355 | w7422);
assign w17767 = v8102;
assign v8103 = ~(w7418 | w7391);
assign w17768 = v8103;
assign w17769 = w7459 & ~w7455;
assign v8104 = ~(w7471 | w7467);
assign w17770 = v8104;
assign w17771 = w7450 & ~w7475;
assign w17772 = w7615 & ~w7611;
assign w17773 = w7606 & ~w7631;
assign w17774 = w7505 & ~w7579;
assign w17775 = (~w8007 & w16550) | (~w8007 & w16549) | (w16550 & w16549);
assign w17776 = (~w8007 & w16550) | (~w8007 & w16548) | (w16550 & w16548);
assign v8105 = ~(w7784 | w7795);
assign w17777 = v8105;
assign v8106 = ~(w8253 | w8221);
assign w17778 = v8106;
assign w17779 = w8016 & ~w8082;
assign v8107 = ~(w8072 | w8075);
assign w17780 = v8107;
assign w17781 = (w16553 & w16554) | (w16553 & w16549) | (w16554 & w16549);
assign w17782 = (w16553 & w16554) | (w16553 & w16548) | (w16554 & w16548);
assign v8108 = ~(w8340 | w8297);
assign w17783 = v8108;
assign v8109 = ~(w8440 | w8405);
assign w17784 = v8109;
assign v8110 = ~(w8283 | w8279);
assign w17785 = v8110;
assign w17786 = w8482 & ~w8478;
assign w17787 = w8473 & ~w8498;
assign w17788 = w8291 & ~w8289;
assign w17789 = (w16557 & w16556) | (w16557 & w16549) | (w16556 & w16549);
assign w17790 = (w16557 & w16556) | (w16557 & w16548) | (w16556 & w16548);
assign v8111 = ~(w8570 | w8573);
assign w17791 = v8111;
assign v8112 = ~(w8549 | w8545);
assign w17792 = v8112;
assign v8113 = ~(w8561 | w8557);
assign w17793 = v8113;
assign w17794 = w9251 & ~w17596;
assign w17795 = w9251 & w9023;
assign w17796 = ~w9251 & w17596;
assign v8114 = ~(w9251 | w9023);
assign w17797 = v8114;
assign w17798 = w8971 & ~w8967;
assign v8115 = ~(w8999 | w9029);
assign w17799 = v8115;
assign v8116 = ~(w9042 | w17598);
assign w17800 = v8116;
assign v8117 = ~(w9042 | w17597);
assign w17801 = v8117;
assign v8118 = ~(w9071 | w9094);
assign w17802 = v8118;
assign w17803 = w9051 & ~w9054;
assign v8119 = ~(w9286 | w17604);
assign w17804 = v8119;
assign v8120 = ~(w9286 | w17603);
assign w17805 = v8120;
assign v8121 = ~(w9437 | w9440);
assign w17806 = v8121;
assign v8122 = ~(w9482 | w9519);
assign w17807 = v8122;
assign v8123 = ~(w9620 | w9571);
assign w17808 = v8123;
assign w17809 = w9543 & ~w9565;
assign v8124 = ~(w9771 | w17606);
assign w17810 = v8124;
assign v8125 = ~(w9771 | w17605);
assign w17811 = v8125;
assign v8126 = ~(w10005 | w17608);
assign w17812 = v8126;
assign v8127 = ~(w10005 | w17607);
assign w17813 = v8127;
assign w17814 = (w16564 & w16565) | (w16564 & ~w17606) | (w16565 & ~w17606);
assign w17815 = (w16564 & w16565) | (w16564 & ~w17605) | (w16565 & ~w17605);
assign w17816 = w10451 & ~w10439;
assign w17817 = w10394 & ~w10385;
assign v8128 = ~(w10471 | w17613);
assign w17818 = v8128;
assign v8129 = ~(w10471 | w17612);
assign w17819 = v8129;
assign v8130 = ~(w10685 | w10560);
assign w17820 = v8130;
assign v8131 = ~(w10826 | w10893);
assign w17821 = v8131;
assign v8132 = ~(w10711 | w10714);
assign w17822 = v8132;
assign v8133 = ~(w10901 | w10764);
assign w17823 = v8133;
assign v8134 = ~(w11059 | w10963);
assign w17824 = v8134;
assign v8135 = ~(w11053 | w11018);
assign w17825 = v8135;
assign w17826 = (w17478 & w17477) | (w17478 & ~w17606) | (w17477 & ~w17606);
assign w17827 = (w17478 & w17477) | (w17478 & ~w17605) | (w17477 & ~w17605);
assign v8136 = ~(w11326 | w11228);
assign w17828 = v8136;
assign w17829 = w11162 & ~w11150;
assign w17830 = w11287 & ~w11275;
assign w17831 = (w17480 & w17479) | (w17480 & w17606) | (w17479 & w17606);
assign w17832 = (w17480 & w17479) | (w17480 & w17605) | (w17479 & w17605);
assign w17833 = w11374 & ~w11363;
assign w17834 = (w17482 & w17481) | (w17482 & ~w17606) | (w17481 & ~w17606);
assign w17835 = (w17482 & w17481) | (w17482 & ~w17605) | (w17481 & ~w17605);
assign w17836 = (w17484 & w17483) | (w17484 & w17606) | (w17483 & w17606);
assign w17837 = (w17484 & w17483) | (w17484 & w17605) | (w17483 & w17605);
assign v8137 = ~(w11824 | w11793);
assign w17838 = v8137;
assign w17839 = w11924 & w12050;
assign v8138 = ~(w11924 | w12050);
assign w17840 = v8138;
assign w17841 = w12041 & ~w12030;
assign w17842 = w12008 & ~w11997;
assign v8139 = ~(w11962 | w11980);
assign w17843 = v8139;
assign v8140 = ~(w12104 | w12082);
assign w17844 = v8140;
assign w17845 = w12108 & ~w12111;
assign w17846 = (w17358 & w17357) | (w17358 & w17606) | (w17357 & w17606);
assign w17847 = (w17358 & w17357) | (w17358 & w17605) | (w17357 & w17605);
assign w17848 = w12240 & ~w12311;
assign w17849 = w12509 & w17486;
assign w17850 = w12509 & w17485;
assign v8141 = ~(w12509 | w17486);
assign w17851 = v8141;
assign v8142 = ~(w12509 | w17485);
assign w17852 = v8142;
assign w17853 = ~w12866 & w17488;
assign w17854 = ~w12866 & w17487;
assign w17855 = w12866 & ~w17488;
assign w17856 = w12866 & ~w17487;
assign w17857 = ~w13365 & w17490;
assign w17858 = ~w13365 & w17489;
assign w17859 = w13365 & ~w17490;
assign w17860 = w13365 & ~w17489;
assign w17861 = ~w13833 & w17492;
assign w17862 = ~w13833 & w17491;
assign w17863 = w13833 & ~w17492;
assign w17864 = w13833 & ~w17491;
assign w17865 = ~w15312 & w17522;
assign w17866 = ~w15312 & w17521;
assign w17867 = w15312 & ~w17522;
assign w17868 = w15312 & ~w17521;
assign w17869 = (w17002 & w17001) | (w17002 & ~w17522) | (w17001 & ~w17522);
assign w17870 = (w17002 & w17001) | (w17002 & ~w17521) | (w17001 & ~w17521);
assign w17871 = (w17004 & w17003) | (w17004 & w17522) | (w17003 & w17522);
assign w17872 = (w17004 & w17003) | (w17004 & w17521) | (w17003 & w17521);
assign w17873 = (w17006 & w17005) | (w17006 & w17522) | (w17005 & w17522);
assign w17874 = (w17006 & w17005) | (w17006 & w17521) | (w17005 & w17521);
assign w17875 = (w17008 & w17007) | (w17008 & ~w17522) | (w17007 & ~w17522);
assign w17876 = (w17008 & w17007) | (w17008 & ~w17521) | (w17007 & ~w17521);
assign w17877 = (w17010 & w17009) | (w17010 & w17522) | (w17009 & w17522);
assign w17878 = (w17010 & w17009) | (w17010 & w17521) | (w17009 & w17521);
assign w17879 = (w17012 & w17011) | (w17012 & ~w17522) | (w17011 & ~w17522);
assign w17880 = (w17012 & w17011) | (w17012 & ~w17521) | (w17011 & ~w17521);
assign w17881 = (w17014 & w17013) | (w17014 & w17522) | (w17013 & w17522);
assign w17882 = (w17014 & w17013) | (w17014 & w17521) | (w17013 & w17521);
assign w17883 = (w17016 & w17015) | (w17016 & ~w17522) | (w17015 & ~w17522);
assign w17884 = (w17016 & w17015) | (w17016 & ~w17521) | (w17015 & ~w17521);
assign w17885 = (w17018 & w17017) | (w17018 & ~w17522) | (w17017 & ~w17522);
assign w17886 = (w17018 & w17017) | (w17018 & ~w17521) | (w17017 & ~w17521);
assign one = 1;
assign po000 = pi00;// level 0
assign po001 = w0;// level 1
assign po002 = w4;// level 3
assign po003 = w10;// level 4
assign po004 = ~w22;// level 7
assign po005 = w38;// level 8
assign po006 = ~w55;// level 9
assign po007 = w83;// level 11
assign po008 = ~w114;// level 12
assign po009 = w151;// level 13
assign po010 = w188;// level 15
assign po011 = ~w234;// level 16
assign po012 = ~w282;// level 16
assign po013 = w336;// level 18
assign po014 = ~w391;// level 19
assign po015 = ~w453;// level 19
assign po016 = w517;// level 21
assign po017 = ~w588;// level 20
assign po018 = ~w660;// level 20
assign po019 = w739;// level 22
assign po020 = ~w820;// level 23
assign po021 = w907;// level 23
assign po022 = w995;// level 23
assign po023 = ~w1092;// level 24
assign po024 = ~w1190;// level 24
assign po025 = w1290;// level 26
assign po026 = ~w1398;// level 26
assign po027 = w1510;// level 26
assign po028 = w1622;// level 26
assign po029 = ~w1744;// level 27
assign po030 = w1867;// level 27
assign po031 = w1992;// level 29
assign po032 = ~w2126;// level 29
assign po033 = w2264;// level 29
assign po034 = w2401;// level 30
assign po035 = ~w2548;// level 30
assign po036 = w2694;// level 29
assign po037 = w2846;// level 31
assign po038 = ~w3002;// level 31
assign po039 = w3164;// level 30
assign po040 = w3327;// level 32
assign po041 = ~w3499;// level 32
assign po042 = ~w3669;// level 32
assign po043 = w3845;// level 33
assign po044 = ~w4028;// level 34
assign po045 = ~w4214;// level 33
assign po046 = ~w4403;// level 34
assign po047 = ~w4599;// level 35
assign po048 = ~w4797;// level 34
assign po049 = w5001;// level 36
assign po050 = ~w5205;// level 36
assign po051 = w5418;// level 35
assign po052 = w5634;// level 36
assign po053 = ~w5851;// level 37
assign po054 = w6074;// level 36
assign po055 = w6302;// level 37
assign po056 = ~w6533;// level 38
assign po057 = w6773;// level 37
assign po058 = w7010;// level 38
assign po059 = ~w7256;// level 39
assign po060 = w7503;// level 38
assign po061 = w7752;// level 39
assign po062 = ~w8011;// level 39
assign po063 = w8274;// level 38
assign po064 = w8534;// level 39
assign po065 = ~w8793;// level 39
assign po066 = ~w9046;// level 38
assign po067 = w9292;// level 39
assign po068 = ~w9539;// level 39
assign po069 = w9777;// level 39
assign po070 = w10012;// level 39
assign po071 = ~w10248;// level 39
assign po072 = ~w10476;// level 39
assign po073 = w10698;// level 39
assign po074 = ~w10915;// level 39
assign po075 = w11125;// level 39
assign po076 = w11339;// level 39
assign po077 = ~w11545;// level 39
assign po078 = ~w11746;// level 39
assign po079 = w11946;// level 39
assign po080 = ~w12139;// level 39
assign po081 = ~w12328;// level 39
assign po082 = w12512;// level 39
assign po083 = ~w12692;// level 39
assign po084 = ~w12869;// level 39
assign po085 = w13040;// level 39
assign po086 = ~w13207;// level 39
assign po087 = ~w13368;// level 39
assign po088 = w13529;// level 39
assign po089 = ~w13684;// level 39
assign po090 = ~w13836;// level 39
assign po091 = w13981;// level 39
assign po092 = ~w14124;// level 39
assign po093 = ~w14261;// level 39
assign po094 = w14393;// level 39
assign po095 = ~w14523;// level 39
assign po096 = ~w14650;// level 39
assign po097 = w14769;// level 39
assign po098 = ~w14888;// level 39
assign po099 = w14999;// level 39
assign po100 = w15108;// level 39
assign po101 = ~w15211;// level 39
assign po102 = ~w15315;// level 39
assign po103 = w15410;// level 39
assign po104 = ~w15503;// level 39
assign po105 = w15591;// level 39
assign po106 = w15675;// level 39
assign po107 = ~w15754;// level 39
assign po108 = ~w15831;// level 39
assign po109 = w15901;// level 39
assign po110 = ~w15970;// level 39
assign po111 = w16032;// level 39
assign po112 = w16093;// level 39
assign po113 = ~w16147;// level 39
assign po114 = ~w16198;// level 39
assign po115 = w16243;// level 39
assign po116 = ~w16287;// level 39
assign po117 = ~w16324;// level 39
assign po118 = w16358;// level 40
assign po119 = ~w16387;// level 40
assign po120 = ~w16414;// level 39
assign po121 = w16434;// level 40
assign po122 = ~w16453;// level 39
assign po123 = ~w16465;// level 39
assign po124 = ~w16473;// level 39
assign po125 = ~w16479;// level 39
assign po126 = w16481;// level 39
endmodule
