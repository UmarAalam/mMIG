//Written by the Majority Logic Package Thu Apr 30 13:39:35 2015
module top (
            pi000, pi001, pi002, pi003, pi004, pi005, pi006, pi007, pi008, pi009, pi010, pi011, pi012, pi013, pi014, pi015, pi016, pi017, pi018, pi019, pi020, pi021, pi022, pi023, pi024, pi025, pi026, pi027, pi028, pi029, pi030, pi031, pi032, pi033, pi034, pi035, pi036, pi037, pi038, pi039, pi040, pi041, pi042, pi043, pi044, pi045, pi046, pi047, pi048, pi049, pi050, pi051, pi052, pi053, pi054, pi055, pi056, pi057, pi058, pi059, pi060, pi061, pi062, pi063, pi064, pi065, pi066, pi067, pi068, pi069, pi070, pi071, pi072, pi073, pi074, pi075, pi076, pi077, pi078, pi079, pi080, pi081, pi082, pi083, pi084, pi085, pi086, pi087, pi088, pi089, pi090, pi091, pi092, pi093, pi094, pi095, pi096, pi097, pi098, pi099, pi100, pi101, pi102, pi103, pi104, pi105, pi106, pi107, pi108, pi109, pi110, pi111, pi112, pi113, pi114, pi115, pi116, pi117, pi118, pi119, pi120, pi121, pi122, pi123, pi124, pi125, pi126, pi127, pi128, pi129, pi130, pi131, pi132, pi133, pi134, pi135, pi136, pi137, pi138, pi139, pi140, pi141, pi142, pi143, pi144, pi145, pi146, pi147, pi148, pi149, pi150, pi151, pi152, pi153, pi154, pi155, pi156, pi157, pi158, pi159, pi160, pi161, pi162, pi163, pi164, pi165, pi166, pi167, pi168, pi169, pi170, pi171, pi172, pi173, pi174, pi175, pi176, pi177, pi178, pi179, pi180, pi181, pi182, pi183, pi184, pi185, pi186, pi187, pi188, pi189, pi190, pi191, pi192, pi193, pi194, pi195, pi196, pi197, pi198, pi199, pi200, pi201, pi202, pi203, pi204, pi205, pi206, pi207, pi208, pi209, pi210, pi211, pi212, pi213, pi214, pi215, pi216, pi217, pi218, pi219, pi220, pi221, pi222, pi223, pi224, pi225, pi226, pi227, pi228, pi229, pi230, pi231, pi232, pi233, pi234, pi235, pi236, pi237, pi238, pi239, pi240, pi241, pi242, pi243, pi244, pi245, pi246, pi247, pi248, pi249, pi250, pi251, pi252, pi253, pi254, pi255, pi256, pi257, pi258, pi259, pi260, pi261, pi262, pi263, pi264, pi265, pi266, pi267, pi268, pi269, pi270, pi271, pi272, pi273, 
            po000, po001, po002, po003, po004, po005, po006, po007, po008, po009, po010, po011, po012, po013, po014, po015, po016, po017, po018, po019, po020, po021, po022, po023, po024, po025, po026, po027, po028, po029, po030, po031, po032, po033, po034, po035, po036, po037, po038, po039, po040, po041, po042, po043, po044, po045, po046, po047, po048, po049, po050, po051, po052, po053, po054, po055, po056, po057, po058, po059, po060, po061, po062, po063, po064, po065, po066, po067, po068, po069, po070, po071, po072, po073, po074, po075, po076, po077, po078, po079, po080, po081, po082, po083, po084, po085, po086, po087, po088, po089, po090, po091, po092, po093, po094, po095, po096, po097, po098, po099, po100, po101, po102, po103, po104, po105, po106, po107, po108, po109, po110, po111, po112, po113, po114, po115, po116, po117, po118, po119, po120, po121, po122, po123, po124, po125, po126, po127, po128, po129, po130, po131, po132, po133, po134, po135, po136, po137, po138, po139, po140, po141, po142, po143, po144, po145, po146, po147, po148, po149, po150, po151, po152, po153, po154, po155, po156, po157, po158, po159, po160, po161, po162, po163, po164, po165, po166, po167, po168, po169, po170, po171, po172, po173, po174, po175, po176, po177, po178, po179, po180, po181, po182, po183, po184, po185, po186, po187, po188, po189, po190, po191, po192, po193, po194, po195, po196, po197, po198, po199, po200, po201, po202, po203, po204, po205, po206, po207, po208, po209, po210, po211, po212, po213, po214, po215, po216, po217, po218, po219, po220, po221, po222, po223, po224, po225, po226, po227, po228, po229, po230, po231, po232, po233, po234, po235, po236, po237, po238, po239, po240, po241, po242, po243, po244, po245, po246, po247, po248, po249, po250, po251, po252, po253, po254, po255, po256, po257, po258, po259, po260, po261, po262, po263, po264, po265, po266, po267, po268, po269, po270, po271, po272, po273, po274, po275);
input pi000, pi001, pi002, pi003, pi004, pi005, pi006, pi007, pi008, pi009, pi010, pi011, pi012, pi013, pi014, pi015, pi016, pi017, pi018, pi019, pi020, pi021, pi022, pi023, pi024, pi025, pi026, pi027, pi028, pi029, pi030, pi031, pi032, pi033, pi034, pi035, pi036, pi037, pi038, pi039, pi040, pi041, pi042, pi043, pi044, pi045, pi046, pi047, pi048, pi049, pi050, pi051, pi052, pi053, pi054, pi055, pi056, pi057, pi058, pi059, pi060, pi061, pi062, pi063, pi064, pi065, pi066, pi067, pi068, pi069, pi070, pi071, pi072, pi073, pi074, pi075, pi076, pi077, pi078, pi079, pi080, pi081, pi082, pi083, pi084, pi085, pi086, pi087, pi088, pi089, pi090, pi091, pi092, pi093, pi094, pi095, pi096, pi097, pi098, pi099, pi100, pi101, pi102, pi103, pi104, pi105, pi106, pi107, pi108, pi109, pi110, pi111, pi112, pi113, pi114, pi115, pi116, pi117, pi118, pi119, pi120, pi121, pi122, pi123, pi124, pi125, pi126, pi127, pi128, pi129, pi130, pi131, pi132, pi133, pi134, pi135, pi136, pi137, pi138, pi139, pi140, pi141, pi142, pi143, pi144, pi145, pi146, pi147, pi148, pi149, pi150, pi151, pi152, pi153, pi154, pi155, pi156, pi157, pi158, pi159, pi160, pi161, pi162, pi163, pi164, pi165, pi166, pi167, pi168, pi169, pi170, pi171, pi172, pi173, pi174, pi175, pi176, pi177, pi178, pi179, pi180, pi181, pi182, pi183, pi184, pi185, pi186, pi187, pi188, pi189, pi190, pi191, pi192, pi193, pi194, pi195, pi196, pi197, pi198, pi199, pi200, pi201, pi202, pi203, pi204, pi205, pi206, pi207, pi208, pi209, pi210, pi211, pi212, pi213, pi214, pi215, pi216, pi217, pi218, pi219, pi220, pi221, pi222, pi223, pi224, pi225, pi226, pi227, pi228, pi229, pi230, pi231, pi232, pi233, pi234, pi235, pi236, pi237, pi238, pi239, pi240, pi241, pi242, pi243, pi244, pi245, pi246, pi247, pi248, pi249, pi250, pi251, pi252, pi253, pi254, pi255, pi256, pi257, pi258, pi259, pi260, pi261, pi262, pi263, pi264, pi265, pi266, pi267, pi268, pi269, pi270, pi271, pi272, pi273;
output po000, po001, po002, po003, po004, po005, po006, po007, po008, po009, po010, po011, po012, po013, po014, po015, po016, po017, po018, po019, po020, po021, po022, po023, po024, po025, po026, po027, po028, po029, po030, po031, po032, po033, po034, po035, po036, po037, po038, po039, po040, po041, po042, po043, po044, po045, po046, po047, po048, po049, po050, po051, po052, po053, po054, po055, po056, po057, po058, po059, po060, po061, po062, po063, po064, po065, po066, po067, po068, po069, po070, po071, po072, po073, po074, po075, po076, po077, po078, po079, po080, po081, po082, po083, po084, po085, po086, po087, po088, po089, po090, po091, po092, po093, po094, po095, po096, po097, po098, po099, po100, po101, po102, po103, po104, po105, po106, po107, po108, po109, po110, po111, po112, po113, po114, po115, po116, po117, po118, po119, po120, po121, po122, po123, po124, po125, po126, po127, po128, po129, po130, po131, po132, po133, po134, po135, po136, po137, po138, po139, po140, po141, po142, po143, po144, po145, po146, po147, po148, po149, po150, po151, po152, po153, po154, po155, po156, po157, po158, po159, po160, po161, po162, po163, po164, po165, po166, po167, po168, po169, po170, po171, po172, po173, po174, po175, po176, po177, po178, po179, po180, po181, po182, po183, po184, po185, po186, po187, po188, po189, po190, po191, po192, po193, po194, po195, po196, po197, po198, po199, po200, po201, po202, po203, po204, po205, po206, po207, po208, po209, po210, po211, po212, po213, po214, po215, po216, po217, po218, po219, po220, po221, po222, po223, po224, po225, po226, po227, po228, po229, po230, po231, po232, po233, po234, po235, po236, po237, po238, po239, po240, po241, po242, po243, po244, po245, po246, po247, po248, po249, po250, po251, po252, po253, po254, po255, po256, po257, po258, po259, po260, po261, po262, po263, po264, po265, po266, po267, po268, po269, po270, po271, po272, po273, po274, po275;
wire one, w0, w1, w2, w3, w4, w5, w6, w7, w8, w9, w10, w11, w12, w13, w14, w15, w16, w17, w18, w19, w20, w21, w22, w23, w24, w25, w26, w27, w28, w29, w30, w31, w32, w33, w34, w35, w36, w37, w38, w39, w40, w41, w42, w43, w44, w45, w46, w47, w48, w49, w50, w51, w52, w53, w54, w55, w56, w57, w58, w59, w60, w61, w62, w63, w64, w65, w66, w67, w68, w69, w70, w71, w72, w73, w74, w75, w76, w77, w78, w79, w80, w81, w82, w83, w84, w85, w86, w87, w88, w89, w90, w91, w92, w93, w94, w95, w96, w97, w98, w99, w100, w101, w102, w103, w104, w105, w106, w107, w108, w109, w110, w111, w112, w113, w114, w115, w116, w117, w118, w119, w120, w121, w122, w123, w124, w125, w126, w127, w128, w129, w130, w131, w132, w133, w134, w135, w136, w137, w138, w139, w140, w141, w142, w143, w144, w145, w146, w147, w148, w149, w150, w151, w152, w153, w154, w155, w156, w157, w158, w159, w160, w161, w162, w163, w164, w165, w166, w167, w168, w169, w170, w171, w172, w173, w174, w175, w176, w177, w178, w179, w180, w181, w182, w183, w184, w185, w186, w187, w188, w189, w190, w191, w192, w193, w194, w195, w196, w197, w198, w199, w200, w201, w202, w203, w204, w205, w206, w207, w208, w209, w210, w211, w212, w213, w214, w215, w216, w217, w218, w219, w220, w221, w222, w223, w224, w225, w226, w227, w228, w229, w230, w231, w232, w233, w234, w235, w236, w237, w238, w239, w240, w241, w242, w243, w244, w245, w246, w247, w248, w249, w250, w251, w252, w253, w254, w255, w256, w257, w258, w259, w260, w261, w262, w263, w264, w265, w266, w267, w268, w269, w270, w271, w272, w273, w274, w275, w276, w277, w278, w279, w280, w281, w282, w283, w284, w285, w286, w287, w288, w289, w290, w291, w292, w293, w294, w295, w296, w297, w298, w299, w300, w301, w302, w303, w304, w305, w306, w307, w308, w309, w310, w311, w312, w313, w314, w315, w316, w317, w318, w319, w320, w321, w322, w323, w324, w325, w326, w327, w328, w329, w330, w331, w332, w333, w334, w335, w336, w337, w338, w339, w340, w341, w342, w343, w344, w345, w346, w347, w348, w349, w350, w351, w352, w353, w354, w355, w356, w357, w358, w359, w360, w361, w362, w363, w364, w365, w366, w367, w368, w369, w370, w371, w372, w373, w374, w375, w376, w377, w378, w379, w380, w381, w382, w383, w384, w385, w386, w387, w388, w389, w390, w391, w392, w393, w394, w395, w396, w397, w398, w399, w400, w401, w402, w403, w404, w405, w406, w407, w408, w409, w410, w411, w412, w413, w414, w415, w416, w417, w418, w419, w420, w421, w422, w423, w424, w425, w426, w427, w428, w429, w430, w431, w432, w433, w434, w435, w436, w437, w438, w439, w440, w441, w442, w443, w444, w445, w446, w447, w448, w449, w450, w451, w452, w453, w454, w455, w456, w457, w458, w459, w460, w461, w462, w463, w464, w465, w466, w467, w468, w469, w470, w471, w472, w473, w474, w475, w476, w477, w478, w479, w480, w481, w482, w483, w484, w485, w486, w487, w488, w489, w490, w491, w492, w493, w494, w495, w496, w497, w498, w499, w500, w501, w502, w503, w504, w505, w506, w507, w508, w509, w510, w511, w512, w513, w514, w515, w516, w517, w518, w519, w520, w521, w522, w523, w524, w525, w526, w527, w528, w529, w530, w531, w532, w533, w534, w535, w536, w537, w538, w539, w540, w541, w542, w543, w544, w545, w546, w547, w548, w549, w550, w551, w552, w553, w554, w555, w556, w557, w558, w559, w560, w561, w562, w563, w564, w565, w566, w567, w568, w569, w570, w571, w572, w573, w574, w575, w576, w577, w578, w579, w580, w581, w582, w583, w584, w585, w586, w587, w588, w589, w590, w591, w592, w593, w594, w595, w596, w597, w598, w599, w600, w601, w602, w603, w604, w605, w606, w607, w608, w609, w610, w611, w612, w613, w614, w615, w616, w617, w618, w619, w620, w621, w622, w623, w624, w625, w626, w627, w628, w629, w630, w631, w632, w633, w634, w635, w636, w637, w638, w639, w640, w641, w642, w643, w644, w645, w646, w647, w648, w649, w650, w651, w652, w653, w654, w655, w656, w657, w658, w659, w660, w661, w662, w663, w664, w665, w666, w667, w668, w669, w670, w671, w672, w673, w674, w675, w676, w677, w678, w679, w680, w681, w682, w683, w684, w685, w686, w687, w688, w689, w690, w691, w692, w693, w694, w695, w696, w697, w698, w699, w700, w701, w702, w703, w704, w705, w706, w707, w708, w709, w710, w711, w712, w713, w714, w715, w716, w717, w718, w719, w720, w721, w722, w723, w724, w725, w726, w727, w728, w729, w730, w731, w732, w733, w734, w735, w736, w737, w738, w739, w740, w741, w742, w743, w744, w745, w746, w747, w748, w749, w750, w751, w752, w753, w754, w755, w756, w757, w758, w759, w760, w761, w762, w763, w764, w765, w766, w767, w768, w769, w770, w771, w772, w773, w774, w775, w776, w777, w778, w779, w780, w781, w782, w783, w784, w785, w786, w787, w788, w789, w790, w791, w792, w793, w794, w795, w796, w797, w798, w799, w800, w801, w802, w803, w804, w805, w806, w807, w808, w809, w810, w811, w812, w813, w814, w815, w816, w817, w818, w819, w820, w821, w822, w823, w824, w825, w826, w827, w828, w829, w830, w831, w832, w833, w834, w835, w836, w837, w838, w839, w840, w841, w842, w843, w844, w845, w846, w847, w848, w849, w850, w851, w852, w853, w854, w855, w856, w857, w858, w859, w860, w861, w862, w863, w864, w865, w866, w867, w868, w869, w870, w871, w872, w873, w874, w875, w876, w877, w878, w879, w880, w881, w882, w883, w884, w885, w886, w887, w888, w889, w890, w891, w892, w893, w894, w895, w896, w897, w898, w899, w900, w901, w902, w903, w904, w905, w906, w907, w908, w909, w910, w911, w912, w913, w914, w915, w916, w917, w918, w919, w920, w921, w922, w923, w924, w925, w926, w927, w928, w929, w930, w931, w932, w933, w934, w935, w936, w937, w938, w939, w940, w941, w942, w943, w944, w945, w946, w947, w948, w949, w950, w951, w952, w953, w954, w955, w956, w957, w958, w959, w960, w961, w962, w963, w964, w965, w966, w967, w968, w969, w970, w971, w972, w973, w974, w975, w976, w977, w978, w979, w980, w981, w982, w983, w984, w985, w986, w987, w988, w989, w990, w991, w992, w993, w994, w995, w996, w997, w998, w999, w1000, w1001, w1002, w1003, w1004, w1005, w1006, w1007, w1008, w1009, w1010, w1011, w1012, w1013, w1014, w1015, w1016, w1017, w1018, w1019, w1020, w1021, w1022, w1023, w1024, w1025, w1026, w1027, w1028, w1029, w1030, w1031, w1032, w1033, w1034, w1035, w1036, w1037, w1038, w1039, w1040, w1041, w1042, w1043, w1044, w1045, w1046, w1047, w1048, w1049, w1050, w1051, w1052, w1053, w1054, w1055, w1056, w1057, w1058, w1059, w1060, w1061, w1062, w1063, w1064, w1065, w1066, w1067, w1068, w1069, w1070, w1071, w1072, w1073, w1074, w1075, w1076, w1077, w1078, w1079, w1080, w1081, w1082, w1083, w1084, w1085, w1086, w1087, w1088, w1089, w1090, w1091, w1092, w1093, w1094, w1095, w1096, w1097, w1098, w1099, w1100, w1101, w1102, w1103, w1104, w1105, w1106, w1107, w1108, w1109, w1110, w1111, w1112, w1113, w1114, w1115, w1116, w1117, w1118, w1119, w1120, w1121, w1122, w1123, w1124, w1125, w1126, w1127, w1128, w1129, w1130, w1131, w1132, w1133, w1134, w1135, w1136, w1137, w1138, w1139, w1140, w1141, w1142, w1143, w1144, w1145, w1146, w1147, w1148, w1149, w1150, w1151, w1152, w1153, w1154, w1155, w1156, w1157, w1158, w1159, w1160, w1161, w1162, w1163, w1164, w1165, w1166, w1167, w1168, w1169, w1170, w1171, w1172, w1173, w1174, w1175, w1176, w1177, w1178, w1179, w1180, w1181, w1182, w1183, w1184, w1185, w1186, w1187, w1188, w1189, w1190, w1191, w1192, w1193, w1194, w1195, w1196, w1197, w1198, w1199, w1200, w1201, w1202, w1203, w1204, w1205, w1206, w1207, w1208, w1209, w1210, w1211, w1212, w1213, w1214, w1215, w1216, w1217, w1218, w1219, w1220, w1221, w1222, w1223, w1224, w1225, w1226, w1227, w1228, w1229, w1230, w1231, w1232, w1233, w1234, w1235, w1236, w1237, w1238, w1239, w1240, w1241, w1242, w1243, w1244, w1245, w1246, w1247, w1248, w1249, w1250, w1251, w1252, w1253, w1254, w1255, w1256, w1257, w1258, w1259, w1260, w1261, w1262, w1263, w1264, w1265, w1266, w1267, w1268, w1269, w1270, w1271, w1272, w1273, w1274, w1275, w1276, w1277, w1278, w1279, w1280, w1281, w1282, w1283, w1284, w1285, w1286, w1287, w1288, w1289, w1290, w1291, w1292, w1293, w1294, w1295, w1296, w1297, w1298, w1299, w1300, w1301, w1302, w1303, w1304, w1305, w1306, w1307, w1308, w1309, w1310, w1311, w1312, w1313, w1314, w1315, w1316, w1317, w1318, w1319, w1320, w1321, w1322, w1323, w1324, w1325, w1326, w1327, w1328, w1329, w1330, w1331, w1332, w1333, w1334, w1335, w1336, w1337, w1338, w1339, w1340, w1341, w1342, w1343, w1344, w1345, w1346, w1347, w1348, w1349, w1350, w1351, w1352, w1353, w1354, w1355, w1356, w1357, w1358, w1359, w1360, w1361, w1362, w1363, w1364, w1365, w1366, w1367, w1368, w1369, w1370, w1371, w1372, w1373, w1374, w1375, w1376, w1377, w1378, w1379, w1380, w1381, w1382, w1383, w1384, w1385, w1386, w1387, w1388, w1389, w1390, w1391, w1392, w1393, w1394, w1395, w1396, w1397, w1398, w1399, w1400, w1401, w1402, w1403, w1404, w1405, w1406, w1407, w1408, w1409, w1410, w1411, w1412, w1413, w1414, w1415, w1416, w1417, w1418, w1419, w1420, w1421, w1422, w1423, w1424, w1425, w1426, w1427, w1428, w1429, w1430, w1431, w1432, w1433, w1434, w1435, w1436, w1437, w1438, w1439, w1440, w1441, w1442, w1443, w1444, w1445, w1446, w1447, w1448, w1449, w1450, w1451, w1452, w1453, w1454, w1455, w1456, w1457, w1458, w1459, w1460, w1461, w1462, w1463, w1464, w1465, w1466, w1467, w1468, w1469, w1470, w1471, w1472, w1473, w1474, w1475, w1476, w1477, w1478, w1479, w1480, w1481, w1482, w1483, w1484, w1485, w1486, w1487, w1488, w1489, w1490, w1491, w1492, w1493, w1494, w1495, w1496, w1497, w1498, w1499, w1500, w1501, w1502, w1503, w1504, w1505, w1506, w1507, w1508, w1509, w1510, w1511, w1512, w1513, w1514, w1515, w1516, w1517, w1518, w1519, w1520, w1521, w1522, w1523, w1524, w1525, w1526, w1527, w1528, w1529, w1530, w1531, w1532, w1533, w1534, w1535, w1536, w1537, w1538, w1539, w1540, w1541, w1542, w1543, w1544, w1545, w1546, w1547, w1548, w1549, w1550, w1551, w1552, w1553, w1554, w1555, w1556, w1557, w1558, w1559, w1560, w1561, w1562, w1563, w1564, w1565, w1566, w1567, w1568, w1569, w1570, w1571, w1572, w1573, w1574, w1575, w1576, w1577, w1578, w1579, w1580, w1581, w1582, w1583, w1584, w1585, w1586, w1587, w1588, w1589, w1590, w1591, w1592, w1593, w1594, w1595, w1596, w1597, w1598, w1599, w1600, w1601, w1602, w1603, w1604, w1605, w1606, w1607, w1608, w1609, w1610, w1611, w1612, w1613, w1614, w1615, w1616, w1617, w1618, w1619, w1620, w1621, w1622, w1623, w1624, w1625, w1626, w1627, w1628, w1629, w1630, w1631, w1632, w1633, w1634, w1635, w1636, w1637, w1638, w1639, w1640, w1641, w1642, w1643, w1644, w1645, w1646, w1647, w1648, w1649, w1650, w1651, w1652, w1653, w1654, w1655, w1656, w1657, w1658, w1659, w1660, w1661, w1662, w1663, w1664, w1665, w1666, w1667, w1668, w1669, w1670, w1671, w1672, w1673, w1674, w1675, w1676, w1677, w1678, w1679, w1680, w1681, w1682, w1683, w1684, w1685, w1686, w1687, w1688, w1689, w1690, w1691, w1692, w1693, w1694, w1695, w1696, w1697, w1698, w1699, w1700, w1701, w1702, w1703, w1704, w1705, w1706, w1707, w1708, w1709, w1710, w1711, w1712, w1713, w1714, w1715, w1716, w1717, w1718, w1719, w1720, w1721, w1722, w1723, w1724, w1725, w1726, w1727, w1728, w1729, w1730, w1731, w1732, w1733, w1734, w1735, w1736, w1737, w1738, w1739, w1740, w1741, w1742, w1743, w1744, w1745, w1746, w1747, w1748, w1749, w1750, w1751, w1752, w1753, w1754, w1755, w1756, w1757, w1758, w1759, w1760, w1761, w1762, w1763, w1764, w1765, w1766, w1767, w1768, w1769, w1770, w1771, w1772, w1773, w1774, w1775, w1776, w1777, w1778, w1779, w1780, w1781, w1782, w1783, w1784, w1785, w1786, w1787, w1788, w1789, w1790, w1791, w1792, w1793, w1794, w1795, w1796, w1797, w1798, w1799, w1800, w1801, w1802, w1803, w1804, w1805, w1806, w1807, w1808, w1809, w1810, w1811, w1812, w1813, w1814, w1815, w1816, w1817, w1818, w1819, w1820, w1821, w1822, w1823, w1824, w1825, w1826, w1827, w1828, w1829, w1830, w1831, w1832, w1833, w1834, w1835, w1836, w1837, w1838, w1839, w1840, w1841, w1842, w1843, w1844, w1845, w1846, w1847, w1848, w1849, w1850, w1851, w1852, w1853, w1854, w1855, w1856, w1857, w1858, w1859, w1860, w1861, w1862, w1863, w1864, w1865, w1866, w1867, w1868, w1869, w1870, w1871, w1872, w1873, w1874, w1875, w1876, w1877, w1878, w1879, w1880, w1881, w1882, w1883, w1884, w1885, w1886, w1887, w1888, w1889, w1890, w1891, w1892, w1893, w1894, w1895, w1896, w1897, w1898, w1899, w1900, w1901, w1902, w1903, w1904, w1905, w1906, w1907, w1908, w1909, w1910, w1911, w1912, w1913, w1914, w1915, w1916, w1917, w1918, w1919, w1920, w1921, w1922, w1923, w1924, w1925, w1926, w1927, w1928, w1929, w1930, w1931, w1932, w1933, w1934, w1935, w1936, w1937, w1938, w1939, w1940, w1941, w1942, w1943, w1944, w1945, w1946, w1947, w1948, w1949, w1950, w1951, w1952, w1953, w1954, w1955, w1956, w1957, w1958, w1959, w1960, w1961, w1962, w1963, w1964, w1965, w1966, w1967, w1968, w1969, w1970, w1971, w1972, w1973, w1974, w1975, w1976, w1977, w1978, w1979, w1980, w1981, w1982, w1983, w1984, w1985, w1986, w1987, w1988, w1989, w1990, w1991, w1992, w1993, w1994, w1995, w1996, w1997, w1998, w1999, w2000, w2001, w2002, w2003, w2004, w2005, w2006, w2007, w2008, w2009, w2010, w2011, w2012, w2013, w2014, w2015, w2016, w2017, w2018, w2019, w2020, w2021, w2022, w2023, w2024, w2025, w2026, w2027, w2028, w2029, w2030, w2031, w2032, w2033, w2034, w2035, w2036, w2037, w2038, w2039, w2040, w2041, w2042, w2043, w2044, w2045, w2046, w2047, w2048, w2049, w2050, w2051, w2052, w2053, w2054, w2055, w2056, w2057, w2058, w2059, w2060, w2061, w2062, w2063, w2064, w2065, w2066, w2067, w2068, w2069, w2070, w2071, w2072, w2073, w2074, w2075, w2076, w2077, w2078, w2079, w2080, w2081, w2082, w2083, w2084, w2085, w2086, w2087, w2088, w2089, w2090, w2091, w2092, w2093, w2094, w2095, w2096, w2097, w2098, w2099, w2100, w2101, w2102, w2103, w2104, w2105, w2106, w2107, w2108, w2109, w2110, w2111, w2112, w2113, w2114, w2115, w2116, w2117, w2118, w2119, w2120, w2121, w2122, w2123, w2124, w2125, w2126, w2127, w2128, w2129, w2130, w2131, w2132, w2133, w2134, w2135, w2136, w2137, w2138, w2139, w2140, w2141, w2142, w2143, w2144, w2145, w2146, w2147, w2148, w2149, w2150, w2151, w2152, w2153, w2154, w2155, w2156, w2157, w2158, w2159, w2160, w2161, w2162, w2163, w2164, w2165, w2166, w2167, w2168, w2169, w2170, w2171, w2172, w2173, w2174, w2175, w2176, w2177, w2178, w2179, w2180, w2181, w2182, w2183, w2184, w2185, w2186, w2187, w2188, w2189, w2190, w2191, w2192, w2193, w2194, w2195, w2196, w2197, w2198, w2199, w2200, w2201, w2202, w2203, w2204, w2205, w2206, w2207, w2208, w2209, w2210, w2211, w2212, w2213, w2214, w2215, w2216, w2217, w2218, w2219, w2220, w2221, w2222, w2223, w2224, w2225, w2226, w2227, w2228, w2229, w2230, w2231, w2232, w2233, w2234, w2235, w2236, w2237, w2238, w2239, w2240, w2241, w2242, w2243, w2244, w2245, w2246, w2247, w2248, w2249, w2250, w2251, w2252, w2253, w2254, w2255, w2256, w2257, w2258, w2259, w2260, w2261, w2262, w2263, w2264, w2265, w2266, w2267, w2268, w2269, w2270, w2271, w2272, w2273, w2274, w2275, w2276, w2277, w2278, w2279, w2280, w2281, w2282, w2283, w2284, w2285, w2286, w2287, w2288, w2289, w2290, w2291, w2292, w2293, w2294, w2295, w2296, w2297, w2298, w2299, w2300, w2301, w2302, w2303, w2304, w2305, w2306, w2307, w2308, w2309, w2310, w2311, w2312, w2313, w2314, w2315, w2316, w2317, w2318, w2319, w2320, w2321, w2322, w2323, w2324, w2325, w2326, w2327, w2328, w2329, w2330, w2331, w2332, w2333, w2334, w2335, w2336, w2337, w2338, w2339, w2340, w2341, w2342, w2343, w2344, w2345, w2346, w2347, w2348, w2349, w2350, w2351, w2352, w2353, w2354, w2355, w2356, w2357, w2358, w2359, w2360, w2361, w2362, w2363, w2364, w2365, w2366, w2367, w2368, w2369, w2370, w2371, w2372, w2373, w2374, w2375, w2376, w2377, w2378, w2379, w2380, w2381, w2382, w2383, w2384, w2385, w2386, w2387, w2388, w2389, w2390, w2391, w2392, w2393, w2394, w2395, w2396, w2397, w2398, w2399, w2400, w2401, w2402, w2403, w2404, w2405, w2406, w2407, w2408, w2409, w2410, w2411, w2412, w2413, w2414, w2415, w2416, w2417, w2418, w2419, w2420, w2421, w2422, w2423, w2424, w2425, w2426, w2427, w2428, w2429, w2430, w2431, w2432, w2433, w2434, w2435, w2436, w2437, w2438, w2439, w2440, w2441, w2442, w2443, w2444, w2445, w2446, w2447, w2448, w2449, w2450, w2451, w2452, w2453, w2454, w2455, w2456, w2457, w2458, w2459, w2460, w2461, w2462, w2463, w2464, w2465, w2466, w2467, w2468, w2469, w2470, w2471, w2472, w2473, w2474, w2475, w2476, w2477, w2478, w2479, w2480, w2481, w2482, w2483, w2484, w2485, w2486, w2487, w2488, w2489, w2490, w2491, w2492, w2493, w2494, w2495, w2496, w2497, w2498, w2499, w2500, w2501, w2502, w2503, w2504, w2505, w2506, w2507, w2508, w2509, w2510, w2511, w2512, w2513, w2514, w2515, w2516, w2517, w2518, w2519, w2520, w2521, w2522, w2523, w2524, w2525, w2526, w2527, w2528, w2529, w2530, w2531, w2532, w2533, w2534, w2535, w2536, w2537, w2538, w2539, w2540, w2541, w2542, w2543, w2544, w2545, w2546, w2547, w2548, w2549, w2550, w2551, w2552, w2553, w2554, w2555, w2556, w2557, w2558, w2559, w2560, w2561, w2562, w2563, w2564, w2565, w2566, w2567, w2568, w2569, w2570, w2571, w2572, w2573, w2574, w2575, w2576, w2577, w2578, w2579, w2580, w2581, w2582, w2583, w2584, w2585, w2586, w2587, w2588, w2589, w2590, w2591, w2592, w2593, w2594, w2595, w2596, w2597, w2598, w2599, w2600, w2601, w2602, w2603, w2604, w2605, w2606, w2607, w2608, w2609, w2610, w2611, w2612, w2613, w2614, w2615, w2616, w2617, w2618, w2619, w2620, w2621, w2622, w2623, w2624, w2625, w2626, w2627, w2628, w2629, w2630, w2631, w2632, w2633, w2634, w2635, w2636, w2637, w2638, w2639, w2640, w2641, w2642, w2643, w2644, w2645, w2646, w2647, w2648, w2649, w2650, w2651, w2652, w2653, w2654, w2655, w2656, w2657, w2658, w2659, w2660, w2661, w2662, w2663, w2664, w2665, w2666, w2667, w2668, w2669, w2670, w2671, w2672, w2673, w2674, w2675, w2676, w2677, w2678, w2679, w2680, w2681, w2682, w2683, w2684, w2685, w2686, w2687, w2688, w2689, w2690, w2691, w2692, w2693, w2694, w2695, w2696, w2697, w2698, w2699, w2700, w2701, w2702, w2703, w2704, w2705, w2706, w2707, w2708, w2709, w2710, w2711, w2712, w2713, w2714, w2715, w2716, w2717, w2718, w2719, w2720, w2721, w2722, w2723, w2724, w2725, w2726, w2727, w2728, w2729, w2730, w2731, w2732, w2733, w2734, w2735, w2736, w2737, w2738, w2739, w2740, w2741, w2742, w2743, w2744, w2745, w2746, w2747, w2748, w2749, w2750, w2751, w2752, w2753, w2754, w2755, w2756, w2757, w2758, w2759, w2760, w2761, w2762, w2763, w2764, w2765, w2766, w2767, w2768, w2769, w2770, w2771, w2772, w2773, w2774, w2775, w2776, w2777, w2778, w2779, w2780, w2781, w2782, w2783, w2784, w2785, w2786, w2787, w2788, w2789, w2790, w2791, w2792, w2793, w2794, w2795, w2796, w2797, w2798, w2799, w2800, w2801, w2802, w2803, w2804, w2805, w2806, w2807, w2808, w2809, w2810, w2811, w2812, w2813, w2814, w2815, w2816, w2817, w2818, w2819, w2820, w2821, w2822, w2823, w2824, w2825, w2826, w2827, w2828, w2829, w2830, w2831, w2832, w2833, w2834, w2835, w2836, w2837, w2838, w2839, w2840, w2841, w2842, w2843, w2844, w2845, w2846, w2847, w2848, w2849, w2850, w2851, w2852, w2853, w2854, w2855, w2856, w2857, w2858, w2859, w2860, w2861, w2862, w2863, w2864, w2865, w2866, w2867, w2868, w2869, w2870, w2871, w2872, w2873, w2874, w2875, w2876, w2877, w2878, w2879, w2880, w2881, w2882, w2883, w2884, w2885, w2886, w2887, w2888, w2889, w2890, w2891, w2892, w2893, w2894, w2895, w2896, w2897, w2898, w2899, w2900, w2901, w2902, w2903, w2904, w2905, w2906, w2907, w2908, w2909, w2910, w2911, w2912, w2913, w2914, w2915, w2916, w2917, w2918, w2919, w2920, w2921, w2922, w2923, w2924, w2925, w2926, w2927, w2928, w2929, w2930, w2931, w2932, w2933, w2934, w2935, w2936, w2937, w2938, w2939, w2940, w2941, w2942, w2943, w2944, w2945, w2946, w2947, w2948, w2949, w2950, w2951, w2952, w2953, w2954, w2955, w2956, w2957, w2958, w2959, w2960, w2961, w2962, w2963, w2964, w2965, w2966, w2967, w2968, w2969, w2970, w2971, w2972, w2973, w2974, w2975, w2976, w2977, w2978, w2979, w2980, w2981, w2982, w2983, w2984, w2985, w2986, w2987, w2988, w2989, w2990, w2991, w2992, w2993, w2994, w2995, w2996, w2997, w2998, w2999, w3000, w3001, w3002, w3003, w3004, w3005, w3006, w3007, w3008, w3009, w3010, w3011, w3012, w3013, w3014, w3015, w3016, w3017, w3018, w3019, w3020, w3021, w3022, w3023, w3024, w3025, w3026, w3027, w3028, w3029, w3030, w3031, w3032, w3033, w3034, w3035, w3036, w3037, w3038, w3039, w3040, w3041, w3042, w3043, w3044, w3045, w3046, w3047, w3048, w3049, w3050, w3051, w3052, w3053, w3054, w3055, w3056, w3057, w3058, w3059, w3060, w3061, w3062, w3063, w3064, w3065, w3066, w3067, w3068, w3069, w3070, w3071, w3072, w3073, w3074, w3075, w3076, w3077, w3078, w3079, w3080, w3081, w3082, w3083, w3084, w3085, w3086, w3087, w3088, w3089, w3090, w3091, w3092, w3093, w3094, w3095, w3096, w3097, w3098, w3099, w3100, w3101, w3102, w3103, w3104, w3105, w3106, w3107, w3108, w3109, w3110, w3111, w3112, w3113, w3114, w3115, w3116, w3117, w3118, w3119, w3120, w3121, w3122, w3123, w3124, w3125, w3126, w3127, w3128, w3129, w3130, w3131, w3132, w3133, w3134, w3135, w3136, w3137, w3138, w3139, w3140, w3141, w3142, w3143, w3144, w3145, w3146, w3147, w3148, w3149, w3150, w3151, w3152, w3153, w3154, w3155, w3156, w3157, w3158, w3159, w3160, w3161, w3162, w3163, w3164, w3165, w3166, w3167, w3168, w3169, w3170, w3171, w3172, w3173, w3174, w3175, w3176, w3177, w3178, w3179, w3180, w3181, w3182, w3183, w3184, w3185, w3186, w3187, w3188, w3189, w3190, w3191, w3192, w3193, w3194, w3195, w3196, w3197, w3198, w3199, w3200, w3201, w3202, w3203, w3204, w3205, w3206, w3207, w3208, w3209, w3210, w3211, w3212, w3213, w3214, w3215, w3216, w3217, w3218, w3219, w3220, w3221, w3222, w3223, w3224, w3225, w3226, w3227, w3228, w3229, w3230, w3231, w3232, w3233, w3234, w3235, w3236, w3237, w3238, w3239, w3240, w3241, w3242, w3243, w3244, w3245, w3246, w3247, w3248, w3249, w3250, w3251, w3252, w3253, w3254, w3255, w3256, w3257, w3258, w3259, w3260, w3261, w3262, w3263, w3264, w3265, w3266, w3267, w3268, w3269, w3270, w3271, w3272, w3273, w3274, w3275, w3276, w3277, w3278, w3279, w3280, w3281, w3282, w3283, w3284, w3285, w3286, w3287, w3288, w3289, w3290, w3291, w3292, w3293, w3294, w3295, w3296, w3297, w3298, w3299, w3300, w3301, w3302, w3303, w3304, w3305, w3306, w3307, w3308, w3309, w3310, w3311, w3312, w3313, w3314, w3315, w3316, w3317, w3318, w3319, w3320, w3321, w3322, w3323, w3324, w3325, w3326, w3327, w3328, w3329, w3330, w3331, w3332, w3333, w3334, w3335, w3336;
assign w0 = ~pi136 & ~pi152;
assign w1 = ~pi196 & ~w0;
assign w2 = ~pi194 & ~w0;
assign w3 = ~pi197 & ~w0;
assign w4 = ~pi193 & ~w0;
assign w5 = ~pi198 & ~w0;
assign w6 = ~pi192 & ~w0;
assign w7 = ~pi199 & ~w0;
assign w8 = ~pi195 & ~w0;
assign w9 = pi187 & pi190;
assign w10 = pi138 & pi148;
assign w11 = w9 & w10;
assign w12 = pi138 & pi190;
assign w13 = (~pi148 & ~w12) | (~pi148 & w2860) | (~w12 & w2860);
assign w14 = ~w11 & ~w13;
assign w15 = pi156 & ~w14;
assign w16 = pi142 & ~pi176;
assign w17 = ~w11 & w16;
assign w18 = ~pi142 & ~pi176;
assign w19 = w11 & w18;
assign w20 = ~w17 & ~w19;
assign w21 = w15 & w20;
assign w22 = pi171 & ~pi187;
assign w23 = ~w12 & w22;
assign w24 = pi171 & pi187;
assign w25 = w12 & w24;
assign w26 = ~w23 & ~w25;
assign w27 = ~pi138 & ~pi190;
assign w28 = ~w12 & ~w27;
assign w29 = ~pi150 & w28;
assign w30 = ~pi171 & ~pi187;
assign w31 = w12 & ~w30;
assign w32 = ~pi171 & pi187;
assign w33 = ~w12 & ~w32;
assign w34 = ~w31 & ~w33;
assign w35 = ~w29 & ~w34;
assign w36 = w26 & ~w35;
assign w37 = ~pi156 & ~w11;
assign w38 = ~w13 & w37;
assign w39 = w20 & ~w38;
assign w40 = ~w36 & w39;
assign w41 = ~w21 & ~w40;
assign w42 = ~pi142 & pi176;
assign w43 = ~w16 & ~w42;
assign w44 = w11 & w43;
assign w45 = ~w11 & ~w43;
assign w46 = ~w44 & ~w45;
assign w47 = pi176 & ~w46;
assign w48 = ~w40 & w2861;
assign w49 = pi142 & w11;
assign w50 = ~pi139 & pi177;
assign w51 = pi139 & ~pi177;
assign w52 = ~w50 & ~w51;
assign w53 = w49 & ~w52;
assign w54 = ~w49 & w52;
assign w55 = ~w53 & ~w54;
assign w56 = ~w48 & w55;
assign w57 = ~w47 & ~w55;
assign w58 = (pi143 & ~w41) | (pi143 & w2862) | (~w41 & w2862);
assign w59 = ~w56 & w58;
assign w60 = pi138 & pi139;
assign w61 = ~pi187 & ~pi190;
assign w62 = ~pi148 & w61;
assign w63 = w61 & w2863;
assign w64 = ~pi139 & w63;
assign w65 = pi139 & ~w63;
assign w66 = ~w64 & ~w65;
assign w67 = ~pi138 & ~w66;
assign w68 = ~pi143 & ~w60;
assign w69 = ~w67 & w68;
assign w70 = ~w59 & ~w69;
assign w71 = ~w14 & w2921;
assign w72 = (pi143 & ~w37) | (pi143 & w2864) | (~w37 & w2864);
assign w73 = ~w36 & w72;
assign w74 = (~w71 & w36) | (~w71 & w2922) | (w36 & w2922);
assign w75 = pi143 & ~w46;
assign w76 = (w75 & w73) | (w75 & w2865) | (w73 & w2865);
assign w77 = w61 & w3237;
assign w78 = pi142 & ~w77;
assign w79 = ~pi143 & ~w63;
assign w80 = (~pi143 & ~w61) | (~pi143 & w2866) | (~w61 & w2866);
assign w81 = ~w79 & ~w80;
assign w82 = ~w78 & ~w81;
assign w83 = ~w75 & ~w82;
assign w84 = w74 & w83;
assign w85 = ~w76 & ~w84;
assign w86 = (w85 & w59) | (w85 & w2923) | (w59 & w2923);
assign w87 = w11 & w2867;
assign w88 = w11 & w3238;
assign w89 = (~pi140 & ~w11) | (~pi140 & w3239) | (~w11 & w3239);
assign w90 = ~w88 & ~w89;
assign w91 = pi161 & ~w90;
assign w92 = ~pi161 & w90;
assign w93 = ~w91 & ~w92;
assign w94 = ~pi139 & ~w49;
assign w95 = ~pi177 & ~w87;
assign w96 = ~w94 & w95;
assign w97 = (~w96 & ~w41) | (~w96 & w2868) | (~w41 & w2868);
assign w98 = w97 & w3240;
assign w99 = pi143 & ~w93;
assign w100 = pi138 & pi140;
assign w101 = w63 & w3241;
assign w102 = pi140 & ~w64;
assign w103 = ~w101 & ~w102;
assign w104 = ~pi138 & ~w103;
assign w105 = ~pi143 & ~w100;
assign w106 = ~w104 & w105;
assign w107 = (~w106 & w97) | (~w106 & w3242) | (w97 & w3242);
assign w108 = ~w98 & w107;
assign w109 = (~w91 & ~w97) | (~w91 & w2924) | (~w97 & w2924);
assign w110 = pi133 & ~pi178;
assign w111 = ~pi133 & pi178;
assign w112 = ~w110 & ~w111;
assign w113 = w88 & w112;
assign w114 = ~w88 & ~w112;
assign w115 = ~w113 & ~w114;
assign w116 = pi143 & ~w115;
assign w117 = pi133 & pi138;
assign w118 = pi133 & ~w101;
assign w119 = ~pi133 & w101;
assign w120 = ~w118 & ~w119;
assign w121 = ~pi138 & ~w120;
assign w122 = ~pi143 & ~w117;
assign w123 = ~w121 & w122;
assign w124 = ~w116 & ~w123;
assign w125 = w109 & ~w124;
assign w126 = pi143 & w115;
assign w127 = ~w123 & ~w126;
assign w128 = ~w109 & ~w127;
assign w129 = ~w125 & ~w128;
assign w130 = w108 & ~w129;
assign w131 = w86 & w130;
assign w132 = pi143 & ~pi150;
assign w133 = w28 & w132;
assign w134 = ~w28 & ~w132;
assign w135 = ~w133 & ~w134;
assign w136 = pi143 & w26;
assign w137 = w35 & w136;
assign w138 = pi187 & ~w27;
assign w139 = w80 & ~w138;
assign w140 = ~w22 & ~w32;
assign w141 = w133 & ~w140;
assign w142 = ~w139 & ~w141;
assign w143 = ~w137 & w142;
assign w144 = ~w135 & w143;
assign w145 = ~w36 & w2869;
assign w146 = pi148 & ~w61;
assign w147 = ~pi143 & ~w146;
assign w148 = ~w10 & ~w77;
assign w149 = w147 & w148;
assign w150 = ~pi148 & pi156;
assign w151 = pi148 & ~pi156;
assign w152 = ~w150 & ~w151;
assign w153 = ~w35 & ~w152;
assign w154 = (~w149 & ~w153) | (~w149 & w3243) | (~w153 & w3243);
assign w155 = ~w145 & w154;
assign w156 = w144 & w155;
assign w157 = pi232 & pi233;
assign w158 = ~pi136 & pi231;
assign w159 = w157 & w158;
assign w160 = pi235 & pi236;
assign w161 = ~pi237 & w160;
assign w162 = w159 & w161;
assign w163 = w156 & ~w162;
assign w164 = w131 & w163;
assign w165 = ~pi000 & ~w164;
assign w166 = ~pi237 & w159;
assign w167 = ~w160 & w166;
assign w168 = ~w165 & ~w167;
assign w169 = pi235 & ~pi236;
assign w170 = ~pi237 & w169;
assign w171 = w159 & w170;
assign w172 = ~pi270 & w171;
assign w173 = ~pi235 & ~pi237;
assign w174 = w159 & w173;
assign w175 = ~w172 & ~w174;
assign w176 = pi000 & ~w175;
assign w177 = pi245 & pi270;
assign w178 = w171 & w177;
assign w179 = ~w176 & ~w178;
assign w180 = ~w168 & w179;
assign w181 = w85 & ~w155;
assign w182 = ~w135 & ~w143;
assign w183 = ~w143 & w2870;
assign w184 = ~w137 & ~w139;
assign w185 = (w135 & w137) | (w135 & w2871) | (w137 & w2871);
assign w186 = pi099 & w185;
assign w187 = w135 & ~w139;
assign w188 = ~w137 & w187;
assign w189 = pi111 & w188;
assign w190 = w143 & w2872;
assign w191 = ~w183 & ~w189;
assign w192 = ~w186 & ~w190;
assign w193 = w191 & w192;
assign w194 = w181 & ~w193;
assign w195 = w85 & w155;
assign w196 = pi113 & w185;
assign w197 = w143 & w2873;
assign w198 = ~w143 & w2874;
assign w199 = pi069 & w188;
assign w200 = ~w196 & ~w199;
assign w201 = ~w197 & ~w198;
assign w202 = w200 & w201;
assign w203 = w195 & ~w202;
assign w204 = ~w85 & ~w155;
assign w205 = ~w143 & w2875;
assign w206 = w143 & w2876;
assign w207 = pi080 & w188;
assign w208 = pi001 & w185;
assign w209 = ~w205 & ~w207;
assign w210 = ~w206 & ~w208;
assign w211 = w209 & w210;
assign w212 = w204 & ~w211;
assign w213 = ~w85 & w155;
assign w214 = pi098 & w185;
assign w215 = ~w143 & w3244;
assign w216 = pi083 & w188;
assign w217 = w143 & w3245;
assign w218 = ~w214 & ~w216;
assign w219 = ~w215 & ~w217;
assign w220 = w218 & w219;
assign w221 = w213 & ~w220;
assign w222 = w70 & ~w194;
assign w223 = ~w203 & ~w212;
assign w224 = ~w221 & w223;
assign w225 = w108 & w222;
assign w226 = w224 & w225;
assign w227 = ~w70 & ~w108;
assign w228 = ~w143 & w3246;
assign w229 = w143 & w3247;
assign w230 = pi101 & w185;
assign w231 = pi109 & w188;
assign w232 = ~w228 & ~w231;
assign w233 = ~w229 & ~w230;
assign w234 = w232 & w233;
assign w235 = w204 & ~w234;
assign w236 = pi074 & w185;
assign w237 = ~w143 & w2877;
assign w238 = w143 & w2878;
assign w239 = pi107 & w188;
assign w240 = ~w236 & ~w239;
assign w241 = ~w237 & ~w238;
assign w242 = w240 & w241;
assign w243 = w195 & ~w242;
assign w244 = pi003 & w185;
assign w245 = w143 & w2879;
assign w246 = pi072 & w188;
assign w247 = ~w143 & w2880;
assign w248 = ~w244 & ~w246;
assign w249 = ~w245 & ~w247;
assign w250 = w248 & w249;
assign w251 = w181 & ~w250;
assign w252 = w143 & w3248;
assign w253 = ~w143 & w3249;
assign w254 = pi077 & w188;
assign w255 = pi112 & w185;
assign w256 = ~w252 & ~w254;
assign w257 = ~w253 & ~w255;
assign w258 = w256 & w257;
assign w259 = w213 & ~w258;
assign w260 = ~w70 & ~w235;
assign w261 = ~w243 & ~w251;
assign w262 = ~w259 & w261;
assign w263 = w260 & w262;
assign w264 = pi051 & w185;
assign w265 = w143 & w2881;
assign w266 = ~w143 & w2882;
assign w267 = pi049 & w188;
assign w268 = ~w264 & ~w267;
assign w269 = ~w265 & ~w266;
assign w270 = w268 & w269;
assign w271 = w204 & ~w270;
assign w272 = w143 & w2883;
assign w273 = ~w143 & w2884;
assign w274 = pi027 & w188;
assign w275 = pi025 & w185;
assign w276 = ~w272 & ~w274;
assign w277 = ~w273 & ~w275;
assign w278 = w276 & w277;
assign w279 = w181 & ~w278;
assign w280 = pi029 & w185;
assign w281 = w143 & w2885;
assign w282 = pi067 & w188;
assign w283 = ~w143 & w2886;
assign w284 = ~w280 & ~w282;
assign w285 = ~w281 & ~w283;
assign w286 = w284 & w285;
assign w287 = w195 & ~w286;
assign w288 = pi053 & w185;
assign w289 = w143 & w2887;
assign w290 = ~w143 & w2888;
assign w291 = pi054 & w188;
assign w292 = ~w288 & ~w291;
assign w293 = ~w289 & ~w290;
assign w294 = w292 & w293;
assign w295 = w213 & ~w294;
assign w296 = ~w271 & ~w279;
assign w297 = ~w287 & ~w295;
assign w298 = w296 & w297;
assign w299 = ~w108 & w298;
assign w300 = ~w226 & ~w227;
assign w301 = ~w263 & ~w299;
assign w302 = w300 & w301;
assign w303 = ~w143 & w3250;
assign w304 = w143 & w3251;
assign w305 = pi018 & w185;
assign w306 = pi019 & w188;
assign w307 = ~w303 & ~w306;
assign w308 = ~w304 & ~w305;
assign w309 = w307 & w308;
assign w310 = w181 & ~w309;
assign w311 = w143 & w3252;
assign w312 = pi022 & w185;
assign w313 = pi056 & w188;
assign w314 = ~w143 & w3253;
assign w315 = ~w311 & ~w313;
assign w316 = ~w312 & ~w314;
assign w317 = w315 & w316;
assign w318 = w204 & ~w317;
assign w319 = w143 & w3254;
assign w320 = ~w143 & w3255;
assign w321 = pi023 & w188;
assign w322 = pi061 & w185;
assign w323 = ~w319 & ~w321;
assign w324 = ~w320 & ~w322;
assign w325 = w323 & w324;
assign w326 = w213 & ~w325;
assign w327 = w143 & w3256;
assign w328 = ~w143 & w3257;
assign w329 = pi020 & w185;
assign w330 = pi060 & w188;
assign w331 = ~w327 & ~w330;
assign w332 = ~w328 & ~w329;
assign w333 = w331 & w332;
assign w334 = w195 & ~w333;
assign w335 = ~w310 & ~w318;
assign w336 = ~w326 & ~w334;
assign w337 = w335 & w336;
assign w338 = w227 & ~w337;
assign w339 = ~w129 & ~w338;
assign w340 = ~w302 & w339;
assign w341 = ~w108 & w129;
assign w342 = pi138 & pi146;
assign w343 = ~pi138 & ~pi145;
assign w344 = ~pi130 & w119;
assign w345 = ~pi129 & w344;
assign w346 = ~w342 & ~w343;
assign w347 = ~w345 & w346;
assign w348 = ~w341 & ~w347;
assign w349 = (~w69 & w84) | (~w69 & w2889) | (w84 & w2889);
assign w350 = ~w59 & w349;
assign w351 = w143 & w2890;
assign w352 = ~pi015 & ~w135;
assign w353 = ~w143 & w352;
assign w354 = ~pi016 & w188;
assign w355 = ~pi031 & w185;
assign w356 = ~w353 & ~w354;
assign w357 = w155 & w356;
assign w358 = ~w351 & ~w355;
assign w359 = w357 & w358;
assign w360 = ~w143 & w2891;
assign w361 = ~pi046 & w188;
assign w362 = ~pi044 & w135;
assign w363 = ~w184 & w362;
assign w364 = w143 & w2892;
assign w365 = ~w361 & ~w363;
assign w366 = ~w155 & w365;
assign w367 = ~w360 & ~w364;
assign w368 = w366 & w367;
assign w369 = ~w359 & ~w368;
assign w370 = ~w59 & w2925;
assign w371 = ~pi040 & w185;
assign w372 = w143 & w2893;
assign w373 = ~pi045 & w188;
assign w374 = ~w143 & w2926;
assign w375 = ~w155 & ~w373;
assign w376 = ~w371 & ~w372;
assign w377 = ~w374 & w376;
assign w378 = w375 & w377;
assign w379 = ~w143 & w2894;
assign w380 = w143 & w2895;
assign w381 = ~pi012 & w188;
assign w382 = ~pi042 & w185;
assign w383 = w155 & ~w381;
assign w384 = ~w379 & ~w380;
assign w385 = ~w382 & w384;
assign w386 = w383 & w385;
assign w387 = ~w378 & ~w386;
assign w388 = w370 & w387;
assign w389 = (~w85 & w59) | (~w85 & w2927) | (w59 & w2927);
assign w390 = w143 & w2896;
assign w391 = ~pi010 & w185;
assign w392 = ~pi048 & w188;
assign w393 = ~w143 & w2928;
assign w394 = w155 & ~w392;
assign w395 = ~w390 & ~w391;
assign w396 = ~w393 & w395;
assign w397 = w394 & w396;
assign w398 = w143 & w2897;
assign w399 = ~w143 & w2898;
assign w400 = ~pi008 & w188;
assign w401 = ~pi037 & w185;
assign w402 = ~w155 & ~w400;
assign w403 = ~w398 & ~w399;
assign w404 = ~w401 & w403;
assign w405 = w402 & w404;
assign w406 = ~w397 & ~w405;
assign w407 = w389 & w406;
assign w408 = w143 & w2899;
assign w409 = pi033 & w185;
assign w410 = pi005 & w188;
assign w411 = ~w143 & w2929;
assign w412 = ~w155 & ~w410;
assign w413 = ~w408 & ~w409;
assign w414 = ~w411 & w413;
assign w415 = w412 & w414;
assign w416 = w143 & w2900;
assign w417 = ~w143 & w2901;
assign w418 = pi036 & w188;
assign w419 = pi006 & w185;
assign w420 = w155 & ~w418;
assign w421 = ~w416 & ~w417;
assign w422 = ~w419 & w421;
assign w423 = w420 & w422;
assign w424 = ~w415 & ~w423;
assign w425 = w86 & ~w424;
assign w426 = (~w347 & ~w369) | (~w347 & w2902) | (~w369 & w2902);
assign w427 = ~w388 & w426;
assign w428 = ~w407 & ~w425;
assign w429 = w427 & w428;
assign w430 = ~w348 & ~w429;
assign w431 = w108 & w129;
assign w432 = ~w143 & w2903;
assign w433 = w143 & w2904;
assign w434 = ~pi095 & w185;
assign w435 = ~pi092 & w188;
assign w436 = w155 & ~w435;
assign w437 = ~w432 & ~w433;
assign w438 = ~w434 & w437;
assign w439 = w436 & w438;
assign w440 = w143 & w2930;
assign w441 = ~pi102 & w185;
assign w442 = ~pi093 & w188;
assign w443 = ~pi088 & w182;
assign w444 = ~w155 & ~w442;
assign w445 = ~w440 & ~w441;
assign w446 = ~w443 & w445;
assign w447 = w444 & w446;
assign w448 = w350 & ~w439;
assign w449 = ~w447 & w448;
assign w450 = w143 & w2905;
assign w451 = ~w143 & w2906;
assign w452 = pi126 & w188;
assign w453 = pi105 & w185;
assign w454 = w155 & ~w452;
assign w455 = ~w450 & ~w451;
assign w456 = ~w453 & w455;
assign w457 = w454 & w456;
assign w458 = ~w143 & w2907;
assign w459 = pi084 & w185;
assign w460 = pi117 & w188;
assign w461 = w143 & w2931;
assign w462 = ~w155 & ~w460;
assign w463 = ~w458 & ~w459;
assign w464 = ~w461 & w463;
assign w465 = w462 & w464;
assign w466 = ~w457 & ~w465;
assign w467 = w389 & ~w466;
assign w468 = ~w143 & w2908;
assign w469 = w143 & w2909;
assign w470 = ~pi120 & w188;
assign w471 = ~pi108 & w185;
assign w472 = w155 & ~w470;
assign w473 = ~w468 & ~w469;
assign w474 = ~w471 & w473;
assign w475 = w472 & w474;
assign w476 = ~w143 & w2910;
assign w477 = w143 & w2911;
assign w478 = ~pi097 & w188;
assign w479 = ~pi086 & w185;
assign w480 = ~w155 & ~w478;
assign w481 = ~w476 & ~w477;
assign w482 = ~w479 & w481;
assign w483 = w480 & w482;
assign w484 = ~w475 & ~w483;
assign w485 = w370 & w484;
assign w486 = ~w143 & w2912;
assign w487 = w143 & w2913;
assign w488 = ~pi123 & w188;
assign w489 = ~pi116 & w185;
assign w490 = w155 & ~w488;
assign w491 = ~w486 & ~w487;
assign w492 = ~w489 & w491;
assign w493 = w490 & w492;
assign w494 = ~w143 & w2914;
assign w495 = w143 & w2915;
assign w496 = ~pi096 & w188;
assign w497 = ~pi118 & w185;
assign w498 = ~w155 & ~w496;
assign w499 = ~w494 & ~w495;
assign w500 = ~w497 & w499;
assign w501 = w498 & w500;
assign w502 = ~w493 & ~w501;
assign w503 = w86 & w502;
assign w504 = ~w449 & ~w467;
assign w505 = ~w485 & ~w503;
assign w506 = w504 & w505;
assign w507 = w431 & ~w506;
assign w508 = ~w430 & ~w507;
assign w509 = pi234 & w347;
assign w510 = w164 & w179;
assign w511 = (w2916 & w2932) | (w2916 & w2933) | (w2932 & w2933);
assign w512 = ~w180 & ~w511;
assign w513 = w130 & w350;
assign w514 = ~w155 & w185;
assign w515 = ~w162 & w514;
assign w516 = w513 & w515;
assign w517 = ~pi001 & ~w516;
assign w518 = ~w167 & ~w517;
assign w519 = ~pi273 & w171;
assign w520 = ~w174 & ~w519;
assign w521 = pi001 & ~w520;
assign w522 = pi262 & pi273;
assign w523 = w171 & w522;
assign w524 = ~w521 & ~w523;
assign w525 = ~w518 & w524;
assign w526 = w516 & w524;
assign w527 = (w2916 & w2934) | (w2916 & w2935) | (w2934 & w2935);
assign w528 = ~w525 & ~w527;
assign w529 = ~pi236 & w166;
assign w530 = pi236 & w166;
assign w531 = w156 & ~w530;
assign w532 = w513 & w531;
assign w533 = ~pi002 & ~w532;
assign w534 = ~w529 & ~w533;
assign w535 = ~pi236 & w174;
assign w536 = ~w519 & ~w535;
assign w537 = pi002 & ~w536;
assign w538 = pi269 & pi273;
assign w539 = w171 & w538;
assign w540 = ~w537 & ~w539;
assign w541 = ~w534 & w540;
assign w542 = w532 & w540;
assign w543 = (w2916 & w2936) | (w2916 & w2937) | (w2936 & w2937);
assign w544 = ~w541 & ~w543;
assign w545 = w131 & w515;
assign w546 = ~pi003 & ~w545;
assign w547 = ~w167 & ~w546;
assign w548 = pi003 & ~w175;
assign w549 = pi238 & pi270;
assign w550 = w171 & w549;
assign w551 = ~w548 & ~w550;
assign w552 = ~w547 & w551;
assign w553 = w545 & w551;
assign w554 = (w2916 & w2938) | (w2916 & w2939) | (w2938 & w2939);
assign w555 = ~w552 & ~w554;
assign w556 = ~w155 & w182;
assign w557 = ~w162 & w556;
assign w558 = w86 & w341;
assign w559 = w557 & w558;
assign w560 = ~pi004 & ~w559;
assign w561 = ~w167 & ~w560;
assign w562 = pi239 & pi270;
assign w563 = pi236 & w174;
assign w564 = w562 & w563;
assign w565 = ~pi270 & w563;
assign w566 = ~w529 & ~w565;
assign w567 = pi004 & ~w566;
assign w568 = ~w564 & ~w567;
assign w569 = ~w561 & w568;
assign w570 = w559 & w568;
assign w571 = (w2916 & w2940) | (w2916 & w2941) | (w2940 & w2941);
assign w572 = ~w569 & ~w571;
assign w573 = w129 & w3258;
assign w574 = ~w70 & w573;
assign w575 = w181 & w188;
assign w576 = w574 & w575;
assign w577 = ~pi005 & ~w576;
assign w578 = ~w167 & ~w577;
assign w579 = pi005 & ~w566;
assign w580 = pi240 & pi270;
assign w581 = w563 & w580;
assign w582 = ~w579 & ~w581;
assign w583 = ~w578 & w582;
assign w584 = w576 & w582;
assign w585 = (w2916 & w2942) | (w2916 & w2943) | (w2942 & w2943);
assign w586 = ~w583 & ~w585;
assign w587 = w185 & w195;
assign w588 = w574 & w587;
assign w589 = ~pi006 & ~w588;
assign w590 = ~w167 & ~w589;
assign w591 = pi006 & ~w566;
assign w592 = pi242 & pi270;
assign w593 = w563 & w592;
assign w594 = ~w591 & ~w593;
assign w595 = ~w590 & w594;
assign w596 = w588 & w594;
assign w597 = (w2916 & w2944) | (w2916 & w2945) | (w2944 & w2945);
assign w598 = ~w595 & ~w597;
assign w599 = w163 & w558;
assign w600 = ~pi007 & ~w599;
assign w601 = ~w167 & ~w600;
assign w602 = w177 & w563;
assign w603 = pi007 & ~w566;
assign w604 = ~w602 & ~w603;
assign w605 = ~w601 & w604;
assign w606 = w599 & w604;
assign w607 = (w2916 & w2946) | (w2916 & w2947) | (w2946 & w2947);
assign w608 = ~w605 & ~w607;
assign w609 = ~w155 & w188;
assign w610 = w389 & w573;
assign w611 = w609 & w610;
assign w612 = ~pi008 & ~w611;
assign w613 = ~w167 & ~w612;
assign w614 = ~pi271 & w563;
assign w615 = ~w529 & ~w614;
assign w616 = pi008 & ~w615;
assign w617 = pi248 & pi271;
assign w618 = w563 & w617;
assign w619 = ~w616 & ~w618;
assign w620 = ~w613 & w619;
assign w621 = w611 & w619;
assign w622 = (w2916 & w2948) | (w2916 & w2949) | (w2948 & w2949);
assign w623 = ~w620 & ~w622;
assign w624 = w144 & ~w155;
assign w625 = w610 & w624;
assign w626 = ~pi009 & ~w625;
assign w627 = ~w167 & ~w626;
assign w628 = pi009 & ~w615;
assign w629 = pi249 & pi271;
assign w630 = w563 & w629;
assign w631 = ~w628 & ~w630;
assign w632 = ~w627 & w631;
assign w633 = w625 & w631;
assign w634 = (w2916 & w2950) | (w2916 & w2951) | (w2950 & w2951);
assign w635 = ~w632 & ~w634;
assign w636 = w155 & w185;
assign w637 = w610 & w636;
assign w638 = ~pi010 & ~w637;
assign w639 = ~w167 & ~w638;
assign w640 = pi010 & ~w615;
assign w641 = pi250 & pi271;
assign w642 = w563 & w641;
assign w643 = ~w640 & ~w642;
assign w644 = ~w639 & w643;
assign w645 = w637 & w643;
assign w646 = (w2916 & w2952) | (w2916 & w2953) | (w2952 & w2953);
assign w647 = ~w644 & ~w646;
assign w648 = w155 & w182;
assign w649 = ~w162 & w648;
assign w650 = w341 & w370;
assign w651 = w649 & w650;
assign w652 = ~pi011 & ~w651;
assign w653 = ~w167 & ~w652;
assign w654 = ~pi272 & w563;
assign w655 = ~w529 & ~w654;
assign w656 = pi011 & ~w655;
assign w657 = pi259 & pi272;
assign w658 = w563 & w657;
assign w659 = ~w656 & ~w658;
assign w660 = ~w653 & w659;
assign w661 = w651 & w659;
assign w662 = (w2916 & w2954) | (w2916 & w2955) | (w2954 & w2955);
assign w663 = ~w660 & ~w662;
assign w664 = w155 & w188;
assign w665 = w573 & w664;
assign w666 = w370 & w665;
assign w667 = ~pi012 & ~w666;
assign w668 = ~w167 & ~w667;
assign w669 = pi012 & ~w655;
assign w670 = pi272 & w563;
assign w671 = pi260 & w670;
assign w672 = ~w669 & ~w671;
assign w673 = ~w668 & w672;
assign w674 = w666 & w672;
assign w675 = (w2916 & w2956) | (w2916 & w2957) | (w2956 & w2957);
assign w676 = ~w673 & ~w675;
assign w677 = w163 & w650;
assign w678 = ~pi013 & ~w677;
assign w679 = ~w167 & ~w678;
assign w680 = pi013 & ~w655;
assign w681 = pi261 & pi272;
assign w682 = w563 & w681;
assign w683 = ~w680 & ~w682;
assign w684 = ~w679 & w683;
assign w685 = w677 & w683;
assign w686 = (w2916 & w2958) | (w2916 & w2959) | (w2958 & w2959);
assign w687 = ~w684 & ~w686;
assign w688 = ~pi273 & w563;
assign w689 = ~w529 & ~w688;
assign w690 = pi014 & ~w689;
assign w691 = pi265 & pi273;
assign w692 = w563 & w691;
assign w693 = ~w690 & ~w692;
assign w694 = w350 & w573;
assign w695 = w624 & w694;
assign w696 = w693 & w695;
assign w697 = (w2916 & w2960) | (w2916 & w2961) | (w2960 & w2961);
assign w698 = ~pi014 & ~w695;
assign w699 = ~w167 & ~w698;
assign w700 = w693 & ~w699;
assign w701 = ~w697 & ~w700;
assign w702 = pi015 & ~w689;
assign w703 = pi267 & pi273;
assign w704 = w563 & w703;
assign w705 = ~w702 & ~w704;
assign w706 = w648 & w694;
assign w707 = w705 & w706;
assign w708 = (w2916 & w2962) | (w2916 & w2963) | (w2962 & w2963);
assign w709 = ~pi015 & ~w706;
assign w710 = ~w167 & ~w709;
assign w711 = w705 & ~w710;
assign w712 = ~w708 & ~w711;
assign w713 = w350 & w665;
assign w714 = ~pi016 & ~w713;
assign w715 = ~w167 & ~w714;
assign w716 = pi016 & ~w689;
assign w717 = pi268 & pi273;
assign w718 = w563 & w717;
assign w719 = ~w716 & ~w718;
assign w720 = ~w715 & w719;
assign w721 = w713 & w719;
assign w722 = (w2916 & w2964) | (w2916 & w2965) | (w2964 & w2965);
assign w723 = ~w720 & ~w722;
assign w724 = w538 & w563;
assign w725 = pi017 & ~w689;
assign w726 = ~w724 & ~w725;
assign w727 = w156 & w694;
assign w728 = w726 & w727;
assign w729 = (w2916 & w2966) | (w2916 & w2967) | (w2966 & w2967);
assign w730 = ~pi017 & ~w727;
assign w731 = ~w167 & ~w730;
assign w732 = w726 & ~w731;
assign w733 = ~w729 & ~w732;
assign w734 = ~w108 & ~w129;
assign w735 = ~w129 & w3259;
assign w736 = ~w166 & w735;
assign w737 = w514 & w736;
assign w738 = pi018 & ~w737;
assign w739 = ~w535 & ~w738;
assign w740 = pi018 & ~pi270;
assign w741 = ~w549 & ~w740;
assign w742 = w535 & w741;
assign w743 = ~w739 & ~w742;
assign w744 = ~w171 & ~w563;
assign w745 = w735 & w744;
assign w746 = w515 & ~w742;
assign w747 = w745 & w746;
assign w748 = (~w2916 & w2968) | (~w2916 & w2969) | (w2968 & w2969);
assign w749 = ~w743 & ~w748;
assign w750 = w609 & w736;
assign w751 = pi019 & ~w750;
assign w752 = ~w535 & ~w751;
assign w753 = pi019 & ~pi270;
assign w754 = ~w580 & ~w753;
assign w755 = w535 & w754;
assign w756 = ~w752 & ~w755;
assign w757 = ~w162 & w745;
assign w758 = w609 & ~w755;
assign w759 = w757 & w758;
assign w760 = (~w2916 & w2970) | (~w2916 & w2971) | (w2970 & w2971);
assign w761 = ~w756 & ~w760;
assign w762 = w636 & w736;
assign w763 = pi020 & ~w762;
assign w764 = ~w535 & ~w763;
assign w765 = pi020 & ~pi270;
assign w766 = ~w592 & ~w765;
assign w767 = w535 & w766;
assign w768 = ~w764 & ~w767;
assign w769 = w636 & ~w767;
assign w770 = w757 & w769;
assign w771 = (~w2916 & w2972) | (~w2916 & w2973) | (w2972 & w2973);
assign w772 = ~w768 & ~w771;
assign w773 = w156 & ~w166;
assign w774 = w735 & w773;
assign w775 = (~w2916 & w2974) | (~w2916 & w2975) | (w2974 & w2975);
assign w776 = ~pi235 & pi270;
assign w777 = w529 & ~w776;
assign w778 = ~w529 & ~w774;
assign w779 = ~w777 & ~w778;
assign w780 = pi021 & ~w779;
assign w781 = w177 & w535;
assign w782 = ~w780 & ~w781;
assign w783 = ~w775 & w782;
assign w784 = ~w129 & w3260;
assign w785 = ~w166 & w514;
assign w786 = w784 & w785;
assign w787 = pi022 & ~w786;
assign w788 = ~w535 & ~w787;
assign w789 = pi022 & ~pi271;
assign w790 = pi246 & pi271;
assign w791 = ~w789 & ~w790;
assign w792 = w535 & w791;
assign w793 = ~w788 & ~w792;
assign w794 = w744 & w784;
assign w795 = w515 & ~w792;
assign w796 = w794 & w795;
assign w797 = (~w2916 & w2976) | (~w2916 & w2977) | (w2976 & w2977);
assign w798 = ~w793 & ~w797;
assign w799 = ~w166 & w664;
assign w800 = w784 & w799;
assign w801 = (~w2916 & w2978) | (~w2916 & w2979) | (w2978 & w2979);
assign w802 = pi271 & w535;
assign w803 = pi252 & w802;
assign w804 = pi023 & ~w802;
assign w805 = ~w800 & w804;
assign w806 = ~w803 & ~w805;
assign w807 = ~w801 & w806;
assign w808 = w773 & w784;
assign w809 = pi024 & ~w808;
assign w810 = ~w535 & ~w809;
assign w811 = pi024 & ~pi271;
assign w812 = pi253 & pi271;
assign w813 = ~w811 & ~w812;
assign w814 = w535 & w813;
assign w815 = ~w810 & ~w814;
assign w816 = w163 & ~w814;
assign w817 = w794 & w816;
assign w818 = (~w2916 & w2980) | (~w2916 & w2981) | (w2980 & w2981);
assign w819 = ~w815 & ~w818;
assign w820 = w370 & w734;
assign w821 = w785 & w820;
assign w822 = pi025 & ~w821;
assign w823 = ~w535 & ~w822;
assign w824 = pi025 & ~pi272;
assign w825 = pi254 & pi272;
assign w826 = ~w824 & ~w825;
assign w827 = w535 & w826;
assign w828 = ~w823 & ~w827;
assign w829 = w744 & w820;
assign w830 = w515 & ~w827;
assign w831 = w829 & w830;
assign w832 = (~w2916 & w2982) | (~w2916 & w2983) | (w2982 & w2983);
assign w833 = ~w828 & ~w832;
assign w834 = ~w166 & w556;
assign w835 = w820 & w834;
assign w836 = (~w2916 & w2984) | (~w2916 & w2985) | (w2984 & w2985);
assign w837 = pi272 & w535;
assign w838 = ~pi255 & w837;
assign w839 = pi026 & ~w835;
assign w840 = ~w837 & ~w839;
assign w841 = ~w838 & ~w840;
assign w842 = ~w836 & ~w841;
assign w843 = ~w166 & w609;
assign w844 = w820 & w843;
assign w845 = (~w2916 & w2986) | (~w2916 & w2987) | (w2986 & w2987);
assign w846 = ~pi256 & w837;
assign w847 = pi027 & ~w844;
assign w848 = ~w837 & ~w847;
assign w849 = ~w846 & ~w848;
assign w850 = ~w845 & ~w849;
assign w851 = w745 & w834;
assign w852 = pi028 & ~w851;
assign w853 = ~w535 & ~w852;
assign w854 = pi028 & ~pi270;
assign w855 = ~w562 & ~w854;
assign w856 = w535 & w855;
assign w857 = ~w853 & ~w856;
assign w858 = w557 & ~w856;
assign w859 = w745 & w858;
assign w860 = (~w2916 & w2988) | (~w2916 & w2989) | (w2988 & w2989);
assign w861 = ~w857 & ~w860;
assign w862 = ~w166 & w636;
assign w863 = w820 & w862;
assign w864 = (~w2916 & w2990) | (~w2916 & w2991) | (w2990 & w2991);
assign w865 = ~pi258 & w837;
assign w866 = pi029 & ~w863;
assign w867 = ~w837 & ~w866;
assign w868 = ~w865 & ~w867;
assign w869 = ~w864 & ~w868;
assign w870 = w773 & w820;
assign w871 = pi030 & ~w870;
assign w872 = ~w535 & ~w871;
assign w873 = pi030 & ~pi272;
assign w874 = ~w681 & ~w873;
assign w875 = w535 & w874;
assign w876 = ~w872 & ~w875;
assign w877 = w163 & ~w875;
assign w878 = w829 & w877;
assign w879 = (~w2916 & w2992) | (~w2916 & w2993) | (w2992 & w2993);
assign w880 = ~w876 & ~w879;
assign w881 = pi031 & ~w689;
assign w882 = pi266 & pi273;
assign w883 = w563 & w882;
assign w884 = ~w881 & ~w883;
assign w885 = w636 & w694;
assign w886 = w884 & w885;
assign w887 = (w2916 & w2994) | (w2916 & w2995) | (w2994 & w2995);
assign w888 = ~pi031 & ~w885;
assign w889 = ~w167 & ~w888;
assign w890 = w884 & ~w889;
assign w891 = ~w887 & ~w890;
assign w892 = pi032 & ~w689;
assign w893 = pi263 & pi273;
assign w894 = w563 & w893;
assign w895 = ~w892 & ~w894;
assign w896 = w556 & w694;
assign w897 = w895 & w896;
assign w898 = (w2916 & w2996) | (w2916 & w2997) | (w2996 & w2997);
assign w899 = ~pi032 & ~w896;
assign w900 = ~w167 & ~w899;
assign w901 = w895 & ~w900;
assign w902 = ~w898 & ~w901;
assign w903 = w515 & w558;
assign w904 = ~pi033 & ~w903;
assign w905 = ~w167 & ~w904;
assign w906 = w549 & w563;
assign w907 = pi033 & ~w566;
assign w908 = ~w906 & ~w907;
assign w909 = ~w905 & w908;
assign w910 = w903 & w908;
assign w911 = (w2916 & w2998) | (w2916 & w2999) | (w2998 & w2999);
assign w912 = ~w909 & ~w911;
assign w913 = ~w162 & w624;
assign w914 = w558 & w913;
assign w915 = ~pi034 & ~w914;
assign w916 = ~w167 & ~w915;
assign w917 = pi034 & ~w566;
assign w918 = pi241 & pi270;
assign w919 = w563 & w918;
assign w920 = ~w917 & ~w919;
assign w921 = ~w916 & w920;
assign w922 = w914 & w920;
assign w923 = (w2916 & w3000) | (w2916 & w3001) | (w3000 & w3001);
assign w924 = ~w921 & ~w923;
assign w925 = w558 & w649;
assign w926 = ~pi035 & ~w925;
assign w927 = ~w167 & ~w926;
assign w928 = pi035 & ~w566;
assign w929 = pi243 & pi270;
assign w930 = w563 & w929;
assign w931 = ~w928 & ~w930;
assign w932 = ~w927 & w931;
assign w933 = w925 & w931;
assign w934 = (w2916 & w3002) | (w2916 & w3003) | (w3002 & w3003);
assign w935 = ~w932 & ~w934;
assign w936 = w86 & w665;
assign w937 = pi036 & ~w566;
assign w938 = pi244 & pi270;
assign w939 = w563 & w938;
assign w940 = ~w937 & ~w939;
assign w941 = w936 & w940;
assign w942 = (w2916 & w3004) | (w2916 & w3005) | (w3004 & w3005);
assign w943 = pi036 & w744;
assign w944 = ~w167 & w936;
assign w945 = w940 & ~w943;
assign w946 = ~w944 & w945;
assign w947 = ~w942 & ~w946;
assign w948 = w514 & w610;
assign w949 = ~pi037 & ~w948;
assign w950 = ~w167 & ~w949;
assign w951 = pi037 & ~w615;
assign w952 = w563 & w790;
assign w953 = ~w951 & ~w952;
assign w954 = ~w950 & w953;
assign w955 = w948 & w953;
assign w956 = (w2916 & w3006) | (w2916 & w3007) | (w3006 & w3007);
assign w957 = ~w954 & ~w956;
assign w958 = w556 & w610;
assign w959 = ~pi038 & ~w958;
assign w960 = ~w167 & ~w959;
assign w961 = pi038 & ~w615;
assign w962 = pi247 & pi271;
assign w963 = w563 & w962;
assign w964 = ~w961 & ~w963;
assign w965 = ~w960 & w964;
assign w966 = w958 & w964;
assign w967 = (w2916 & w3008) | (w2916 & w3009) | (w3008 & w3009);
assign w968 = ~w965 & ~w967;
assign w969 = w610 & w648;
assign w970 = ~pi039 & ~w969;
assign w971 = ~w167 & ~w970;
assign w972 = pi039 & ~w615;
assign w973 = pi251 & pi271;
assign w974 = w563 & w973;
assign w975 = ~w972 & ~w974;
assign w976 = ~w971 & w975;
assign w977 = w969 & w975;
assign w978 = (w2916 & w3010) | (w2916 & w3011) | (w3010 & w3011);
assign w979 = ~w976 & ~w978;
assign w980 = w515 & w650;
assign w981 = ~pi040 & ~w980;
assign w982 = ~w167 & ~w981;
assign w983 = pi040 & ~w655;
assign w984 = w563 & w825;
assign w985 = ~w983 & ~w984;
assign w986 = ~w982 & w985;
assign w987 = w980 & w985;
assign w988 = (w2916 & w3012) | (w2916 & w3013) | (w3012 & w3013);
assign w989 = ~w986 & ~w988;
assign w990 = w650 & w913;
assign w991 = ~pi041 & ~w990;
assign w992 = ~w167 & ~w991;
assign w993 = pi041 & ~w655;
assign w994 = pi257 & w670;
assign w995 = ~w993 & ~w994;
assign w996 = ~w992 & w995;
assign w997 = w990 & w995;
assign w998 = (w2916 & w3014) | (w2916 & w3015) | (w3014 & w3015);
assign w999 = ~w996 & ~w998;
assign w1000 = w70 & w573;
assign w1001 = w587 & w1000;
assign w1002 = ~pi042 & ~w1001;
assign w1003 = ~w167 & ~w1002;
assign w1004 = pi042 & ~w655;
assign w1005 = pi258 & w670;
assign w1006 = ~w1004 & ~w1005;
assign w1007 = ~w1003 & w1006;
assign w1008 = w1001 & w1006;
assign w1009 = (w2916 & w3016) | (w2916 & w3017) | (w3016 & w3017);
assign w1010 = ~w1007 & ~w1009;
assign w1011 = w557 & w650;
assign w1012 = ~pi043 & ~w1011;
assign w1013 = ~w167 & ~w1012;
assign w1014 = pi043 & ~w655;
assign w1015 = pi255 & w670;
assign w1016 = ~w1014 & ~w1015;
assign w1017 = ~w1013 & w1016;
assign w1018 = w1011 & w1016;
assign w1019 = (w2916 & w3018) | (w2916 & w3019) | (w3018 & w3019);
assign w1020 = ~w1017 & ~w1019;
assign w1021 = w522 & w563;
assign w1022 = pi044 & ~w689;
assign w1023 = ~w1021 & ~w1022;
assign w1024 = w514 & w694;
assign w1025 = w1023 & w1024;
assign w1026 = (w2916 & w3020) | (w2916 & w3021) | (w3020 & w3021);
assign w1027 = ~pi044 & ~w1024;
assign w1028 = ~w167 & ~w1027;
assign w1029 = w1023 & ~w1028;
assign w1030 = ~w1026 & ~w1029;
assign w1031 = w575 & w1000;
assign w1032 = ~pi045 & ~w1031;
assign w1033 = ~w167 & ~w1032;
assign w1034 = pi045 & ~w655;
assign w1035 = pi256 & w670;
assign w1036 = ~w1034 & ~w1035;
assign w1037 = ~w1033 & w1036;
assign w1038 = w1031 & w1036;
assign w1039 = (w2916 & w3022) | (w2916 & w3023) | (w3022 & w3023);
assign w1040 = ~w1037 & ~w1039;
assign w1041 = pi046 & ~w689;
assign w1042 = pi264 & pi273;
assign w1043 = w563 & w1042;
assign w1044 = ~w1041 & ~w1043;
assign w1045 = w609 & w694;
assign w1046 = w1044 & w1045;
assign w1047 = (w2916 & w3024) | (w2916 & w3025) | (w3024 & w3025);
assign w1048 = ~pi046 & ~w1045;
assign w1049 = ~w167 & ~w1048;
assign w1050 = w1044 & ~w1049;
assign w1051 = ~w1047 & ~w1050;
assign w1052 = w156 & w610;
assign w1053 = ~pi047 & ~w1052;
assign w1054 = ~w167 & ~w1053;
assign w1055 = pi047 & ~w615;
assign w1056 = w563 & w812;
assign w1057 = ~w1055 & ~w1056;
assign w1058 = ~w1054 & w1057;
assign w1059 = w1052 & w1057;
assign w1060 = (w2916 & w3026) | (w2916 & w3027) | (w3026 & w3027);
assign w1061 = ~w1058 & ~w1060;
assign w1062 = w610 & w664;
assign w1063 = ~pi048 & ~w1062;
assign w1064 = ~w167 & ~w1063;
assign w1065 = pi048 & ~w615;
assign w1066 = pi252 & pi271;
assign w1067 = w563 & w1066;
assign w1068 = ~w1065 & ~w1067;
assign w1069 = ~w1064 & w1068;
assign w1070 = w1062 & w1068;
assign w1071 = (w2916 & w3028) | (w2916 & w3029) | (w3028 & w3029);
assign w1072 = ~w1069 & ~w1071;
assign w1073 = w350 & w734;
assign w1074 = w843 & w1073;
assign w1075 = (~w2916 & w3030) | (~w2916 & w3031) | (w3030 & w3031);
assign w1076 = pi273 & w535;
assign w1077 = pi264 & w1076;
assign w1078 = pi049 & ~w1076;
assign w1079 = ~w1074 & w1078;
assign w1080 = ~w1077 & ~w1079;
assign w1081 = ~w1075 & w1080;
assign w1082 = ~w166 & w624;
assign w1083 = w1073 & w1082;
assign w1084 = (~w2916 & w3032) | (~w2916 & w3033) | (w3032 & w3033);
assign w1085 = pi265 & w1076;
assign w1086 = pi050 & ~w1076;
assign w1087 = ~w1083 & w1086;
assign w1088 = ~w1085 & ~w1087;
assign w1089 = ~w1084 & w1088;
assign w1090 = w785 & w1073;
assign w1091 = (~w2916 & w3034) | (~w2916 & w3035) | (w3034 & w3035);
assign w1092 = pi051 & ~w1076;
assign w1093 = ~w1090 & w1092;
assign w1094 = pi262 & w1076;
assign w1095 = ~w1093 & ~w1094;
assign w1096 = ~w1091 & w1095;
assign w1097 = ~w166 & w648;
assign w1098 = w1073 & w1097;
assign w1099 = (~w2916 & w3036) | (~w2916 & w3037) | (w3036 & w3037);
assign w1100 = pi267 & w1076;
assign w1101 = pi052 & ~w1076;
assign w1102 = ~w1098 & w1101;
assign w1103 = ~w1100 & ~w1102;
assign w1104 = ~w1099 & w1103;
assign w1105 = w862 & w1073;
assign w1106 = (~w2916 & w3038) | (~w2916 & w3039) | (w3038 & w3039);
assign w1107 = pi266 & w1076;
assign w1108 = pi053 & ~w1076;
assign w1109 = ~w1105 & w1108;
assign w1110 = ~w1107 & ~w1109;
assign w1111 = ~w1106 & w1110;
assign w1112 = w799 & w1073;
assign w1113 = (~w2916 & w3040) | (~w2916 & w3041) | (w3040 & w3041);
assign w1114 = pi268 & w1076;
assign w1115 = pi054 & ~w1076;
assign w1116 = ~w1112 & w1115;
assign w1117 = ~w1114 & ~w1116;
assign w1118 = ~w1113 & w1117;
assign w1119 = w773 & w1073;
assign w1120 = (~w2916 & w3042) | (~w2916 & w3043) | (w3042 & w3043);
assign w1121 = pi269 & w1076;
assign w1122 = pi055 & ~w1076;
assign w1123 = ~w1119 & w1122;
assign w1124 = ~w1121 & ~w1123;
assign w1125 = ~w1120 & w1124;
assign w1126 = w784 & w843;
assign w1127 = ~pi056 & ~w802;
assign w1128 = ~w1126 & w1127;
assign w1129 = ~w529 & ~w1128;
assign w1130 = (~w2916 & w3044) | (~w2916 & w3045) | (w3044 & w3045);
assign w1131 = ~pi248 & w802;
assign w1132 = ~w1127 & ~w1131;
assign w1133 = ~w1126 & w1132;
assign w1134 = ~w1130 & ~w1133;
assign w1135 = w735 & w1082;
assign w1136 = (~w2916 & w3046) | (~w2916 & w3047) | (w3046 & w3047);
assign w1137 = ~w529 & ~w1135;
assign w1138 = ~w777 & ~w1137;
assign w1139 = pi057 & ~w1138;
assign w1140 = w535 & w918;
assign w1141 = ~w1139 & ~w1140;
assign w1142 = ~w1136 & w1141;
assign w1143 = w735 & w1097;
assign w1144 = (~w2916 & w3048) | (~w2916 & w3049) | (w3048 & w3049);
assign w1145 = ~w529 & ~w1143;
assign w1146 = ~w777 & ~w1145;
assign w1147 = pi058 & ~w1146;
assign w1148 = w535 & w929;
assign w1149 = ~w1147 & ~w1148;
assign w1150 = ~w1144 & w1149;
assign w1151 = w834 & w1073;
assign w1152 = (~w2916 & w3050) | (~w2916 & w3051) | (w3050 & w3051);
assign w1153 = pi263 & w1076;
assign w1154 = pi059 & ~w1076;
assign w1155 = ~w1151 & w1154;
assign w1156 = ~w1153 & ~w1155;
assign w1157 = ~w1152 & w1156;
assign w1158 = w735 & w799;
assign w1159 = (~w2916 & w3052) | (~w2916 & w3053) | (w3052 & w3053);
assign w1160 = ~w529 & ~w1158;
assign w1161 = ~w777 & ~w1160;
assign w1162 = pi060 & ~w1161;
assign w1163 = w535 & w938;
assign w1164 = ~w1162 & ~w1163;
assign w1165 = ~w1159 & w1164;
assign w1166 = w784 & w862;
assign w1167 = (~w2916 & w3054) | (~w2916 & w3055) | (w3054 & w3055);
assign w1168 = pi250 & w802;
assign w1169 = pi061 & ~w802;
assign w1170 = ~w1166 & w1169;
assign w1171 = ~w1168 & ~w1170;
assign w1172 = ~w1167 & w1171;
assign w1173 = w784 & w1097;
assign w1174 = (~w2916 & w3056) | (~w2916 & w3057) | (w3056 & w3057);
assign w1175 = pi062 & ~w802;
assign w1176 = ~w1173 & w1175;
assign w1177 = pi251 & w802;
assign w1178 = ~w1176 & ~w1177;
assign w1179 = ~w1174 & w1178;
assign w1180 = w784 & w1082;
assign w1181 = (~w2916 & w3058) | (~w2916 & w3059) | (w3058 & w3059);
assign w1182 = pi249 & w802;
assign w1183 = pi063 & ~w802;
assign w1184 = ~w1180 & w1183;
assign w1185 = ~w1182 & ~w1184;
assign w1186 = ~w1181 & w1185;
assign w1187 = w784 & w834;
assign w1188 = (~w2916 & w3060) | (~w2916 & w3061) | (w3060 & w3061);
assign w1189 = pi247 & w802;
assign w1190 = pi064 & ~w802;
assign w1191 = ~w1187 & w1190;
assign w1192 = ~w1189 & ~w1191;
assign w1193 = ~w1188 & w1192;
assign w1194 = w820 & w1082;
assign w1195 = (~w2916 & w3062) | (~w2916 & w3063) | (w3062 & w3063);
assign w1196 = ~pi257 & w837;
assign w1197 = pi065 & ~w1194;
assign w1198 = ~w837 & ~w1197;
assign w1199 = ~w1196 & ~w1198;
assign w1200 = ~w1195 & ~w1199;
assign w1201 = w820 & w1097;
assign w1202 = (~w2916 & w3064) | (~w2916 & w3065) | (w3064 & w3065);
assign w1203 = pi259 & w837;
assign w1204 = pi066 & ~w837;
assign w1205 = ~w1201 & w1204;
assign w1206 = ~w1203 & ~w1205;
assign w1207 = ~w1202 & w1206;
assign w1208 = w799 & w820;
assign w1209 = (~w2916 & w3066) | (~w2916 & w3067) | (w3066 & w3067);
assign w1210 = ~pi260 & w837;
assign w1211 = pi067 & ~w1208;
assign w1212 = ~w837 & ~w1211;
assign w1213 = ~w1210 & ~w1212;
assign w1214 = ~w1209 & ~w1213;
assign w1215 = w130 & w370;
assign w1216 = w1097 & w1215;
assign w1217 = (~w2916 & w3068) | (~w2916 & w3069) | (w3068 & w3069);
assign w1218 = pi272 & w171;
assign w1219 = pi259 & w1218;
assign w1220 = pi068 & ~w1218;
assign w1221 = ~w1216 & w1220;
assign w1222 = ~w1219 & ~w1221;
assign w1223 = ~w1217 & w1222;
assign w1224 = w799 & w1215;
assign w1225 = (~w2916 & w3070) | (~w2916 & w3071) | (w3070 & w3071);
assign w1226 = ~pi260 & w1218;
assign w1227 = pi069 & ~w1224;
assign w1228 = ~w1218 & ~w1227;
assign w1229 = ~w1226 & ~w1228;
assign w1230 = ~w1225 & ~w1229;
assign w1231 = w1082 & w1215;
assign w1232 = (~w2916 & w3072) | (~w2916 & w3073) | (w3072 & w3073);
assign w1233 = ~pi257 & w1218;
assign w1234 = pi070 & ~w1231;
assign w1235 = ~w1218 & ~w1234;
assign w1236 = ~w1233 & ~w1235;
assign w1237 = ~w1232 & ~w1236;
assign w1238 = ~w530 & w556;
assign w1239 = w131 & w1238;
assign w1240 = ~pi071 & ~w1239;
assign w1241 = ~w529 & ~w1240;
assign w1242 = w171 & w562;
assign w1243 = ~w172 & ~w535;
assign w1244 = pi071 & ~w1243;
assign w1245 = ~w1242 & ~w1244;
assign w1246 = ~w1241 & w1245;
assign w1247 = w1239 & w1245;
assign w1248 = (w2916 & w3074) | (w2916 & w3075) | (w3074 & w3075);
assign w1249 = ~w1246 & ~w1248;
assign w1250 = ~w530 & w609;
assign w1251 = w131 & w1250;
assign w1252 = ~pi072 & ~w1251;
assign w1253 = ~w529 & ~w1252;
assign w1254 = w171 & w580;
assign w1255 = pi072 & ~w1243;
assign w1256 = ~w1254 & ~w1255;
assign w1257 = ~w1253 & w1256;
assign w1258 = w1251 & w1256;
assign w1259 = (w2916 & w3076) | (w2916 & w3077) | (w3076 & w3077);
assign w1260 = ~w1257 & ~w1259;
assign w1261 = ~w530 & w624;
assign w1262 = w131 & w1261;
assign w1263 = ~pi073 & ~w1262;
assign w1264 = ~w529 & ~w1263;
assign w1265 = w171 & w918;
assign w1266 = pi073 & ~w1243;
assign w1267 = ~w1265 & ~w1266;
assign w1268 = ~w1264 & w1267;
assign w1269 = w1262 & w1267;
assign w1270 = (w2916 & w3078) | (w2916 & w3079) | (w3078 & w3079);
assign w1271 = ~w1268 & ~w1270;
assign w1272 = ~w530 & w636;
assign w1273 = w131 & w1272;
assign w1274 = ~pi074 & ~w1273;
assign w1275 = ~w529 & ~w1274;
assign w1276 = w171 & w592;
assign w1277 = pi074 & ~w1243;
assign w1278 = ~w1276 & ~w1277;
assign w1279 = ~w1275 & w1278;
assign w1280 = w1273 & w1278;
assign w1281 = (w2916 & w3080) | (w2916 & w3081) | (w3080 & w3081);
assign w1282 = ~w1279 & ~w1281;
assign w1283 = w130 & w389;
assign w1284 = w1082 & w1283;
assign w1285 = (~w2916 & w3082) | (~w2916 & w3083) | (w3082 & w3083);
assign w1286 = pi271 & w171;
assign w1287 = pi249 & w1286;
assign w1288 = pi075 & ~w1286;
assign w1289 = ~w1284 & w1288;
assign w1290 = ~w1287 & ~w1289;
assign w1291 = ~w1285 & w1290;
assign w1292 = w1097 & w1283;
assign w1293 = (~w2916 & w3084) | (~w2916 & w3085) | (w3084 & w3085);
assign w1294 = pi251 & w1286;
assign w1295 = pi076 & ~w1286;
assign w1296 = ~w1292 & w1295;
assign w1297 = ~w1294 & ~w1296;
assign w1298 = ~w1293 & w1297;
assign w1299 = w799 & w1283;
assign w1300 = (~w2916 & w3086) | (~w2916 & w3087) | (w3086 & w3087);
assign w1301 = pi252 & w1286;
assign w1302 = pi077 & ~w1286;
assign w1303 = ~w1299 & w1302;
assign w1304 = ~w1301 & ~w1303;
assign w1305 = ~w1300 & w1304;
assign w1306 = w773 & w1283;
assign w1307 = (~w2916 & w3088) | (~w2916 & w3089) | (w3088 & w3089);
assign w1308 = pi253 & w1286;
assign w1309 = pi078 & ~w1286;
assign w1310 = ~w1306 & w1309;
assign w1311 = ~w1308 & ~w1310;
assign w1312 = ~w1307 & w1311;
assign w1313 = w513 & w1238;
assign w1314 = ~pi079 & ~w1313;
assign w1315 = ~w529 & ~w1314;
assign w1316 = pi079 & ~w536;
assign w1317 = w171 & w893;
assign w1318 = ~w1316 & ~w1317;
assign w1319 = ~w1315 & w1318;
assign w1320 = w1313 & w1318;
assign w1321 = (w2916 & w3090) | (w2916 & w3091) | (w3090 & w3091);
assign w1322 = ~w1319 & ~w1321;
assign w1323 = w513 & w1250;
assign w1324 = ~pi080 & ~w1323;
assign w1325 = ~w529 & ~w1324;
assign w1326 = pi080 & ~w536;
assign w1327 = w171 & w1042;
assign w1328 = ~w1326 & ~w1327;
assign w1329 = ~w1325 & w1328;
assign w1330 = w1323 & w1328;
assign w1331 = (w2916 & w3092) | (w2916 & w3093) | (w3092 & w3093);
assign w1332 = ~w1329 & ~w1331;
assign w1333 = w513 & w1261;
assign w1334 = ~pi081 & ~w1333;
assign w1335 = ~w529 & ~w1334;
assign w1336 = pi081 & ~w536;
assign w1337 = w171 & w691;
assign w1338 = ~w1336 & ~w1337;
assign w1339 = ~w1335 & w1338;
assign w1340 = w1333 & w1338;
assign w1341 = (w2916 & w3094) | (w2916 & w3095) | (w3094 & w3095);
assign w1342 = ~w1339 & ~w1341;
assign w1343 = ~w530 & w648;
assign w1344 = w513 & w1343;
assign w1345 = ~pi082 & ~w1344;
assign w1346 = ~w529 & ~w1345;
assign w1347 = pi082 & ~w536;
assign w1348 = w171 & w703;
assign w1349 = ~w1347 & ~w1348;
assign w1350 = ~w1346 & w1349;
assign w1351 = w1344 & w1349;
assign w1352 = (w2916 & w3096) | (w2916 & w3097) | (w3096 & w3097);
assign w1353 = ~w1350 & ~w1352;
assign w1354 = ~w530 & w664;
assign w1355 = w513 & w1354;
assign w1356 = ~pi083 & ~w1355;
assign w1357 = ~w529 & ~w1356;
assign w1358 = pi083 & ~w536;
assign w1359 = w171 & w717;
assign w1360 = ~w1358 & ~w1359;
assign w1361 = ~w1357 & w1360;
assign w1362 = w1355 & w1360;
assign w1363 = (w2916 & w3098) | (w2916 & w3099) | (w3098 & w3099);
assign w1364 = ~w1361 & ~w1363;
assign w1365 = w389 & w431;
assign w1366 = w514 & ~w529;
assign w1367 = w1365 & w1366;
assign w1368 = ~pi084 & ~w1367;
assign w1369 = ~w530 & ~w1368;
assign w1370 = pi271 & w160;
assign w1371 = w166 & ~w1370;
assign w1372 = pi084 & w1371;
assign w1373 = w166 & w1370;
assign w1374 = pi246 & w1373;
assign w1375 = ~w1372 & ~w1374;
assign w1376 = ~w1369 & w1375;
assign w1377 = w514 & w1375;
assign w1378 = w1365 & w1377;
assign w1379 = (w2916 & w3100) | (w2916 & w3101) | (w3100 & w3101);
assign w1380 = ~w1376 & ~w1379;
assign w1381 = pi085 & w1371;
assign w1382 = pi253 & w1373;
assign w1383 = ~w1381 & ~w1382;
assign w1384 = w156 & w1383;
assign w1385 = w1365 & w1384;
assign w1386 = (w2916 & w3102) | (w2916 & w3103) | (w3102 & w3103);
assign w1387 = pi085 & ~w530;
assign w1388 = w773 & w1365;
assign w1389 = w1383 & ~w1387;
assign w1390 = ~w1388 & w1389;
assign w1391 = ~w1386 & ~w1390;
assign w1392 = w370 & w431;
assign w1393 = w1366 & w1392;
assign w1394 = ~pi086 & ~w1393;
assign w1395 = ~w530 & ~w1394;
assign w1396 = pi272 & w160;
assign w1397 = w166 & ~w1396;
assign w1398 = pi086 & w1397;
assign w1399 = w166 & w1396;
assign w1400 = pi254 & w1399;
assign w1401 = ~w1398 & ~w1400;
assign w1402 = ~w1395 & w1401;
assign w1403 = w514 & w1401;
assign w1404 = w1392 & w1403;
assign w1405 = (w2916 & w3104) | (w2916 & w3105) | (w3104 & w3105);
assign w1406 = ~w1402 & ~w1405;
assign w1407 = pi087 & w1397;
assign w1408 = pi261 & w1399;
assign w1409 = ~w1407 & ~w1408;
assign w1410 = w156 & w1409;
assign w1411 = w1392 & w1410;
assign w1412 = (w2916 & w3106) | (w2916 & w3107) | (w3106 & w3107);
assign w1413 = pi087 & ~w530;
assign w1414 = w773 & w1392;
assign w1415 = w1409 & ~w1413;
assign w1416 = ~w1414 & w1415;
assign w1417 = ~w1412 & ~w1416;
assign w1418 = w129 & w3261;
assign w1419 = pi273 & w160;
assign w1420 = w166 & ~w1419;
assign w1421 = pi088 & w1420;
assign w1422 = w162 & w893;
assign w1423 = ~w1421 & ~w1422;
assign w1424 = w556 & w1423;
assign w1425 = w1418 & w1424;
assign w1426 = (w2916 & w3108) | (w2916 & w3109) | (w3108 & w3109);
assign w1427 = pi088 & ~w530;
assign w1428 = w834 & w1418;
assign w1429 = w1423 & ~w1427;
assign w1430 = ~w1428 & w1429;
assign w1431 = ~w1426 & ~w1430;
assign w1432 = w86 & w431;
assign w1433 = pi270 & w160;
assign w1434 = w166 & ~w1433;
assign w1435 = pi089 & w1434;
assign w1436 = w162 & w562;
assign w1437 = ~w1435 & ~w1436;
assign w1438 = w556 & w1437;
assign w1439 = w1432 & w1438;
assign w1440 = (w2916 & w3110) | (w2916 & w3111) | (w3110 & w3111);
assign w1441 = pi089 & ~w530;
assign w1442 = w834 & w1432;
assign w1443 = w1437 & ~w1441;
assign w1444 = ~w1442 & w1443;
assign w1445 = ~w1440 & ~w1444;
assign w1446 = pi090 & w1420;
assign w1447 = w162 & w691;
assign w1448 = ~w1446 & ~w1447;
assign w1449 = w624 & w1448;
assign w1450 = w1418 & w1449;
assign w1451 = (w2916 & w3112) | (w2916 & w3113) | (w3112 & w3113);
assign w1452 = pi090 & ~w530;
assign w1453 = w1082 & w1418;
assign w1454 = w1448 & ~w1452;
assign w1455 = ~w1453 & w1454;
assign w1456 = ~w1451 & ~w1455;
assign w1457 = pi091 & w1420;
assign w1458 = w162 & w703;
assign w1459 = ~w1457 & ~w1458;
assign w1460 = w648 & w1459;
assign w1461 = w1418 & w1460;
assign w1462 = (w2916 & w3114) | (w2916 & w3115) | (w3114 & w3115);
assign w1463 = pi091 & ~w530;
assign w1464 = w1097 & w1418;
assign w1465 = w1459 & ~w1463;
assign w1466 = ~w1464 & w1465;
assign w1467 = ~w1462 & ~w1466;
assign w1468 = pi092 & w1420;
assign w1469 = w162 & w717;
assign w1470 = ~w1468 & ~w1469;
assign w1471 = w664 & w1470;
assign w1472 = w1418 & w1471;
assign w1473 = (w2916 & w3116) | (w2916 & w3117) | (w3116 & w3117);
assign w1474 = pi092 & ~w530;
assign w1475 = w799 & w1418;
assign w1476 = w1470 & ~w1474;
assign w1477 = ~w1475 & w1476;
assign w1478 = ~w1473 & ~w1477;
assign w1479 = pi093 & w1420;
assign w1480 = w162 & w1042;
assign w1481 = ~w1479 & ~w1480;
assign w1482 = w609 & w1481;
assign w1483 = w1418 & w1482;
assign w1484 = (w2916 & w3118) | (w2916 & w3119) | (w3118 & w3119);
assign w1485 = pi093 & ~w530;
assign w1486 = w843 & w1418;
assign w1487 = w1481 & ~w1485;
assign w1488 = ~w1486 & w1487;
assign w1489 = ~w1484 & ~w1488;
assign w1490 = pi094 & w1420;
assign w1491 = w162 & w538;
assign w1492 = ~w1490 & ~w1491;
assign w1493 = w156 & w1492;
assign w1494 = w1418 & w1493;
assign w1495 = (w2916 & w3120) | (w2916 & w3121) | (w3120 & w3121);
assign w1496 = pi094 & ~w530;
assign w1497 = w773 & w1418;
assign w1498 = w1492 & ~w1496;
assign w1499 = ~w1497 & w1498;
assign w1500 = ~w1495 & ~w1499;
assign w1501 = pi095 & w1420;
assign w1502 = w162 & w882;
assign w1503 = ~w1501 & ~w1502;
assign w1504 = w636 & w1503;
assign w1505 = w1418 & w1504;
assign w1506 = (w2916 & w3122) | (w2916 & w3123) | (w3122 & w3123);
assign w1507 = pi095 & ~w530;
assign w1508 = w862 & w1418;
assign w1509 = w1503 & ~w1507;
assign w1510 = ~w1508 & w1509;
assign w1511 = ~w1506 & ~w1510;
assign w1512 = pi096 & w1434;
assign w1513 = w162 & w580;
assign w1514 = ~w1512 & ~w1513;
assign w1515 = w609 & w1514;
assign w1516 = w1432 & w1515;
assign w1517 = (w2916 & w3124) | (w2916 & w3125) | (w3124 & w3125);
assign w1518 = pi096 & ~w530;
assign w1519 = w843 & w1432;
assign w1520 = w1514 & ~w1518;
assign w1521 = ~w1519 & w1520;
assign w1522 = ~w1517 & ~w1521;
assign w1523 = pi097 & w1397;
assign w1524 = pi256 & w1399;
assign w1525 = ~w1523 & ~w1524;
assign w1526 = w609 & w1525;
assign w1527 = w1392 & w1526;
assign w1528 = (w2916 & w3126) | (w2916 & w3127) | (w3126 & w3127);
assign w1529 = pi097 & ~w530;
assign w1530 = w843 & w1392;
assign w1531 = w1525 & ~w1529;
assign w1532 = ~w1530 & w1531;
assign w1533 = ~w1528 & ~w1532;
assign w1534 = w513 & w1272;
assign w1535 = ~pi098 & ~w1534;
assign w1536 = ~w529 & ~w1535;
assign w1537 = pi098 & ~w536;
assign w1538 = w171 & w882;
assign w1539 = ~w1537 & ~w1538;
assign w1540 = ~w1536 & w1539;
assign w1541 = w1534 & w1539;
assign w1542 = (w2916 & w3128) | (w2916 & w3129) | (w3128 & w3129);
assign w1543 = ~w1540 & ~w1542;
assign w1544 = w785 & w1215;
assign w1545 = (~w2916 & w3130) | (~w2916 & w3131) | (w3130 & w3131);
assign w1546 = pi254 & w1218;
assign w1547 = pi099 & ~w1218;
assign w1548 = ~w1544 & w1547;
assign w1549 = ~w1546 & ~w1548;
assign w1550 = ~w1545 & w1549;
assign w1551 = w834 & w1283;
assign w1552 = (~w2916 & w3132) | (~w2916 & w3133) | (w3132 & w3133);
assign w1553 = pi247 & w1286;
assign w1554 = pi100 & ~w1286;
assign w1555 = ~w1551 & w1554;
assign w1556 = ~w1553 & ~w1555;
assign w1557 = ~w1552 & w1556;
assign w1558 = w785 & w1283;
assign w1559 = (~w2916 & w3134) | (~w2916 & w3135) | (w3134 & w3135);
assign w1560 = pi246 & w1286;
assign w1561 = pi101 & ~w1286;
assign w1562 = ~w1558 & w1561;
assign w1563 = ~w1560 & ~w1562;
assign w1564 = ~w1559 & w1563;
assign w1565 = w514 & w1418;
assign w1566 = ~w530 & ~w1565;
assign w1567 = ~w1420 & ~w1566;
assign w1568 = pi102 & ~w1567;
assign w1569 = w162 & w522;
assign w1570 = ~w166 & w1565;
assign w1571 = (~w2916 & w3136) | (~w2916 & w3137) | (w3136 & w3137);
assign w1572 = ~w1568 & ~w1569;
assign w1573 = ~w1571 & w1572;
assign w1574 = pi103 & w1371;
assign w1575 = pi247 & w1373;
assign w1576 = ~w1574 & ~w1575;
assign w1577 = w556 & w1576;
assign w1578 = w1365 & w1577;
assign w1579 = (w2916 & w3138) | (w2916 & w3139) | (w3138 & w3139);
assign w1580 = pi103 & ~w530;
assign w1581 = w834 & w1365;
assign w1582 = w1576 & ~w1580;
assign w1583 = ~w1581 & w1582;
assign w1584 = ~w1579 & ~w1583;
assign w1585 = pi104 & w1397;
assign w1586 = pi255 & w1399;
assign w1587 = ~w1585 & ~w1586;
assign w1588 = w556 & w1587;
assign w1589 = w1392 & w1588;
assign w1590 = (w2916 & w3140) | (w2916 & w3141) | (w3140 & w3141);
assign w1591 = pi104 & ~w530;
assign w1592 = w834 & w1392;
assign w1593 = w1587 & ~w1591;
assign w1594 = ~w1592 & w1593;
assign w1595 = ~w1590 & ~w1594;
assign w1596 = pi105 & w1371;
assign w1597 = pi250 & w1373;
assign w1598 = ~w1596 & ~w1597;
assign w1599 = w636 & w1598;
assign w1600 = w1365 & w1599;
assign w1601 = (w2916 & w3142) | (w2916 & w3143) | (w3142 & w3143);
assign w1602 = pi105 & ~w530;
assign w1603 = w862 & w1365;
assign w1604 = w1598 & ~w1602;
assign w1605 = ~w1603 & w1604;
assign w1606 = ~w1601 & ~w1605;
assign w1607 = w131 & w1343;
assign w1608 = ~pi106 & ~w1607;
assign w1609 = ~w529 & ~w1608;
assign w1610 = w171 & w929;
assign w1611 = pi106 & ~w1243;
assign w1612 = ~w1610 & ~w1611;
assign w1613 = ~w1609 & w1612;
assign w1614 = w1607 & w1612;
assign w1615 = (w2916 & w3144) | (w2916 & w3145) | (w3144 & w3145);
assign w1616 = ~w1613 & ~w1615;
assign w1617 = w131 & w1354;
assign w1618 = ~pi107 & ~w1617;
assign w1619 = ~w529 & ~w1618;
assign w1620 = w171 & w938;
assign w1621 = pi107 & ~w1243;
assign w1622 = ~w1620 & ~w1621;
assign w1623 = ~w1619 & w1622;
assign w1624 = w1617 & w1622;
assign w1625 = (w2916 & w3146) | (w2916 & w3147) | (w3146 & w3147);
assign w1626 = ~w1623 & ~w1625;
assign w1627 = pi108 & w1397;
assign w1628 = pi258 & w1399;
assign w1629 = ~w1627 & ~w1628;
assign w1630 = w636 & w1629;
assign w1631 = w1392 & w1630;
assign w1632 = (w2916 & w3148) | (w2916 & w3149) | (w3148 & w3149);
assign w1633 = pi108 & ~w530;
assign w1634 = w862 & w1392;
assign w1635 = w1629 & ~w1633;
assign w1636 = ~w1634 & w1635;
assign w1637 = ~w1632 & ~w1636;
assign w1638 = w843 & w1283;
assign w1639 = (~w2916 & w3150) | (~w2916 & w3151) | (w3150 & w3151);
assign w1640 = pi109 & ~w1286;
assign w1641 = ~w1638 & w1640;
assign w1642 = pi248 & w1286;
assign w1643 = ~w1641 & ~w1642;
assign w1644 = ~w1639 & w1643;
assign w1645 = w834 & w1215;
assign w1646 = (~w2916 & w3152) | (~w2916 & w3153) | (w3152 & w3153);
assign w1647 = ~pi255 & w1218;
assign w1648 = pi110 & ~w1645;
assign w1649 = ~w1218 & ~w1648;
assign w1650 = ~w1647 & ~w1649;
assign w1651 = ~w1646 & ~w1650;
assign w1652 = w843 & w1215;
assign w1653 = (~w2916 & w3154) | (~w2916 & w3155) | (w3154 & w3155);
assign w1654 = ~pi256 & w1218;
assign w1655 = pi111 & ~w1652;
assign w1656 = ~w1218 & ~w1655;
assign w1657 = ~w1654 & ~w1656;
assign w1658 = ~w1653 & ~w1657;
assign w1659 = w862 & w1283;
assign w1660 = (~w2916 & w3156) | (~w2916 & w3157) | (w3156 & w3157);
assign w1661 = pi250 & w1286;
assign w1662 = pi112 & ~w1286;
assign w1663 = ~w1659 & w1662;
assign w1664 = ~w1661 & ~w1663;
assign w1665 = ~w1660 & w1664;
assign w1666 = w862 & w1215;
assign w1667 = (~w2916 & w3158) | (~w2916 & w3159) | (w3158 & w3159);
assign w1668 = ~pi258 & w1218;
assign w1669 = pi113 & ~w1666;
assign w1670 = ~w1218 & ~w1669;
assign w1671 = ~w1668 & ~w1670;
assign w1672 = ~w1667 & ~w1671;
assign w1673 = w773 & w1215;
assign w1674 = (~w2916 & w3160) | (~w2916 & w3161) | (w3160 & w3161);
assign w1675 = pi261 & w1218;
assign w1676 = pi114 & ~w1218;
assign w1677 = ~w1673 & w1676;
assign w1678 = ~w1675 & ~w1677;
assign w1679 = ~w1674 & w1678;
assign w1680 = w773 & w1432;
assign w1681 = (~w2916 & w3162) | (~w2916 & w3163) | (w3162 & w3163);
assign w1682 = pi270 & w162;
assign w1683 = pi115 & ~w1682;
assign w1684 = ~w1680 & w1683;
assign w1685 = pi245 & w1682;
assign w1686 = ~w1684 & ~w1685;
assign w1687 = ~w1681 & w1686;
assign w1688 = pi116 & w1434;
assign w1689 = w162 & w592;
assign w1690 = ~w1688 & ~w1689;
assign w1691 = w636 & w1690;
assign w1692 = w1432 & w1691;
assign w1693 = (w2916 & w3164) | (w2916 & w3165) | (w3164 & w3165);
assign w1694 = pi116 & ~w530;
assign w1695 = w862 & w1432;
assign w1696 = w1690 & ~w1694;
assign w1697 = ~w1695 & w1696;
assign w1698 = ~w1693 & ~w1697;
assign w1699 = pi117 & w1371;
assign w1700 = pi248 & w1373;
assign w1701 = ~w1699 & ~w1700;
assign w1702 = w609 & w1701;
assign w1703 = w1365 & w1702;
assign w1704 = (w2916 & w3166) | (w2916 & w3167) | (w3166 & w3167);
assign w1705 = pi117 & ~w530;
assign w1706 = w843 & w1365;
assign w1707 = w1701 & ~w1705;
assign w1708 = ~w1706 & w1707;
assign w1709 = ~w1704 & ~w1708;
assign w1710 = pi118 & w1434;
assign w1711 = w162 & w549;
assign w1712 = ~w1710 & ~w1711;
assign w1713 = w514 & w1712;
assign w1714 = w1432 & w1713;
assign w1715 = (w2916 & w3168) | (w2916 & w3169) | (w3168 & w3169);
assign w1716 = pi118 & ~w530;
assign w1717 = w785 & w1432;
assign w1718 = w1712 & ~w1716;
assign w1719 = ~w1717 & w1718;
assign w1720 = ~w1715 & ~w1719;
assign w1721 = pi119 & w1434;
assign w1722 = w162 & w918;
assign w1723 = ~w1721 & ~w1722;
assign w1724 = w624 & w1723;
assign w1725 = w1432 & w1724;
assign w1726 = (w2916 & w3170) | (w2916 & w3171) | (w3170 & w3171);
assign w1727 = pi119 & ~w530;
assign w1728 = w1082 & w1432;
assign w1729 = w1723 & ~w1727;
assign w1730 = ~w1728 & w1729;
assign w1731 = ~w1726 & ~w1730;
assign w1732 = pi120 & w1397;
assign w1733 = pi260 & w1399;
assign w1734 = ~w1732 & ~w1733;
assign w1735 = w664 & w1734;
assign w1736 = w1392 & w1735;
assign w1737 = (w2916 & w3172) | (w2916 & w3173) | (w3172 & w3173);
assign w1738 = pi120 & ~w530;
assign w1739 = w799 & w1392;
assign w1740 = w1734 & ~w1738;
assign w1741 = ~w1739 & w1740;
assign w1742 = ~w1737 & ~w1741;
assign w1743 = w1082 & w1392;
assign w1744 = (~w2916 & w3174) | (~w2916 & w3175) | (w3174 & w3175);
assign w1745 = ~pi257 & w1399;
assign w1746 = pi121 & ~w1743;
assign w1747 = ~w1399 & ~w1746;
assign w1748 = ~w1745 & ~w1747;
assign w1749 = ~w1744 & ~w1748;
assign w1750 = w1097 & w1432;
assign w1751 = (~w2916 & w3176) | (~w2916 & w3177) | (w3176 & w3177);
assign w1752 = ~pi243 & w1682;
assign w1753 = pi122 & ~w1750;
assign w1754 = ~w1682 & ~w1753;
assign w1755 = ~w1752 & ~w1754;
assign w1756 = ~w1751 & ~w1755;
assign w1757 = w799 & w1432;
assign w1758 = (~w2916 & w3178) | (~w2916 & w3179) | (w3178 & w3179);
assign w1759 = ~pi244 & w1682;
assign w1760 = pi123 & ~w1757;
assign w1761 = ~w1682 & ~w1760;
assign w1762 = ~w1759 & ~w1761;
assign w1763 = ~w1758 & ~w1762;
assign w1764 = pi124 & w1371;
assign w1765 = pi249 & w1373;
assign w1766 = ~w1764 & ~w1765;
assign w1767 = w624 & w1766;
assign w1768 = w1365 & w1767;
assign w1769 = (w2916 & w3180) | (w2916 & w3181) | (w3180 & w3181);
assign w1770 = pi124 & ~w530;
assign w1771 = w1082 & w1365;
assign w1772 = w1766 & ~w1770;
assign w1773 = ~w1771 & w1772;
assign w1774 = ~w1769 & ~w1773;
assign w1775 = w1097 & w1365;
assign w1776 = (~w2916 & w3182) | (~w2916 & w3183) | (w3182 & w3183);
assign w1777 = ~pi251 & w1373;
assign w1778 = pi125 & ~w1775;
assign w1779 = ~w1373 & ~w1778;
assign w1780 = ~w1777 & ~w1779;
assign w1781 = ~w1776 & ~w1780;
assign w1782 = w799 & w1365;
assign w1783 = (~w2916 & w3184) | (~w2916 & w3185) | (w3184 & w3185);
assign w1784 = ~pi252 & w1373;
assign w1785 = pi126 & ~w1782;
assign w1786 = ~w1373 & ~w1785;
assign w1787 = ~w1784 & ~w1786;
assign w1788 = ~w1783 & ~w1787;
assign w1789 = pi127 & w1397;
assign w1790 = w162 & w657;
assign w1791 = ~w1789 & ~w1790;
assign w1792 = w648 & w1791;
assign w1793 = w1392 & w1792;
assign w1794 = (w2916 & w3186) | (w2916 & w3187) | (w3186 & w3187);
assign w1795 = pi127 & ~w530;
assign w1796 = w1097 & w1392;
assign w1797 = w1791 & ~w1795;
assign w1798 = ~w1796 & w1797;
assign w1799 = ~w1794 & ~w1798;
assign w1800 = pi144 & pi146;
assign w1801 = ~pi144 & ~pi145;
assign w1802 = ~w1800 & ~w1801;
assign w1803 = ~w344 & w1802;
assign w1804 = pi136 & ~w1803;
assign w1805 = ~pi128 & w1804;
assign w1806 = ~pi143 & w103;
assign w1807 = pi140 & ~pi161;
assign w1808 = ~pi140 & pi161;
assign w1809 = ~w1807 & ~w1808;
assign w1810 = ~pi150 & pi190;
assign w1811 = (~w32 & ~w140) | (~w32 & w2917) | (~w140 & w2917);
assign w1812 = (~w151 & w1811) | (~w151 & w2918) | (w1811 & w2918);
assign w1813 = (~w16 & w1812) | (~w16 & w3188) | (w1812 & w3188);
assign w1814 = w52 & ~w1813;
assign w1815 = ~w51 & ~w1814;
assign w1816 = w1809 & ~w1815;
assign w1817 = ~w1809 & w1815;
assign w1818 = pi143 & ~w1816;
assign w1819 = ~w1817 & w1818;
assign w1820 = ~w1806 & ~w1819;
assign w1821 = ~w1807 & ~w1816;
assign w1822 = pi143 & ~w1821;
assign w1823 = pi143 & ~w112;
assign w1824 = ~pi143 & ~w120;
assign w1825 = ~w1823 & ~w1824;
assign w1826 = ~w1822 & w1825;
assign w1827 = ~w112 & w1822;
assign w1828 = ~w1826 & ~w1827;
assign w1829 = pi142 & ~w62;
assign w1830 = w79 & ~w1829;
assign w1831 = ~w43 & w1812;
assign w1832 = (pi143 & w1812) | (pi143 & w3189) | (w1812 & w3189);
assign w1833 = ~w1831 & w1832;
assign w1834 = ~w1830 & ~w1833;
assign w1835 = ~w62 & w147;
assign w1836 = ~w152 & w1811;
assign w1837 = (pi143 & w1811) | (pi143 & w2919) | (w1811 & w2919);
assign w1838 = ~w1836 & w1837;
assign w1839 = ~w1835 & ~w1838;
assign w1840 = ~w1834 & w1839;
assign w1841 = pi190 & ~w132;
assign w1842 = ~pi190 & w132;
assign w1843 = ~w1841 & ~w1842;
assign w1844 = ~w140 & ~w1810;
assign w1845 = (pi143 & ~w140) | (pi143 & w2920) | (~w140 & w2920);
assign w1846 = ~w1844 & w1845;
assign w1847 = ~pi143 & ~w9;
assign w1848 = ~w61 & w1847;
assign w1849 = ~w1846 & ~w1848;
assign w1850 = (~pi035 & w1846) | (~pi035 & w3190) | (w1846 & w3190);
assign w1851 = ~pi007 & w1849;
assign w1852 = w1843 & ~w1850;
assign w1853 = ~w1851 & w1852;
assign w1854 = (~pi006 & w1846) | (~pi006 & w3191) | (w1846 & w3191);
assign w1855 = ~pi036 & w1849;
assign w1856 = ~w1843 & ~w1854;
assign w1857 = ~w1855 & w1856;
assign w1858 = ~w1853 & ~w1857;
assign w1859 = w1840 & ~w1858;
assign w1860 = ~w1834 & ~w1839;
assign w1861 = (~pi004 & w1846) | (~pi004 & w3192) | (w1846 & w3192);
assign w1862 = ~pi034 & w1849;
assign w1863 = w1843 & ~w1861;
assign w1864 = ~w1862 & w1863;
assign w1865 = (~pi033 & w1846) | (~pi033 & w3193) | (w1846 & w3193);
assign w1866 = ~pi005 & w1849;
assign w1867 = ~w1843 & ~w1865;
assign w1868 = ~w1866 & w1867;
assign w1869 = ~w1864 & ~w1868;
assign w1870 = w1860 & ~w1869;
assign w1871 = ~pi143 & w66;
assign w1872 = ~w52 & w1813;
assign w1873 = pi143 & ~w1814;
assign w1874 = ~w1872 & w1873;
assign w1875 = ~w1871 & ~w1874;
assign w1876 = ~pi037 & ~w1843;
assign w1877 = ~pi038 & w1843;
assign w1878 = ~w1876 & ~w1877;
assign w1879 = ~w1839 & w1878;
assign w1880 = ~pi010 & ~w1843;
assign w1881 = ~pi039 & w1843;
assign w1882 = ~w1880 & ~w1881;
assign w1883 = w1839 & w1882;
assign w1884 = ~w1849 & ~w1879;
assign w1885 = ~w1883 & w1884;
assign w1886 = ~pi048 & ~w1843;
assign w1887 = ~pi047 & w1843;
assign w1888 = ~w1886 & ~w1887;
assign w1889 = w1839 & w1888;
assign w1890 = ~pi008 & ~w1843;
assign w1891 = ~pi009 & w1843;
assign w1892 = ~w1890 & ~w1891;
assign w1893 = ~w1839 & w1892;
assign w1894 = w1849 & ~w1889;
assign w1895 = ~w1893 & w1894;
assign w1896 = w1834 & ~w1885;
assign w1897 = ~w1895 & w1896;
assign w1898 = ~w1859 & ~w1870;
assign w1899 = ~w1875 & w1898;
assign w1900 = ~w1897 & w1899;
assign w1901 = ~w1838 & w3194;
assign w1902 = pi014 & ~w1839;
assign w1903 = w1843 & ~w1901;
assign w1904 = ~w1902 & w1903;
assign w1905 = ~w1838 & w3195;
assign w1906 = pi046 & ~w1839;
assign w1907 = ~w1843 & ~w1905;
assign w1908 = ~w1906 & w1907;
assign w1909 = ~w1904 & ~w1908;
assign w1910 = w1849 & ~w1909;
assign w1911 = ~pi031 & ~w1843;
assign w1912 = ~pi015 & w1843;
assign w1913 = ~w1911 & ~w1912;
assign w1914 = w1839 & w1913;
assign w1915 = ~pi044 & ~w1843;
assign w1916 = ~pi032 & w1843;
assign w1917 = ~w1915 & ~w1916;
assign w1918 = ~w1839 & w1917;
assign w1919 = ~w1849 & ~w1914;
assign w1920 = ~w1918 & w1919;
assign w1921 = w1834 & ~w1920;
assign w1922 = ~w1910 & w1921;
assign w1923 = (~pi011 & w1846) | (~pi011 & w3196) | (w1846 & w3196);
assign w1924 = ~pi013 & w1849;
assign w1925 = w1843 & ~w1923;
assign w1926 = ~w1924 & w1925;
assign w1927 = (~pi042 & w1846) | (~pi042 & w3197) | (w1846 & w3197);
assign w1928 = ~pi012 & w1849;
assign w1929 = ~w1843 & ~w1927;
assign w1930 = ~w1928 & w1929;
assign w1931 = ~w1926 & ~w1930;
assign w1932 = w1840 & ~w1931;
assign w1933 = ~pi043 & ~w1849;
assign w1934 = ~pi041 & w1849;
assign w1935 = w1843 & ~w1933;
assign w1936 = ~w1934 & w1935;
assign w1937 = ~pi040 & ~w1849;
assign w1938 = ~pi045 & w1849;
assign w1939 = ~w1843 & ~w1937;
assign w1940 = ~w1938 & w1939;
assign w1941 = ~w1936 & ~w1940;
assign w1942 = w1860 & ~w1941;
assign w1943 = w1875 & ~w1932;
assign w1944 = ~w1942 & w1943;
assign w1945 = ~w1922 & w1944;
assign w1946 = ~w1820 & w1828;
assign w1947 = ~w1900 & ~w1945;
assign w1948 = w1946 & w1947;
assign w1949 = ~w1838 & w3198;
assign w1950 = pi103 & ~w1839;
assign w1951 = ~w1849 & ~w1949;
assign w1952 = ~w1950 & w1951;
assign w1953 = ~w1838 & w3199;
assign w1954 = pi124 & ~w1839;
assign w1955 = w1849 & ~w1953;
assign w1956 = ~w1954 & w1955;
assign w1957 = ~w1952 & ~w1956;
assign w1958 = w1843 & ~w1957;
assign w1959 = (~pi105 & w1846) | (~pi105 & w3200) | (w1846 & w3200);
assign w1960 = ~w1846 & w3201;
assign w1961 = ~w1959 & ~w1960;
assign w1962 = w1839 & w1961;
assign w1963 = ~pi084 & ~w1849;
assign w1964 = ~pi117 & w1849;
assign w1965 = ~w1963 & ~w1964;
assign w1966 = ~w1839 & w1965;
assign w1967 = ~w1843 & ~w1962;
assign w1968 = ~w1966 & w1967;
assign w1969 = w1834 & ~w1968;
assign w1970 = ~w1958 & w1969;
assign w1971 = (~pi122 & w1846) | (~pi122 & w3202) | (w1846 & w3202);
assign w1972 = ~pi115 & w1849;
assign w1973 = w1843 & ~w1971;
assign w1974 = ~w1972 & w1973;
assign w1975 = (~pi116 & w1846) | (~pi116 & w3203) | (w1846 & w3203);
assign w1976 = ~pi123 & w1849;
assign w1977 = ~w1843 & ~w1975;
assign w1978 = ~w1976 & w1977;
assign w1979 = ~w1974 & ~w1978;
assign w1980 = w1840 & ~w1979;
assign w1981 = ~pi089 & ~w1849;
assign w1982 = ~pi119 & w1849;
assign w1983 = w1843 & ~w1981;
assign w1984 = ~w1982 & w1983;
assign w1985 = ~pi118 & ~w1849;
assign w1986 = ~pi096 & w1849;
assign w1987 = ~w1843 & ~w1985;
assign w1988 = ~w1986 & w1987;
assign w1989 = ~w1984 & ~w1988;
assign w1990 = w1860 & ~w1989;
assign w1991 = ~w1875 & ~w1980;
assign w1992 = ~w1990 & w1991;
assign w1993 = ~w1970 & w1992;
assign w1994 = ~w1838 & w3204;
assign w1995 = pi090 & ~w1839;
assign w1996 = w1843 & ~w1994;
assign w1997 = ~w1995 & w1996;
assign w1998 = ~w1838 & w3205;
assign w1999 = pi093 & ~w1839;
assign w2000 = ~w1843 & ~w1998;
assign w2001 = ~w1999 & w2000;
assign w2002 = ~w1997 & ~w2001;
assign w2003 = w1849 & ~w2002;
assign w2004 = ~pi095 & ~w1843;
assign w2005 = ~pi091 & w1843;
assign w2006 = ~w2004 & ~w2005;
assign w2007 = w1839 & w2006;
assign w2008 = ~pi102 & ~w1843;
assign w2009 = ~pi088 & w1843;
assign w2010 = ~w2008 & ~w2009;
assign w2011 = ~w1839 & w2010;
assign w2012 = ~w1849 & ~w2007;
assign w2013 = ~w2011 & w2012;
assign w2014 = w1834 & ~w2013;
assign w2015 = ~w2003 & w2014;
assign w2016 = (~pi127 & w1846) | (~pi127 & w3206) | (w1846 & w3206);
assign w2017 = ~pi087 & w1849;
assign w2018 = w1843 & ~w2016;
assign w2019 = ~w2017 & w2018;
assign w2020 = (~pi108 & w1846) | (~pi108 & w3207) | (w1846 & w3207);
assign w2021 = ~pi120 & w1849;
assign w2022 = ~w1843 & ~w2020;
assign w2023 = ~w2021 & w2022;
assign w2024 = ~w2019 & ~w2023;
assign w2025 = w1840 & ~w2024;
assign w2026 = ~pi104 & ~w1849;
assign w2027 = ~pi121 & w1849;
assign w2028 = w1843 & ~w2026;
assign w2029 = ~w2027 & w2028;
assign w2030 = ~pi086 & ~w1849;
assign w2031 = ~pi097 & w1849;
assign w2032 = ~w1843 & ~w2030;
assign w2033 = ~w2031 & w2032;
assign w2034 = ~w2029 & ~w2033;
assign w2035 = w1860 & ~w2034;
assign w2036 = w1875 & ~w2025;
assign w2037 = ~w2035 & w2036;
assign w2038 = ~w2015 & w2037;
assign w2039 = w1820 & w1828;
assign w2040 = ~w1993 & ~w2038;
assign w2041 = w2039 & w2040;
assign w2042 = (~pi106 & w1846) | (~pi106 & w3208) | (w1846 & w3208);
assign w2043 = ~pi000 & w1849;
assign w2044 = w1843 & ~w2042;
assign w2045 = ~w2043 & w2044;
assign w2046 = (~pi074 & w1846) | (~pi074 & w3209) | (w1846 & w3209);
assign w2047 = ~pi107 & w1849;
assign w2048 = ~w1843 & ~w2046;
assign w2049 = ~w2047 & w2048;
assign w2050 = ~w2045 & ~w2049;
assign w2051 = w1840 & ~w2050;
assign w2052 = ~pi071 & ~w1849;
assign w2053 = ~pi073 & w1849;
assign w2054 = w1843 & ~w2052;
assign w2055 = ~w2053 & w2054;
assign w2056 = ~pi003 & ~w1849;
assign w2057 = ~pi072 & w1849;
assign w2058 = ~w1843 & ~w2056;
assign w2059 = ~w2057 & w2058;
assign w2060 = ~w2055 & ~w2059;
assign w2061 = w1860 & ~w2060;
assign w2062 = ~pi101 & ~w1843;
assign w2063 = ~pi100 & w1843;
assign w2064 = ~w2062 & ~w2063;
assign w2065 = ~w1839 & w2064;
assign w2066 = ~pi112 & ~w1843;
assign w2067 = ~pi076 & w1843;
assign w2068 = ~w2066 & ~w2067;
assign w2069 = w1839 & w2068;
assign w2070 = ~w1849 & ~w2065;
assign w2071 = ~w2069 & w2070;
assign w2072 = ~pi077 & ~w1843;
assign w2073 = ~pi078 & w1843;
assign w2074 = ~w2072 & ~w2073;
assign w2075 = w1839 & w2074;
assign w2076 = ~pi109 & ~w1843;
assign w2077 = ~pi075 & w1843;
assign w2078 = ~w2076 & ~w2077;
assign w2079 = ~w1839 & w2078;
assign w2080 = w1849 & ~w2075;
assign w2081 = ~w2079 & w2080;
assign w2082 = w1834 & ~w2071;
assign w2083 = ~w2081 & w2082;
assign w2084 = ~w1875 & ~w2051;
assign w2085 = ~w2061 & w2084;
assign w2086 = ~w2083 & w2085;
assign w2087 = (~pi110 & w1846) | (~pi110 & w3210) | (w1846 & w3210);
assign w2088 = ~pi070 & w1849;
assign w2089 = w1843 & ~w2087;
assign w2090 = ~w2088 & w2089;
assign w2091 = (~pi099 & w1846) | (~pi099 & w3211) | (w1846 & w3211);
assign w2092 = ~pi111 & w1849;
assign w2093 = ~w1843 & ~w2091;
assign w2094 = ~w2092 & w2093;
assign w2095 = ~w2090 & ~w2094;
assign w2096 = w1860 & ~w2095;
assign w2097 = ~pi068 & ~w1849;
assign w2098 = ~pi114 & w1849;
assign w2099 = w1843 & ~w2097;
assign w2100 = ~w2098 & w2099;
assign w2101 = ~pi113 & ~w1849;
assign w2102 = ~pi069 & w1849;
assign w2103 = ~w1843 & ~w2101;
assign w2104 = ~w2102 & w2103;
assign w2105 = ~w2100 & ~w2104;
assign w2106 = w1840 & ~w2105;
assign w2107 = ~pi001 & ~w1843;
assign w2108 = ~pi079 & w1843;
assign w2109 = ~w2107 & ~w2108;
assign w2110 = ~w1839 & w2109;
assign w2111 = ~pi098 & ~w1843;
assign w2112 = ~pi082 & w1843;
assign w2113 = ~w2111 & ~w2112;
assign w2114 = w1839 & w2113;
assign w2115 = ~w1849 & ~w2110;
assign w2116 = ~w2114 & w2115;
assign w2117 = ~pi083 & ~w1843;
assign w2118 = ~pi002 & w1843;
assign w2119 = ~w2117 & ~w2118;
assign w2120 = w1839 & w2119;
assign w2121 = ~pi080 & ~w1843;
assign w2122 = ~pi081 & w1843;
assign w2123 = ~w2121 & ~w2122;
assign w2124 = ~w1839 & w2123;
assign w2125 = w1849 & ~w2120;
assign w2126 = ~w2124 & w2125;
assign w2127 = w1834 & ~w2116;
assign w2128 = ~w2126 & w2127;
assign w2129 = w1875 & ~w2096;
assign w2130 = ~w2106 & w2129;
assign w2131 = ~w2128 & w2130;
assign w2132 = w1820 & ~w1828;
assign w2133 = ~w2086 & ~w2131;
assign w2134 = w2132 & w2133;
assign w2135 = ~pi053 & ~w1843;
assign w2136 = ~pi052 & w1843;
assign w2137 = ~w2135 & ~w2136;
assign w2138 = w1839 & w2137;
assign w2139 = ~pi051 & ~w1843;
assign w2140 = ~pi059 & w1843;
assign w2141 = ~w2139 & ~w2140;
assign w2142 = ~w1839 & w2141;
assign w2143 = ~w1849 & ~w2138;
assign w2144 = ~w2142 & w2143;
assign w2145 = ~pi050 & ~w1839;
assign w2146 = ~pi055 & w1839;
assign w2147 = w1843 & ~w2145;
assign w2148 = ~w2146 & w2147;
assign w2149 = ~pi049 & ~w1839;
assign w2150 = ~pi054 & w1839;
assign w2151 = ~w1843 & ~w2149;
assign w2152 = ~w2150 & w2151;
assign w2153 = w1849 & ~w2148;
assign w2154 = ~w2152 & w2153;
assign w2155 = w1834 & ~w2144;
assign w2156 = ~w2154 & w2155;
assign w2157 = ~pi066 & ~w1849;
assign w2158 = ~pi030 & w1849;
assign w2159 = w1843 & ~w2157;
assign w2160 = ~w2158 & w2159;
assign w2161 = ~pi029 & ~w1849;
assign w2162 = ~pi067 & w1849;
assign w2163 = ~w1843 & ~w2161;
assign w2164 = ~w2162 & w2163;
assign w2165 = ~w2160 & ~w2164;
assign w2166 = w1840 & ~w2165;
assign w2167 = ~pi026 & ~w1849;
assign w2168 = ~pi065 & w1849;
assign w2169 = w1843 & ~w2167;
assign w2170 = ~w2168 & w2169;
assign w2171 = ~pi025 & ~w1849;
assign w2172 = ~pi027 & w1849;
assign w2173 = ~w1843 & ~w2171;
assign w2174 = ~w2172 & w2173;
assign w2175 = ~w2170 & ~w2174;
assign w2176 = w1860 & ~w2175;
assign w2177 = w1875 & ~w2166;
assign w2178 = ~w2176 & w2177;
assign w2179 = ~w2156 & w2178;
assign w2180 = ~pi022 & ~w1839;
assign w2181 = ~pi061 & w1839;
assign w2182 = ~w1849 & ~w2180;
assign w2183 = ~w2181 & w2182;
assign w2184 = ~pi056 & ~w1839;
assign w2185 = ~pi023 & w1839;
assign w2186 = w1849 & ~w2184;
assign w2187 = ~w2185 & w2186;
assign w2188 = ~w1843 & ~w2183;
assign w2189 = ~w2187 & w2188;
assign w2190 = ~pi063 & ~w1839;
assign w2191 = ~pi024 & w1839;
assign w2192 = w1849 & ~w2190;
assign w2193 = ~w2191 & w2192;
assign w2194 = ~pi064 & ~w1839;
assign w2195 = ~pi062 & w1839;
assign w2196 = ~w1849 & ~w2194;
assign w2197 = ~w2195 & w2196;
assign w2198 = w1843 & ~w2193;
assign w2199 = ~w2197 & w2198;
assign w2200 = w1834 & ~w2189;
assign w2201 = ~w2199 & w2200;
assign w2202 = ~pi058 & ~w1849;
assign w2203 = ~pi021 & w1849;
assign w2204 = w1843 & ~w2202;
assign w2205 = ~w2203 & w2204;
assign w2206 = ~pi020 & ~w1849;
assign w2207 = ~pi060 & w1849;
assign w2208 = ~w1843 & ~w2206;
assign w2209 = ~w2207 & w2208;
assign w2210 = ~w2205 & ~w2209;
assign w2211 = w1840 & ~w2210;
assign w2212 = ~pi028 & ~w1849;
assign w2213 = ~pi057 & w1849;
assign w2214 = w1843 & ~w2212;
assign w2215 = ~w2213 & w2214;
assign w2216 = ~pi018 & ~w1849;
assign w2217 = ~pi019 & w1849;
assign w2218 = ~w1843 & ~w2216;
assign w2219 = ~w2217 & w2218;
assign w2220 = ~w2215 & ~w2219;
assign w2221 = w1860 & ~w2220;
assign w2222 = ~w1875 & ~w2211;
assign w2223 = ~w2221 & w2222;
assign w2224 = ~w2201 & w2223;
assign w2225 = ~w1820 & ~w1828;
assign w2226 = ~w2179 & w2225;
assign w2227 = ~w2224 & w2226;
assign w2228 = ~w1804 & ~w1948;
assign w2229 = ~w2041 & ~w2134;
assign w2230 = w2228 & w2229;
assign w2231 = ~w2227 & w2230;
assign w2232 = ~w1805 & ~w2231;
assign w2233 = ~pi165 & ~pi170;
assign w2234 = ~pi162 & ~pi164;
assign w2235 = ~pi166 & ~pi167;
assign w2236 = ~pi168 & ~pi186;
assign w2237 = w2235 & w2236;
assign w2238 = w2234 & w2237;
assign w2239 = w2233 & w2238;
assign w2240 = ~pi191 & w2239;
assign w2241 = ~pi169 & w2240;
assign w2242 = ~pi159 & w2241;
assign w2243 = ~pi141 & w2242;
assign w2244 = ~pi154 & w2243;
assign w2245 = ~pi149 & w2244;
assign w2246 = ~pi147 & w2245;
assign w2247 = ~pi132 & w2246;
assign w2248 = pi136 & w2247;
assign w2249 = pi129 & ~w2248;
assign w2250 = ~pi129 & pi136;
assign w2251 = ~w344 & w2250;
assign w2252 = w2247 & w2251;
assign w2253 = ~w2249 & ~w2252;
assign w2254 = pi145 & w61;
assign w2255 = ~pi148 & w2254;
assign w2256 = ~pi142 & w2255;
assign w2257 = ~pi139 & w2256;
assign w2258 = ~pi140 & w2257;
assign w2259 = ~pi133 & w2258;
assign w2260 = ~pi130 & w2259;
assign w2261 = pi136 & ~w2260;
assign w2262 = pi130 & ~w2259;
assign w2263 = w2261 & ~w2262;
assign w2264 = ~pi150 & ~pi156;
assign w2265 = ~pi161 & ~pi171;
assign w2266 = ~pi176 & ~pi177;
assign w2267 = ~pi178 & w2266;
assign w2268 = w2264 & w2265;
assign w2269 = w2267 & w2268;
assign w2270 = ~pi136 & ~w2269;
assign w2271 = ~w2263 & ~w2270;
assign w2272 = ~pi235 & pi237;
assign w2273 = ~pi236 & w2272;
assign w2274 = w159 & w2273;
assign w2275 = pi136 & w2260;
assign w2276 = ~pi131 & ~w2275;
assign w2277 = ~w2274 & ~w2276;
assign w2278 = ~pi131 & ~pi271;
assign w2279 = ~w790 & ~w2278;
assign w2280 = w2274 & w2279;
assign w2281 = ~w2277 & ~w2280;
assign w2282 = pi136 & ~w2247;
assign w2283 = pi157 & ~w2282;
assign w2284 = pi136 & ~w2246;
assign w2285 = pi132 & w2284;
assign w2286 = ~w2283 & ~w2285;
assign w2287 = ~pi136 & ~pi178;
assign w2288 = pi133 & ~w2258;
assign w2289 = pi136 & ~w2259;
assign w2290 = ~w2288 & w2289;
assign w2291 = ~w2287 & ~w2290;
assign w2292 = pi134 & ~pi228;
assign w2293 = ~pi151 & w2275;
assign w2294 = ~w2292 & ~w2293;
assign w2295 = pi236 & w173;
assign w2296 = pi038 & w2295;
assign w2297 = pi100 & w170;
assign w2298 = pi103 & w161;
assign w2299 = pi138 & w2273;
assign w2300 = ~pi236 & w173;
assign w2301 = pi064 & w2300;
assign w2302 = pi237 & w169;
assign w2303 = pi185 & w2302;
assign w2304 = ~w2296 & ~w2297;
assign w2305 = ~w2298 & ~w2299;
assign w2306 = ~w2301 & ~w2303;
assign w2307 = w2305 & w2306;
assign w2308 = w2304 & w2307;
assign w2309 = ~pi131 & ~pi136;
assign w2310 = ~w2261 & ~w2309;
assign w2311 = pi143 & w2273;
assign w2312 = pi124 & w161;
assign w2313 = pi075 & w170;
assign w2314 = pi009 & w2295;
assign w2315 = pi063 & w2300;
assign w2316 = pi153 & w2302;
assign w2317 = ~w2311 & ~w2312;
assign w2318 = ~w2313 & ~w2314;
assign w2319 = ~w2315 & ~w2316;
assign w2320 = w2318 & w2319;
assign w2321 = w2317 & w2320;
assign w2322 = pi271 & w2274;
assign w2323 = pi138 & ~w2322;
assign w2324 = w962 & w2274;
assign w2325 = ~w2323 & ~w2324;
assign w2326 = pi139 & ~w2256;
assign w2327 = ~w2257 & ~w2326;
assign w2328 = pi136 & ~w2327;
assign w2329 = ~pi136 & pi177;
assign w2330 = ~w2328 & ~w2329;
assign w2331 = ~pi136 & ~pi161;
assign w2332 = pi140 & ~w2257;
assign w2333 = pi136 & ~w2258;
assign w2334 = ~w2332 & w2333;
assign w2335 = ~w2331 & ~w2334;
assign w2336 = pi141 & ~w2242;
assign w2337 = ~w2243 & ~w2336;
assign w2338 = w2282 & ~w2337;
assign w2339 = pi153 & ~w2282;
assign w2340 = ~w2338 & ~w2339;
assign w2341 = ~pi136 & ~pi176;
assign w2342 = pi142 & ~w2255;
assign w2343 = pi136 & ~w2256;
assign w2344 = ~w2342 & w2343;
assign w2345 = ~w2341 & ~w2344;
assign w2346 = pi143 & ~w2322;
assign w2347 = w629 & w2274;
assign w2348 = ~w2346 & ~w2347;
assign w2349 = pi144 & ~w2322;
assign w2350 = w617 & w2274;
assign w2351 = ~w2349 & ~w2350;
assign w2352 = ~pi129 & ~w2309;
assign w2353 = ~pi153 & ~pi155;
assign w2354 = ~pi157 & ~pi160;
assign w2355 = ~pi163 & ~pi172;
assign w2356 = ~pi173 & ~pi174;
assign w2357 = ~pi175 & ~pi179;
assign w2358 = ~pi180 & ~pi181;
assign w2359 = ~pi182 & ~pi183;
assign w2360 = ~pi184 & ~pi185;
assign w2361 = w2359 & w2360;
assign w2362 = w2357 & w2358;
assign w2363 = w2355 & w2356;
assign w2364 = w2353 & w2354;
assign w2365 = w2363 & w2364;
assign w2366 = w2361 & w2362;
assign w2367 = w2365 & w2366;
assign w2368 = ~w2352 & w2367;
assign w2369 = ~pi132 & ~pi141;
assign w2370 = ~pi147 & ~pi149;
assign w2371 = ~pi154 & ~pi159;
assign w2372 = pi165 & ~pi169;
assign w2373 = ~pi170 & ~pi191;
assign w2374 = w2372 & w2373;
assign w2375 = w2370 & w2371;
assign w2376 = w2369 & w2375;
assign w2377 = w2374 & w2376;
assign w2378 = w2238 & w2377;
assign w2379 = w2250 & w2378;
assign w2380 = ~w2368 & ~w2379;
assign w2381 = w2250 & w2367;
assign w2382 = pi129 & pi136;
assign w2383 = w2378 & w2382;
assign w2384 = ~w2381 & ~w2383;
assign w2385 = pi147 & ~w2245;
assign w2386 = w2284 & ~w2385;
assign w2387 = ~pi180 & ~w2282;
assign w2388 = ~w2386 & ~w2387;
assign w2389 = ~pi136 & ~pi156;
assign w2390 = pi148 & ~w2254;
assign w2391 = pi136 & ~w2255;
assign w2392 = ~w2390 & w2391;
assign w2393 = ~w2389 & ~w2392;
assign w2394 = pi149 & ~w2244;
assign w2395 = ~w2245 & ~w2394;
assign w2396 = w2282 & ~w2395;
assign w2397 = pi163 & ~w2282;
assign w2398 = ~w2396 & ~w2397;
assign w2399 = w549 & w2274;
assign w2400 = ~pi150 & ~w2399;
assign w2401 = ~pi151 & ~w2322;
assign w2402 = w641 & w2274;
assign w2403 = ~w2401 & ~w2402;
assign w2404 = ~pi152 & ~w2322;
assign w2405 = w973 & w2274;
assign w2406 = ~w2404 & ~w2405;
assign w2407 = w159 & w2302;
assign w2408 = pi271 & w2407;
assign w2409 = pi153 & ~w2408;
assign w2410 = w629 & w2407;
assign w2411 = ~w2409 & ~w2410;
assign w2412 = ~pi172 & ~w2282;
assign w2413 = pi154 & ~w2243;
assign w2414 = pi136 & ~w2244;
assign w2415 = ~w2413 & w2414;
assign w2416 = ~w2412 & ~w2415;
assign w2417 = pi270 & w2407;
assign w2418 = pi155 & ~w2417;
assign w2419 = w592 & w2407;
assign w2420 = ~w2418 & ~w2419;
assign w2421 = pi270 & w2274;
assign w2422 = pi156 & ~w2421;
assign w2423 = w580 & w2274;
assign w2424 = ~w2422 & ~w2423;
assign w2425 = pi157 & ~w2408;
assign w2426 = w812 & w2407;
assign w2427 = ~w2425 & ~w2426;
assign w2428 = ~pi158 & ~w2421;
assign w2429 = w177 & w2274;
assign w2430 = ~w2428 & ~w2429;
assign w2431 = pi159 & ~w2241;
assign w2432 = ~w2242 & ~w2431;
assign w2433 = w2282 & ~w2432;
assign w2434 = pi173 & ~w2282;
assign w2435 = ~w2433 & ~w2434;
assign w2436 = pi160 & ~w2408;
assign w2437 = w790 & w2407;
assign w2438 = ~w2436 & ~w2437;
assign w2439 = pi161 & ~w2421;
assign w2440 = w929 & w2274;
assign w2441 = ~w2439 & ~w2440;
assign w2442 = ~pi166 & w2233;
assign w2443 = ~pi162 & w2442;
assign w2444 = pi162 & ~w2442;
assign w2445 = ~w2443 & ~w2444;
assign w2446 = w2282 & ~w2445;
assign w2447 = pi181 & ~w2282;
assign w2448 = ~w2446 & ~w2447;
assign w2449 = pi163 & ~w2408;
assign w2450 = w973 & w2407;
assign w2451 = ~w2449 & ~w2450;
assign w2452 = ~pi186 & w2443;
assign w2453 = pi164 & ~w2452;
assign w2454 = ~pi164 & w2452;
assign w2455 = ~w2453 & ~w2454;
assign w2456 = w2282 & ~w2455;
assign w2457 = pi182 & ~w2282;
assign w2458 = ~w2456 & ~w2457;
assign w2459 = pi136 & pi165;
assign w2460 = ~pi179 & ~w2282;
assign w2461 = ~w2459 & ~w2460;
assign w2462 = pi166 & ~w2233;
assign w2463 = ~w2442 & ~w2462;
assign w2464 = w2282 & ~w2463;
assign w2465 = pi175 & ~w2282;
assign w2466 = ~w2464 & ~w2465;
assign w2467 = ~pi184 & ~w2282;
assign w2468 = ~pi168 & w2454;
assign w2469 = pi167 & ~w2468;
assign w2470 = ~w2239 & ~w2469;
assign w2471 = w2282 & w2470;
assign w2472 = ~w2467 & ~w2471;
assign w2473 = pi168 & ~w2454;
assign w2474 = ~w2468 & ~w2473;
assign w2475 = w2282 & ~w2474;
assign w2476 = pi183 & ~w2282;
assign w2477 = ~w2475 & ~w2476;
assign w2478 = ~pi185 & ~w2282;
assign w2479 = pi169 & ~w2240;
assign w2480 = pi136 & ~w2241;
assign w2481 = ~w2479 & w2480;
assign w2482 = ~w2478 & ~w2481;
assign w2483 = ~pi174 & ~w2282;
assign w2484 = pi165 & pi170;
assign w2485 = pi136 & ~w2233;
assign w2486 = ~w2484 & w2485;
assign w2487 = ~w2483 & ~w2486;
assign w2488 = pi171 & ~w2421;
assign w2489 = w562 & w2274;
assign w2490 = ~w2488 & ~w2489;
assign w2491 = pi172 & ~w2408;
assign w2492 = w641 & w2407;
assign w2493 = ~w2491 & ~w2492;
assign w2494 = pi173 & ~w2408;
assign w2495 = w617 & w2407;
assign w2496 = ~w2494 & ~w2495;
assign w2497 = pi174 & ~w2417;
assign w2498 = w562 & w2407;
assign w2499 = ~w2497 & ~w2498;
assign w2500 = pi175 & ~w2417;
assign w2501 = w580 & w2407;
assign w2502 = ~w2500 & ~w2501;
assign w2503 = pi176 & ~w2421;
assign w2504 = w918 & w2274;
assign w2505 = ~w2503 & ~w2504;
assign w2506 = pi177 & ~w2421;
assign w2507 = w592 & w2274;
assign w2508 = ~w2506 & ~w2507;
assign w2509 = pi178 & ~w2421;
assign w2510 = w938 & w2274;
assign w2511 = ~w2509 & ~w2510;
assign w2512 = pi179 & ~w2417;
assign w2513 = w549 & w2407;
assign w2514 = ~w2512 & ~w2513;
assign w2515 = pi180 & ~w2408;
assign w2516 = w1066 & w2407;
assign w2517 = ~w2515 & ~w2516;
assign w2518 = pi181 & ~w2417;
assign w2519 = w918 & w2407;
assign w2520 = ~w2518 & ~w2519;
assign w2521 = pi182 & ~w2417;
assign w2522 = w929 & w2407;
assign w2523 = ~w2521 & ~w2522;
assign w2524 = pi183 & ~w2417;
assign w2525 = w938 & w2407;
assign w2526 = ~w2524 & ~w2525;
assign w2527 = pi184 & ~w2417;
assign w2528 = w177 & w2407;
assign w2529 = ~w2527 & ~w2528;
assign w2530 = pi185 & ~w2408;
assign w2531 = w962 & w2407;
assign w2532 = ~w2530 & ~w2531;
assign w2533 = pi186 & ~w2443;
assign w2534 = ~w2452 & ~w2533;
assign w2535 = w2282 & ~w2534;
assign w2536 = pi155 & ~w2282;
assign w2537 = ~w2535 & ~w2536;
assign w2538 = pi145 & ~pi190;
assign w2539 = pi187 & ~w2538;
assign w2540 = ~w2254 & ~w2539;
assign w2541 = pi136 & ~w2540;
assign w2542 = ~pi136 & pi171;
assign w2543 = ~w2541 & ~w2542;
assign w2544 = pi236 & w2272;
assign w2545 = ~pi195 & w2544;
assign w2546 = pi021 & w2300;
assign w2547 = ~pi158 & w2273;
assign w2548 = pi115 & w161;
assign w2549 = pi184 & w2302;
assign w2550 = pi000 & w170;
assign w2551 = pi007 & w2295;
assign w2552 = ~w2545 & ~w2546;
assign w2553 = ~w2547 & ~w2548;
assign w2554 = ~w2549 & ~w2550;
assign w2555 = ~w2551 & w2554;
assign w2556 = w2552 & w2553;
assign w2557 = w2555 & w2556;
assign w2558 = pi073 & w170;
assign w2559 = pi057 & w2300;
assign w2560 = pi034 & w2295;
assign w2561 = pi119 & w161;
assign w2562 = pi176 & w2273;
assign w2563 = ~pi193 & w2544;
assign w2564 = pi181 & w2302;
assign w2565 = ~w2558 & ~w2559;
assign w2566 = ~w2560 & ~w2561;
assign w2567 = ~w2562 & ~w2563;
assign w2568 = ~w2564 & w2567;
assign w2569 = w2565 & w2566;
assign w2570 = w2568 & w2569;
assign w2571 = ~pi145 & pi190;
assign w2572 = ~w2538 & ~w2571;
assign w2573 = pi136 & ~w2572;
assign w2574 = ~pi136 & pi150;
assign w2575 = ~w2573 & ~w2574;
assign w2576 = pi191 & ~w2239;
assign w2577 = ~w2240 & ~w2576;
assign w2578 = w2282 & ~w2577;
assign w2579 = pi160 & ~w2282;
assign w2580 = ~w2578 & ~w2579;
assign w2581 = w159 & w2544;
assign w2582 = pi270 & w2581;
assign w2583 = ~pi192 & ~w2582;
assign w2584 = w929 & w2581;
assign w2585 = ~w2583 & ~w2584;
assign w2586 = ~pi193 & ~w2582;
assign w2587 = w918 & w2581;
assign w2588 = ~w2586 & ~w2587;
assign w2589 = ~pi194 & ~w2582;
assign w2590 = w562 & w2581;
assign w2591 = ~w2589 & ~w2590;
assign w2592 = ~pi195 & ~w2582;
assign w2593 = w177 & w2581;
assign w2594 = ~w2592 & ~w2593;
assign w2595 = ~pi196 & ~w2582;
assign w2596 = w549 & w2581;
assign w2597 = ~w2595 & ~w2596;
assign w2598 = ~pi197 & ~w2582;
assign w2599 = w580 & w2581;
assign w2600 = ~w2598 & ~w2599;
assign w2601 = ~pi198 & ~w2582;
assign w2602 = w592 & w2581;
assign w2603 = ~w2601 & ~w2602;
assign w2604 = ~pi199 & ~w2582;
assign w2605 = w938 & w2581;
assign w2606 = ~w2604 & ~w2605;
assign w2607 = pi020 & w2300;
assign w2608 = pi006 & w2295;
assign w2609 = pi177 & w2273;
assign w2610 = pi116 & w161;
assign w2611 = pi074 & w170;
assign w2612 = ~pi198 & w2544;
assign w2613 = pi155 & w2302;
assign w2614 = ~w2607 & ~w2608;
assign w2615 = ~w2609 & ~w2610;
assign w2616 = ~w2611 & ~w2612;
assign w2617 = ~w2613 & w2616;
assign w2618 = w2614 & w2615;
assign w2619 = w2617 & w2618;
assign w2620 = pi058 & w2300;
assign w2621 = pi035 & w2295;
assign w2622 = ~pi192 & w2544;
assign w2623 = pi182 & w2302;
assign w2624 = pi161 & w2273;
assign w2625 = pi122 & w161;
assign w2626 = pi106 & w170;
assign w2627 = ~w2620 & ~w2621;
assign w2628 = ~w2622 & ~w2623;
assign w2629 = ~w2624 & ~w2625;
assign w2630 = ~w2626 & w2629;
assign w2631 = w2627 & w2628;
assign w2632 = w2630 & w2631;
assign w2633 = pi033 & w2295;
assign w2634 = pi003 & w170;
assign w2635 = pi118 & w161;
assign w2636 = pi018 & w2300;
assign w2637 = pi179 & w2302;
assign w2638 = ~pi196 & w2544;
assign w2639 = pi150 & w2273;
assign w2640 = ~w2633 & ~w2634;
assign w2641 = ~w2635 & ~w2636;
assign w2642 = ~w2637 & ~w2638;
assign w2643 = ~w2639 & w2642;
assign w2644 = w2640 & w2641;
assign w2645 = w2643 & w2644;
assign w2646 = pi174 & w2302;
assign w2647 = pi089 & w161;
assign w2648 = pi028 & w2300;
assign w2649 = pi071 & w170;
assign w2650 = pi171 & w2273;
assign w2651 = ~pi194 & w2544;
assign w2652 = pi004 & w2295;
assign w2653 = ~w2646 & ~w2647;
assign w2654 = ~w2648 & ~w2649;
assign w2655 = ~w2650 & ~w2651;
assign w2656 = ~w2652 & w2655;
assign w2657 = w2653 & w2654;
assign w2658 = w2656 & w2657;
assign w2659 = pi183 & w2302;
assign w2660 = ~pi199 & w2544;
assign w2661 = pi178 & w2273;
assign w2662 = pi036 & w2295;
assign w2663 = pi107 & w170;
assign w2664 = pi123 & w161;
assign w2665 = pi060 & w2300;
assign w2666 = ~w2659 & ~w2660;
assign w2667 = ~w2661 & ~w2662;
assign w2668 = ~w2663 & ~w2664;
assign w2669 = ~w2665 & w2668;
assign w2670 = w2666 & w2667;
assign w2671 = w2669 & w2670;
assign w2672 = pi096 & w161;
assign w2673 = ~pi197 & w2544;
assign w2674 = pi072 & w170;
assign w2675 = pi005 & w2295;
assign w2676 = pi019 & w2300;
assign w2677 = pi175 & w2302;
assign w2678 = pi156 & w2273;
assign w2679 = ~w2672 & ~w2673;
assign w2680 = ~w2674 & ~w2675;
assign w2681 = ~w2676 & ~w2677;
assign w2682 = ~w2678 & w2681;
assign w2683 = w2679 & w2680;
assign w2684 = w2682 & w2683;
assign w2685 = pi144 & w2273;
assign w2686 = pi117 & w161;
assign w2687 = pi109 & w170;
assign w2688 = pi008 & w2295;
assign w2689 = pi056 & w2300;
assign w2690 = pi173 & w2302;
assign w2691 = ~w2685 & ~w2686;
assign w2692 = ~w2687 & ~w2688;
assign w2693 = ~w2689 & ~w2690;
assign w2694 = w2692 & w2693;
assign w2695 = w2691 & w2694;
assign w2696 = pi125 & w161;
assign w2697 = pi062 & w2300;
assign w2698 = pi076 & w170;
assign w2699 = pi039 & w2295;
assign w2700 = pi163 & w2302;
assign w2701 = ~pi152 & w2273;
assign w2702 = ~w2696 & ~w2697;
assign w2703 = ~w2698 & ~w2699;
assign w2704 = ~w2700 & ~w2701;
assign w2705 = w2703 & w2704;
assign w2706 = w2702 & w2705;
assign w2707 = pi048 & w2295;
assign w2708 = pi126 & w161;
assign w2709 = pi077 & w170;
assign w2710 = pi180 & w2302;
assign w2711 = pi023 & w2300;
assign w2712 = ~w2707 & ~w2708;
assign w2713 = ~w2709 & ~w2710;
assign w2714 = ~w2711 & w2713;
assign w2715 = w2712 & w2714;
assign w2716 = pi105 & w161;
assign w2717 = pi112 & w170;
assign w2718 = pi172 & w2302;
assign w2719 = ~pi151 & w2273;
assign w2720 = pi061 & w2300;
assign w2721 = pi010 & w2295;
assign w2722 = ~w2716 & ~w2717;
assign w2723 = ~w2718 & ~w2719;
assign w2724 = ~w2720 & ~w2721;
assign w2725 = w2723 & w2724;
assign w2726 = w2722 & w2725;
assign w2727 = pi084 & w161;
assign w2728 = ~pi131 & w2273;
assign w2729 = pi037 & w2295;
assign w2730 = pi101 & w170;
assign w2731 = pi160 & w2302;
assign w2732 = pi022 & w2300;
assign w2733 = ~w2727 & ~w2728;
assign w2734 = ~w2729 & ~w2730;
assign w2735 = ~w2731 & ~w2732;
assign w2736 = w2734 & w2735;
assign w2737 = w2733 & w2736;
assign w2738 = pi047 & w2295;
assign w2739 = pi078 & w170;
assign w2740 = pi157 & w2302;
assign w2741 = pi085 & w161;
assign w2742 = pi024 & w2300;
assign w2743 = ~w2738 & ~w2739;
assign w2744 = ~w2740 & ~w2741;
assign w2745 = ~w2742 & w2744;
assign w2746 = w2743 & w2745;
assign w2747 = pi080 & w170;
assign w2748 = pi049 & w2300;
assign w2749 = pi046 & w2295;
assign w2750 = pi093 & w161;
assign w2751 = ~w2747 & ~w2748;
assign w2752 = ~w2749 & ~w2750;
assign w2753 = w2751 & w2752;
assign w2754 = pi086 & w161;
assign w2755 = pi040 & w2295;
assign w2756 = pi099 & w170;
assign w2757 = pi025 & w2300;
assign w2758 = ~w2754 & ~w2755;
assign w2759 = ~w2756 & ~w2757;
assign w2760 = w2758 & w2759;
assign w2761 = pi097 & w161;
assign w2762 = pi111 & w170;
assign w2763 = pi027 & w2300;
assign w2764 = pi045 & w2295;
assign w2765 = ~w2761 & ~w2762;
assign w2766 = ~w2763 & ~w2764;
assign w2767 = w2765 & w2766;
assign w2768 = pi110 & w170;
assign w2769 = pi026 & w2300;
assign w2770 = pi043 & w2295;
assign w2771 = pi104 & w161;
assign w2772 = ~w2768 & ~w2769;
assign w2773 = ~w2770 & ~w2771;
assign w2774 = w2772 & w2773;
assign w2775 = pi070 & w170;
assign w2776 = pi041 & w2295;
assign w2777 = pi065 & w2300;
assign w2778 = pi121 & w161;
assign w2779 = ~w2775 & ~w2776;
assign w2780 = ~w2777 & ~w2778;
assign w2781 = w2779 & w2780;
assign w2782 = pi067 & w2300;
assign w2783 = pi120 & w161;
assign w2784 = pi012 & w2295;
assign w2785 = pi069 & w170;
assign w2786 = ~w2782 & ~w2783;
assign w2787 = ~w2784 & ~w2785;
assign w2788 = w2786 & w2787;
assign w2789 = pi050 & w2300;
assign w2790 = pi081 & w170;
assign w2791 = pi090 & w161;
assign w2792 = pi014 & w2295;
assign w2793 = ~w2789 & ~w2790;
assign w2794 = ~w2791 & ~w2792;
assign w2795 = w2793 & w2794;
assign w2796 = pi011 & w2295;
assign w2797 = pi127 & w161;
assign w2798 = pi068 & w170;
assign w2799 = pi066 & w2300;
assign w2800 = ~w2796 & ~w2797;
assign w2801 = ~w2798 & ~w2799;
assign w2802 = w2800 & w2801;
assign w2803 = pi094 & w161;
assign w2804 = pi017 & w2295;
assign w2805 = pi055 & w2300;
assign w2806 = pi002 & w170;
assign w2807 = ~w2803 & ~w2804;
assign w2808 = ~w2805 & ~w2806;
assign w2809 = w2807 & w2808;
assign w2810 = pi031 & w2295;
assign w2811 = pi098 & w170;
assign w2812 = pi053 & w2300;
assign w2813 = pi095 & w161;
assign w2814 = ~w2810 & ~w2811;
assign w2815 = ~w2812 & ~w2813;
assign w2816 = w2814 & w2815;
assign w2817 = pi044 & w2295;
assign w2818 = pi102 & w161;
assign w2819 = pi001 & w170;
assign w2820 = pi051 & w2300;
assign w2821 = ~w2817 & ~w2818;
assign w2822 = ~w2819 & ~w2820;
assign w2823 = w2821 & w2822;
assign w2824 = pi087 & w161;
assign w2825 = pi013 & w2295;
assign w2826 = pi114 & w170;
assign w2827 = pi030 & w2300;
assign w2828 = ~w2824 & ~w2825;
assign w2829 = ~w2826 & ~w2827;
assign w2830 = w2828 & w2829;
assign w2831 = pi016 & w2295;
assign w2832 = pi092 & w161;
assign w2833 = pi054 & w2300;
assign w2834 = pi083 & w170;
assign w2835 = ~w2831 & ~w2832;
assign w2836 = ~w2833 & ~w2834;
assign w2837 = w2835 & w2836;
assign w2838 = pi108 & w161;
assign w2839 = pi042 & w2295;
assign w2840 = pi113 & w170;
assign w2841 = pi029 & w2300;
assign w2842 = ~w2838 & ~w2839;
assign w2843 = ~w2840 & ~w2841;
assign w2844 = w2842 & w2843;
assign w2845 = pi015 & w2295;
assign w2846 = pi091 & w161;
assign w2847 = pi052 & w2300;
assign w2848 = pi082 & w170;
assign w2849 = ~w2845 & ~w2846;
assign w2850 = ~w2847 & ~w2848;
assign w2851 = w2849 & w2850;
assign w2852 = pi088 & w161;
assign w2853 = pi079 & w170;
assign w2854 = pi059 & w2300;
assign w2855 = pi032 & w2295;
assign w2856 = ~w2852 & ~w2853;
assign w2857 = ~w2854 & ~w2855;
assign w2858 = w2856 & w2857;
assign w2859 = ~pi228 & w157;
assign w2860 = ~pi187 & ~pi148;
assign w2861 = ~w21 & ~w47;
assign w2862 = ~w57 & pi143;
assign w2863 = ~pi148 & ~pi142;
assign w2864 = w13 & pi143;
assign w2865 = w71 & w75;
assign w2866 = pi138 & ~pi143;
assign w2867 = pi142 & pi139;
assign w2868 = ~w57 & ~w96;
assign w2869 = w72 & ~w15;
assign w2870 = ~w135 & pi110;
assign w2871 = w139 & w135;
assign w2872 = ~w135 & pi070;
assign w2873 = ~w135 & pi114;
assign w2874 = ~w135 & pi068;
assign w2875 = ~w135 & pi079;
assign w2876 = ~w135 & pi081;
assign w2877 = ~w135 & pi106;
assign w2878 = ~w135 & pi000;
assign w2879 = ~w135 & pi073;
assign w2880 = ~w135 & pi071;
assign w2881 = ~w135 & pi050;
assign w2882 = ~w135 & pi059;
assign w2883 = ~w135 & pi065;
assign w2884 = ~w135 & pi026;
assign w2885 = ~w135 & pi030;
assign w2886 = ~w135 & pi066;
assign w2887 = ~w135 & pi055;
assign w2888 = ~w135 & pi052;
assign w2889 = w76 & ~w69;
assign w2890 = ~w135 & ~pi017;
assign w2891 = ~w135 & ~pi032;
assign w2892 = ~w135 & ~pi014;
assign w2893 = ~w135 & ~pi041;
assign w2894 = ~w135 & ~pi011;
assign w2895 = ~w135 & ~pi013;
assign w2896 = ~w135 & ~pi047;
assign w2897 = ~w135 & ~pi009;
assign w2898 = ~w135 & ~pi038;
assign w2899 = ~w135 & pi034;
assign w2900 = ~w135 & pi007;
assign w2901 = ~w135 & pi035;
assign w2902 = ~w350 & ~w347;
assign w2903 = ~w135 & ~pi091;
assign w2904 = ~w135 & ~pi094;
assign w2905 = ~w135 & pi085;
assign w2906 = ~w135 & pi125;
assign w2907 = ~w135 & pi103;
assign w2908 = ~w135 & ~pi127;
assign w2909 = ~w135 & ~pi087;
assign w2910 = ~w135 & ~pi104;
assign w2911 = ~w135 & ~pi121;
assign w2912 = ~w135 & ~pi122;
assign w2913 = ~w135 & ~pi115;
assign w2914 = ~w135 & ~pi089;
assign w2915 = ~w135 & ~pi119;
assign w2916 = ~w508 & ~w509;
assign w2917 = ~w1810 & ~w32;
assign w2918 = ~w152 & ~w151;
assign w2919 = ~w152 & pi143;
assign w2920 = ~w1810 & pi143;
assign w2921 = pi156 & pi143;
assign w2922 = ~w72 & ~w71;
assign w2923 = w69 & w85;
assign w2924 = ~w93 & ~w91;
assign w2925 = ~w69 & w85;
assign w2926 = ~w135 & ~pi043;
assign w2927 = w69 & ~w85;
assign w2928 = ~w135 & ~pi039;
assign w2929 = ~w135 & pi004;
assign w2930 = ~w135 & ~pi090;
assign w2931 = ~w135 & pi124;
assign w2932 = w510 & ~w509;
assign w2933 = w510 & w340;
assign w2934 = w526 & ~w509;
assign w2935 = w526 & w340;
assign w2936 = w542 & ~w509;
assign w2937 = w542 & w340;
assign w2938 = w553 & ~w509;
assign w2939 = w553 & w340;
assign w2940 = w570 & ~w509;
assign w2941 = w570 & w340;
assign w2942 = w576 & w3212;
assign w2943 = w584 & w340;
assign w2944 = w588 & w3213;
assign w2945 = w596 & w340;
assign w2946 = w606 & ~w509;
assign w2947 = w606 & w340;
assign w2948 = w611 & w3214;
assign w2949 = w621 & w340;
assign w2950 = w625 & w3215;
assign w2951 = w633 & w340;
assign w2952 = w637 & w3216;
assign w2953 = w645 & w340;
assign w2954 = w661 & ~w509;
assign w2955 = w661 & w340;
assign w2956 = w666 & w3217;
assign w2957 = w674 & w340;
assign w2958 = w685 & ~w509;
assign w2959 = w685 & w340;
assign w2960 = w695 & w3218;
assign w2961 = w696 & w340;
assign w2962 = w706 & w3219;
assign w2963 = w707 & w340;
assign w2964 = w713 & w3220;
assign w2965 = w721 & w340;
assign w2966 = w727 & w3221;
assign w2967 = w728 & w340;
assign w2968 = w747 & w509;
assign w2969 = (w747 & w302) | (w747 & w3262) | (w302 & w3262);
assign w2970 = w757 & w3222;
assign w2971 = w759 & ~w340;
assign w2972 = w757 & w3223;
assign w2973 = w770 & ~w340;
assign w2974 = w774 & w509;
assign w2975 = (w774 & w302) | (w774 & w3263) | (w302 & w3263);
assign w2976 = w796 & w509;
assign w2977 = (w796 & w302) | (w796 & w3264) | (w302 & w3264);
assign w2978 = w800 & w509;
assign w2979 = (w800 & w302) | (w800 & w3265) | (w302 & w3265);
assign w2980 = w817 & w509;
assign w2981 = (w817 & w302) | (w817 & w3266) | (w302 & w3266);
assign w2982 = w831 & w509;
assign w2983 = w831 & ~w340;
assign w2984 = w835 & w509;
assign w2985 = (w835 & w302) | (w835 & w3267) | (w302 & w3267);
assign w2986 = w844 & w509;
assign w2987 = (w844 & w302) | (w844 & w3268) | (w302 & w3268);
assign w2988 = w859 & w509;
assign w2989 = (w859 & w302) | (w859 & w3269) | (w302 & w3269);
assign w2990 = w863 & w509;
assign w2991 = (w863 & w302) | (w863 & w3270) | (w302 & w3270);
assign w2992 = w878 & w509;
assign w2993 = w878 & ~w340;
assign w2994 = w885 & w3224;
assign w2995 = w886 & w340;
assign w2996 = w896 & w3225;
assign w2997 = w897 & w340;
assign w2998 = w910 & ~w509;
assign w2999 = w910 & w340;
assign w3000 = w922 & ~w509;
assign w3001 = w922 & w340;
assign w3002 = w933 & ~w509;
assign w3003 = w933 & w340;
assign w3004 = w936 & w3226;
assign w3005 = w941 & w340;
assign w3006 = w948 & w3227;
assign w3007 = w955 & w340;
assign w3008 = w958 & w3228;
assign w3009 = w966 & w340;
assign w3010 = w969 & w3229;
assign w3011 = w977 & w340;
assign w3012 = w987 & ~w509;
assign w3013 = w987 & w340;
assign w3014 = w997 & ~w509;
assign w3015 = w997 & w340;
assign w3016 = w1001 & w3230;
assign w3017 = w1008 & w340;
assign w3018 = w1018 & ~w509;
assign w3019 = w1018 & w340;
assign w3020 = w1024 & w3231;
assign w3021 = w1025 & w340;
assign w3022 = w1031 & w3232;
assign w3023 = w1038 & w340;
assign w3024 = w1045 & w3233;
assign w3025 = w1046 & w340;
assign w3026 = w1052 & w3234;
assign w3027 = w1059 & w340;
assign w3028 = w1062 & w3235;
assign w3029 = w1070 & w340;
assign w3030 = w1074 & w509;
assign w3031 = (w1074 & w302) | (w1074 & w3271) | (w302 & w3271);
assign w3032 = w1083 & w509;
assign w3033 = (w1083 & w302) | (w1083 & w3272) | (w302 & w3272);
assign w3034 = w1090 & w509;
assign w3035 = (w1090 & w302) | (w1090 & w3273) | (w302 & w3273);
assign w3036 = w1098 & w509;
assign w3037 = (w1098 & w302) | (w1098 & w3274) | (w302 & w3274);
assign w3038 = w1105 & w509;
assign w3039 = (w1105 & w302) | (w1105 & w3275) | (w302 & w3275);
assign w3040 = w1112 & w509;
assign w3041 = (w1112 & w302) | (w1112 & w3276) | (w302 & w3276);
assign w3042 = w1119 & w509;
assign w3043 = (w1119 & w302) | (w1119 & w3277) | (w302 & w3277);
assign w3044 = ~w1128 & w3236;
assign w3045 = w1129 & ~w340;
assign w3046 = w1135 & w509;
assign w3047 = (w1135 & w302) | (w1135 & w3278) | (w302 & w3278);
assign w3048 = w1143 & w509;
assign w3049 = (w1143 & w302) | (w1143 & w3279) | (w302 & w3279);
assign w3050 = w1151 & w509;
assign w3051 = (w1151 & w302) | (w1151 & w3280) | (w302 & w3280);
assign w3052 = w1158 & w509;
assign w3053 = (w1158 & w302) | (w1158 & w3281) | (w302 & w3281);
assign w3054 = w1166 & w509;
assign w3055 = (w1166 & w302) | (w1166 & w3282) | (w302 & w3282);
assign w3056 = w1173 & w509;
assign w3057 = (w1173 & w302) | (w1173 & w3283) | (w302 & w3283);
assign w3058 = w1180 & w509;
assign w3059 = (w1180 & w302) | (w1180 & w3284) | (w302 & w3284);
assign w3060 = w1187 & w509;
assign w3061 = (w1187 & w302) | (w1187 & w3285) | (w302 & w3285);
assign w3062 = w1194 & w509;
assign w3063 = (w1194 & w302) | (w1194 & w3286) | (w302 & w3286);
assign w3064 = w1201 & w509;
assign w3065 = (w1201 & w302) | (w1201 & w3287) | (w302 & w3287);
assign w3066 = w1208 & w509;
assign w3067 = (w1208 & w302) | (w1208 & w3288) | (w302 & w3288);
assign w3068 = w1216 & w509;
assign w3069 = (w1216 & w302) | (w1216 & w3289) | (w302 & w3289);
assign w3070 = w1224 & w509;
assign w3071 = (w1224 & w302) | (w1224 & w3290) | (w302 & w3290);
assign w3072 = w1231 & w509;
assign w3073 = (w1231 & w302) | (w1231 & w3291) | (w302 & w3291);
assign w3074 = w1247 & ~w509;
assign w3075 = w1247 & w340;
assign w3076 = w1258 & ~w509;
assign w3077 = w1258 & w340;
assign w3078 = w1269 & ~w509;
assign w3079 = w1269 & w340;
assign w3080 = w1280 & ~w509;
assign w3081 = w1280 & w340;
assign w3082 = w1284 & w509;
assign w3083 = (w1284 & w302) | (w1284 & w3292) | (w302 & w3292);
assign w3084 = w1292 & w509;
assign w3085 = (w1292 & w302) | (w1292 & w3293) | (w302 & w3293);
assign w3086 = w1299 & w509;
assign w3087 = (w1299 & w302) | (w1299 & w3294) | (w302 & w3294);
assign w3088 = w1306 & w509;
assign w3089 = (w1306 & w302) | (w1306 & w3295) | (w302 & w3295);
assign w3090 = w1320 & ~w509;
assign w3091 = w1320 & w340;
assign w3092 = w1330 & ~w509;
assign w3093 = w1330 & w340;
assign w3094 = w1340 & ~w509;
assign w3095 = w1340 & w340;
assign w3096 = w1351 & ~w509;
assign w3097 = w1351 & w340;
assign w3098 = w1362 & ~w509;
assign w3099 = w1362 & w340;
assign w3100 = w1378 & ~w509;
assign w3101 = ~w302 & w3296;
assign w3102 = w1385 & ~w509;
assign w3103 = ~w302 & w3297;
assign w3104 = w1404 & ~w509;
assign w3105 = ~w302 & w3298;
assign w3106 = w1411 & ~w509;
assign w3107 = ~w302 & w3299;
assign w3108 = w1425 & ~w509;
assign w3109 = ~w302 & w3300;
assign w3110 = w1439 & ~w509;
assign w3111 = ~w302 & w3301;
assign w3112 = w1450 & ~w509;
assign w3113 = ~w302 & w3302;
assign w3114 = w1461 & ~w509;
assign w3115 = ~w302 & w3303;
assign w3116 = w1472 & ~w509;
assign w3117 = ~w302 & w3304;
assign w3118 = w1483 & ~w509;
assign w3119 = ~w302 & w3305;
assign w3120 = w1494 & ~w509;
assign w3121 = ~w302 & w3306;
assign w3122 = w1505 & ~w509;
assign w3123 = ~w302 & w3307;
assign w3124 = w1516 & ~w509;
assign w3125 = ~w302 & w3308;
assign w3126 = w1527 & ~w509;
assign w3127 = ~w302 & w3309;
assign w3128 = w1541 & ~w509;
assign w3129 = w1541 & w340;
assign w3130 = w1544 & w509;
assign w3131 = (w1544 & w302) | (w1544 & w3310) | (w302 & w3310);
assign w3132 = w1551 & w509;
assign w3133 = (w1551 & w302) | (w1551 & w3311) | (w302 & w3311);
assign w3134 = w1558 & w509;
assign w3135 = (w1558 & w302) | (w1558 & w3312) | (w302 & w3312);
assign w3136 = w1570 & w509;
assign w3137 = (w1570 & w302) | (w1570 & w3313) | (w302 & w3313);
assign w3138 = w1578 & ~w509;
assign w3139 = ~w302 & w3314;
assign w3140 = w1589 & ~w509;
assign w3141 = ~w302 & w3315;
assign w3142 = w1600 & ~w509;
assign w3143 = ~w302 & w3316;
assign w3144 = w1614 & ~w509;
assign w3145 = w1614 & w340;
assign w3146 = w1624 & ~w509;
assign w3147 = w1624 & w340;
assign w3148 = w1631 & ~w509;
assign w3149 = ~w302 & w3317;
assign w3150 = w1638 & w509;
assign w3151 = (w1638 & w302) | (w1638 & w3318) | (w302 & w3318);
assign w3152 = w1645 & w509;
assign w3153 = (w1645 & w302) | (w1645 & w3319) | (w302 & w3319);
assign w3154 = w1652 & w509;
assign w3155 = (w1652 & w302) | (w1652 & w3320) | (w302 & w3320);
assign w3156 = w1659 & w509;
assign w3157 = (w1659 & w302) | (w1659 & w3321) | (w302 & w3321);
assign w3158 = w1666 & w509;
assign w3159 = (w1666 & w302) | (w1666 & w3322) | (w302 & w3322);
assign w3160 = w1673 & w509;
assign w3161 = (w1673 & w302) | (w1673 & w3323) | (w302 & w3323);
assign w3162 = w1680 & w509;
assign w3163 = (w1680 & w302) | (w1680 & w3324) | (w302 & w3324);
assign w3164 = w1692 & ~w509;
assign w3165 = ~w302 & w3325;
assign w3166 = w1703 & ~w509;
assign w3167 = ~w302 & w3326;
assign w3168 = w1714 & ~w509;
assign w3169 = ~w302 & w3327;
assign w3170 = w1725 & ~w509;
assign w3171 = ~w302 & w3328;
assign w3172 = w1736 & ~w509;
assign w3173 = ~w302 & w3329;
assign w3174 = w1743 & w509;
assign w3175 = (w1743 & w302) | (w1743 & w3330) | (w302 & w3330);
assign w3176 = w1750 & w509;
assign w3177 = (w1750 & w302) | (w1750 & w3331) | (w302 & w3331);
assign w3178 = w1757 & w509;
assign w3179 = (w1757 & w302) | (w1757 & w3332) | (w302 & w3332);
assign w3180 = w1768 & ~w509;
assign w3181 = ~w302 & w3333;
assign w3182 = w1775 & w509;
assign w3183 = (w1775 & w302) | (w1775 & w3334) | (w302 & w3334);
assign w3184 = w1782 & w509;
assign w3185 = (w1782 & w302) | (w1782 & w3335) | (w302 & w3335);
assign w3186 = w1793 & ~w509;
assign w3187 = ~w302 & w3336;
assign w3188 = ~w43 & ~w16;
assign w3189 = ~w43 & pi143;
assign w3190 = w1848 & ~pi035;
assign w3191 = w1848 & ~pi006;
assign w3192 = w1848 & ~pi004;
assign w3193 = w1848 & ~pi033;
assign w3194 = ~w1835 & pi017;
assign w3195 = ~w1835 & pi016;
assign w3196 = w1848 & ~pi011;
assign w3197 = w1848 & ~pi042;
assign w3198 = ~w1835 & pi125;
assign w3199 = ~w1835 & pi085;
assign w3200 = w1848 & ~pi105;
assign w3201 = ~w1848 & ~pi126;
assign w3202 = w1848 & ~pi122;
assign w3203 = w1848 & ~pi116;
assign w3204 = ~w1835 & pi094;
assign w3205 = ~w1835 & pi092;
assign w3206 = w1848 & ~pi127;
assign w3207 = w1848 & ~pi108;
assign w3208 = w1848 & ~pi106;
assign w3209 = w1848 & ~pi074;
assign w3210 = w1848 & ~pi110;
assign w3211 = w1848 & ~pi099;
assign w3212 = w582 & ~w509;
assign w3213 = w594 & ~w509;
assign w3214 = w619 & ~w509;
assign w3215 = w631 & ~w509;
assign w3216 = w643 & ~w509;
assign w3217 = w672 & ~w509;
assign w3218 = w693 & ~w509;
assign w3219 = w705 & ~w509;
assign w3220 = w719 & ~w509;
assign w3221 = w726 & ~w509;
assign w3222 = w758 & w509;
assign w3223 = w769 & w509;
assign w3224 = w884 & ~w509;
assign w3225 = w895 & ~w509;
assign w3226 = w940 & ~w509;
assign w3227 = w953 & ~w509;
assign w3228 = w964 & ~w509;
assign w3229 = w975 & ~w509;
assign w3230 = w1006 & ~w509;
assign w3231 = w1023 & ~w509;
assign w3232 = w1036 & ~w509;
assign w3233 = w1044 & ~w509;
assign w3234 = w1057 & ~w509;
assign w3235 = w1068 & ~w509;
assign w3236 = ~w529 & w509;
assign w3237 = ~pi138 & ~pi148;
assign w3238 = w2867 & pi140;
assign w3239 = ~w2867 & ~pi140;
assign w3240 = w93 & pi143;
assign w3241 = ~pi139 & ~pi140;
assign w3242 = ~w99 & ~w106;
assign w3243 = ~w136 & ~w149;
assign w3244 = ~w135 & pi082;
assign w3245 = ~w135 & pi002;
assign w3246 = ~w135 & pi100;
assign w3247 = ~w135 & pi075;
assign w3248 = ~w135 & pi078;
assign w3249 = ~w135 & pi076;
assign w3250 = ~w135 & pi028;
assign w3251 = ~w135 & pi057;
assign w3252 = ~w135 & pi063;
assign w3253 = ~w135 & pi064;
assign w3254 = ~w135 & pi024;
assign w3255 = ~w135 & pi062;
assign w3256 = ~w135 & pi021;
assign w3257 = ~w135 & pi058;
assign w3258 = ~w108 & ~w162;
assign w3259 = ~w108 & w86;
assign w3260 = ~w108 & w389;
assign w3261 = w108 & w350;
assign w3262 = ~w339 & w747;
assign w3263 = ~w339 & w774;
assign w3264 = ~w339 & w796;
assign w3265 = ~w339 & w800;
assign w3266 = ~w339 & w817;
assign w3267 = ~w339 & w835;
assign w3268 = ~w339 & w844;
assign w3269 = ~w339 & w859;
assign w3270 = ~w339 & w863;
assign w3271 = ~w339 & w1074;
assign w3272 = ~w339 & w1083;
assign w3273 = ~w339 & w1090;
assign w3274 = ~w339 & w1098;
assign w3275 = ~w339 & w1105;
assign w3276 = ~w339 & w1112;
assign w3277 = ~w339 & w1119;
assign w3278 = ~w339 & w1135;
assign w3279 = ~w339 & w1143;
assign w3280 = ~w339 & w1151;
assign w3281 = ~w339 & w1158;
assign w3282 = ~w339 & w1166;
assign w3283 = ~w339 & w1173;
assign w3284 = ~w339 & w1180;
assign w3285 = ~w339 & w1187;
assign w3286 = ~w339 & w1194;
assign w3287 = ~w339 & w1201;
assign w3288 = ~w339 & w1208;
assign w3289 = ~w339 & w1216;
assign w3290 = ~w339 & w1224;
assign w3291 = ~w339 & w1231;
assign w3292 = ~w339 & w1284;
assign w3293 = ~w339 & w1292;
assign w3294 = ~w339 & w1299;
assign w3295 = ~w339 & w1306;
assign w3296 = w339 & w1378;
assign w3297 = w339 & w1385;
assign w3298 = w339 & w1404;
assign w3299 = w339 & w1411;
assign w3300 = w339 & w1425;
assign w3301 = w339 & w1439;
assign w3302 = w339 & w1450;
assign w3303 = w339 & w1461;
assign w3304 = w339 & w1472;
assign w3305 = w339 & w1483;
assign w3306 = w339 & w1494;
assign w3307 = w339 & w1505;
assign w3308 = w339 & w1516;
assign w3309 = w339 & w1527;
assign w3310 = ~w339 & w1544;
assign w3311 = ~w339 & w1551;
assign w3312 = ~w339 & w1558;
assign w3313 = ~w339 & w1570;
assign w3314 = w339 & w1578;
assign w3315 = w339 & w1589;
assign w3316 = w339 & w1600;
assign w3317 = w339 & w1631;
assign w3318 = ~w339 & w1638;
assign w3319 = ~w339 & w1645;
assign w3320 = ~w339 & w1652;
assign w3321 = ~w339 & w1659;
assign w3322 = ~w339 & w1666;
assign w3323 = ~w339 & w1673;
assign w3324 = ~w339 & w1680;
assign w3325 = w339 & w1692;
assign w3326 = w339 & w1703;
assign w3327 = w339 & w1714;
assign w3328 = w339 & w1725;
assign w3329 = w339 & w1736;
assign w3330 = ~w339 & w1743;
assign w3331 = ~w339 & w1750;
assign w3332 = ~w339 & w1757;
assign w3333 = w339 & w1768;
assign w3334 = ~w339 & w1775;
assign w3335 = ~w339 & w1782;
assign w3336 = w339 & w1793;
assign one = 1;
assign po000 = pi202;// level 0
assign po001 = pi203;// level 0
assign po002 = pi205;// level 0
assign po003 = pi189;// level 0
assign po004 = pi200;// level 0
assign po005 = pi201;// level 0
assign po006 = pi204;// level 0
assign po007 = pi188;// level 0
assign po008 = pi210;// level 0
assign po009 = pi135;// level 0
assign po010 = pi206;// level 0
assign po011 = pi137;// level 0
assign po012 = pi209;// level 0
assign po013 = pi207;// level 0
assign po014 = pi208;// level 0
assign po015 = pi211;// level 0
assign po016 = pi213;// level 0
assign po017 = pi215;// level 0
assign po018 = pi214;// level 0
assign po019 = pi216;// level 0
assign po020 = pi225;// level 0
assign po021 = pi219;// level 0
assign po022 = pi217;// level 0
assign po023 = pi223;// level 0
assign po024 = pi222;// level 0
assign po025 = pi227;// level 0
assign po026 = pi212;// level 0
assign po027 = pi218;// level 0
assign po028 = pi221;// level 0
assign po029 = pi226;// level 0
assign po030 = pi224;// level 0
assign po031 = pi220;// level 0
assign po032 = pi228;// level 0
assign po033 = pi134;// level 0
assign po034 = pi129;// level 0
assign po035 = pi128;// level 0
assign po036 = ~w1;// level 2
assign po037 = ~w2;// level 2
assign po038 = ~w3;// level 2
assign po039 = ~w4;// level 2
assign po040 = ~w5;// level 2
assign po041 = ~w6;// level 2
assign po042 = ~w7;// level 2
assign po043 = ~w8;// level 2
assign po044 = ~pi230;// level 0
assign po045 = one;// level 0
assign po046 = pi229;// level 0
assign po047 = w512;// level 19
assign po048 = w528;// level 19
assign po049 = w544;// level 19
assign po050 = w555;// level 19
assign po051 = w572;// level 19
assign po052 = w586;// level 19
assign po053 = w598;// level 19
assign po054 = w608;// level 19
assign po055 = w623;// level 19
assign po056 = w635;// level 19
assign po057 = w647;// level 19
assign po058 = w663;// level 19
assign po059 = w676;// level 19
assign po060 = w687;// level 19
assign po061 = w701;// level 19
assign po062 = w712;// level 19
assign po063 = w723;// level 19
assign po064 = w733;// level 19
assign po065 = ~w749;// level 19
assign po066 = ~w761;// level 19
assign po067 = ~w772;// level 19
assign po068 = ~w783;// level 19
assign po069 = ~w798;// level 19
assign po070 = ~w807;// level 19
assign po071 = ~w819;// level 19
assign po072 = ~w833;// level 19
assign po073 = ~w842;// level 19
assign po074 = ~w850;// level 19
assign po075 = ~w861;// level 19
assign po076 = ~w869;// level 19
assign po077 = ~w880;// level 19
assign po078 = w891;// level 19
assign po079 = w902;// level 19
assign po080 = w912;// level 19
assign po081 = w924;// level 19
assign po082 = w935;// level 19
assign po083 = w947;// level 19
assign po084 = w957;// level 19
assign po085 = w968;// level 19
assign po086 = w979;// level 19
assign po087 = w989;// level 19
assign po088 = w999;// level 19
assign po089 = w1010;// level 19
assign po090 = w1020;// level 19
assign po091 = w1030;// level 19
assign po092 = w1040;// level 19
assign po093 = w1051;// level 19
assign po094 = w1061;// level 19
assign po095 = w1072;// level 19
assign po096 = ~w1081;// level 19
assign po097 = ~w1089;// level 19
assign po098 = ~w1096;// level 19
assign po099 = ~w1104;// level 19
assign po100 = ~w1111;// level 19
assign po101 = ~w1118;// level 19
assign po102 = ~w1125;// level 19
assign po103 = ~w1134;// level 19
assign po104 = ~w1142;// level 19
assign po105 = ~w1150;// level 19
assign po106 = ~w1157;// level 19
assign po107 = ~w1165;// level 19
assign po108 = ~w1172;// level 19
assign po109 = ~w1179;// level 19
assign po110 = ~w1186;// level 19
assign po111 = ~w1193;// level 19
assign po112 = ~w1200;// level 19
assign po113 = ~w1207;// level 19
assign po114 = ~w1214;// level 19
assign po115 = ~w1223;// level 19
assign po116 = ~w1230;// level 19
assign po117 = ~w1237;// level 19
assign po118 = w1249;// level 19
assign po119 = w1260;// level 19
assign po120 = w1271;// level 19
assign po121 = w1282;// level 19
assign po122 = ~w1291;// level 19
assign po123 = ~w1298;// level 19
assign po124 = ~w1305;// level 19
assign po125 = ~w1312;// level 19
assign po126 = w1322;// level 19
assign po127 = w1332;// level 19
assign po128 = w1342;// level 19
assign po129 = w1353;// level 19
assign po130 = w1364;// level 19
assign po131 = w1380;// level 19
assign po132 = w1391;// level 19
assign po133 = w1406;// level 19
assign po134 = w1417;// level 19
assign po135 = w1431;// level 19
assign po136 = w1445;// level 19
assign po137 = w1456;// level 19
assign po138 = w1467;// level 19
assign po139 = w1478;// level 19
assign po140 = w1489;// level 19
assign po141 = w1500;// level 19
assign po142 = w1511;// level 19
assign po143 = w1522;// level 19
assign po144 = w1533;// level 19
assign po145 = w1543;// level 19
assign po146 = ~w1550;// level 19
assign po147 = ~w1557;// level 19
assign po148 = ~w1564;// level 19
assign po149 = ~w1573;// level 19
assign po150 = w1584;// level 19
assign po151 = w1595;// level 19
assign po152 = w1606;// level 19
assign po153 = w1616;// level 19
assign po154 = w1626;// level 19
assign po155 = w1637;// level 19
assign po156 = ~w1644;// level 19
assign po157 = ~w1651;// level 19
assign po158 = ~w1658;// level 19
assign po159 = ~w1665;// level 19
assign po160 = ~w1672;// level 19
assign po161 = ~w1679;// level 19
assign po162 = ~w1687;// level 19
assign po163 = w1698;// level 19
assign po164 = w1709;// level 19
assign po165 = w1720;// level 19
assign po166 = w1731;// level 19
assign po167 = w1742;// level 19
assign po168 = ~w1749;// level 19
assign po169 = ~w1756;// level 19
assign po170 = ~w1763;// level 19
assign po171 = w1774;// level 19
assign po172 = ~w1781;// level 19
assign po173 = ~w1788;// level 19
assign po174 = w1799;// level 19
assign po175 = w2232;// level 18
assign po176 = ~w2253;// level 15
assign po177 = w2271;// level 11
assign po178 = w2281;// level 12
assign po179 = ~w2286;// level 15
assign po180 = w2291;// level 10
assign po181 = ~w2294;// level 11
assign po182 = ~w2308;// level 6
assign po183 = ~w2310;// level 10
assign po184 = ~w2321;// level 6
assign po185 = ~w2325;// level 6
assign po186 = ~w2330;// level 8
assign po187 = w2335;// level 9
assign po188 = ~w2340;// level 15
assign po189 = w2345;// level 7
assign po190 = ~w2348;// level 6
assign po191 = ~w2351;// level 6
assign po192 = ~w2380;// level 7
assign po193 = ~w2384;// level 7
assign po194 = w2388;// level 15
assign po195 = w2393;// level 6
assign po196 = ~w2398;// level 15
assign po197 = ~w2400;// level 5
assign po198 = ~w2403;// level 6
assign po199 = ~w2406;// level 6
assign po200 = ~w2411;// level 6
assign po201 = w2416;// level 15
assign po202 = ~w2420;// level 6
assign po203 = ~w2424;// level 6
assign po204 = ~w2427;// level 6
assign po205 = ~w2430;// level 6
assign po206 = ~w2435;// level 15
assign po207 = ~w2438;// level 6
assign po208 = ~w2441;// level 6
assign po209 = ~w2448;// level 15
assign po210 = ~w2451;// level 6
assign po211 = ~w2458;// level 15
assign po212 = w2461;// level 15
assign po213 = ~w2466;// level 15
assign po214 = w2472;// level 15
assign po215 = ~w2477;// level 15
assign po216 = w2482;// level 15
assign po217 = w2487;// level 15
assign po218 = ~w2490;// level 6
assign po219 = ~w2493;// level 6
assign po220 = ~w2496;// level 6
assign po221 = ~w2499;// level 6
assign po222 = ~w2502;// level 6
assign po223 = ~w2505;// level 6
assign po224 = ~w2508;// level 6
assign po225 = ~w2511;// level 6
assign po226 = ~w2514;// level 6
assign po227 = ~w2517;// level 6
assign po228 = ~w2520;// level 6
assign po229 = ~w2523;// level 6
assign po230 = ~w2526;// level 6
assign po231 = ~w2529;// level 6
assign po232 = ~w2532;// level 6
assign po233 = ~w2537;// level 15
assign po234 = ~w2543;// level 5
assign po235 = ~w2557;// level 6
assign po236 = ~w2570;// level 6
assign po237 = ~w2575;// level 4
assign po238 = ~w2580;// level 15
assign po239 = ~w2585;// level 6
assign po240 = ~w2588;// level 6
assign po241 = ~w2591;// level 6
assign po242 = ~w2594;// level 6
assign po243 = ~w2597;// level 6
assign po244 = ~w2600;// level 6
assign po245 = ~w2603;// level 6
assign po246 = ~w2606;// level 6
assign po247 = ~w2619;// level 6
assign po248 = ~w2632;// level 6
assign po249 = ~w2645;// level 6
assign po250 = ~w2658;// level 6
assign po251 = ~w2671;// level 6
assign po252 = ~w2684;// level 6
assign po253 = ~w2695;// level 6
assign po254 = ~w2706;// level 6
assign po255 = ~w2715;// level 6
assign po256 = ~w2726;// level 6
assign po257 = ~w2737;// level 6
assign po258 = ~w2746;// level 6
assign po259 = ~w2753;// level 5
assign po260 = ~w2760;// level 5
assign po261 = ~w2767;// level 5
assign po262 = ~w2774;// level 5
assign po263 = ~w2781;// level 5
assign po264 = ~w2788;// level 5
assign po265 = ~w2795;// level 5
assign po266 = ~w2802;// level 5
assign po267 = ~w2809;// level 5
assign po268 = ~w2816;// level 5
assign po269 = ~w2823;// level 5
assign po270 = ~w2830;// level 5
assign po271 = ~w2837;// level 5
assign po272 = ~w2844;// level 5
assign po273 = ~w2851;// level 5
assign po274 = ~w2858;// level 5
assign po275 = w2859;// level 2
endmodule
