// Benchmark "sasc" written by ABC on Wed Apr 29 13:50:37 2015

module sasc ( 
    pi000, pi001, pi002, pi003, pi004, pi005, pi006, pi007, pi008, pi009,
    pi010, pi011, pi012, pi013, pi014, pi015, pi016, pi017, pi018, pi019,
    pi020, pi021, pi022, pi023, pi024, pi025, pi026, pi027, pi028, pi029,
    pi030, pi031, pi032, pi033, pi034, pi035, pi036, pi037, pi038, pi039,
    pi040, pi041, pi042, pi043, pi044, pi045, pi046, pi047, pi048, pi049,
    pi050, pi051, pi052, pi053, pi054, pi055, pi056, pi057, pi058, pi059,
    pi060, pi061, pi062, pi063, pi064, pi065, pi066, pi067, pi068, pi069,
    pi070, pi071, pi072, pi073, pi074, pi075, pi076, pi077, pi078, pi079,
    pi080, pi081, pi082, pi083, pi084, pi085, pi086, pi087, pi088, pi089,
    pi090, pi091, pi092, pi093, pi094, pi095, pi096, pi097, pi098, pi099,
    pi100, pi101, pi102, pi103, pi104, pi105, pi106, pi107, pi108, pi109,
    pi110, pi111, pi112, pi113, pi114, pi115, pi116, pi117, pi118, pi119,
    pi120, pi121, pi122, pi123, pi124, pi125, pi126, pi127, pi128, pi129,
    pi130, pi131, pi132,
    po000, po001, po002, po003, po004, po005, po006, po007, po008, po009,
    po010, po011, po012, po013, po014, po015, po016, po017, po018, po019,
    po020, po021, po022, po023, po024, po025, po026, po027, po028, po029,
    po030, po031, po032, po033, po034, po035, po036, po037, po038, po039,
    po040, po041, po042, po043, po044, po045, po046, po047, po048, po049,
    po050, po051, po052, po053, po054, po055, po056, po057, po058, po059,
    po060, po061, po062, po063, po064, po065, po066, po067, po068, po069,
    po070, po071, po072, po073, po074, po075, po076, po077, po078, po079,
    po080, po081, po082, po083, po084, po085, po086, po087, po088, po089,
    po090, po091, po092, po093, po094, po095, po096, po097, po098, po099,
    po100, po101, po102, po103, po104, po105, po106, po107, po108, po109,
    po110, po111, po112, po113, po114, po115, po116, po117, po118, po119,
    po120, po121, po122, po123, po124, po125, po126, po127, po128, po129,
    po130, po131  );
  input  pi000, pi001, pi002, pi003, pi004, pi005, pi006, pi007, pi008,
    pi009, pi010, pi011, pi012, pi013, pi014, pi015, pi016, pi017, pi018,
    pi019, pi020, pi021, pi022, pi023, pi024, pi025, pi026, pi027, pi028,
    pi029, pi030, pi031, pi032, pi033, pi034, pi035, pi036, pi037, pi038,
    pi039, pi040, pi041, pi042, pi043, pi044, pi045, pi046, pi047, pi048,
    pi049, pi050, pi051, pi052, pi053, pi054, pi055, pi056, pi057, pi058,
    pi059, pi060, pi061, pi062, pi063, pi064, pi065, pi066, pi067, pi068,
    pi069, pi070, pi071, pi072, pi073, pi074, pi075, pi076, pi077, pi078,
    pi079, pi080, pi081, pi082, pi083, pi084, pi085, pi086, pi087, pi088,
    pi089, pi090, pi091, pi092, pi093, pi094, pi095, pi096, pi097, pi098,
    pi099, pi100, pi101, pi102, pi103, pi104, pi105, pi106, pi107, pi108,
    pi109, pi110, pi111, pi112, pi113, pi114, pi115, pi116, pi117, pi118,
    pi119, pi120, pi121, pi122, pi123, pi124, pi125, pi126, pi127, pi128,
    pi129, pi130, pi131, pi132;
  output po000, po001, po002, po003, po004, po005, po006, po007, po008, po009,
    po010, po011, po012, po013, po014, po015, po016, po017, po018, po019,
    po020, po021, po022, po023, po024, po025, po026, po027, po028, po029,
    po030, po031, po032, po033, po034, po035, po036, po037, po038, po039,
    po040, po041, po042, po043, po044, po045, po046, po047, po048, po049,
    po050, po051, po052, po053, po054, po055, po056, po057, po058, po059,
    po060, po061, po062, po063, po064, po065, po066, po067, po068, po069,
    po070, po071, po072, po073, po074, po075, po076, po077, po078, po079,
    po080, po081, po082, po083, po084, po085, po086, po087, po088, po089,
    po090, po091, po092, po093, po094, po095, po096, po097, po098, po099,
    po100, po101, po102, po103, po104, po105, po106, po107, po108, po109,
    po110, po111, po112, po113, po114, po115, po116, po117, po118, po119,
    po120, po121, po122, po123, po124, po125, po126, po127, po128, po129,
    po130, po131;
  wire n267, n268, n269, n270, n271, n272, n273, n275, n276, n277, n278,
    n279, n280, n281, n283, n284, n285, n286, n287, n288, n289, n290, n291,
    n292, n294, n295, n296, n297, n298, n299, n301, n302, n303, n304, n305,
    n306, n308, n309, n310, n311, n312, n313, n315, n316, n317, n318, n319,
    n320, n322, n323, n324, n325, n326, n327, n329, n330, n331, n332, n333,
    n334, n336, n337, n338, n339, n340, n341, n343, n344, n345, n346, n347,
    n348, n349, n350, n351, n352, n353, n354, n355, n356, n358, n359, n360,
    n361, n362, n363, n365, n366, n368, n369, n370, n371, n372, n374, n375,
    n376, n377, n378, n380, n381, n382, n383, n384, n386, n387, n388, n389,
    n390, n392, n393, n394, n395, n396, n398, n399, n400, n401, n402, n404,
    n405, n406, n407, n408, n410, n411, n412, n413, n414, n416, n417, n418,
    n419, n420, n422, n423, n424, n425, n426, n428, n429, n430, n431, n432,
    n434, n435, n436, n437, n438, n440, n441, n442, n443, n444, n446, n447,
    n448, n449, n450, n452, n453, n454, n455, n456, n458, n459, n460, n461,
    n462, n464, n465, n466, n467, n468, n469, n471, n472, n473, n474, n475,
    n477, n478, n479, n480, n481, n483, n484, n485, n486, n487, n489, n490,
    n491, n492, n493, n495, n496, n497, n498, n499, n501, n502, n503, n504,
    n505, n507, n508, n509, n510, n511, n513, n514, n515, n516, n517, n518,
    n520, n521, n522, n523, n524, n526, n527, n528, n529, n530, n532, n533,
    n534, n535, n536, n538, n539, n540, n541, n542, n544, n545, n546, n547,
    n548, n550, n551, n552, n553, n554, n556, n557, n558, n559, n560, n562,
    n563, n564, n565, n566, n567, n568, n569, n570, n571, n573, n574, n576,
    n577, n578, n579, n580, n581, n582, n583, n584, n586, n587, n588, n589,
    n591, n592, n593, n594, n595, n596, n598, n599, n601, n602, n604, n605,
    n607, n608, n610, n611, n613, n614, n616, n617, n619, n620, n622, n623,
    n624, n625, n626, n627, n628, n629, n630, n631, n632, n634, n635, n636,
    n637, n638, n639, n640, n641, n642, n643, n645, n646, n647, n648, n649,
    n650, n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n662,
    n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, n673, n675,
    n676, n677, n678, n679, n680, n681, n682, n683, n684, n685, n686, n688,
    n689, n690, n691, n692, n693, n694, n695, n696, n697, n698, n699, n701,
    n702, n703, n704, n705, n706, n707, n708, n709, n710, n711, n712, n714,
    n715, n716, n717, n718, n719, n720, n721, n722, n723, n724, n725, n727,
    n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738, n740,
    n741, n742, n743, n744, n745, n746, n748, n749, n750, n751, n752, n753,
    n754, n755, n756, n757, n758, n759, n761, n762, n763, n764, n766, n767,
    n768, n769, n770, n772, n773, n774, n776, n777, n778, n779, n780, n781,
    n782, n784, n785, n786, n787, n789, n790, n791, n792, n793, n795, n796,
    n797, n798, n799, n801, n802, n803, n804, n805, n807, n808, n809, n810,
    n811, n813, n814, n815, n816, n817, n819, n820, n821, n822, n823, n825,
    n826, n827, n828, n829, n831, n832, n833, n834, n835, n837, n838, n839,
    n840, n841, n843, n844, n845, n846, n847, n849, n850, n851, n852, n853,
    n855, n856, n857, n858, n859, n861, n862, n863, n864, n865, n867, n868,
    n869, n870, n871, n873, n874, n875, n877, n878, n879, n881, n882, n883,
    n884, n885, n887, n888, n889, n890, n891, n893, n894, n895, n896, n897,
    n898, n900, n901, n902, n903, n904, n906, n907, n908, n909, n910, n912,
    n913, n914, n915, n916, n917, n919, n920, n921, n922, n923, n924, n926,
    n927, n928, n929, n930, n932, n933, n934, n935, n936, n938, n939, n940,
    n941, n942, n944, n945, n946, n947, n948, n950, n951, n952, n953, n954,
    n956, n957, n958, n959, n960, n962, n963, n964, n965, n966, n968, n969,
    n970, n971, n972, n974, n975, n976, n977, n978, n980, n981, n982, n984,
    n986, n987, n988, n989, n990, n992, n993, n994, n995, n996, n998, n999,
    n1000, n1001, n1002, n1004, n1005, n1006, n1007, n1008, n1009, n1012,
    n1013, n1015, n1016, n1018, n1019, n1021, n1022, n1024, n1025, n1027,
    n1028, n1030, n1031, n1033, n1035, n1036, n1038;
  assign n267 = ~pi077 & pi104;
  assign n268 = pi077 & ~pi104;
  assign n269 = ~n267 & ~n268;
  assign n270 = ~pi109 & ~pi112;
  assign n271 = pi109 & pi112;
  assign n272 = ~n270 & ~n271;
  assign n273 = n269 & ~n272;
  assign po002 = ~pi048 & n273;
  assign n275 = pi035 & ~pi096;
  assign n276 = ~pi035 & pi096;
  assign n277 = ~n275 & ~n276;
  assign n278 = pi001 & pi107;
  assign n279 = ~pi001 & ~pi107;
  assign n280 = ~n278 & ~n279;
  assign n281 = n277 & ~n280;
  assign po003 = ~pi000 & n281;
  assign n283 = pi096 & ~pi107;
  assign n284 = pi004 & n283;
  assign n285 = pi096 & pi107;
  assign n286 = pi018 & n285;
  assign n287 = ~n284 & ~n286;
  assign n288 = ~pi096 & pi107;
  assign n289 = pi012 & n288;
  assign n290 = ~pi096 & ~pi107;
  assign n291 = pi026 & n290;
  assign n292 = ~n289 & ~n291;
  assign po004 = ~n287 | ~n292;
  assign n294 = pi005 & n283;
  assign n295 = pi019 & n285;
  assign n296 = ~n294 & ~n295;
  assign n297 = pi013 & n288;
  assign n298 = pi027 & n290;
  assign n299 = ~n297 & ~n298;
  assign po005 = ~n296 | ~n299;
  assign n301 = pi006 & n283;
  assign n302 = pi020 & n285;
  assign n303 = ~n301 & ~n302;
  assign n304 = pi014 & n288;
  assign n305 = pi028 & n290;
  assign n306 = ~n304 & ~n305;
  assign po006 = ~n303 | ~n306;
  assign n308 = pi007 & n283;
  assign n309 = pi021 & n285;
  assign n310 = ~n308 & ~n309;
  assign n311 = pi015 & n288;
  assign n312 = pi029 & n290;
  assign n313 = ~n311 & ~n312;
  assign po007 = ~n310 | ~n313;
  assign n315 = pi008 & n283;
  assign n316 = pi022 & n285;
  assign n317 = ~n315 & ~n316;
  assign n318 = pi016 & n288;
  assign n319 = pi030 & n290;
  assign n320 = ~n318 & ~n319;
  assign po008 = ~n317 | ~n320;
  assign n322 = pi009 & n283;
  assign n323 = pi023 & n285;
  assign n324 = ~n322 & ~n323;
  assign n325 = pi017 & n288;
  assign n326 = pi031 & n290;
  assign n327 = ~n325 & ~n326;
  assign po009 = ~n324 | ~n327;
  assign n329 = pi002 & n288;
  assign n330 = pi032 & n290;
  assign n331 = ~n329 & ~n330;
  assign n332 = pi010 & n283;
  assign n333 = pi024 & n285;
  assign n334 = ~n332 & ~n333;
  assign po010 = ~n331 | ~n334;
  assign n336 = pi003 & n288;
  assign n337 = pi033 & n290;
  assign n338 = ~n336 & ~n337;
  assign n339 = pi011 & n283;
  assign n340 = pi025 & n285;
  assign n341 = ~n339 & ~n340;
  assign po011 = ~n338 | ~n341;
  assign n343 = pi001 & ~pi107;
  assign n344 = ~pi001 & pi107;
  assign n345 = ~n343 & ~n344;
  assign n346 = ~pi001 & pi035;
  assign n347 = pi001 & ~pi035;
  assign n348 = ~n346 & ~n347;
  assign n349 = pi096 & ~n348;
  assign n350 = ~pi096 & n348;
  assign n351 = ~n349 & ~n350;
  assign n352 = ~pi035 & ~pi096;
  assign n353 = pi000 & n352;
  assign n354 = pi035 & pi096;
  assign n355 = pi000 & n354;
  assign n356 = ~n353 & ~n355;
  assign po076 = ~n280 & ~n356;
  assign n358 = pi083 & pi106;
  assign n359 = ~po076 & n358;
  assign n360 = ~n351 & n359;
  assign n361 = ~n345 & n360;
  assign n362 = pi000 & ~pi123;
  assign n363 = ~n361 & ~n362;
  assign po014 = pi118 & ~n363;
  assign n365 = pi001 & ~n359;
  assign n366 = ~pi001 & n359;
  assign po016 = n365 | n366;
  assign n368 = pi045 & n347;
  assign n369 = pi002 & ~n347;
  assign n370 = ~n368 & ~n369;
  assign n371 = n359 & ~n370;
  assign n372 = pi002 & ~n359;
  assign po017 = n371 | n372;
  assign n374 = pi040 & n347;
  assign n375 = pi003 & ~n347;
  assign n376 = ~n374 & ~n375;
  assign n377 = n359 & ~n376;
  assign n378 = pi003 & ~n359;
  assign po018 = n377 | n378;
  assign n380 = pi041 & n346;
  assign n381 = pi004 & ~n346;
  assign n382 = ~n380 & ~n381;
  assign n383 = n359 & ~n382;
  assign n384 = pi004 & ~n359;
  assign po019 = n383 | n384;
  assign n386 = pi039 & n346;
  assign n387 = pi005 & ~n346;
  assign n388 = ~n386 & ~n387;
  assign n389 = n359 & ~n388;
  assign n390 = pi005 & ~n359;
  assign po020 = n389 | n390;
  assign n392 = pi042 & n346;
  assign n393 = pi006 & ~n346;
  assign n394 = ~n392 & ~n393;
  assign n395 = n359 & ~n394;
  assign n396 = pi006 & ~n359;
  assign po021 = n395 | n396;
  assign n398 = pi043 & n346;
  assign n399 = pi007 & ~n346;
  assign n400 = ~n398 & ~n399;
  assign n401 = n359 & ~n400;
  assign n402 = pi007 & ~n359;
  assign po022 = n401 | n402;
  assign n404 = pi044 & n346;
  assign n405 = pi008 & ~n346;
  assign n406 = ~n404 & ~n405;
  assign n407 = n359 & ~n406;
  assign n408 = pi008 & ~n359;
  assign po023 = n407 | n408;
  assign n410 = pi046 & n346;
  assign n411 = pi009 & ~n346;
  assign n412 = ~n410 & ~n411;
  assign n413 = n359 & ~n412;
  assign n414 = pi009 & ~n359;
  assign po024 = n413 | n414;
  assign n416 = pi045 & n346;
  assign n417 = pi010 & ~n346;
  assign n418 = ~n416 & ~n417;
  assign n419 = n359 & ~n418;
  assign n420 = pi010 & ~n359;
  assign po025 = n419 | n420;
  assign n422 = pi040 & n346;
  assign n423 = pi011 & ~n346;
  assign n424 = ~n422 & ~n423;
  assign n425 = n359 & ~n424;
  assign n426 = pi011 & ~n359;
  assign po026 = n425 | n426;
  assign n428 = pi041 & n347;
  assign n429 = pi012 & ~n347;
  assign n430 = ~n428 & ~n429;
  assign n431 = n359 & ~n430;
  assign n432 = pi012 & ~n359;
  assign po027 = n431 | n432;
  assign n434 = pi039 & n347;
  assign n435 = pi013 & ~n347;
  assign n436 = ~n434 & ~n435;
  assign n437 = n359 & ~n436;
  assign n438 = pi013 & ~n359;
  assign po028 = n437 | n438;
  assign n440 = pi042 & n347;
  assign n441 = pi014 & ~n347;
  assign n442 = ~n440 & ~n441;
  assign n443 = n359 & ~n442;
  assign n444 = pi014 & ~n359;
  assign po029 = n443 | n444;
  assign n446 = pi043 & n347;
  assign n447 = pi015 & ~n347;
  assign n448 = ~n446 & ~n447;
  assign n449 = n359 & ~n448;
  assign n450 = pi015 & ~n359;
  assign po030 = n449 | n450;
  assign n452 = pi044 & n347;
  assign n453 = pi016 & ~n347;
  assign n454 = ~n452 & ~n453;
  assign n455 = n359 & ~n454;
  assign n456 = pi016 & ~n359;
  assign po031 = n455 | n456;
  assign n458 = pi046 & n347;
  assign n459 = pi017 & ~n347;
  assign n460 = ~n458 & ~n459;
  assign n461 = n359 & ~n460;
  assign n462 = pi017 & ~n359;
  assign po032 = n461 | n462;
  assign n464 = pi001 & pi035;
  assign n465 = pi041 & n464;
  assign n466 = pi018 & ~n464;
  assign n467 = ~n465 & ~n466;
  assign n468 = n359 & ~n467;
  assign n469 = pi018 & ~n359;
  assign po033 = n468 | n469;
  assign n471 = pi039 & n464;
  assign n472 = pi019 & ~n464;
  assign n473 = ~n471 & ~n472;
  assign n474 = n359 & ~n473;
  assign n475 = pi019 & ~n359;
  assign po034 = n474 | n475;
  assign n477 = pi042 & n464;
  assign n478 = pi020 & ~n464;
  assign n479 = ~n477 & ~n478;
  assign n480 = n359 & ~n479;
  assign n481 = pi020 & ~n359;
  assign po035 = n480 | n481;
  assign n483 = pi043 & n464;
  assign n484 = pi021 & ~n464;
  assign n485 = ~n483 & ~n484;
  assign n486 = n359 & ~n485;
  assign n487 = pi021 & ~n359;
  assign po036 = n486 | n487;
  assign n489 = pi044 & n464;
  assign n490 = pi022 & ~n464;
  assign n491 = ~n489 & ~n490;
  assign n492 = n359 & ~n491;
  assign n493 = pi022 & ~n359;
  assign po037 = n492 | n493;
  assign n495 = pi046 & n464;
  assign n496 = pi023 & ~n464;
  assign n497 = ~n495 & ~n496;
  assign n498 = n359 & ~n497;
  assign n499 = pi023 & ~n359;
  assign po038 = n498 | n499;
  assign n501 = pi045 & n464;
  assign n502 = pi024 & ~n464;
  assign n503 = ~n501 & ~n502;
  assign n504 = n359 & ~n503;
  assign n505 = pi024 & ~n359;
  assign po039 = n504 | n505;
  assign n507 = pi040 & n464;
  assign n508 = pi025 & ~n464;
  assign n509 = ~n507 & ~n508;
  assign n510 = n359 & ~n509;
  assign n511 = pi025 & ~n359;
  assign po040 = n510 | n511;
  assign n513 = ~pi001 & ~pi035;
  assign n514 = pi026 & ~n513;
  assign n515 = pi041 & n513;
  assign n516 = ~n514 & ~n515;
  assign n517 = n359 & ~n516;
  assign n518 = pi026 & ~n359;
  assign po041 = n517 | n518;
  assign n520 = pi027 & ~n513;
  assign n521 = pi039 & n513;
  assign n522 = ~n520 & ~n521;
  assign n523 = n359 & ~n522;
  assign n524 = pi027 & ~n359;
  assign po042 = n523 | n524;
  assign n526 = pi028 & ~n513;
  assign n527 = pi042 & n513;
  assign n528 = ~n526 & ~n527;
  assign n529 = n359 & ~n528;
  assign n530 = pi028 & ~n359;
  assign po043 = n529 | n530;
  assign n532 = pi029 & ~n513;
  assign n533 = pi043 & n513;
  assign n534 = ~n532 & ~n533;
  assign n535 = n359 & ~n534;
  assign n536 = pi029 & ~n359;
  assign po044 = n535 | n536;
  assign n538 = pi030 & ~n513;
  assign n539 = pi044 & n513;
  assign n540 = ~n538 & ~n539;
  assign n541 = n359 & ~n540;
  assign n542 = pi030 & ~n359;
  assign po045 = n541 | n542;
  assign n544 = pi031 & ~n513;
  assign n545 = pi046 & n513;
  assign n546 = ~n544 & ~n545;
  assign n547 = n359 & ~n546;
  assign n548 = pi031 & ~n359;
  assign po046 = n547 | n548;
  assign n550 = pi032 & ~n513;
  assign n551 = pi045 & n513;
  assign n552 = ~n550 & ~n551;
  assign n553 = n359 & ~n552;
  assign n554 = pi032 & ~n359;
  assign po047 = n553 | n554;
  assign n556 = pi033 & ~n513;
  assign n557 = pi040 & n513;
  assign n558 = ~n556 & ~n557;
  assign n559 = n359 & ~n558;
  assign n560 = pi033 & ~n359;
  assign po048 = n559 | n560;
  assign n562 = ~pi108 & ~pi116;
  assign n563 = ~pi115 & n562;
  assign n564 = ~pi034 & pi037;
  assign n565 = pi034 & ~pi037;
  assign n566 = ~n564 & ~n565;
  assign n567 = pi102 & pi108;
  assign n568 = ~n566 & n567;
  assign n569 = pi034 & ~n567;
  assign n570 = ~n568 & ~n569;
  assign n571 = ~n563 & ~n570;
  assign po049 = ~pi118 | n571;
  assign n573 = ~n348 & n359;
  assign n574 = pi035 & ~n359;
  assign po050 = n573 | n574;
  assign n576 = pi034 & pi037;
  assign n577 = pi038 & n576;
  assign n578 = pi036 & n577;
  assign n579 = ~pi036 & ~n577;
  assign n580 = ~n578 & ~n579;
  assign n581 = n567 & n580;
  assign n582 = pi036 & ~n567;
  assign n583 = ~n581 & ~n582;
  assign n584 = ~n563 & ~n583;
  assign po051 = ~pi118 | n584;
  assign n586 = ~pi037 & n567;
  assign n587 = pi037 & ~n567;
  assign n588 = ~n586 & ~n587;
  assign n589 = pi118 & ~n563;
  assign po052 = ~n588 & n589;
  assign n591 = ~pi038 & n576;
  assign n592 = pi038 & ~n576;
  assign n593 = ~n591 & ~n592;
  assign n594 = n567 & ~n593;
  assign n595 = pi038 & ~n567;
  assign n596 = ~n594 & ~n595;
  assign po053 = n589 & ~n596;
  assign n598 = pi042 & n567;
  assign n599 = pi039 & ~n567;
  assign po054 = n598 | n599;
  assign n601 = pi116 & n567;
  assign n602 = pi040 & ~n567;
  assign po055 = n601 | n602;
  assign n604 = pi039 & n567;
  assign n605 = pi041 & ~n567;
  assign po056 = n604 | n605;
  assign n607 = pi043 & n567;
  assign n608 = pi042 & ~n567;
  assign po057 = n607 | n608;
  assign n610 = pi044 & n567;
  assign n611 = pi043 & ~n567;
  assign po058 = n610 | n611;
  assign n613 = pi046 & n567;
  assign n614 = pi044 & ~n567;
  assign po059 = n613 | n614;
  assign n616 = pi040 & n567;
  assign n617 = pi045 & ~n567;
  assign po060 = n616 | n617;
  assign n619 = pi045 & n567;
  assign n620 = pi046 & ~n567;
  assign po061 = n619 | n620;
  assign n622 = pi113 & pi121;
  assign n623 = pi062 & pi101;
  assign n624 = pi056 & n623;
  assign n625 = pi047 & n624;
  assign n626 = ~pi047 & ~n624;
  assign n627 = ~n625 & ~n626;
  assign n628 = n622 & n627;
  assign n629 = pi047 & ~n622;
  assign n630 = ~n628 & ~n629;
  assign n631 = pi110 & pi121;
  assign n632 = ~n630 & ~n631;
  assign po062 = ~pi118 | n632;
  assign n634 = ~pi048 & ~n631;
  assign n635 = ~pi104 & pi112;
  assign n636 = pi104 & ~pi112;
  assign n637 = ~n635 & ~n636;
  assign n638 = ~pi077 & n637;
  assign n639 = pi077 & ~n637;
  assign n640 = ~n638 & ~n639;
  assign n641 = n272 & ~n640;
  assign n642 = pi124 & n641;
  assign n643 = ~n634 & ~n642;
  assign po063 = pi118 & ~n643;
  assign n645 = ~pi050 & n622;
  assign n646 = ~pi049 & ~n622;
  assign n647 = ~n645 & ~n646;
  assign n648 = ~n631 & ~n647;
  assign n649 = ~pi077 & pi109;
  assign n650 = pi079 & n649;
  assign n651 = pi077 & ~pi109;
  assign n652 = pi080 & n651;
  assign n653 = ~n650 & ~n652;
  assign n654 = ~pi077 & ~pi109;
  assign n655 = pi099 & n654;
  assign n656 = pi077 & pi109;
  assign n657 = pi084 & n656;
  assign n658 = ~n655 & ~n657;
  assign n659 = n653 & n658;
  assign n660 = n631 & ~n659;
  assign po064 = n648 | n660;
  assign n662 = ~pi051 & n622;
  assign n663 = ~pi050 & ~n622;
  assign n664 = ~n662 & ~n663;
  assign n665 = ~n631 & ~n664;
  assign n666 = pi082 & n656;
  assign n667 = pi068 & n649;
  assign n668 = ~n666 & ~n667;
  assign n669 = pi098 & n654;
  assign n670 = pi074 & n651;
  assign n671 = ~n669 & ~n670;
  assign n672 = n668 & n671;
  assign n673 = n631 & ~n672;
  assign po065 = n665 | n673;
  assign n675 = pi097 & n622;
  assign n676 = ~pi051 & ~n622;
  assign n677 = ~n675 & ~n676;
  assign n678 = ~n631 & ~n677;
  assign n679 = pi089 & n654;
  assign n680 = pi069 & n649;
  assign n681 = ~n679 & ~n680;
  assign n682 = pi095 & n656;
  assign n683 = pi075 & n651;
  assign n684 = ~n682 & ~n683;
  assign n685 = n681 & n684;
  assign n686 = n631 & ~n685;
  assign po066 = n678 | n686;
  assign n688 = ~pi053 & n622;
  assign n689 = ~pi052 & ~n622;
  assign n690 = ~n688 & ~n689;
  assign n691 = ~n631 & ~n690;
  assign n692 = pi091 & n656;
  assign n693 = pi070 & n651;
  assign n694 = ~n692 & ~n693;
  assign n695 = pi086 & n654;
  assign n696 = pi063 & n649;
  assign n697 = ~n695 & ~n696;
  assign n698 = n694 & n697;
  assign n699 = n631 & ~n698;
  assign po067 = n691 | n699;
  assign n701 = ~pi054 & n622;
  assign n702 = ~pi053 & ~n622;
  assign n703 = ~n701 & ~n702;
  assign n704 = ~n631 & ~n703;
  assign n705 = pi081 & n656;
  assign n706 = pi059 & n651;
  assign n707 = ~n705 & ~n706;
  assign n708 = pi100 & n654;
  assign n709 = pi064 & n649;
  assign n710 = ~n708 & ~n709;
  assign n711 = n707 & n710;
  assign n712 = n631 & ~n711;
  assign po068 = n704 | n712;
  assign n714 = ~pi055 & n622;
  assign n715 = ~pi054 & ~n622;
  assign n716 = ~n714 & ~n715;
  assign n717 = ~n631 & ~n716;
  assign n718 = pi092 & n656;
  assign n719 = pi065 & n649;
  assign n720 = ~n718 & ~n719;
  assign n721 = pi090 & n654;
  assign n722 = pi071 & n651;
  assign n723 = ~n721 & ~n722;
  assign n724 = n720 & n723;
  assign n725 = n631 & ~n724;
  assign po069 = n717 | n725;
  assign n727 = ~pi057 & n622;
  assign n728 = ~pi055 & ~n622;
  assign n729 = ~n727 & ~n728;
  assign n730 = ~n631 & ~n729;
  assign n731 = pi087 & n654;
  assign n732 = pi066 & n649;
  assign n733 = ~n731 & ~n732;
  assign n734 = pi093 & n656;
  assign n735 = pi072 & n651;
  assign n736 = ~n734 & ~n735;
  assign n737 = n733 & n736;
  assign n738 = n631 & ~n737;
  assign po070 = n730 | n738;
  assign n740 = ~pi056 & n623;
  assign n741 = pi056 & ~n623;
  assign n742 = ~n740 & ~n741;
  assign n743 = n622 & ~n742;
  assign n744 = pi056 & ~n622;
  assign n745 = ~n743 & ~n744;
  assign n746 = pi118 & ~n631;
  assign po071 = ~n745 & n746;
  assign n748 = ~pi049 & n622;
  assign n749 = ~pi057 & ~n622;
  assign n750 = ~n748 & ~n749;
  assign n751 = ~n631 & ~n750;
  assign n752 = pi088 & n654;
  assign n753 = pi073 & n651;
  assign n754 = ~n752 & ~n753;
  assign n755 = pi094 & n656;
  assign n756 = pi067 & n649;
  assign n757 = ~n755 & ~n756;
  assign n758 = n754 & n757;
  assign n759 = n631 & ~n758;
  assign po072 = n751 | n759;
  assign n761 = pi048 & pi121;
  assign n762 = n273 & n761;
  assign n763 = ~pi058 & ~pi121;
  assign n764 = ~n762 & ~n763;
  assign po073 = ~pi118 | ~n764;
  assign n766 = pi059 & ~pi124;
  assign n767 = pi126 & n636;
  assign n768 = pi059 & ~n636;
  assign n769 = ~n767 & ~n768;
  assign n770 = pi124 & ~n769;
  assign po074 = n766 | n770;
  assign n772 = ~pi085 & pi122;
  assign n773 = ~pi060 & ~pi105;
  assign n774 = n772 & n773;
  assign po129 = pi060 & ~pi105;
  assign n776 = pi122 & po129;
  assign n777 = pi085 & n776;
  assign n778 = ~n774 & ~n777;
  assign n779 = pi105 & n772;
  assign n780 = ~pi060 & n779;
  assign n781 = pi060 & ~pi122;
  assign n782 = ~n780 & ~n781;
  assign po075 = ~n778 | ~n782;
  assign n784 = ~pi062 & n622;
  assign n785 = pi062 & ~n622;
  assign n786 = ~n784 & ~n785;
  assign n787 = ~n631 & ~n786;
  assign po077 = ~pi118 | n787;
  assign n789 = pi063 & ~pi124;
  assign n790 = pi125 & n635;
  assign n791 = pi063 & ~n635;
  assign n792 = ~n790 & ~n791;
  assign n793 = pi124 & ~n792;
  assign po078 = n789 | n793;
  assign n795 = pi064 & ~pi124;
  assign n796 = pi126 & n635;
  assign n797 = pi064 & ~n635;
  assign n798 = ~n796 & ~n797;
  assign n799 = pi124 & ~n798;
  assign po079 = n795 | n799;
  assign n801 = pi065 & ~pi124;
  assign n802 = pi127 & n635;
  assign n803 = pi065 & ~n635;
  assign n804 = ~n802 & ~n803;
  assign n805 = pi124 & ~n804;
  assign po080 = n801 | n805;
  assign n807 = pi066 & ~pi124;
  assign n808 = pi128 & n635;
  assign n809 = pi066 & ~n635;
  assign n810 = ~n808 & ~n809;
  assign n811 = pi124 & ~n810;
  assign po081 = n807 | n811;
  assign n813 = pi067 & ~pi124;
  assign n814 = pi129 & n635;
  assign n815 = pi067 & ~n635;
  assign n816 = ~n814 & ~n815;
  assign n817 = pi124 & ~n816;
  assign po082 = n813 | n817;
  assign n819 = pi068 & ~pi124;
  assign n820 = pi131 & n635;
  assign n821 = pi068 & ~n635;
  assign n822 = ~n820 & ~n821;
  assign n823 = pi124 & ~n822;
  assign po083 = n819 | n823;
  assign n825 = pi069 & ~pi124;
  assign n826 = pi132 & n635;
  assign n827 = pi069 & ~n635;
  assign n828 = ~n826 & ~n827;
  assign n829 = pi124 & ~n828;
  assign po084 = n825 | n829;
  assign n831 = pi070 & ~pi124;
  assign n832 = pi125 & n636;
  assign n833 = pi070 & ~n636;
  assign n834 = ~n832 & ~n833;
  assign n835 = pi124 & ~n834;
  assign po085 = n831 | n835;
  assign n837 = pi071 & ~pi124;
  assign n838 = pi127 & n636;
  assign n839 = pi071 & ~n636;
  assign n840 = ~n838 & ~n839;
  assign n841 = pi124 & ~n840;
  assign po086 = n837 | n841;
  assign n843 = pi072 & ~pi124;
  assign n844 = pi128 & n636;
  assign n845 = pi072 & ~n636;
  assign n846 = ~n844 & ~n845;
  assign n847 = pi124 & ~n846;
  assign po087 = n843 | n847;
  assign n849 = pi073 & ~pi124;
  assign n850 = pi129 & n636;
  assign n851 = pi073 & ~n636;
  assign n852 = ~n850 & ~n851;
  assign n853 = pi124 & ~n852;
  assign po088 = n849 | n853;
  assign n855 = pi074 & ~pi124;
  assign n856 = pi131 & n636;
  assign n857 = pi074 & ~n636;
  assign n858 = ~n856 & ~n857;
  assign n859 = pi124 & ~n858;
  assign po089 = n855 | n859;
  assign n861 = pi075 & ~pi124;
  assign n862 = pi132 & n636;
  assign n863 = pi075 & ~n636;
  assign n864 = ~n862 & ~n863;
  assign n865 = pi124 & ~n864;
  assign po090 = n861 | n865;
  assign n867 = ~pi103 & ~pi113;
  assign n868 = ~pi078 & ~n867;
  assign n869 = pi121 & ~n868;
  assign n870 = pi076 & ~pi121;
  assign n871 = ~n869 & ~n870;
  assign po091 = ~pi118 | ~n871;
  assign n873 = pi077 & ~n631;
  assign n874 = ~n649 & ~n651;
  assign n875 = n631 & ~n874;
  assign po092 = n873 | n875;
  assign n877 = pi078 & ~n622;
  assign n878 = ~pi052 & n622;
  assign n879 = ~n877 & ~n878;
  assign po093 = ~n631 & ~n879;
  assign n881 = pi079 & ~pi124;
  assign n882 = pi130 & n635;
  assign n883 = pi079 & ~n635;
  assign n884 = ~n882 & ~n883;
  assign n885 = pi124 & ~n884;
  assign po094 = n881 | n885;
  assign n887 = pi080 & ~pi124;
  assign n888 = pi130 & n636;
  assign n889 = pi080 & ~n636;
  assign n890 = ~n888 & ~n889;
  assign n891 = pi124 & ~n890;
  assign po095 = n887 | n891;
  assign n893 = pi081 & ~pi124;
  assign n894 = pi104 & pi112;
  assign n895 = pi126 & n894;
  assign n896 = pi081 & ~n894;
  assign n897 = ~n895 & ~n896;
  assign n898 = pi124 & ~n897;
  assign po096 = n893 | n898;
  assign n900 = pi082 & ~pi124;
  assign n901 = pi131 & n894;
  assign n902 = pi082 & ~n894;
  assign n903 = ~n901 & ~n902;
  assign n904 = pi124 & ~n903;
  assign po097 = n900 | n904;
  assign n906 = pi084 & ~pi124;
  assign n907 = pi130 & n894;
  assign n908 = pi084 & ~n894;
  assign n909 = ~n907 & ~n908;
  assign n910 = pi124 & ~n909;
  assign po099 = n906 | n910;
  assign n912 = pi085 & ~pi122;
  assign n913 = pi118 & n912;
  assign n914 = ~pi115 & pi116;
  assign n915 = pi115 & ~pi116;
  assign n916 = ~n914 & ~n915;
  assign n917 = pi118 & n916;
  assign po100 = n913 | n917;
  assign n919 = pi086 & ~pi124;
  assign n920 = ~pi104 & ~pi112;
  assign n921 = pi086 & ~n920;
  assign n922 = pi125 & n920;
  assign n923 = ~n921 & ~n922;
  assign n924 = pi124 & ~n923;
  assign po101 = n919 | n924;
  assign n926 = pi087 & ~pi124;
  assign n927 = pi087 & ~n920;
  assign n928 = pi128 & n920;
  assign n929 = ~n927 & ~n928;
  assign n930 = pi124 & ~n929;
  assign po102 = n926 | n930;
  assign n932 = pi088 & ~pi124;
  assign n933 = pi088 & ~n920;
  assign n934 = pi129 & n920;
  assign n935 = ~n933 & ~n934;
  assign n936 = pi124 & ~n935;
  assign po103 = n932 | n936;
  assign n938 = pi089 & ~pi124;
  assign n939 = pi089 & ~n920;
  assign n940 = pi132 & n920;
  assign n941 = ~n939 & ~n940;
  assign n942 = pi124 & ~n941;
  assign po104 = n938 | n942;
  assign n944 = pi090 & ~pi124;
  assign n945 = pi090 & ~n920;
  assign n946 = pi127 & n920;
  assign n947 = ~n945 & ~n946;
  assign n948 = pi124 & ~n947;
  assign po105 = n944 | n948;
  assign n950 = pi091 & ~pi124;
  assign n951 = pi125 & n894;
  assign n952 = pi091 & ~n894;
  assign n953 = ~n951 & ~n952;
  assign n954 = pi124 & ~n953;
  assign po106 = n950 | n954;
  assign n956 = pi092 & ~pi124;
  assign n957 = pi127 & n894;
  assign n958 = pi092 & ~n894;
  assign n959 = ~n957 & ~n958;
  assign n960 = pi124 & ~n959;
  assign po107 = n956 | n960;
  assign n962 = pi093 & ~pi124;
  assign n963 = pi128 & n894;
  assign n964 = pi093 & ~n894;
  assign n965 = ~n963 & ~n964;
  assign n966 = pi124 & ~n965;
  assign po108 = n962 | n966;
  assign n968 = pi094 & ~pi124;
  assign n969 = pi129 & n894;
  assign n970 = pi094 & ~n894;
  assign n971 = ~n969 & ~n970;
  assign n972 = pi124 & ~n971;
  assign po109 = n968 | n972;
  assign n974 = pi095 & ~pi124;
  assign n975 = pi132 & n894;
  assign n976 = pi095 & ~n894;
  assign n977 = ~n975 & ~n976;
  assign n978 = pi124 & ~n977;
  assign po110 = n974 | n978;
  assign n980 = pi096 & ~pi123;
  assign n981 = ~n283 & ~n288;
  assign n982 = pi123 & ~n981;
  assign po111 = n980 | n982;
  assign n984 = ~n622 & ~n631;
  assign po112 = pi097 | ~n984;
  assign n986 = pi098 & ~pi124;
  assign n987 = pi098 & ~n920;
  assign n988 = pi131 & n920;
  assign n989 = ~n987 & ~n988;
  assign n990 = pi124 & ~n989;
  assign po113 = n986 | n990;
  assign n992 = pi099 & ~pi124;
  assign n993 = pi099 & ~n920;
  assign n994 = pi130 & n920;
  assign n995 = ~n993 & ~n994;
  assign n996 = pi124 & ~n995;
  assign po114 = n992 | n996;
  assign n998 = pi100 & ~pi124;
  assign n999 = pi100 & ~n920;
  assign n1000 = pi126 & n920;
  assign n1001 = ~n999 & ~n1000;
  assign n1002 = pi124 & ~n1001;
  assign po115 = n998 | n1002;
  assign n1004 = pi062 & ~pi101;
  assign n1005 = ~pi062 & pi101;
  assign n1006 = ~n1004 & ~n1005;
  assign n1007 = n622 & ~n1006;
  assign n1008 = pi101 & ~n622;
  assign n1009 = ~n1007 & ~n1008;
  assign po116 = n746 & ~n1009;
  assign po117 = ~pi111 & ~pi114;
  assign n1012 = pi103 & ~pi121;
  assign n1013 = ~n622 & ~n1012;
  assign po118 = pi118 & ~n1013;
  assign n1015 = pi104 & ~pi124;
  assign n1016 = pi124 & ~n637;
  assign po119 = n1015 | n1016;
  assign n1018 = pi105 & ~pi122;
  assign n1019 = ~n776 & ~n1018;
  assign po120 = n780 | ~n1019;
  assign n1021 = ~pi034 & ~pi038;
  assign n1022 = pi036 & pi037;
  assign po121 = n1021 & n1022;
  assign n1024 = ~pi107 & pi123;
  assign n1025 = pi107 & ~pi123;
  assign po122 = n1024 | n1025;
  assign n1027 = pi034 & ~pi038;
  assign n1028 = pi036 & n1027;
  assign po123 = pi037 | ~n1028;
  assign n1030 = pi109 & ~n631;
  assign n1031 = ~pi109 & n631;
  assign po124 = n1030 | n1031;
  assign n1033 = pi058 & ~pi113;
  assign po125 = ~pi120 & n1033;
  assign n1035 = pi112 & ~pi124;
  assign n1036 = ~pi112 & pi124;
  assign po127 = n1035 | n1036;
  assign n1038 = pi047 & ~pi056;
  assign po128 = ~n1004 | ~n1038;
  assign po012 = 1'b1;
  assign po126 = ~pi114;
  assign po000 = pi076;
  assign po001 = pi061;
  assign po013 = pi117;
  assign po015 = pi118;
  assign po098 = pi106;
  assign po130 = pi116;
  assign po131 = pi119;
endmodule


