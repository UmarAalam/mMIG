//Written by the Majority Logic Package Thu Apr 30 13:14:51 2015
module top (
            pi000, pi001, pi002, pi003, pi004, pi005, pi006, pi007, pi008, pi009, pi010, pi011, pi012, pi013, pi014, pi015, pi016, pi017, pi018, pi019, pi020, pi021, pi022, pi023, pi024, pi025, pi026, pi027, pi028, pi029, pi030, pi031, pi032, pi033, pi034, pi035, pi036, pi037, pi038, pi039, pi040, pi041, pi042, pi043, pi044, pi045, pi046, pi047, pi048, pi049, pi050, pi051, pi052, pi053, pi054, pi055, pi056, pi057, pi058, pi059, pi060, pi061, pi062, pi063, pi064, pi065, pi066, pi067, pi068, pi069, pi070, pi071, pi072, pi073, pi074, pi075, pi076, pi077, pi078, pi079, pi080, pi081, pi082, pi083, pi084, pi085, pi086, pi087, pi088, pi089, pi090, pi091, pi092, pi093, pi094, pi095, pi096, pi097, pi098, pi099, pi100, pi101, pi102, pi103, pi104, pi105, pi106, pi107, pi108, pi109, pi110, pi111, pi112, pi113, pi114, pi115, pi116, pi117, pi118, pi119, pi120, pi121, pi122, pi123, pi124, pi125, pi126, pi127, pi128, pi129, pi130, pi131, pi132, 
            po000, po001, po002, po003, po004, po005, po006, po007, po008, po009, po010, po011, po012, po013, po014, po015, po016, po017, po018, po019, po020, po021, po022, po023, po024, po025, po026, po027, po028, po029, po030, po031, po032, po033, po034, po035, po036, po037, po038, po039, po040, po041, po042, po043, po044, po045, po046, po047, po048, po049, po050, po051, po052, po053, po054, po055, po056, po057, po058, po059, po060, po061, po062, po063, po064, po065, po066, po067, po068, po069, po070, po071, po072, po073, po074, po075, po076, po077, po078, po079, po080, po081, po082, po083, po084, po085, po086, po087, po088, po089, po090, po091, po092, po093, po094, po095, po096, po097, po098, po099, po100, po101, po102, po103, po104, po105, po106, po107, po108, po109, po110, po111, po112, po113, po114, po115, po116, po117, po118, po119, po120, po121, po122, po123, po124, po125, po126, po127, po128, po129, po130, po131);
input pi000, pi001, pi002, pi003, pi004, pi005, pi006, pi007, pi008, pi009, pi010, pi011, pi012, pi013, pi014, pi015, pi016, pi017, pi018, pi019, pi020, pi021, pi022, pi023, pi024, pi025, pi026, pi027, pi028, pi029, pi030, pi031, pi032, pi033, pi034, pi035, pi036, pi037, pi038, pi039, pi040, pi041, pi042, pi043, pi044, pi045, pi046, pi047, pi048, pi049, pi050, pi051, pi052, pi053, pi054, pi055, pi056, pi057, pi058, pi059, pi060, pi061, pi062, pi063, pi064, pi065, pi066, pi067, pi068, pi069, pi070, pi071, pi072, pi073, pi074, pi075, pi076, pi077, pi078, pi079, pi080, pi081, pi082, pi083, pi084, pi085, pi086, pi087, pi088, pi089, pi090, pi091, pi092, pi093, pi094, pi095, pi096, pi097, pi098, pi099, pi100, pi101, pi102, pi103, pi104, pi105, pi106, pi107, pi108, pi109, pi110, pi111, pi112, pi113, pi114, pi115, pi116, pi117, pi118, pi119, pi120, pi121, pi122, pi123, pi124, pi125, pi126, pi127, pi128, pi129, pi130, pi131, pi132;
output po000, po001, po002, po003, po004, po005, po006, po007, po008, po009, po010, po011, po012, po013, po014, po015, po016, po017, po018, po019, po020, po021, po022, po023, po024, po025, po026, po027, po028, po029, po030, po031, po032, po033, po034, po035, po036, po037, po038, po039, po040, po041, po042, po043, po044, po045, po046, po047, po048, po049, po050, po051, po052, po053, po054, po055, po056, po057, po058, po059, po060, po061, po062, po063, po064, po065, po066, po067, po068, po069, po070, po071, po072, po073, po074, po075, po076, po077, po078, po079, po080, po081, po082, po083, po084, po085, po086, po087, po088, po089, po090, po091, po092, po093, po094, po095, po096, po097, po098, po099, po100, po101, po102, po103, po104, po105, po106, po107, po108, po109, po110, po111, po112, po113, po114, po115, po116, po117, po118, po119, po120, po121, po122, po123, po124, po125, po126, po127, po128, po129, po130, po131;
wire one, v0, v1, v2, v3, v4, v5, v6, v7, v8, v9, v10, v11, v12, v13, v14, v15, v16, v17, v18, v19, v20, v21, v22, v23, v24, v25, v26, v27, v28, v29, v30, v31, v32, v33, v34, v35, v36, v37, v38, v39, v40, v41, v42, v43, v44, v45, v46, v47, v48, v49, v50, v51, v52, v53, v54, v55, v56, v57, v58, v59, v60, v61, v62, v63, v64, v65, v66, v67, v68, v69, v70, v71, v72, v73, v74, v75, v76, v77, v78, v79, v80, v81, v82, v83, v84, v85, v86, v87, v88, v89, v90, v91, v92, v93, v94, v95, v96, v97, v98, v99, v100, v101, v102, v103, v104, v105, v106, v107, v108, v109, v110, v111, v112, v113, v114, v115, v116, v117, v118, v119, v120, v121, v122, v123, v124, v125, v126, v127, v128, v129, v130, v131, v132, v133, v134, v135, v136, v137, v138, v139, v140, v141, v142, v143, v144, v145, v146, v147, v148, v149, v150, v151, v152, v153, v154, v155, v156, v157, v158, v159, v160, v161, v162, v163, v164, v165, v166, v167, 
 w0, w1, w2, w3, w4, w5, w6, w7, w8, w9, w10, w11, w12, w13, w14, w15, w16, w17, w18, w19, w20, w21, w22, w23, w24, w25, w26, w27, w28, w29, w30, w31, w32, w33, w34, w35, w36, w37, w38, w39, w40, w41, w42, w43, w44, w45, w46, w47, w48, w49, w50, w51, w52, w53, w54, w55, w56, w57, w58, w59, w60, w61, w62, w63, w64, w65, w66, w67, w68, w69, w70, w71, w72, w73, w74, w75, w76, w77, w78, w79, w80, w81, w82, w83, w84, w85, w86, w87, w88, w89, w90, w91, w92, w93, w94, w95, w96, w97, w98, w99, w100, w101, w102, w103, w104, w105, w106, w107, w108, w109, w110, w111, w112, w113, w114, w115, w116, w117, w118, w119, w120, w121, w122, w123, w124, w125, w126, w127, w128, w129, w130, w131, w132, w133, w134, w135, w136, w137, w138, w139, w140, w141, w142, w143, w144, w145, w146, w147, w148, w149, w150, w151, w152, w153, w154, w155, w156, w157, w158, w159, w160, w161, w162, w163, w164, w165, w166, w167, w168, w169, w170, w171, w172, w173, w174, w175, w176, w177, w178, w179, w180, w181, w182, w183, w184, w185, w186, w187, w188, w189, w190, w191, w192, w193, w194, w195, w196, w197, w198, w199, w200, w201, w202, w203, w204, w205, w206, w207, w208, w209, w210, w211, w212, w213, w214, w215, w216, w217, w218, w219, w220, w221, w222, w223, w224, w225, w226, w227, w228, w229, w230, w231, w232, w233, w234, w235, w236, w237, w238, w239, w240, w241, w242, w243, w244, w245, w246, w247, w248, w249, w250, w251, w252, w253, w254, w255, w256, w257, w258, w259, w260, w261, w262, w263, w264, w265, w266, w267, w268, w269, w270, w271, w272, w273, w274, w275, w276, w277, w278, w279, w280, w281, w282, w283, w284, w285, w286, w287, w288, w289, w290, w291, w292, w293, w294, w295, w296, w297, w298, w299, w300, w301, w302, w303, w304, w305, w306, w307, w308, w309, w310, w311, w312, w313, w314, w315, w316, w317, w318, w319, w320, w321, w322, w323, w324, w325, w326, w327, w328, w329, w330, w331, w332, w333, w334, w335, w336, w337, w338, w339, w340, w341, w342, w343, w344, w345, w346, w347, w348, w349, w350, w351, w352, w353, w354, w355, w356, w357, w358, w359, w360, w361, w362, w363, w364, w365, w366, w367, w368, w369, w370, w371, w372, w373, w374, w375, w376, w377, w378, w379, w380, w381, w382, w383, w384, w385, w386, w387, w388, w389, w390, w391, w392, w393, w394, w395, w396, w397, w398, w399, w400, w401, w402, w403, w404, w405, w406, w407, w408, w409, w410, w411, w412, w413, w414, w415, w416, w417, w418, w419, w420, w421, w422, w423, w424, w425, w426, w427, w428, w429, w430, w431, w432, w433, w434, w435, w436, w437, w438, w439, w440, w441, w442, w443, w444, w445, w446, w447, w448, w449, w450, w451, w452, w453, w454, w455, w456, w457, w458, w459, w460, w461, w462, w463, w464, w465, w466, w467, w468, w469, w470, w471, w472, w473, w474, w475, w476, w477, w478, w479, w480, w481, w482, w483, w484, w485, w486, w487, w488, w489, w490, w491, w492, w493, w494, w495, w496, w497, w498, w499, w500, w501, w502, w503, w504, w505, w506, w507, w508, w509, w510, w511, w512, w513, w514, w515, w516, w517, w518, w519, w520, w521, w522, w523, w524, w525, w526, w527, w528, w529, w530, w531, w532, w533, w534, w535, w536, w537, w538, w539, w540, w541, w542, w543, w544, w545, w546, w547, w548, w549, w550, w551, w552, w553, w554, w555, w556, w557, w558, w559, w560, w561, w562, w563, w564, w565, w566, w567, w568, w569, w570, w571, w572, w573, w574, w575, w576, w577, w578, w579, w580, w581, w582, w583, w584, w585, w586, w587, w588, w589, w590, w591, w592, w593, w594, w595, w596, w597, w598, w599, w600, w601, w602, w603, w604, w605, w606, w607, w608, w609, w610, w611, w612, w613, w614, w615, w616, w617, w618, w619, w620;
assign w0 = ~pi109 & pi112;
assign w1 = pi109 & ~pi112;
assign w2 = pi077 & ~pi104;
assign w3 = ~pi077 & pi104;
assign v0 = ~(w2 | w3);
assign w4 = v0;
assign w5 = ~w1 & w4;
assign w6 = ~w0 & w5;
assign w7 = ~pi048 & w6;
assign w8 = ~pi001 & pi107;
assign w9 = pi035 & ~pi096;
assign w10 = ~pi035 & pi096;
assign v1 = ~(w9 | w10);
assign w11 = v1;
assign w12 = ~w8 & w11;
assign w13 = pi001 & ~pi107;
assign v2 = ~(pi000 | w13);
assign w14 = v2;
assign w15 = w12 & w14;
assign w16 = pi096 & pi107;
assign w17 = pi018 & w16;
assign v3 = ~(pi096 | pi107);
assign w18 = v3;
assign w19 = pi026 & w18;
assign v4 = ~(w17 | w19);
assign w20 = v4;
assign w21 = ~pi096 & pi107;
assign w22 = pi012 & w21;
assign w23 = pi096 & ~pi107;
assign w24 = pi004 & w23;
assign v5 = ~(w22 | w24);
assign w25 = v5;
assign w26 = w20 & w25;
assign w27 = pi005 & w23;
assign w28 = pi027 & w18;
assign v6 = ~(w27 | w28);
assign w29 = v6;
assign w30 = pi019 & w16;
assign w31 = pi013 & w21;
assign v7 = ~(w30 | w31);
assign w32 = v7;
assign w33 = w29 & w32;
assign w34 = pi028 & w18;
assign w35 = pi020 & w16;
assign v8 = ~(w34 | w35);
assign w36 = v8;
assign w37 = pi014 & w21;
assign w38 = pi006 & w23;
assign v9 = ~(w37 | w38);
assign w39 = v9;
assign w40 = w36 & w39;
assign w41 = pi021 & w16;
assign w42 = pi015 & w21;
assign v10 = ~(w41 | w42);
assign w43 = v10;
assign w44 = pi007 & w23;
assign w45 = pi029 & w18;
assign v11 = ~(w44 | w45);
assign w46 = v11;
assign w47 = w43 & w46;
assign w48 = pi022 & w16;
assign w49 = pi008 & w23;
assign v12 = ~(w48 | w49);
assign w50 = v12;
assign w51 = pi016 & w21;
assign w52 = pi030 & w18;
assign v13 = ~(w51 | w52);
assign w53 = v13;
assign w54 = w50 & w53;
assign w55 = pi031 & w18;
assign w56 = pi017 & w21;
assign v14 = ~(w55 | w56);
assign w57 = v14;
assign w58 = pi023 & w16;
assign w59 = pi009 & w23;
assign v15 = ~(w58 | w59);
assign w60 = v15;
assign w61 = w57 & w60;
assign w62 = pi032 & w18;
assign w63 = pi002 & w21;
assign v16 = ~(w62 | w63);
assign w64 = v16;
assign w65 = pi010 & w23;
assign w66 = pi024 & w16;
assign v17 = ~(w65 | w66);
assign w67 = v17;
assign w68 = w64 & w67;
assign w69 = pi003 & w21;
assign w70 = pi025 & w16;
assign v18 = ~(w69 | w70);
assign w71 = v18;
assign w72 = pi033 & w18;
assign w73 = pi011 & w23;
assign v19 = ~(w72 | w73);
assign w74 = v19;
assign w75 = w71 & w74;
assign w76 = pi000 & ~pi123;
assign v20 = ~(w11 | w13);
assign w77 = v20;
assign w78 = pi083 & pi106;
assign w79 = (w78 & ~w11) | (w78 & w548) | (~w11 & w548);
assign w80 = ~w77 & w79;
assign v21 = ~(w76 | w80);
assign w81 = v21;
assign w82 = pi118 & ~w81;
assign w83 = pi000 & ~w13;
assign w84 = w12 & w83;
assign w85 = (w78 & ~w12) | (w78 & w542) | (~w12 & w542);
assign v22 = ~(pi001 | w85);
assign w86 = v22;
assign w87 = pi001 & w85;
assign v23 = ~(w86 | w87);
assign w88 = v23;
assign w89 = w85 & w543;
assign w90 = (pi002 & ~w85) | (pi002 & w549) | (~w85 & w549);
assign w91 = w85 & w550;
assign v24 = ~(w90 | w91);
assign w92 = v24;
assign w93 = (pi003 & ~w85) | (pi003 & w551) | (~w85 & w551);
assign w94 = w85 & w552;
assign v25 = ~(w93 | w94);
assign w95 = v25;
assign w96 = ~pi001 & pi035;
assign w97 = (pi004 & ~w85) | (pi004 & w553) | (~w85 & w553);
assign w98 = w85 & w554;
assign v26 = ~(w97 | w98);
assign w99 = v26;
assign w100 = (pi005 & ~w85) | (pi005 & w555) | (~w85 & w555);
assign w101 = w85 & w556;
assign v27 = ~(w100 | w101);
assign w102 = v27;
assign w103 = (pi006 & ~w85) | (pi006 & w557) | (~w85 & w557);
assign w104 = w85 & w558;
assign v28 = ~(w103 | w104);
assign w105 = v28;
assign w106 = (pi007 & ~w85) | (pi007 & w559) | (~w85 & w559);
assign w107 = w85 & w560;
assign v29 = ~(w106 | w107);
assign w108 = v29;
assign w109 = (pi008 & ~w85) | (pi008 & w561) | (~w85 & w561);
assign w110 = w85 & w562;
assign v30 = ~(w109 | w110);
assign w111 = v30;
assign w112 = (pi009 & ~w85) | (pi009 & w563) | (~w85 & w563);
assign w113 = w85 & w564;
assign v31 = ~(w112 | w113);
assign w114 = v31;
assign w115 = (pi010 & ~w85) | (pi010 & w565) | (~w85 & w565);
assign w116 = w85 & w566;
assign v32 = ~(w115 | w116);
assign w117 = v32;
assign w118 = (pi011 & ~w85) | (pi011 & w567) | (~w85 & w567);
assign w119 = w85 & w568;
assign v33 = ~(w118 | w119);
assign w120 = v33;
assign w121 = (pi012 & ~w85) | (pi012 & w569) | (~w85 & w569);
assign w122 = w85 & w570;
assign v34 = ~(w121 | w122);
assign w123 = v34;
assign w124 = (pi013 & ~w85) | (pi013 & w571) | (~w85 & w571);
assign w125 = w85 & w572;
assign v35 = ~(w124 | w125);
assign w126 = v35;
assign w127 = (pi014 & ~w85) | (pi014 & w573) | (~w85 & w573);
assign w128 = w85 & w574;
assign v36 = ~(w127 | w128);
assign w129 = v36;
assign w130 = (pi015 & ~w85) | (pi015 & w575) | (~w85 & w575);
assign w131 = w85 & w576;
assign v37 = ~(w130 | w131);
assign w132 = v37;
assign w133 = (pi016 & ~w85) | (pi016 & w577) | (~w85 & w577);
assign w134 = w85 & w578;
assign v38 = ~(w133 | w134);
assign w135 = v38;
assign w136 = (pi017 & ~w85) | (pi017 & w579) | (~w85 & w579);
assign w137 = w85 & w580;
assign v39 = ~(w136 | w137);
assign w138 = v39;
assign w139 = (pi018 & ~w85) | (pi018 & w581) | (~w85 & w581);
assign w140 = w85 & w582;
assign v40 = ~(w139 | w140);
assign w141 = v40;
assign w142 = (pi019 & ~w85) | (pi019 & w583) | (~w85 & w583);
assign w143 = w85 & w584;
assign v41 = ~(w142 | w143);
assign w144 = v41;
assign w145 = (pi020 & ~w85) | (pi020 & w585) | (~w85 & w585);
assign w146 = w85 & w586;
assign v42 = ~(w145 | w146);
assign w147 = v42;
assign w148 = (pi021 & ~w85) | (pi021 & w587) | (~w85 & w587);
assign w149 = w85 & w588;
assign v43 = ~(w148 | w149);
assign w150 = v43;
assign w151 = (pi022 & ~w85) | (pi022 & w589) | (~w85 & w589);
assign w152 = w85 & w590;
assign v44 = ~(w151 | w152);
assign w153 = v44;
assign w154 = (pi023 & ~w85) | (pi023 & w591) | (~w85 & w591);
assign w155 = w85 & w592;
assign v45 = ~(w154 | w155);
assign w156 = v45;
assign w157 = (pi024 & ~w85) | (pi024 & w593) | (~w85 & w593);
assign w158 = w85 & w594;
assign v46 = ~(w157 | w158);
assign w159 = v46;
assign w160 = (pi025 & ~w85) | (pi025 & w595) | (~w85 & w595);
assign w161 = w85 & w596;
assign v47 = ~(w160 | w161);
assign w162 = v47;
assign v48 = ~(pi001 | pi035);
assign w163 = v48;
assign w164 = (pi026 & ~w85) | (pi026 & w597) | (~w85 & w597);
assign w165 = w85 & w598;
assign v49 = ~(w164 | w165);
assign w166 = v49;
assign w167 = (pi027 & ~w85) | (pi027 & w599) | (~w85 & w599);
assign w168 = w85 & w600;
assign v50 = ~(w167 | w168);
assign w169 = v50;
assign w170 = (pi028 & ~w85) | (pi028 & w601) | (~w85 & w601);
assign w171 = w85 & w602;
assign v51 = ~(w170 | w171);
assign w172 = v51;
assign w173 = (pi029 & ~w85) | (pi029 & w603) | (~w85 & w603);
assign w174 = w85 & w604;
assign v52 = ~(w173 | w174);
assign w175 = v52;
assign w176 = (pi030 & ~w85) | (pi030 & w605) | (~w85 & w605);
assign w177 = w85 & w606;
assign v53 = ~(w176 | w177);
assign w178 = v53;
assign w179 = (pi031 & ~w85) | (pi031 & w607) | (~w85 & w607);
assign w180 = w85 & w608;
assign v54 = ~(w179 | w180);
assign w181 = v54;
assign w182 = (pi032 & ~w85) | (pi032 & w609) | (~w85 & w609);
assign w183 = w85 & w610;
assign v55 = ~(w182 | w183);
assign w184 = v55;
assign w185 = (pi033 & ~w85) | (pi033 & w611) | (~w85 & w611);
assign w186 = w85 & w612;
assign v56 = ~(w185 | w186);
assign w187 = v56;
assign w188 = pi102 & pi108;
assign w189 = pi037 & w188;
assign w190 = w188 & w545;
assign w191 = (~pi034 & ~w188) | (~pi034 & w619) | (~w188 & w619);
assign v57 = ~(pi115 | pi116);
assign w192 = v57;
assign w193 = ~pi108 & w192;
assign v58 = ~(w191 | w193);
assign w194 = v58;
assign w195 = ~w190 & w194;
assign w196 = pi118 & ~w195;
assign w197 = (pi035 & ~w85) | (pi035 & w96) | (~w85 & w96);
assign v59 = ~(w89 | w197);
assign w198 = v59;
assign w199 = pi038 & w190;
assign w200 = w190 & w620;
assign w201 = (~pi036 & ~w190) | (~pi036 & w613) | (~w190 & w613);
assign v60 = ~(w193 | w201);
assign w202 = v60;
assign w203 = ~w200 & w202;
assign w204 = pi118 & ~w203;
assign w205 = pi118 & ~w193;
assign v61 = ~(pi037 | w188);
assign w206 = v61;
assign v62 = ~(w189 | w206);
assign w207 = v62;
assign w208 = w205 & w207;
assign v63 = ~(pi038 | w190);
assign w209 = v63;
assign w210 = ~w199 & w205;
assign w211 = ~w209 & w210;
assign w212 = pi039 & ~w188;
assign w213 = pi042 & w188;
assign v64 = ~(w212 | w213);
assign w214 = v64;
assign w215 = pi040 & ~w188;
assign w216 = pi116 & w188;
assign v65 = ~(w215 | w216);
assign w217 = v65;
assign w218 = pi041 & ~w188;
assign w219 = pi039 & w188;
assign v66 = ~(w218 | w219);
assign w220 = v66;
assign w221 = pi042 & ~w188;
assign w222 = pi043 & w188;
assign v67 = ~(w221 | w222);
assign w223 = v67;
assign w224 = pi043 & ~w188;
assign w225 = pi044 & w188;
assign v68 = ~(w224 | w225);
assign w226 = v68;
assign w227 = pi044 & ~w188;
assign w228 = pi046 & w188;
assign v69 = ~(w227 | w228);
assign w229 = v69;
assign w230 = pi045 & ~w188;
assign w231 = pi040 & w188;
assign v70 = ~(w230 | w231);
assign w232 = v70;
assign w233 = pi046 & ~w188;
assign w234 = pi045 & w188;
assign v71 = ~(w233 | w234);
assign w235 = v71;
assign w236 = pi113 & pi121;
assign w237 = pi062 & w236;
assign w238 = w236 & w546;
assign w239 = pi056 & w238;
assign w240 = w238 & w614;
assign w241 = pi110 & pi121;
assign w242 = (w238 & w615) | (w238 & w616) | (w615 & w616);
assign w243 = ~w240 & w242;
assign w244 = pi118 & ~w243;
assign w245 = pi118 & ~w241;
assign w246 = ~pi048 & w245;
assign v72 = ~(w0 | w4);
assign w247 = v72;
assign w248 = pi118 & pi124;
assign w249 = (w248 & ~w4) | (w248 & w617) | (~w4 & w617);
assign w250 = ~w247 & w249;
assign v73 = ~(w246 | w250);
assign w251 = v73;
assign w252 = pi077 & ~pi109;
assign w253 = pi080 & w252;
assign w254 = pi077 & pi109;
assign w255 = pi084 & w254;
assign v74 = ~(w253 | w255);
assign w256 = v74;
assign v75 = ~(pi077 | pi109);
assign w257 = v75;
assign w258 = pi099 & w257;
assign w259 = ~pi077 & pi109;
assign w260 = pi079 & w259;
assign v76 = ~(w258 | w260);
assign w261 = v76;
assign w262 = w256 & w261;
assign w263 = w241 & ~w262;
assign w264 = pi049 & ~w236;
assign w265 = pi050 & w236;
assign v77 = ~(w241 | w265);
assign w266 = v77;
assign w267 = ~w264 & w266;
assign v78 = ~(w263 | w267);
assign w268 = v78;
assign w269 = pi082 & w254;
assign w270 = pi068 & w259;
assign v79 = ~(w269 | w270);
assign w271 = v79;
assign w272 = pi074 & w252;
assign w273 = pi098 & w257;
assign v80 = ~(w272 | w273);
assign w274 = v80;
assign w275 = w271 & w274;
assign w276 = w241 & ~w275;
assign w277 = pi050 & ~w236;
assign w278 = pi051 & w236;
assign v81 = ~(w241 | w278);
assign w279 = v81;
assign w280 = ~w277 & w279;
assign v82 = ~(w276 | w280);
assign w281 = v82;
assign w282 = ~pi097 & w236;
assign v83 = ~(w241 | w282);
assign w283 = v83;
assign w284 = pi051 & ~w236;
assign w285 = w283 & ~w284;
assign w286 = pi089 & w257;
assign w287 = pi095 & w254;
assign v84 = ~(w286 | w287);
assign w288 = v84;
assign w289 = pi069 & w259;
assign w290 = pi075 & w252;
assign v85 = ~(w289 | w290);
assign w291 = v85;
assign w292 = w288 & w291;
assign w293 = w241 & ~w292;
assign v86 = ~(w285 | w293);
assign w294 = v86;
assign w295 = pi070 & w252;
assign w296 = pi063 & w259;
assign v87 = ~(w295 | w296);
assign w297 = v87;
assign w298 = pi091 & w254;
assign w299 = pi086 & w257;
assign v88 = ~(w298 | w299);
assign w300 = v88;
assign w301 = w297 & w300;
assign w302 = w241 & ~w301;
assign w303 = pi052 & ~w236;
assign w304 = pi053 & w236;
assign v89 = ~(w241 | w304);
assign w305 = v89;
assign w306 = ~w303 & w305;
assign v90 = ~(w302 | w306);
assign w307 = v90;
assign w308 = pi064 & w259;
assign w309 = pi081 & w254;
assign v91 = ~(w308 | w309);
assign w310 = v91;
assign w311 = pi100 & w257;
assign w312 = pi059 & w252;
assign v92 = ~(w311 | w312);
assign w313 = v92;
assign w314 = w310 & w313;
assign w315 = w241 & ~w314;
assign w316 = pi053 & ~w236;
assign w317 = pi054 & w236;
assign v93 = ~(w241 | w317);
assign w318 = v93;
assign w319 = ~w316 & w318;
assign v94 = ~(w315 | w319);
assign w320 = v94;
assign w321 = pi071 & w252;
assign w322 = pi092 & w254;
assign v95 = ~(w321 | w322);
assign w323 = v95;
assign w324 = pi065 & w259;
assign w325 = pi090 & w257;
assign v96 = ~(w324 | w325);
assign w326 = v96;
assign w327 = w323 & w326;
assign w328 = w241 & ~w327;
assign w329 = pi054 & ~w236;
assign w330 = pi055 & w236;
assign v97 = ~(w241 | w330);
assign w331 = v97;
assign w332 = ~w329 & w331;
assign v98 = ~(w328 | w332);
assign w333 = v98;
assign w334 = pi093 & w254;
assign w335 = pi066 & w259;
assign v99 = ~(w334 | w335);
assign w336 = v99;
assign w337 = pi087 & w257;
assign w338 = pi072 & w252;
assign v100 = ~(w337 | w338);
assign w339 = v100;
assign w340 = w336 & w339;
assign w341 = w241 & ~w340;
assign w342 = pi055 & ~w236;
assign w343 = pi057 & w236;
assign v101 = ~(w241 | w343);
assign w344 = v101;
assign w345 = ~w342 & w344;
assign v102 = ~(w341 | w345);
assign w346 = v102;
assign v103 = ~(pi056 | w238);
assign w347 = v103;
assign w348 = ~w239 & w245;
assign w349 = ~w347 & w348;
assign w350 = pi094 & w254;
assign w351 = pi067 & w259;
assign v104 = ~(w350 | w351);
assign w352 = v104;
assign w353 = pi088 & w257;
assign w354 = pi073 & w252;
assign v105 = ~(w353 | w354);
assign w355 = v105;
assign w356 = w352 & w355;
assign w357 = w241 & ~w356;
assign w358 = pi057 & ~w236;
assign w359 = pi049 & w236;
assign v106 = ~(w241 | w359);
assign w360 = v106;
assign w361 = ~w358 & w360;
assign v107 = ~(w357 | w361);
assign w362 = v107;
assign w363 = pi048 & pi121;
assign w364 = w5 & w618;
assign v108 = ~(pi058 | pi121);
assign w365 = v108;
assign w366 = pi118 & ~w365;
assign w367 = ~w364 & w366;
assign w368 = ~pi112 & pi124;
assign w369 = pi104 & w368;
assign w370 = pi059 & ~w369;
assign w371 = pi126 & w369;
assign v109 = ~(w370 | w371);
assign w372 = v109;
assign v110 = ~(pi060 | pi122);
assign w373 = v110;
assign v111 = ~(pi060 | pi085);
assign w374 = v111;
assign w375 = pi122 & ~w374;
assign w376 = pi060 & ~pi105;
assign w377 = pi085 & w376;
assign w378 = w375 & ~w377;
assign v112 = ~(w373 | w378);
assign w379 = v112;
assign v113 = ~(pi062 | w236);
assign w380 = v113;
assign v114 = ~(w237 | w241);
assign w381 = v114;
assign w382 = ~w380 & w381;
assign w383 = pi118 & ~w382;
assign w384 = ~pi104 & pi112;
assign w385 = pi124 & w384;
assign w386 = pi063 & ~w385;
assign w387 = pi124 & pi125;
assign w388 = w384 & w387;
assign v115 = ~(w386 | w388);
assign w389 = v115;
assign w390 = pi064 & ~w385;
assign w391 = pi124 & pi126;
assign w392 = w384 & w391;
assign v116 = ~(w390 | w392);
assign w393 = v116;
assign w394 = pi065 & ~w385;
assign w395 = pi124 & pi127;
assign w396 = w384 & w395;
assign v117 = ~(w394 | w396);
assign w397 = v117;
assign w398 = pi066 & ~w385;
assign w399 = pi124 & pi128;
assign w400 = w384 & w399;
assign v118 = ~(w398 | w400);
assign w401 = v118;
assign w402 = pi067 & ~w385;
assign w403 = pi124 & pi129;
assign w404 = w384 & w403;
assign v119 = ~(w402 | w404);
assign w405 = v119;
assign w406 = pi068 & ~w385;
assign w407 = pi124 & pi131;
assign w408 = w384 & w407;
assign v120 = ~(w406 | w408);
assign w409 = v120;
assign w410 = pi069 & ~w385;
assign w411 = pi124 & pi132;
assign w412 = w384 & w411;
assign v121 = ~(w410 | w412);
assign w413 = v121;
assign w414 = pi070 & ~w369;
assign w415 = pi125 & w369;
assign v122 = ~(w414 | w415);
assign w416 = v122;
assign w417 = pi071 & ~w369;
assign w418 = pi127 & w369;
assign v123 = ~(w417 | w418);
assign w419 = v123;
assign w420 = pi072 & ~w369;
assign w421 = pi128 & w369;
assign v124 = ~(w420 | w421);
assign w422 = v124;
assign w423 = pi073 & ~w369;
assign w424 = pi129 & w369;
assign v125 = ~(w423 | w424);
assign w425 = v125;
assign w426 = pi074 & ~w369;
assign w427 = pi131 & w369;
assign v126 = ~(w426 | w427);
assign w428 = v126;
assign w429 = pi075 & ~w369;
assign w430 = pi132 & w369;
assign v127 = ~(w429 | w430);
assign w431 = v127;
assign v128 = ~(pi103 | pi113);
assign w432 = v128;
assign v129 = ~(pi078 | w432);
assign w433 = v129;
assign w434 = pi121 & ~w433;
assign w435 = pi076 & ~pi121;
assign w436 = pi118 & ~w435;
assign w437 = ~w434 & w436;
assign w438 = pi109 & w241;
assign v130 = ~(pi077 | w438);
assign w439 = v130;
assign w440 = pi077 & w438;
assign v131 = ~(w439 | w440);
assign w441 = v131;
assign w442 = pi052 & w236;
assign v132 = ~(pi078 | w236);
assign w443 = v132;
assign v133 = ~(w241 | w443);
assign w444 = v133;
assign w445 = ~w442 & w444;
assign w446 = pi079 & ~w385;
assign w447 = pi124 & pi130;
assign w448 = w384 & w447;
assign v134 = ~(w446 | w448);
assign w449 = v134;
assign w450 = pi080 & ~w369;
assign w451 = pi130 & w369;
assign v135 = ~(w450 | w451);
assign w452 = v135;
assign w453 = pi104 & pi112;
assign w454 = pi124 & w453;
assign w455 = pi081 & ~w454;
assign w456 = w391 & w453;
assign v136 = ~(w455 | w456);
assign w457 = v136;
assign w458 = pi082 & ~w454;
assign w459 = w407 & w453;
assign v137 = ~(w458 | w459);
assign w460 = v137;
assign w461 = pi084 & ~w454;
assign w462 = w447 & w453;
assign v138 = ~(w461 | w462);
assign w463 = v138;
assign w464 = pi085 & ~pi122;
assign w465 = pi115 & pi116;
assign v139 = ~(w192 | w465);
assign w466 = v139;
assign w467 = ~w464 & w466;
assign w468 = pi118 & ~w467;
assign w469 = ~pi104 & w368;
assign w470 = pi086 & ~w469;
assign w471 = pi125 & w469;
assign v140 = ~(w470 | w471);
assign w472 = v140;
assign w473 = pi087 & ~w469;
assign w474 = pi128 & w469;
assign v141 = ~(w473 | w474);
assign w475 = v141;
assign w476 = pi088 & ~w469;
assign w477 = pi129 & w469;
assign v142 = ~(w476 | w477);
assign w478 = v142;
assign w479 = pi089 & ~w469;
assign w480 = pi132 & w469;
assign v143 = ~(w479 | w480);
assign w481 = v143;
assign w482 = pi090 & ~w469;
assign w483 = pi127 & w469;
assign v144 = ~(w482 | w483);
assign w484 = v144;
assign w485 = pi091 & ~w454;
assign w486 = w387 & w453;
assign v145 = ~(w485 | w486);
assign w487 = v145;
assign w488 = pi092 & ~w454;
assign w489 = w395 & w453;
assign v146 = ~(w488 | w489);
assign w490 = v146;
assign w491 = pi093 & ~w454;
assign w492 = w399 & w453;
assign v147 = ~(w491 | w492);
assign w493 = v147;
assign w494 = pi094 & ~w454;
assign w495 = w403 & w453;
assign v148 = ~(w494 | w495);
assign w496 = v148;
assign w497 = pi095 & ~w454;
assign w498 = w411 & w453;
assign v149 = ~(w497 | w498);
assign w499 = v149;
assign w500 = pi107 & pi123;
assign w501 = pi096 & ~w500;
assign w502 = ~pi096 & w500;
assign v150 = ~(w501 | w502);
assign w503 = v150;
assign w504 = ~pi097 & w283;
assign w505 = pi098 & ~w469;
assign w506 = pi131 & w469;
assign v151 = ~(w505 | w506);
assign w507 = v151;
assign w508 = pi099 & ~w469;
assign w509 = pi130 & w469;
assign v152 = ~(w508 | w509);
assign w510 = v152;
assign w511 = pi100 & ~w469;
assign w512 = pi126 & w469;
assign v153 = ~(w511 | w512);
assign w513 = v153;
assign v154 = ~(pi101 | w237);
assign w514 = v154;
assign w515 = ~w238 & w245;
assign w516 = ~w514 & w515;
assign v155 = ~(pi111 | pi114);
assign w517 = v155;
assign w518 = pi103 & ~pi121;
assign v156 = ~(w236 | w518);
assign w519 = v156;
assign w520 = pi118 & ~w519;
assign w521 = pi104 & ~w454;
assign v157 = ~(w385 | w521);
assign w522 = v157;
assign w523 = pi122 & w376;
assign w524 = pi105 & ~w375;
assign v158 = ~(w523 | w524);
assign w525 = v158;
assign w526 = pi036 & ~pi038;
assign w527 = ~pi034 & pi037;
assign w528 = w526 & w527;
assign v159 = ~(pi107 | pi123);
assign w529 = v159;
assign v160 = ~(w500 | w529);
assign w530 = v160;
assign w531 = pi034 & ~pi037;
assign w532 = w526 & w531;
assign v161 = ~(pi109 | w241);
assign w533 = v161;
assign v162 = ~(w438 | w533);
assign w534 = v162;
assign w535 = pi058 & ~pi113;
assign w536 = ~pi120 & w535;
assign w537 = pi112 & ~pi124;
assign v163 = ~(w368 | w537);
assign w538 = v163;
assign w539 = pi047 & ~pi056;
assign w540 = pi062 & ~pi101;
assign w541 = w539 & w540;
assign w542 = ~w83 & w78;
assign w543 = pi001 & ~pi035;
assign w544 = pi001 & pi035;
assign w545 = pi037 & pi034;
assign w546 = pi062 & pi101;
assign v164 = ~(pi056 | pi047);
assign w547 = v164;
assign w548 = w8 & w78;
assign w549 = ~w543 & pi002;
assign w550 = w543 & pi045;
assign w551 = ~w543 & pi003;
assign w552 = w543 & pi040;
assign w553 = ~w96 & pi004;
assign w554 = w96 & pi041;
assign w555 = ~w96 & pi005;
assign w556 = w96 & pi039;
assign w557 = ~w96 & pi006;
assign w558 = w96 & pi042;
assign w559 = ~w96 & pi007;
assign w560 = w96 & pi043;
assign w561 = ~w96 & pi008;
assign w562 = w96 & pi044;
assign w563 = ~w96 & pi009;
assign w564 = w96 & pi046;
assign w565 = ~w96 & pi010;
assign w566 = w96 & pi045;
assign w567 = ~w96 & pi011;
assign w568 = w96 & pi040;
assign w569 = ~w543 & pi012;
assign w570 = w543 & pi041;
assign w571 = ~w543 & pi013;
assign w572 = w543 & pi039;
assign w573 = ~w543 & pi014;
assign w574 = w543 & pi042;
assign w575 = ~w543 & pi015;
assign w576 = w543 & pi043;
assign w577 = ~w543 & pi016;
assign w578 = w543 & pi044;
assign w579 = ~w543 & pi017;
assign w580 = w543 & pi046;
assign w581 = ~w544 & pi018;
assign w582 = w544 & pi041;
assign w583 = ~w544 & pi019;
assign w584 = w544 & pi039;
assign w585 = ~w544 & pi020;
assign w586 = w544 & pi042;
assign w587 = ~w544 & pi021;
assign w588 = w544 & pi043;
assign w589 = ~w544 & pi022;
assign w590 = w544 & pi044;
assign w591 = ~w544 & pi023;
assign w592 = w544 & pi046;
assign w593 = ~w544 & pi024;
assign w594 = w544 & pi045;
assign w595 = ~w544 & pi025;
assign w596 = w544 & pi040;
assign w597 = ~w163 & pi026;
assign w598 = w163 & pi041;
assign w599 = ~w163 & pi027;
assign w600 = w163 & pi039;
assign w601 = ~w163 & pi028;
assign w602 = w163 & pi042;
assign w603 = ~w163 & pi029;
assign w604 = w163 & pi043;
assign w605 = ~w163 & pi030;
assign w606 = w163 & pi044;
assign w607 = ~w163 & pi031;
assign w608 = w163 & pi046;
assign w609 = ~w163 & pi032;
assign w610 = w163 & pi045;
assign w611 = ~w163 & pi033;
assign w612 = w163 & pi040;
assign v165 = ~(pi038 | pi036);
assign w613 = v165;
assign w614 = pi056 & pi047;
assign w615 = ~w241 & pi047;
assign v166 = ~(w241 | w547);
assign w616 = v166;
assign w617 = w1 & w248;
assign w618 = ~w0 & w363;
assign v167 = ~(pi037 | pi034);
assign w619 = v167;
assign w620 = pi038 & pi036;
assign one = 1;
assign po000 = pi076;// level 0
assign po001 = pi061;// level 0
assign po002 = w7;// level 5
assign po003 = w15;// level 4
assign po004 = ~w26;// level 4
assign po005 = ~w33;// level 4
assign po006 = ~w40;// level 4
assign po007 = ~w47;// level 4
assign po008 = ~w54;// level 4
assign po009 = ~w61;// level 4
assign po010 = ~w68;// level 4
assign po011 = ~w75;// level 4
assign po012 = one;// level 0
assign po013 = pi117;// level 0
assign po014 = w82;// level 6
assign po015 = pi118;// level 0
assign po016 = w88;// level 6
assign po017 = ~w92;// level 6
assign po018 = ~w95;// level 6
assign po019 = ~w99;// level 6
assign po020 = ~w102;// level 6
assign po021 = ~w105;// level 6
assign po022 = ~w108;// level 6
assign po023 = ~w111;// level 6
assign po024 = ~w114;// level 6
assign po025 = ~w117;// level 6
assign po026 = ~w120;// level 6
assign po027 = ~w123;// level 6
assign po028 = ~w126;// level 6
assign po029 = ~w129;// level 6
assign po030 = ~w132;// level 6
assign po031 = ~w135;// level 6
assign po032 = ~w138;// level 6
assign po033 = ~w141;// level 6
assign po034 = ~w144;// level 6
assign po035 = ~w147;// level 6
assign po036 = ~w150;// level 6
assign po037 = ~w153;// level 6
assign po038 = ~w156;// level 6
assign po039 = ~w159;// level 6
assign po040 = ~w162;// level 6
assign po041 = ~w166;// level 6
assign po042 = ~w169;// level 6
assign po043 = ~w172;// level 6
assign po044 = ~w175;// level 6
assign po045 = ~w178;// level 6
assign po046 = ~w181;// level 6
assign po047 = ~w184;// level 6
assign po048 = ~w187;// level 6
assign po049 = ~w196;// level 5
assign po050 = ~w198;// level 6
assign po051 = ~w204;// level 6
assign po052 = w208;// level 4
assign po053 = w211;// level 5
assign po054 = ~w214;// level 3
assign po055 = ~w217;// level 3
assign po056 = ~w220;// level 3
assign po057 = ~w223;// level 3
assign po058 = ~w226;// level 3
assign po059 = ~w229;// level 3
assign po060 = ~w232;// level 3
assign po061 = ~w235;// level 3
assign po062 = ~w244;// level 5
assign po063 = ~w251;// level 5
assign po064 = ~w268;// level 6
assign po065 = ~w281;// level 6
assign po066 = ~w294;// level 6
assign po067 = ~w307;// level 6
assign po068 = ~w320;// level 6
assign po069 = ~w333;// level 6
assign po070 = ~w346;// level 6
assign po071 = w349;// level 5
assign po072 = ~w362;// level 6
assign po073 = ~w367;// level 5
assign po074 = ~w372;// level 4
assign po075 = w379;// level 4
assign po076 = w84;// level 4
assign po077 = ~w383;// level 5
assign po078 = ~w389;// level 4
assign po079 = ~w393;// level 4
assign po080 = ~w397;// level 4
assign po081 = ~w401;// level 4
assign po082 = ~w405;// level 4
assign po083 = ~w409;// level 4
assign po084 = ~w413;// level 4
assign po085 = ~w416;// level 4
assign po086 = ~w419;// level 4
assign po087 = ~w422;// level 4
assign po088 = ~w425;// level 4
assign po089 = ~w428;// level 4
assign po090 = ~w431;// level 4
assign po091 = ~w437;// level 4
assign po092 = w441;// level 4
assign po093 = w445;// level 4
assign po094 = ~w449;// level 4
assign po095 = ~w452;// level 4
assign po096 = ~w457;// level 4
assign po097 = ~w460;// level 4
assign po098 = pi106;// level 0
assign po099 = ~w463;// level 4
assign po100 = w468;// level 4
assign po101 = ~w472;// level 4
assign po102 = ~w475;// level 4
assign po103 = ~w478;// level 4
assign po104 = ~w481;// level 4
assign po105 = ~w484;// level 4
assign po106 = ~w487;// level 4
assign po107 = ~w490;// level 4
assign po108 = ~w493;// level 4
assign po109 = ~w496;// level 4
assign po110 = ~w499;// level 4
assign po111 = ~w503;// level 3
assign po112 = ~w504;// level 4
assign po113 = ~w507;// level 4
assign po114 = ~w510;// level 4
assign po115 = ~w513;// level 4
assign po116 = w516;// level 4
assign po117 = w517;// level 1
assign po118 = w520;// level 3
assign po119 = ~w522;// level 4
assign po120 = ~w525;// level 4
assign po121 = w528;// level 2
assign po122 = w530;// level 2
assign po123 = ~w532;// level 2
assign po124 = w534;// level 3
assign po125 = w536;// level 2
assign po126 = ~pi114;// level 0
assign po127 = ~w538;// level 2
assign po128 = ~w541;// level 2
assign po129 = w376;// level 1
assign po130 = pi116;// level 0
assign po131 = pi119;// level 0
endmodule
