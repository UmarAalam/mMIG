//Written by the Majority Logic Package Thu Apr 30 16:14:57 2015
module top (
            pi0000, pi0001, pi0002, pi0003, pi0004, pi0005, pi0006, pi0007, pi0008, pi0009, pi0010, pi0011, pi0012, pi0013, pi0014, pi0015, pi0016, pi0017, pi0018, pi0019, pi0020, pi0021, pi0022, pi0023, pi0024, pi0025, pi0026, pi0027, pi0028, pi0029, pi0030, pi0031, pi0032, pi0033, pi0034, pi0035, pi0036, pi0037, pi0038, pi0039, pi0040, pi0041, pi0042, pi0043, pi0044, pi0045, pi0046, pi0047, pi0048, pi0049, pi0050, pi0051, pi0052, pi0053, pi0054, pi0055, pi0056, pi0057, pi0058, pi0059, pi0060, pi0061, pi0062, pi0063, pi0064, pi0065, pi0066, pi0067, pi0068, pi0069, pi0070, pi0071, pi0072, pi0073, pi0074, pi0075, pi0076, pi0077, pi0078, pi0079, pi0080, pi0081, pi0082, pi0083, pi0084, pi0085, pi0086, pi0087, pi0088, pi0089, pi0090, pi0091, pi0092, pi0093, pi0094, pi0095, pi0096, pi0097, pi0098, pi0099, pi0100, pi0101, pi0102, pi0103, pi0104, pi0105, pi0106, pi0107, pi0108, pi0109, pi0110, pi0111, pi0112, pi0113, pi0114, pi0115, pi0116, pi0117, pi0118, pi0119, pi0120, pi0121, pi0122, pi0123, pi0124, pi0125, pi0126, pi0127, pi0128, pi0129, pi0130, pi0131, pi0132, pi0133, pi0134, pi0135, pi0136, pi0137, pi0138, pi0139, pi0140, pi0141, pi0142, pi0143, pi0144, pi0145, pi0146, pi0147, pi0148, pi0149, pi0150, pi0151, pi0152, pi0153, pi0154, pi0155, pi0156, pi0157, pi0158, pi0159, pi0160, pi0161, pi0162, pi0163, pi0164, pi0165, pi0166, pi0167, pi0168, pi0169, pi0170, pi0171, pi0172, pi0173, pi0174, pi0175, pi0176, pi0177, pi0178, pi0179, pi0180, pi0181, pi0182, pi0183, pi0184, pi0185, pi0186, pi0187, pi0188, pi0189, pi0190, pi0191, pi0192, pi0193, pi0194, pi0195, pi0196, pi0197, pi0198, pi0199, pi0200, pi0201, pi0202, pi0203, pi0204, pi0205, pi0206, pi0207, pi0208, pi0209, pi0210, pi0211, pi0212, pi0213, pi0214, pi0215, pi0216, pi0217, pi0218, pi0219, pi0220, pi0221, pi0222, pi0223, pi0224, pi0225, pi0226, pi0227, pi0228, pi0229, pi0230, pi0231, pi0232, pi0233, pi0234, pi0235, pi0236, pi0237, pi0238, pi0239, pi0240, pi0241, pi0242, pi0243, pi0244, pi0245, pi0246, pi0247, pi0248, pi0249, pi0250, pi0251, pi0252, pi0253, pi0254, pi0255, pi0256, pi0257, pi0258, pi0259, pi0260, pi0261, pi0262, pi0263, pi0264, pi0265, pi0266, pi0267, pi0268, pi0269, pi0270, pi0271, pi0272, pi0273, pi0274, pi0275, pi0276, pi0277, pi0278, pi0279, pi0280, pi0281, pi0282, pi0283, pi0284, pi0285, pi0286, pi0287, pi0288, pi0289, pi0290, pi0291, pi0292, pi0293, pi0294, pi0295, pi0296, pi0297, pi0298, pi0299, pi0300, pi0301, pi0302, pi0303, pi0304, pi0305, pi0306, pi0307, pi0308, pi0309, pi0310, pi0311, pi0312, pi0313, pi0314, pi0315, pi0316, pi0317, pi0318, pi0319, pi0320, pi0321, pi0322, pi0323, pi0324, pi0325, pi0326, pi0327, pi0328, pi0329, pi0330, pi0331, pi0332, pi0333, pi0334, pi0335, pi0336, pi0337, pi0338, pi0339, pi0340, pi0341, pi0342, pi0343, pi0344, pi0345, pi0346, pi0347, pi0348, pi0349, pi0350, pi0351, pi0352, pi0353, pi0354, pi0355, pi0356, pi0357, pi0358, pi0359, pi0360, pi0361, pi0362, pi0363, pi0364, pi0365, pi0366, pi0367, pi0368, pi0369, pi0370, pi0371, pi0372, pi0373, pi0374, pi0375, pi0376, pi0377, pi0378, pi0379, pi0380, pi0381, pi0382, pi0383, pi0384, pi0385, pi0386, pi0387, pi0388, pi0389, pi0390, pi0391, pi0392, pi0393, pi0394, pi0395, pi0396, pi0397, pi0398, pi0399, pi0400, pi0401, pi0402, pi0403, pi0404, pi0405, pi0406, pi0407, pi0408, pi0409, pi0410, pi0411, pi0412, pi0413, pi0414, pi0415, pi0416, pi0417, pi0418, pi0419, pi0420, pi0421, pi0422, pi0423, pi0424, pi0425, pi0426, pi0427, pi0428, pi0429, pi0430, pi0431, pi0432, pi0433, pi0434, pi0435, pi0436, pi0437, pi0438, pi0439, pi0440, pi0441, pi0442, pi0443, pi0444, pi0445, pi0446, pi0447, pi0448, pi0449, pi0450, pi0451, pi0452, pi0453, pi0454, pi0455, pi0456, pi0457, pi0458, pi0459, pi0460, pi0461, pi0462, pi0463, pi0464, pi0465, pi0466, pi0467, pi0468, pi0469, pi0470, pi0471, pi0472, pi0473, pi0474, pi0475, pi0476, pi0477, pi0478, pi0479, pi0480, pi0481, pi0482, pi0483, pi0484, pi0485, pi0486, pi0487, pi0488, pi0489, pi0490, pi0491, pi0492, pi0493, pi0494, pi0495, pi0496, pi0497, pi0498, pi0499, pi0500, pi0501, pi0502, pi0503, pi0504, pi0505, pi0506, pi0507, pi0508, pi0509, pi0510, pi0511, pi0512, pi0513, pi0514, pi0515, pi0516, pi0517, pi0518, pi0519, pi0520, pi0521, pi0522, pi0523, pi0524, pi0525, pi0526, pi0527, pi0528, pi0529, pi0530, pi0531, pi0532, pi0533, pi0534, pi0535, pi0536, pi0537, pi0538, pi0539, pi0540, pi0541, pi0542, pi0543, pi0544, pi0545, pi0546, pi0547, pi0548, pi0549, pi0550, pi0551, pi0552, pi0553, pi0554, pi0555, pi0556, pi0557, pi0558, pi0559, pi0560, pi0561, pi0562, pi0563, pi0564, pi0565, pi0566, pi0567, pi0568, pi0569, pi0570, pi0571, pi0572, pi0573, pi0574, pi0575, pi0576, pi0577, pi0578, pi0579, pi0580, pi0581, pi0582, pi0583, pi0584, pi0585, pi0586, pi0587, pi0588, pi0589, pi0590, pi0591, pi0592, pi0593, pi0594, pi0595, pi0596, pi0597, pi0598, pi0599, pi0600, pi0601, pi0602, pi0603, pi0604, pi0605, pi0606, pi0607, pi0608, pi0609, pi0610, pi0611, pi0612, pi0613, pi0614, pi0615, pi0616, pi0617, pi0618, pi0619, pi0620, pi0621, pi0622, pi0623, pi0624, pi0625, pi0626, pi0627, pi0628, pi0629, pi0630, pi0631, pi0632, pi0633, pi0634, pi0635, pi0636, pi0637, pi0638, pi0639, pi0640, pi0641, pi0642, pi0643, pi0644, pi0645, pi0646, pi0647, pi0648, pi0649, pi0650, pi0651, pi0652, pi0653, pi0654, pi0655, pi0656, pi0657, pi0658, pi0659, pi0660, pi0661, pi0662, pi0663, pi0664, pi0665, pi0666, pi0667, pi0668, pi0669, pi0670, pi0671, pi0672, pi0673, pi0674, pi0675, pi0676, pi0677, pi0678, pi0679, pi0680, pi0681, pi0682, pi0683, pi0684, pi0685, pi0686, pi0687, pi0688, pi0689, pi0690, pi0691, pi0692, pi0693, pi0694, pi0695, pi0696, pi0697, pi0698, pi0699, pi0700, pi0701, pi0702, pi0703, pi0704, pi0705, pi0706, pi0707, pi0708, pi0709, pi0710, pi0711, pi0712, pi0713, pi0714, pi0715, pi0716, pi0717, pi0718, pi0719, pi0720, pi0721, pi0722, pi0723, pi0724, pi0725, pi0726, pi0727, pi0728, pi0729, pi0730, pi0731, pi0732, pi0733, pi0734, pi0735, pi0736, pi0737, pi0738, pi0739, pi0740, pi0741, pi0742, pi0743, pi0744, pi0745, pi0746, pi0747, pi0748, pi0749, pi0750, pi0751, pi0752, pi0753, pi0754, pi0755, pi0756, pi0757, pi0758, pi0759, pi0760, pi0761, pi0762, pi0763, pi0764, pi0765, pi0766, pi0767, pi0768, pi0769, pi0770, pi0771, pi0772, pi0773, pi0774, pi0775, pi0776, pi0777, pi0778, pi0779, pi0780, pi0781, pi0782, pi0783, pi0784, pi0785, pi0786, pi0787, pi0788, pi0789, pi0790, pi0791, pi0792, pi0793, pi0794, pi0795, pi0796, pi0797, pi0798, pi0799, pi0800, pi0801, pi0802, pi0803, pi0804, pi0805, pi0806, pi0807, pi0808, pi0809, pi0810, pi0811, pi0812, pi0813, pi0814, pi0815, pi0816, pi0817, pi0818, pi0819, pi0820, pi0821, pi0822, pi0823, pi0824, pi0825, pi0826, pi0827, pi0828, pi0829, pi0830, pi0831, pi0832, pi0833, pi0834, pi0835, pi0836, pi0837, pi0838, pi0839, pi0840, pi0841, pi0842, pi0843, pi0844, pi0845, pi0846, pi0847, pi0848, pi0849, pi0850, pi0851, pi0852, pi0853, pi0854, pi0855, pi0856, pi0857, pi0858, pi0859, pi0860, pi0861, pi0862, pi0863, pi0864, pi0865, pi0866, pi0867, pi0868, pi0869, pi0870, pi0871, pi0872, pi0873, pi0874, pi0875, pi0876, pi0877, pi0878, pi0879, pi0880, pi0881, pi0882, pi0883, pi0884, pi0885, pi0886, pi0887, pi0888, pi0889, pi0890, pi0891, pi0892, pi0893, pi0894, pi0895, pi0896, pi0897, pi0898, pi0899, pi0900, pi0901, pi0902, pi0903, pi0904, pi0905, pi0906, pi0907, pi0908, pi0909, pi0910, pi0911, pi0912, pi0913, pi0914, pi0915, pi0916, pi0917, pi0918, pi0919, pi0920, pi0921, pi0922, pi0923, pi0924, pi0925, pi0926, pi0927, pi0928, pi0929, pi0930, pi0931, pi0932, pi0933, pi0934, pi0935, pi0936, pi0937, pi0938, pi0939, pi0940, pi0941, pi0942, pi0943, pi0944, pi0945, pi0946, pi0947, pi0948, pi0949, pi0950, pi0951, pi0952, pi0953, pi0954, pi0955, pi0956, pi0957, pi0958, pi0959, pi0960, pi0961, pi0962, pi0963, pi0964, pi0965, pi0966, pi0967, pi0968, pi0969, pi0970, pi0971, pi0972, pi0973, pi0974, pi0975, pi0976, pi0977, pi0978, pi0979, pi0980, pi0981, pi0982, pi0983, pi0984, pi0985, pi0986, pi0987, pi0988, pi0989, pi0990, pi0991, pi0992, pi0993, pi0994, pi0995, pi0996, pi0997, pi0998, pi0999, pi1000, pi1001, pi1002, pi1003, pi1004, pi1005, pi1006, pi1007, pi1008, pi1009, pi1010, pi1011, pi1012, pi1013, pi1014, pi1015, pi1016, pi1017, pi1018, pi1019, pi1020, pi1021, pi1022, pi1023, pi1024, pi1025, pi1026, pi1027, pi1028, pi1029, pi1030, pi1031, pi1032, pi1033, pi1034, pi1035, pi1036, pi1037, pi1038, pi1039, pi1040, pi1041, pi1042, pi1043, pi1044, pi1045, pi1046, pi1047, pi1048, pi1049, pi1050, pi1051, pi1052, pi1053, pi1054, pi1055, pi1056, pi1057, pi1058, pi1059, pi1060, pi1061, pi1062, pi1063, pi1064, pi1065, pi1066, pi1067, pi1068, pi1069, pi1070, pi1071, pi1072, pi1073, pi1074, pi1075, pi1076, pi1077, pi1078, pi1079, pi1080, pi1081, pi1082, pi1083, pi1084, pi1085, pi1086, pi1087, pi1088, pi1089, pi1090, pi1091, pi1092, pi1093, pi1094, pi1095, pi1096, pi1097, pi1098, pi1099, pi1100, pi1101, pi1102, pi1103, pi1104, pi1105, pi1106, pi1107, pi1108, pi1109, pi1110, pi1111, pi1112, pi1113, pi1114, pi1115, pi1116, pi1117, pi1118, pi1119, pi1120, pi1121, pi1122, pi1123, pi1124, pi1125, pi1126, pi1127, pi1128, pi1129, pi1130, pi1131, pi1132, pi1133, pi1134, pi1135, pi1136, pi1137, pi1138, pi1139, pi1140, pi1141, pi1142, pi1143, pi1144, pi1145, pi1146, pi1147, pi1148, pi1149, pi1150, pi1151, pi1152, pi1153, pi1154, pi1155, pi1156, pi1157, pi1158, pi1159, pi1160, pi1161, pi1162, pi1163, pi1164, pi1165, pi1166, pi1167, pi1168, pi1169, pi1170, pi1171, pi1172, pi1173, pi1174, pi1175, pi1176, pi1177, pi1178, pi1179, pi1180, pi1181, pi1182, pi1183, pi1184, pi1185, pi1186, pi1187, pi1188, pi1189, pi1190, pi1191, pi1192, pi1193, pi1194, pi1195, pi1196, pi1197, pi1198, pi1199, pi1200, pi1201, pi1202, pi1203, pi1204, pi1205, pi1206, pi1207, pi1208, pi1209, pi1210, pi1211, pi1212, pi1213, pi1214, pi1215, pi1216, pi1217, pi1218, pi1219, pi1220, pi1221, pi1222, pi1223, pi1224, pi1225, pi1226, pi1227, pi1228, pi1229, pi1230, pi1231, pi1232, pi1233, pi1234, pi1235, pi1236, pi1237, pi1238, pi1239, pi1240, pi1241, pi1242, pi1243, pi1244, pi1245, pi1246, pi1247, pi1248, pi1249, pi1250, pi1251, pi1252, pi1253, pi1254, pi1255, pi1256, pi1257, pi1258, pi1259, pi1260, pi1261, pi1262, pi1263, pi1264, pi1265, pi1266, pi1267, pi1268, pi1269, pi1270, pi1271, pi1272, pi1273, pi1274, pi1275, pi1276, pi1277, pi1278, pi1279, pi1280, pi1281, pi1282, pi1283, pi1284, pi1285, pi1286, pi1287, pi1288, pi1289, pi1290, pi1291, pi1292, pi1293, pi1294, pi1295, pi1296, pi1297, pi1298, pi1299, pi1300, pi1301, pi1302, pi1303, pi1304, pi1305, pi1306, pi1307, pi1308, pi1309, pi1310, pi1311, pi1312, pi1313, pi1314, pi1315, pi1316, pi1317, pi1318, pi1319, pi1320, pi1321, pi1322, pi1323, pi1324, pi1325, pi1326, pi1327, pi1328, pi1329, pi1330, pi1331, pi1332, pi1333, pi1334, pi1335, pi1336, pi1337, pi1338, pi1339, pi1340, pi1341, pi1342, pi1343, pi1344, pi1345, pi1346, pi1347, pi1348, pi1349, pi1350, pi1351, pi1352, pi1353, pi1354, pi1355, pi1356, pi1357, pi1358, pi1359, pi1360, pi1361, pi1362, pi1363, pi1364, pi1365, pi1366, pi1367, pi1368, pi1369, pi1370, pi1371, pi1372, pi1373, pi1374, pi1375, pi1376, pi1377, pi1378, pi1379, pi1380, pi1381, pi1382, pi1383, pi1384, pi1385, pi1386, pi1387, pi1388, pi1389, pi1390, pi1391, pi1392, pi1393, pi1394, pi1395, pi1396, pi1397, pi1398, pi1399, pi1400, pi1401, pi1402, pi1403, pi1404, pi1405, pi1406, pi1407, pi1408, pi1409, pi1410, pi1411, pi1412, pi1413, pi1414, pi1415, pi1416, pi1417, pi1418, pi1419, pi1420, pi1421, pi1422, pi1423, pi1424, pi1425, pi1426, pi1427, pi1428, pi1429, pi1430, pi1431, pi1432, pi1433, pi1434, pi1435, pi1436, pi1437, pi1438, pi1439, pi1440, pi1441, pi1442, pi1443, pi1444, pi1445, pi1446, pi1447, pi1448, pi1449, pi1450, pi1451, pi1452, pi1453, pi1454, pi1455, pi1456, pi1457, pi1458, pi1459, pi1460, pi1461, pi1462, pi1463, pi1464, pi1465, pi1466, pi1467, pi1468, pi1469, pi1470, pi1471, pi1472, pi1473, pi1474, pi1475, pi1476, pi1477, pi1478, pi1479, pi1480, pi1481, pi1482, pi1483, pi1484, pi1485, pi1486, pi1487, pi1488, pi1489, pi1490, pi1491, pi1492, pi1493, pi1494, pi1495, pi1496, pi1497, pi1498, pi1499, pi1500, pi1501, pi1502, pi1503, pi1504, pi1505, pi1506, pi1507, pi1508, pi1509, pi1510, pi1511, pi1512, pi1513, pi1514, pi1515, pi1516, pi1517, pi1518, pi1519, pi1520, pi1521, pi1522, pi1523, pi1524, pi1525, pi1526, pi1527, pi1528, pi1529, pi1530, pi1531, pi1532, pi1533, pi1534, pi1535, pi1536, pi1537, pi1538, pi1539, pi1540, pi1541, pi1542, pi1543, pi1544, pi1545, pi1546, pi1547, pi1548, pi1549, pi1550, pi1551, pi1552, pi1553, pi1554, pi1555, pi1556, pi1557, pi1558, pi1559, pi1560, pi1561, pi1562, pi1563, pi1564, pi1565, pi1566, pi1567, pi1568, pi1569, pi1570, pi1571, pi1572, pi1573, pi1574, pi1575, pi1576, pi1577, pi1578, pi1579, pi1580, pi1581, pi1582, pi1583, pi1584, pi1585, pi1586, pi1587, pi1588, pi1589, pi1590, pi1591, pi1592, pi1593, pi1594, pi1595, pi1596, pi1597, pi1598, pi1599, pi1600, pi1601, pi1602, pi1603, pi1604, pi1605, pi1606, pi1607, pi1608, pi1609, pi1610, pi1611, pi1612, pi1613, pi1614, pi1615, pi1616, pi1617, pi1618, pi1619, pi1620, pi1621, pi1622, pi1623, pi1624, pi1625, pi1626, pi1627, pi1628, pi1629, pi1630, pi1631, pi1632, pi1633, pi1634, pi1635, pi1636, pi1637, pi1638, pi1639, pi1640, pi1641, pi1642, pi1643, pi1644, pi1645, pi1646, pi1647, pi1648, pi1649, pi1650, pi1651, pi1652, pi1653, pi1654, pi1655, pi1656, pi1657, pi1658, pi1659, pi1660, pi1661, pi1662, pi1663, pi1664, pi1665, pi1666, pi1667, pi1668, pi1669, pi1670, pi1671, pi1672, pi1673, pi1674, pi1675, pi1676, pi1677, pi1678, pi1679, pi1680, pi1681, pi1682, pi1683, pi1684, pi1685, pi1686, pi1687, pi1688, pi1689, pi1690, pi1691, pi1692, pi1693, pi1694, pi1695, pi1696, pi1697, pi1698, pi1699, pi1700, pi1701, pi1702, pi1703, pi1704, pi1705, pi1706, pi1707, pi1708, pi1709, pi1710, pi1711, pi1712, pi1713, pi1714, pi1715, pi1716, pi1717, pi1718, pi1719, pi1720, pi1721, pi1722, pi1723, pi1724, pi1725, pi1726, pi1727, pi1728, pi1729, pi1730, pi1731, pi1732, pi1733, pi1734, pi1735, pi1736, pi1737, pi1738, pi1739, pi1740, pi1741, pi1742, pi1743, pi1744, pi1745, pi1746, pi1747, pi1748, pi1749, pi1750, pi1751, pi1752, pi1753, pi1754, pi1755, pi1756, pi1757, pi1758, pi1759, pi1760, pi1761, pi1762, pi1763, pi1764, pi1765, pi1766, pi1767, pi1768, pi1769, pi1770, pi1771, pi1772, pi1773, pi1774, pi1775, pi1776, pi1777, pi1778, pi1779, pi1780, pi1781, pi1782, pi1783, pi1784, pi1785, pi1786, pi1787, pi1788, pi1789, pi1790, pi1791, pi1792, pi1793, pi1794, pi1795, pi1796, pi1797, pi1798, pi1799, pi1800, pi1801, pi1802, pi1803, pi1804, pi1805, pi1806, pi1807, pi1808, pi1809, pi1810, pi1811, pi1812, pi1813, pi1814, pi1815, pi1816, pi1817, pi1818, pi1819, pi1820, pi1821, pi1822, pi1823, pi1824, pi1825, pi1826, pi1827, pi1828, pi1829, pi1830, pi1831, pi1832, pi1833, pi1834, pi1835, pi1836, pi1837, pi1838, pi1839, pi1840, pi1841, pi1842, pi1843, pi1844, pi1845, pi1846, pi1847, pi1848, pi1849, pi1850, pi1851, pi1852, pi1853, pi1854, pi1855, pi1856, pi1857, pi1858, pi1859, 
            po0000, po0001, po0002, po0003, po0004, po0005, po0006, po0007, po0008, po0009, po0010, po0011, po0012, po0013, po0014, po0015, po0016, po0017, po0018, po0019, po0020, po0021, po0022, po0023, po0024, po0025, po0026, po0027, po0028, po0029, po0030, po0031, po0032, po0033, po0034, po0035, po0036, po0037, po0038, po0039, po0040, po0041, po0042, po0043, po0044, po0045, po0046, po0047, po0048, po0049, po0050, po0051, po0052, po0053, po0054, po0055, po0056, po0057, po0058, po0059, po0060, po0061, po0062, po0063, po0064, po0065, po0066, po0067, po0068, po0069, po0070, po0071, po0072, po0073, po0074, po0075, po0076, po0077, po0078, po0079, po0080, po0081, po0082, po0083, po0084, po0085, po0086, po0087, po0088, po0089, po0090, po0091, po0092, po0093, po0094, po0095, po0096, po0097, po0098, po0099, po0100, po0101, po0102, po0103, po0104, po0105, po0106, po0107, po0108, po0109, po0110, po0111, po0112, po0113, po0114, po0115, po0116, po0117, po0118, po0119, po0120, po0121, po0122, po0123, po0124, po0125, po0126, po0127, po0128, po0129, po0130, po0131, po0132, po0133, po0134, po0135, po0136, po0137, po0138, po0139, po0140, po0141, po0142, po0143, po0144, po0145, po0146, po0147, po0148, po0149, po0150, po0151, po0152, po0153, po0154, po0155, po0156, po0157, po0158, po0159, po0160, po0161, po0162, po0163, po0164, po0165, po0166, po0167, po0168, po0169, po0170, po0171, po0172, po0173, po0174, po0175, po0176, po0177, po0178, po0179, po0180, po0181, po0182, po0183, po0184, po0185, po0186, po0187, po0188, po0189, po0190, po0191, po0192, po0193, po0194, po0195, po0196, po0197, po0198, po0199, po0200, po0201, po0202, po0203, po0204, po0205, po0206, po0207, po0208, po0209, po0210, po0211, po0212, po0213, po0214, po0215, po0216, po0217, po0218, po0219, po0220, po0221, po0222, po0223, po0224, po0225, po0226, po0227, po0228, po0229, po0230, po0231, po0232, po0233, po0234, po0235, po0236, po0237, po0238, po0239, po0240, po0241, po0242, po0243, po0244, po0245, po0246, po0247, po0248, po0249, po0250, po0251, po0252, po0253, po0254, po0255, po0256, po0257, po0258, po0259, po0260, po0261, po0262, po0263, po0264, po0265, po0266, po0267, po0268, po0269, po0270, po0271, po0272, po0273, po0274, po0275, po0276, po0277, po0278, po0279, po0280, po0281, po0282, po0283, po0284, po0285, po0286, po0287, po0288, po0289, po0290, po0291, po0292, po0293, po0294, po0295, po0296, po0297, po0298, po0299, po0300, po0301, po0302, po0303, po0304, po0305, po0306, po0307, po0308, po0309, po0310, po0311, po0312, po0313, po0314, po0315, po0316, po0317, po0318, po0319, po0320, po0321, po0322, po0323, po0324, po0325, po0326, po0327, po0328, po0329, po0330, po0331, po0332, po0333, po0334, po0335, po0336, po0337, po0338, po0339, po0340, po0341, po0342, po0343, po0344, po0345, po0346, po0347, po0348, po0349, po0350, po0351, po0352, po0353, po0354, po0355, po0356, po0357, po0358, po0359, po0360, po0361, po0362, po0363, po0364, po0365, po0366, po0367, po0368, po0369, po0370, po0371, po0372, po0373, po0374, po0375, po0376, po0377, po0378, po0379, po0380, po0381, po0382, po0383, po0384, po0385, po0386, po0387, po0388, po0389, po0390, po0391, po0392, po0393, po0394, po0395, po0396, po0397, po0398, po0399, po0400, po0401, po0402, po0403, po0404, po0405, po0406, po0407, po0408, po0409, po0410, po0411, po0412, po0413, po0414, po0415, po0416, po0417, po0418, po0419, po0420, po0421, po0422, po0423, po0424, po0425, po0426, po0427, po0428, po0429, po0430, po0431, po0432, po0433, po0434, po0435, po0436, po0437, po0438, po0439, po0440, po0441, po0442, po0443, po0444, po0445, po0446, po0447, po0448, po0449, po0450, po0451, po0452, po0453, po0454, po0455, po0456, po0457, po0458, po0459, po0460, po0461, po0462, po0463, po0464, po0465, po0466, po0467, po0468, po0469, po0470, po0471, po0472, po0473, po0474, po0475, po0476, po0477, po0478, po0479, po0480, po0481, po0482, po0483, po0484, po0485, po0486, po0487, po0488, po0489, po0490, po0491, po0492, po0493, po0494, po0495, po0496, po0497, po0498, po0499, po0500, po0501, po0502, po0503, po0504, po0505, po0506, po0507, po0508, po0509, po0510, po0511, po0512, po0513, po0514, po0515, po0516, po0517, po0518, po0519, po0520, po0521, po0522, po0523, po0524, po0525, po0526, po0527, po0528, po0529, po0530, po0531, po0532, po0533, po0534, po0535, po0536, po0537, po0538, po0539, po0540, po0541, po0542, po0543, po0544, po0545, po0546, po0547, po0548, po0549, po0550, po0551, po0552, po0553, po0554, po0555, po0556, po0557, po0558, po0559, po0560, po0561, po0562, po0563, po0564, po0565, po0566, po0567, po0568, po0569, po0570, po0571, po0572, po0573, po0574, po0575, po0576, po0577, po0578, po0579, po0580, po0581, po0582, po0583, po0584, po0585, po0586, po0587, po0588, po0589, po0590, po0591, po0592, po0593, po0594, po0595, po0596, po0597, po0598, po0599, po0600, po0601, po0602, po0603, po0604, po0605, po0606, po0607, po0608, po0609, po0610, po0611, po0612, po0613, po0614, po0615, po0616, po0617, po0618, po0619, po0620, po0621, po0622, po0623, po0624, po0625, po0626, po0627, po0628, po0629, po0630, po0631, po0632, po0633, po0634, po0635, po0636, po0637, po0638, po0639, po0640, po0641, po0642, po0643, po0644, po0645, po0646, po0647, po0648, po0649, po0650, po0651, po0652, po0653, po0654, po0655, po0656, po0657, po0658, po0659, po0660, po0661, po0662, po0663, po0664, po0665, po0666, po0667, po0668, po0669, po0670, po0671, po0672, po0673, po0674, po0675, po0676, po0677, po0678, po0679, po0680, po0681, po0682, po0683, po0684, po0685, po0686, po0687, po0688, po0689, po0690, po0691, po0692, po0693, po0694, po0695, po0696, po0697, po0698, po0699, po0700, po0701, po0702, po0703, po0704, po0705, po0706, po0707, po0708, po0709, po0710, po0711, po0712, po0713, po0714, po0715, po0716, po0717, po0718, po0719, po0720, po0721, po0722, po0723, po0724, po0725, po0726, po0727, po0728, po0729, po0730, po0731, po0732, po0733, po0734, po0735, po0736, po0737, po0738, po0739, po0740, po0741, po0742, po0743, po0744, po0745, po0746, po0747, po0748, po0749, po0750, po0751, po0752, po0753, po0754, po0755, po0756, po0757, po0758, po0759, po0760, po0761, po0762, po0763, po0764, po0765, po0766, po0767, po0768, po0769, po0770, po0771, po0772, po0773, po0774, po0775, po0776, po0777, po0778, po0779, po0780, po0781, po0782, po0783, po0784, po0785, po0786, po0787, po0788, po0789, po0790, po0791, po0792, po0793, po0794, po0795, po0796, po0797, po0798, po0799, po0800, po0801, po0802, po0803, po0804, po0805, po0806, po0807, po0808, po0809, po0810, po0811, po0812, po0813, po0814, po0815, po0816, po0817, po0818, po0819, po0820, po0821, po0822, po0823, po0824, po0825, po0826, po0827, po0828, po0829, po0830, po0831, po0832, po0833, po0834, po0835, po0836, po0837, po0838, po0839, po0840, po0841, po0842, po0843, po0844, po0845, po0846, po0847, po0848, po0849, po0850, po0851, po0852, po0853, po0854, po0855, po0856, po0857, po0858, po0859, po0860, po0861, po0862, po0863, po0864, po0865, po0866, po0867, po0868, po0869, po0870, po0871, po0872, po0873, po0874, po0875, po0876, po0877, po0878, po0879, po0880, po0881, po0882, po0883, po0884, po0885, po0886, po0887, po0888, po0889, po0890, po0891, po0892, po0893, po0894, po0895, po0896, po0897, po0898, po0899, po0900, po0901, po0902, po0903, po0904, po0905, po0906, po0907, po0908, po0909, po0910, po0911, po0912, po0913, po0914, po0915, po0916, po0917, po0918, po0919, po0920, po0921, po0922, po0923, po0924, po0925, po0926, po0927, po0928, po0929, po0930, po0931, po0932, po0933, po0934, po0935, po0936, po0937, po0938, po0939, po0940, po0941, po0942, po0943, po0944, po0945, po0946, po0947, po0948, po0949, po0950, po0951, po0952, po0953, po0954, po0955, po0956, po0957, po0958, po0959, po0960, po0961, po0962, po0963, po0964, po0965, po0966, po0967, po0968, po0969, po0970, po0971, po0972, po0973, po0974, po0975, po0976, po0977, po0978, po0979, po0980, po0981, po0982, po0983, po0984, po0985, po0986, po0987, po0988, po0989, po0990, po0991, po0992, po0993, po0994, po0995, po0996, po0997, po0998, po0999, po1000, po1001, po1002, po1003, po1004, po1005, po1006, po1007, po1008, po1009, po1010, po1011, po1012, po1013, po1014, po1015, po1016, po1017, po1018, po1019, po1020, po1021, po1022, po1023, po1024, po1025, po1026, po1027, po1028, po1029, po1030, po1031, po1032, po1033, po1034, po1035, po1036, po1037, po1038, po1039, po1040, po1041, po1042, po1043, po1044, po1045, po1046, po1047, po1048, po1049, po1050, po1051, po1052, po1053, po1054, po1055, po1056, po1057, po1058, po1059, po1060, po1061, po1062, po1063, po1064, po1065, po1066, po1067, po1068, po1069, po1070, po1071, po1072, po1073, po1074, po1075, po1076, po1077, po1078, po1079, po1080, po1081, po1082, po1083, po1084, po1085, po1086, po1087, po1088, po1089, po1090, po1091, po1092, po1093, po1094, po1095, po1096, po1097, po1098, po1099, po1100, po1101, po1102, po1103, po1104, po1105, po1106, po1107, po1108, po1109, po1110, po1111, po1112, po1113, po1114, po1115, po1116, po1117, po1118, po1119, po1120, po1121, po1122, po1123, po1124, po1125, po1126, po1127, po1128, po1129, po1130, po1131, po1132, po1133, po1134, po1135, po1136, po1137, po1138, po1139, po1140, po1141, po1142, po1143, po1144, po1145, po1146, po1147, po1148, po1149, po1150, po1151, po1152, po1153, po1154, po1155, po1156, po1157, po1158, po1159, po1160, po1161, po1162, po1163, po1164, po1165, po1166, po1167, po1168, po1169, po1170, po1171, po1172, po1173, po1174, po1175, po1176, po1177, po1178, po1179, po1180, po1181, po1182, po1183, po1184, po1185, po1186, po1187, po1188, po1189, po1190, po1191, po1192, po1193, po1194, po1195, po1196, po1197, po1198, po1199, po1200, po1201, po1202, po1203, po1204, po1205, po1206, po1207, po1208, po1209, po1210, po1211, po1212, po1213, po1214, po1215, po1216, po1217, po1218, po1219, po1220, po1221, po1222, po1223, po1224, po1225, po1226, po1227, po1228, po1229, po1230, po1231, po1232, po1233, po1234, po1235, po1236, po1237, po1238, po1239, po1240, po1241, po1242, po1243, po1244, po1245, po1246, po1247, po1248, po1249, po1250, po1251, po1252, po1253, po1254, po1255, po1256, po1257, po1258, po1259, po1260, po1261, po1262, po1263, po1264, po1265, po1266, po1267, po1268, po1269, po1270, po1271, po1272, po1273, po1274, po1275, po1276, po1277, po1278, po1279, po1280, po1281, po1282, po1283, po1284, po1285, po1286, po1287, po1288, po1289, po1290, po1291, po1292, po1293, po1294, po1295, po1296, po1297, po1298, po1299, po1300, po1301, po1302, po1303, po1304, po1305, po1306, po1307, po1308, po1309, po1310, po1311, po1312, po1313, po1314, po1315, po1316, po1317, po1318, po1319, po1320, po1321, po1322, po1323, po1324, po1325, po1326, po1327, po1328, po1329, po1330, po1331, po1332, po1333, po1334, po1335, po1336, po1337, po1338, po1339, po1340, po1341, po1342, po1343, po1344, po1345, po1346, po1347, po1348, po1349, po1350, po1351, po1352, po1353, po1354, po1355, po1356, po1357, po1358, po1359, po1360, po1361, po1362, po1363, po1364, po1365, po1366, po1367, po1368, po1369, po1370, po1371, po1372, po1373, po1374, po1375, po1376, po1377, po1378, po1379, po1380, po1381, po1382, po1383, po1384, po1385, po1386, po1387, po1388, po1389, po1390, po1391, po1392, po1393, po1394, po1395, po1396, po1397, po1398, po1399, po1400, po1401, po1402, po1403, po1404, po1405, po1406, po1407, po1408, po1409, po1410, po1411, po1412, po1413, po1414, po1415, po1416, po1417, po1418, po1419, po1420, po1421, po1422, po1423, po1424, po1425, po1426, po1427, po1428, po1429, po1430, po1431, po1432, po1433, po1434, po1435, po1436, po1437, po1438, po1439, po1440, po1441, po1442, po1443, po1444, po1445, po1446, po1447, po1448, po1449, po1450, po1451, po1452, po1453, po1454, po1455, po1456, po1457, po1458, po1459, po1460, po1461, po1462, po1463, po1464, po1465, po1466, po1467, po1468, po1469, po1470, po1471, po1472, po1473, po1474, po1475, po1476, po1477, po1478, po1479, po1480, po1481, po1482, po1483, po1484, po1485, po1486, po1487, po1488, po1489, po1490, po1491, po1492, po1493, po1494, po1495, po1496, po1497, po1498, po1499, po1500, po1501, po1502, po1503, po1504, po1505, po1506, po1507, po1508, po1509, po1510, po1511, po1512, po1513, po1514, po1515, po1516, po1517, po1518, po1519, po1520, po1521, po1522, po1523, po1524, po1525, po1526, po1527, po1528, po1529, po1530, po1531, po1532, po1533, po1534, po1535, po1536, po1537, po1538, po1539, po1540, po1541, po1542, po1543, po1544, po1545, po1546, po1547, po1548, po1549, po1550, po1551, po1552, po1553, po1554, po1555, po1556, po1557, po1558, po1559, po1560, po1561, po1562, po1563, po1564, po1565, po1566, po1567, po1568, po1569, po1570, po1571, po1572, po1573, po1574, po1575, po1576, po1577, po1578, po1579, po1580, po1581, po1582, po1583, po1584, po1585, po1586, po1587, po1588, po1589, po1590, po1591, po1592, po1593, po1594, po1595, po1596, po1597, po1598, po1599, po1600, po1601, po1602, po1603, po1604, po1605, po1606, po1607, po1608, po1609, po1610, po1611, po1612, po1613, po1614, po1615, po1616, po1617, po1618, po1619, po1620, po1621, po1622, po1623, po1624, po1625, po1626, po1627, po1628, po1629, po1630, po1631, po1632, po1633, po1634, po1635, po1636, po1637, po1638, po1639, po1640, po1641, po1642, po1643, po1644, po1645, po1646, po1647, po1648, po1649, po1650, po1651, po1652, po1653, po1654, po1655, po1656, po1657, po1658, po1659, po1660, po1661, po1662, po1663, po1664, po1665, po1666, po1667, po1668, po1669, po1670, po1671, po1672, po1673, po1674, po1675, po1676, po1677, po1678, po1679, po1680, po1681, po1682, po1683, po1684, po1685, po1686, po1687, po1688, po1689, po1690, po1691, po1692, po1693, po1694, po1695, po1696, po1697, po1698, po1699, po1700, po1701, po1702, po1703, po1704, po1705, po1706, po1707, po1708, po1709, po1710, po1711, po1712, po1713, po1714, po1715, po1716, po1717, po1718, po1719, po1720, po1721, po1722, po1723, po1724, po1725, po1726, po1727, po1728, po1729, po1730, po1731, po1732, po1733, po1734, po1735, po1736, po1737, po1738, po1739, po1740, po1741, po1742, po1743, po1744, po1745, po1746, po1747, po1748, po1749, po1750, po1751, po1752, po1753, po1754, po1755, po1756, po1757, po1758, po1759, po1760, po1761, po1762, po1763, po1764, po1765, po1766, po1767, po1768, po1769, po1770, po1771, po1772, po1773, po1774, po1775, po1776, po1777, po1778, po1779, po1780, po1781, po1782, po1783, po1784, po1785, po1786, po1787, po1788, po1789, po1790, po1791, po1792, po1793, po1794, po1795, po1796, po1797, po1798, po1799, po1800, po1801, po1802, po1803, po1804, po1805, po1806, po1807, po1808, po1809, po1810, po1811, po1812, po1813, po1814, po1815, po1816, po1817, po1818, po1819, po1820, po1821, po1822, po1823, po1824, po1825, po1826, po1827, po1828, po1829, po1830, po1831, po1832, po1833, po1834, po1835, po1836, po1837, po1838, po1839, po1840, po1841, po1842, po1843, po1844, po1845);
input pi0000, pi0001, pi0002, pi0003, pi0004, pi0005, pi0006, pi0007, pi0008, pi0009, pi0010, pi0011, pi0012, pi0013, pi0014, pi0015, pi0016, pi0017, pi0018, pi0019, pi0020, pi0021, pi0022, pi0023, pi0024, pi0025, pi0026, pi0027, pi0028, pi0029, pi0030, pi0031, pi0032, pi0033, pi0034, pi0035, pi0036, pi0037, pi0038, pi0039, pi0040, pi0041, pi0042, pi0043, pi0044, pi0045, pi0046, pi0047, pi0048, pi0049, pi0050, pi0051, pi0052, pi0053, pi0054, pi0055, pi0056, pi0057, pi0058, pi0059, pi0060, pi0061, pi0062, pi0063, pi0064, pi0065, pi0066, pi0067, pi0068, pi0069, pi0070, pi0071, pi0072, pi0073, pi0074, pi0075, pi0076, pi0077, pi0078, pi0079, pi0080, pi0081, pi0082, pi0083, pi0084, pi0085, pi0086, pi0087, pi0088, pi0089, pi0090, pi0091, pi0092, pi0093, pi0094, pi0095, pi0096, pi0097, pi0098, pi0099, pi0100, pi0101, pi0102, pi0103, pi0104, pi0105, pi0106, pi0107, pi0108, pi0109, pi0110, pi0111, pi0112, pi0113, pi0114, pi0115, pi0116, pi0117, pi0118, pi0119, pi0120, pi0121, pi0122, pi0123, pi0124, pi0125, pi0126, pi0127, pi0128, pi0129, pi0130, pi0131, pi0132, pi0133, pi0134, pi0135, pi0136, pi0137, pi0138, pi0139, pi0140, pi0141, pi0142, pi0143, pi0144, pi0145, pi0146, pi0147, pi0148, pi0149, pi0150, pi0151, pi0152, pi0153, pi0154, pi0155, pi0156, pi0157, pi0158, pi0159, pi0160, pi0161, pi0162, pi0163, pi0164, pi0165, pi0166, pi0167, pi0168, pi0169, pi0170, pi0171, pi0172, pi0173, pi0174, pi0175, pi0176, pi0177, pi0178, pi0179, pi0180, pi0181, pi0182, pi0183, pi0184, pi0185, pi0186, pi0187, pi0188, pi0189, pi0190, pi0191, pi0192, pi0193, pi0194, pi0195, pi0196, pi0197, pi0198, pi0199, pi0200, pi0201, pi0202, pi0203, pi0204, pi0205, pi0206, pi0207, pi0208, pi0209, pi0210, pi0211, pi0212, pi0213, pi0214, pi0215, pi0216, pi0217, pi0218, pi0219, pi0220, pi0221, pi0222, pi0223, pi0224, pi0225, pi0226, pi0227, pi0228, pi0229, pi0230, pi0231, pi0232, pi0233, pi0234, pi0235, pi0236, pi0237, pi0238, pi0239, pi0240, pi0241, pi0242, pi0243, pi0244, pi0245, pi0246, pi0247, pi0248, pi0249, pi0250, pi0251, pi0252, pi0253, pi0254, pi0255, pi0256, pi0257, pi0258, pi0259, pi0260, pi0261, pi0262, pi0263, pi0264, pi0265, pi0266, pi0267, pi0268, pi0269, pi0270, pi0271, pi0272, pi0273, pi0274, pi0275, pi0276, pi0277, pi0278, pi0279, pi0280, pi0281, pi0282, pi0283, pi0284, pi0285, pi0286, pi0287, pi0288, pi0289, pi0290, pi0291, pi0292, pi0293, pi0294, pi0295, pi0296, pi0297, pi0298, pi0299, pi0300, pi0301, pi0302, pi0303, pi0304, pi0305, pi0306, pi0307, pi0308, pi0309, pi0310, pi0311, pi0312, pi0313, pi0314, pi0315, pi0316, pi0317, pi0318, pi0319, pi0320, pi0321, pi0322, pi0323, pi0324, pi0325, pi0326, pi0327, pi0328, pi0329, pi0330, pi0331, pi0332, pi0333, pi0334, pi0335, pi0336, pi0337, pi0338, pi0339, pi0340, pi0341, pi0342, pi0343, pi0344, pi0345, pi0346, pi0347, pi0348, pi0349, pi0350, pi0351, pi0352, pi0353, pi0354, pi0355, pi0356, pi0357, pi0358, pi0359, pi0360, pi0361, pi0362, pi0363, pi0364, pi0365, pi0366, pi0367, pi0368, pi0369, pi0370, pi0371, pi0372, pi0373, pi0374, pi0375, pi0376, pi0377, pi0378, pi0379, pi0380, pi0381, pi0382, pi0383, pi0384, pi0385, pi0386, pi0387, pi0388, pi0389, pi0390, pi0391, pi0392, pi0393, pi0394, pi0395, pi0396, pi0397, pi0398, pi0399, pi0400, pi0401, pi0402, pi0403, pi0404, pi0405, pi0406, pi0407, pi0408, pi0409, pi0410, pi0411, pi0412, pi0413, pi0414, pi0415, pi0416, pi0417, pi0418, pi0419, pi0420, pi0421, pi0422, pi0423, pi0424, pi0425, pi0426, pi0427, pi0428, pi0429, pi0430, pi0431, pi0432, pi0433, pi0434, pi0435, pi0436, pi0437, pi0438, pi0439, pi0440, pi0441, pi0442, pi0443, pi0444, pi0445, pi0446, pi0447, pi0448, pi0449, pi0450, pi0451, pi0452, pi0453, pi0454, pi0455, pi0456, pi0457, pi0458, pi0459, pi0460, pi0461, pi0462, pi0463, pi0464, pi0465, pi0466, pi0467, pi0468, pi0469, pi0470, pi0471, pi0472, pi0473, pi0474, pi0475, pi0476, pi0477, pi0478, pi0479, pi0480, pi0481, pi0482, pi0483, pi0484, pi0485, pi0486, pi0487, pi0488, pi0489, pi0490, pi0491, pi0492, pi0493, pi0494, pi0495, pi0496, pi0497, pi0498, pi0499, pi0500, pi0501, pi0502, pi0503, pi0504, pi0505, pi0506, pi0507, pi0508, pi0509, pi0510, pi0511, pi0512, pi0513, pi0514, pi0515, pi0516, pi0517, pi0518, pi0519, pi0520, pi0521, pi0522, pi0523, pi0524, pi0525, pi0526, pi0527, pi0528, pi0529, pi0530, pi0531, pi0532, pi0533, pi0534, pi0535, pi0536, pi0537, pi0538, pi0539, pi0540, pi0541, pi0542, pi0543, pi0544, pi0545, pi0546, pi0547, pi0548, pi0549, pi0550, pi0551, pi0552, pi0553, pi0554, pi0555, pi0556, pi0557, pi0558, pi0559, pi0560, pi0561, pi0562, pi0563, pi0564, pi0565, pi0566, pi0567, pi0568, pi0569, pi0570, pi0571, pi0572, pi0573, pi0574, pi0575, pi0576, pi0577, pi0578, pi0579, pi0580, pi0581, pi0582, pi0583, pi0584, pi0585, pi0586, pi0587, pi0588, pi0589, pi0590, pi0591, pi0592, pi0593, pi0594, pi0595, pi0596, pi0597, pi0598, pi0599, pi0600, pi0601, pi0602, pi0603, pi0604, pi0605, pi0606, pi0607, pi0608, pi0609, pi0610, pi0611, pi0612, pi0613, pi0614, pi0615, pi0616, pi0617, pi0618, pi0619, pi0620, pi0621, pi0622, pi0623, pi0624, pi0625, pi0626, pi0627, pi0628, pi0629, pi0630, pi0631, pi0632, pi0633, pi0634, pi0635, pi0636, pi0637, pi0638, pi0639, pi0640, pi0641, pi0642, pi0643, pi0644, pi0645, pi0646, pi0647, pi0648, pi0649, pi0650, pi0651, pi0652, pi0653, pi0654, pi0655, pi0656, pi0657, pi0658, pi0659, pi0660, pi0661, pi0662, pi0663, pi0664, pi0665, pi0666, pi0667, pi0668, pi0669, pi0670, pi0671, pi0672, pi0673, pi0674, pi0675, pi0676, pi0677, pi0678, pi0679, pi0680, pi0681, pi0682, pi0683, pi0684, pi0685, pi0686, pi0687, pi0688, pi0689, pi0690, pi0691, pi0692, pi0693, pi0694, pi0695, pi0696, pi0697, pi0698, pi0699, pi0700, pi0701, pi0702, pi0703, pi0704, pi0705, pi0706, pi0707, pi0708, pi0709, pi0710, pi0711, pi0712, pi0713, pi0714, pi0715, pi0716, pi0717, pi0718, pi0719, pi0720, pi0721, pi0722, pi0723, pi0724, pi0725, pi0726, pi0727, pi0728, pi0729, pi0730, pi0731, pi0732, pi0733, pi0734, pi0735, pi0736, pi0737, pi0738, pi0739, pi0740, pi0741, pi0742, pi0743, pi0744, pi0745, pi0746, pi0747, pi0748, pi0749, pi0750, pi0751, pi0752, pi0753, pi0754, pi0755, pi0756, pi0757, pi0758, pi0759, pi0760, pi0761, pi0762, pi0763, pi0764, pi0765, pi0766, pi0767, pi0768, pi0769, pi0770, pi0771, pi0772, pi0773, pi0774, pi0775, pi0776, pi0777, pi0778, pi0779, pi0780, pi0781, pi0782, pi0783, pi0784, pi0785, pi0786, pi0787, pi0788, pi0789, pi0790, pi0791, pi0792, pi0793, pi0794, pi0795, pi0796, pi0797, pi0798, pi0799, pi0800, pi0801, pi0802, pi0803, pi0804, pi0805, pi0806, pi0807, pi0808, pi0809, pi0810, pi0811, pi0812, pi0813, pi0814, pi0815, pi0816, pi0817, pi0818, pi0819, pi0820, pi0821, pi0822, pi0823, pi0824, pi0825, pi0826, pi0827, pi0828, pi0829, pi0830, pi0831, pi0832, pi0833, pi0834, pi0835, pi0836, pi0837, pi0838, pi0839, pi0840, pi0841, pi0842, pi0843, pi0844, pi0845, pi0846, pi0847, pi0848, pi0849, pi0850, pi0851, pi0852, pi0853, pi0854, pi0855, pi0856, pi0857, pi0858, pi0859, pi0860, pi0861, pi0862, pi0863, pi0864, pi0865, pi0866, pi0867, pi0868, pi0869, pi0870, pi0871, pi0872, pi0873, pi0874, pi0875, pi0876, pi0877, pi0878, pi0879, pi0880, pi0881, pi0882, pi0883, pi0884, pi0885, pi0886, pi0887, pi0888, pi0889, pi0890, pi0891, pi0892, pi0893, pi0894, pi0895, pi0896, pi0897, pi0898, pi0899, pi0900, pi0901, pi0902, pi0903, pi0904, pi0905, pi0906, pi0907, pi0908, pi0909, pi0910, pi0911, pi0912, pi0913, pi0914, pi0915, pi0916, pi0917, pi0918, pi0919, pi0920, pi0921, pi0922, pi0923, pi0924, pi0925, pi0926, pi0927, pi0928, pi0929, pi0930, pi0931, pi0932, pi0933, pi0934, pi0935, pi0936, pi0937, pi0938, pi0939, pi0940, pi0941, pi0942, pi0943, pi0944, pi0945, pi0946, pi0947, pi0948, pi0949, pi0950, pi0951, pi0952, pi0953, pi0954, pi0955, pi0956, pi0957, pi0958, pi0959, pi0960, pi0961, pi0962, pi0963, pi0964, pi0965, pi0966, pi0967, pi0968, pi0969, pi0970, pi0971, pi0972, pi0973, pi0974, pi0975, pi0976, pi0977, pi0978, pi0979, pi0980, pi0981, pi0982, pi0983, pi0984, pi0985, pi0986, pi0987, pi0988, pi0989, pi0990, pi0991, pi0992, pi0993, pi0994, pi0995, pi0996, pi0997, pi0998, pi0999, pi1000, pi1001, pi1002, pi1003, pi1004, pi1005, pi1006, pi1007, pi1008, pi1009, pi1010, pi1011, pi1012, pi1013, pi1014, pi1015, pi1016, pi1017, pi1018, pi1019, pi1020, pi1021, pi1022, pi1023, pi1024, pi1025, pi1026, pi1027, pi1028, pi1029, pi1030, pi1031, pi1032, pi1033, pi1034, pi1035, pi1036, pi1037, pi1038, pi1039, pi1040, pi1041, pi1042, pi1043, pi1044, pi1045, pi1046, pi1047, pi1048, pi1049, pi1050, pi1051, pi1052, pi1053, pi1054, pi1055, pi1056, pi1057, pi1058, pi1059, pi1060, pi1061, pi1062, pi1063, pi1064, pi1065, pi1066, pi1067, pi1068, pi1069, pi1070, pi1071, pi1072, pi1073, pi1074, pi1075, pi1076, pi1077, pi1078, pi1079, pi1080, pi1081, pi1082, pi1083, pi1084, pi1085, pi1086, pi1087, pi1088, pi1089, pi1090, pi1091, pi1092, pi1093, pi1094, pi1095, pi1096, pi1097, pi1098, pi1099, pi1100, pi1101, pi1102, pi1103, pi1104, pi1105, pi1106, pi1107, pi1108, pi1109, pi1110, pi1111, pi1112, pi1113, pi1114, pi1115, pi1116, pi1117, pi1118, pi1119, pi1120, pi1121, pi1122, pi1123, pi1124, pi1125, pi1126, pi1127, pi1128, pi1129, pi1130, pi1131, pi1132, pi1133, pi1134, pi1135, pi1136, pi1137, pi1138, pi1139, pi1140, pi1141, pi1142, pi1143, pi1144, pi1145, pi1146, pi1147, pi1148, pi1149, pi1150, pi1151, pi1152, pi1153, pi1154, pi1155, pi1156, pi1157, pi1158, pi1159, pi1160, pi1161, pi1162, pi1163, pi1164, pi1165, pi1166, pi1167, pi1168, pi1169, pi1170, pi1171, pi1172, pi1173, pi1174, pi1175, pi1176, pi1177, pi1178, pi1179, pi1180, pi1181, pi1182, pi1183, pi1184, pi1185, pi1186, pi1187, pi1188, pi1189, pi1190, pi1191, pi1192, pi1193, pi1194, pi1195, pi1196, pi1197, pi1198, pi1199, pi1200, pi1201, pi1202, pi1203, pi1204, pi1205, pi1206, pi1207, pi1208, pi1209, pi1210, pi1211, pi1212, pi1213, pi1214, pi1215, pi1216, pi1217, pi1218, pi1219, pi1220, pi1221, pi1222, pi1223, pi1224, pi1225, pi1226, pi1227, pi1228, pi1229, pi1230, pi1231, pi1232, pi1233, pi1234, pi1235, pi1236, pi1237, pi1238, pi1239, pi1240, pi1241, pi1242, pi1243, pi1244, pi1245, pi1246, pi1247, pi1248, pi1249, pi1250, pi1251, pi1252, pi1253, pi1254, pi1255, pi1256, pi1257, pi1258, pi1259, pi1260, pi1261, pi1262, pi1263, pi1264, pi1265, pi1266, pi1267, pi1268, pi1269, pi1270, pi1271, pi1272, pi1273, pi1274, pi1275, pi1276, pi1277, pi1278, pi1279, pi1280, pi1281, pi1282, pi1283, pi1284, pi1285, pi1286, pi1287, pi1288, pi1289, pi1290, pi1291, pi1292, pi1293, pi1294, pi1295, pi1296, pi1297, pi1298, pi1299, pi1300, pi1301, pi1302, pi1303, pi1304, pi1305, pi1306, pi1307, pi1308, pi1309, pi1310, pi1311, pi1312, pi1313, pi1314, pi1315, pi1316, pi1317, pi1318, pi1319, pi1320, pi1321, pi1322, pi1323, pi1324, pi1325, pi1326, pi1327, pi1328, pi1329, pi1330, pi1331, pi1332, pi1333, pi1334, pi1335, pi1336, pi1337, pi1338, pi1339, pi1340, pi1341, pi1342, pi1343, pi1344, pi1345, pi1346, pi1347, pi1348, pi1349, pi1350, pi1351, pi1352, pi1353, pi1354, pi1355, pi1356, pi1357, pi1358, pi1359, pi1360, pi1361, pi1362, pi1363, pi1364, pi1365, pi1366, pi1367, pi1368, pi1369, pi1370, pi1371, pi1372, pi1373, pi1374, pi1375, pi1376, pi1377, pi1378, pi1379, pi1380, pi1381, pi1382, pi1383, pi1384, pi1385, pi1386, pi1387, pi1388, pi1389, pi1390, pi1391, pi1392, pi1393, pi1394, pi1395, pi1396, pi1397, pi1398, pi1399, pi1400, pi1401, pi1402, pi1403, pi1404, pi1405, pi1406, pi1407, pi1408, pi1409, pi1410, pi1411, pi1412, pi1413, pi1414, pi1415, pi1416, pi1417, pi1418, pi1419, pi1420, pi1421, pi1422, pi1423, pi1424, pi1425, pi1426, pi1427, pi1428, pi1429, pi1430, pi1431, pi1432, pi1433, pi1434, pi1435, pi1436, pi1437, pi1438, pi1439, pi1440, pi1441, pi1442, pi1443, pi1444, pi1445, pi1446, pi1447, pi1448, pi1449, pi1450, pi1451, pi1452, pi1453, pi1454, pi1455, pi1456, pi1457, pi1458, pi1459, pi1460, pi1461, pi1462, pi1463, pi1464, pi1465, pi1466, pi1467, pi1468, pi1469, pi1470, pi1471, pi1472, pi1473, pi1474, pi1475, pi1476, pi1477, pi1478, pi1479, pi1480, pi1481, pi1482, pi1483, pi1484, pi1485, pi1486, pi1487, pi1488, pi1489, pi1490, pi1491, pi1492, pi1493, pi1494, pi1495, pi1496, pi1497, pi1498, pi1499, pi1500, pi1501, pi1502, pi1503, pi1504, pi1505, pi1506, pi1507, pi1508, pi1509, pi1510, pi1511, pi1512, pi1513, pi1514, pi1515, pi1516, pi1517, pi1518, pi1519, pi1520, pi1521, pi1522, pi1523, pi1524, pi1525, pi1526, pi1527, pi1528, pi1529, pi1530, pi1531, pi1532, pi1533, pi1534, pi1535, pi1536, pi1537, pi1538, pi1539, pi1540, pi1541, pi1542, pi1543, pi1544, pi1545, pi1546, pi1547, pi1548, pi1549, pi1550, pi1551, pi1552, pi1553, pi1554, pi1555, pi1556, pi1557, pi1558, pi1559, pi1560, pi1561, pi1562, pi1563, pi1564, pi1565, pi1566, pi1567, pi1568, pi1569, pi1570, pi1571, pi1572, pi1573, pi1574, pi1575, pi1576, pi1577, pi1578, pi1579, pi1580, pi1581, pi1582, pi1583, pi1584, pi1585, pi1586, pi1587, pi1588, pi1589, pi1590, pi1591, pi1592, pi1593, pi1594, pi1595, pi1596, pi1597, pi1598, pi1599, pi1600, pi1601, pi1602, pi1603, pi1604, pi1605, pi1606, pi1607, pi1608, pi1609, pi1610, pi1611, pi1612, pi1613, pi1614, pi1615, pi1616, pi1617, pi1618, pi1619, pi1620, pi1621, pi1622, pi1623, pi1624, pi1625, pi1626, pi1627, pi1628, pi1629, pi1630, pi1631, pi1632, pi1633, pi1634, pi1635, pi1636, pi1637, pi1638, pi1639, pi1640, pi1641, pi1642, pi1643, pi1644, pi1645, pi1646, pi1647, pi1648, pi1649, pi1650, pi1651, pi1652, pi1653, pi1654, pi1655, pi1656, pi1657, pi1658, pi1659, pi1660, pi1661, pi1662, pi1663, pi1664, pi1665, pi1666, pi1667, pi1668, pi1669, pi1670, pi1671, pi1672, pi1673, pi1674, pi1675, pi1676, pi1677, pi1678, pi1679, pi1680, pi1681, pi1682, pi1683, pi1684, pi1685, pi1686, pi1687, pi1688, pi1689, pi1690, pi1691, pi1692, pi1693, pi1694, pi1695, pi1696, pi1697, pi1698, pi1699, pi1700, pi1701, pi1702, pi1703, pi1704, pi1705, pi1706, pi1707, pi1708, pi1709, pi1710, pi1711, pi1712, pi1713, pi1714, pi1715, pi1716, pi1717, pi1718, pi1719, pi1720, pi1721, pi1722, pi1723, pi1724, pi1725, pi1726, pi1727, pi1728, pi1729, pi1730, pi1731, pi1732, pi1733, pi1734, pi1735, pi1736, pi1737, pi1738, pi1739, pi1740, pi1741, pi1742, pi1743, pi1744, pi1745, pi1746, pi1747, pi1748, pi1749, pi1750, pi1751, pi1752, pi1753, pi1754, pi1755, pi1756, pi1757, pi1758, pi1759, pi1760, pi1761, pi1762, pi1763, pi1764, pi1765, pi1766, pi1767, pi1768, pi1769, pi1770, pi1771, pi1772, pi1773, pi1774, pi1775, pi1776, pi1777, pi1778, pi1779, pi1780, pi1781, pi1782, pi1783, pi1784, pi1785, pi1786, pi1787, pi1788, pi1789, pi1790, pi1791, pi1792, pi1793, pi1794, pi1795, pi1796, pi1797, pi1798, pi1799, pi1800, pi1801, pi1802, pi1803, pi1804, pi1805, pi1806, pi1807, pi1808, pi1809, pi1810, pi1811, pi1812, pi1813, pi1814, pi1815, pi1816, pi1817, pi1818, pi1819, pi1820, pi1821, pi1822, pi1823, pi1824, pi1825, pi1826, pi1827, pi1828, pi1829, pi1830, pi1831, pi1832, pi1833, pi1834, pi1835, pi1836, pi1837, pi1838, pi1839, pi1840, pi1841, pi1842, pi1843, pi1844, pi1845, pi1846, pi1847, pi1848, pi1849, pi1850, pi1851, pi1852, pi1853, pi1854, pi1855, pi1856, pi1857, pi1858, pi1859;
output po0000, po0001, po0002, po0003, po0004, po0005, po0006, po0007, po0008, po0009, po0010, po0011, po0012, po0013, po0014, po0015, po0016, po0017, po0018, po0019, po0020, po0021, po0022, po0023, po0024, po0025, po0026, po0027, po0028, po0029, po0030, po0031, po0032, po0033, po0034, po0035, po0036, po0037, po0038, po0039, po0040, po0041, po0042, po0043, po0044, po0045, po0046, po0047, po0048, po0049, po0050, po0051, po0052, po0053, po0054, po0055, po0056, po0057, po0058, po0059, po0060, po0061, po0062, po0063, po0064, po0065, po0066, po0067, po0068, po0069, po0070, po0071, po0072, po0073, po0074, po0075, po0076, po0077, po0078, po0079, po0080, po0081, po0082, po0083, po0084, po0085, po0086, po0087, po0088, po0089, po0090, po0091, po0092, po0093, po0094, po0095, po0096, po0097, po0098, po0099, po0100, po0101, po0102, po0103, po0104, po0105, po0106, po0107, po0108, po0109, po0110, po0111, po0112, po0113, po0114, po0115, po0116, po0117, po0118, po0119, po0120, po0121, po0122, po0123, po0124, po0125, po0126, po0127, po0128, po0129, po0130, po0131, po0132, po0133, po0134, po0135, po0136, po0137, po0138, po0139, po0140, po0141, po0142, po0143, po0144, po0145, po0146, po0147, po0148, po0149, po0150, po0151, po0152, po0153, po0154, po0155, po0156, po0157, po0158, po0159, po0160, po0161, po0162, po0163, po0164, po0165, po0166, po0167, po0168, po0169, po0170, po0171, po0172, po0173, po0174, po0175, po0176, po0177, po0178, po0179, po0180, po0181, po0182, po0183, po0184, po0185, po0186, po0187, po0188, po0189, po0190, po0191, po0192, po0193, po0194, po0195, po0196, po0197, po0198, po0199, po0200, po0201, po0202, po0203, po0204, po0205, po0206, po0207, po0208, po0209, po0210, po0211, po0212, po0213, po0214, po0215, po0216, po0217, po0218, po0219, po0220, po0221, po0222, po0223, po0224, po0225, po0226, po0227, po0228, po0229, po0230, po0231, po0232, po0233, po0234, po0235, po0236, po0237, po0238, po0239, po0240, po0241, po0242, po0243, po0244, po0245, po0246, po0247, po0248, po0249, po0250, po0251, po0252, po0253, po0254, po0255, po0256, po0257, po0258, po0259, po0260, po0261, po0262, po0263, po0264, po0265, po0266, po0267, po0268, po0269, po0270, po0271, po0272, po0273, po0274, po0275, po0276, po0277, po0278, po0279, po0280, po0281, po0282, po0283, po0284, po0285, po0286, po0287, po0288, po0289, po0290, po0291, po0292, po0293, po0294, po0295, po0296, po0297, po0298, po0299, po0300, po0301, po0302, po0303, po0304, po0305, po0306, po0307, po0308, po0309, po0310, po0311, po0312, po0313, po0314, po0315, po0316, po0317, po0318, po0319, po0320, po0321, po0322, po0323, po0324, po0325, po0326, po0327, po0328, po0329, po0330, po0331, po0332, po0333, po0334, po0335, po0336, po0337, po0338, po0339, po0340, po0341, po0342, po0343, po0344, po0345, po0346, po0347, po0348, po0349, po0350, po0351, po0352, po0353, po0354, po0355, po0356, po0357, po0358, po0359, po0360, po0361, po0362, po0363, po0364, po0365, po0366, po0367, po0368, po0369, po0370, po0371, po0372, po0373, po0374, po0375, po0376, po0377, po0378, po0379, po0380, po0381, po0382, po0383, po0384, po0385, po0386, po0387, po0388, po0389, po0390, po0391, po0392, po0393, po0394, po0395, po0396, po0397, po0398, po0399, po0400, po0401, po0402, po0403, po0404, po0405, po0406, po0407, po0408, po0409, po0410, po0411, po0412, po0413, po0414, po0415, po0416, po0417, po0418, po0419, po0420, po0421, po0422, po0423, po0424, po0425, po0426, po0427, po0428, po0429, po0430, po0431, po0432, po0433, po0434, po0435, po0436, po0437, po0438, po0439, po0440, po0441, po0442, po0443, po0444, po0445, po0446, po0447, po0448, po0449, po0450, po0451, po0452, po0453, po0454, po0455, po0456, po0457, po0458, po0459, po0460, po0461, po0462, po0463, po0464, po0465, po0466, po0467, po0468, po0469, po0470, po0471, po0472, po0473, po0474, po0475, po0476, po0477, po0478, po0479, po0480, po0481, po0482, po0483, po0484, po0485, po0486, po0487, po0488, po0489, po0490, po0491, po0492, po0493, po0494, po0495, po0496, po0497, po0498, po0499, po0500, po0501, po0502, po0503, po0504, po0505, po0506, po0507, po0508, po0509, po0510, po0511, po0512, po0513, po0514, po0515, po0516, po0517, po0518, po0519, po0520, po0521, po0522, po0523, po0524, po0525, po0526, po0527, po0528, po0529, po0530, po0531, po0532, po0533, po0534, po0535, po0536, po0537, po0538, po0539, po0540, po0541, po0542, po0543, po0544, po0545, po0546, po0547, po0548, po0549, po0550, po0551, po0552, po0553, po0554, po0555, po0556, po0557, po0558, po0559, po0560, po0561, po0562, po0563, po0564, po0565, po0566, po0567, po0568, po0569, po0570, po0571, po0572, po0573, po0574, po0575, po0576, po0577, po0578, po0579, po0580, po0581, po0582, po0583, po0584, po0585, po0586, po0587, po0588, po0589, po0590, po0591, po0592, po0593, po0594, po0595, po0596, po0597, po0598, po0599, po0600, po0601, po0602, po0603, po0604, po0605, po0606, po0607, po0608, po0609, po0610, po0611, po0612, po0613, po0614, po0615, po0616, po0617, po0618, po0619, po0620, po0621, po0622, po0623, po0624, po0625, po0626, po0627, po0628, po0629, po0630, po0631, po0632, po0633, po0634, po0635, po0636, po0637, po0638, po0639, po0640, po0641, po0642, po0643, po0644, po0645, po0646, po0647, po0648, po0649, po0650, po0651, po0652, po0653, po0654, po0655, po0656, po0657, po0658, po0659, po0660, po0661, po0662, po0663, po0664, po0665, po0666, po0667, po0668, po0669, po0670, po0671, po0672, po0673, po0674, po0675, po0676, po0677, po0678, po0679, po0680, po0681, po0682, po0683, po0684, po0685, po0686, po0687, po0688, po0689, po0690, po0691, po0692, po0693, po0694, po0695, po0696, po0697, po0698, po0699, po0700, po0701, po0702, po0703, po0704, po0705, po0706, po0707, po0708, po0709, po0710, po0711, po0712, po0713, po0714, po0715, po0716, po0717, po0718, po0719, po0720, po0721, po0722, po0723, po0724, po0725, po0726, po0727, po0728, po0729, po0730, po0731, po0732, po0733, po0734, po0735, po0736, po0737, po0738, po0739, po0740, po0741, po0742, po0743, po0744, po0745, po0746, po0747, po0748, po0749, po0750, po0751, po0752, po0753, po0754, po0755, po0756, po0757, po0758, po0759, po0760, po0761, po0762, po0763, po0764, po0765, po0766, po0767, po0768, po0769, po0770, po0771, po0772, po0773, po0774, po0775, po0776, po0777, po0778, po0779, po0780, po0781, po0782, po0783, po0784, po0785, po0786, po0787, po0788, po0789, po0790, po0791, po0792, po0793, po0794, po0795, po0796, po0797, po0798, po0799, po0800, po0801, po0802, po0803, po0804, po0805, po0806, po0807, po0808, po0809, po0810, po0811, po0812, po0813, po0814, po0815, po0816, po0817, po0818, po0819, po0820, po0821, po0822, po0823, po0824, po0825, po0826, po0827, po0828, po0829, po0830, po0831, po0832, po0833, po0834, po0835, po0836, po0837, po0838, po0839, po0840, po0841, po0842, po0843, po0844, po0845, po0846, po0847, po0848, po0849, po0850, po0851, po0852, po0853, po0854, po0855, po0856, po0857, po0858, po0859, po0860, po0861, po0862, po0863, po0864, po0865, po0866, po0867, po0868, po0869, po0870, po0871, po0872, po0873, po0874, po0875, po0876, po0877, po0878, po0879, po0880, po0881, po0882, po0883, po0884, po0885, po0886, po0887, po0888, po0889, po0890, po0891, po0892, po0893, po0894, po0895, po0896, po0897, po0898, po0899, po0900, po0901, po0902, po0903, po0904, po0905, po0906, po0907, po0908, po0909, po0910, po0911, po0912, po0913, po0914, po0915, po0916, po0917, po0918, po0919, po0920, po0921, po0922, po0923, po0924, po0925, po0926, po0927, po0928, po0929, po0930, po0931, po0932, po0933, po0934, po0935, po0936, po0937, po0938, po0939, po0940, po0941, po0942, po0943, po0944, po0945, po0946, po0947, po0948, po0949, po0950, po0951, po0952, po0953, po0954, po0955, po0956, po0957, po0958, po0959, po0960, po0961, po0962, po0963, po0964, po0965, po0966, po0967, po0968, po0969, po0970, po0971, po0972, po0973, po0974, po0975, po0976, po0977, po0978, po0979, po0980, po0981, po0982, po0983, po0984, po0985, po0986, po0987, po0988, po0989, po0990, po0991, po0992, po0993, po0994, po0995, po0996, po0997, po0998, po0999, po1000, po1001, po1002, po1003, po1004, po1005, po1006, po1007, po1008, po1009, po1010, po1011, po1012, po1013, po1014, po1015, po1016, po1017, po1018, po1019, po1020, po1021, po1022, po1023, po1024, po1025, po1026, po1027, po1028, po1029, po1030, po1031, po1032, po1033, po1034, po1035, po1036, po1037, po1038, po1039, po1040, po1041, po1042, po1043, po1044, po1045, po1046, po1047, po1048, po1049, po1050, po1051, po1052, po1053, po1054, po1055, po1056, po1057, po1058, po1059, po1060, po1061, po1062, po1063, po1064, po1065, po1066, po1067, po1068, po1069, po1070, po1071, po1072, po1073, po1074, po1075, po1076, po1077, po1078, po1079, po1080, po1081, po1082, po1083, po1084, po1085, po1086, po1087, po1088, po1089, po1090, po1091, po1092, po1093, po1094, po1095, po1096, po1097, po1098, po1099, po1100, po1101, po1102, po1103, po1104, po1105, po1106, po1107, po1108, po1109, po1110, po1111, po1112, po1113, po1114, po1115, po1116, po1117, po1118, po1119, po1120, po1121, po1122, po1123, po1124, po1125, po1126, po1127, po1128, po1129, po1130, po1131, po1132, po1133, po1134, po1135, po1136, po1137, po1138, po1139, po1140, po1141, po1142, po1143, po1144, po1145, po1146, po1147, po1148, po1149, po1150, po1151, po1152, po1153, po1154, po1155, po1156, po1157, po1158, po1159, po1160, po1161, po1162, po1163, po1164, po1165, po1166, po1167, po1168, po1169, po1170, po1171, po1172, po1173, po1174, po1175, po1176, po1177, po1178, po1179, po1180, po1181, po1182, po1183, po1184, po1185, po1186, po1187, po1188, po1189, po1190, po1191, po1192, po1193, po1194, po1195, po1196, po1197, po1198, po1199, po1200, po1201, po1202, po1203, po1204, po1205, po1206, po1207, po1208, po1209, po1210, po1211, po1212, po1213, po1214, po1215, po1216, po1217, po1218, po1219, po1220, po1221, po1222, po1223, po1224, po1225, po1226, po1227, po1228, po1229, po1230, po1231, po1232, po1233, po1234, po1235, po1236, po1237, po1238, po1239, po1240, po1241, po1242, po1243, po1244, po1245, po1246, po1247, po1248, po1249, po1250, po1251, po1252, po1253, po1254, po1255, po1256, po1257, po1258, po1259, po1260, po1261, po1262, po1263, po1264, po1265, po1266, po1267, po1268, po1269, po1270, po1271, po1272, po1273, po1274, po1275, po1276, po1277, po1278, po1279, po1280, po1281, po1282, po1283, po1284, po1285, po1286, po1287, po1288, po1289, po1290, po1291, po1292, po1293, po1294, po1295, po1296, po1297, po1298, po1299, po1300, po1301, po1302, po1303, po1304, po1305, po1306, po1307, po1308, po1309, po1310, po1311, po1312, po1313, po1314, po1315, po1316, po1317, po1318, po1319, po1320, po1321, po1322, po1323, po1324, po1325, po1326, po1327, po1328, po1329, po1330, po1331, po1332, po1333, po1334, po1335, po1336, po1337, po1338, po1339, po1340, po1341, po1342, po1343, po1344, po1345, po1346, po1347, po1348, po1349, po1350, po1351, po1352, po1353, po1354, po1355, po1356, po1357, po1358, po1359, po1360, po1361, po1362, po1363, po1364, po1365, po1366, po1367, po1368, po1369, po1370, po1371, po1372, po1373, po1374, po1375, po1376, po1377, po1378, po1379, po1380, po1381, po1382, po1383, po1384, po1385, po1386, po1387, po1388, po1389, po1390, po1391, po1392, po1393, po1394, po1395, po1396, po1397, po1398, po1399, po1400, po1401, po1402, po1403, po1404, po1405, po1406, po1407, po1408, po1409, po1410, po1411, po1412, po1413, po1414, po1415, po1416, po1417, po1418, po1419, po1420, po1421, po1422, po1423, po1424, po1425, po1426, po1427, po1428, po1429, po1430, po1431, po1432, po1433, po1434, po1435, po1436, po1437, po1438, po1439, po1440, po1441, po1442, po1443, po1444, po1445, po1446, po1447, po1448, po1449, po1450, po1451, po1452, po1453, po1454, po1455, po1456, po1457, po1458, po1459, po1460, po1461, po1462, po1463, po1464, po1465, po1466, po1467, po1468, po1469, po1470, po1471, po1472, po1473, po1474, po1475, po1476, po1477, po1478, po1479, po1480, po1481, po1482, po1483, po1484, po1485, po1486, po1487, po1488, po1489, po1490, po1491, po1492, po1493, po1494, po1495, po1496, po1497, po1498, po1499, po1500, po1501, po1502, po1503, po1504, po1505, po1506, po1507, po1508, po1509, po1510, po1511, po1512, po1513, po1514, po1515, po1516, po1517, po1518, po1519, po1520, po1521, po1522, po1523, po1524, po1525, po1526, po1527, po1528, po1529, po1530, po1531, po1532, po1533, po1534, po1535, po1536, po1537, po1538, po1539, po1540, po1541, po1542, po1543, po1544, po1545, po1546, po1547, po1548, po1549, po1550, po1551, po1552, po1553, po1554, po1555, po1556, po1557, po1558, po1559, po1560, po1561, po1562, po1563, po1564, po1565, po1566, po1567, po1568, po1569, po1570, po1571, po1572, po1573, po1574, po1575, po1576, po1577, po1578, po1579, po1580, po1581, po1582, po1583, po1584, po1585, po1586, po1587, po1588, po1589, po1590, po1591, po1592, po1593, po1594, po1595, po1596, po1597, po1598, po1599, po1600, po1601, po1602, po1603, po1604, po1605, po1606, po1607, po1608, po1609, po1610, po1611, po1612, po1613, po1614, po1615, po1616, po1617, po1618, po1619, po1620, po1621, po1622, po1623, po1624, po1625, po1626, po1627, po1628, po1629, po1630, po1631, po1632, po1633, po1634, po1635, po1636, po1637, po1638, po1639, po1640, po1641, po1642, po1643, po1644, po1645, po1646, po1647, po1648, po1649, po1650, po1651, po1652, po1653, po1654, po1655, po1656, po1657, po1658, po1659, po1660, po1661, po1662, po1663, po1664, po1665, po1666, po1667, po1668, po1669, po1670, po1671, po1672, po1673, po1674, po1675, po1676, po1677, po1678, po1679, po1680, po1681, po1682, po1683, po1684, po1685, po1686, po1687, po1688, po1689, po1690, po1691, po1692, po1693, po1694, po1695, po1696, po1697, po1698, po1699, po1700, po1701, po1702, po1703, po1704, po1705, po1706, po1707, po1708, po1709, po1710, po1711, po1712, po1713, po1714, po1715, po1716, po1717, po1718, po1719, po1720, po1721, po1722, po1723, po1724, po1725, po1726, po1727, po1728, po1729, po1730, po1731, po1732, po1733, po1734, po1735, po1736, po1737, po1738, po1739, po1740, po1741, po1742, po1743, po1744, po1745, po1746, po1747, po1748, po1749, po1750, po1751, po1752, po1753, po1754, po1755, po1756, po1757, po1758, po1759, po1760, po1761, po1762, po1763, po1764, po1765, po1766, po1767, po1768, po1769, po1770, po1771, po1772, po1773, po1774, po1775, po1776, po1777, po1778, po1779, po1780, po1781, po1782, po1783, po1784, po1785, po1786, po1787, po1788, po1789, po1790, po1791, po1792, po1793, po1794, po1795, po1796, po1797, po1798, po1799, po1800, po1801, po1802, po1803, po1804, po1805, po1806, po1807, po1808, po1809, po1810, po1811, po1812, po1813, po1814, po1815, po1816, po1817, po1818, po1819, po1820, po1821, po1822, po1823, po1824, po1825, po1826, po1827, po1828, po1829, po1830, po1831, po1832, po1833, po1834, po1835, po1836, po1837, po1838, po1839, po1840, po1841, po1842, po1843, po1844, po1845;
wire one, w0, w1, w2, w3, w4, w5, w6, w7, w8, w9, w10, w11, w12, w13, w14, w15, w16, w17, w18, w19, w20, w21, w22, w23, w24, w25, w26, w27, w28, w29, w30, w31, w32, w33, w34, w35, w36, w37, w38, w39, w40, w41, w42, w43, w44, w45, w46, w47, w48, w49, w50, w51, w52, w53, w54, w55, w56, w57, w58, w59, w60, w61, w62, w63, w64, w65, w66, w67, w68, w69, w70, w71, w72, w73, w74, w75, w76, w77, w78, w79, w80, w81, w82, w83, w84, w85, w86, w87, w88, w89, w90, w91, w92, w93, w94, w95, w96, w97, w98, w99, w100, w101, w102, w103, w104, w105, w106, w107, w108, w109, w110, w111, w112, w113, w114, w115, w116, w117, w118, w119, w120, w121, w122, w123, w124, w125, w126, w127, w128, w129, w130, w131, w132, w133, w134, w135, w136, w137, w138, w139, w140, w141, w142, w143, w144, w145, w146, w147, w148, w149, w150, w151, w152, w153, w154, w155, w156, w157, w158, w159, w160, w161, w162, w163, w164, w165, w166, w167, w168, w169, w170, w171, w172, w173, w174, w175, w176, w177, w178, w179, w180, w181, w182, w183, w184, w185, w186, w187, w188, w189, w190, w191, w192, w193, w194, w195, w196, w197, w198, w199, w200, w201, w202, w203, w204, w205, w206, w207, w208, w209, w210, w211, w212, w213, w214, w215, w216, w217, w218, w219, w220, w221, w222, w223, w224, w225, w226, w227, w228, w229, w230, w231, w232, w233, w234, w235, w236, w237, w238, w239, w240, w241, w242, w243, w244, w245, w246, w247, w248, w249, w250, w251, w252, w253, w254, w255, w256, w257, w258, w259, w260, w261, w262, w263, w264, w265, w266, w267, w268, w269, w270, w271, w272, w273, w274, w275, w276, w277, w278, w279, w280, w281, w282, w283, w284, w285, w286, w287, w288, w289, w290, w291, w292, w293, w294, w295, w296, w297, w298, w299, w300, w301, w302, w303, w304, w305, w306, w307, w308, w309, w310, w311, w312, w313, w314, w315, w316, w317, w318, w319, w320, w321, w322, w323, w324, w325, w326, w327, w328, w329, w330, w331, w332, w333, w334, w335, w336, w337, w338, w339, w340, w341, w342, w343, w344, w345, w346, w347, w348, w349, w350, w351, w352, w353, w354, w355, w356, w357, w358, w359, w360, w361, w362, w363, w364, w365, w366, w367, w368, w369, w370, w371, w372, w373, w374, w375, w376, w377, w378, w379, w380, w381, w382, w383, w384, w385, w386, w387, w388, w389, w390, w391, w392, w393, w394, w395, w396, w397, w398, w399, w400, w401, w402, w403, w404, w405, w406, w407, w408, w409, w410, w411, w412, w413, w414, w415, w416, w417, w418, w419, w420, w421, w422, w423, w424, w425, w426, w427, w428, w429, w430, w431, w432, w433, w434, w435, w436, w437, w438, w439, w440, w441, w442, w443, w444, w445, w446, w447, w448, w449, w450, w451, w452, w453, w454, w455, w456, w457, w458, w459, w460, w461, w462, w463, w464, w465, w466, w467, w468, w469, w470, w471, w472, w473, w474, w475, w476, w477, w478, w479, w480, w481, w482, w483, w484, w485, w486, w487, w488, w489, w490, w491, w492, w493, w494, w495, w496, w497, w498, w499, w500, w501, w502, w503, w504, w505, w506, w507, w508, w509, w510, w511, w512, w513, w514, w515, w516, w517, w518, w519, w520, w521, w522, w523, w524, w525, w526, w527, w528, w529, w530, w531, w532, w533, w534, w535, w536, w537, w538, w539, w540, w541, w542, w543, w544, w545, w546, w547, w548, w549, w550, w551, w552, w553, w554, w555, w556, w557, w558, w559, w560, w561, w562, w563, w564, w565, w566, w567, w568, w569, w570, w571, w572, w573, w574, w575, w576, w577, w578, w579, w580, w581, w582, w583, w584, w585, w586, w587, w588, w589, w590, w591, w592, w593, w594, w595, w596, w597, w598, w599, w600, w601, w602, w603, w604, w605, w606, w607, w608, w609, w610, w611, w612, w613, w614, w615, w616, w617, w618, w619, w620, w621, w622, w623, w624, w625, w626, w627, w628, w629, w630, w631, w632, w633, w634, w635, w636, w637, w638, w639, w640, w641, w642, w643, w644, w645, w646, w647, w648, w649, w650, w651, w652, w653, w654, w655, w656, w657, w658, w659, w660, w661, w662, w663, w664, w665, w666, w667, w668, w669, w670, w671, w672, w673, w674, w675, w676, w677, w678, w679, w680, w681, w682, w683, w684, w685, w686, w687, w688, w689, w690, w691, w692, w693, w694, w695, w696, w697, w698, w699, w700, w701, w702, w703, w704, w705, w706, w707, w708, w709, w710, w711, w712, w713, w714, w715, w716, w717, w718, w719, w720, w721, w722, w723, w724, w725, w726, w727, w728, w729, w730, w731, w732, w733, w734, w735, w736, w737, w738, w739, w740, w741, w742, w743, w744, w745, w746, w747, w748, w749, w750, w751, w752, w753, w754, w755, w756, w757, w758, w759, w760, w761, w762, w763, w764, w765, w766, w767, w768, w769, w770, w771, w772, w773, w774, w775, w776, w777, w778, w779, w780, w781, w782, w783, w784, w785, w786, w787, w788, w789, w790, w791, w792, w793, w794, w795, w796, w797, w798, w799, w800, w801, w802, w803, w804, w805, w806, w807, w808, w809, w810, w811, w812, w813, w814, w815, w816, w817, w818, w819, w820, w821, w822, w823, w824, w825, w826, w827, w828, w829, w830, w831, w832, w833, w834, w835, w836, w837, w838, w839, w840, w841, w842, w843, w844, w845, w846, w847, w848, w849, w850, w851, w852, w853, w854, w855, w856, w857, w858, w859, w860, w861, w862, w863, w864, w865, w866, w867, w868, w869, w870, w871, w872, w873, w874, w875, w876, w877, w878, w879, w880, w881, w882, w883, w884, w885, w886, w887, w888, w889, w890, w891, w892, w893, w894, w895, w896, w897, w898, w899, w900, w901, w902, w903, w904, w905, w906, w907, w908, w909, w910, w911, w912, w913, w914, w915, w916, w917, w918, w919, w920, w921, w922, w923, w924, w925, w926, w927, w928, w929, w930, w931, w932, w933, w934, w935, w936, w937, w938, w939, w940, w941, w942, w943, w944, w945, w946, w947, w948, w949, w950, w951, w952, w953, w954, w955, w956, w957, w958, w959, w960, w961, w962, w963, w964, w965, w966, w967, w968, w969, w970, w971, w972, w973, w974, w975, w976, w977, w978, w979, w980, w981, w982, w983, w984, w985, w986, w987, w988, w989, w990, w991, w992, w993, w994, w995, w996, w997, w998, w999, w1000, w1001, w1002, w1003, w1004, w1005, w1006, w1007, w1008, w1009, w1010, w1011, w1012, w1013, w1014, w1015, w1016, w1017, w1018, w1019, w1020, w1021, w1022, w1023, w1024, w1025, w1026, w1027, w1028, w1029, w1030, w1031, w1032, w1033, w1034, w1035, w1036, w1037, w1038, w1039, w1040, w1041, w1042, w1043, w1044, w1045, w1046, w1047, w1048, w1049, w1050, w1051, w1052, w1053, w1054, w1055, w1056, w1057, w1058, w1059, w1060, w1061, w1062, w1063, w1064, w1065, w1066, w1067, w1068, w1069, w1070, w1071, w1072, w1073, w1074, w1075, w1076, w1077, w1078, w1079, w1080, w1081, w1082, w1083, w1084, w1085, w1086, w1087, w1088, w1089, w1090, w1091, w1092, w1093, w1094, w1095, w1096, w1097, w1098, w1099, w1100, w1101, w1102, w1103, w1104, w1105, w1106, w1107, w1108, w1109, w1110, w1111, w1112, w1113, w1114, w1115, w1116, w1117, w1118, w1119, w1120, w1121, w1122, w1123, w1124, w1125, w1126, w1127, w1128, w1129, w1130, w1131, w1132, w1133, w1134, w1135, w1136, w1137, w1138, w1139, w1140, w1141, w1142, w1143, w1144, w1145, w1146, w1147, w1148, w1149, w1150, w1151, w1152, w1153, w1154, w1155, w1156, w1157, w1158, w1159, w1160, w1161, w1162, w1163, w1164, w1165, w1166, w1167, w1168, w1169, w1170, w1171, w1172, w1173, w1174, w1175, w1176, w1177, w1178, w1179, w1180, w1181, w1182, w1183, w1184, w1185, w1186, w1187, w1188, w1189, w1190, w1191, w1192, w1193, w1194, w1195, w1196, w1197, w1198, w1199, w1200, w1201, w1202, w1203, w1204, w1205, w1206, w1207, w1208, w1209, w1210, w1211, w1212, w1213, w1214, w1215, w1216, w1217, w1218, w1219, w1220, w1221, w1222, w1223, w1224, w1225, w1226, w1227, w1228, w1229, w1230, w1231, w1232, w1233, w1234, w1235, w1236, w1237, w1238, w1239, w1240, w1241, w1242, w1243, w1244, w1245, w1246, w1247, w1248, w1249, w1250, w1251, w1252, w1253, w1254, w1255, w1256, w1257, w1258, w1259, w1260, w1261, w1262, w1263, w1264, w1265, w1266, w1267, w1268, w1269, w1270, w1271, w1272, w1273, w1274, w1275, w1276, w1277, w1278, w1279, w1280, w1281, w1282, w1283, w1284, w1285, w1286, w1287, w1288, w1289, w1290, w1291, w1292, w1293, w1294, w1295, w1296, w1297, w1298, w1299, w1300, w1301, w1302, w1303, w1304, w1305, w1306, w1307, w1308, w1309, w1310, w1311, w1312, w1313, w1314, w1315, w1316, w1317, w1318, w1319, w1320, w1321, w1322, w1323, w1324, w1325, w1326, w1327, w1328, w1329, w1330, w1331, w1332, w1333, w1334, w1335, w1336, w1337, w1338, w1339, w1340, w1341, w1342, w1343, w1344, w1345, w1346, w1347, w1348, w1349, w1350, w1351, w1352, w1353, w1354, w1355, w1356, w1357, w1358, w1359, w1360, w1361, w1362, w1363, w1364, w1365, w1366, w1367, w1368, w1369, w1370, w1371, w1372, w1373, w1374, w1375, w1376, w1377, w1378, w1379, w1380, w1381, w1382, w1383, w1384, w1385, w1386, w1387, w1388, w1389, w1390, w1391, w1392, w1393, w1394, w1395, w1396, w1397, w1398, w1399, w1400, w1401, w1402, w1403, w1404, w1405, w1406, w1407, w1408, w1409, w1410, w1411, w1412, w1413, w1414, w1415, w1416, w1417, w1418, w1419, w1420, w1421, w1422, w1423, w1424, w1425, w1426, w1427, w1428, w1429, w1430, w1431, w1432, w1433, w1434, w1435, w1436, w1437, w1438, w1439, w1440, w1441, w1442, w1443, w1444, w1445, w1446, w1447, w1448, w1449, w1450, w1451, w1452, w1453, w1454, w1455, w1456, w1457, w1458, w1459, w1460, w1461, w1462, w1463, w1464, w1465, w1466, w1467, w1468, w1469, w1470, w1471, w1472, w1473, w1474, w1475, w1476, w1477, w1478, w1479, w1480, w1481, w1482, w1483, w1484, w1485, w1486, w1487, w1488, w1489, w1490, w1491, w1492, w1493, w1494, w1495, w1496, w1497, w1498, w1499, w1500, w1501, w1502, w1503, w1504, w1505, w1506, w1507, w1508, w1509, w1510, w1511, w1512, w1513, w1514, w1515, w1516, w1517, w1518, w1519, w1520, w1521, w1522, w1523, w1524, w1525, w1526, w1527, w1528, w1529, w1530, w1531, w1532, w1533, w1534, w1535, w1536, w1537, w1538, w1539, w1540, w1541, w1542, w1543, w1544, w1545, w1546, w1547, w1548, w1549, w1550, w1551, w1552, w1553, w1554, w1555, w1556, w1557, w1558, w1559, w1560, w1561, w1562, w1563, w1564, w1565, w1566, w1567, w1568, w1569, w1570, w1571, w1572, w1573, w1574, w1575, w1576, w1577, w1578, w1579, w1580, w1581, w1582, w1583, w1584, w1585, w1586, w1587, w1588, w1589, w1590, w1591, w1592, w1593, w1594, w1595, w1596, w1597, w1598, w1599, w1600, w1601, w1602, w1603, w1604, w1605, w1606, w1607, w1608, w1609, w1610, w1611, w1612, w1613, w1614, w1615, w1616, w1617, w1618, w1619, w1620, w1621, w1622, w1623, w1624, w1625, w1626, w1627, w1628, w1629, w1630, w1631, w1632, w1633, w1634, w1635, w1636, w1637, w1638, w1639, w1640, w1641, w1642, w1643, w1644, w1645, w1646, w1647, w1648, w1649, w1650, w1651, w1652, w1653, w1654, w1655, w1656, w1657, w1658, w1659, w1660, w1661, w1662, w1663, w1664, w1665, w1666, w1667, w1668, w1669, w1670, w1671, w1672, w1673, w1674, w1675, w1676, w1677, w1678, w1679, w1680, w1681, w1682, w1683, w1684, w1685, w1686, w1687, w1688, w1689, w1690, w1691, w1692, w1693, w1694, w1695, w1696, w1697, w1698, w1699, w1700, w1701, w1702, w1703, w1704, w1705, w1706, w1707, w1708, w1709, w1710, w1711, w1712, w1713, w1714, w1715, w1716, w1717, w1718, w1719, w1720, w1721, w1722, w1723, w1724, w1725, w1726, w1727, w1728, w1729, w1730, w1731, w1732, w1733, w1734, w1735, w1736, w1737, w1738, w1739, w1740, w1741, w1742, w1743, w1744, w1745, w1746, w1747, w1748, w1749, w1750, w1751, w1752, w1753, w1754, w1755, w1756, w1757, w1758, w1759, w1760, w1761, w1762, w1763, w1764, w1765, w1766, w1767, w1768, w1769, w1770, w1771, w1772, w1773, w1774, w1775, w1776, w1777, w1778, w1779, w1780, w1781, w1782, w1783, w1784, w1785, w1786, w1787, w1788, w1789, w1790, w1791, w1792, w1793, w1794, w1795, w1796, w1797, w1798, w1799, w1800, w1801, w1802, w1803, w1804, w1805, w1806, w1807, w1808, w1809, w1810, w1811, w1812, w1813, w1814, w1815, w1816, w1817, w1818, w1819, w1820, w1821, w1822, w1823, w1824, w1825, w1826, w1827, w1828, w1829, w1830, w1831, w1832, w1833, w1834, w1835, w1836, w1837, w1838, w1839, w1840, w1841, w1842, w1843, w1844, w1845, w1846, w1847, w1848, w1849, w1850, w1851, w1852, w1853, w1854, w1855, w1856, w1857, w1858, w1859, w1860, w1861, w1862, w1863, w1864, w1865, w1866, w1867, w1868, w1869, w1870, w1871, w1872, w1873, w1874, w1875, w1876, w1877, w1878, w1879, w1880, w1881, w1882, w1883, w1884, w1885, w1886, w1887, w1888, w1889, w1890, w1891, w1892, w1893, w1894, w1895, w1896, w1897, w1898, w1899, w1900, w1901, w1902, w1903, w1904, w1905, w1906, w1907, w1908, w1909, w1910, w1911, w1912, w1913, w1914, w1915, w1916, w1917, w1918, w1919, w1920, w1921, w1922, w1923, w1924, w1925, w1926, w1927, w1928, w1929, w1930, w1931, w1932, w1933, w1934, w1935, w1936, w1937, w1938, w1939, w1940, w1941, w1942, w1943, w1944, w1945, w1946, w1947, w1948, w1949, w1950, w1951, w1952, w1953, w1954, w1955, w1956, w1957, w1958, w1959, w1960, w1961, w1962, w1963, w1964, w1965, w1966, w1967, w1968, w1969, w1970, w1971, w1972, w1973, w1974, w1975, w1976, w1977, w1978, w1979, w1980, w1981, w1982, w1983, w1984, w1985, w1986, w1987, w1988, w1989, w1990, w1991, w1992, w1993, w1994, w1995, w1996, w1997, w1998, w1999, w2000, w2001, w2002, w2003, w2004, w2005, w2006, w2007, w2008, w2009, w2010, w2011, w2012, w2013, w2014, w2015, w2016, w2017, w2018, w2019, w2020, w2021, w2022, w2023, w2024, w2025, w2026, w2027, w2028, w2029, w2030, w2031, w2032, w2033, w2034, w2035, w2036, w2037, w2038, w2039, w2040, w2041, w2042, w2043, w2044, w2045, w2046, w2047, w2048, w2049, w2050, w2051, w2052, w2053, w2054, w2055, w2056, w2057, w2058, w2059, w2060, w2061, w2062, w2063, w2064, w2065, w2066, w2067, w2068, w2069, w2070, w2071, w2072, w2073, w2074, w2075, w2076, w2077, w2078, w2079, w2080, w2081, w2082, w2083, w2084, w2085, w2086, w2087, w2088, w2089, w2090, w2091, w2092, w2093, w2094, w2095, w2096, w2097, w2098, w2099, w2100, w2101, w2102, w2103, w2104, w2105, w2106, w2107, w2108, w2109, w2110, w2111, w2112, w2113, w2114, w2115, w2116, w2117, w2118, w2119, w2120, w2121, w2122, w2123, w2124, w2125, w2126, w2127, w2128, w2129, w2130, w2131, w2132, w2133, w2134, w2135, w2136, w2137, w2138, w2139, w2140, w2141, w2142, w2143, w2144, w2145, w2146, w2147, w2148, w2149, w2150, w2151, w2152, w2153, w2154, w2155, w2156, w2157, w2158, w2159, w2160, w2161, w2162, w2163, w2164, w2165, w2166, w2167, w2168, w2169, w2170, w2171, w2172, w2173, w2174, w2175, w2176, w2177, w2178, w2179, w2180, w2181, w2182, w2183, w2184, w2185, w2186, w2187, w2188, w2189, w2190, w2191, w2192, w2193, w2194, w2195, w2196, w2197, w2198, w2199, w2200, w2201, w2202, w2203, w2204, w2205, w2206, w2207, w2208, w2209, w2210, w2211, w2212, w2213, w2214, w2215, w2216, w2217, w2218, w2219, w2220, w2221, w2222, w2223, w2224, w2225, w2226, w2227, w2228, w2229, w2230, w2231, w2232, w2233, w2234, w2235, w2236, w2237, w2238, w2239, w2240, w2241, w2242, w2243, w2244, w2245, w2246, w2247, w2248, w2249, w2250, w2251, w2252, w2253, w2254, w2255, w2256, w2257, w2258, w2259, w2260, w2261, w2262, w2263, w2264, w2265, w2266, w2267, w2268, w2269, w2270, w2271, w2272, w2273, w2274, w2275, w2276, w2277, w2278, w2279, w2280, w2281, w2282, w2283, w2284, w2285, w2286, w2287, w2288, w2289, w2290, w2291, w2292, w2293, w2294, w2295, w2296, w2297, w2298, w2299, w2300, w2301, w2302, w2303, w2304, w2305, w2306, w2307, w2308, w2309, w2310, w2311, w2312, w2313, w2314, w2315, w2316, w2317, w2318, w2319, w2320, w2321, w2322, w2323, w2324, w2325, w2326, w2327, w2328, w2329, w2330, w2331, w2332, w2333, w2334, w2335, w2336, w2337, w2338, w2339, w2340, w2341, w2342, w2343, w2344, w2345, w2346, w2347, w2348, w2349, w2350, w2351, w2352, w2353, w2354, w2355, w2356, w2357, w2358, w2359, w2360, w2361, w2362, w2363, w2364, w2365, w2366, w2367, w2368, w2369, w2370, w2371, w2372, w2373, w2374, w2375, w2376, w2377, w2378, w2379, w2380, w2381, w2382, w2383, w2384, w2385, w2386, w2387, w2388, w2389, w2390, w2391, w2392, w2393, w2394, w2395, w2396, w2397, w2398, w2399, w2400, w2401, w2402, w2403, w2404, w2405, w2406, w2407, w2408, w2409, w2410, w2411, w2412, w2413, w2414, w2415, w2416, w2417, w2418, w2419, w2420, w2421, w2422, w2423, w2424, w2425, w2426, w2427, w2428, w2429, w2430, w2431, w2432, w2433, w2434, w2435, w2436, w2437, w2438, w2439, w2440, w2441, w2442, w2443, w2444, w2445, w2446, w2447, w2448, w2449, w2450, w2451, w2452, w2453, w2454, w2455, w2456, w2457, w2458, w2459, w2460, w2461, w2462, w2463, w2464, w2465, w2466, w2467, w2468, w2469, w2470, w2471, w2472, w2473, w2474, w2475, w2476, w2477, w2478, w2479, w2480, w2481, w2482, w2483, w2484, w2485, w2486, w2487, w2488, w2489, w2490, w2491, w2492, w2493, w2494, w2495, w2496, w2497, w2498, w2499, w2500, w2501, w2502, w2503, w2504, w2505, w2506, w2507, w2508, w2509, w2510, w2511, w2512, w2513, w2514, w2515, w2516, w2517, w2518, w2519, w2520, w2521, w2522, w2523, w2524, w2525, w2526, w2527, w2528, w2529, w2530, w2531, w2532, w2533, w2534, w2535, w2536, w2537, w2538, w2539, w2540, w2541, w2542, w2543, w2544, w2545, w2546, w2547, w2548, w2549, w2550, w2551, w2552, w2553, w2554, w2555, w2556, w2557, w2558, w2559, w2560, w2561, w2562, w2563, w2564, w2565, w2566, w2567, w2568, w2569, w2570, w2571, w2572, w2573, w2574, w2575, w2576, w2577, w2578, w2579, w2580, w2581, w2582, w2583, w2584, w2585, w2586, w2587, w2588, w2589, w2590, w2591, w2592, w2593, w2594, w2595, w2596, w2597, w2598, w2599, w2600, w2601, w2602, w2603, w2604, w2605, w2606, w2607, w2608, w2609, w2610, w2611, w2612, w2613, w2614, w2615, w2616, w2617, w2618, w2619, w2620, w2621, w2622, w2623, w2624, w2625, w2626, w2627, w2628, w2629, w2630, w2631, w2632, w2633, w2634, w2635, w2636, w2637, w2638, w2639, w2640, w2641, w2642, w2643, w2644, w2645, w2646, w2647, w2648, w2649, w2650, w2651, w2652, w2653, w2654, w2655, w2656, w2657, w2658, w2659, w2660, w2661, w2662, w2663, w2664, w2665, w2666, w2667, w2668, w2669, w2670, w2671, w2672, w2673, w2674, w2675, w2676, w2677, w2678, w2679, w2680, w2681, w2682, w2683, w2684, w2685, w2686, w2687, w2688, w2689, w2690, w2691, w2692, w2693, w2694, w2695, w2696, w2697, w2698, w2699, w2700, w2701, w2702, w2703, w2704, w2705, w2706, w2707, w2708, w2709, w2710, w2711, w2712, w2713, w2714, w2715, w2716, w2717, w2718, w2719, w2720, w2721, w2722, w2723, w2724, w2725, w2726, w2727, w2728, w2729, w2730, w2731, w2732, w2733, w2734, w2735, w2736, w2737, w2738, w2739, w2740, w2741, w2742, w2743, w2744, w2745, w2746, w2747, w2748, w2749, w2750, w2751, w2752, w2753, w2754, w2755, w2756, w2757, w2758, w2759, w2760, w2761, w2762, w2763, w2764, w2765, w2766, w2767, w2768, w2769, w2770, w2771, w2772, w2773, w2774, w2775, w2776, w2777, w2778, w2779, w2780, w2781, w2782, w2783, w2784, w2785, w2786, w2787, w2788, w2789, w2790, w2791, w2792, w2793, w2794, w2795, w2796, w2797, w2798, w2799, w2800, w2801, w2802, w2803, w2804, w2805, w2806, w2807, w2808, w2809, w2810, w2811, w2812, w2813, w2814, w2815, w2816, w2817, w2818, w2819, w2820, w2821, w2822, w2823, w2824, w2825, w2826, w2827, w2828, w2829, w2830, w2831, w2832, w2833, w2834, w2835, w2836, w2837, w2838, w2839, w2840, w2841, w2842, w2843, w2844, w2845, w2846, w2847, w2848, w2849, w2850, w2851, w2852, w2853, w2854, w2855, w2856, w2857, w2858, w2859, w2860, w2861, w2862, w2863, w2864, w2865, w2866, w2867, w2868, w2869, w2870, w2871, w2872, w2873, w2874, w2875, w2876, w2877, w2878, w2879, w2880, w2881, w2882, w2883, w2884, w2885, w2886, w2887, w2888, w2889, w2890, w2891, w2892, w2893, w2894, w2895, w2896, w2897, w2898, w2899, w2900, w2901, w2902, w2903, w2904, w2905, w2906, w2907, w2908, w2909, w2910, w2911, w2912, w2913, w2914, w2915, w2916, w2917, w2918, w2919, w2920, w2921, w2922, w2923, w2924, w2925, w2926, w2927, w2928, w2929, w2930, w2931, w2932, w2933, w2934, w2935, w2936, w2937, w2938, w2939, w2940, w2941, w2942, w2943, w2944, w2945, w2946, w2947, w2948, w2949, w2950, w2951, w2952, w2953, w2954, w2955, w2956, w2957, w2958, w2959, w2960, w2961, w2962, w2963, w2964, w2965, w2966, w2967, w2968, w2969, w2970, w2971, w2972, w2973, w2974, w2975, w2976, w2977, w2978, w2979, w2980, w2981, w2982, w2983, w2984, w2985, w2986, w2987, w2988, w2989, w2990, w2991, w2992, w2993, w2994, w2995, w2996, w2997, w2998, w2999, w3000, w3001, w3002, w3003, w3004, w3005, w3006, w3007, w3008, w3009, w3010, w3011, w3012, w3013, w3014, w3015, w3016, w3017, w3018, w3019, w3020, w3021, w3022, w3023, w3024, w3025, w3026, w3027, w3028, w3029, w3030, w3031, w3032, w3033, w3034, w3035, w3036, w3037, w3038, w3039, w3040, w3041, w3042, w3043, w3044, w3045, w3046, w3047, w3048, w3049, w3050, w3051, w3052, w3053, w3054, w3055, w3056, w3057, w3058, w3059, w3060, w3061, w3062, w3063, w3064, w3065, w3066, w3067, w3068, w3069, w3070, w3071, w3072, w3073, w3074, w3075, w3076, w3077, w3078, w3079, w3080, w3081, w3082, w3083, w3084, w3085, w3086, w3087, w3088, w3089, w3090, w3091, w3092, w3093, w3094, w3095, w3096, w3097, w3098, w3099, w3100, w3101, w3102, w3103, w3104, w3105, w3106, w3107, w3108, w3109, w3110, w3111, w3112, w3113, w3114, w3115, w3116, w3117, w3118, w3119, w3120, w3121, w3122, w3123, w3124, w3125, w3126, w3127, w3128, w3129, w3130, w3131, w3132, w3133, w3134, w3135, w3136, w3137, w3138, w3139, w3140, w3141, w3142, w3143, w3144, w3145, w3146, w3147, w3148, w3149, w3150, w3151, w3152, w3153, w3154, w3155, w3156, w3157, w3158, w3159, w3160, w3161, w3162, w3163, w3164, w3165, w3166, w3167, w3168, w3169, w3170, w3171, w3172, w3173, w3174, w3175, w3176, w3177, w3178, w3179, w3180, w3181, w3182, w3183, w3184, w3185, w3186, w3187, w3188, w3189, w3190, w3191, w3192, w3193, w3194, w3195, w3196, w3197, w3198, w3199, w3200, w3201, w3202, w3203, w3204, w3205, w3206, w3207, w3208, w3209, w3210, w3211, w3212, w3213, w3214, w3215, w3216, w3217, w3218, w3219, w3220, w3221, w3222, w3223, w3224, w3225, w3226, w3227, w3228, w3229, w3230, w3231, w3232, w3233, w3234, w3235, w3236, w3237, w3238, w3239, w3240, w3241, w3242, w3243, w3244, w3245, w3246, w3247, w3248, w3249, w3250, w3251, w3252, w3253, w3254, w3255, w3256, w3257, w3258, w3259, w3260, w3261, w3262, w3263, w3264, w3265, w3266, w3267, w3268, w3269, w3270, w3271, w3272, w3273, w3274, w3275, w3276, w3277, w3278, w3279, w3280, w3281, w3282, w3283, w3284, w3285, w3286, w3287, w3288, w3289, w3290, w3291, w3292, w3293, w3294, w3295, w3296, w3297, w3298, w3299, w3300, w3301, w3302, w3303, w3304, w3305, w3306, w3307, w3308, w3309, w3310, w3311, w3312, w3313, w3314, w3315, w3316, w3317, w3318, w3319, w3320, w3321, w3322, w3323, w3324, w3325, w3326, w3327, w3328, w3329, w3330, w3331, w3332, w3333, w3334, w3335, w3336, w3337, w3338, w3339, w3340, w3341, w3342, w3343, w3344, w3345, w3346, w3347, w3348, w3349, w3350, w3351, w3352, w3353, w3354, w3355, w3356, w3357, w3358, w3359, w3360, w3361, w3362, w3363, w3364, w3365, w3366, w3367, w3368, w3369, w3370, w3371, w3372, w3373, w3374, w3375, w3376, w3377, w3378, w3379, w3380, w3381, w3382, w3383, w3384, w3385, w3386, w3387, w3388, w3389, w3390, w3391, w3392, w3393, w3394, w3395, w3396, w3397, w3398, w3399, w3400, w3401, w3402, w3403, w3404, w3405, w3406, w3407, w3408, w3409, w3410, w3411, w3412, w3413, w3414, w3415, w3416, w3417, w3418, w3419, w3420, w3421, w3422, w3423, w3424, w3425, w3426, w3427, w3428, w3429, w3430, w3431, w3432, w3433, w3434, w3435, w3436, w3437, w3438, w3439, w3440, w3441, w3442, w3443, w3444, w3445, w3446, w3447, w3448, w3449, w3450, w3451, w3452, w3453, w3454, w3455, w3456, w3457, w3458, w3459, w3460, w3461, w3462, w3463, w3464, w3465, w3466, w3467, w3468, w3469, w3470, w3471, w3472, w3473, w3474, w3475, w3476, w3477, w3478, w3479, w3480, w3481, w3482, w3483, w3484, w3485, w3486, w3487, w3488, w3489, w3490, w3491, w3492, w3493, w3494, w3495, w3496, w3497, w3498, w3499, w3500, w3501, w3502, w3503, w3504, w3505, w3506, w3507, w3508, w3509, w3510, w3511, w3512, w3513, w3514, w3515, w3516, w3517, w3518, w3519, w3520, w3521, w3522, w3523, w3524, w3525, w3526, w3527, w3528, w3529, w3530, w3531, w3532, w3533, w3534, w3535, w3536, w3537, w3538, w3539, w3540, w3541, w3542, w3543, w3544, w3545, w3546, w3547, w3548, w3549, w3550, w3551, w3552, w3553, w3554, w3555, w3556, w3557, w3558, w3559, w3560, w3561, w3562, w3563, w3564, w3565, w3566, w3567, w3568, w3569, w3570, w3571, w3572, w3573, w3574, w3575, w3576, w3577, w3578, w3579, w3580, w3581, w3582, w3583, w3584, w3585, w3586, w3587, w3588, w3589, w3590, w3591, w3592, w3593, w3594, w3595, w3596, w3597, w3598, w3599, w3600, w3601, w3602, w3603, w3604, w3605, w3606, w3607, w3608, w3609, w3610, w3611, w3612, w3613, w3614, w3615, w3616, w3617, w3618, w3619, w3620, w3621, w3622, w3623, w3624, w3625, w3626, w3627, w3628, w3629, w3630, w3631, w3632, w3633, w3634, w3635, w3636, w3637, w3638, w3639, w3640, w3641, w3642, w3643, w3644, w3645, w3646, w3647, w3648, w3649, w3650, w3651, w3652, w3653, w3654, w3655, w3656, w3657, w3658, w3659, w3660, w3661, w3662, w3663, w3664, w3665, w3666, w3667, w3668, w3669, w3670, w3671, w3672, w3673, w3674, w3675, w3676, w3677, w3678, w3679, w3680, w3681, w3682, w3683, w3684, w3685, w3686, w3687, w3688, w3689, w3690, w3691, w3692, w3693, w3694, w3695, w3696, w3697, w3698, w3699, w3700, w3701, w3702, w3703, w3704, w3705, w3706, w3707, w3708, w3709, w3710, w3711, w3712, w3713, w3714, w3715, w3716, w3717, w3718, w3719, w3720, w3721, w3722, w3723, w3724, w3725, w3726, w3727, w3728, w3729, w3730, w3731, w3732, w3733, w3734, w3735, w3736, w3737, w3738, w3739, w3740, w3741, w3742, w3743, w3744, w3745, w3746, w3747, w3748, w3749, w3750, w3751, w3752, w3753, w3754, w3755, w3756, w3757, w3758, w3759, w3760, w3761, w3762, w3763, w3764, w3765, w3766, w3767, w3768, w3769, w3770, w3771, w3772, w3773, w3774, w3775, w3776, w3777, w3778, w3779, w3780, w3781, w3782, w3783, w3784, w3785, w3786, w3787, w3788, w3789, w3790, w3791, w3792, w3793, w3794, w3795, w3796, w3797, w3798, w3799, w3800, w3801, w3802, w3803, w3804, w3805, w3806, w3807, w3808, w3809, w3810, w3811, w3812, w3813, w3814, w3815, w3816, w3817, w3818, w3819, w3820, w3821, w3822, w3823, w3824, w3825, w3826, w3827, w3828, w3829, w3830, w3831, w3832, w3833, w3834, w3835, w3836, w3837, w3838, w3839, w3840, w3841, w3842, w3843, w3844, w3845, w3846, w3847, w3848, w3849, w3850, w3851, w3852, w3853, w3854, w3855, w3856, w3857, w3858, w3859, w3860, w3861, w3862, w3863, w3864, w3865, w3866, w3867, w3868, w3869, w3870, w3871, w3872, w3873, w3874, w3875, w3876, w3877, w3878, w3879, w3880, w3881, w3882, w3883, w3884, w3885, w3886, w3887, w3888, w3889, w3890, w3891, w3892, w3893, w3894, w3895, w3896, w3897, w3898, w3899, w3900, w3901, w3902, w3903, w3904, w3905, w3906, w3907, w3908, w3909, w3910, w3911, w3912, w3913, w3914, w3915, w3916, w3917, w3918, w3919, w3920, w3921, w3922, w3923, w3924, w3925, w3926, w3927, w3928, w3929, w3930, w3931, w3932, w3933, w3934, w3935, w3936, w3937, w3938, w3939, w3940, w3941, w3942, w3943, w3944, w3945, w3946, w3947, w3948, w3949, w3950, w3951, w3952, w3953, w3954, w3955, w3956, w3957, w3958, w3959, w3960, w3961, w3962, w3963, w3964, w3965, w3966, w3967, w3968, w3969, w3970, w3971, w3972, w3973, w3974, w3975, w3976, w3977, w3978, w3979, w3980, w3981, w3982, w3983, w3984, w3985, w3986, w3987, w3988, w3989, w3990, w3991, w3992, w3993, w3994, w3995, w3996, w3997, w3998, w3999, w4000, w4001, w4002, w4003, w4004, w4005, w4006, w4007, w4008, w4009, w4010, w4011, w4012, w4013, w4014, w4015, w4016, w4017, w4018, w4019, w4020, w4021, w4022, w4023, w4024, w4025, w4026, w4027, w4028, w4029, w4030, w4031, w4032, w4033, w4034, w4035, w4036, w4037, w4038, w4039, w4040, w4041, w4042, w4043, w4044, w4045, w4046, w4047, w4048, w4049, w4050, w4051, w4052, w4053, w4054, w4055, w4056, w4057, w4058, w4059, w4060, w4061, w4062, w4063, w4064, w4065, w4066, w4067, w4068, w4069, w4070, w4071, w4072, w4073, w4074, w4075, w4076, w4077, w4078, w4079, w4080, w4081, w4082, w4083, w4084, w4085, w4086, w4087, w4088, w4089, w4090, w4091, w4092, w4093, w4094, w4095, w4096, w4097, w4098, w4099, w4100, w4101, w4102, w4103, w4104, w4105, w4106, w4107, w4108, w4109, w4110, w4111, w4112, w4113, w4114, w4115, w4116, w4117, w4118, w4119, w4120, w4121, w4122, w4123, w4124, w4125, w4126, w4127, w4128, w4129, w4130, w4131, w4132, w4133, w4134, w4135, w4136, w4137, w4138, w4139, w4140, w4141, w4142, w4143, w4144, w4145, w4146, w4147, w4148, w4149, w4150, w4151, w4152, w4153, w4154, w4155, w4156, w4157, w4158, w4159, w4160, w4161, w4162, w4163, w4164, w4165, w4166, w4167, w4168, w4169, w4170, w4171, w4172, w4173, w4174, w4175, w4176, w4177, w4178, w4179, w4180, w4181, w4182, w4183, w4184, w4185, w4186, w4187, w4188, w4189, w4190, w4191, w4192, w4193, w4194, w4195, w4196, w4197, w4198, w4199, w4200, w4201, w4202, w4203, w4204, w4205, w4206, w4207, w4208, w4209, w4210, w4211, w4212, w4213, w4214, w4215, w4216, w4217, w4218, w4219, w4220, w4221, w4222, w4223, w4224, w4225, w4226, w4227, w4228, w4229, w4230, w4231, w4232, w4233, w4234, w4235, w4236, w4237, w4238, w4239, w4240, w4241, w4242, w4243, w4244, w4245, w4246, w4247, w4248, w4249, w4250, w4251, w4252, w4253, w4254, w4255, w4256, w4257, w4258, w4259, w4260, w4261, w4262, w4263, w4264, w4265, w4266, w4267, w4268, w4269, w4270, w4271, w4272, w4273, w4274, w4275, w4276, w4277, w4278, w4279, w4280, w4281, w4282, w4283, w4284, w4285, w4286, w4287, w4288, w4289, w4290, w4291, w4292, w4293, w4294, w4295, w4296, w4297, w4298, w4299, w4300, w4301, w4302, w4303, w4304, w4305, w4306, w4307, w4308, w4309, w4310, w4311, w4312, w4313, w4314, w4315, w4316, w4317, w4318, w4319, w4320, w4321, w4322, w4323, w4324, w4325, w4326, w4327, w4328, w4329, w4330, w4331, w4332, w4333, w4334, w4335, w4336, w4337, w4338, w4339, w4340, w4341, w4342, w4343, w4344, w4345, w4346, w4347, w4348, w4349, w4350, w4351, w4352, w4353, w4354, w4355, w4356, w4357, w4358, w4359, w4360, w4361, w4362, w4363, w4364, w4365, w4366, w4367, w4368, w4369, w4370, w4371, w4372, w4373, w4374, w4375, w4376, w4377, w4378, w4379, w4380, w4381, w4382, w4383, w4384, w4385, w4386, w4387, w4388, w4389, w4390, w4391, w4392, w4393, w4394, w4395, w4396, w4397, w4398, w4399, w4400, w4401, w4402, w4403, w4404, w4405, w4406, w4407, w4408, w4409, w4410, w4411, w4412, w4413, w4414, w4415, w4416, w4417, w4418, w4419, w4420, w4421, w4422, w4423, w4424, w4425, w4426, w4427, w4428, w4429, w4430, w4431, w4432, w4433, w4434, w4435, w4436, w4437, w4438, w4439, w4440, w4441, w4442, w4443, w4444, w4445, w4446, w4447, w4448, w4449, w4450, w4451, w4452, w4453, w4454, w4455, w4456, w4457, w4458, w4459, w4460, w4461, w4462, w4463, w4464, w4465, w4466, w4467, w4468, w4469, w4470, w4471, w4472, w4473, w4474, w4475, w4476, w4477, w4478, w4479, w4480, w4481, w4482, w4483, w4484, w4485, w4486, w4487, w4488, w4489, w4490, w4491, w4492, w4493, w4494, w4495, w4496, w4497, w4498, w4499, w4500, w4501, w4502, w4503, w4504, w4505, w4506, w4507, w4508, w4509, w4510, w4511, w4512, w4513, w4514, w4515, w4516, w4517, w4518, w4519, w4520, w4521, w4522, w4523, w4524, w4525, w4526, w4527, w4528, w4529, w4530, w4531, w4532, w4533, w4534, w4535, w4536, w4537, w4538, w4539, w4540, w4541, w4542, w4543, w4544, w4545, w4546, w4547, w4548, w4549, w4550, w4551, w4552, w4553, w4554, w4555, w4556, w4557, w4558, w4559, w4560, w4561, w4562, w4563, w4564, w4565, w4566, w4567, w4568, w4569, w4570, w4571, w4572, w4573, w4574, w4575, w4576, w4577, w4578, w4579, w4580, w4581, w4582, w4583, w4584, w4585, w4586, w4587, w4588, w4589, w4590, w4591, w4592, w4593, w4594, w4595, w4596, w4597, w4598, w4599, w4600, w4601, w4602, w4603, w4604, w4605, w4606, w4607, w4608, w4609, w4610, w4611, w4612, w4613, w4614, w4615, w4616, w4617, w4618, w4619, w4620, w4621, w4622, w4623, w4624, w4625, w4626, w4627, w4628, w4629, w4630, w4631, w4632, w4633, w4634, w4635, w4636, w4637, w4638, w4639, w4640, w4641, w4642, w4643, w4644, w4645, w4646, w4647, w4648, w4649, w4650, w4651, w4652, w4653, w4654, w4655, w4656, w4657, w4658, w4659, w4660, w4661, w4662, w4663, w4664, w4665, w4666, w4667, w4668, w4669, w4670, w4671, w4672, w4673, w4674, w4675, w4676, w4677, w4678, w4679, w4680, w4681, w4682, w4683, w4684, w4685, w4686, w4687, w4688, w4689, w4690, w4691, w4692, w4693, w4694, w4695, w4696, w4697, w4698, w4699, w4700, w4701, w4702, w4703, w4704, w4705, w4706, w4707, w4708, w4709, w4710, w4711, w4712, w4713, w4714, w4715, w4716, w4717, w4718, w4719, w4720, w4721, w4722, w4723, w4724, w4725, w4726, w4727, w4728, w4729, w4730, w4731, w4732, w4733, w4734, w4735, w4736, w4737, w4738, w4739, w4740, w4741, w4742, w4743, w4744, w4745, w4746, w4747, w4748, w4749, w4750, w4751, w4752, w4753, w4754, w4755, w4756, w4757, w4758, w4759, w4760, w4761, w4762, w4763, w4764, w4765, w4766, w4767, w4768, w4769, w4770, w4771, w4772, w4773, w4774, w4775, w4776, w4777, w4778, w4779, w4780, w4781, w4782, w4783, w4784, w4785, w4786, w4787, w4788, w4789, w4790, w4791, w4792, w4793, w4794, w4795, w4796, w4797, w4798, w4799, w4800, w4801, w4802, w4803, w4804, w4805, w4806, w4807, w4808, w4809, w4810, w4811, w4812, w4813, w4814, w4815, w4816, w4817, w4818, w4819, w4820, w4821, w4822, w4823, w4824, w4825, w4826, w4827, w4828, w4829, w4830, w4831, w4832, w4833, w4834, w4835, w4836, w4837, w4838, w4839, w4840, w4841, w4842, w4843, w4844, w4845, w4846, w4847, w4848, w4849, w4850, w4851, w4852, w4853, w4854, w4855, w4856, w4857, w4858, w4859, w4860, w4861, w4862, w4863, w4864, w4865, w4866, w4867, w4868, w4869, w4870, w4871, w4872, w4873, w4874, w4875, w4876, w4877, w4878, w4879, w4880, w4881, w4882, w4883, w4884, w4885, w4886, w4887, w4888, w4889, w4890, w4891, w4892, w4893, w4894, w4895, w4896, w4897, w4898, w4899, w4900, w4901, w4902, w4903, w4904, w4905, w4906, w4907, w4908, w4909, w4910, w4911, w4912, w4913, w4914, w4915, w4916, w4917, w4918, w4919, w4920, w4921, w4922, w4923, w4924, w4925, w4926, w4927, w4928, w4929, w4930, w4931, w4932, w4933, w4934, w4935, w4936, w4937, w4938, w4939, w4940, w4941, w4942, w4943, w4944, w4945, w4946, w4947, w4948, w4949, w4950, w4951, w4952, w4953, w4954, w4955, w4956, w4957, w4958, w4959, w4960, w4961, w4962, w4963, w4964, w4965, w4966, w4967, w4968, w4969, w4970, w4971, w4972, w4973, w4974, w4975, w4976, w4977, w4978, w4979, w4980, w4981, w4982, w4983, w4984, w4985, w4986, w4987, w4988, w4989, w4990, w4991, w4992, w4993, w4994, w4995, w4996, w4997, w4998, w4999, w5000, w5001, w5002, w5003, w5004, w5005, w5006, w5007, w5008, w5009, w5010, w5011, w5012, w5013, w5014, w5015, w5016, w5017, w5018, w5019, w5020, w5021, w5022, w5023, w5024, w5025, w5026, w5027, w5028, w5029, w5030, w5031, w5032, w5033, w5034, w5035, w5036, w5037, w5038, w5039, w5040, w5041, w5042, w5043, w5044, w5045, w5046, w5047, w5048, w5049, w5050, w5051, w5052, w5053, w5054, w5055, w5056, w5057, w5058, w5059, w5060, w5061, w5062, w5063, w5064, w5065, w5066, w5067, w5068, w5069, w5070, w5071, w5072, w5073, w5074, w5075, w5076, w5077, w5078, w5079, w5080, w5081, w5082, w5083, w5084, w5085, w5086, w5087, w5088, w5089, w5090, w5091, w5092, w5093, w5094, w5095, w5096, w5097, w5098, w5099, w5100, w5101, w5102, w5103, w5104, w5105, w5106, w5107, w5108, w5109, w5110, w5111, w5112, w5113, w5114, w5115, w5116, w5117, w5118, w5119, w5120, w5121, w5122, w5123, w5124, w5125, w5126, w5127, w5128, w5129, w5130, w5131, w5132, w5133, w5134, w5135, w5136, w5137, w5138, w5139, w5140, w5141, w5142, w5143, w5144, w5145, w5146, w5147, w5148, w5149, w5150, w5151, w5152, w5153, w5154, w5155, w5156, w5157, w5158, w5159, w5160, w5161, w5162, w5163, w5164, w5165, w5166, w5167, w5168, w5169, w5170, w5171, w5172, w5173, w5174, w5175, w5176, w5177, w5178, w5179, w5180, w5181, w5182, w5183, w5184, w5185, w5186, w5187, w5188, w5189, w5190, w5191, w5192, w5193, w5194, w5195, w5196, w5197, w5198, w5199, w5200, w5201, w5202, w5203, w5204, w5205, w5206, w5207, w5208, w5209, w5210, w5211, w5212, w5213, w5214, w5215, w5216, w5217, w5218, w5219, w5220, w5221, w5222, w5223, w5224, w5225, w5226, w5227, w5228, w5229, w5230, w5231, w5232, w5233, w5234, w5235, w5236, w5237, w5238, w5239, w5240, w5241, w5242, w5243, w5244, w5245, w5246, w5247, w5248, w5249, w5250, w5251, w5252, w5253, w5254, w5255, w5256, w5257, w5258, w5259, w5260, w5261, w5262, w5263, w5264, w5265, w5266, w5267, w5268, w5269, w5270, w5271, w5272, w5273, w5274, w5275, w5276, w5277, w5278, w5279, w5280, w5281, w5282, w5283, w5284, w5285, w5286, w5287, w5288, w5289, w5290, w5291, w5292, w5293, w5294, w5295, w5296, w5297, w5298, w5299, w5300, w5301, w5302, w5303, w5304, w5305, w5306, w5307, w5308, w5309, w5310, w5311, w5312, w5313, w5314, w5315, w5316, w5317, w5318, w5319, w5320, w5321, w5322, w5323, w5324, w5325, w5326, w5327, w5328, w5329, w5330, w5331, w5332, w5333, w5334, w5335, w5336, w5337, w5338, w5339, w5340, w5341, w5342, w5343, w5344, w5345, w5346, w5347, w5348, w5349, w5350, w5351, w5352, w5353, w5354, w5355, w5356, w5357, w5358, w5359, w5360, w5361, w5362, w5363, w5364, w5365, w5366, w5367, w5368, w5369, w5370, w5371, w5372, w5373, w5374, w5375, w5376, w5377, w5378, w5379, w5380, w5381, w5382, w5383, w5384, w5385, w5386, w5387, w5388, w5389, w5390, w5391, w5392, w5393, w5394, w5395, w5396, w5397, w5398, w5399, w5400, w5401, w5402, w5403, w5404, w5405, w5406, w5407, w5408, w5409, w5410, w5411, w5412, w5413, w5414, w5415, w5416, w5417, w5418, w5419, w5420, w5421, w5422, w5423, w5424, w5425, w5426, w5427, w5428, w5429, w5430, w5431, w5432, w5433, w5434, w5435, w5436, w5437, w5438, w5439, w5440, w5441, w5442, w5443, w5444, w5445, w5446, w5447, w5448, w5449, w5450, w5451, w5452, w5453, w5454, w5455, w5456, w5457, w5458, w5459, w5460, w5461, w5462, w5463, w5464, w5465, w5466, w5467, w5468, w5469, w5470, w5471, w5472, w5473, w5474, w5475, w5476, w5477, w5478, w5479, w5480, w5481, w5482, w5483, w5484, w5485, w5486, w5487, w5488, w5489, w5490, w5491, w5492, w5493, w5494, w5495, w5496, w5497, w5498, w5499, w5500, w5501, w5502, w5503, w5504, w5505, w5506, w5507, w5508, w5509, w5510, w5511, w5512, w5513, w5514, w5515, w5516, w5517, w5518, w5519, w5520, w5521, w5522, w5523, w5524, w5525, w5526, w5527, w5528, w5529, w5530, w5531, w5532, w5533, w5534, w5535, w5536, w5537, w5538, w5539, w5540, w5541, w5542, w5543, w5544, w5545, w5546, w5547, w5548, w5549, w5550, w5551, w5552, w5553, w5554, w5555, w5556, w5557, w5558, w5559, w5560, w5561, w5562, w5563, w5564, w5565, w5566, w5567, w5568, w5569, w5570, w5571, w5572, w5573, w5574, w5575, w5576, w5577, w5578, w5579, w5580, w5581, w5582, w5583, w5584, w5585, w5586, w5587, w5588, w5589, w5590, w5591, w5592, w5593, w5594, w5595, w5596, w5597, w5598, w5599, w5600, w5601, w5602, w5603, w5604, w5605, w5606, w5607, w5608, w5609, w5610, w5611, w5612, w5613, w5614, w5615, w5616, w5617, w5618, w5619, w5620, w5621, w5622, w5623, w5624, w5625, w5626, w5627, w5628, w5629, w5630, w5631, w5632, w5633, w5634, w5635, w5636, w5637, w5638, w5639, w5640, w5641, w5642, w5643, w5644, w5645, w5646, w5647, w5648, w5649, w5650, w5651, w5652, w5653, w5654, w5655, w5656, w5657, w5658, w5659, w5660, w5661, w5662, w5663, w5664, w5665, w5666, w5667, w5668, w5669, w5670, w5671, w5672, w5673, w5674, w5675, w5676, w5677, w5678, w5679, w5680, w5681, w5682, w5683, w5684, w5685, w5686, w5687, w5688, w5689, w5690, w5691, w5692, w5693, w5694, w5695, w5696, w5697, w5698, w5699, w5700, w5701, w5702, w5703, w5704, w5705, w5706, w5707, w5708, w5709, w5710, w5711, w5712, w5713, w5714, w5715, w5716, w5717, w5718, w5719, w5720, w5721, w5722, w5723, w5724, w5725, w5726, w5727, w5728, w5729, w5730, w5731, w5732, w5733, w5734, w5735, w5736, w5737, w5738, w5739, w5740, w5741, w5742, w5743, w5744, w5745, w5746, w5747, w5748, w5749, w5750, w5751, w5752, w5753, w5754, w5755, w5756, w5757, w5758, w5759, w5760, w5761, w5762, w5763, w5764, w5765, w5766, w5767, w5768, w5769, w5770, w5771, w5772, w5773, w5774, w5775, w5776, w5777, w5778, w5779, w5780, w5781, w5782, w5783, w5784, w5785, w5786, w5787, w5788, w5789, w5790, w5791, w5792, w5793, w5794, w5795, w5796, w5797, w5798, w5799, w5800, w5801, w5802, w5803, w5804, w5805, w5806, w5807, w5808, w5809, w5810, w5811, w5812, w5813, w5814, w5815, w5816, w5817, w5818, w5819, w5820, w5821, w5822, w5823, w5824, w5825, w5826, w5827, w5828, w5829, w5830, w5831, w5832, w5833, w5834, w5835, w5836, w5837, w5838, w5839, w5840, w5841, w5842, w5843, w5844, w5845, w5846, w5847, w5848, w5849, w5850, w5851, w5852, w5853, w5854, w5855, w5856, w5857, w5858, w5859, w5860, w5861, w5862, w5863, w5864, w5865, w5866, w5867, w5868, w5869, w5870, w5871, w5872, w5873, w5874, w5875, w5876, w5877, w5878, w5879, w5880, w5881, w5882, w5883, w5884, w5885, w5886, w5887, w5888, w5889, w5890, w5891, w5892, w5893, w5894, w5895, w5896, w5897, w5898, w5899, w5900, w5901, w5902, w5903, w5904, w5905, w5906, w5907, w5908, w5909, w5910, w5911, w5912, w5913, w5914, w5915, w5916, w5917, w5918, w5919, w5920, w5921, w5922, w5923, w5924, w5925, w5926, w5927, w5928, w5929, w5930, w5931, w5932, w5933, w5934, w5935, w5936, w5937, w5938, w5939, w5940, w5941, w5942, w5943, w5944, w5945, w5946, w5947, w5948, w5949, w5950, w5951, w5952, w5953, w5954, w5955, w5956, w5957, w5958, w5959, w5960, w5961, w5962, w5963, w5964, w5965, w5966, w5967, w5968, w5969, w5970, w5971, w5972, w5973, w5974, w5975, w5976, w5977, w5978, w5979, w5980, w5981, w5982, w5983, w5984, w5985, w5986, w5987, w5988, w5989, w5990, w5991, w5992, w5993, w5994, w5995, w5996, w5997, w5998, w5999, w6000, w6001, w6002, w6003, w6004, w6005, w6006, w6007, w6008, w6009, w6010, w6011, w6012, w6013, w6014, w6015, w6016, w6017, w6018, w6019, w6020, w6021, w6022, w6023, w6024, w6025, w6026, w6027, w6028, w6029, w6030, w6031, w6032, w6033, w6034, w6035, w6036, w6037, w6038, w6039, w6040, w6041, w6042, w6043, w6044, w6045, w6046, w6047, w6048, w6049, w6050, w6051, w6052, w6053, w6054, w6055, w6056, w6057, w6058, w6059, w6060, w6061, w6062, w6063, w6064, w6065, w6066, w6067, w6068, w6069, w6070, w6071, w6072, w6073, w6074, w6075, w6076, w6077, w6078, w6079, w6080, w6081, w6082, w6083, w6084, w6085, w6086, w6087, w6088, w6089, w6090, w6091, w6092, w6093, w6094, w6095, w6096, w6097, w6098, w6099, w6100, w6101, w6102, w6103, w6104, w6105, w6106, w6107, w6108, w6109, w6110, w6111, w6112, w6113, w6114, w6115, w6116, w6117, w6118, w6119, w6120, w6121, w6122, w6123, w6124, w6125, w6126, w6127, w6128, w6129, w6130, w6131, w6132, w6133, w6134, w6135, w6136, w6137, w6138, w6139, w6140, w6141, w6142, w6143, w6144, w6145, w6146, w6147, w6148, w6149, w6150, w6151, w6152, w6153, w6154, w6155, w6156, w6157, w6158, w6159, w6160, w6161, w6162, w6163, w6164, w6165, w6166, w6167, w6168, w6169, w6170, w6171, w6172, w6173, w6174, w6175, w6176, w6177, w6178, w6179, w6180, w6181, w6182, w6183, w6184, w6185, w6186, w6187, w6188, w6189, w6190, w6191, w6192, w6193, w6194, w6195, w6196, w6197, w6198, w6199, w6200, w6201, w6202, w6203, w6204, w6205, w6206, w6207, w6208, w6209, w6210, w6211, w6212, w6213, w6214, w6215, w6216, w6217, w6218, w6219, w6220, w6221, w6222, w6223, w6224, w6225, w6226, w6227, w6228, w6229, w6230, w6231, w6232, w6233, w6234, w6235, w6236, w6237, w6238, w6239, w6240, w6241, w6242, w6243, w6244, w6245, w6246, w6247, w6248, w6249, w6250, w6251, w6252, w6253, w6254, w6255, w6256, w6257, w6258, w6259, w6260, w6261, w6262, w6263, w6264, w6265, w6266, w6267, w6268, w6269, w6270, w6271, w6272, w6273, w6274, w6275, w6276, w6277, w6278, w6279, w6280, w6281, w6282, w6283, w6284, w6285, w6286, w6287, w6288, w6289, w6290, w6291, w6292, w6293, w6294, w6295, w6296, w6297, w6298, w6299, w6300, w6301, w6302, w6303, w6304, w6305, w6306, w6307, w6308, w6309, w6310, w6311, w6312, w6313, w6314, w6315, w6316, w6317, w6318, w6319, w6320, w6321, w6322, w6323, w6324, w6325, w6326, w6327, w6328, w6329, w6330, w6331, w6332, w6333, w6334, w6335, w6336, w6337, w6338, w6339, w6340, w6341, w6342, w6343, w6344, w6345, w6346, w6347, w6348, w6349, w6350, w6351, w6352, w6353, w6354, w6355, w6356, w6357, w6358, w6359, w6360, w6361, w6362, w6363, w6364, w6365, w6366, w6367, w6368, w6369, w6370, w6371, w6372, w6373, w6374, w6375, w6376, w6377, w6378, w6379, w6380, w6381, w6382, w6383, w6384, w6385, w6386, w6387, w6388, w6389, w6390, w6391, w6392, w6393, w6394, w6395, w6396, w6397, w6398, w6399, w6400, w6401, w6402, w6403, w6404, w6405, w6406, w6407, w6408, w6409, w6410, w6411, w6412, w6413, w6414, w6415, w6416, w6417, w6418, w6419, w6420, w6421, w6422, w6423, w6424, w6425, w6426, w6427, w6428, w6429, w6430, w6431, w6432, w6433, w6434, w6435, w6436, w6437, w6438, w6439, w6440, w6441, w6442, w6443, w6444, w6445, w6446, w6447, w6448, w6449, w6450, w6451, w6452, w6453, w6454, w6455, w6456, w6457, w6458, w6459, w6460, w6461, w6462, w6463, w6464, w6465, w6466, w6467, w6468, w6469, w6470, w6471, w6472, w6473, w6474, w6475, w6476, w6477, w6478, w6479, w6480, w6481, w6482, w6483, w6484, w6485, w6486, w6487, w6488, w6489, w6490, w6491, w6492, w6493, w6494, w6495, w6496, w6497, w6498, w6499, w6500, w6501, w6502, w6503, w6504, w6505, w6506, w6507, w6508, w6509, w6510, w6511, w6512, w6513, w6514, w6515, w6516, w6517, w6518, w6519, w6520, w6521, w6522, w6523, w6524, w6525, w6526, w6527, w6528, w6529, w6530, w6531, w6532, w6533, w6534, w6535, w6536, w6537, w6538, w6539, w6540, w6541, w6542, w6543, w6544, w6545, w6546, w6547, w6548, w6549, w6550, w6551, w6552, w6553, w6554, w6555, w6556, w6557, w6558, w6559, w6560, w6561, w6562, w6563, w6564, w6565, w6566, w6567, w6568, w6569, w6570, w6571, w6572, w6573, w6574, w6575, w6576, w6577, w6578, w6579, w6580, w6581, w6582, w6583, w6584, w6585, w6586, w6587, w6588, w6589, w6590, w6591, w6592, w6593, w6594, w6595, w6596, w6597, w6598, w6599, w6600, w6601, w6602, w6603, w6604, w6605, w6606, w6607, w6608, w6609, w6610, w6611, w6612, w6613, w6614, w6615, w6616, w6617, w6618, w6619, w6620, w6621, w6622, w6623, w6624, w6625, w6626, w6627, w6628, w6629, w6630, w6631, w6632, w6633, w6634, w6635, w6636, w6637, w6638, w6639, w6640, w6641, w6642, w6643, w6644, w6645, w6646, w6647, w6648, w6649, w6650, w6651, w6652, w6653, w6654, w6655, w6656, w6657, w6658, w6659, w6660, w6661, w6662, w6663, w6664, w6665, w6666, w6667, w6668, w6669, w6670, w6671, w6672, w6673, w6674, w6675, w6676, w6677, w6678, w6679, w6680, w6681, w6682, w6683, w6684, w6685, w6686, w6687, w6688, w6689, w6690, w6691, w6692, w6693, w6694, w6695, w6696, w6697, w6698, w6699, w6700, w6701, w6702, w6703, w6704, w6705, w6706, w6707, w6708, w6709, w6710, w6711, w6712, w6713, w6714, w6715, w6716, w6717, w6718, w6719, w6720, w6721, w6722, w6723, w6724, w6725, w6726, w6727, w6728, w6729, w6730, w6731, w6732, w6733, w6734, w6735, w6736, w6737, w6738, w6739, w6740, w6741, w6742, w6743, w6744, w6745, w6746, w6747, w6748, w6749, w6750, w6751, w6752, w6753, w6754, w6755, w6756, w6757, w6758, w6759, w6760, w6761, w6762, w6763, w6764, w6765, w6766, w6767, w6768, w6769, w6770, w6771, w6772, w6773, w6774, w6775, w6776, w6777, w6778, w6779, w6780, w6781, w6782, w6783, w6784, w6785, w6786, w6787, w6788, w6789, w6790, w6791, w6792, w6793, w6794, w6795, w6796, w6797, w6798, w6799, w6800, w6801, w6802, w6803, w6804, w6805, w6806, w6807, w6808, w6809, w6810, w6811, w6812, w6813, w6814, w6815, w6816, w6817, w6818, w6819, w6820, w6821, w6822, w6823, w6824, w6825, w6826, w6827, w6828, w6829, w6830, w6831, w6832, w6833, w6834, w6835, w6836, w6837, w6838, w6839, w6840, w6841, w6842, w6843, w6844, w6845, w6846, w6847, w6848, w6849, w6850, w6851, w6852, w6853, w6854, w6855, w6856, w6857, w6858, w6859, w6860, w6861, w6862, w6863, w6864, w6865, w6866, w6867, w6868, w6869, w6870, w6871, w6872, w6873, w6874, w6875, w6876, w6877, w6878, w6879, w6880, w6881, w6882, w6883, w6884, w6885, w6886, w6887, w6888, w6889, w6890, w6891, w6892, w6893, w6894, w6895, w6896, w6897, w6898, w6899, w6900, w6901, w6902, w6903, w6904, w6905, w6906, w6907, w6908, w6909, w6910, w6911, w6912, w6913, w6914, w6915, w6916, w6917, w6918, w6919, w6920, w6921, w6922, w6923, w6924, w6925, w6926, w6927, w6928, w6929, w6930, w6931, w6932, w6933, w6934, w6935, w6936, w6937, w6938, w6939, w6940, w6941, w6942, w6943, w6944, w6945, w6946, w6947, w6948, w6949, w6950, w6951, w6952, w6953, w6954, w6955, w6956, w6957, w6958, w6959, w6960, w6961, w6962, w6963, w6964, w6965, w6966, w6967, w6968, w6969, w6970, w6971, w6972, w6973, w6974, w6975, w6976, w6977, w6978, w6979, w6980, w6981, w6982, w6983, w6984, w6985, w6986, w6987, w6988, w6989, w6990, w6991, w6992, w6993, w6994, w6995, w6996, w6997, w6998, w6999, w7000, w7001, w7002, w7003, w7004, w7005, w7006, w7007, w7008, w7009, w7010, w7011, w7012, w7013, w7014, w7015, w7016, w7017, w7018, w7019, w7020, w7021, w7022, w7023, w7024, w7025, w7026, w7027, w7028, w7029, w7030, w7031, w7032, w7033, w7034, w7035, w7036, w7037, w7038, w7039, w7040, w7041, w7042, w7043, w7044, w7045, w7046, w7047, w7048, w7049, w7050, w7051, w7052, w7053, w7054, w7055, w7056, w7057, w7058, w7059, w7060, w7061, w7062, w7063, w7064, w7065, w7066, w7067, w7068, w7069, w7070, w7071, w7072, w7073, w7074, w7075, w7076, w7077, w7078, w7079, w7080, w7081, w7082, w7083, w7084, w7085, w7086, w7087, w7088, w7089, w7090, w7091, w7092, w7093, w7094, w7095, w7096, w7097, w7098, w7099, w7100, w7101, w7102, w7103, w7104, w7105, w7106, w7107, w7108, w7109, w7110, w7111, w7112, w7113, w7114, w7115, w7116, w7117, w7118, w7119, w7120, w7121, w7122, w7123, w7124, w7125, w7126, w7127, w7128, w7129, w7130, w7131, w7132, w7133, w7134, w7135, w7136, w7137, w7138, w7139, w7140, w7141, w7142, w7143, w7144, w7145, w7146, w7147, w7148, w7149, w7150, w7151, w7152, w7153, w7154, w7155, w7156, w7157, w7158, w7159, w7160, w7161, w7162, w7163, w7164, w7165, w7166, w7167, w7168, w7169, w7170, w7171, w7172, w7173, w7174, w7175, w7176, w7177, w7178, w7179, w7180, w7181, w7182, w7183, w7184, w7185, w7186, w7187, w7188, w7189, w7190, w7191, w7192, w7193, w7194, w7195, w7196, w7197, w7198, w7199, w7200, w7201, w7202, w7203, w7204, w7205, w7206, w7207, w7208, w7209, w7210, w7211, w7212, w7213, w7214, w7215, w7216, w7217, w7218, w7219, w7220, w7221, w7222, w7223, w7224, w7225, w7226, w7227, w7228, w7229, w7230, w7231, w7232, w7233, w7234, w7235, w7236, w7237, w7238, w7239, w7240, w7241, w7242, w7243, w7244, w7245, w7246, w7247, w7248, w7249, w7250, w7251, w7252, w7253, w7254, w7255, w7256, w7257, w7258, w7259, w7260, w7261, w7262, w7263, w7264, w7265, w7266, w7267, w7268, w7269, w7270, w7271, w7272, w7273, w7274, w7275, w7276, w7277, w7278, w7279, w7280, w7281, w7282, w7283, w7284, w7285, w7286, w7287, w7288, w7289, w7290, w7291, w7292, w7293, w7294, w7295, w7296, w7297, w7298, w7299, w7300, w7301, w7302, w7303, w7304, w7305, w7306, w7307, w7308, w7309, w7310, w7311, w7312, w7313, w7314, w7315, w7316, w7317, w7318, w7319, w7320, w7321, w7322, w7323, w7324, w7325, w7326, w7327, w7328, w7329, w7330, w7331, w7332, w7333, w7334, w7335, w7336, w7337, w7338, w7339, w7340, w7341, w7342, w7343, w7344, w7345, w7346, w7347, w7348, w7349, w7350, w7351, w7352, w7353, w7354, w7355, w7356, w7357, w7358, w7359, w7360, w7361, w7362, w7363, w7364, w7365, w7366, w7367, w7368, w7369, w7370, w7371, w7372, w7373, w7374, w7375, w7376, w7377, w7378, w7379, w7380, w7381, w7382, w7383, w7384, w7385, w7386, w7387, w7388, w7389, w7390, w7391, w7392, w7393, w7394, w7395, w7396, w7397, w7398, w7399, w7400, w7401, w7402, w7403, w7404, w7405, w7406, w7407, w7408, w7409, w7410, w7411, w7412, w7413, w7414, w7415, w7416, w7417, w7418, w7419, w7420, w7421, w7422, w7423, w7424, w7425, w7426, w7427, w7428, w7429, w7430, w7431, w7432, w7433, w7434, w7435, w7436, w7437, w7438, w7439, w7440, w7441, w7442, w7443, w7444, w7445, w7446, w7447, w7448, w7449, w7450, w7451, w7452, w7453, w7454, w7455, w7456, w7457, w7458, w7459, w7460, w7461, w7462, w7463, w7464, w7465, w7466, w7467, w7468, w7469, w7470, w7471, w7472, w7473, w7474, w7475, w7476, w7477, w7478, w7479, w7480, w7481, w7482, w7483, w7484, w7485, w7486, w7487, w7488, w7489, w7490, w7491, w7492, w7493, w7494, w7495, w7496, w7497, w7498, w7499, w7500, w7501, w7502, w7503, w7504, w7505, w7506, w7507, w7508, w7509, w7510, w7511, w7512, w7513, w7514, w7515, w7516, w7517, w7518, w7519, w7520, w7521, w7522, w7523, w7524, w7525, w7526, w7527, w7528, w7529, w7530, w7531, w7532, w7533, w7534, w7535, w7536, w7537, w7538, w7539, w7540, w7541, w7542, w7543, w7544, w7545, w7546, w7547, w7548, w7549, w7550, w7551, w7552, w7553, w7554, w7555, w7556, w7557, w7558, w7559, w7560, w7561, w7562, w7563, w7564, w7565, w7566, w7567, w7568, w7569, w7570, w7571, w7572, w7573, w7574, w7575, w7576, w7577, w7578, w7579, w7580, w7581, w7582, w7583, w7584, w7585, w7586, w7587, w7588, w7589, w7590, w7591, w7592, w7593, w7594, w7595, w7596, w7597, w7598, w7599, w7600, w7601, w7602, w7603, w7604, w7605, w7606, w7607, w7608, w7609, w7610, w7611, w7612, w7613, w7614, w7615, w7616, w7617, w7618, w7619, w7620, w7621, w7622, w7623, w7624, w7625, w7626, w7627, w7628, w7629, w7630, w7631, w7632, w7633, w7634, w7635, w7636, w7637, w7638, w7639, w7640, w7641, w7642, w7643, w7644, w7645, w7646, w7647, w7648, w7649, w7650, w7651, w7652, w7653, w7654, w7655, w7656, w7657, w7658, w7659, w7660, w7661, w7662, w7663, w7664, w7665, w7666, w7667, w7668, w7669, w7670, w7671, w7672, w7673, w7674, w7675, w7676, w7677, w7678, w7679, w7680, w7681, w7682, w7683, w7684, w7685, w7686, w7687, w7688, w7689, w7690, w7691, w7692, w7693, w7694, w7695, w7696, w7697, w7698, w7699, w7700, w7701, w7702, w7703, w7704, w7705, w7706, w7707, w7708, w7709, w7710, w7711, w7712, w7713, w7714, w7715, w7716, w7717, w7718, w7719, w7720, w7721, w7722, w7723, w7724, w7725, w7726, w7727, w7728, w7729, w7730, w7731, w7732, w7733, w7734, w7735, w7736, w7737, w7738, w7739, w7740, w7741, w7742, w7743, w7744, w7745, w7746, w7747, w7748, w7749, w7750, w7751, w7752, w7753, w7754, w7755, w7756, w7757, w7758, w7759, w7760, w7761, w7762, w7763, w7764, w7765, w7766, w7767, w7768, w7769, w7770, w7771, w7772, w7773, w7774, w7775, w7776, w7777, w7778, w7779, w7780, w7781, w7782, w7783, w7784, w7785, w7786, w7787, w7788, w7789, w7790, w7791, w7792, w7793, w7794, w7795, w7796, w7797, w7798, w7799, w7800, w7801, w7802, w7803, w7804, w7805, w7806, w7807, w7808, w7809, w7810, w7811, w7812, w7813, w7814, w7815, w7816, w7817, w7818, w7819, w7820, w7821, w7822, w7823, w7824, w7825, w7826, w7827, w7828, w7829, w7830, w7831, w7832, w7833, w7834, w7835, w7836, w7837, w7838, w7839, w7840, w7841, w7842, w7843, w7844, w7845, w7846, w7847, w7848, w7849, w7850, w7851, w7852, w7853, w7854, w7855, w7856, w7857, w7858, w7859, w7860, w7861, w7862, w7863, w7864, w7865, w7866, w7867, w7868, w7869, w7870, w7871, w7872, w7873, w7874, w7875, w7876, w7877, w7878, w7879, w7880, w7881, w7882, w7883, w7884, w7885, w7886, w7887, w7888, w7889, w7890, w7891, w7892, w7893, w7894, w7895, w7896, w7897, w7898, w7899, w7900, w7901, w7902, w7903, w7904, w7905, w7906, w7907, w7908, w7909, w7910, w7911, w7912, w7913, w7914, w7915, w7916, w7917, w7918, w7919, w7920, w7921, w7922, w7923, w7924, w7925, w7926, w7927, w7928, w7929, w7930, w7931, w7932, w7933, w7934, w7935, w7936, w7937, w7938, w7939, w7940, w7941, w7942, w7943, w7944, w7945, w7946, w7947, w7948, w7949, w7950, w7951, w7952, w7953, w7954, w7955, w7956, w7957, w7958, w7959, w7960, w7961, w7962, w7963, w7964, w7965, w7966, w7967, w7968, w7969, w7970, w7971, w7972, w7973, w7974, w7975, w7976, w7977, w7978, w7979, w7980, w7981, w7982, w7983, w7984, w7985, w7986, w7987, w7988, w7989, w7990, w7991, w7992, w7993, w7994, w7995, w7996, w7997, w7998, w7999, w8000, w8001, w8002, w8003, w8004, w8005, w8006, w8007, w8008, w8009, w8010, w8011, w8012, w8013, w8014, w8015, w8016, w8017, w8018, w8019, w8020, w8021, w8022, w8023, w8024, w8025, w8026, w8027, w8028, w8029, w8030, w8031, w8032, w8033, w8034, w8035, w8036, w8037, w8038, w8039, w8040, w8041, w8042, w8043, w8044, w8045, w8046, w8047, w8048, w8049, w8050, w8051, w8052, w8053, w8054, w8055, w8056, w8057, w8058, w8059, w8060, w8061, w8062, w8063, w8064, w8065, w8066, w8067, w8068, w8069, w8070, w8071, w8072, w8073, w8074, w8075, w8076, w8077, w8078, w8079, w8080, w8081, w8082, w8083, w8084, w8085, w8086, w8087, w8088, w8089, w8090, w8091, w8092, w8093, w8094, w8095, w8096, w8097, w8098, w8099, w8100, w8101, w8102, w8103, w8104, w8105, w8106, w8107, w8108, w8109, w8110, w8111, w8112, w8113, w8114, w8115, w8116, w8117, w8118, w8119, w8120, w8121, w8122, w8123, w8124, w8125, w8126, w8127, w8128, w8129, w8130, w8131, w8132, w8133, w8134, w8135, w8136, w8137, w8138, w8139, w8140, w8141, w8142, w8143, w8144, w8145, w8146, w8147, w8148, w8149, w8150, w8151, w8152, w8153, w8154, w8155, w8156, w8157, w8158, w8159, w8160, w8161, w8162, w8163, w8164, w8165, w8166, w8167, w8168, w8169, w8170, w8171, w8172, w8173, w8174, w8175, w8176, w8177, w8178, w8179, w8180, w8181, w8182, w8183, w8184, w8185, w8186, w8187, w8188, w8189, w8190, w8191, w8192, w8193, w8194, w8195, w8196, w8197, w8198, w8199, w8200, w8201, w8202, w8203, w8204, w8205, w8206, w8207, w8208, w8209, w8210, w8211, w8212, w8213, w8214, w8215, w8216, w8217, w8218, w8219, w8220, w8221, w8222, w8223, w8224, w8225, w8226, w8227, w8228, w8229, w8230, w8231, w8232, w8233, w8234, w8235, w8236, w8237, w8238, w8239, w8240, w8241, w8242, w8243, w8244, w8245, w8246, w8247, w8248, w8249, w8250, w8251, w8252, w8253, w8254, w8255, w8256, w8257, w8258, w8259, w8260, w8261, w8262, w8263, w8264, w8265, w8266, w8267, w8268, w8269, w8270, w8271, w8272, w8273, w8274, w8275, w8276, w8277, w8278, w8279, w8280, w8281, w8282, w8283, w8284, w8285, w8286, w8287, w8288, w8289, w8290, w8291, w8292, w8293, w8294, w8295, w8296, w8297, w8298, w8299, w8300, w8301, w8302, w8303, w8304, w8305, w8306, w8307, w8308, w8309, w8310, w8311, w8312, w8313, w8314, w8315, w8316, w8317, w8318, w8319, w8320, w8321, w8322, w8323, w8324, w8325, w8326, w8327, w8328, w8329, w8330, w8331, w8332, w8333, w8334, w8335, w8336, w8337, w8338, w8339, w8340, w8341, w8342, w8343, w8344, w8345, w8346, w8347, w8348, w8349, w8350, w8351, w8352, w8353, w8354, w8355, w8356, w8357, w8358, w8359, w8360, w8361, w8362, w8363, w8364, w8365, w8366, w8367, w8368, w8369, w8370, w8371, w8372, w8373, w8374, w8375, w8376, w8377, w8378, w8379, w8380, w8381, w8382, w8383, w8384, w8385, w8386, w8387, w8388, w8389, w8390, w8391, w8392, w8393, w8394, w8395, w8396, w8397, w8398, w8399, w8400, w8401, w8402, w8403, w8404, w8405, w8406, w8407, w8408, w8409, w8410, w8411, w8412, w8413, w8414, w8415, w8416, w8417, w8418, w8419, w8420, w8421, w8422, w8423, w8424, w8425, w8426, w8427, w8428, w8429, w8430, w8431, w8432, w8433, w8434, w8435, w8436, w8437, w8438, w8439, w8440, w8441, w8442, w8443, w8444, w8445, w8446, w8447, w8448, w8449, w8450, w8451, w8452, w8453, w8454, w8455, w8456, w8457, w8458, w8459, w8460, w8461, w8462, w8463, w8464, w8465, w8466, w8467, w8468, w8469, w8470, w8471, w8472, w8473, w8474, w8475, w8476, w8477, w8478, w8479, w8480, w8481, w8482, w8483, w8484, w8485, w8486, w8487, w8488, w8489, w8490, w8491, w8492, w8493, w8494, w8495, w8496, w8497, w8498, w8499, w8500, w8501, w8502, w8503, w8504, w8505, w8506, w8507, w8508, w8509, w8510, w8511, w8512, w8513, w8514, w8515, w8516, w8517, w8518, w8519, w8520, w8521, w8522, w8523, w8524, w8525, w8526, w8527, w8528, w8529, w8530, w8531, w8532, w8533, w8534, w8535, w8536, w8537, w8538, w8539, w8540, w8541, w8542, w8543, w8544, w8545, w8546, w8547, w8548, w8549, w8550, w8551, w8552, w8553, w8554, w8555, w8556, w8557, w8558, w8559, w8560, w8561, w8562, w8563, w8564, w8565, w8566, w8567, w8568, w8569, w8570, w8571, w8572, w8573, w8574, w8575, w8576, w8577, w8578, w8579, w8580, w8581, w8582, w8583, w8584, w8585, w8586, w8587, w8588, w8589, w8590, w8591, w8592, w8593, w8594, w8595, w8596, w8597, w8598, w8599, w8600, w8601, w8602, w8603, w8604, w8605, w8606, w8607, w8608, w8609, w8610, w8611, w8612, w8613, w8614, w8615, w8616, w8617, w8618, w8619, w8620, w8621, w8622, w8623, w8624, w8625, w8626, w8627, w8628, w8629, w8630, w8631, w8632, w8633, w8634, w8635, w8636, w8637, w8638, w8639, w8640, w8641, w8642, w8643, w8644, w8645, w8646, w8647, w8648, w8649, w8650, w8651, w8652, w8653, w8654, w8655, w8656, w8657, w8658, w8659, w8660, w8661, w8662, w8663, w8664, w8665, w8666, w8667, w8668, w8669, w8670, w8671, w8672, w8673, w8674, w8675, w8676, w8677, w8678, w8679, w8680, w8681, w8682, w8683, w8684, w8685, w8686, w8687, w8688, w8689, w8690, w8691, w8692, w8693, w8694, w8695, w8696, w8697, w8698, w8699, w8700, w8701, w8702, w8703, w8704, w8705, w8706, w8707, w8708, w8709, w8710, w8711, w8712, w8713, w8714, w8715, w8716, w8717, w8718, w8719, w8720, w8721, w8722, w8723, w8724, w8725, w8726, w8727, w8728, w8729, w8730, w8731, w8732, w8733, w8734, w8735, w8736, w8737, w8738, w8739, w8740, w8741, w8742, w8743, w8744, w8745, w8746, w8747, w8748, w8749, w8750, w8751, w8752, w8753, w8754, w8755, w8756, w8757, w8758, w8759, w8760, w8761, w8762, w8763, w8764, w8765, w8766, w8767, w8768, w8769, w8770, w8771, w8772, w8773, w8774, w8775, w8776, w8777, w8778, w8779, w8780, w8781, w8782, w8783, w8784, w8785, w8786, w8787, w8788, w8789, w8790, w8791, w8792, w8793, w8794, w8795, w8796, w8797, w8798, w8799, w8800, w8801, w8802, w8803, w8804, w8805, w8806, w8807, w8808, w8809, w8810, w8811, w8812, w8813, w8814, w8815, w8816, w8817, w8818, w8819, w8820, w8821, w8822, w8823, w8824, w8825, w8826, w8827, w8828, w8829, w8830, w8831, w8832, w8833, w8834, w8835, w8836, w8837, w8838, w8839, w8840, w8841, w8842, w8843, w8844, w8845, w8846, w8847, w8848, w8849, w8850, w8851, w8852, w8853, w8854, w8855, w8856, w8857, w8858, w8859, w8860, w8861, w8862, w8863, w8864, w8865, w8866, w8867, w8868, w8869, w8870, w8871, w8872, w8873, w8874, w8875, w8876, w8877, w8878, w8879, w8880, w8881, w8882, w8883, w8884, w8885, w8886, w8887, w8888, w8889, w8890, w8891, w8892, w8893, w8894, w8895, w8896, w8897, w8898, w8899, w8900, w8901, w8902, w8903, w8904, w8905, w8906, w8907, w8908, w8909, w8910, w8911, w8912, w8913, w8914, w8915, w8916, w8917, w8918, w8919, w8920, w8921, w8922, w8923, w8924, w8925, w8926, w8927, w8928, w8929, w8930, w8931, w8932, w8933, w8934, w8935, w8936, w8937, w8938, w8939, w8940, w8941, w8942, w8943, w8944, w8945, w8946, w8947, w8948, w8949, w8950, w8951, w8952, w8953, w8954, w8955, w8956, w8957, w8958, w8959, w8960, w8961, w8962, w8963, w8964, w8965, w8966, w8967, w8968, w8969, w8970, w8971, w8972, w8973, w8974, w8975, w8976, w8977, w8978, w8979, w8980, w8981, w8982, w8983, w8984, w8985, w8986, w8987, w8988, w8989, w8990, w8991, w8992, w8993, w8994, w8995, w8996, w8997, w8998, w8999, w9000, w9001, w9002, w9003, w9004, w9005, w9006, w9007, w9008, w9009, w9010, w9011, w9012, w9013, w9014, w9015, w9016, w9017, w9018, w9019, w9020, w9021, w9022, w9023, w9024, w9025, w9026, w9027, w9028, w9029, w9030, w9031, w9032, w9033, w9034, w9035, w9036, w9037, w9038, w9039, w9040, w9041, w9042, w9043, w9044, w9045, w9046, w9047, w9048, w9049, w9050, w9051, w9052, w9053, w9054, w9055, w9056, w9057, w9058, w9059, w9060, w9061, w9062, w9063, w9064, w9065, w9066, w9067, w9068, w9069, w9070, w9071, w9072, w9073, w9074, w9075, w9076, w9077, w9078, w9079, w9080, w9081, w9082, w9083, w9084, w9085, w9086, w9087, w9088, w9089, w9090, w9091, w9092, w9093, w9094, w9095, w9096, w9097, w9098, w9099, w9100, w9101, w9102, w9103, w9104, w9105, w9106, w9107, w9108, w9109, w9110, w9111, w9112, w9113, w9114, w9115, w9116, w9117, w9118, w9119, w9120, w9121, w9122, w9123, w9124, w9125, w9126, w9127, w9128, w9129, w9130, w9131, w9132, w9133, w9134, w9135, w9136, w9137, w9138, w9139, w9140, w9141, w9142, w9143, w9144, w9145, w9146, w9147, w9148, w9149, w9150, w9151, w9152, w9153, w9154, w9155, w9156, w9157, w9158, w9159, w9160, w9161, w9162, w9163, w9164, w9165, w9166, w9167, w9168, w9169, w9170, w9171, w9172, w9173, w9174, w9175, w9176, w9177, w9178, w9179, w9180, w9181, w9182, w9183, w9184, w9185, w9186, w9187, w9188, w9189, w9190, w9191, w9192, w9193, w9194, w9195, w9196, w9197, w9198, w9199, w9200, w9201, w9202, w9203, w9204, w9205, w9206, w9207, w9208, w9209, w9210, w9211, w9212, w9213, w9214, w9215, w9216, w9217, w9218, w9219, w9220, w9221, w9222, w9223, w9224, w9225, w9226, w9227, w9228, w9229, w9230, w9231, w9232, w9233, w9234, w9235, w9236, w9237, w9238, w9239, w9240, w9241, w9242, w9243, w9244, w9245, w9246, w9247, w9248, w9249, w9250, w9251, w9252, w9253, w9254, w9255, w9256, w9257, w9258, w9259, w9260, w9261, w9262, w9263, w9264, w9265, w9266, w9267, w9268, w9269, w9270, w9271, w9272, w9273, w9274, w9275, w9276, w9277, w9278, w9279, w9280, w9281, w9282, w9283, w9284, w9285, w9286, w9287, w9288, w9289, w9290, w9291, w9292, w9293, w9294, w9295, w9296, w9297, w9298, w9299, w9300, w9301, w9302, w9303, w9304, w9305, w9306, w9307, w9308, w9309, w9310, w9311, w9312, w9313, w9314, w9315, w9316, w9317, w9318, w9319, w9320, w9321, w9322, w9323, w9324, w9325, w9326, w9327, w9328, w9329, w9330, w9331, w9332, w9333, w9334, w9335, w9336, w9337, w9338, w9339, w9340, w9341, w9342, w9343, w9344, w9345, w9346, w9347, w9348, w9349, w9350, w9351, w9352, w9353, w9354, w9355, w9356, w9357, w9358, w9359, w9360, w9361, w9362, w9363, w9364, w9365, w9366, w9367, w9368, w9369, w9370, w9371, w9372, w9373, w9374, w9375, w9376, w9377, w9378, w9379, w9380, w9381, w9382, w9383, w9384, w9385, w9386, w9387, w9388, w9389, w9390, w9391, w9392, w9393, w9394, w9395, w9396, w9397, w9398, w9399, w9400, w9401, w9402, w9403, w9404, w9405, w9406, w9407, w9408, w9409, w9410, w9411, w9412, w9413, w9414, w9415, w9416, w9417, w9418, w9419, w9420, w9421, w9422, w9423, w9424, w9425, w9426, w9427, w9428, w9429, w9430, w9431, w9432, w9433, w9434, w9435, w9436, w9437, w9438, w9439, w9440, w9441, w9442, w9443, w9444, w9445, w9446, w9447, w9448, w9449, w9450, w9451, w9452, w9453, w9454, w9455, w9456, w9457, w9458, w9459, w9460, w9461, w9462, w9463, w9464, w9465, w9466, w9467, w9468, w9469, w9470, w9471, w9472, w9473, w9474, w9475, w9476, w9477, w9478, w9479, w9480, w9481, w9482, w9483, w9484, w9485, w9486, w9487, w9488, w9489, w9490, w9491, w9492, w9493, w9494, w9495, w9496, w9497, w9498, w9499, w9500, w9501, w9502, w9503, w9504, w9505, w9506, w9507, w9508, w9509, w9510, w9511, w9512, w9513, w9514, w9515, w9516, w9517, w9518, w9519, w9520, w9521, w9522, w9523, w9524, w9525, w9526, w9527, w9528, w9529, w9530, w9531, w9532, w9533, w9534, w9535, w9536, w9537, w9538, w9539, w9540, w9541, w9542, w9543, w9544, w9545, w9546, w9547, w9548, w9549, w9550, w9551, w9552, w9553, w9554, w9555, w9556, w9557, w9558, w9559, w9560, w9561, w9562, w9563, w9564, w9565, w9566, w9567, w9568, w9569, w9570, w9571, w9572, w9573, w9574, w9575, w9576, w9577, w9578, w9579, w9580, w9581, w9582, w9583, w9584, w9585, w9586, w9587, w9588, w9589, w9590, w9591, w9592, w9593, w9594, w9595, w9596, w9597, w9598, w9599, w9600, w9601, w9602, w9603, w9604, w9605, w9606, w9607, w9608, w9609, w9610, w9611, w9612, w9613, w9614, w9615, w9616, w9617, w9618, w9619, w9620, w9621, w9622, w9623, w9624, w9625, w9626, w9627, w9628, w9629, w9630, w9631, w9632, w9633, w9634, w9635, w9636, w9637, w9638, w9639, w9640, w9641, w9642, w9643, w9644, w9645, w9646, w9647, w9648, w9649, w9650, w9651, w9652, w9653, w9654, w9655, w9656, w9657, w9658, w9659, w9660, w9661, w9662, w9663, w9664, w9665, w9666, w9667, w9668, w9669, w9670, w9671, w9672, w9673, w9674, w9675, w9676, w9677, w9678, w9679, w9680, w9681, w9682, w9683, w9684, w9685, w9686, w9687, w9688, w9689, w9690, w9691, w9692, w9693, w9694, w9695, w9696, w9697, w9698, w9699, w9700, w9701, w9702, w9703, w9704, w9705, w9706, w9707, w9708, w9709, w9710, w9711, w9712, w9713, w9714, w9715, w9716, w9717, w9718, w9719, w9720, w9721, w9722, w9723, w9724, w9725, w9726, w9727, w9728, w9729, w9730, w9731, w9732, w9733, w9734, w9735, w9736, w9737, w9738, w9739, w9740, w9741, w9742, w9743, w9744, w9745, w9746, w9747, w9748, w9749, w9750, w9751, w9752, w9753, w9754, w9755, w9756, w9757, w9758, w9759, w9760, w9761, w9762, w9763, w9764, w9765, w9766, w9767, w9768, w9769, w9770, w9771, w9772, w9773, w9774, w9775, w9776, w9777, w9778, w9779, w9780, w9781, w9782, w9783, w9784, w9785, w9786, w9787, w9788, w9789, w9790, w9791, w9792, w9793, w9794, w9795, w9796, w9797, w9798, w9799, w9800, w9801, w9802, w9803, w9804, w9805, w9806, w9807, w9808, w9809, w9810, w9811, w9812, w9813, w9814, w9815, w9816, w9817, w9818, w9819, w9820, w9821, w9822, w9823, w9824, w9825, w9826, w9827, w9828, w9829, w9830, w9831, w9832, w9833, w9834, w9835, w9836, w9837, w9838, w9839, w9840, w9841, w9842, w9843, w9844, w9845, w9846, w9847, w9848, w9849, w9850, w9851, w9852, w9853, w9854, w9855, w9856, w9857, w9858, w9859, w9860, w9861, w9862, w9863, w9864, w9865, w9866, w9867, w9868, w9869, w9870, w9871, w9872, w9873, w9874, w9875, w9876, w9877, w9878, w9879, w9880, w9881, w9882, w9883, w9884, w9885, w9886, w9887, w9888, w9889, w9890, w9891, w9892, w9893, w9894, w9895, w9896, w9897, w9898, w9899, w9900, w9901, w9902, w9903, w9904, w9905, w9906, w9907, w9908, w9909, w9910, w9911, w9912, w9913, w9914, w9915, w9916, w9917, w9918, w9919, w9920, w9921, w9922, w9923, w9924, w9925, w9926, w9927, w9928, w9929, w9930, w9931, w9932, w9933, w9934, w9935, w9936, w9937, w9938, w9939, w9940, w9941, w9942, w9943, w9944, w9945, w9946, w9947, w9948, w9949, w9950, w9951, w9952, w9953, w9954, w9955, w9956, w9957, w9958, w9959, w9960, w9961, w9962, w9963, w9964, w9965, w9966, w9967, w9968, w9969, w9970, w9971, w9972, w9973, w9974, w9975, w9976, w9977, w9978, w9979, w9980, w9981, w9982, w9983, w9984, w9985, w9986, w9987, w9988, w9989, w9990, w9991, w9992, w9993, w9994, w9995, w9996, w9997, w9998, w9999, w10000, w10001, w10002, w10003, w10004, w10005, w10006, w10007, w10008, w10009, w10010, w10011, w10012, w10013, w10014, w10015, w10016, w10017, w10018, w10019, w10020, w10021, w10022, w10023, w10024, w10025, w10026, w10027, w10028, w10029, w10030, w10031, w10032, w10033, w10034, w10035, w10036, w10037, w10038, w10039, w10040, w10041, w10042, w10043, w10044, w10045, w10046, w10047, w10048, w10049, w10050, w10051, w10052, w10053, w10054, w10055, w10056, w10057, w10058, w10059, w10060, w10061, w10062, w10063, w10064, w10065, w10066, w10067, w10068, w10069, w10070, w10071, w10072, w10073, w10074, w10075, w10076, w10077, w10078, w10079, w10080, w10081, w10082, w10083, w10084, w10085, w10086, w10087, w10088, w10089, w10090, w10091, w10092, w10093, w10094, w10095, w10096, w10097, w10098, w10099, w10100, w10101, w10102, w10103, w10104, w10105, w10106, w10107, w10108, w10109, w10110, w10111, w10112, w10113, w10114, w10115, w10116, w10117, w10118, w10119, w10120, w10121, w10122, w10123, w10124, w10125, w10126, w10127, w10128, w10129, w10130, w10131, w10132, w10133, w10134, w10135, w10136, w10137, w10138, w10139, w10140, w10141, w10142, w10143, w10144, w10145, w10146, w10147, w10148, w10149, w10150, w10151, w10152, w10153, w10154, w10155, w10156, w10157, w10158, w10159, w10160, w10161, w10162, w10163, w10164, w10165, w10166, w10167, w10168, w10169, w10170, w10171, w10172, w10173, w10174, w10175, w10176, w10177, w10178, w10179, w10180, w10181, w10182, w10183, w10184, w10185, w10186, w10187, w10188, w10189, w10190, w10191, w10192, w10193, w10194, w10195, w10196, w10197, w10198, w10199, w10200, w10201, w10202, w10203, w10204, w10205, w10206, w10207, w10208, w10209, w10210, w10211, w10212, w10213, w10214, w10215, w10216, w10217, w10218, w10219, w10220, w10221, w10222, w10223, w10224, w10225, w10226, w10227, w10228, w10229, w10230, w10231, w10232, w10233, w10234, w10235, w10236, w10237, w10238, w10239, w10240, w10241, w10242, w10243, w10244, w10245, w10246, w10247, w10248, w10249, w10250, w10251, w10252, w10253, w10254, w10255, w10256, w10257, w10258, w10259, w10260, w10261, w10262, w10263, w10264, w10265, w10266, w10267, w10268, w10269, w10270, w10271, w10272, w10273, w10274, w10275, w10276, w10277, w10278, w10279, w10280, w10281, w10282, w10283, w10284, w10285, w10286, w10287, w10288, w10289, w10290, w10291, w10292, w10293, w10294, w10295, w10296, w10297, w10298, w10299, w10300, w10301, w10302, w10303, w10304, w10305, w10306, w10307, w10308, w10309, w10310, w10311, w10312, w10313, w10314, w10315, w10316, w10317, w10318, w10319, w10320, w10321, w10322, w10323, w10324, w10325, w10326, w10327, w10328, w10329, w10330, w10331, w10332, w10333, w10334, w10335, w10336, w10337, w10338, w10339, w10340, w10341, w10342, w10343, w10344, w10345, w10346, w10347, w10348, w10349, w10350, w10351, w10352, w10353, w10354, w10355, w10356, w10357, w10358, w10359, w10360, w10361, w10362, w10363, w10364, w10365, w10366, w10367, w10368, w10369, w10370, w10371, w10372, w10373, w10374, w10375, w10376, w10377, w10378, w10379, w10380, w10381, w10382, w10383, w10384, w10385, w10386, w10387, w10388, w10389, w10390, w10391, w10392, w10393, w10394, w10395, w10396, w10397, w10398, w10399, w10400, w10401, w10402, w10403, w10404, w10405, w10406, w10407, w10408, w10409, w10410, w10411, w10412, w10413, w10414, w10415, w10416, w10417, w10418, w10419, w10420, w10421, w10422, w10423, w10424, w10425, w10426, w10427, w10428, w10429, w10430, w10431, w10432, w10433, w10434, w10435, w10436, w10437, w10438, w10439, w10440, w10441, w10442, w10443, w10444, w10445, w10446, w10447, w10448, w10449, w10450, w10451, w10452, w10453, w10454, w10455, w10456, w10457, w10458, w10459, w10460, w10461, w10462, w10463, w10464, w10465, w10466, w10467, w10468, w10469, w10470, w10471, w10472, w10473, w10474, w10475, w10476, w10477, w10478, w10479, w10480, w10481, w10482, w10483, w10484, w10485, w10486, w10487, w10488, w10489, w10490, w10491, w10492, w10493, w10494, w10495, w10496, w10497, w10498, w10499, w10500, w10501, w10502, w10503, w10504, w10505, w10506, w10507, w10508, w10509, w10510, w10511, w10512, w10513, w10514, w10515, w10516, w10517, w10518, w10519, w10520, w10521, w10522, w10523, w10524, w10525, w10526, w10527, w10528, w10529, w10530, w10531, w10532, w10533, w10534, w10535, w10536, w10537, w10538, w10539, w10540, w10541, w10542, w10543, w10544, w10545, w10546, w10547, w10548, w10549, w10550, w10551, w10552, w10553, w10554, w10555, w10556, w10557, w10558, w10559, w10560, w10561, w10562, w10563, w10564, w10565, w10566, w10567, w10568, w10569, w10570, w10571, w10572, w10573, w10574, w10575, w10576, w10577, w10578, w10579, w10580, w10581, w10582, w10583, w10584, w10585, w10586, w10587, w10588, w10589, w10590, w10591, w10592, w10593, w10594, w10595, w10596, w10597, w10598, w10599, w10600, w10601, w10602, w10603, w10604, w10605, w10606, w10607, w10608, w10609, w10610, w10611, w10612, w10613, w10614, w10615, w10616, w10617, w10618, w10619, w10620, w10621, w10622, w10623, w10624, w10625, w10626, w10627, w10628, w10629, w10630, w10631, w10632, w10633, w10634, w10635, w10636, w10637, w10638, w10639, w10640, w10641, w10642, w10643, w10644, w10645, w10646, w10647, w10648, w10649, w10650, w10651, w10652, w10653, w10654, w10655, w10656, w10657, w10658, w10659, w10660, w10661, w10662, w10663, w10664, w10665, w10666, w10667, w10668, w10669, w10670, w10671, w10672, w10673, w10674, w10675, w10676, w10677, w10678, w10679, w10680, w10681, w10682, w10683, w10684, w10685, w10686, w10687, w10688, w10689, w10690, w10691, w10692, w10693, w10694, w10695, w10696, w10697, w10698, w10699, w10700, w10701, w10702, w10703, w10704, w10705, w10706, w10707, w10708, w10709, w10710, w10711, w10712, w10713, w10714, w10715, w10716, w10717, w10718, w10719, w10720, w10721, w10722, w10723, w10724, w10725, w10726, w10727, w10728, w10729, w10730, w10731, w10732, w10733, w10734, w10735, w10736, w10737, w10738, w10739, w10740, w10741, w10742, w10743, w10744, w10745, w10746, w10747, w10748, w10749, w10750, w10751, w10752, w10753, w10754, w10755, w10756, w10757, w10758, w10759, w10760, w10761, w10762, w10763, w10764, w10765, w10766, w10767, w10768, w10769, w10770, w10771, w10772, w10773, w10774, w10775, w10776, w10777, w10778, w10779, w10780, w10781, w10782, w10783, w10784, w10785, w10786, w10787, w10788, w10789, w10790, w10791, w10792, w10793, w10794, w10795, w10796, w10797, w10798, w10799, w10800, w10801, w10802, w10803, w10804, w10805, w10806, w10807, w10808, w10809, w10810, w10811, w10812, w10813, w10814, w10815, w10816, w10817, w10818, w10819, w10820, w10821, w10822, w10823, w10824, w10825, w10826, w10827, w10828, w10829, w10830, w10831, w10832, w10833, w10834, w10835, w10836, w10837, w10838, w10839, w10840, w10841, w10842, w10843, w10844, w10845, w10846, w10847, w10848, w10849, w10850, w10851, w10852, w10853, w10854, w10855, w10856, w10857, w10858, w10859, w10860, w10861, w10862, w10863, w10864, w10865, w10866, w10867, w10868, w10869, w10870, w10871, w10872, w10873, w10874, w10875, w10876, w10877, w10878, w10879, w10880, w10881, w10882, w10883, w10884, w10885, w10886, w10887, w10888, w10889, w10890, w10891, w10892, w10893, w10894, w10895, w10896, w10897, w10898, w10899, w10900, w10901, w10902, w10903, w10904, w10905, w10906, w10907, w10908, w10909, w10910, w10911, w10912, w10913, w10914, w10915, w10916, w10917, w10918, w10919, w10920, w10921, w10922, w10923, w10924, w10925, w10926, w10927, w10928, w10929, w10930, w10931, w10932, w10933, w10934, w10935, w10936, w10937, w10938, w10939, w10940, w10941, w10942, w10943, w10944, w10945, w10946, w10947, w10948, w10949, w10950, w10951, w10952, w10953, w10954, w10955, w10956, w10957, w10958, w10959, w10960, w10961, w10962, w10963, w10964, w10965, w10966, w10967, w10968, w10969, w10970, w10971, w10972, w10973, w10974, w10975, w10976, w10977, w10978, w10979, w10980, w10981, w10982, w10983, w10984, w10985, w10986, w10987, w10988, w10989, w10990, w10991, w10992, w10993, w10994, w10995, w10996, w10997, w10998, w10999, w11000, w11001, w11002, w11003, w11004, w11005, w11006, w11007, w11008, w11009, w11010, w11011, w11012, w11013, w11014, w11015, w11016, w11017, w11018, w11019, w11020, w11021, w11022, w11023, w11024, w11025, w11026, w11027, w11028, w11029, w11030, w11031, w11032, w11033, w11034, w11035, w11036, w11037, w11038, w11039, w11040, w11041, w11042, w11043, w11044, w11045, w11046, w11047, w11048, w11049, w11050, w11051, w11052, w11053, w11054, w11055, w11056, w11057, w11058, w11059, w11060, w11061, w11062, w11063, w11064, w11065, w11066, w11067, w11068, w11069, w11070, w11071, w11072, w11073, w11074, w11075, w11076, w11077, w11078, w11079, w11080, w11081, w11082, w11083, w11084, w11085, w11086, w11087, w11088, w11089, w11090, w11091, w11092, w11093, w11094, w11095, w11096, w11097, w11098, w11099, w11100, w11101, w11102, w11103, w11104, w11105, w11106, w11107, w11108, w11109, w11110, w11111, w11112, w11113, w11114, w11115, w11116, w11117, w11118, w11119, w11120, w11121, w11122, w11123, w11124, w11125, w11126, w11127, w11128, w11129, w11130, w11131, w11132, w11133, w11134, w11135, w11136, w11137, w11138, w11139, w11140, w11141, w11142, w11143, w11144, w11145, w11146, w11147, w11148, w11149, w11150, w11151, w11152, w11153, w11154, w11155, w11156, w11157, w11158, w11159, w11160, w11161, w11162, w11163, w11164, w11165, w11166, w11167, w11168, w11169, w11170, w11171, w11172, w11173, w11174, w11175, w11176, w11177, w11178, w11179, w11180, w11181, w11182, w11183, w11184, w11185, w11186, w11187, w11188, w11189, w11190, w11191, w11192, w11193, w11194, w11195, w11196, w11197, w11198, w11199, w11200, w11201, w11202, w11203, w11204, w11205, w11206, w11207, w11208, w11209, w11210, w11211, w11212, w11213, w11214, w11215, w11216, w11217, w11218, w11219, w11220, w11221, w11222, w11223, w11224, w11225, w11226, w11227, w11228, w11229, w11230, w11231, w11232, w11233, w11234, w11235, w11236, w11237, w11238, w11239, w11240, w11241, w11242, w11243, w11244, w11245, w11246, w11247, w11248, w11249, w11250, w11251, w11252, w11253, w11254, w11255, w11256, w11257, w11258, w11259, w11260, w11261, w11262, w11263, w11264, w11265, w11266, w11267, w11268, w11269, w11270, w11271, w11272, w11273, w11274, w11275, w11276, w11277, w11278, w11279, w11280, w11281, w11282, w11283, w11284, w11285, w11286, w11287, w11288, w11289, w11290, w11291, w11292, w11293, w11294, w11295, w11296, w11297, w11298, w11299, w11300, w11301, w11302, w11303, w11304, w11305, w11306, w11307, w11308, w11309, w11310, w11311, w11312, w11313, w11314, w11315, w11316, w11317, w11318, w11319, w11320, w11321, w11322, w11323, w11324, w11325, w11326, w11327, w11328, w11329, w11330, w11331, w11332, w11333, w11334, w11335, w11336, w11337, w11338, w11339, w11340, w11341, w11342, w11343, w11344, w11345, w11346, w11347, w11348, w11349, w11350, w11351, w11352, w11353, w11354, w11355, w11356, w11357, w11358, w11359, w11360, w11361, w11362, w11363, w11364, w11365, w11366, w11367, w11368, w11369, w11370, w11371, w11372, w11373, w11374, w11375, w11376, w11377, w11378, w11379, w11380, w11381, w11382, w11383, w11384, w11385, w11386, w11387, w11388, w11389, w11390, w11391, w11392, w11393, w11394, w11395, w11396, w11397, w11398, w11399, w11400, w11401, w11402, w11403, w11404, w11405, w11406, w11407, w11408, w11409, w11410, w11411, w11412, w11413, w11414, w11415, w11416, w11417, w11418, w11419, w11420, w11421, w11422, w11423, w11424, w11425, w11426, w11427, w11428, w11429, w11430, w11431, w11432, w11433, w11434, w11435, w11436, w11437, w11438, w11439, w11440, w11441, w11442, w11443, w11444, w11445, w11446, w11447, w11448, w11449, w11450, w11451, w11452, w11453, w11454, w11455, w11456, w11457, w11458, w11459, w11460, w11461, w11462, w11463, w11464, w11465, w11466, w11467, w11468, w11469, w11470, w11471, w11472, w11473, w11474, w11475, w11476, w11477, w11478, w11479, w11480, w11481, w11482, w11483, w11484, w11485, w11486, w11487, w11488, w11489, w11490, w11491, w11492, w11493, w11494, w11495, w11496, w11497, w11498, w11499, w11500, w11501, w11502, w11503, w11504, w11505, w11506, w11507, w11508, w11509, w11510, w11511, w11512, w11513, w11514, w11515, w11516, w11517, w11518, w11519, w11520, w11521, w11522, w11523, w11524, w11525, w11526, w11527, w11528, w11529, w11530, w11531, w11532, w11533, w11534, w11535, w11536, w11537, w11538, w11539, w11540, w11541, w11542, w11543, w11544, w11545, w11546, w11547, w11548, w11549, w11550, w11551, w11552, w11553, w11554, w11555, w11556, w11557, w11558, w11559, w11560, w11561, w11562, w11563, w11564, w11565, w11566, w11567, w11568, w11569, w11570, w11571, w11572, w11573, w11574, w11575, w11576, w11577, w11578, w11579, w11580, w11581, w11582, w11583, w11584, w11585, w11586, w11587, w11588, w11589, w11590, w11591, w11592, w11593, w11594, w11595, w11596, w11597, w11598, w11599, w11600, w11601, w11602, w11603, w11604, w11605, w11606, w11607, w11608, w11609, w11610, w11611, w11612, w11613, w11614, w11615, w11616, w11617, w11618, w11619, w11620, w11621, w11622, w11623, w11624, w11625, w11626, w11627, w11628, w11629, w11630, w11631, w11632, w11633, w11634, w11635, w11636, w11637, w11638, w11639, w11640, w11641, w11642, w11643, w11644, w11645, w11646, w11647, w11648, w11649, w11650, w11651, w11652, w11653, w11654, w11655, w11656, w11657, w11658, w11659, w11660, w11661, w11662, w11663, w11664, w11665, w11666, w11667, w11668, w11669, w11670, w11671, w11672, w11673, w11674, w11675, w11676, w11677, w11678, w11679, w11680, w11681, w11682, w11683, w11684, w11685, w11686, w11687, w11688, w11689, w11690, w11691, w11692, w11693, w11694, w11695, w11696, w11697, w11698, w11699, w11700, w11701, w11702, w11703, w11704, w11705, w11706, w11707, w11708, w11709, w11710, w11711, w11712, w11713, w11714, w11715, w11716, w11717, w11718, w11719, w11720, w11721, w11722, w11723, w11724, w11725, w11726, w11727, w11728, w11729, w11730, w11731, w11732, w11733, w11734, w11735, w11736, w11737, w11738, w11739, w11740, w11741, w11742, w11743, w11744, w11745, w11746, w11747, w11748, w11749, w11750, w11751, w11752, w11753, w11754, w11755, w11756, w11757, w11758, w11759, w11760, w11761, w11762, w11763, w11764, w11765, w11766, w11767, w11768, w11769, w11770, w11771, w11772, w11773, w11774, w11775, w11776, w11777, w11778, w11779, w11780, w11781, w11782, w11783, w11784, w11785, w11786, w11787, w11788, w11789, w11790, w11791, w11792, w11793, w11794, w11795, w11796, w11797, w11798, w11799, w11800, w11801, w11802, w11803, w11804, w11805, w11806, w11807, w11808, w11809, w11810, w11811, w11812, w11813, w11814, w11815, w11816, w11817, w11818, w11819, w11820, w11821, w11822, w11823, w11824, w11825, w11826, w11827, w11828, w11829, w11830, w11831, w11832, w11833, w11834, w11835, w11836, w11837, w11838, w11839, w11840, w11841, w11842, w11843, w11844, w11845, w11846, w11847, w11848, w11849, w11850, w11851, w11852, w11853, w11854, w11855, w11856, w11857, w11858, w11859, w11860, w11861, w11862, w11863, w11864, w11865, w11866, w11867, w11868, w11869, w11870, w11871, w11872, w11873, w11874, w11875, w11876, w11877, w11878, w11879, w11880, w11881, w11882, w11883, w11884, w11885, w11886, w11887, w11888, w11889, w11890, w11891, w11892, w11893, w11894, w11895, w11896, w11897, w11898, w11899, w11900, w11901, w11902, w11903, w11904, w11905, w11906, w11907, w11908, w11909, w11910, w11911, w11912, w11913, w11914, w11915, w11916, w11917, w11918, w11919, w11920, w11921, w11922, w11923, w11924, w11925, w11926, w11927, w11928, w11929, w11930, w11931, w11932, w11933, w11934, w11935, w11936, w11937, w11938, w11939, w11940, w11941, w11942, w11943, w11944, w11945, w11946, w11947, w11948, w11949, w11950, w11951, w11952, w11953, w11954, w11955, w11956, w11957, w11958, w11959, w11960, w11961, w11962, w11963, w11964, w11965, w11966, w11967, w11968, w11969, w11970, w11971, w11972, w11973, w11974, w11975, w11976, w11977, w11978, w11979, w11980, w11981, w11982, w11983, w11984, w11985, w11986, w11987, w11988, w11989, w11990, w11991, w11992, w11993, w11994, w11995, w11996, w11997, w11998, w11999, w12000, w12001, w12002, w12003, w12004, w12005, w12006, w12007, w12008, w12009, w12010, w12011, w12012, w12013, w12014, w12015, w12016, w12017, w12018, w12019, w12020, w12021, w12022, w12023, w12024, w12025, w12026, w12027, w12028, w12029, w12030, w12031, w12032, w12033, w12034, w12035, w12036, w12037, w12038, w12039, w12040, w12041, w12042, w12043, w12044, w12045, w12046, w12047, w12048, w12049, w12050, w12051, w12052, w12053, w12054, w12055, w12056, w12057, w12058, w12059, w12060, w12061, w12062, w12063, w12064, w12065, w12066, w12067, w12068, w12069, w12070, w12071, w12072, w12073, w12074, w12075, w12076, w12077, w12078, w12079, w12080, w12081, w12082, w12083, w12084, w12085, w12086, w12087, w12088, w12089, w12090, w12091, w12092, w12093, w12094, w12095, w12096, w12097, w12098, w12099, w12100, w12101, w12102, w12103, w12104, w12105, w12106, w12107, w12108, w12109, w12110, w12111, w12112, w12113, w12114, w12115, w12116, w12117, w12118, w12119, w12120, w12121, w12122, w12123, w12124, w12125, w12126, w12127, w12128, w12129, w12130, w12131, w12132, w12133, w12134, w12135, w12136, w12137, w12138, w12139, w12140, w12141, w12142, w12143, w12144, w12145, w12146, w12147, w12148, w12149, w12150, w12151, w12152, w12153, w12154, w12155, w12156, w12157, w12158, w12159, w12160, w12161, w12162, w12163, w12164, w12165, w12166, w12167, w12168, w12169, w12170, w12171, w12172, w12173, w12174, w12175, w12176, w12177, w12178, w12179, w12180, w12181, w12182, w12183, w12184, w12185, w12186, w12187, w12188, w12189, w12190, w12191, w12192, w12193, w12194, w12195, w12196, w12197, w12198, w12199, w12200, w12201, w12202, w12203, w12204, w12205, w12206, w12207, w12208, w12209, w12210, w12211, w12212, w12213, w12214, w12215, w12216, w12217, w12218, w12219, w12220, w12221, w12222, w12223, w12224, w12225, w12226, w12227, w12228, w12229, w12230, w12231, w12232, w12233, w12234, w12235, w12236, w12237, w12238, w12239, w12240, w12241, w12242, w12243, w12244, w12245, w12246, w12247, w12248, w12249, w12250, w12251, w12252, w12253, w12254, w12255, w12256, w12257, w12258, w12259, w12260, w12261, w12262, w12263, w12264, w12265, w12266, w12267, w12268, w12269, w12270, w12271, w12272, w12273, w12274, w12275, w12276, w12277, w12278, w12279, w12280, w12281, w12282, w12283, w12284, w12285, w12286, w12287, w12288, w12289, w12290, w12291, w12292, w12293, w12294, w12295, w12296, w12297, w12298, w12299, w12300, w12301, w12302, w12303, w12304, w12305, w12306, w12307, w12308, w12309, w12310, w12311, w12312, w12313, w12314, w12315, w12316, w12317, w12318, w12319, w12320, w12321, w12322, w12323, w12324, w12325, w12326, w12327, w12328, w12329, w12330, w12331, w12332, w12333, w12334, w12335, w12336, w12337, w12338, w12339, w12340, w12341, w12342, w12343, w12344, w12345, w12346, w12347, w12348, w12349, w12350, w12351, w12352, w12353, w12354, w12355, w12356, w12357, w12358, w12359, w12360, w12361, w12362, w12363, w12364, w12365, w12366, w12367, w12368, w12369, w12370, w12371, w12372, w12373, w12374, w12375, w12376, w12377, w12378, w12379, w12380, w12381, w12382, w12383, w12384, w12385, w12386, w12387, w12388, w12389, w12390, w12391, w12392, w12393, w12394, w12395, w12396, w12397, w12398, w12399, w12400, w12401, w12402, w12403, w12404, w12405, w12406, w12407, w12408, w12409, w12410, w12411, w12412, w12413, w12414, w12415, w12416, w12417, w12418, w12419, w12420, w12421, w12422, w12423, w12424, w12425, w12426, w12427, w12428, w12429, w12430, w12431, w12432, w12433, w12434, w12435, w12436, w12437, w12438, w12439, w12440, w12441, w12442, w12443, w12444, w12445, w12446, w12447, w12448, w12449, w12450, w12451, w12452, w12453, w12454, w12455, w12456, w12457, w12458, w12459, w12460, w12461, w12462, w12463, w12464, w12465, w12466, w12467, w12468, w12469, w12470, w12471, w12472, w12473, w12474, w12475, w12476, w12477, w12478, w12479, w12480, w12481, w12482, w12483, w12484, w12485, w12486, w12487, w12488, w12489, w12490, w12491, w12492, w12493, w12494, w12495, w12496, w12497, w12498, w12499, w12500, w12501, w12502, w12503, w12504, w12505, w12506, w12507, w12508, w12509, w12510, w12511, w12512, w12513, w12514, w12515, w12516, w12517, w12518, w12519, w12520, w12521, w12522, w12523, w12524, w12525, w12526, w12527, w12528, w12529, w12530, w12531, w12532, w12533, w12534, w12535, w12536, w12537, w12538, w12539, w12540, w12541, w12542, w12543, w12544, w12545, w12546, w12547, w12548, w12549, w12550, w12551, w12552, w12553, w12554, w12555, w12556, w12557, w12558, w12559, w12560, w12561, w12562, w12563, w12564, w12565, w12566, w12567, w12568, w12569, w12570, w12571, w12572, w12573, w12574, w12575, w12576, w12577, w12578, w12579, w12580, w12581, w12582, w12583, w12584, w12585, w12586, w12587, w12588, w12589, w12590, w12591, w12592, w12593, w12594, w12595, w12596, w12597, w12598, w12599, w12600, w12601, w12602, w12603, w12604, w12605, w12606, w12607, w12608, w12609, w12610, w12611, w12612, w12613, w12614, w12615, w12616, w12617, w12618, w12619, w12620, w12621, w12622, w12623, w12624, w12625, w12626, w12627, w12628, w12629, w12630, w12631, w12632, w12633, w12634, w12635, w12636, w12637, w12638, w12639, w12640, w12641, w12642, w12643, w12644, w12645, w12646, w12647, w12648, w12649, w12650, w12651, w12652, w12653, w12654, w12655, w12656, w12657, w12658, w12659, w12660, w12661, w12662, w12663, w12664, w12665, w12666, w12667, w12668, w12669, w12670, w12671, w12672, w12673, w12674, w12675, w12676, w12677, w12678, w12679, w12680, w12681, w12682, w12683, w12684, w12685, w12686, w12687, w12688, w12689, w12690, w12691, w12692, w12693, w12694, w12695, w12696, w12697, w12698, w12699, w12700, w12701, w12702, w12703, w12704, w12705, w12706, w12707, w12708, w12709, w12710, w12711, w12712, w12713, w12714, w12715, w12716, w12717, w12718, w12719, w12720, w12721, w12722, w12723, w12724, w12725, w12726, w12727, w12728, w12729, w12730, w12731, w12732, w12733, w12734, w12735, w12736, w12737, w12738, w12739, w12740, w12741, w12742, w12743, w12744, w12745, w12746, w12747, w12748, w12749, w12750, w12751, w12752, w12753, w12754, w12755, w12756, w12757, w12758, w12759, w12760, w12761, w12762, w12763, w12764, w12765, w12766, w12767, w12768, w12769, w12770, w12771, w12772, w12773, w12774, w12775, w12776, w12777, w12778, w12779, w12780, w12781, w12782, w12783, w12784, w12785, w12786, w12787, w12788, w12789, w12790, w12791, w12792, w12793, w12794, w12795, w12796, w12797, w12798, w12799, w12800, w12801, w12802, w12803, w12804, w12805, w12806, w12807, w12808, w12809, w12810, w12811, w12812, w12813, w12814, w12815, w12816, w12817, w12818, w12819, w12820, w12821, w12822, w12823, w12824, w12825, w12826, w12827, w12828, w12829, w12830, w12831, w12832, w12833, w12834, w12835, w12836, w12837, w12838, w12839, w12840, w12841, w12842, w12843, w12844, w12845, w12846, w12847, w12848, w12849, w12850, w12851, w12852, w12853, w12854, w12855, w12856, w12857, w12858, w12859, w12860, w12861, w12862, w12863, w12864, w12865, w12866, w12867, w12868, w12869, w12870, w12871, w12872, w12873, w12874, w12875, w12876, w12877, w12878, w12879, w12880, w12881, w12882, w12883, w12884, w12885, w12886, w12887, w12888, w12889, w12890, w12891, w12892, w12893, w12894, w12895, w12896, w12897, w12898, w12899, w12900, w12901, w12902, w12903, w12904, w12905, w12906, w12907, w12908, w12909, w12910, w12911, w12912, w12913, w12914, w12915, w12916, w12917, w12918, w12919, w12920, w12921, w12922, w12923, w12924, w12925, w12926, w12927, w12928, w12929, w12930, w12931, w12932, w12933, w12934, w12935, w12936, w12937, w12938, w12939, w12940, w12941, w12942, w12943, w12944, w12945, w12946, w12947, w12948, w12949, w12950, w12951, w12952, w12953, w12954, w12955, w12956, w12957, w12958, w12959, w12960, w12961, w12962, w12963, w12964, w12965, w12966, w12967, w12968, w12969, w12970, w12971, w12972, w12973, w12974, w12975, w12976, w12977, w12978, w12979, w12980, w12981, w12982, w12983, w12984, w12985, w12986, w12987, w12988, w12989, w12990, w12991, w12992, w12993, w12994;
assign w0 = ~pi0138 & pi1090;
assign w1 = ~pi1101 & w0;
assign w2 = ~pi1088 & ~pi1091;
assign w3 = ~pi0336 & ~pi0409;
assign w4 = ~pi0660 & w3;
assign w5 = w2 & w4;
assign w6 = w4 & w11198;
assign w7 = ~pi0309 & w6;
assign w8 = w6 & w11199;
assign w9 = pi1088 & pi1091;
assign w10 = ~pi0309 & ~pi1090;
assign w11 = ~pi1370 & w10;
assign w12 = w4 & ~w9;
assign w13 = w11 & w12;
assign w14 = w12 & w11200;
assign w15 = ~pi1101 & w14;
assign w16 = ~pi0196 & ~w8;
assign w17 = ~w15 & w16;
assign w18 = pi0646 & w17;
assign w19 = ~pi0634 & pi1688;
assign w20 = ~pi0702 & ~pi0716;
assign w21 = ~pi0677 & w20;
assign w22 = w20 & w11201;
assign w23 = pi0619 & pi1773;
assign w24 = w22 & w11202;
assign w25 = ~pi0619 & ~pi0634;
assign w26 = ~pi1401 & w25;
assign w27 = w25 & w11201;
assign w28 = pi0702 & ~pi0716;
assign w29 = ~pi0702 & pi0716;
assign w30 = ~w28 & ~w29;
assign w31 = ~pi0646 & ~w30;
assign w32 = w27 & w31;
assign w33 = ~w24 & ~w32;
assign w34 = w17 & ~w33;
assign w35 = ~w18 & ~w34;
assign w36 = pi1774 & ~w35;
assign w37 = pi0156 & w35;
assign w38 = ~w36 & ~w37;
assign w39 = pi1775 & ~w35;
assign w40 = pi0146 & w35;
assign w41 = ~w39 & ~w40;
assign w42 = pi1776 & ~w35;
assign w43 = pi0175 & w35;
assign w44 = ~w42 & ~w43;
assign w45 = pi1777 & ~w35;
assign w46 = pi0177 & w35;
assign w47 = ~w45 & ~w46;
assign w48 = pi1778 & ~w35;
assign w49 = pi0178 & w35;
assign w50 = ~w48 & ~w49;
assign w51 = pi1779 & ~w35;
assign w52 = pi0144 & w35;
assign w53 = ~w51 & ~w52;
assign w54 = pi1780 & ~w35;
assign w55 = pi0179 & w35;
assign w56 = ~w54 & ~w55;
assign w57 = pi1781 & ~w35;
assign w58 = pi0180 & w35;
assign w59 = ~w57 & ~w58;
assign w60 = pi1782 & ~w35;
assign w61 = pi0181 & w35;
assign w62 = ~w60 & ~w61;
assign w63 = pi1783 & ~w35;
assign w64 = pi0182 & w35;
assign w65 = ~w63 & ~w64;
assign w66 = pi1784 & ~w35;
assign w67 = pi0157 & w35;
assign w68 = ~w66 & ~w67;
assign w69 = pi1785 & ~w35;
assign w70 = pi0159 & w35;
assign w71 = ~w69 & ~w70;
assign w72 = pi1786 & ~w35;
assign w73 = pi0158 & w35;
assign w74 = ~w72 & ~w73;
assign w75 = pi1787 & ~w35;
assign w76 = pi0160 & w35;
assign w77 = ~w75 & ~w76;
assign w78 = pi1788 & ~w35;
assign w79 = pi0161 & w35;
assign w80 = ~w78 & ~w79;
assign w81 = pi1789 & ~w35;
assign w82 = pi0162 & w35;
assign w83 = ~w81 & ~w82;
assign w84 = pi1790 & ~w35;
assign w85 = pi0147 & w35;
assign w86 = ~w84 & ~w85;
assign w87 = pi1791 & ~w35;
assign w88 = pi0163 & w35;
assign w89 = ~w87 & ~w88;
assign w90 = pi1792 & ~w35;
assign w91 = pi0164 & w35;
assign w92 = ~w90 & ~w91;
assign w93 = pi1793 & ~w35;
assign w94 = pi0165 & w35;
assign w95 = ~w93 & ~w94;
assign w96 = pi1794 & ~w35;
assign w97 = pi0166 & w35;
assign w98 = ~w96 & ~w97;
assign w99 = pi1795 & ~w35;
assign w100 = pi0167 & w35;
assign w101 = ~w99 & ~w100;
assign w102 = pi1796 & ~w35;
assign w103 = pi0168 & w35;
assign w104 = ~w102 & ~w103;
assign w105 = pi1797 & ~w35;
assign w106 = pi0169 & w35;
assign w107 = ~w105 & ~w106;
assign w108 = pi1798 & ~w35;
assign w109 = pi0170 & w35;
assign w110 = ~w108 & ~w109;
assign w111 = pi1799 & ~w35;
assign w112 = pi0171 & w35;
assign w113 = ~w111 & ~w112;
assign w114 = pi1800 & ~w35;
assign w115 = pi0172 & w35;
assign w116 = ~w114 & ~w115;
assign w117 = pi1801 & ~w35;
assign w118 = pi0145 & w35;
assign w119 = ~w117 & ~w118;
assign w120 = pi1802 & ~w35;
assign w121 = pi0173 & w35;
assign w122 = ~w120 & ~w121;
assign w123 = pi1803 & ~w35;
assign w124 = pi0174 & w35;
assign w125 = ~w123 & ~w124;
assign w126 = pi1804 & ~w35;
assign w127 = pi0141 & w35;
assign w128 = ~w126 & ~w127;
assign w129 = pi1805 & ~w35;
assign w130 = pi0176 & w35;
assign w131 = ~w129 & ~w130;
assign w132 = pi1038 & pi1683;
assign w133 = ~pi1858 & pi1859;
assign w134 = ~w132 & ~w133;
assign w135 = ~pi1669 & ~w17;
assign w136 = ~pi0716 & pi1748;
assign w137 = ~pi0702 & ~w136;
assign w138 = w17 & w11203;
assign w139 = ~w135 & ~w138;
assign w140 = pi1758 & ~w35;
assign w141 = pi0038 & w35;
assign w142 = ~w140 & ~w141;
assign w143 = pi1759 & ~w35;
assign w144 = pi0044 & w35;
assign w145 = ~w143 & ~w144;
assign w146 = pi1760 & ~w35;
assign w147 = pi0040 & w35;
assign w148 = ~w146 & ~w147;
assign w149 = pi1761 & ~w35;
assign w150 = pi0039 & w35;
assign w151 = ~w149 & ~w150;
assign w152 = pi1762 & ~w35;
assign w153 = pi0041 & w35;
assign w154 = ~w152 & ~w153;
assign w155 = pi1763 & ~w35;
assign w156 = pi0034 & w35;
assign w157 = ~w155 & ~w156;
assign w158 = pi1764 & ~w35;
assign w159 = pi0035 & w35;
assign w160 = ~w158 & ~w159;
assign w161 = pi1765 & ~w35;
assign w162 = pi0036 & w35;
assign w163 = ~w161 & ~w162;
assign w164 = pi1766 & ~w35;
assign w165 = pi0037 & w35;
assign w166 = ~w164 & ~w165;
assign w167 = pi1767 & ~w35;
assign w168 = pi0045 & w35;
assign w169 = ~w167 & ~w168;
assign w170 = pi1768 & ~w35;
assign w171 = pi0042 & w35;
assign w172 = ~w170 & ~w171;
assign w173 = pi1769 & ~w35;
assign w174 = pi0031 & w35;
assign w175 = ~w173 & ~w174;
assign w176 = pi1770 & ~w35;
assign w177 = pi0043 & w35;
assign w178 = ~w176 & ~w177;
assign w179 = pi1771 & ~w35;
assign w180 = pi0032 & w35;
assign w181 = ~w179 & ~w180;
assign w182 = pi1772 & ~w35;
assign w183 = pi0033 & w35;
assign w184 = ~w182 & ~w183;
assign w185 = ~pi0096 & ~pi1018;
assign w186 = pi0093 & w185;
assign w187 = (pi0068 & ~w185) | (pi0068 & w11204) | (~w185 & w11204);
assign w188 = ~pi1753 & ~w187;
assign w189 = ~pi0065 & pi0093;
assign w190 = (~w189 & w187) | (~w189 & w11205) | (w187 & w11205);
assign w191 = ~pi0005 & w190;
assign w192 = w190 & w11206;
assign w193 = ~w187 & w11208;
assign w194 = pi0005 & w190;
assign w195 = w190 & w11209;
assign w196 = (w189 & w187) | (w189 & w11210) | (w187 & w11210);
assign w197 = ~pi0059 & ~pi0061;
assign w198 = ~pi0055 & ~pi1429;
assign w199 = pi1422 & w197;
assign w200 = w198 & w199;
assign w201 = w199 & w11211;
assign w202 = ~pi1422 & w197;
assign w203 = ~pi0055 & pi1429;
assign w204 = w202 & w203;
assign w205 = ~w201 & ~w204;
assign w206 = pi0058 & pi1692;
assign w207 = w185 & w206;
assign w208 = pi0055 & ~pi1429;
assign w209 = w202 & w208;
assign w210 = w207 & w209;
assign w211 = w199 & w11212;
assign w212 = ~pi1422 & w198;
assign w213 = ~pi0059 & pi0061;
assign w214 = w212 & w213;
assign w215 = ~w210 & w11213;
assign w216 = pi0059 & ~pi0061;
assign w217 = w212 & w11214;
assign w218 = w215 & w11215;
assign w219 = pi0152 & pi0874;
assign w220 = pi0055 & pi0152;
assign w221 = w206 & w220;
assign w222 = ~w219 & ~w221;
assign w223 = ~w221 & w11216;
assign w224 = pi0055 & w206;
assign w225 = (~pi0874 & ~w206) | (~pi0874 & w11217) | (~w206 & w11217);
assign w226 = pi0152 & pi0199;
assign w227 = ~w225 & w226;
assign w228 = ~w223 & ~w227;
assign w229 = pi0193 & ~w226;
assign w230 = pi0193 & ~pi0874;
assign w231 = ~w224 & w230;
assign w232 = ~w229 & ~w231;
assign w233 = ~pi0193 & w226;
assign w234 = ~w225 & w233;
assign w235 = w232 & ~w234;
assign w236 = ~w235 & w11218;
assign w237 = ~pi0152 & w225;
assign w238 = w222 & ~w237;
assign w239 = ~w223 & ~w232;
assign w240 = ~w232 & w11219;
assign w241 = w228 & w11220;
assign w242 = ~w228 & w235;
assign w243 = w235 & w11221;
assign w244 = ~w238 & ~w240;
assign w245 = ~w236 & w244;
assign w246 = ~w241 & ~w243;
assign w247 = w245 & w246;
assign w248 = ~w235 & w11222;
assign w249 = ~w232 & w11223;
assign w250 = w228 & w11224;
assign w251 = w235 & w11225;
assign w252 = w238 & ~w249;
assign w253 = ~w248 & w252;
assign w254 = ~w250 & ~w251;
assign w255 = w253 & w254;
assign w256 = ~w247 & ~w255;
assign w257 = pi1422 & pi1692;
assign w258 = (~w257 & ~w202) | (~w257 & w11226) | (~w202 & w11226);
assign w259 = pi0052 & ~w258;
assign w260 = ~pi0982 & w217;
assign w261 = w215 & w11227;
assign w262 = (~w259 & w215) | (~w259 & w11228) | (w215 & w11228);
assign w263 = ~w261 & w262;
assign w264 = w196 & ~w263;
assign w265 = (w264 & w256) | (w264 & w11229) | (w256 & w11229);
assign w266 = ~w192 & ~w193;
assign w267 = ~w195 & w266;
assign w268 = ~w265 & w267;
assign w269 = w190 & w11230;
assign w270 = ~w232 & w11231;
assign w271 = w235 & w11232;
assign w272 = w228 & w11233;
assign w273 = ~w235 & w11234;
assign w274 = ~w238 & ~w270;
assign w275 = ~w271 & w274;
assign w276 = ~w272 & ~w273;
assign w277 = w275 & w276;
assign w278 = ~w232 & w11235;
assign w279 = w235 & w11236;
assign w280 = w228 & w11237;
assign w281 = ~w235 & w11238;
assign w282 = w238 & ~w278;
assign w283 = ~w279 & w282;
assign w284 = ~w280 & ~w281;
assign w285 = w283 & w284;
assign w286 = ~w277 & ~w285;
assign w287 = ~pi0013 & ~w258;
assign w288 = (~w287 & w215) | (~w287 & w11239) | (w215 & w11239);
assign w289 = ~w261 & w288;
assign w290 = (~w289 & ~w286) | (~w289 & w11240) | (~w286 & w11240);
assign w291 = w196 & ~w290;
assign w292 = ~w187 & w11241;
assign w293 = w190 & w11242;
assign w294 = ~w269 & ~w292;
assign w295 = ~w293 & w294;
assign w296 = ~w291 & w295;
assign w297 = ~w187 & w11243;
assign w298 = ~w232 & w11244;
assign w299 = ~w235 & w11245;
assign w300 = w228 & w11246;
assign w301 = w235 & w11247;
assign w302 = ~w238 & ~w298;
assign w303 = ~w299 & w302;
assign w304 = ~w300 & ~w301;
assign w305 = w303 & w304;
assign w306 = ~w232 & w11248;
assign w307 = ~w235 & w11249;
assign w308 = w228 & w11250;
assign w309 = w235 & w11251;
assign w310 = w238 & ~w306;
assign w311 = ~w307 & w310;
assign w312 = ~w308 & ~w309;
assign w313 = w311 & w312;
assign w314 = ~w305 & ~w313;
assign w315 = ~pi1016 & w217;
assign w316 = w215 & w11252;
assign w317 = pi0060 & ~w258;
assign w318 = (~w317 & w215) | (~w317 & w11253) | (w215 & w11253);
assign w319 = ~w316 & w318;
assign w320 = w196 & ~w319;
assign w321 = (w320 & w314) | (w320 & w11254) | (w314 & w11254);
assign w322 = ~w191 & ~w297;
assign w323 = ~w321 & w322;
assign w324 = ~w187 & w11255;
assign w325 = ~w235 & w11256;
assign w326 = ~w232 & w11257;
assign w327 = w228 & w11258;
assign w328 = w235 & w11259;
assign w329 = w238 & ~w326;
assign w330 = ~w325 & w329;
assign w331 = ~w327 & ~w328;
assign w332 = w330 & w331;
assign w333 = ~w235 & w11260;
assign w334 = ~w232 & w11261;
assign w335 = w228 & w11262;
assign w336 = w235 & w11263;
assign w337 = ~w238 & ~w334;
assign w338 = ~w333 & w337;
assign w339 = ~w335 & ~w336;
assign w340 = w338 & w339;
assign w341 = ~w332 & ~w340;
assign w342 = ~pi0010 & ~w258;
assign w343 = (~w342 & w215) | (~w342 & w11264) | (w215 & w11264);
assign w344 = ~w316 & w343;
assign w345 = (~w344 & ~w341) | (~w344 & w11265) | (~w341 & w11265);
assign w346 = w196 & ~w345;
assign w347 = ~w194 & ~w324;
assign w348 = ~w346 & w347;
assign w349 = pi0110 & ~pi0138;
assign w350 = ~pi0725 & ~pi0743;
assign w351 = pi0006 & pi0008;
assign w352 = ~pi0625 & pi1479;
assign w353 = w351 & w352;
assign w354 = (w349 & w353) | (w349 & w11266) | (w353 & w11266);
assign w355 = pi1227 & ~pi1228;
assign w356 = pi1229 & ~pi1236;
assign w357 = w355 & w356;
assign w358 = pi0352 & ~w357;
assign w359 = ~pi0780 & pi0798;
assign w360 = ~w357 & w11267;
assign w361 = ~pi0092 & ~pi0108;
assign w362 = ~pi0088 & ~pi0112;
assign w363 = ~pi0110 & w362;
assign w364 = w362 & w11268;
assign w365 = ~pi0095 & w364;
assign w366 = w364 & w11269;
assign w367 = w366 & w11270;
assign w368 = w360 & w367;
assign w369 = pi0780 & ~pi0798;
assign w370 = ~pi0771 & ~pi0801;
assign w371 = ~pi1229 & w355;
assign w372 = w355 & w11271;
assign w373 = w370 & w372;
assign w374 = ~pi0771 & pi0801;
assign w375 = ~pi0385 & w374;
assign w376 = pi0771 & ~pi0801;
assign w377 = ~pi0125 & w376;
assign w378 = ~w375 & ~w377;
assign w379 = (~pi1470 & w378) | (~pi1470 & w11272) | (w378 & w11272);
assign w380 = ~w373 & w379;
assign w381 = w355 & w1709;
assign w382 = w370 & w381;
assign w383 = (~pi1471 & w378) | (~pi1471 & w393) | (w378 & w393);
assign w384 = ~w382 & w383;
assign w385 = ~w380 & ~w384;
assign w386 = w385 & w11273;
assign w387 = ~w354 & ~w386;
assign w388 = w367 & w11274;
assign w389 = w349 & w350;
assign w390 = w353 & w389;
assign w391 = ~w388 & ~w390;
assign w392 = ~pi0767 & ~pi1470;
assign w393 = ~pi0796 & ~pi1471;
assign w394 = ~w392 & w393;
assign w395 = ~w370 & ~w394;
assign w396 = ~pi1458 & w370;
assign w397 = ~w395 & ~w396;
assign w398 = pi0796 & ~w370;
assign w399 = (pi0024 & w370) | (pi0024 & w11275) | (w370 & w11275);
assign w400 = (w399 & w395) | (w399 & w11276) | (w395 & w11276);
assign w401 = ~w395 & w11277;
assign w402 = w379 & ~w400;
assign w403 = ~w401 & w402;
assign w404 = pi0796 & w376;
assign w405 = ~pi0801 & ~pi1458;
assign w406 = ~pi0771 & ~w405;
assign w407 = ~w404 & ~w406;
assign w408 = pi0237 & w407;
assign w409 = w376 & w11278;
assign w410 = ~w405 & w11279;
assign w411 = ~w409 & ~w410;
assign w412 = (pi0946 & w408) | (pi0946 & w11280) | (w408 & w11280);
assign w413 = ~w408 & w11281;
assign w414 = pi0257 & w407;
assign w415 = w376 & w11282;
assign w416 = ~w405 & w11283;
assign w417 = ~w415 & ~w416;
assign w418 = ~w414 & w417;
assign w419 = (~pi0895 & w414) | (~pi0895 & w11284) | (w414 & w11284);
assign w420 = ~w413 & w419;
assign w421 = (pi0940 & w420) | (pi0940 & w11285) | (w420 & w11285);
assign w422 = ~pi0940 & ~w412;
assign w423 = ~w420 & w422;
assign w424 = w376 & w11286;
assign w425 = (~w424 & ~w407) | (~w424 & w11287) | (~w407 & w11287);
assign w426 = pi0150 & w406;
assign w427 = w425 & ~w426;
assign w428 = ~w423 & ~w427;
assign w429 = w376 & w11288;
assign w430 = (~w429 & ~w407) | (~w429 & w11289) | (~w407 & w11289);
assign w431 = pi0188 & w406;
assign w432 = (pi0742 & ~w430) | (pi0742 & w11290) | (~w430 & w11290);
assign w433 = w376 & w11291;
assign w434 = (~w433 & ~w407) | (~w433 & w11292) | (~w407 & w11292);
assign w435 = pi0149 & w406;
assign w436 = w434 & w11293;
assign w437 = (pi0741 & ~w434) | (pi0741 & w11294) | (~w434 & w11294);
assign w438 = ~w436 & ~w437;
assign w439 = ~w432 & w438;
assign w440 = ~w428 & w11295;
assign w441 = w430 & w11296;
assign w442 = ~w432 & w436;
assign w443 = ~w441 & ~w442;
assign w444 = (~pi0945 & w440) | (~pi0945 & w11297) | (w440 & w11297);
assign w445 = w376 & w11298;
assign w446 = (~w445 & ~w407) | (~w445 & w11299) | (~w407 & w11299);
assign w447 = pi0151 & w406;
assign w448 = w446 & ~w447;
assign w449 = (~w440 & w11300) | (~w440 & w11301) | (w11300 & w11301);
assign w450 = w376 & w11302;
assign w451 = (~w450 & ~w407) | (~w450 & w11303) | (~w407 & w11303);
assign w452 = pi0133 & w406;
assign w453 = w451 & w11304;
assign w454 = (pi0867 & ~w451) | (pi0867 & w11305) | (~w451 & w11305);
assign w455 = ~w453 & ~w454;
assign w456 = ~w440 & w11306;
assign w457 = w455 & ~w456;
assign w458 = w376 & w11307;
assign w459 = (~w458 & ~w407) | (~w458 & w11308) | (~w407 & w11308);
assign w460 = pi0189 & w406;
assign w461 = w459 & w11309;
assign w462 = ~w405 & w11310;
assign w463 = ~pi0864 & ~w462;
assign w464 = ~w461 & ~w463;
assign w465 = w376 & w11311;
assign w466 = (~w465 & ~w407) | (~w465 & w11312) | (~w407 & w11312);
assign w467 = pi0134 & w406;
assign w468 = w466 & w11313;
assign w469 = w376 & w11314;
assign w470 = (~w469 & ~w407) | (~w469 & w11315) | (~w407 & w11315);
assign w471 = pi0132 & w406;
assign w472 = (pi0868 & ~w470) | (pi0868 & w11316) | (~w470 & w11316);
assign w473 = w470 & w11317;
assign w474 = ~w472 & ~w473;
assign w475 = ~w453 & w474;
assign w476 = w376 & w11318;
assign w477 = (~w476 & ~w407) | (~w476 & w11319) | (~w407 & w11319);
assign w478 = pi0135 & w406;
assign w479 = (pi0875 & ~w477) | (pi0875 & w11320) | (~w477 & w11320);
assign w480 = w477 & w11321;
assign w481 = ~w479 & ~w480;
assign w482 = ~w468 & w481;
assign w483 = w475 & w482;
assign w484 = w464 & w483;
assign w485 = (w484 & ~w457) | (w484 & w11322) | (~w457 & w11322);
assign w486 = (pi0869 & ~w466) | (pi0869 & w11323) | (~w466 & w11323);
assign w487 = ~w472 & ~w486;
assign w488 = ~w468 & ~w487;
assign w489 = w481 & w488;
assign w490 = w488 & w11324;
assign w491 = pi0864 & w462;
assign w492 = (pi0739 & ~w459) | (pi0739 & w11325) | (~w459 & w11325);
assign w493 = ~w479 & ~w492;
assign w494 = w464 & ~w493;
assign w495 = ~w491 & ~w494;
assign w496 = ~w405 & w11327;
assign w497 = pi0774 & ~w496;
assign w498 = ~pi0815 & pi1099;
assign w499 = (~w498 & w496) | (~w498 & w11328) | (w496 & w11328);
assign w500 = ~pi0774 & w496;
assign w501 = ~w405 & w11330;
assign w502 = pi0740 & w501;
assign w503 = ~pi0740 & ~w501;
assign w504 = ~w502 & ~w503;
assign w505 = w504 & w11331;
assign w506 = ~w498 & ~w505;
assign w507 = (~w485 & w11332) | (~w485 & w11333) | (w11332 & w11333);
assign w508 = ~w497 & ~w500;
assign w509 = (~pi1099 & w496) | (~pi1099 & w11335) | (w496 & w11335);
assign w510 = ~w504 & w509;
assign w511 = (w510 & w485) | (w510 & w11336) | (w485 & w11336);
assign w512 = ~w507 & ~w511;
assign w513 = ~w395 & w11337;
assign w514 = (pi0672 & w395) | (pi0672 & w11338) | (w395 & w11338);
assign w515 = ~pi1471 & ~w513;
assign w516 = ~w514 & w515;
assign w517 = ~pi0778 & ~w314;
assign w518 = pi0778 & w314;
assign w519 = ~w517 & ~w518;
assign w520 = ~w235 & w11339;
assign w521 = ~w232 & w11340;
assign w522 = w228 & w11341;
assign w523 = w235 & w11342;
assign w524 = w238 & ~w521;
assign w525 = ~w520 & w524;
assign w526 = ~w522 & ~w523;
assign w527 = w525 & w526;
assign w528 = ~w235 & w11343;
assign w529 = ~w232 & w11344;
assign w530 = w228 & w11345;
assign w531 = w235 & w11346;
assign w532 = ~w238 & ~w529;
assign w533 = ~w528 & w532;
assign w534 = ~w530 & ~w531;
assign w535 = w533 & w534;
assign w536 = ~w527 & ~w535;
assign w537 = ~pi0878 & ~w536;
assign w538 = pi0878 & w536;
assign w539 = ~w537 & ~w538;
assign w540 = ~pi0779 & ~w256;
assign w541 = pi0779 & w256;
assign w542 = ~w540 & ~w541;
assign w543 = w539 & ~w542;
assign w544 = ~w539 & w542;
assign w545 = ~w543 & ~w544;
assign w546 = w519 & w545;
assign w547 = ~w519 & ~w545;
assign w548 = ~w546 & ~w547;
assign w549 = w235 & w11347;
assign w550 = ~w232 & w11348;
assign w551 = ~w235 & w11349;
assign w552 = w228 & w11350;
assign w553 = ~w238 & ~w550;
assign w554 = ~w549 & w553;
assign w555 = ~w551 & ~w552;
assign w556 = w554 & w555;
assign w557 = w235 & w11351;
assign w558 = ~w232 & w11352;
assign w559 = ~w235 & w11353;
assign w560 = w228 & w11354;
assign w561 = w238 & ~w558;
assign w562 = ~w557 & w561;
assign w563 = ~w559 & ~w560;
assign w564 = w562 & w563;
assign w565 = ~w556 & ~w564;
assign w566 = ~pi0009 & ~w565;
assign w567 = pi0009 & w565;
assign w568 = ~w566 & ~w567;
assign w569 = w235 & w11355;
assign w570 = ~w232 & w11356;
assign w571 = ~w235 & w11357;
assign w572 = w228 & w11358;
assign w573 = w238 & ~w570;
assign w574 = ~w569 & w573;
assign w575 = ~w571 & ~w572;
assign w576 = w574 & w575;
assign w577 = w235 & w11359;
assign w578 = ~w232 & w11360;
assign w579 = ~w235 & w11361;
assign w580 = w228 & w11362;
assign w581 = ~w238 & ~w578;
assign w582 = ~w577 & w581;
assign w583 = ~w579 & ~w580;
assign w584 = w582 & w583;
assign w585 = ~w576 & ~w584;
assign w586 = ~pi0747 & ~w585;
assign w587 = pi0747 & w585;
assign w588 = ~w586 & ~w587;
assign w589 = w568 & ~w588;
assign w590 = ~w568 & w588;
assign w591 = ~w589 & ~w590;
assign w592 = ~pi0054 & ~w341;
assign w593 = pi0054 & w341;
assign w594 = ~w592 & ~w593;
assign w595 = ~w235 & w11363;
assign w596 = ~w232 & w11364;
assign w597 = w228 & w11365;
assign w598 = w235 & w11366;
assign w599 = w238 & ~w596;
assign w600 = ~w595 & w599;
assign w601 = ~w597 & ~w598;
assign w602 = w600 & w601;
assign w603 = ~w235 & w11367;
assign w604 = w228 & w11368;
assign w605 = (~w238 & ~w239) | (~w238 & w11369) | (~w239 & w11369);
assign w606 = ~w603 & w605;
assign w607 = (~w604 & ~w242) | (~w604 & w11370) | (~w242 & w11370);
assign w608 = w606 & w607;
assign w609 = ~w602 & ~w608;
assign w610 = ~pi0777 & ~w609;
assign w611 = pi0777 & w609;
assign w612 = ~w610 & ~w611;
assign w613 = w594 & ~w612;
assign w614 = ~w594 & w612;
assign w615 = ~w613 & ~w614;
assign w616 = w591 & w615;
assign w617 = ~w591 & ~w615;
assign w618 = ~w616 & ~w617;
assign w619 = w548 & w618;
assign w620 = ~w548 & ~w618;
assign w621 = ~w619 & ~w620;
assign w622 = ~pi0066 & pi1542;
assign w623 = ~pi1625 & w622;
assign w624 = (~w623 & ~w215) | (~w623 & w11371) | (~w215 & w11371);
assign w625 = ~w621 & ~w624;
assign w626 = ~pi0025 & ~w286;
assign w627 = pi0025 & w286;
assign w628 = ~w626 & ~w627;
assign w629 = ~pi0053 & ~w628;
assign w630 = pi0053 & w628;
assign w631 = ~w629 & ~w630;
assign w632 = ~w621 & w11372;
assign w633 = ~w624 & ~w631;
assign w634 = pi1625 & ~w185;
assign w635 = (w215 & w11375) | (w215 & w11376) | (w11375 & w11376);
assign w636 = (w635 & ~w621) | (w635 & w12976) | (~w621 & w12976);
assign w637 = ~w632 & w636;
assign w638 = (w215 & w11379) | (w215 & w11380) | (w11379 & w11380);
assign w639 = ~w625 & w638;
assign w640 = (~w503 & ~w504) | (~w503 & w11381) | (~w504 & w11381);
assign w641 = w495 & ~w640;
assign w642 = ~w485 & w11382;
assign w643 = w497 & ~w502;
assign w644 = ~w503 & ~w643;
assign w645 = ~pi0870 & pi1099;
assign w646 = ~pi0865 & ~w645;
assign w647 = (~w485 & w11384) | (~w485 & w11385) | (w11384 & w11385);
assign w648 = ~pi1099 & w641;
assign w649 = ~w485 & w11386;
assign w650 = pi0865 & w644;
assign w651 = (w644 & w11388) | (w644 & w11389) | (w11388 & w11389);
assign w652 = ~w649 & w651;
assign w653 = ~w647 & ~w652;
assign w654 = (pi0024 & w405) | (pi0024 & w11390) | (w405 & w11390);
assign w655 = ~w405 & w11391;
assign w656 = ~w654 & ~w655;
assign w657 = ~w621 & w11392;
assign w658 = ~w624 & ~w628;
assign w659 = (w215 & w11395) | (w215 & w11396) | (w11395 & w11396);
assign w660 = (w659 & ~w621) | (w659 & w12977) | (~w621 & w12977);
assign w661 = ~w657 & w660;
assign w662 = pi0814 & pi1099;
assign w663 = ~w500 & w509;
assign w664 = (w663 & w485) | (w663 & w11397) | (w485 & w11397);
assign w665 = ~pi1099 & ~w508;
assign w666 = ~w485 & w11398;
assign w667 = ~w662 & ~w664;
assign w668 = ~w666 & w667;
assign w669 = (~pi1099 & ~w644) | (~pi1099 & w11400) | (~w644 & w11400);
assign w670 = pi0817 & pi1099;
assign w671 = ~pi0775 & ~pi1099;
assign w672 = ~w670 & ~w671;
assign w673 = ~w649 & w11401;
assign w674 = (pi0775 & w649) | (pi0775 & w11402) | (w649 & w11402);
assign w675 = ~w673 & ~w674;
assign w676 = pi0812 & pi1099;
assign w677 = (w483 & ~w457) | (w483 & w11403) | (~w457 & w11403);
assign w678 = ~w489 & ~w677;
assign w679 = ~w461 & ~w492;
assign w680 = ~pi1099 & ~w679;
assign w681 = ~w677 & w11405;
assign w682 = ~pi1099 & w679;
assign w683 = (w682 & w677) | (w682 & w11406) | (w677 & w11406);
assign w684 = ~w676 & ~w681;
assign w685 = ~w683 & w684;
assign w686 = ~w187 & w11407;
assign w687 = pi0051 & ~w205;
assign w688 = ~pi0878 & ~w215;
assign w689 = ~w687 & ~w688;
assign w690 = (w689 & ~w536) | (w689 & w11408) | (~w536 & w11408);
assign w691 = ~w188 & ~w690;
assign w692 = ~w190 & ~w686;
assign w693 = ~w691 & w692;
assign w694 = ~pi0816 & pi1099;
assign w695 = ~w649 & w11409;
assign w696 = ~pi0866 & ~w694;
assign w697 = (w696 & w642) | (w696 & w11410) | (w642 & w11410);
assign w698 = ~w695 & ~w697;
assign w699 = (~w461 & w677) | (~w461 & w11412) | (w677 & w11412);
assign w700 = ~w463 & ~w491;
assign w701 = ~pi0813 & pi1099;
assign w702 = (~w701 & w700) | (~w701 & w11413) | (w700 & w11413);
assign w703 = w699 & ~w702;
assign w704 = (~w701 & ~w700) | (~w701 & w11413) | (~w700 & w11413);
assign w705 = ~w699 & ~w704;
assign w706 = ~w703 & ~w705;
assign w707 = ~w187 & w11414;
assign w708 = pi0747 & ~w215;
assign w709 = (~w188 & w205) | (~w188 & w11415) | (w205 & w11415);
assign w710 = ~w708 & w709;
assign w711 = (w710 & w585) | (w710 & w11416) | (w585 & w11416);
assign w712 = ~w190 & ~w707;
assign w713 = ~w711 & w712;
assign w714 = ~w187 & w11417;
assign w715 = pi0009 & ~w215;
assign w716 = (w196 & w205) | (w196 & w11418) | (w205 & w11418);
assign w717 = ~w715 & w716;
assign w718 = (w717 & w565) | (w717 & w11419) | (w565 & w11419);
assign w719 = ~w714 & ~w718;
assign w720 = ~pi0834 & pi1099;
assign w721 = (w475 & ~w457) | (w475 & w11420) | (~w457 & w11420);
assign w722 = ~w481 & ~w488;
assign w723 = (w722 & ~w721) | (w722 & w11421) | (~w721 & w11421);
assign w724 = ~pi1099 & w678;
assign w725 = ~w723 & w724;
assign w726 = ~w720 & ~w725;
assign w727 = pi0832 & pi1099;
assign w728 = ~w449 & ~w456;
assign w729 = ~w455 & ~w728;
assign w730 = (~pi1099 & ~w457) | (~pi1099 & w11422) | (~w457 & w11422);
assign w731 = ~w729 & w730;
assign w732 = ~w727 & ~w731;
assign w733 = pi0280 & pi0759;
assign w734 = pi0218 & pi0877;
assign w735 = ~pi0280 & ~pi0759;
assign w736 = ~pi0353 & ~pi0810;
assign w737 = pi0355 & pi0809;
assign w738 = pi0353 & pi0810;
assign w739 = ~pi0355 & ~pi0809;
assign w740 = ~pi0431 & ~pi0808;
assign w741 = ~pi0333 & pi0755;
assign w742 = pi0431 & pi0808;
assign w743 = pi0333 & ~pi0755;
assign w744 = pi0620 & ~pi0807;
assign w745 = pi0545 & pi0806;
assign w746 = ~pi0620 & pi0807;
assign w747 = ~pi0545 & ~pi0806;
assign w748 = ~pi0673 & ~pi0804;
assign w749 = pi0726 & pi0750;
assign w750 = pi0673 & pi0804;
assign w751 = ~pi0726 & ~pi0750;
assign w752 = pi0859 & ~pi1358;
assign w753 = ~w751 & w752;
assign w754 = ~w749 & ~w750;
assign w755 = ~w753 & w754;
assign w756 = ~w747 & ~w748;
assign w757 = ~w745 & ~w746;
assign w758 = (w757 & w755) | (w757 & w11423) | (w755 & w11423);
assign w759 = ~w743 & ~w744;
assign w760 = ~w741 & ~w742;
assign w761 = ~w739 & ~w740;
assign w762 = (~w758 & w11425) | (~w758 & w11426) | (w11425 & w11426);
assign w763 = ~w737 & ~w738;
assign w764 = ~w735 & ~w736;
assign w765 = ~w733 & ~w734;
assign w766 = (~w762 & w11428) | (~w762 & w11429) | (w11428 & w11429);
assign w767 = ~pi0218 & ~pi0877;
assign w768 = pi0086 & pi0200;
assign w769 = pi0281 & w768;
assign w770 = ~w767 & w769;
assign w771 = ~w766 & w770;
assign w772 = pi0013 & ~w591;
assign w773 = ~pi0013 & w591;
assign w774 = ~w772 & ~w773;
assign w775 = ~w624 & ~w774;
assign w776 = (w215 & w11432) | (w215 & w11433) | (w11432 & w11433);
assign w777 = ~w775 & w776;
assign w778 = ~w187 & w11434;
assign w779 = ~pi0777 & ~w215;
assign w780 = pi0050 & ~w205;
assign w781 = ~w779 & ~w780;
assign w782 = (w781 & ~w609) | (w781 & w11435) | (~w609 & w11435);
assign w783 = w196 & ~w782;
assign w784 = ~w778 & ~w783;
assign w785 = ~w468 & ~w486;
assign w786 = ~w721 & w11436;
assign w787 = (~w785 & w721) | (~w785 & w11437) | (w721 & w11437);
assign w788 = ~w786 & ~w787;
assign w789 = ~pi1099 & ~w788;
assign w790 = ~pi0833 & pi1099;
assign w791 = ~w789 & ~w790;
assign w792 = ~w444 & ~w456;
assign w793 = ~w448 & ~w792;
assign w794 = w448 & w792;
assign w795 = ~w793 & ~w794;
assign w796 = ~pi1099 & ~w795;
assign w797 = ~pi0831 & pi1099;
assign w798 = ~w796 & ~w797;
assign w799 = pi0218 & pi0280;
assign w800 = ~pi0333 & pi0353;
assign w801 = pi0355 & pi0431;
assign w802 = pi0545 & ~pi0620;
assign w803 = pi0673 & pi0726;
assign w804 = ~pi1358 & w803;
assign w805 = w801 & w802;
assign w806 = w799 & w800;
assign w807 = w805 & w806;
assign w808 = w769 & w804;
assign w809 = w807 & w808;
assign w810 = pi0757 & pi1099;
assign w811 = (~w453 & ~w457) | (~w453 & w11438) | (~w457 & w11438);
assign w812 = ~w474 & ~w811;
assign w813 = (~pi1099 & w812) | (~pi1099 & w11439) | (w812 & w11439);
assign w814 = ~w810 & ~w813;
assign w815 = ~pi0097 & ~pi0121;
assign w816 = pi1001 & ~w815;
assign w817 = pi0038 & pi1101;
assign w818 = pi1579 & w817;
assign w819 = w817 & w11440;
assign w820 = pi0040 & w819;
assign w821 = w819 & w11441;
assign w822 = w819 & w11442;
assign w823 = pi0034 & w822;
assign w824 = w822 & w11443;
assign w825 = w822 & w11444;
assign w826 = w822 & w11445;
assign w827 = pi0045 & w826;
assign w828 = w826 & w11446;
assign w829 = w826 & w11447;
assign w830 = (~pi0031 & ~w826) | (~pi0031 & w11448) | (~w826 & w11448);
assign w831 = ~w829 & ~w830;
assign w832 = pi1101 & pi1579;
assign w833 = ~pi0038 & ~w832;
assign w834 = ~w818 & ~w833;
assign w835 = pi0701 & ~w834;
assign w836 = ~pi0701 & w834;
assign w837 = ~w835 & ~w836;
assign w838 = (~pi0044 & ~w817) | (~pi0044 & w11449) | (~w817 & w11449);
assign w839 = ~w819 & ~w838;
assign w840 = pi0361 & ~w839;
assign w841 = ~pi0361 & w839;
assign w842 = ~w840 & ~w841;
assign w843 = ~pi0040 & ~w819;
assign w844 = ~w820 & ~w843;
assign w845 = pi0260 & ~w844;
assign w846 = ~pi0260 & w844;
assign w847 = ~w845 & ~w846;
assign w848 = (~pi0039 & ~w819) | (~pi0039 & w11450) | (~w819 & w11450);
assign w849 = ~w821 & ~w848;
assign w850 = pi0282 & ~w849;
assign w851 = ~pi0282 & w849;
assign w852 = ~w850 & ~w851;
assign w853 = (~pi0041 & ~w819) | (~pi0041 & w11451) | (~w819 & w11451);
assign w854 = ~w822 & ~w853;
assign w855 = pi0215 & ~w854;
assign w856 = ~pi0215 & w854;
assign w857 = ~w855 & ~w856;
assign w858 = ~pi0034 & ~w822;
assign w859 = ~w823 & ~w858;
assign w860 = pi0216 & ~w859;
assign w861 = ~pi0216 & w859;
assign w862 = ~w860 & ~w861;
assign w863 = (~pi0035 & ~w822) | (~pi0035 & w11452) | (~w822 & w11452);
assign w864 = ~w824 & ~w863;
assign w865 = pi0140 & ~w864;
assign w866 = ~pi0140 & w864;
assign w867 = ~w865 & ~w866;
assign w868 = (~pi0036 & ~w822) | (~pi0036 & w11453) | (~w822 & w11453);
assign w869 = ~w825 & ~w868;
assign w870 = pi0245 & ~w869;
assign w871 = ~pi0245 & w869;
assign w872 = ~w870 & ~w871;
assign w873 = (~pi0037 & ~w822) | (~pi0037 & w11454) | (~w822 & w11454);
assign w874 = ~w826 & ~w873;
assign w875 = pi0139 & ~w874;
assign w876 = ~pi0139 & w874;
assign w877 = ~w875 & ~w876;
assign w878 = ~pi0045 & ~w826;
assign w879 = ~w827 & ~w878;
assign w880 = ~pi0120 & w879;
assign w881 = pi0120 & ~w879;
assign w882 = ~w880 & ~w881;
assign w883 = (~pi0042 & ~w826) | (~pi0042 & w11455) | (~w826 & w11455);
assign w884 = ~w828 & ~w883;
assign w885 = pi0102 & ~w884;
assign w886 = ~pi0102 & w884;
assign w887 = ~w885 & ~w886;
assign w888 = pi0122 & ~w831;
assign w889 = ~pi0122 & w831;
assign w890 = ~w888 & ~w889;
assign w891 = pi0043 & ~pi0113;
assign w892 = ~pi0043 & pi0113;
assign w893 = ~w891 & ~w892;
assign w894 = (w893 & ~w826) | (w893 & w11456) | (~w826 & w11456);
assign w895 = w826 & w11457;
assign w896 = ~w894 & ~w895;
assign w897 = pi0031 & pi0043;
assign w898 = w826 & w11459;
assign w899 = pi0033 & ~pi0091;
assign w900 = ~pi0033 & pi0091;
assign w901 = ~w899 & ~w900;
assign w902 = w826 & w11460;
assign w903 = (w901 & ~w826) | (w901 & w11461) | (~w826 & w11461);
assign w904 = ~w902 & ~w903;
assign w905 = (~pi0032 & ~w826) | (~pi0032 & w11462) | (~w826 & w11462);
assign w906 = ~w898 & ~w905;
assign w907 = ~pi0090 & ~w906;
assign w908 = pi0090 & w906;
assign w909 = ~w907 & ~w908;
assign w910 = w398 & ~w837;
assign w911 = ~w842 & w910;
assign w912 = w911 & w11463;
assign w913 = w912 & w11464;
assign w914 = w913 & w11465;
assign w915 = w914 & w11466;
assign w916 = ~w890 & ~w904;
assign w917 = w915 & w11468;
assign w918 = w815 & w831;
assign w919 = (w918 & ~w917) | (w918 & w11469) | (~w917 & w11469);
assign w920 = ~w816 & ~w919;
assign w921 = ~pi1003 & ~w815;
assign w922 = w815 & w906;
assign w923 = (w922 & ~w917) | (w922 & w11470) | (~w917 & w11470);
assign w924 = ~w921 & ~w923;
assign w925 = ~pi1004 & ~w815;
assign w926 = w826 & w11471;
assign w927 = (~pi0033 & ~w826) | (~pi0033 & w11472) | (~w826 & w11472);
assign w928 = w815 & ~w926;
assign w929 = ~w927 & w928;
assign w930 = (w929 & ~w917) | (w929 & w11473) | (~w917 & w11473);
assign w931 = ~w925 & ~w930;
assign w932 = ~pi1009 & ~w815;
assign w933 = w815 & w859;
assign w934 = (w933 & ~w917) | (w933 & w11474) | (~w917 & w11474);
assign w935 = ~w932 & ~w934;
assign w936 = ~pi1010 & ~w815;
assign w937 = w815 & w864;
assign w938 = (w937 & ~w917) | (w937 & w11475) | (~w917 & w11475);
assign w939 = ~w936 & ~w938;
assign w940 = ~pi1011 & ~w815;
assign w941 = w815 & w869;
assign w942 = (w941 & ~w917) | (w941 & w11476) | (~w917 & w11476);
assign w943 = ~w940 & ~w942;
assign w944 = pi1012 & ~w815;
assign w945 = w815 & w874;
assign w946 = (w945 & ~w917) | (w945 & w11477) | (~w917 & w11477);
assign w947 = ~w944 & ~w946;
assign w948 = pi0999 & ~w815;
assign w949 = w815 & w834;
assign w950 = (w949 & ~w917) | (w949 & w11478) | (~w917 & w11478);
assign w951 = ~w948 & ~w950;
assign w952 = pi1007 & ~w815;
assign w953 = w815 & w849;
assign w954 = (w953 & ~w917) | (w953 & w11479) | (~w917 & w11479);
assign w955 = ~w952 & ~w954;
assign w956 = pi1006 & ~w815;
assign w957 = w815 & w844;
assign w958 = (w957 & ~w917) | (w957 & w11480) | (~w917 & w11480);
assign w959 = ~w956 & ~w958;
assign w960 = ~pi1008 & ~w815;
assign w961 = w815 & w854;
assign w962 = (w961 & ~w917) | (w961 & w11481) | (~w917 & w11481);
assign w963 = ~w960 & ~w962;
assign w964 = ~pi1000 & ~w815;
assign w965 = w815 & w884;
assign w966 = (w965 & ~w917) | (w965 & w11482) | (~w917 & w11482);
assign w967 = ~w964 & ~w966;
assign w968 = ~pi1002 & ~w815;
assign w969 = (~pi0043 & ~w826) | (~pi0043 & w11483) | (~w826 & w11483);
assign w970 = (w815 & ~w826) | (w815 & w11484) | (~w826 & w11484);
assign w971 = ~w969 & w970;
assign w972 = (w971 & ~w917) | (w971 & w11485) | (~w917 & w11485);
assign w973 = ~w968 & ~w972;
assign w974 = pi1005 & ~w815;
assign w975 = w815 & w839;
assign w976 = (w975 & ~w917) | (w975 & w11486) | (~w917 & w11486);
assign w977 = ~w974 & ~w976;
assign w978 = ~pi1013 & ~w815;
assign w979 = w815 & w879;
assign w980 = (w979 & ~w917) | (w979 & w11487) | (~w917 & w11487);
assign w981 = ~w978 & ~w980;
assign w982 = ~w432 & ~w441;
assign w983 = ~w428 & w11488;
assign w984 = (w982 & w983) | (w982 & w11489) | (w983 & w11489);
assign w985 = ~w983 & w11490;
assign w986 = ~w984 & ~w985;
assign w987 = ~pi1099 & ~w986;
assign w988 = ~pi0830 & pi1099;
assign w989 = ~w987 & ~w988;
assign w990 = ~w200 & ~w209;
assign w991 = w990 & w11491;
assign w992 = ~pi1692 & w204;
assign w993 = pi0047 & pi1549;
assign w994 = ~pi1753 & w993;
assign w995 = pi0093 & pi1667;
assign w996 = ~w994 & w995;
assign w997 = ~w992 & w996;
assign w998 = w991 & w997;
assign w999 = pi1747 & ~w998;
assign w1000 = w519 & ~w542;
assign w1001 = ~w519 & w542;
assign w1002 = ~w1000 & ~w1001;
assign w1003 = ~w624 & ~w1002;
assign w1004 = (w215 & w11494) | (w215 & w11495) | (w11494 & w11495);
assign w1005 = ~w1003 & w1004;
assign w1006 = ~w370 & w11496;
assign w1007 = pi0095 & ~w1006;
assign w1008 = (w1006 & w11498) | (w1006 & w11499) | (w11498 & w11499);
assign w1009 = (w1006 & w11500) | (w1006 & w11501) | (w11500 & w11501);
assign w1010 = (~w438 & w428) | (~w438 & w11502) | (w428 & w11502);
assign w1011 = ~w983 & w1007;
assign w1012 = ~w1010 & w1011;
assign w1013 = ~w1008 & ~w1009;
assign w1014 = ~w1012 & w1013;
assign w1015 = ~w594 & ~w628;
assign w1016 = w594 & w628;
assign w1017 = ~w1015 & ~w1016;
assign w1018 = ~w624 & ~w1017;
assign w1019 = (w215 & w11505) | (w215 & w11506) | (w11505 & w11506);
assign w1020 = ~w1018 & w1019;
assign w1021 = ~w615 & ~w624;
assign w1022 = (w215 & w11509) | (w215 & w11510) | (w11509 & w11510);
assign w1023 = ~w1021 & w1022;
assign w1024 = w539 & ~w612;
assign w1025 = ~w539 & w612;
assign w1026 = ~w1024 & ~w1025;
assign w1027 = ~w624 & ~w1026;
assign w1028 = (w215 & w11513) | (w215 & w11514) | (w11513 & w11514);
assign w1029 = ~w1027 & w1028;
assign w1030 = w519 & ~w588;
assign w1031 = ~w519 & w588;
assign w1032 = ~w1030 & ~w1031;
assign w1033 = ~w624 & ~w1032;
assign w1034 = (w215 & w11517) | (w215 & w11518) | (w11517 & w11518);
assign w1035 = ~w1033 & w1034;
assign w1036 = ~pi0010 & ~w568;
assign w1037 = pi0010 & w568;
assign w1038 = ~w1036 & ~w1037;
assign w1039 = ~w624 & ~w1038;
assign w1040 = (w215 & w11521) | (w215 & w11522) | (w11521 & w11522);
assign w1041 = ~w1039 & w1040;
assign w1042 = ~w207 & w209;
assign w1043 = pi0094 & w217;
assign w1044 = ~w1042 & ~w1043;
assign w1045 = pi1747 & ~w1044;
assign w1046 = (w1006 & w11523) | (w1006 & w11524) | (w11523 & w11524);
assign w1047 = (w1006 & w11525) | (w1006 & w11526) | (w11525 & w11526);
assign w1048 = ~w421 & ~w423;
assign w1049 = w427 & ~w1048;
assign w1050 = (w1007 & ~w428) | (w1007 & w11527) | (~w428 & w11527);
assign w1051 = ~w1049 & w1050;
assign w1052 = ~w1046 & ~w1047;
assign w1053 = ~w1051 & w1052;
assign w1054 = (w1006 & w11528) | (w1006 & w11529) | (w11528 & w11529);
assign w1055 = ~w412 & ~w413;
assign w1056 = w419 & w1007;
assign w1057 = ~w1055 & w1056;
assign w1058 = ~w419 & w1007;
assign w1059 = w1055 & w1058;
assign w1060 = ~pi0095 & ~pi1099;
assign w1061 = ~w398 & w1060;
assign w1062 = pi0012 & pi0767;
assign w1063 = pi0805 & ~w1062;
assign w1064 = ~pi0805 & w1062;
assign w1065 = ~w1063 & ~w1064;
assign w1066 = w1061 & w1065;
assign w1067 = ~w1054 & ~w1066;
assign w1068 = ~w1057 & w1067;
assign w1069 = ~w1059 & w1068;
assign w1070 = w212 & w11530;
assign w1071 = pi1692 & w204;
assign w1072 = pi1747 & ~w1070;
assign w1073 = ~w1071 & w1072;
assign w1074 = ~w545 & ~w624;
assign w1075 = (w215 & w11533) | (w215 & w11534) | (w11533 & w11534);
assign w1076 = ~w1074 & w1075;
assign w1077 = ~pi0094 & pi1747;
assign w1078 = w217 & w1077;
assign w1079 = ~pi0086 & ~pi1099;
assign w1080 = (w1006 & w11535) | (w1006 & w11536) | (w11535 & w11536);
assign w1081 = pi0895 & w418;
assign w1082 = w1058 & ~w1081;
assign w1083 = ~pi0012 & ~pi0767;
assign w1084 = ~w1062 & ~w1083;
assign w1085 = w1061 & w1084;
assign w1086 = ~w1080 & ~w1085;
assign w1087 = ~w1082 & w1086;
assign w1088 = pi0065 & ~pi1692;
assign w1089 = pi0093 & ~w1088;
assign w1090 = pi1747 & ~w1089;
assign w1091 = ~w185 & w11537;
assign w1092 = ~w201 & ~w992;
assign w1093 = (~pi0066 & w185) | (~pi0066 & w11538) | (w185 & w11538);
assign w1094 = pi1747 & ~w1091;
assign w1095 = ~w1093 & w1094;
assign w1096 = w1092 & w1095;
assign w1097 = ~pi0067 & ~pi0089;
assign w1098 = pi0109 & w1097;
assign w1099 = w366 & w11539;
assign w1100 = ~pi1049 & ~pi1096;
assign w1101 = pi1049 & pi1096;
assign w1102 = ~w1100 & ~w1101;
assign w1103 = ~pi1017 & ~pi1317;
assign w1104 = pi1017 & pi1317;
assign w1105 = ~w1103 & ~w1104;
assign w1106 = pi1042 & ~pi1285;
assign w1107 = ~pi1042 & pi1285;
assign w1108 = ~w1106 & ~w1107;
assign w1109 = pi1039 & ~pi1041;
assign w1110 = ~pi1039 & pi1041;
assign w1111 = ~w1109 & ~w1110;
assign w1112 = w1108 & ~w1111;
assign w1113 = ~w1108 & w1111;
assign w1114 = ~w1112 & ~w1113;
assign w1115 = ~w1105 & w1114;
assign w1116 = w1105 & ~w1114;
assign w1117 = ~w1115 & ~w1116;
assign w1118 = pi1313 & ~pi1334;
assign w1119 = ~pi1313 & pi1334;
assign w1120 = ~w1118 & ~w1119;
assign w1121 = pi1017 & ~pi1043;
assign w1122 = ~pi1017 & pi1043;
assign w1123 = ~w1121 & ~w1122;
assign w1124 = w1120 & w1123;
assign w1125 = ~w1120 & ~w1123;
assign w1126 = ~w1124 & ~w1125;
assign w1127 = ~pi1049 & w1126;
assign w1128 = pi1049 & ~w1126;
assign w1129 = ~w1127 & ~w1128;
assign w1130 = ~pi1039 & ~pi1040;
assign w1131 = pi1039 & pi1040;
assign w1132 = ~w1130 & ~w1131;
assign w1133 = pi1042 & ~pi1318;
assign w1134 = ~pi1042 & pi1318;
assign w1135 = ~w1133 & ~w1134;
assign w1136 = pi1044 & ~w1135;
assign w1137 = ~pi1044 & w1135;
assign w1138 = ~w1136 & ~w1137;
assign w1139 = pi1043 & ~pi1337;
assign w1140 = ~pi1043 & pi1337;
assign w1141 = ~w1139 & ~w1140;
assign w1142 = w1138 & w1141;
assign w1143 = ~w1138 & ~w1141;
assign w1144 = ~w1142 & ~w1143;
assign w1145 = ~w1132 & w1144;
assign w1146 = w1129 & ~w1145;
assign w1147 = w1132 & ~w1144;
assign w1148 = ~w1129 & ~w1147;
assign w1149 = pi1044 & ~pi1335;
assign w1150 = ~pi1044 & pi1335;
assign w1151 = ~w1149 & ~w1150;
assign w1152 = w1105 & w1151;
assign w1153 = ~w1105 & ~w1151;
assign w1154 = ~w1152 & ~w1153;
assign w1155 = pi1313 & ~pi1336;
assign w1156 = ~pi1313 & pi1336;
assign w1157 = ~w1155 & ~w1156;
assign w1158 = w1138 & w1157;
assign w1159 = ~w1138 & ~w1157;
assign w1160 = ~w1158 & ~w1159;
assign w1161 = w1154 & w1160;
assign w1162 = pi1049 & ~w1132;
assign w1163 = (~w1162 & ~w1126) | (~w1162 & w11540) | (~w1126 & w11540);
assign w1164 = ~pi1041 & w1163;
assign w1165 = pi1041 & ~w1163;
assign w1166 = ~w1164 & ~w1165;
assign w1167 = ~w1160 & ~w1166;
assign w1168 = ~w1154 & w1166;
assign w1169 = ~w1117 & ~w1161;
assign w1170 = ~w1146 & w1169;
assign w1171 = ~w1148 & w1170;
assign w1172 = ~w1167 & ~w1168;
assign w1173 = w1171 & w1172;
assign w1174 = w1171 & w11541;
assign w1175 = pi1039 & ~pi1094;
assign w1176 = pi1041 & ~pi1069;
assign w1177 = ~pi1041 & pi1069;
assign w1178 = pi1017 & ~pi1098;
assign w1179 = ~pi1039 & pi1094;
assign w1180 = pi1040 & ~pi1095;
assign w1181 = ~pi1040 & pi1095;
assign w1182 = pi1042 & ~pi1097;
assign w1183 = pi1043 & ~pi1068;
assign w1184 = ~pi1043 & pi1068;
assign w1185 = ~pi1017 & pi1098;
assign w1186 = ~pi1042 & pi1097;
assign w1187 = pi1229 & ~pi1479;
assign w1188 = ~pi1228 & ~pi1236;
assign w1189 = ~w1187 & w1188;
assign w1190 = ~pi1227 & ~w1189;
assign w1191 = pi1234 & ~w1175;
assign w1192 = ~w1176 & ~w1177;
assign w1193 = ~w1178 & ~w1179;
assign w1194 = ~w1180 & ~w1181;
assign w1195 = ~w1182 & ~w1183;
assign w1196 = ~w1184 & ~w1185;
assign w1197 = ~w1186 & w1196;
assign w1198 = w1194 & w1195;
assign w1199 = w1192 & w1193;
assign w1200 = ~w1102 & w1191;
assign w1201 = w1199 & w1200;
assign w1202 = w1197 & w1198;
assign w1203 = ~w1190 & w1202;
assign w1204 = w1201 & w1203;
assign w1205 = w1174 & w1204;
assign w1206 = (pi1747 & ~w1174) | (pi1747 & w11542) | (~w1174 & w11542);
assign w1207 = w366 & w11543;
assign w1208 = ~pi1227 & ~pi1228;
assign w1209 = w356 & w1208;
assign w1210 = (~w369 & ~w1209) | (~w369 & w11544) | (~w1209 & w11544);
assign w1211 = (~w374 & ~w372) | (~w374 & w11545) | (~w372 & w11545);
assign w1212 = pi1229 & pi1236;
assign w1213 = w355 & w1212;
assign w1214 = ~pi0771 & ~w1213;
assign w1215 = (~pi0801 & ~w1214) | (~pi0801 & w11546) | (~w1214 & w11546);
assign w1216 = w1211 & ~w1215;
assign w1217 = ~w385 & w11547;
assign w1218 = (w1207 & w1217) | (w1207 & w11548) | (w1217 & w11548);
assign w1219 = ~pi0067 & pi0089;
assign w1220 = w366 & w11549;
assign w1221 = ~pi1416 & w1220;
assign w1222 = ~pi0092 & pi0108;
assign w1223 = ~pi0109 & w1097;
assign w1224 = w365 & w1223;
assign w1225 = pi1417 & w1222;
assign w1226 = w365 & w11550;
assign w1227 = ~w1221 & ~w1226;
assign w1228 = ~pi1626 & ~pi1627;
assign w1229 = ~pi0695 & ~pi0696;
assign w1230 = ~pi0382 & pi0647;
assign w1231 = w1229 & w1230;
assign w1232 = ~w1228 & w1231;
assign w1233 = ~pi0722 & ~pi0723;
assign w1234 = pi0727 & pi0729;
assign w1235 = ~pi0730 & ~pi0731;
assign w1236 = ~pi0732 & pi0733;
assign w1237 = ~pi0734 & ~pi0735;
assign w1238 = ~pi0736 & ~pi0737;
assign w1239 = ~pi0738 & ~pi0744;
assign w1240 = ~pi0745 & pi0746;
assign w1241 = w1239 & w1240;
assign w1242 = w1237 & w1238;
assign w1243 = w1235 & w1236;
assign w1244 = w1233 & w1234;
assign w1245 = w1243 & w1244;
assign w1246 = w1241 & w1242;
assign w1247 = w1245 & w1246;
assign w1248 = w1232 & ~w1247;
assign w1249 = (~pi0138 & w1247) | (~pi0138 & w11551) | (w1247 & w11551);
assign w1250 = w1220 & ~w1249;
assign w1251 = w361 & w1223;
assign w1252 = (~pi0111 & ~w389) | (~pi0111 & w11552) | (~w389 & w11552);
assign w1253 = pi0110 & ~w362;
assign w1254 = pi0088 & pi0112;
assign w1255 = ~pi0095 & ~w1254;
assign w1256 = ~w363 & w1255;
assign w1257 = ~w1253 & w1256;
assign w1258 = w1257 & w11553;
assign w1259 = ~w1099 & ~w1258;
assign w1260 = ~w1250 & w1259;
assign w1261 = w1227 & w1260;
assign w1262 = ~w1218 & w1261;
assign w1263 = w1206 & w1262;
assign w1264 = ~w385 & w11554;
assign w1265 = ~w1211 & w1264;
assign w1266 = (~pi0121 & ~w1264) | (~pi0121 & w11555) | (~w1264 & w11555);
assign w1267 = (w1264 & w11556) | (w1264 & w11557) | (w11556 & w11557);
assign w1268 = (pi0762 & w395) | (pi0762 & w11558) | (w395 & w11558);
assign w1269 = ~w395 & w11559;
assign w1270 = ~w1268 & ~w1269;
assign w1271 = (pi0768 & w395) | (pi0768 & w11560) | (w395 & w11560);
assign w1272 = ~w395 & w11561;
assign w1273 = ~w1271 & ~w1272;
assign w1274 = (pi0827 & w395) | (pi0827 & w11562) | (w395 & w11562);
assign w1275 = ~w395 & w11563;
assign w1276 = ~w1274 & ~w1275;
assign w1277 = w1270 & w1273;
assign w1278 = w1276 & w1277;
assign w1279 = (pi0826 & w395) | (pi0826 & w11564) | (w395 & w11564);
assign w1280 = ~w395 & w11565;
assign w1281 = ~w1279 & ~w1280;
assign w1282 = w1277 & w11566;
assign w1283 = pi0877 & ~w1282;
assign w1284 = w1267 & ~w1283;
assign w1285 = (~w1264 & w11567) | (~w1264 & w11568) | (w11567 & w11568);
assign w1286 = ~pi0071 & ~pi0076;
assign w1287 = ~pi0077 & ~pi0078;
assign w1288 = ~pi0079 & w1287;
assign w1289 = w1286 & w1288;
assign w1290 = pi1091 & pi1101;
assign w1291 = ~pi0069 & ~pi0070;
assign w1292 = ~pi0074 & ~pi0080;
assign w1293 = ~pi0081 & ~pi0082;
assign w1294 = ~pi0083 & w1293;
assign w1295 = w1291 & w1292;
assign w1296 = w1294 & w1295;
assign w1297 = w1289 & w1296;
assign w1298 = ~pi0075 & w1297;
assign w1299 = (w1297 & w11570) | (w1297 & w11571) | (w11570 & w11571);
assign w1300 = ~w1299 & w11572;
assign w1301 = ~w1299 & w11573;
assign w1302 = ~pi0081 & w1301;
assign w1303 = w1301 & w1293;
assign w1304 = w1301 & w1294;
assign w1305 = (pi0069 & ~w1301) | (pi0069 & w11574) | (~w1301 & w11574);
assign w1306 = w1301 & w11575;
assign w1307 = w1285 & w11576;
assign w1308 = ~w1284 & ~w1307;
assign w1309 = w1301 & w11577;
assign w1310 = (pi0070 & ~w1301) | (pi0070 & w11578) | (~w1301 & w11578);
assign w1311 = ~w1299 & w11579;
assign w1312 = ~w1310 & ~w1311;
assign w1313 = w1266 & ~w1312;
assign w1314 = pi1747 & ~w1313;
assign w1315 = (pi0751 & ~w370) | (pi0751 & w11580) | (~w370 & w11580);
assign w1316 = ~w395 & w1315;
assign w1317 = ~w370 & w394;
assign w1318 = (pi0770 & ~w370) | (pi0770 & w11581) | (~w370 & w11581);
assign w1319 = ~w1317 & w1318;
assign w1320 = ~w1316 & ~w1319;
assign w1321 = ~pi0877 & ~w1281;
assign w1322 = w1278 & ~w1321;
assign w1323 = pi0877 & w1281;
assign w1324 = (pi0825 & w395) | (pi0825 & w11582) | (w395 & w11582);
assign w1325 = ~w395 & w11583;
assign w1326 = ~w1324 & ~w1325;
assign w1327 = ~pi0759 & ~w1326;
assign w1328 = ~w1323 & w1327;
assign w1329 = w1322 & ~w1328;
assign w1330 = (pi0772 & w395) | (pi0772 & w11584) | (w395 & w11584);
assign w1331 = ~w395 & w11585;
assign w1332 = ~w1330 & ~w1331;
assign w1333 = pi0810 & w1332;
assign w1334 = pi0759 & w1326;
assign w1335 = (pi0871 & ~w370) | (pi0871 & w11586) | (~w370 & w11586);
assign w1336 = ~w1317 & w1335;
assign w1337 = (pi0754 & ~w370) | (pi0754 & w11587) | (~w370 & w11587);
assign w1338 = ~w395 & w1337;
assign w1339 = ~w1336 & ~w1338;
assign w1340 = pi0750 & w1339;
assign w1341 = (pi0818 & ~w370) | (pi0818 & w11588) | (~w370 & w11588);
assign w1342 = ~w1317 & w1341;
assign w1343 = (pi0841 & ~w370) | (pi0841 & w11589) | (~w370 & w11589);
assign w1344 = ~w395 & w1343;
assign w1345 = ~w1342 & ~w1344;
assign w1346 = pi0859 & w1345;
assign w1347 = ~w1340 & ~w1346;
assign w1348 = ~pi0750 & ~w1339;
assign w1349 = (pi0842 & ~w370) | (pi0842 & w11590) | (~w370 & w11590);
assign w1350 = ~w395 & w1349;
assign w1351 = (pi0819 & ~w370) | (pi0819 & w11591) | (~w370 & w11591);
assign w1352 = ~w1317 & w1351;
assign w1353 = ~w1350 & ~w1352;
assign w1354 = ~pi0804 & ~w1353;
assign w1355 = ~w1348 & ~w1354;
assign w1356 = ~w1347 & w1355;
assign w1357 = (pi0821 & w395) | (pi0821 & w11592) | (w395 & w11592);
assign w1358 = ~w395 & w11593;
assign w1359 = ~w1357 & ~w1358;
assign w1360 = pi0806 & w1359;
assign w1361 = pi0804 & w1353;
assign w1362 = ~w1360 & ~w1361;
assign w1363 = ~pi0807 & ~w1320;
assign w1364 = ~pi0806 & ~w1359;
assign w1365 = ~w1363 & ~w1364;
assign w1366 = (w1365 & w1356) | (w1365 & w11594) | (w1356 & w11594);
assign w1367 = pi0807 & w1320;
assign w1368 = (pi0822 & w395) | (pi0822 & w11595) | (w395 & w11595);
assign w1369 = ~w395 & w11596;
assign w1370 = ~w1368 & ~w1369;
assign w1371 = pi0755 & w1370;
assign w1372 = ~w1367 & ~w1371;
assign w1373 = ~pi0755 & ~w1370;
assign w1374 = (pi0823 & w395) | (pi0823 & w11597) | (w395 & w11597);
assign w1375 = ~w395 & w11598;
assign w1376 = ~w1374 & ~w1375;
assign w1377 = ~pi0808 & ~w1376;
assign w1378 = ~w1373 & ~w1377;
assign w1379 = pi0808 & w1376;
assign w1380 = (pi0824 & w395) | (pi0824 & w11600) | (w395 & w11600);
assign w1381 = ~w395 & w11601;
assign w1382 = ~w1380 & ~w1381;
assign w1383 = pi0809 & w1382;
assign w1384 = ~w1379 & ~w1383;
assign w1385 = (~w1366 & w11602) | (~w1366 & w11603) | (w11602 & w11603);
assign w1386 = ~pi0809 & ~w1382;
assign w1387 = ~pi0810 & ~w1332;
assign w1388 = ~w1386 & ~w1387;
assign w1389 = ~w1323 & ~w1333;
assign w1390 = ~w1334 & w1389;
assign w1391 = (w1390 & w1385) | (w1390 & w11604) | (w1385 & w11604);
assign w1392 = ~w1391 & w11605;
assign w1393 = (pi0807 & w1391) | (pi0807 & w11606) | (w1391 & w11606);
assign w1394 = ~w1392 & ~w1393;
assign w1395 = w1267 & w1394;
assign w1396 = ~w1299 & w11607;
assign w1397 = ~w1299 & w11608;
assign w1398 = ~w1299 & w11609;
assign w1399 = (pi0071 & w1299) | (pi0071 & w11610) | (w1299 & w11610);
assign w1400 = ~w1299 & w11611;
assign w1401 = (~w1264 & w11612) | (~w1264 & w11613) | (w11612 & w11613);
assign w1402 = ~w1400 & w1401;
assign w1403 = ~w1395 & ~w1402;
assign w1404 = ~pi0711 & ~pi1608;
assign w1405 = ~pi1080 & pi1132;
assign w1406 = pi0137 & pi1492;
assign w1407 = ~w1405 & w1406;
assign w1408 = (pi1839 & ~w1405) | (pi1839 & w11614) | (~w1405 & w11614);
assign w1409 = ~w1407 & w1408;
assign w1410 = (~w1404 & w1409) | (~w1404 & w11615) | (w1409 & w11615);
assign w1411 = pi1747 & ~w1410;
assign w1412 = ~w1391 & w11616;
assign w1413 = (pi0859 & w1391) | (pi0859 & w11617) | (w1391 & w11617);
assign w1414 = ~w1412 & ~w1413;
assign w1415 = w1267 & w1414;
assign w1416 = (pi0073 & ~w206) | (pi0073 & w11618) | (~w206 & w11618);
assign w1417 = ~w1290 & w1416;
assign w1418 = (~w1417 & w1299) | (~w1417 & w11619) | (w1299 & w11619);
assign w1419 = (~w1264 & w11620) | (~w1264 & w11621) | (w11620 & w11621);
assign w1420 = ~w1415 & ~w1419;
assign w1421 = (pi0074 & ~w1301) | (pi0074 & w11622) | (~w1301 & w11622);
assign w1422 = ~w1309 & ~w1421;
assign w1423 = w1266 & ~w1422;
assign w1424 = pi1747 & ~w1423;
assign w1425 = pi0075 & w1311;
assign w1426 = ~pi0075 & ~w1311;
assign w1427 = ~w1425 & ~w1426;
assign w1428 = w1266 & w1427;
assign w1429 = pi1747 & ~w1428;
assign w1430 = ~w1391 & w11623;
assign w1431 = (pi0750 & w1391) | (pi0750 & w11624) | (w1391 & w11624);
assign w1432 = ~w1430 & ~w1431;
assign w1433 = w1267 & w1432;
assign w1434 = (pi0076 & w1299) | (pi0076 & w11625) | (w1299 & w11625);
assign w1435 = ~w1396 & ~w1434;
assign w1436 = w1285 & w1435;
assign w1437 = ~w1433 & ~w1436;
assign w1438 = ~w1391 & w11626;
assign w1439 = (pi0804 & w1391) | (pi0804 & w11627) | (w1391 & w11627);
assign w1440 = ~w1438 & ~w1439;
assign w1441 = w1267 & w1440;
assign w1442 = (pi0077 & w1299) | (pi0077 & w11628) | (w1299 & w11628);
assign w1443 = ~w1397 & ~w1442;
assign w1444 = w1285 & w1443;
assign w1445 = ~w1441 & ~w1444;
assign w1446 = ~w1391 & w11629;
assign w1447 = (pi0806 & w1391) | (pi0806 & w11630) | (w1391 & w11630);
assign w1448 = ~w1446 & ~w1447;
assign w1449 = w1267 & w1448;
assign w1450 = (pi0078 & w1299) | (pi0078 & w11631) | (w1299 & w11631);
assign w1451 = ~w1398 & ~w1450;
assign w1452 = w1285 & w1451;
assign w1453 = ~w1449 & ~w1452;
assign w1454 = ~w1391 & w11632;
assign w1455 = (pi0755 & w1391) | (pi0755 & w11633) | (w1391 & w11633);
assign w1456 = ~w1454 & ~w1455;
assign w1457 = w1267 & w1456;
assign w1458 = (pi0079 & w1299) | (pi0079 & w11634) | (w1299 & w11634);
assign w1459 = (~w1264 & w11635) | (~w1264 & w11636) | (w11635 & w11636);
assign w1460 = ~w1458 & w1459;
assign w1461 = ~w1457 & ~w1460;
assign w1462 = ~w1391 & w11637;
assign w1463 = (pi0808 & w1391) | (pi0808 & w11638) | (w1391 & w11638);
assign w1464 = ~w1462 & ~w1463;
assign w1465 = w1267 & w1464;
assign w1466 = (pi0080 & w1299) | (pi0080 & w11639) | (w1299 & w11639);
assign w1467 = ~w1301 & ~w1466;
assign w1468 = w1285 & w1467;
assign w1469 = ~w1465 & ~w1468;
assign w1470 = ~w1391 & w11640;
assign w1471 = (pi0809 & w1391) | (pi0809 & w11641) | (w1391 & w11641);
assign w1472 = ~w1470 & ~w1471;
assign w1473 = w1267 & w1472;
assign w1474 = pi0081 & ~w1301;
assign w1475 = ~w1302 & ~w1474;
assign w1476 = w1285 & w1475;
assign w1477 = ~w1473 & ~w1476;
assign w1478 = ~w1391 & w11642;
assign w1479 = (pi0810 & w1391) | (pi0810 & w11643) | (w1391 & w11643);
assign w1480 = ~w1478 & ~w1479;
assign w1481 = w1267 & w1480;
assign w1482 = (pi0082 & ~w1301) | (pi0082 & w11644) | (~w1301 & w11644);
assign w1483 = w1285 & w11645;
assign w1484 = ~w1481 & ~w1483;
assign w1485 = (pi0759 & ~w1278) | (pi0759 & w11646) | (~w1278 & w11646);
assign w1486 = w1322 & w11647;
assign w1487 = ~w1485 & ~w1486;
assign w1488 = ~w1486 & w11648;
assign w1489 = (pi0083 & ~w1301) | (pi0083 & w11649) | (~w1301 & w11649);
assign w1490 = w1285 & w11650;
assign w1491 = ~w1488 & ~w1490;
assign w1492 = ~pi0713 & ~pi1583;
assign w1493 = ~pi1144 & pi1259;
assign w1494 = pi0142 & pi1491;
assign w1495 = ~w1493 & w1494;
assign w1496 = (pi1840 & ~w1493) | (pi1840 & w11651) | (~w1493 & w11651);
assign w1497 = ~w1495 & w1496;
assign w1498 = (~w1492 & w1497) | (~w1492 & w11652) | (w1497 & w11652);
assign w1499 = pi1747 & ~w1498;
assign w1500 = ~pi0676 & ~pi1607;
assign w1501 = ~pi1256 & pi1257;
assign w1502 = pi0143 & pi1477;
assign w1503 = ~w1501 & w1502;
assign w1504 = (pi1838 & ~w1501) | (pi1838 & w11653) | (~w1501 & w11653);
assign w1505 = ~w1503 & w1504;
assign w1506 = (~w1500 & w1505) | (~w1500 & w11654) | (w1505 & w11654);
assign w1507 = pi1747 & ~w1506;
assign w1508 = pi0117 & ~w1320;
assign w1509 = ~pi0117 & w1320;
assign w1510 = ~w1508 & ~w1509;
assign w1511 = pi0105 & ~w1353;
assign w1512 = ~pi0103 & w1345;
assign w1513 = (pi0104 & ~w1345) | (pi0104 & w11655) | (~w1345 & w11655);
assign w1514 = w1345 & w11656;
assign w1515 = ~w1339 & ~w1514;
assign w1516 = ~w1513 & ~w1515;
assign w1517 = ~w1515 & w11657;
assign w1518 = ~pi0105 & w1353;
assign w1519 = (pi0106 & ~w1353) | (pi0106 & w11658) | (~w1353 & w11658);
assign w1520 = ~w1517 & w1519;
assign w1521 = ~w1517 & w11659;
assign w1522 = ~w1511 & ~w1518;
assign w1523 = ~w1516 & w1522;
assign w1524 = (~pi0106 & w1353) | (~pi0106 & w11660) | (w1353 & w11660);
assign w1525 = (w1524 & w1516) | (w1524 & w11661) | (w1516 & w11661);
assign w1526 = ~w1359 & w1510;
assign w1527 = ~w1525 & w1526;
assign w1528 = ~w1521 & ~w1527;
assign w1529 = ~w1527 & w11662;
assign w1530 = ~pi0098 & w1376;
assign w1531 = pi0099 & ~w1382;
assign w1532 = ~pi0099 & w1382;
assign w1533 = ~w1531 & ~w1532;
assign w1534 = ~w1530 & w1533;
assign w1535 = pi0107 & ~w1370;
assign w1536 = ~pi0107 & w1370;
assign w1537 = ~w1535 & ~w1536;
assign w1538 = w1534 & w1537;
assign w1539 = pi0101 & ~w1326;
assign w1540 = ~pi0100 & w1332;
assign w1541 = w1539 & w1540;
assign w1542 = w1534 & w11663;
assign w1543 = pi0100 & ~w1332;
assign w1544 = pi0098 & ~w1376;
assign w1545 = ~w1535 & ~w1544;
assign w1546 = w1534 & ~w1545;
assign w1547 = ~w1531 & ~w1543;
assign w1548 = (w1547 & ~w1534) | (w1547 & w11664) | (~w1534 & w11664);
assign w1549 = (w1539 & w1548) | (w1539 & w1541) | (w1548 & w1541);
assign w1550 = (w1549 & w1529) | (w1549 & w11665) | (w1529 & w11665);
assign w1551 = ~pi0101 & ~w1326;
assign w1552 = ~w1548 & w1553;
assign w1553 = ~w1540 & w1551;
assign w1554 = w1534 & w11666;
assign w1555 = (~w1552 & w1529) | (~w1552 & w11667) | (w1529 & w11667);
assign w1556 = ~w1550 & w1555;
assign w1557 = pi0119 & ~w1281;
assign w1558 = (pi0101 & ~w1332) | (pi0101 & w11668) | (~w1332 & w11668);
assign w1559 = w1534 & w11669;
assign w1560 = ~w1548 & w1558;
assign w1561 = (~w1560 & w1529) | (~w1560 & w11670) | (w1529 & w11670);
assign w1562 = ~w1557 & w1561;
assign w1563 = w1556 & w1562;
assign w1564 = ~pi0119 & w1281;
assign w1565 = pi0126 & ~w1276;
assign w1566 = ~pi0126 & w1276;
assign w1567 = ~w1565 & ~w1566;
assign w1568 = ~w1564 & w1567;
assign w1569 = pi0127 & ~w1270;
assign w1570 = ~pi0127 & w1270;
assign w1571 = ~w1569 & ~w1570;
assign w1572 = w1568 & w1571;
assign w1573 = ~w1563 & w1572;
assign w1574 = w1565 & w1571;
assign w1575 = (~w1569 & ~w1571) | (~w1569 & w11671) | (~w1571 & w11671);
assign w1576 = pi0123 & ~w1575;
assign w1577 = ~pi0123 & w1575;
assign w1578 = ~w1576 & ~w1577;
assign w1579 = w1273 & ~w1578;
assign w1580 = ~w1273 & w1578;
assign w1581 = ~w1579 & ~w1580;
assign w1582 = ~w1563 & w11672;
assign w1583 = (~w1581 & w1563) | (~w1581 & w11673) | (w1563 & w11673);
assign w1584 = ~w1582 & ~w1583;
assign w1585 = ~pi0721 & ~pi1604;
assign w1586 = ~pi1112 & pi1113;
assign w1587 = pi0184 & pi1520;
assign w1588 = ~w1586 & w1587;
assign w1589 = (pi1841 & ~w1586) | (pi1841 & w11674) | (~w1586 & w11674);
assign w1590 = ~w1588 & w1589;
assign w1591 = (~w1585 & w1590) | (~w1585 & w11675) | (w1590 & w11675);
assign w1592 = pi1747 & ~w1591;
assign w1593 = (~w1174 & w11676) | (~w1174 & w11677) | (w11676 & w11677);
assign w1594 = (w368 & w385) | (w368 & w11678) | (w385 & w11678);
assign w1595 = w1593 & w1594;
assign w1596 = w1215 & w1264;
assign w1597 = (~w1174 & w11679) | (~w1174 & w11680) | (w11679 & w11680);
assign w1598 = ~pi0138 & pi1416;
assign w1599 = w366 & w11681;
assign w1600 = (~w1174 & w11684) | (~w1174 & w11685) | (w11684 & w11685);
assign w1601 = ~w1597 & ~w1600;
assign w1602 = pi0999 & ~w1353;
assign w1603 = (~pi1005 & w1353) | (~pi1005 & w11686) | (w1353 & w11686);
assign w1604 = ~w1359 & ~w1603;
assign w1605 = ~pi0999 & w1353;
assign w1606 = ~w1602 & ~w1605;
assign w1607 = ~pi0998 & w1339;
assign w1608 = pi0998 & ~w1339;
assign w1609 = pi0997 & ~w1345;
assign w1610 = ~w1608 & ~w1609;
assign w1611 = ~w1607 & ~w1610;
assign w1612 = ~w1359 & w1606;
assign w1613 = w1611 & w1612;
assign w1614 = ~w1604 & ~w1613;
assign w1615 = ~pi1006 & w1320;
assign w1616 = pi1006 & ~w1320;
assign w1617 = ~w1615 & ~w1616;
assign w1618 = (pi1005 & ~w1353) | (pi1005 & w11687) | (~w1353 & w11687);
assign w1619 = w1617 & ~w1618;
assign w1620 = ~w1602 & w1617;
assign w1621 = ~w1611 & w1620;
assign w1622 = ~w1619 & ~w1621;
assign w1623 = w1614 & ~w1622;
assign w1624 = pi1008 & w1376;
assign w1625 = pi1009 & w1382;
assign w1626 = ~w1624 & ~w1625;
assign w1627 = pi1007 & ~w1370;
assign w1628 = ~pi1007 & w1370;
assign w1629 = ~w1627 & ~w1628;
assign w1630 = ~w1615 & w1629;
assign w1631 = w1626 & w1630;
assign w1632 = ~pi1011 & ~w1326;
assign w1633 = ~w1326 & w11688;
assign w1634 = ~pi1010 & ~w1332;
assign w1635 = ~pi1008 & ~w1376;
assign w1636 = ~w1627 & ~w1635;
assign w1637 = w1626 & ~w1636;
assign w1638 = ~pi1009 & ~w1382;
assign w1639 = ~w1637 & ~w1638;
assign w1640 = ~w1637 & w11689;
assign w1641 = ~w1637 & w11690;
assign w1642 = pi1011 & w1326;
assign w1643 = ~w1632 & ~w1642;
assign w1644 = pi1010 & w1332;
assign w1645 = w1643 & ~w1644;
assign w1646 = (~w1632 & ~w1643) | (~w1632 & w11692) | (~w1643 & w11692);
assign w1647 = pi1012 & ~w1646;
assign w1648 = (~w1623 & w11693) | (~w1623 & w11694) | (w11693 & w11694);
assign w1649 = ~pi1012 & ~w1632;
assign w1650 = (~w1281 & w1632) | (~w1281 & w11695) | (w1632 & w11695);
assign w1651 = w1643 & w11696;
assign w1652 = ~w1640 & w1651;
assign w1653 = w1631 & w1651;
assign w1654 = (~w1652 & w1623) | (~w1652 & w11697) | (w1623 & w11697);
assign w1655 = ~w1650 & w1654;
assign w1656 = (~pi1013 & ~w1655) | (~pi1013 & w11698) | (~w1655 & w11698);
assign w1657 = ~pi1000 & ~w1270;
assign w1658 = ~w1270 & w11699;
assign w1659 = w1276 & ~w1658;
assign w1660 = ~w1656 & w1659;
assign w1661 = pi1013 & ~w1650;
assign w1662 = w1654 & w1661;
assign w1663 = ~w1648 & w1662;
assign w1664 = w1662 & w11700;
assign w1665 = pi1000 & w1270;
assign w1666 = (pi1001 & ~w1270) | (pi1001 & w11699) | (~w1270 & w11699);
assign w1667 = ~w1664 & w1666;
assign w1668 = ~w1660 & w1667;
assign w1669 = (~pi1001 & w1270) | (~pi1001 & w11701) | (w1270 & w11701);
assign w1670 = w1276 & w1669;
assign w1671 = ~w1656 & w1670;
assign w1672 = (~w1665 & ~w1662) | (~w1665 & w11702) | (~w1662 & w11702);
assign w1673 = w1669 & ~w1672;
assign w1674 = ~w1671 & ~w1673;
assign w1675 = ~w1668 & w1674;
assign w1676 = w1273 & ~w1675;
assign w1677 = ~w1273 & w1675;
assign w1678 = ~w1676 & ~w1677;
assign w1679 = ~w1273 & w1674;
assign w1680 = ~pi1002 & ~w1668;
assign w1681 = ~w1679 & w1680;
assign w1682 = pi1002 & w1668;
assign w1683 = pi1002 & ~w1273;
assign w1684 = w1674 & w1683;
assign w1685 = ~w1682 & ~w1684;
assign w1686 = ~w1681 & w1685;
assign w1687 = (~w1174 & w11703) | (~w1174 & w11704) | (w11703 & w11704);
assign w1688 = (~w1174 & w11705) | (~w1174 & w11706) | (w11705 & w11706);
assign w1689 = pi0092 & ~pi0108;
assign w1690 = pi1251 & w1689;
assign w1691 = (~w1174 & w11707) | (~w1174 & w11708) | (w11707 & w11708);
assign w1692 = ~w1687 & ~w1691;
assign w1693 = ~w389 & ~w1594;
assign w1694 = ~pi0750 & ~pi0755;
assign w1695 = ~pi0759 & ~pi0804;
assign w1696 = ~pi0806 & ~pi0807;
assign w1697 = ~pi0808 & ~pi0809;
assign w1698 = ~pi0810 & ~pi0859;
assign w1699 = ~pi0877 & w1698;
assign w1700 = w1696 & w1697;
assign w1701 = w1694 & w1695;
assign w1702 = w1700 & w1701;
assign w1703 = w1699 & w1702;
assign w1704 = w1265 & w1703;
assign w1705 = pi0799 & ~pi0800;
assign w1706 = ~pi1251 & w1689;
assign w1707 = w1705 & w1706;
assign w1708 = ~pi1227 & pi1228;
assign w1709 = ~pi1229 & ~pi1236;
assign w1710 = w1708 & w1709;
assign w1711 = pi1233 & w1710;
assign w1712 = ~pi1417 & w1222;
assign w1713 = w1711 & w1712;
assign w1714 = ~w1707 & ~w1713;
assign w1715 = w1223 & w11709;
assign w1716 = ~w1252 & w1715;
assign w1717 = (~w1716 & w1714) | (~w1716 & w11710) | (w1714 & w11710);
assign w1718 = pi0110 & pi0111;
assign w1719 = ~pi0095 & ~w1718;
assign w1720 = ~w1717 & w1719;
assign w1721 = w1206 & w1720;
assign w1722 = w406 & ~w1464;
assign w1723 = w451 & ~w1722;
assign w1724 = w406 & ~w1472;
assign w1725 = w470 & ~w1724;
assign w1726 = w406 & ~w1480;
assign w1727 = w466 & ~w1726;
assign w1728 = (w406 & w1486) | (w406 & w11711) | (w1486 & w11711);
assign w1729 = w477 & ~w1728;
assign w1730 = (w1639 & w1623) | (w1639 & w11712) | (w1623 & w11712);
assign w1731 = (w1645 & ~w1730) | (w1645 & w11713) | (~w1730 & w11713);
assign w1732 = (~w1648 & w1731) | (~w1648 & w11714) | (w1731 & w11714);
assign w1733 = ~w1281 & w1732;
assign w1734 = w1281 & ~w1732;
assign w1735 = ~w1733 & ~w1734;
assign w1736 = w406 & ~w1414;
assign w1737 = (~w415 & ~w407) | (~w415 & w11715) | (~w407 & w11715);
assign w1738 = ~w1736 & w1737;
assign w1739 = w406 & ~w1432;
assign w1740 = (~w409 & ~w407) | (~w409 & w11716) | (~w407 & w11716);
assign w1741 = ~w1739 & w1740;
assign w1742 = w406 & ~w1440;
assign w1743 = w425 & ~w1742;
assign w1744 = w406 & ~w1448;
assign w1745 = w434 & ~w1744;
assign w1746 = w406 & ~w1456;
assign w1747 = w446 & ~w1746;
assign w1748 = ~w1705 & w1706;
assign w1749 = ~w1711 & w1712;
assign w1750 = ~w1748 & ~w1749;
assign w1751 = w1688 & ~w1750;
assign w1752 = w1232 & w1247;
assign w1753 = (~w1174 & w11717) | (~w1174 & w11718) | (w11717 & w11718);
assign w1754 = ~w1705 & w1753;
assign w1755 = ~pi0138 & pi1747;
assign w1756 = w366 & w11719;
assign w1757 = ~w1205 & w1756;
assign w1758 = w1705 & w1753;
assign w1759 = pi0095 & w364;
assign w1760 = w1251 & w1759;
assign w1761 = w1206 & w1760;
assign w1762 = ~w1657 & ~w1665;
assign w1763 = ~w1656 & ~w1663;
assign w1764 = ~w1276 & w1763;
assign w1765 = (~w1656 & ~w1763) | (~w1656 & w11720) | (~w1763 & w11720);
assign w1766 = ~w1762 & w1765;
assign w1767 = w1762 & ~w1765;
assign w1768 = ~w1766 & ~w1767;
assign w1769 = pi1439 & pi1747;
assign w1770 = pi0198 & pi1459;
assign w1771 = ~pi0114 & ~w1770;
assign w1772 = w1769 & ~w1771;
assign w1773 = pi1473 & pi1747;
assign w1774 = pi0198 & pi1480;
assign w1775 = ~pi0115 & ~w1774;
assign w1776 = w1773 & ~w1775;
assign w1777 = pi1440 & pi1747;
assign w1778 = pi0198 & pi1430;
assign w1779 = ~pi0116 & ~w1778;
assign w1780 = w1777 & ~w1779;
assign w1781 = w406 & ~w1394;
assign w1782 = w430 & ~w1781;
assign w1783 = pi1437 & pi1747;
assign w1784 = pi0198 & pi1447;
assign w1785 = ~pi0118 & ~w1784;
assign w1786 = w1783 & ~w1785;
assign w1787 = ~w1282 & w11721;
assign w1788 = w459 & ~w1787;
assign w1789 = ~w1634 & ~w1644;
assign w1790 = (~w1623 & w11722) | (~w1623 & w11723) | (w11722 & w11723);
assign w1791 = ~w1634 & ~w1643;
assign w1792 = ~w1790 & w1791;
assign w1793 = ~w1731 & ~w1792;
assign w1794 = w1276 & ~w1763;
assign w1795 = ~w1764 & ~w1794;
assign w1796 = pi0236 & pi1099;
assign w1797 = ~pi0218 & ~pi1099;
assign w1798 = ~w1796 & ~w1797;
assign w1799 = ~pi1260 & ~pi1313;
assign w1800 = pi1260 & pi1313;
assign w1801 = ~w1799 & ~w1800;
assign w1802 = pi1123 & ~pi1317;
assign w1803 = ~pi1123 & pi1317;
assign w1804 = pi1026 & ~pi1044;
assign w1805 = ~pi1026 & pi1044;
assign w1806 = ~pi1262 & ~pi1318;
assign w1807 = pi1262 & pi1318;
assign w1808 = ~w1806 & ~w1807;
assign w1809 = ~w1802 & ~w1803;
assign w1810 = ~w1804 & ~w1805;
assign w1811 = w1809 & w1810;
assign w1812 = ~w1801 & ~w1808;
assign w1813 = w1811 & w1812;
assign w1814 = ~pi1134 & ~pi1313;
assign w1815 = pi1134 & pi1313;
assign w1816 = ~w1814 & ~w1815;
assign w1817 = pi1135 & ~pi1317;
assign w1818 = ~pi1135 & pi1317;
assign w1819 = pi1044 & ~pi1054;
assign w1820 = ~pi1044 & pi1054;
assign w1821 = ~pi1136 & ~pi1318;
assign w1822 = pi1136 & pi1318;
assign w1823 = ~w1821 & ~w1822;
assign w1824 = ~w1817 & ~w1818;
assign w1825 = ~w1819 & ~w1820;
assign w1826 = w1824 & w1825;
assign w1827 = ~w1816 & ~w1823;
assign w1828 = w1826 & w1827;
assign w1829 = ~w1813 & ~w1828;
assign w1830 = ~pi1253 & ~pi1313;
assign w1831 = pi1253 & pi1313;
assign w1832 = ~w1830 & ~w1831;
assign w1833 = pi1148 & ~pi1317;
assign w1834 = ~pi1148 & pi1317;
assign w1835 = pi1044 & ~pi1146;
assign w1836 = ~pi1044 & pi1146;
assign w1837 = ~pi1147 & ~pi1318;
assign w1838 = pi1147 & pi1318;
assign w1839 = ~w1837 & ~w1838;
assign w1840 = ~w1833 & ~w1834;
assign w1841 = ~w1835 & ~w1836;
assign w1842 = w1840 & w1841;
assign w1843 = ~w1832 & ~w1839;
assign w1844 = w1842 & w1843;
assign w1845 = ~pi1044 & ~pi1115;
assign w1846 = pi1044 & pi1115;
assign w1847 = ~w1845 & ~w1846;
assign w1848 = pi1070 & ~pi1318;
assign w1849 = ~pi1070 & pi1318;
assign w1850 = pi1117 & ~pi1317;
assign w1851 = ~pi1117 & pi1317;
assign w1852 = ~pi1116 & ~pi1313;
assign w1853 = pi1116 & pi1313;
assign w1854 = ~w1852 & ~w1853;
assign w1855 = ~w1848 & ~w1849;
assign w1856 = ~w1850 & ~w1851;
assign w1857 = w1855 & w1856;
assign w1858 = ~w1847 & ~w1854;
assign w1859 = w1857 & w1858;
assign w1860 = w1829 & w11724;
assign w1861 = pi0125 & w1860;
assign w1862 = w1829 & w1844;
assign w1863 = w1829 & w11725;
assign w1864 = pi0264 & w1813;
assign w1865 = w1829 & w11726;
assign w1866 = pi0266 & w1865;
assign w1867 = ~w1813 & w1828;
assign w1868 = pi0249 & w1867;
assign w1869 = ~w1864 & ~w1868;
assign w1870 = ~w1863 & w1869;
assign w1871 = ~w1861 & w1870;
assign w1872 = ~w1866 & w1871;
assign w1873 = pi0259 & pi1459;
assign w1874 = ~pi0128 & ~w1873;
assign w1875 = w1769 & ~w1874;
assign w1876 = pi0259 & pi1480;
assign w1877 = ~pi0129 & ~w1876;
assign w1878 = w1773 & ~w1877;
assign w1879 = pi0259 & pi1430;
assign w1880 = ~pi0130 & ~w1879;
assign w1881 = w1777 & ~w1880;
assign w1882 = pi0259 & pi1447;
assign w1883 = ~pi0131 & ~w1882;
assign w1884 = w1783 & ~w1883;
assign w1885 = pi1424 & pi1747;
assign w1886 = ~pi0136 & pi0222;
assign w1887 = w1885 & ~w1886;
assign w1888 = pi0468 & pi1421;
assign w1889 = pi0380 & pi1468;
assign w1890 = pi0562 & pi1456;
assign w1891 = ~pi0380 & ~pi1468;
assign w1892 = ~pi0533 & ~pi1455;
assign w1893 = pi0533 & pi1455;
assign w1894 = pi0483 & pi1454;
assign w1895 = ~pi0485 & ~pi1490;
assign w1896 = ~pi0483 & ~pi1454;
assign w1897 = pi0485 & pi1490;
assign w1898 = pi0549 & pi1513;
assign w1899 = ~pi0549 & ~pi1513;
assign w1900 = ~pi0567 & ~pi1488;
assign w1901 = pi0567 & pi1488;
assign w1902 = pi0622 & pi1482;
assign w1903 = ~pi0622 & ~pi1482;
assign w1904 = ~pi0587 & ~pi1489;
assign w1905 = pi0587 & pi1489;
assign w1906 = ~pi0618 & ~pi1637;
assign w1907 = ~pi0506 & ~pi1678;
assign w1908 = ~w1906 & ~w1907;
assign w1909 = pi0618 & pi1637;
assign w1910 = ~w1905 & ~w1909;
assign w1911 = ~w1908 & w1910;
assign w1912 = ~w1903 & ~w1904;
assign w1913 = ~w1901 & ~w1902;
assign w1914 = (w1913 & w1911) | (w1913 & w11727) | (w1911 & w11727);
assign w1915 = ~w1899 & ~w1900;
assign w1916 = ~w1897 & ~w1898;
assign w1917 = ~w1895 & ~w1896;
assign w1918 = (~w1914 & w11729) | (~w1914 & w11730) | (w11729 & w11730);
assign w1919 = ~w1893 & ~w1894;
assign w1920 = ~w1891 & ~w1892;
assign w1921 = ~w1889 & ~w1890;
assign w1922 = ~pi0468 & ~pi1421;
assign w1923 = ~pi0562 & ~pi1456;
assign w1924 = ~w1922 & ~w1923;
assign w1925 = (w1918 & w11734) | (w1918 & w11735) | (w11734 & w11735);
assign w1926 = ~w1888 & ~w1925;
assign w1927 = pi0352 & pi0725;
assign w1928 = w1174 & w11736;
assign w1929 = pi0244 & ~w1927;
assign w1930 = ~w1928 & w1929;
assign w1931 = (w1623 & w11737) | (w1623 & w11738) | (w11737 & w11738);
assign w1932 = ~w1790 & ~w1931;
assign w1933 = ~w1624 & ~w1635;
assign w1934 = ~w1623 & w1630;
assign w1935 = (w1623 & w11740) | (w1623 & w11741) | (w11740 & w11741);
assign w1936 = (~w1623 & w11742) | (~w1623 & w11743) | (w11742 & w11743);
assign w1937 = ~w1935 & ~w1936;
assign w1938 = ~pi0213 & ~pi0261;
assign w1939 = ~pi0141 & pi0261;
assign w1940 = ~w1938 & ~w1939;
assign w1941 = ~pi0621 & ~pi1449;
assign w1942 = ~pi0645 & ~pi1441;
assign w1943 = pi0358 & pi1436;
assign w1944 = ~pi0358 & ~pi1436;
assign w1945 = ~pi0623 & ~pi1486;
assign w1946 = pi0566 & pi1484;
assign w1947 = pi0623 & pi1486;
assign w1948 = ~pi0566 & ~pi1484;
assign w1949 = ~pi0569 & ~pi1475;
assign w1950 = pi0648 & pi1515;
assign w1951 = pi0569 & pi1475;
assign w1952 = ~pi0648 & ~pi1515;
assign w1953 = ~pi0650 & ~pi1535;
assign w1954 = pi0654 & pi1525;
assign w1955 = pi0650 & pi1535;
assign w1956 = ~pi0654 & ~pi1525;
assign w1957 = ~pi0653 & ~pi1536;
assign w1958 = pi0662 & pi1567;
assign w1959 = pi0653 & pi1536;
assign w1960 = ~pi0662 & ~pi1567;
assign w1961 = ~pi0586 & ~pi1703;
assign w1962 = ~w1960 & ~w1961;
assign w1963 = ~w1958 & ~w1959;
assign w1964 = ~w1962 & w1963;
assign w1965 = ~w1956 & ~w1957;
assign w1966 = ~w1954 & ~w1955;
assign w1967 = (w1966 & w1964) | (w1966 & w11744) | (w1964 & w11744);
assign w1968 = ~w1952 & ~w1953;
assign w1969 = ~w1950 & ~w1951;
assign w1970 = ~w1948 & ~w1949;
assign w1971 = (~w1967 & w11746) | (~w1967 & w11747) | (w11746 & w11747);
assign w1972 = ~w1946 & ~w1947;
assign w1973 = ~w1944 & ~w1945;
assign w1974 = (w1973 & w1971) | (w1973 & w11748) | (w1971 & w11748);
assign w1975 = pi0621 & pi1449;
assign w1976 = pi0645 & pi1441;
assign w1977 = ~w1975 & ~w1976;
assign w1978 = (~w1974 & w11750) | (~w1974 & w11751) | (w11750 & w11751);
assign w1979 = ~w1941 & ~w1978;
assign w1980 = pi0381 & pi1434;
assign w1981 = pi0470 & pi1438;
assign w1982 = ~pi0379 & ~pi1435;
assign w1983 = pi0379 & pi1435;
assign w1984 = pi0466 & pi1462;
assign w1985 = ~pi0466 & ~pi1462;
assign w1986 = ~pi0386 & ~pi1461;
assign w1987 = pi0386 & pi1461;
assign w1988 = pi0387 & pi1474;
assign w1989 = ~pi0480 & ~pi1512;
assign w1990 = ~pi0387 & ~pi1474;
assign w1991 = pi0480 & pi1512;
assign w1992 = pi0484 & pi1507;
assign w1993 = ~pi0509 & ~pi1497;
assign w1994 = ~pi0484 & ~pi1507;
assign w1995 = pi0509 & pi1497;
assign w1996 = pi0508 & pi1509;
assign w1997 = ~pi0508 & ~pi1509;
assign w1998 = ~pi0507 & ~pi1565;
assign w1999 = pi0507 & pi1565;
assign w2000 = ~pi0408 & ~pi1702;
assign w2001 = ~w1999 & w2000;
assign w2002 = ~w1997 & ~w1998;
assign w2003 = ~w2001 & w2002;
assign w2004 = ~w1995 & ~w1996;
assign w2005 = ~w1993 & ~w1994;
assign w2006 = (w2005 & w2003) | (w2005 & w11752) | (w2003 & w11752);
assign w2007 = ~w1991 & ~w1992;
assign w2008 = ~w1989 & ~w1990;
assign w2009 = ~w1987 & ~w1988;
assign w2010 = (~w2006 & w11754) | (~w2006 & w11755) | (w11754 & w11755);
assign w2011 = ~w1985 & ~w1986;
assign w2012 = ~w1983 & ~w1984;
assign w2013 = (w2012 & w2010) | (w2012 & w11756) | (w2010 & w11756);
assign w2014 = ~pi0381 & ~pi1434;
assign w2015 = ~pi0470 & ~pi1438;
assign w2016 = ~w2014 & ~w2015;
assign w2017 = (~w2013 & w11758) | (~w2013 & w11759) | (w11758 & w11759);
assign w2018 = ~w1980 & ~w2017;
assign w2019 = ~pi0232 & ~pi0261;
assign w2020 = ~pi0144 & pi0261;
assign w2021 = ~w2019 & ~w2020;
assign w2022 = ~pi0211 & ~pi0261;
assign w2023 = ~pi0145 & pi0261;
assign w2024 = ~w2022 & ~w2023;
assign w2025 = ~pi0230 & ~pi0261;
assign w2026 = ~pi0146 & pi0261;
assign w2027 = ~w2025 & ~w2026;
assign w2028 = ~pi0220 & ~pi0261;
assign w2029 = ~pi0147 & pi0261;
assign w2030 = ~w2028 & ~w2029;
assign w2031 = ~pi0097 & pi1747;
assign w2032 = ~pi0121 & w2031;
assign w2033 = w238 & w2032;
assign w2034 = ~w815 & w11760;
assign w2035 = ~w2033 & ~w2034;
assign w2036 = ~pi0429 & pi1747;
assign w2037 = pi0706 & pi1747;
assign w2038 = ~w2036 & ~w2037;
assign w2039 = pi0186 & ~pi0429;
assign w2040 = pi0153 & w2039;
assign w2041 = ~pi0153 & ~w2039;
assign w2042 = ~w2038 & ~w2040;
assign w2043 = ~w2041 & w2042;
assign w2044 = pi0224 & pi1099;
assign w2045 = ~pi0353 & ~pi1099;
assign w2046 = ~w2044 & ~w2045;
assign w2047 = pi0243 & pi1099;
assign w2048 = ~pi0280 & ~pi1099;
assign w2049 = ~w2047 & ~w2048;
assign w2050 = ~pi0229 & ~pi0261;
assign w2051 = ~pi0156 & pi0261;
assign w2052 = ~w2050 & ~w2051;
assign w2053 = ~pi0201 & ~pi0261;
assign w2054 = ~pi0157 & pi0261;
assign w2055 = ~w2053 & ~w2054;
assign w2056 = ~pi0197 & ~pi0261;
assign w2057 = ~pi0158 & pi0261;
assign w2058 = ~w2056 & ~w2057;
assign w2059 = ~pi0202 & ~pi0261;
assign w2060 = ~pi0159 & pi0261;
assign w2061 = ~w2059 & ~w2060;
assign w2062 = ~pi0203 & ~pi0261;
assign w2063 = ~pi0160 & pi0261;
assign w2064 = ~w2062 & ~w2063;
assign w2065 = ~pi0204 & ~pi0261;
assign w2066 = ~pi0161 & pi0261;
assign w2067 = ~w2065 & ~w2066;
assign w2068 = ~pi0205 & ~pi0261;
assign w2069 = ~pi0162 & pi0261;
assign w2070 = ~w2068 & ~w2069;
assign w2071 = ~pi0206 & ~pi0261;
assign w2072 = ~pi0163 & pi0261;
assign w2073 = ~w2071 & ~w2072;
assign w2074 = ~pi0225 & ~pi0261;
assign w2075 = ~pi0164 & pi0261;
assign w2076 = ~w2074 & ~w2075;
assign w2077 = ~pi0219 & ~pi0261;
assign w2078 = ~pi0165 & pi0261;
assign w2079 = ~w2077 & ~w2078;
assign w2080 = ~pi0226 & ~pi0261;
assign w2081 = ~pi0166 & pi0261;
assign w2082 = ~w2080 & ~w2081;
assign w2083 = ~pi0227 & ~pi0261;
assign w2084 = ~pi0167 & pi0261;
assign w2085 = ~w2083 & ~w2084;
assign w2086 = ~pi0246 & ~pi0261;
assign w2087 = ~pi0168 & pi0261;
assign w2088 = ~w2086 & ~w2087;
assign w2089 = ~pi0207 & ~pi0261;
assign w2090 = ~pi0169 & pi0261;
assign w2091 = ~w2089 & ~w2090;
assign w2092 = ~pi0209 & ~pi0261;
assign w2093 = ~pi0170 & pi0261;
assign w2094 = ~w2092 & ~w2093;
assign w2095 = ~pi0208 & ~pi0261;
assign w2096 = ~pi0171 & pi0261;
assign w2097 = ~w2095 & ~w2096;
assign w2098 = ~pi0210 & ~pi0261;
assign w2099 = ~pi0172 & pi0261;
assign w2100 = ~w2098 & ~w2099;
assign w2101 = ~pi0217 & ~pi0261;
assign w2102 = ~pi0173 & pi0261;
assign w2103 = ~w2101 & ~w2102;
assign w2104 = ~pi0212 & ~pi0261;
assign w2105 = ~pi0174 & pi0261;
assign w2106 = ~w2104 & ~w2105;
assign w2107 = ~pi0247 & ~pi0261;
assign w2108 = ~pi0175 & pi0261;
assign w2109 = ~w2107 & ~w2108;
assign w2110 = ~pi0214 & ~pi0261;
assign w2111 = ~pi0176 & pi0261;
assign w2112 = ~w2110 & ~w2111;
assign w2113 = ~pi0235 & ~pi0261;
assign w2114 = ~pi0177 & pi0261;
assign w2115 = ~w2113 & ~w2114;
assign w2116 = ~pi0231 & ~pi0261;
assign w2117 = ~pi0178 & pi0261;
assign w2118 = ~w2116 & ~w2117;
assign w2119 = ~pi0233 & ~pi0261;
assign w2120 = ~pi0179 & pi0261;
assign w2121 = ~w2119 & ~w2120;
assign w2122 = ~pi0234 & ~pi0261;
assign w2123 = ~pi0180 & pi0261;
assign w2124 = ~w2122 & ~w2123;
assign w2125 = ~pi0248 & ~pi0261;
assign w2126 = ~pi0181 & pi0261;
assign w2127 = ~w2125 & ~w2126;
assign w2128 = ~pi0228 & ~pi0261;
assign w2129 = ~pi0182 & pi0261;
assign w2130 = ~w2128 & ~w2129;
assign w2131 = pi0284 & pi0306;
assign w2132 = pi1737 & ~pi1739;
assign w2133 = pi1629 & w2132;
assign w2134 = w2132 & w11761;
assign w2135 = ~pi0984 & ~pi1045;
assign w2136 = ~pi0773 & ~pi0937;
assign w2137 = ~pi0954 & ~pi1021;
assign w2138 = w2137 & w11762;
assign w2139 = ~pi0760 & w2138;
assign w2140 = w2138 & w11763;
assign w2141 = ~pi0916 & ~pi1046;
assign w2142 = w2140 & w11764;
assign w2143 = w2140 & w11765;
assign w2144 = pi0971 & ~pi1019;
assign w2145 = w2143 & w11766;
assign w2146 = w2143 & w11767;
assign w2147 = ~pi0971 & ~pi1019;
assign w2148 = w2147 & w11768;
assign w2149 = w2135 & w2148;
assign w2150 = w2140 & w2149;
assign w2151 = ~pi0916 & pi1046;
assign w2152 = pi0276 & w2151;
assign w2153 = w2133 & w2152;
assign w2154 = pi0916 & ~pi1046;
assign w2155 = pi0724 & pi0960;
assign w2156 = ~pi1345 & w2155;
assign w2157 = w2155 & w11769;
assign w2158 = w2154 & w2157;
assign w2159 = ~w2153 & ~w2158;
assign w2160 = w2150 & ~w2159;
assign w2161 = ~w2146 & ~w2160;
assign w2162 = ~pi0971 & pi1019;
assign w2163 = w2143 & w11770;
assign w2164 = pi0262 & w2163;
assign w2165 = w2148 & w11764;
assign w2166 = w2136 & w2165;
assign w2167 = w2165 & w11763;
assign w2168 = w2165 & w11771;
assign w2169 = ~pi1677 & w2168;
assign w2170 = pi0954 & ~pi1021;
assign w2171 = w2168 & w11772;
assign w2172 = w2168 & w11773;
assign w2173 = w2137 & w2168;
assign w2174 = w2168 & w11774;
assign w2175 = w2147 & w11775;
assign w2176 = w2142 & w2175;
assign w2177 = w2142 & w11776;
assign w2178 = pi0785 & pi0916;
assign w2179 = pi1479 & w2178;
assign w2180 = w2178 & w11777;
assign w2181 = w2150 & w2180;
assign w2182 = ~w2177 & ~w2181;
assign w2183 = ~w2174 & w2182;
assign w2184 = w2183 & w11778;
assign w2185 = w2161 & w2184;
assign w2186 = ~pi0300 & ~pi0301;
assign w2187 = ~pi0302 & pi0303;
assign w2188 = ~pi0304 & ~pi0305;
assign w2189 = w2187 & w2188;
assign w2190 = w2131 & w2186;
assign w2191 = w2189 & w2190;
assign w2192 = w2185 & w2191;
assign w2193 = pi0665 & pi1448;
assign w2194 = pi0664 & pi1469;
assign w2195 = pi0712 & pi1485;
assign w2196 = pi0359 & pi1467;
assign w2197 = ~pi0675 & ~pi1483;
assign w2198 = ~pi0712 & ~pi1485;
assign w2199 = pi0678 & pi1514;
assign w2200 = pi0675 & pi1483;
assign w2201 = ~pi0678 & ~pi1514;
assign w2202 = ~pi0714 & ~pi1537;
assign w2203 = pi0714 & pi1537;
assign w2204 = pi0717 & pi1533;
assign w2205 = ~pi0717 & ~pi1533;
assign w2206 = ~pi0708 & ~pi1524;
assign w2207 = pi0708 & pi1524;
assign w2208 = pi0719 & pi1545;
assign w2209 = ~pi0719 & ~pi1545;
assign w2210 = ~pi0718 & ~pi1566;
assign w2211 = pi0718 & pi1566;
assign w2212 = ~pi0697 & ~pi1704;
assign w2213 = ~w2211 & w2212;
assign w2214 = ~w2209 & ~w2210;
assign w2215 = ~w2213 & w2214;
assign w2216 = ~w2207 & ~w2208;
assign w2217 = ~w2205 & ~w2206;
assign w2218 = (w2217 & w2215) | (w2217 & w11779) | (w2215 & w11779);
assign w2219 = ~w2203 & ~w2204;
assign w2220 = ~w2201 & ~w2202;
assign w2221 = ~w2199 & ~w2200;
assign w2222 = (~w2218 & w11781) | (~w2218 & w11782) | (w11781 & w11782);
assign w2223 = ~w2197 & ~w2198;
assign w2224 = ~w2195 & ~w2196;
assign w2225 = ~pi0359 & ~pi1467;
assign w2226 = (~w2222 & w11784) | (~w2222 & w11785) | (w11784 & w11785);
assign w2227 = ~pi0665 & ~pi1448;
assign w2228 = ~pi0664 & ~pi1469;
assign w2229 = ~w2227 & ~w2228;
assign w2230 = (w2229 & w2226) | (w2229 & w11786) | (w2226 & w11786);
assign w2231 = ~w2193 & ~w2230;
assign w2232 = w2039 & w11787;
assign w2233 = ~pi0185 & ~w2232;
assign w2234 = pi0185 & w2232;
assign w2235 = ~w2038 & ~w2233;
assign w2236 = ~w2234 & w2235;
assign w2237 = ~pi0186 & ~w2036;
assign w2238 = ~w2038 & ~w2039;
assign w2239 = ~w2237 & w2238;
assign w2240 = (w2032 & ~w232) | (w2032 & w11788) | (~w232 & w11788);
assign w2241 = ~w815 & w11789;
assign w2242 = ~w2240 & ~w2241;
assign w2243 = ~pi0281 & ~pi1099;
assign w2244 = (~pi0195 & ~w2039) | (~pi0195 & w11790) | (~w2039 & w11790);
assign w2245 = ~w2038 & ~w2232;
assign w2246 = ~w2244 & w2245;
assign w2247 = ~pi0196 & ~pi0261;
assign w2248 = (pi1579 & ~w219) | (pi1579 & w11791) | (~w219 & w11791);
assign w2249 = w219 & w11792;
assign w2250 = ~pi1709 & w2249;
assign w2251 = ~pi1579 & pi1818;
assign w2252 = (~w2251 & ~w2248) | (~w2251 & w11793) | (~w2248 & w11793);
assign w2253 = ~w2250 & w2252;
assign w2254 = pi1570 & w374;
assign w2255 = pi1570 & pi1580;
assign w2256 = ~pi0771 & ~w2255;
assign w2257 = ~pi0801 & pi1568;
assign w2258 = pi1582 & w2257;
assign w2259 = ~w2256 & w2258;
assign w2260 = ~w2254 & ~w2259;
assign w2261 = w358 & ~w2260;
assign w2262 = w228 & w2032;
assign w2263 = ~w815 & w11794;
assign w2264 = ~w2262 & ~w2263;
assign w2265 = ~w1563 & w1568;
assign w2266 = (~w1567 & w1563) | (~w1567 & w11795) | (w1563 & w11795);
assign w2267 = ~w2265 & ~w2266;
assign w2268 = pi0201 & w2248;
assign w2269 = ~pi1579 & pi1816;
assign w2270 = (~w2269 & ~w2249) | (~w2269 & w11796) | (~w2249 & w11796);
assign w2271 = ~w2268 & w2270;
assign w2272 = ~pi1714 & w2249;
assign w2273 = ~pi1579 & pi1817;
assign w2274 = (~w2273 & ~w2248) | (~w2273 & w11797) | (~w2248 & w11797);
assign w2275 = ~w2272 & w2274;
assign w2276 = ~pi1717 & w2249;
assign w2277 = ~pi1579 & pi1819;
assign w2278 = (~w2277 & ~w2248) | (~w2277 & w11798) | (~w2248 & w11798);
assign w2279 = ~w2276 & w2278;
assign w2280 = pi0204 & w2248;
assign w2281 = ~pi1579 & pi1820;
assign w2282 = (~w2281 & ~w2249) | (~w2281 & w11799) | (~w2249 & w11799);
assign w2283 = ~w2280 & w2282;
assign w2284 = pi0205 & w2248;
assign w2285 = ~pi1579 & pi1821;
assign w2286 = (~w2285 & ~w2249) | (~w2285 & w11800) | (~w2249 & w11800);
assign w2287 = ~w2284 & w2286;
assign w2288 = ~pi0152 & pi0199;
assign w2289 = w2288 & w11801;
assign w2290 = (pi1579 & ~w2288) | (pi1579 & w11802) | (~w2288 & w11802);
assign w2291 = pi0206 & w2290;
assign w2292 = ~pi1579 & pi1823;
assign w2293 = (~w2292 & ~w2289) | (~w2292 & w11803) | (~w2289 & w11803);
assign w2294 = ~w2291 & w2293;
assign w2295 = ~pi1711 & w2289;
assign w2296 = ~pi1579 & pi1829;
assign w2297 = (~w2296 & ~w2290) | (~w2296 & w11804) | (~w2290 & w11804);
assign w2298 = ~w2295 & w2297;
assign w2299 = pi0874 & w226;
assign w2300 = w226 & w11801;
assign w2301 = (pi1579 & ~w226) | (pi1579 & w11802) | (~w226 & w11802);
assign w2302 = pi0208 & w2301;
assign w2303 = ~pi1579 & pi1831;
assign w2304 = (~w2303 & ~w2300) | (~w2303 & w11805) | (~w2300 & w11805);
assign w2305 = ~w2302 & w2304;
assign w2306 = ~pi1712 & w2300;
assign w2307 = ~pi1579 & pi1830;
assign w2308 = (~w2307 & ~w2301) | (~w2307 & w11806) | (~w2301 & w11806);
assign w2309 = ~w2306 & w2308;
assign w2310 = pi0210 & w2301;
assign w2311 = ~pi1579 & pi1832;
assign w2312 = (~w2311 & ~w2300) | (~w2311 & w11807) | (~w2300 & w11807);
assign w2313 = ~w2310 & w2312;
assign w2314 = pi0211 & w2301;
assign w2315 = ~pi1579 & pi1833;
assign w2316 = (~w2315 & ~w2300) | (~w2315 & w11808) | (~w2300 & w11808);
assign w2317 = ~w2314 & w2316;
assign w2318 = ~pi1717 & w2300;
assign w2319 = ~pi1579 & pi1835;
assign w2320 = (~w2319 & ~w2301) | (~w2319 & w11809) | (~w2301 & w11809);
assign w2321 = ~w2318 & w2320;
assign w2322 = pi0213 & w2301;
assign w2323 = ~pi1579 & pi1836;
assign w2324 = (~w2323 & ~w2300) | (~w2323 & w11810) | (~w2300 & w11810);
assign w2325 = ~w2322 & w2324;
assign w2326 = pi0214 & w2301;
assign w2327 = ~pi1579 & pi1837;
assign w2328 = (~w2327 & ~w2300) | (~w2327 & w11811) | (~w2300 & w11811);
assign w2329 = ~w2326 & w2328;
assign w2330 = (~w1602 & w1610) | (~w1602 & w11812) | (w1610 & w11812);
assign w2331 = w1618 & ~w2330;
assign w2332 = (~w1617 & ~w1614) | (~w1617 & w11813) | (~w1614 & w11813);
assign w2333 = ~w1623 & ~w2332;
assign w2334 = (~w1629 & w1623) | (~w1629 & w11814) | (w1623 & w11814);
assign w2335 = ~w1934 & ~w2334;
assign w2336 = pi0217 & w2301;
assign w2337 = ~pi1579 & pi1834;
assign w2338 = (~w2337 & ~w2300) | (~w2337 & w11815) | (~w2300 & w11815);
assign w2339 = ~w2336 & w2338;
assign w2340 = ~w1557 & ~w1564;
assign w2341 = w1556 & w11816;
assign w2342 = (~w2340 & ~w1556) | (~w2340 & w11817) | (~w1556 & w11817);
assign w2343 = ~w2341 & ~w2342;
assign w2344 = ~pi1714 & w2289;
assign w2345 = ~pi1579 & pi1825;
assign w2346 = (~w2345 & ~w2290) | (~w2345 & w11818) | (~w2290 & w11818);
assign w2347 = ~w2344 & w2346;
assign w2348 = pi0220 & w2290;
assign w2349 = ~pi1579 & pi1822;
assign w2350 = (~w2349 & ~w2289) | (~w2349 & w11819) | (~w2289 & w11819);
assign w2351 = ~w2348 & w2350;
assign w2352 = pi0257 & pi0874;
assign w2353 = pi0237 & w2352;
assign w2354 = w2352 & w11820;
assign w2355 = w2354 & w11821;
assign w2356 = (~pi0221 & ~w2354) | (~pi0221 & w11822) | (~w2354 & w11822);
assign w2357 = w2354 & w11823;
assign w2358 = w2031 & ~w2356;
assign w2359 = ~w2357 & w2358;
assign w2360 = pi0242 & pi1099;
assign w2361 = ~pi0355 & ~pi1099;
assign w2362 = ~w2360 & ~w2361;
assign w2363 = w2357 & w11824;
assign w2364 = w2357 & w11826;
assign w2365 = (w2357 & w11827) | (w2357 & w11828) | (w11827 & w11828);
assign w2366 = ~w2364 & w2365;
assign w2367 = pi0225 & w2290;
assign w2368 = ~pi1579 & pi1824;
assign w2369 = (~w2368 & ~w2289) | (~w2368 & w11829) | (~w2289 & w11829);
assign w2370 = ~w2367 & w2369;
assign w2371 = ~pi1709 & w2289;
assign w2372 = ~pi1579 & pi1826;
assign w2373 = (~w2372 & ~w2290) | (~w2372 & w11830) | (~w2290 & w11830);
assign w2374 = ~w2371 & w2373;
assign w2375 = ~pi1717 & w2289;
assign w2376 = ~pi1579 & pi1827;
assign w2377 = (~w2376 & ~w2290) | (~w2376 & w11831) | (~w2290 & w11831);
assign w2378 = ~w2375 & w2377;
assign w2379 = pi0228 & w2248;
assign w2380 = ~pi1579 & pi1815;
assign w2381 = (~w2380 & ~w2249) | (~w2380 & w11832) | (~w2249 & w11832);
assign w2382 = ~w2379 & w2381;
assign w2383 = ~pi0152 & ~pi0199;
assign w2384 = w2383 & w11801;
assign w2385 = (pi1579 & ~w2383) | (pi1579 & w11802) | (~w2383 & w11802);
assign w2386 = pi0229 & w2385;
assign w2387 = ~pi1579 & pi1806;
assign w2388 = (~w2387 & ~w2384) | (~w2387 & w11833) | (~w2384 & w11833);
assign w2389 = ~w2386 & w2388;
assign w2390 = ~pi1716 & w2384;
assign w2391 = ~pi1579 & pi1807;
assign w2392 = (~w2391 & ~w2385) | (~w2391 & w11834) | (~w2385 & w11834);
assign w2393 = ~w2390 & w2392;
assign w2394 = ~pi1709 & w2384;
assign w2395 = ~pi1579 & pi1810;
assign w2396 = (~w2395 & ~w2385) | (~w2395 & w11835) | (~w2385 & w11835);
assign w2397 = ~w2394 & w2396;
assign w2398 = ~pi1717 & w2384;
assign w2399 = ~pi1579 & pi1811;
assign w2400 = (~w2399 & ~w2385) | (~w2399 & w11836) | (~w2385 & w11836);
assign w2401 = ~w2398 & w2400;
assign w2402 = pi0233 & w2385;
assign w2403 = ~pi1579 & pi1812;
assign w2404 = (~w2403 & ~w2384) | (~w2403 & w11837) | (~w2384 & w11837);
assign w2405 = ~w2402 & w2404;
assign w2406 = ~pi1711 & w2384;
assign w2407 = ~pi1579 & pi1813;
assign w2408 = (~w2407 & ~w2385) | (~w2407 & w11838) | (~w2385 & w11838);
assign w2409 = ~w2406 & w2408;
assign w2410 = pi0235 & w2385;
assign w2411 = ~pi1579 & pi1809;
assign w2412 = (~w2411 & ~w2384) | (~w2411 & w11839) | (~w2384 & w11839);
assign w2413 = ~w2410 & w2412;
assign w2414 = w2357 & w11840;
assign w2415 = pi0236 & w2414;
assign w2416 = (w2031 & w2414) | (w2031 & w11841) | (w2414 & w11841);
assign w2417 = ~w2415 & w2416;
assign w2418 = ~pi0237 & ~w2352;
assign w2419 = w2031 & ~w2353;
assign w2420 = ~w2418 & w2419;
assign w2421 = (~pi0238 & ~w2352) | (~pi0238 & w11842) | (~w2352 & w11842);
assign w2422 = w2031 & ~w2354;
assign w2423 = ~w2421 & w2422;
assign w2424 = ~pi0239 & ~w2354;
assign w2425 = (w2031 & ~w2354) | (w2031 & w11843) | (~w2354 & w11843);
assign w2426 = ~w2424 & w2425;
assign w2427 = (~pi0240 & ~w2354) | (~pi0240 & w11844) | (~w2354 & w11844);
assign w2428 = w2031 & ~w2355;
assign w2429 = ~w2427 & w2428;
assign w2430 = ~pi0241 & ~w2357;
assign w2431 = (w2031 & ~w2357) | (w2031 & w11845) | (~w2357 & w11845);
assign w2432 = ~w2430 & w2431;
assign w2433 = (~pi0242 & ~w2357) | (~pi0242 & w11846) | (~w2357 & w11846);
assign w2434 = w2031 & ~w2363;
assign w2435 = ~w2433 & w2434;
assign w2436 = (~pi0243 & ~w2357) | (~pi0243 & w11847) | (~w2357 & w11847);
assign w2437 = w2031 & ~w2414;
assign w2438 = ~w2436 & w2437;
assign w2439 = pi0236 & w1281;
assign w2440 = pi0243 & w1326;
assign w2441 = ~pi0224 & ~w1332;
assign w2442 = ~pi0243 & ~w1326;
assign w2443 = pi0242 & w1382;
assign w2444 = pi0224 & w1332;
assign w2445 = ~pi0241 & ~w1376;
assign w2446 = ~pi0242 & ~w1382;
assign w2447 = ~pi0221 & ~w1370;
assign w2448 = ~pi0240 & ~w1320;
assign w2449 = pi0239 & w1359;
assign w2450 = pi0240 & w1320;
assign w2451 = ~pi0239 & ~w1359;
assign w2452 = ~pi0238 & ~w1353;
assign w2453 = pi0238 & w1353;
assign w2454 = pi0237 & w1339;
assign w2455 = ~pi0237 & ~w1339;
assign w2456 = pi0257 & w1345;
assign w2457 = ~w2455 & w2456;
assign w2458 = ~w2453 & ~w2454;
assign w2459 = ~w2457 & w2458;
assign w2460 = ~w2451 & ~w2452;
assign w2461 = ~w2449 & ~w2450;
assign w2462 = (w2461 & w2459) | (w2461 & w11848) | (w2459 & w11848);
assign w2463 = ~w2447 & ~w2448;
assign w2464 = pi0241 & w1376;
assign w2465 = pi0221 & w1370;
assign w2466 = ~w2464 & ~w2465;
assign w2467 = ~w2445 & ~w2446;
assign w2468 = (~w2462 & w11850) | (~w2462 & w11851) | (w11850 & w11851);
assign w2469 = ~w2443 & ~w2444;
assign w2470 = ~w2441 & ~w2442;
assign w2471 = ~w2439 & ~w2440;
assign w2472 = (~w2468 & w11853) | (~w2468 & w11854) | (w11853 & w11854);
assign w2473 = (pi0974 & w1281) | (pi0974 & w11855) | (w1281 & w11855);
assign w2474 = w1278 & w2473;
assign w2475 = ~w2472 & w2474;
assign w2476 = ~w1625 & ~w1638;
assign w2477 = (w1623 & w11856) | (w1623 & w11857) | (w11856 & w11857);
assign w2478 = ~w2476 & w2477;
assign w2479 = w2476 & ~w2477;
assign w2480 = ~w2478 & ~w2479;
assign w2481 = pi0246 & w2290;
assign w2482 = ~pi1579 & pi1828;
assign w2483 = (~w2482 & ~w2289) | (~w2482 & w11858) | (~w2289 & w11858);
assign w2484 = ~w2481 & w2483;
assign w2485 = ~pi1713 & w2384;
assign w2486 = ~pi1579 & pi1808;
assign w2487 = (~w2486 & ~w2385) | (~w2486 & w11859) | (~w2385 & w11859);
assign w2488 = ~w2485 & w2487;
assign w2489 = ~pi1712 & w2249;
assign w2490 = ~pi1579 & pi1814;
assign w2491 = (~w2490 & ~w2248) | (~w2490 & w11860) | (~w2248 & w11860);
assign w2492 = ~w2489 & w2491;
assign w2493 = ~pi1127 & ~pi1308;
assign w2494 = pi1127 & pi1308;
assign w2495 = pi1029 & ~pi1420;
assign w2496 = ~pi1029 & pi1420;
assign w2497 = ~pi1076 & pi1444;
assign w2498 = pi1130 & pi1452;
assign w2499 = pi1076 & ~pi1444;
assign w2500 = ~pi1130 & ~pi1452;
assign w2501 = ~pi1083 & ~pi1500;
assign w2502 = pi1083 & pi1500;
assign w2503 = pi1028 & pi1530;
assign w2504 = ~pi1028 & ~pi1530;
assign w2505 = ~pi1129 & pi1552;
assign w2506 = pi1129 & ~pi1552;
assign w2507 = pi1310 & pi1558;
assign w2508 = ~pi1310 & ~pi1558;
assign w2509 = pi1027 & pi1630;
assign w2510 = ~w2508 & w2509;
assign w2511 = ~w2506 & ~w2507;
assign w2512 = ~w2510 & w2511;
assign w2513 = ~w2504 & ~w2505;
assign w2514 = ~w2502 & ~w2503;
assign w2515 = (w2514 & w2512) | (w2514 & w11861) | (w2512 & w11861);
assign w2516 = ~w2500 & ~w2501;
assign w2517 = ~w2498 & ~w2499;
assign w2518 = ~w2496 & ~w2497;
assign w2519 = (~w2515 & w11863) | (~w2515 & w11864) | (w11863 & w11864);
assign w2520 = ~w2494 & ~w2495;
assign w2521 = ~w2519 & w2520;
assign w2522 = ~pi0949 & ~pi0980;
assign w2523 = pi1341 & w2522;
assign w2524 = ~w2493 & w2523;
assign w2525 = ~w2521 & w2524;
assign w2526 = pi0250 & w2037;
assign w2527 = ~pi0706 & pi1747;
assign w2528 = pi1318 & w2527;
assign w2529 = ~w2526 & ~w2528;
assign w2530 = pi0251 & w2037;
assign w2531 = pi1042 & w2527;
assign w2532 = ~w2530 & ~w2531;
assign w2533 = pi0252 & w2037;
assign w2534 = pi1044 & w2527;
assign w2535 = ~w2533 & ~w2534;
assign w2536 = pi0253 & w2037;
assign w2537 = pi1313 & w2527;
assign w2538 = ~w2536 & ~w2537;
assign w2539 = pi0241 & pi1099;
assign w2540 = ~pi0431 & ~pi1099;
assign w2541 = ~w2539 & ~w2540;
assign w2542 = pi0255 & w2037;
assign w2543 = pi1317 & w2527;
assign w2544 = ~w2542 & ~w2543;
assign w2545 = ~pi0256 & pi0354;
assign w2546 = pi0630 & w2545;
assign w2547 = ~pi0257 & ~pi0874;
assign w2548 = w2031 & ~w2352;
assign w2549 = ~w2547 & w2548;
assign w2550 = w2 & w11;
assign w2551 = pi0660 & w3;
assign w2552 = w2550 & w2551;
assign w2553 = w2550 & w11865;
assign w2554 = ~pi0138 & w2553;
assign w2555 = w11 & w11866;
assign w2556 = pi0336 & ~pi0409;
assign w2557 = w2555 & w2556;
assign w2558 = ~w2554 & ~w2557;
assign w2559 = ~pi0874 & ~w2383;
assign w2560 = ~w2558 & w2559;
assign w2561 = pi0089 & pi0625;
assign w2562 = w1598 & w2561;
assign w2563 = w1705 & w2562;
assign w2564 = w1752 & w2563;
assign w2565 = w1606 & w1611;
assign w2566 = ~w1606 & ~w1611;
assign w2567 = ~w2565 & ~w2566;
assign w2568 = ~pi0258 & ~w2299;
assign w2569 = pi0300 & pi0301;
assign w2570 = (pi0303 & w2569) | (pi0303 & w11867) | (w2569 & w11867);
assign w2571 = pi0304 & pi0305;
assign w2572 = w2131 & w2571;
assign w2573 = ~w2570 & w2572;
assign w2574 = w2185 & ~w2573;
assign w2575 = pi0263 & w2037;
assign w2576 = pi1043 & w2527;
assign w2577 = ~w2575 & ~w2576;
assign w2578 = ~pi1119 & ~pi1307;
assign w2579 = pi1119 & pi1307;
assign w2580 = pi1267 & ~pi1432;
assign w2581 = ~pi1267 & pi1432;
assign w2582 = ~pi1270 & pi1443;
assign w2583 = pi1274 & pi1450;
assign w2584 = pi1270 & ~pi1443;
assign w2585 = ~pi1274 & ~pi1450;
assign w2586 = ~pi1121 & ~pi1499;
assign w2587 = pi1272 & pi1529;
assign w2588 = pi1121 & pi1499;
assign w2589 = ~pi1272 & ~pi1529;
assign w2590 = ~pi1023 & pi1553;
assign w2591 = pi1023 & ~pi1553;
assign w2592 = pi1277 & pi1559;
assign w2593 = ~pi1277 & ~pi1559;
assign w2594 = pi1022 & pi1624;
assign w2595 = ~w2593 & w2594;
assign w2596 = ~w2591 & ~w2592;
assign w2597 = ~w2595 & w2596;
assign w2598 = ~w2589 & ~w2590;
assign w2599 = ~w2587 & ~w2588;
assign w2600 = (w2599 & w2597) | (w2599 & w11868) | (w2597 & w11868);
assign w2601 = ~w2585 & ~w2586;
assign w2602 = ~w2583 & ~w2584;
assign w2603 = ~w2581 & ~w2582;
assign w2604 = (~w2600 & w11870) | (~w2600 & w11871) | (w11870 & w11871);
assign w2605 = ~w2579 & ~w2580;
assign w2606 = ~w2604 & w2605;
assign w2607 = ~pi0948 & ~pi0979;
assign w2608 = pi1340 & w2607;
assign w2609 = ~w2578 & w2608;
assign w2610 = ~w2606 & w2609;
assign w2611 = ~pi1139 & ~pi1309;
assign w2612 = pi1139 & pi1309;
assign w2613 = pi1034 & ~pi1433;
assign w2614 = ~pi1034 & pi1433;
assign w2615 = ~pi1265 & pi1446;
assign w2616 = pi1265 & ~pi1446;
assign w2617 = pi1142 & pi1453;
assign w2618 = ~pi1142 & ~pi1453;
assign w2619 = ~pi1033 & ~pi1501;
assign w2620 = pi1033 & pi1501;
assign w2621 = pi1258 & pi1531;
assign w2622 = ~pi1258 & ~pi1531;
assign w2623 = ~pi1141 & pi1555;
assign w2624 = pi1141 & ~pi1555;
assign w2625 = pi1342 & pi1557;
assign w2626 = ~pi1342 & ~pi1557;
assign w2627 = pi1032 & pi1623;
assign w2628 = ~w2626 & w2627;
assign w2629 = ~w2624 & ~w2625;
assign w2630 = ~w2628 & w2629;
assign w2631 = ~w2622 & ~w2623;
assign w2632 = ~w2620 & ~w2621;
assign w2633 = (w2632 & w2630) | (w2632 & w11872) | (w2630 & w11872);
assign w2634 = ~w2618 & ~w2619;
assign w2635 = ~w2616 & ~w2617;
assign w2636 = ~w2614 & ~w2615;
assign w2637 = (~w2633 & w11874) | (~w2633 & w11875) | (w11874 & w11875);
assign w2638 = ~w2612 & ~w2613;
assign w2639 = ~w2637 & w2638;
assign w2640 = ~pi0950 & ~pi0981;
assign w2641 = pi1399 & w2640;
assign w2642 = ~w2611 & w2641;
assign w2643 = ~w2639 & w2642;
assign w2644 = ~pi1102 & ~pi1306;
assign w2645 = pi1102 & pi1306;
assign w2646 = pi1110 & ~pi1431;
assign w2647 = ~pi1110 & pi1431;
assign w2648 = ~pi1109 & pi1442;
assign w2649 = pi1081 & pi1451;
assign w2650 = pi1109 & ~pi1442;
assign w2651 = ~pi1081 & ~pi1451;
assign w2652 = ~pi1108 & ~pi1498;
assign w2653 = pi1108 & pi1498;
assign w2654 = pi1107 & pi1528;
assign w2655 = ~pi1107 & ~pi1528;
assign w2656 = ~pi1106 & pi1554;
assign w2657 = pi1106 & ~pi1554;
assign w2658 = pi1338 & pi1560;
assign w2659 = ~pi1338 & ~pi1560;
assign w2660 = pi1105 & pi1622;
assign w2661 = ~w2659 & w2660;
assign w2662 = ~w2657 & ~w2658;
assign w2663 = ~w2661 & w2662;
assign w2664 = ~w2655 & ~w2656;
assign w2665 = ~w2653 & ~w2654;
assign w2666 = (w2665 & w2663) | (w2665 & w11876) | (w2663 & w11876);
assign w2667 = ~w2651 & ~w2652;
assign w2668 = ~w2649 & ~w2650;
assign w2669 = ~w2647 & ~w2648;
assign w2670 = (~w2666 & w11878) | (~w2666 & w11879) | (w11878 & w11879);
assign w2671 = ~w2645 & ~w2646;
assign w2672 = ~w2670 & w2671;
assign w2673 = ~pi0947 & ~pi0978;
assign w2674 = pi1398 & w2673;
assign w2675 = ~w2644 & w2674;
assign w2676 = ~w2672 & w2675;
assign w2677 = w355 & ~w356;
assign w2678 = pi1233 & w2677;
assign w2679 = ~w1205 & w2678;
assign w2680 = ~pi0268 & ~pi0331;
assign w2681 = ~pi1671 & w2037;
assign w2682 = pi0268 & pi0331;
assign w2683 = ~w2680 & ~w2682;
assign w2684 = w2681 & w2683;
assign w2685 = pi0269 & w2037;
assign w2686 = pi1039 & w2527;
assign w2687 = ~w2685 & ~w2686;
assign w2688 = pi0270 & w2037;
assign w2689 = pi1041 & w2527;
assign w2690 = ~w2688 & ~w2689;
assign w2691 = pi0271 & w2037;
assign w2692 = pi1040 & w2527;
assign w2693 = ~w2691 & ~w2692;
assign w2694 = pi0272 & w2037;
assign w2695 = pi1049 & w2527;
assign w2696 = ~w2694 & ~w2695;
assign w2697 = pi0273 & w2037;
assign w2698 = pi1017 & w2527;
assign w2699 = ~w2697 & ~w2698;
assign w2700 = ~pi0274 & ~w2682;
assign w2701 = pi0274 & w2682;
assign w2702 = w2681 & ~w2700;
assign w2703 = ~w2701 & w2702;
assign w2704 = (~pi0275 & ~w2682) | (~pi0275 & w11880) | (~w2682 & w11880);
assign w2705 = w2682 & w11192;
assign w2706 = w2681 & ~w2704;
assign w2707 = ~w2705 & w2706;
assign w2708 = pi0287 & pi0288;
assign w2709 = (pi0290 & ~w2708) | (pi0290 & w11881) | (~w2708 & w11881);
assign w2710 = pi0291 & ~w2709;
assign w2711 = pi0292 & pi0293;
assign w2712 = (~w2709 & w11883) | (~w2709 & w11884) | (w11883 & w11884);
assign w2713 = w2185 & ~w2712;
assign w2714 = ~w2569 & w11885;
assign w2715 = w2572 & w2714;
assign w2716 = w2185 & ~w2715;
assign w2717 = ~pi0279 & ~pi0294;
assign w2718 = w2184 & w11886;
assign w2719 = pi0279 & pi0294;
assign w2720 = ~w2717 & ~w2719;
assign w2721 = w2718 & w2720;
assign w2722 = ~w1529 & w11887;
assign w2723 = (~pi0101 & w1548) | (~pi0101 & w11888) | (w1548 & w11888);
assign w2724 = ~w2722 & w2723;
assign w2725 = (w1326 & w2724) | (w1326 & w11889) | (w2724 & w11889);
assign w2726 = w1556 & ~w2725;
assign w2727 = ~w1565 & ~w1571;
assign w2728 = ~w1574 & ~w2727;
assign w2729 = (~w2728 & w1563) | (~w2728 & w11890) | (w1563 & w11890);
assign w2730 = ~w1573 & ~w2729;
assign w2731 = (w1603 & ~w1611) | (w1603 & w11891) | (~w1611 & w11891);
assign w2732 = ~w2331 & ~w2731;
assign w2733 = ~w1359 & w2732;
assign w2734 = w1359 & ~w2732;
assign w2735 = ~w2733 & ~w2734;
assign w2736 = ~pi0287 & pi1621;
assign w2737 = ~pi0288 & w2736;
assign w2738 = w2736 & w11892;
assign w2739 = pi0290 & w2738;
assign w2740 = w2738 & w11893;
assign w2741 = w2738 & w11894;
assign w2742 = w2184 & w11895;
assign w2743 = (pi0283 & ~w2738) | (pi0283 & w11896) | (~w2738 & w11896);
assign w2744 = ~w2741 & ~w2743;
assign w2745 = w2742 & w2744;
assign w2746 = pi0183 & pi1534;
assign w2747 = pi0300 & w2746;
assign w2748 = w2746 & w2569;
assign w2749 = pi0302 & w2748;
assign w2750 = w2748 & w11867;
assign w2751 = w2748 & w11897;
assign w2752 = (pi0284 & ~w2748) | (pi0284 & w11898) | (~w2748 & w11898);
assign w2753 = ~w2751 & ~w2752;
assign w2754 = w2185 & w2753;
assign w2755 = ~pi0285 & ~w2705;
assign w2756 = pi0285 & w2705;
assign w2757 = w2681 & ~w2755;
assign w2758 = ~w2756 & w2757;
assign w2759 = ~pi0620 & ~pi1099;
assign w2760 = ~pi0240 & pi1099;
assign w2761 = ~w2759 & ~w2760;
assign w2762 = pi0287 & ~pi1621;
assign w2763 = ~w2736 & ~w2762;
assign w2764 = w2742 & w2763;
assign w2765 = pi0288 & ~w2736;
assign w2766 = ~w2737 & ~w2765;
assign w2767 = w2742 & w2766;
assign w2768 = (pi0289 & ~w2736) | (pi0289 & w11899) | (~w2736 & w11899);
assign w2769 = ~w2738 & ~w2768;
assign w2770 = w2742 & w2769;
assign w2771 = ~pi0290 & ~w2738;
assign w2772 = ~w2739 & ~w2771;
assign w2773 = w2742 & w2772;
assign w2774 = (pi0291 & ~w2738) | (pi0291 & w11900) | (~w2738 & w11900);
assign w2775 = ~w2740 & ~w2774;
assign w2776 = w2742 & w2775;
assign w2777 = ~pi0292 & w2741;
assign w2778 = pi0292 & ~w2741;
assign w2779 = ~w2777 & ~w2778;
assign w2780 = w2742 & w2779;
assign w2781 = (pi0293 & ~w2741) | (pi0293 & w2711) | (~w2741 & w2711);
assign w2782 = w2741 & w10789;
assign w2783 = ~w2781 & ~w2782;
assign w2784 = w2742 & w2783;
assign w2785 = pi0294 & w2718;
assign w2786 = ~pi0295 & w2717;
assign w2787 = pi0295 & ~w2717;
assign w2788 = ~w2786 & ~w2787;
assign w2789 = w2718 & w2788;
assign w2790 = w2717 & w11901;
assign w2791 = ~pi0296 & w2790;
assign w2792 = pi0296 & ~w2790;
assign w2793 = ~w2791 & ~w2792;
assign w2794 = w2718 & w2793;
assign w2795 = w2790 & w11902;
assign w2796 = (pi0297 & ~w2790) | (pi0297 & w11903) | (~w2790 & w11903);
assign w2797 = ~w2795 & ~w2796;
assign w2798 = w2718 & w2797;
assign w2799 = w2790 & w11904;
assign w2800 = (pi0298 & ~w2790) | (pi0298 & w11905) | (~w2790 & w11905);
assign w2801 = ~w2799 & ~w2800;
assign w2802 = w2718 & w2801;
assign w2803 = pi0239 & pi1099;
assign w2804 = ~pi0545 & ~pi1099;
assign w2805 = ~w2803 & ~w2804;
assign w2806 = ~pi0300 & ~w2746;
assign w2807 = ~w2747 & ~w2806;
assign w2808 = w2185 & w2807;
assign w2809 = (~pi0301 & ~w2746) | (~pi0301 & w2186) | (~w2746 & w2186);
assign w2810 = ~w2748 & ~w2809;
assign w2811 = w2185 & w2810;
assign w2812 = ~pi0302 & ~w2748;
assign w2813 = ~w2749 & ~w2812;
assign w2814 = w2185 & w2813;
assign w2815 = (~pi0303 & ~w2748) | (~pi0303 & w11885) | (~w2748 & w11885);
assign w2816 = ~w2750 & ~w2815;
assign w2817 = w2185 & w2816;
assign w2818 = ~pi0306 & w2751;
assign w2819 = w2751 & w11906;
assign w2820 = (pi0304 & ~w2751) | (pi0304 & w11907) | (~w2751 & w11907);
assign w2821 = ~w2819 & ~w2820;
assign w2822 = w2185 & w2821;
assign w2823 = (pi0305 & ~w2751) | (pi0305 & w11908) | (~w2751 & w11908);
assign w2824 = w2751 & w11909;
assign w2825 = ~w2823 & ~w2824;
assign w2826 = w2185 & w2825;
assign w2827 = pi0306 & ~w2751;
assign w2828 = ~w2818 & ~w2827;
assign w2829 = w2185 & w2828;
assign w2830 = (pi0307 & ~w2717) | (pi0307 & w11910) | (~w2717 & w11910);
assign w2831 = ~w2790 & ~w2830;
assign w2832 = w2718 & w2831;
assign w2833 = pi0308 & ~w2799;
assign w2834 = ~pi0308 & w2799;
assign w2835 = ~w2833 & ~w2834;
assign w2836 = w2718 & w2835;
assign w2837 = w2555 & w11912;
assign w2838 = ~pi0096 & pi0121;
assign w2839 = pi0309 & ~pi1090;
assign w2840 = w6 & w2839;
assign w2841 = w6 & w11913;
assign w2842 = w6 & w11914;
assign w2843 = ~pi0138 & ~w2842;
assign w2844 = ~w2842 & w11915;
assign w2845 = pi1370 & w10;
assign w2846 = w5 & w2845;
assign w2847 = ~w2844 & w2846;
assign w2848 = ~pi0336 & pi0409;
assign w2849 = w2555 & w2848;
assign w2850 = (pi1747 & ~w2555) | (pi1747 & w11917) | (~w2555 & w11917);
assign w2851 = pi1090 & w7;
assign w2852 = ~w14 & ~w2552;
assign w2853 = ~w2557 & ~w2840;
assign w2854 = w2852 & w2853;
assign w2855 = (~w2843 & ~w2854) | (~w2843 & w11918) | (~w2854 & w11918);
assign w2856 = ~w2837 & w2850;
assign w2857 = ~w2855 & w2856;
assign w2858 = ~w2847 & w2857;
assign w2859 = pi0237 & pi1099;
assign w2860 = ~pi0726 & ~pi1099;
assign w2861 = ~w2859 & ~w2860;
assign w2862 = pi1759 & ~pi1760;
assign w2863 = ~pi1763 & ~pi1764;
assign w2864 = ~pi1761 & w2863;
assign w2865 = ~pi1758 & pi1762;
assign w2866 = w2864 & w11919;
assign w2867 = w22 & w11920;
assign w2868 = pi1748 & w2867;
assign w2869 = w2866 & w2868;
assign w2870 = (pi1430 & ~w2868) | (pi1430 & w11921) | (~w2868 & w11921);
assign w2871 = pi1047 & ~pi1526;
assign w2872 = w2870 & w11922;
assign w2873 = ~pi1047 & ~pi1526;
assign w2874 = pi1430 & ~w2873;
assign w2875 = (~w2874 & ~w2868) | (~w2874 & w11923) | (~w2868 & w11923);
assign w2876 = ~pi0311 & w2875;
assign w2877 = w2868 & w11924;
assign w2878 = pi1747 & ~w2877;
assign w2879 = w2870 & w11925;
assign w2880 = ~w2876 & w2878;
assign w2881 = ~w2872 & w2880;
assign w2882 = ~w2879 & w2881;
assign w2883 = w2870 & w11926;
assign w2884 = ~pi0312 & w2875;
assign w2885 = w2868 & w11927;
assign w2886 = pi1747 & ~w2885;
assign w2887 = w2870 & w11928;
assign w2888 = ~w2884 & w2886;
assign w2889 = ~w2883 & w2888;
assign w2890 = ~w2887 & w2889;
assign w2891 = w2870 & w11929;
assign w2892 = ~pi0313 & w2875;
assign w2893 = w2868 & w11930;
assign w2894 = pi1747 & ~w2893;
assign w2895 = w2870 & w11931;
assign w2896 = ~w2892 & w2894;
assign w2897 = ~w2891 & w2896;
assign w2898 = ~w2895 & w2897;
assign w2899 = w2870 & w11932;
assign w2900 = ~pi0314 & w2875;
assign w2901 = w2868 & w11933;
assign w2902 = pi1747 & ~w2901;
assign w2903 = w2870 & w11934;
assign w2904 = ~w2900 & w2902;
assign w2905 = ~w2899 & w2904;
assign w2906 = ~w2903 & w2905;
assign w2907 = w2870 & w11935;
assign w2908 = ~pi0315 & w2875;
assign w2909 = w2868 & w11936;
assign w2910 = pi1747 & ~w2909;
assign w2911 = w2870 & w11937;
assign w2912 = ~w2908 & w2910;
assign w2913 = ~w2907 & w2912;
assign w2914 = ~w2911 & w2913;
assign w2915 = w2870 & w11938;
assign w2916 = ~pi0316 & w2875;
assign w2917 = w2868 & w11939;
assign w2918 = pi1747 & ~w2917;
assign w2919 = w2870 & w11940;
assign w2920 = ~w2916 & w2918;
assign w2921 = ~w2915 & w2920;
assign w2922 = ~w2919 & w2921;
assign w2923 = w2870 & w11941;
assign w2924 = ~pi0317 & w2875;
assign w2925 = w2868 & w11942;
assign w2926 = pi1747 & ~w2925;
assign w2927 = w2870 & w11943;
assign w2928 = ~w2924 & w2926;
assign w2929 = ~w2923 & w2928;
assign w2930 = ~w2927 & w2929;
assign w2931 = pi1758 & pi1762;
assign w2932 = w2864 & w11944;
assign w2933 = w2868 & w11945;
assign w2934 = ~pi0996 & ~pi1729;
assign w2935 = pi1430 & ~w2934;
assign w2936 = (~w2935 & ~w2868) | (~w2935 & w11946) | (~w2868 & w11946);
assign w2937 = ~pi0318 & w2936;
assign w2938 = (w2935 & ~w2868) | (w2935 & w11947) | (~w2868 & w11947);
assign w2939 = pi0011 & w2938;
assign w2940 = pi1747 & ~w2933;
assign w2941 = ~w2937 & w2940;
assign w2942 = ~w2939 & w2941;
assign w2943 = w2870 & w11948;
assign w2944 = ~pi0319 & w2875;
assign w2945 = w2868 & w11949;
assign w2946 = pi1747 & ~w2945;
assign w2947 = w2870 & w11950;
assign w2948 = ~w2944 & w2946;
assign w2949 = ~w2943 & w2948;
assign w2950 = ~w2947 & w2949;
assign w2951 = w2870 & w11951;
assign w2952 = ~pi0320 & w2875;
assign w2953 = w2868 & w11952;
assign w2954 = pi1747 & ~w2953;
assign w2955 = w2870 & w11953;
assign w2956 = ~w2952 & w2954;
assign w2957 = ~w2951 & w2956;
assign w2958 = ~w2955 & w2957;
assign w2959 = w2870 & w11954;
assign w2960 = ~pi0321 & w2875;
assign w2961 = w2868 & w11955;
assign w2962 = pi1747 & ~w2961;
assign w2963 = w2870 & w11956;
assign w2964 = ~w2960 & w2962;
assign w2965 = ~w2959 & w2964;
assign w2966 = ~w2963 & w2965;
assign w2967 = w2868 & w11957;
assign w2968 = ~pi0322 & w2936;
assign w2969 = pi0016 & w2938;
assign w2970 = pi1747 & ~w2967;
assign w2971 = ~w2968 & w2970;
assign w2972 = ~w2969 & w2971;
assign w2973 = w2868 & w11958;
assign w2974 = pi0007 & w2938;
assign w2975 = ~pi0323 & w2936;
assign w2976 = pi1747 & ~w2973;
assign w2977 = ~w2974 & w2976;
assign w2978 = ~w2975 & w2977;
assign w2979 = w2870 & w11959;
assign w2980 = ~pi0324 & w2875;
assign w2981 = w2868 & w11960;
assign w2982 = pi1747 & ~w2981;
assign w2983 = w2870 & w11961;
assign w2984 = ~w2980 & w2982;
assign w2985 = ~w2979 & w2984;
assign w2986 = ~w2983 & w2985;
assign w2987 = w2868 & w11962;
assign w2988 = pi0019 & w2938;
assign w2989 = ~pi0325 & w2936;
assign w2990 = pi1747 & ~w2987;
assign w2991 = ~w2988 & w2990;
assign w2992 = ~w2989 & w2991;
assign w2993 = w2868 & w11963;
assign w2994 = pi0018 & w2938;
assign w2995 = ~pi0326 & w2936;
assign w2996 = pi1747 & ~w2993;
assign w2997 = ~w2994 & w2996;
assign w2998 = ~w2995 & w2997;
assign w2999 = w2868 & w11964;
assign w3000 = pi0023 & w2938;
assign w3001 = ~pi0327 & w2936;
assign w3002 = pi1747 & ~w2999;
assign w3003 = ~w3000 & w3002;
assign w3004 = ~w3001 & w3003;
assign w3005 = w2868 & w11965;
assign w3006 = pi0046 & w2938;
assign w3007 = ~pi0328 & w2936;
assign w3008 = pi1747 & ~w3005;
assign w3009 = ~w3006 & w3008;
assign w3010 = ~w3007 & w3009;
assign w3011 = w2868 & w11966;
assign w3012 = ~pi0329 & w2936;
assign w3013 = pi0028 & w2938;
assign w3014 = pi1747 & ~w3011;
assign w3015 = ~w3012 & w3014;
assign w3016 = ~w3013 & w3015;
assign w3017 = w2868 & w11967;
assign w3018 = ~pi0330 & w2936;
assign w3019 = pi0030 & w2938;
assign w3020 = pi1747 & ~w3017;
assign w3021 = ~w3018 & w3020;
assign w3022 = ~w3019 & w3021;
assign w3023 = ~pi0331 & w2681;
assign w3024 = pi0238 & pi1099;
assign w3025 = ~pi0673 & ~pi1099;
assign w3026 = ~w3024 & ~w3025;
assign w3027 = ~w1529 & w1537;
assign w3028 = w1529 & ~w1537;
assign w3029 = ~w3027 & ~w3028;
assign w3030 = w2868 & w11968;
assign w3031 = ~pi1672 & w2938;
assign w3032 = ~pi0334 & w2936;
assign w3033 = pi1747 & ~w3030;
assign w3034 = ~w3031 & w3033;
assign w3035 = ~w3032 & w3034;
assign w3036 = w2868 & w11969;
assign w3037 = ~pi1666 & w2938;
assign w3038 = ~pi0335 & w2936;
assign w3039 = pi1747 & ~w3036;
assign w3040 = ~w3037 & w3039;
assign w3041 = ~w3038 & w3040;
assign w3042 = w2555 & w11970;
assign w3043 = ~w2553 & ~w3042;
assign w3044 = w1755 & ~w3043;
assign w3045 = w2870 & w11971;
assign w3046 = ~pi0337 & w2875;
assign w3047 = w2868 & w11972;
assign w3048 = pi1747 & ~w3047;
assign w3049 = w2870 & w11973;
assign w3050 = ~w3046 & w3048;
assign w3051 = ~w3045 & w3050;
assign w3052 = ~w3049 & w3051;
assign w3053 = w2870 & w11974;
assign w3054 = ~pi0338 & w2875;
assign w3055 = w2868 & w11975;
assign w3056 = pi1747 & ~w3055;
assign w3057 = w2870 & w11976;
assign w3058 = ~w3054 & w3056;
assign w3059 = ~w3053 & w3058;
assign w3060 = ~w3057 & w3059;
assign w3061 = w2870 & w11977;
assign w3062 = ~pi0339 & w2875;
assign w3063 = w2868 & w11978;
assign w3064 = pi1747 & ~w3063;
assign w3065 = w2870 & w11979;
assign w3066 = ~w3062 & w3064;
assign w3067 = ~w3061 & w3066;
assign w3068 = ~w3065 & w3067;
assign w3069 = w2870 & w11980;
assign w3070 = ~pi0340 & w2875;
assign w3071 = w2868 & w11981;
assign w3072 = pi1747 & ~w3071;
assign w3073 = w2870 & w11982;
assign w3074 = ~w3070 & w3072;
assign w3075 = ~w3069 & w3074;
assign w3076 = ~w3073 & w3075;
assign w3077 = w2870 & w11983;
assign w3078 = ~pi0341 & w2875;
assign w3079 = w2868 & w11984;
assign w3080 = pi1747 & ~w3079;
assign w3081 = w2870 & w11985;
assign w3082 = ~w3078 & w3080;
assign w3083 = ~w3077 & w3082;
assign w3084 = ~w3081 & w3083;
assign w3085 = w2870 & w11986;
assign w3086 = ~pi0342 & w2875;
assign w3087 = w2868 & w11987;
assign w3088 = pi1747 & ~w3087;
assign w3089 = w2870 & w11988;
assign w3090 = ~w3086 & w3088;
assign w3091 = ~w3085 & w3090;
assign w3092 = ~w3089 & w3091;
assign w3093 = w2870 & w11989;
assign w3094 = ~pi0343 & w2875;
assign w3095 = w2868 & w11990;
assign w3096 = pi1747 & ~w3095;
assign w3097 = w2870 & w11991;
assign w3098 = ~w3094 & w3096;
assign w3099 = ~w3093 & w3098;
assign w3100 = ~w3097 & w3099;
assign w3101 = w2870 & w11992;
assign w3102 = ~pi0344 & w2875;
assign w3103 = w2868 & w11993;
assign w3104 = pi1747 & ~w3103;
assign w3105 = w2870 & w11994;
assign w3106 = ~w3102 & w3104;
assign w3107 = ~w3101 & w3106;
assign w3108 = ~w3105 & w3107;
assign w3109 = w2870 & w11995;
assign w3110 = ~pi0345 & w2875;
assign w3111 = w2868 & w11996;
assign w3112 = pi1747 & ~w3111;
assign w3113 = w2870 & w11997;
assign w3114 = ~w3110 & w3112;
assign w3115 = ~w3109 & w3114;
assign w3116 = ~w3113 & w3115;
assign w3117 = w2870 & w11998;
assign w3118 = ~pi0346 & w2875;
assign w3119 = w2868 & w11999;
assign w3120 = pi1747 & ~w3119;
assign w3121 = w2870 & w12000;
assign w3122 = ~w3118 & w3120;
assign w3123 = ~w3117 & w3122;
assign w3124 = ~w3121 & w3123;
assign w3125 = w2870 & w12001;
assign w3126 = ~pi0347 & w2875;
assign w3127 = w2868 & w12002;
assign w3128 = pi1747 & ~w3127;
assign w3129 = w2870 & w12003;
assign w3130 = ~w3126 & w3128;
assign w3131 = ~w3125 & w3130;
assign w3132 = ~w3129 & w3131;
assign w3133 = w2870 & w12004;
assign w3134 = ~pi0348 & w2875;
assign w3135 = w2868 & w12005;
assign w3136 = pi1747 & ~w3135;
assign w3137 = w2870 & w12006;
assign w3138 = ~w3134 & w3136;
assign w3139 = ~w3133 & w3138;
assign w3140 = ~w3137 & w3139;
assign w3141 = w2870 & w12007;
assign w3142 = ~pi0349 & w2875;
assign w3143 = w2868 & w12008;
assign w3144 = pi1747 & ~w3143;
assign w3145 = w2870 & w12009;
assign w3146 = ~w3142 & w3144;
assign w3147 = ~w3141 & w3146;
assign w3148 = ~w3145 & w3147;
assign w3149 = pi1759 & pi1760;
assign w3150 = w2864 & w12010;
assign w3151 = w2868 & w3150;
assign w3152 = (pi1447 & ~w2868) | (pi1447 & w12011) | (~w2868 & w12011);
assign w3153 = w3152 & w11922;
assign w3154 = pi1447 & ~w2873;
assign w3155 = (~w3154 & ~w2868) | (~w3154 & w12012) | (~w2868 & w12012);
assign w3156 = ~pi0350 & w3155;
assign w3157 = w2868 & w12013;
assign w3158 = pi1747 & ~w3157;
assign w3159 = w3152 & w12014;
assign w3160 = ~w3156 & w3158;
assign w3161 = ~w3153 & w3160;
assign w3162 = ~w3159 & w3161;
assign w3163 = w3152 & w11926;
assign w3164 = ~pi0351 & w3155;
assign w3165 = w2868 & w12015;
assign w3166 = pi1747 & ~w3165;
assign w3167 = w3152 & w12016;
assign w3168 = ~w3164 & w3166;
assign w3169 = ~w3163 & w3168;
assign w3170 = ~w3167 & w3169;
assign w3171 = ~w1540 & ~w1543;
assign w3172 = (~w1546 & w1529) | (~w1546 & w12017) | (w1529 & w12017);
assign w3173 = (w3171 & ~w3172) | (w3171 & w12018) | (~w3172 & w12018);
assign w3174 = w3172 & w12019;
assign w3175 = ~w3173 & ~w3174;
assign w3176 = ~w1530 & ~w1544;
assign w3177 = (w1529 & w12021) | (w1529 & w12022) | (w12021 & w12022);
assign w3178 = (w1529 & w12025) | (w1529 & w12026) | (w12025 & w12026);
assign w3179 = w3172 & ~w3178;
assign w3180 = w3152 & w12027;
assign w3181 = ~pi0356 & w3155;
assign w3182 = w2868 & w12028;
assign w3183 = pi1747 & ~w3182;
assign w3184 = w3152 & w12007;
assign w3185 = ~w3181 & w3183;
assign w3186 = ~w3180 & w3185;
assign w3187 = ~w3184 & w3186;
assign w3188 = w2864 & w12029;
assign w3189 = w2868 & w12030;
assign w3190 = pi1447 & ~w2934;
assign w3191 = (w3190 & ~w2868) | (w3190 & w12031) | (~w2868 & w12031);
assign w3192 = pi0023 & w3191;
assign w3193 = (~w3190 & ~w2868) | (~w3190 & w12032) | (~w2868 & w12032);
assign w3194 = ~pi0357 & w3193;
assign w3195 = pi1747 & ~w3189;
assign w3196 = ~w3192 & w3195;
assign w3197 = ~w3194 & w3196;
assign w3198 = pi0586 & ~pi1697;
assign w3199 = pi0662 & w3198;
assign w3200 = w3198 & w12033;
assign w3201 = pi0654 & w3200;
assign w3202 = w3200 & w12034;
assign w3203 = w3200 & w12035;
assign w3204 = pi0569 & w3203;
assign w3205 = w3203 & w12036;
assign w3206 = w3203 & w12037;
assign w3207 = pi0623 & ~pi1139;
assign w3208 = ~pi0623 & pi1139;
assign w3209 = ~w3207 & ~w3208;
assign w3210 = ~pi0566 & pi1034;
assign w3211 = pi0566 & ~pi1034;
assign w3212 = ~w3210 & ~w3211;
assign w3213 = ~pi0569 & pi1265;
assign w3214 = pi0569 & ~pi1265;
assign w3215 = ~w3213 & ~w3214;
assign w3216 = ~pi0648 & pi1142;
assign w3217 = pi0648 & ~pi1142;
assign w3218 = ~w3216 & ~w3217;
assign w3219 = ~pi0650 & pi1033;
assign w3220 = pi0650 & ~pi1033;
assign w3221 = ~w3219 & ~w3220;
assign w3222 = ~pi0654 & pi1258;
assign w3223 = pi0654 & ~pi1258;
assign w3224 = ~w3222 & ~w3223;
assign w3225 = pi0653 & ~pi1141;
assign w3226 = ~pi0653 & pi1141;
assign w3227 = pi0662 & ~pi1342;
assign w3228 = ~pi0662 & pi1342;
assign w3229 = ~pi0586 & pi1032;
assign w3230 = ~w3228 & ~w3229;
assign w3231 = ~w3227 & ~w3230;
assign w3232 = (~w3226 & w3230) | (~w3226 & w12038) | (w3230 & w12038);
assign w3233 = ~w3232 & w12039;
assign w3234 = (w3221 & w3233) | (w3221 & w12040) | (w3233 & w12040);
assign w3235 = (~w3233 & w12041) | (~w3233 & w12042) | (w12041 & w12042);
assign w3236 = w3218 & ~w3235;
assign w3237 = (~w3235 & w12044) | (~w3235 & w12045) | (w12044 & w12045);
assign w3238 = (w3235 & w12046) | (w3235 & w12047) | (w12046 & w12047);
assign w3239 = w3212 & ~w3238;
assign w3240 = (w3238 & w12049) | (w3238 & w12050) | (w12049 & w12050);
assign w3241 = (pi1459 & ~w2873) | (pi1459 & w12051) | (~w2873 & w12051);
assign w3242 = pi1697 & w3241;
assign w3243 = (pi1143 & ~w3241) | (pi1143 & w12052) | (~w3241 & w12052);
assign w3244 = (w3241 & w12053) | (w3241 & w12054) | (w12053 & w12054);
assign w3245 = (w3238 & w12057) | (w3238 & w12058) | (w12057 & w12058);
assign w3246 = w3203 & w12059;
assign w3247 = pi1143 & ~w3246;
assign w3248 = (w3247 & w3245) | (w3247 & w12060) | (w3245 & w12060);
assign w3249 = ~pi0358 & ~w3207;
assign w3250 = (~w3238 & w12061) | (~w3238 & w12062) | (w12061 & w12062);
assign w3251 = w3241 & w5574;
assign w3252 = (~w3238 & w12063) | (~w3238 & w12064) | (w12063 & w12064);
assign w3253 = ~w3248 & ~w3252;
assign w3254 = pi1111 & ~pi1699;
assign w3255 = pi0678 & ~pi1109;
assign w3256 = ~pi0708 & pi1107;
assign w3257 = pi0708 & ~pi1107;
assign w3258 = ~w3256 & ~w3257;
assign w3259 = pi0718 & ~pi1338;
assign w3260 = ~pi0718 & pi1338;
assign w3261 = ~pi0697 & pi1105;
assign w3262 = ~w3260 & ~w3261;
assign w3263 = (~pi1106 & w3262) | (~pi1106 & w12065) | (w3262 & w12065);
assign w3264 = ~w3262 & w12066;
assign w3265 = pi0719 & ~w3264;
assign w3266 = ~w3265 & w12067;
assign w3267 = ~pi1108 & ~w3256;
assign w3268 = (~pi0717 & w3266) | (~pi0717 & w12068) | (w3266 & w12068);
assign w3269 = (~w3256 & w3265) | (~w3256 & w12069) | (w3265 & w12069);
assign w3270 = pi1108 & ~w3257;
assign w3271 = ~w3269 & w3270;
assign w3272 = (~pi1081 & w3269) | (~pi1081 & w12070) | (w3269 & w12070);
assign w3273 = ~w3268 & w3272;
assign w3274 = ~pi0714 & ~w3273;
assign w3275 = ~pi0678 & pi1109;
assign w3276 = ~w3255 & ~w3275;
assign w3277 = ~w3269 & w12071;
assign w3278 = ~pi0717 & pi1081;
assign w3279 = (w3278 & w3266) | (w3278 & w12072) | (w3266 & w12072);
assign w3280 = ~w3277 & ~w3279;
assign w3281 = w3276 & w3280;
assign w3282 = ~w3274 & w3281;
assign w3283 = (~pi1110 & w3282) | (~pi1110 & w12073) | (w3282 & w12073);
assign w3284 = pi1110 & ~w3255;
assign w3285 = ~w3282 & w3284;
assign w3286 = (pi0675 & w3282) | (pi0675 & w12074) | (w3282 & w12074);
assign w3287 = ~w3283 & ~w3286;
assign w3288 = pi1102 & w3287;
assign w3289 = (pi0712 & ~w3287) | (pi0712 & w12075) | (~w3287 & w12075);
assign w3290 = ~pi1102 & ~w3287;
assign w3291 = (pi1480 & ~w2873) | (pi1480 & w12076) | (~w2873 & w12076);
assign w3292 = ~w3290 & w3291;
assign w3293 = (~w3254 & ~w3292) | (~w3254 & w12077) | (~w3292 & w12077);
assign w3294 = pi1111 & pi1699;
assign w3295 = pi0697 & pi0718;
assign w3296 = pi0719 & w3295;
assign w3297 = w3295 & w12078;
assign w3298 = pi0717 & w3297;
assign w3299 = w3297 & w12079;
assign w3300 = pi0675 & pi0678;
assign w3301 = pi0712 & w3300;
assign w3302 = w3299 & w3301;
assign w3303 = (~w3294 & ~w3299) | (~w3294 & w12080) | (~w3299 & w12080);
assign w3304 = ~pi0359 & ~w3303;
assign w3305 = ~w3293 & w3304;
assign w3306 = w3292 & w12081;
assign w3307 = pi0359 & pi1111;
assign w3308 = (w3307 & ~w3302) | (w3307 & w12082) | (~w3302 & w12082);
assign w3309 = ~w3306 & w3308;
assign w3310 = ~w3305 & ~w3309;
assign w3311 = w2868 & w12083;
assign w3312 = pi0049 & w2938;
assign w3313 = ~pi0360 & w2936;
assign w3314 = pi1747 & ~w3311;
assign w3315 = ~w3312 & w3314;
assign w3316 = ~w3313 & w3315;
assign w3317 = ~w1607 & ~w1608;
assign w3318 = w1609 & w3317;
assign w3319 = ~w1609 & ~w3317;
assign w3320 = ~w3318 & ~w3319;
assign w3321 = w3152 & w12084;
assign w3322 = ~pi0362 & w3155;
assign w3323 = w2868 & w12085;
assign w3324 = pi1747 & ~w3323;
assign w3325 = w3152 & w11954;
assign w3326 = ~w3322 & w3324;
assign w3327 = ~w3321 & w3326;
assign w3328 = ~w3325 & w3327;
assign w3329 = w3152 & w12086;
assign w3330 = ~pi0363 & w3155;
assign w3331 = w2868 & w12087;
assign w3332 = pi1747 & ~w3331;
assign w3333 = w3152 & w11935;
assign w3334 = ~w3330 & w3332;
assign w3335 = ~w3329 & w3334;
assign w3336 = ~w3333 & w3335;
assign w3337 = w3152 & w12088;
assign w3338 = ~pi0364 & w3155;
assign w3339 = w2868 & w12089;
assign w3340 = pi1747 & ~w3339;
assign w3341 = w3152 & w11938;
assign w3342 = ~w3338 & w3340;
assign w3343 = ~w3337 & w3342;
assign w3344 = ~w3341 & w3343;
assign w3345 = w3152 & w11941;
assign w3346 = ~pi0365 & w3155;
assign w3347 = w2868 & w12090;
assign w3348 = pi1747 & ~w3347;
assign w3349 = w3152 & w12091;
assign w3350 = ~w3346 & w3348;
assign w3351 = ~w3345 & w3350;
assign w3352 = ~w3349 & w3351;
assign w3353 = w2868 & w12092;
assign w3354 = pi0011 & w3191;
assign w3355 = ~pi0366 & w3193;
assign w3356 = pi1747 & ~w3353;
assign w3357 = ~w3354 & w3356;
assign w3358 = ~w3355 & w3357;
assign w3359 = w3152 & w12093;
assign w3360 = ~pi0367 & w3155;
assign w3361 = w2868 & w12094;
assign w3362 = pi1747 & ~w3361;
assign w3363 = w3152 & w11950;
assign w3364 = ~w3360 & w3362;
assign w3365 = ~w3359 & w3364;
assign w3366 = ~w3363 & w3365;
assign w3367 = w3152 & w12095;
assign w3368 = ~pi0368 & w3155;
assign w3369 = w2868 & w12096;
assign w3370 = pi1747 & ~w3369;
assign w3371 = w3152 & w11951;
assign w3372 = ~w3368 & w3370;
assign w3373 = ~w3367 & w3372;
assign w3374 = ~w3371 & w3373;
assign w3375 = w2868 & w12097;
assign w3376 = pi0016 & w3191;
assign w3377 = ~pi0369 & w3193;
assign w3378 = pi1747 & ~w3375;
assign w3379 = ~w3376 & w3378;
assign w3380 = ~w3377 & w3379;
assign w3381 = w2868 & w12098;
assign w3382 = pi0007 & w3191;
assign w3383 = ~pi0370 & w3193;
assign w3384 = pi1747 & ~w3381;
assign w3385 = ~w3382 & w3384;
assign w3386 = ~w3383 & w3385;
assign w3387 = w3152 & w12099;
assign w3388 = ~pi0371 & w3155;
assign w3389 = w2868 & w12100;
assign w3390 = pi1747 & ~w3389;
assign w3391 = w3152 & w11959;
assign w3392 = ~w3388 & w3390;
assign w3393 = ~w3387 & w3392;
assign w3394 = ~w3391 & w3393;
assign w3395 = w2868 & w12101;
assign w3396 = pi0019 & w3191;
assign w3397 = ~pi0372 & w3193;
assign w3398 = pi1747 & ~w3395;
assign w3399 = ~w3396 & w3398;
assign w3400 = ~w3397 & w3399;
assign w3401 = w2868 & w12102;
assign w3402 = pi0018 & w3191;
assign w3403 = ~pi0373 & w3193;
assign w3404 = pi1747 & ~w3401;
assign w3405 = ~w3402 & w3404;
assign w3406 = ~w3403 & w3405;
assign w3407 = w2868 & w12103;
assign w3408 = pi0046 & w3191;
assign w3409 = ~pi0374 & w3193;
assign w3410 = pi1747 & ~w3407;
assign w3411 = ~w3408 & w3410;
assign w3412 = ~w3409 & w3411;
assign w3413 = w2868 & w12104;
assign w3414 = pi0030 & w3191;
assign w3415 = ~pi0375 & w3193;
assign w3416 = pi1747 & ~w3413;
assign w3417 = ~w3414 & w3416;
assign w3418 = ~w3415 & w3417;
assign w3419 = w2868 & w12105;
assign w3420 = pi0028 & w3191;
assign w3421 = ~pi0376 & w3193;
assign w3422 = pi1747 & ~w3419;
assign w3423 = ~w3420 & w3422;
assign w3424 = ~w3421 & w3423;
assign w3425 = w2868 & w12106;
assign w3426 = ~pi0377 & w2936;
assign w3427 = pi0194 & w2938;
assign w3428 = pi1747 & ~w3425;
assign w3429 = ~w3426 & w3428;
assign w3430 = ~w3427 & w3429;
assign w3431 = w2868 & w12107;
assign w3432 = pi0286 & w2938;
assign w3433 = ~pi0378 & w2936;
assign w3434 = pi1747 & ~w3431;
assign w3435 = ~w3432 & w3434;
assign w3436 = ~w3433 & w3435;
assign w3437 = ~pi0387 & pi1270;
assign w3438 = ~pi0480 & pi1274;
assign w3439 = pi0480 & ~pi1274;
assign w3440 = ~w3438 & ~w3439;
assign w3441 = ~pi0484 & pi1121;
assign w3442 = pi0484 & ~pi1121;
assign w3443 = ~w3441 & ~w3442;
assign w3444 = ~pi0508 & pi1023;
assign w3445 = pi0508 & ~pi1023;
assign w3446 = ~w3444 & ~w3445;
assign w3447 = pi0507 & ~pi1277;
assign w3448 = ~pi0507 & pi1277;
assign w3449 = ~pi0408 & pi1022;
assign w3450 = ~w3448 & ~w3449;
assign w3451 = ~w3447 & ~w3450;
assign w3452 = w3446 & w3451;
assign w3453 = (~w3444 & ~w3451) | (~w3444 & w12108) | (~w3451 & w12108);
assign w3454 = pi1272 & ~w3453;
assign w3455 = ~pi1272 & w3453;
assign w3456 = (~pi0509 & ~w3453) | (~pi0509 & w12109) | (~w3453 & w12109);
assign w3457 = ~w3454 & ~w3456;
assign w3458 = w3443 & ~w3457;
assign w3459 = (~w3457 & w12111) | (~w3457 & w12112) | (w12111 & w12112);
assign w3460 = (w3457 & w12115) | (w3457 & w12116) | (w12115 & w12116);
assign w3461 = pi0387 & ~pi1270;
assign w3462 = pi1267 & ~w3461;
assign w3463 = ~w3460 & w12117;
assign w3464 = (~w3457 & w12118) | (~w3457 & w12119) | (w12118 & w12119);
assign w3465 = ~pi1267 & ~w3437;
assign w3466 = ~w3464 & w3465;
assign w3467 = ~pi0386 & pi1119;
assign w3468 = (w3467 & w3464) | (w3467 & w12120) | (w3464 & w12120);
assign w3469 = ~w3463 & ~w3468;
assign w3470 = pi0466 & w3469;
assign w3471 = (pi1430 & ~w2873) | (pi1430 & w12121) | (~w2873 & w12121);
assign w3472 = pi1690 & w3471;
assign w3473 = (~pi0386 & w3464) | (~pi0386 & w12122) | (w3464 & w12122);
assign w3474 = (~pi1119 & w3460) | (~pi1119 & w12123) | (w3460 & w12123);
assign w3475 = ~w3473 & w3474;
assign w3476 = w3472 & ~w3475;
assign w3477 = ~w3470 & w3476;
assign w3478 = pi0480 & pi0484;
assign w3479 = pi0387 & w3478;
assign w3480 = pi0408 & pi0507;
assign w3481 = pi0508 & w3480;
assign w3482 = w3480 & w12124;
assign w3483 = w3478 & w12125;
assign w3484 = w3482 & w3483;
assign w3485 = w3484 & w12126;
assign w3486 = pi0379 & pi1122;
assign w3487 = ~w3477 & w12127;
assign w3488 = ~pi0379 & pi1122;
assign w3489 = (w3488 & w3477) | (w3488 & w12128) | (w3477 & w12128);
assign w3490 = ~w3487 & ~w3489;
assign w3491 = pi1131 & pi1679;
assign w3492 = pi1131 & ~pi1679;
assign w3493 = pi0485 & pi0549;
assign w3494 = pi0506 & pi0618;
assign w3495 = pi0587 & w3494;
assign w3496 = pi0567 & pi0622;
assign w3497 = w3495 & w3496;
assign w3498 = pi0483 & w3493;
assign w3499 = w3497 & w12129;
assign w3500 = pi0380 & w3499;
assign w3501 = (w3492 & w3499) | (w3492 & w12130) | (w3499 & w12130);
assign w3502 = ~w3500 & w3501;
assign w3503 = ~w3491 & ~w3502;
assign w3504 = pi0533 & ~pi1127;
assign w3505 = ~pi0485 & pi1076;
assign w3506 = pi0567 & ~pi1083;
assign w3507 = ~pi0567 & pi1083;
assign w3508 = ~w3506 & ~w3507;
assign w3509 = pi0618 & ~pi1310;
assign w3510 = ~pi0618 & pi1310;
assign w3511 = ~pi0506 & pi1027;
assign w3512 = ~w3510 & ~w3511;
assign w3513 = (~pi1129 & w3512) | (~pi1129 & w12131) | (w3512 & w12131);
assign w3514 = ~w3512 & w12132;
assign w3515 = pi0587 & ~w3514;
assign w3516 = (~pi1028 & w3515) | (~pi1028 & w12133) | (w3515 & w12133);
assign w3517 = ~w3515 & w12134;
assign w3518 = pi0622 & ~w3517;
assign w3519 = (w3508 & w3518) | (w3508 & w12135) | (w3518 & w12135);
assign w3520 = (~pi1130 & w3519) | (~pi1130 & w12136) | (w3519 & w12136);
assign w3521 = pi1130 & ~w3506;
assign w3522 = ~w3519 & w3521;
assign w3523 = (pi0549 & w3519) | (pi0549 & w12137) | (w3519 & w12137);
assign w3524 = ~w3520 & ~w3523;
assign w3525 = ~pi0483 & pi1029;
assign w3526 = pi0483 & ~pi1029;
assign w3527 = ~w3525 & ~w3526;
assign w3528 = pi0485 & ~pi1076;
assign w3529 = w3527 & ~w3528;
assign w3530 = (w3529 & w3524) | (w3529 & w12138) | (w3524 & w12138);
assign w3531 = pi0533 & ~w3525;
assign w3532 = (w3524 & w12141) | (w3524 & w12142) | (w12141 & w12142);
assign w3533 = ~pi1127 & ~w3525;
assign w3534 = (~w3524 & w12143) | (~w3524 & w12144) | (w12143 & w12144);
assign w3535 = (pi1447 & ~w2873) | (pi1447 & w12145) | (~w2873 & w12145);
assign w3536 = ~w3534 & w3535;
assign w3537 = (pi0380 & ~w3536) | (pi0380 & w12146) | (~w3536 & w12146);
assign w3538 = ~pi0380 & w3535;
assign w3539 = (w3524 & w12147) | (w3524 & w12148) | (w12147 & w12148);
assign w3540 = w3532 & w3539;
assign w3541 = ~w3502 & ~w3540;
assign w3542 = ~w3537 & w3541;
assign w3543 = ~w3503 & ~w3542;
assign w3544 = w3484 & w12149;
assign w3545 = (pi0470 & ~w3484) | (pi0470 & w12150) | (~w3484 & w12150);
assign w3546 = pi1122 & w3545;
assign w3547 = w3545 & w12151;
assign w3548 = w3471 & w12152;
assign w3549 = ~w3475 & w3548;
assign w3550 = ~w3470 & w3549;
assign w3551 = ~pi0470 & pi1122;
assign w3552 = pi0381 & w3551;
assign w3553 = ~w3550 & w3552;
assign w3554 = ~pi0381 & pi1122;
assign w3555 = ~w3545 & w3554;
assign w3556 = (w3555 & w3550) | (w3555 & w12153) | (w3550 & w12153);
assign w3557 = ~w3547 & ~w3553;
assign w3558 = ~w3556 & w3557;
assign w3559 = ~pi1626 & pi1628;
assign w3560 = ~pi1627 & w3559;
assign w3561 = ~w355 & ~w1209;
assign w3562 = ~pi0382 & ~pi0647;
assign w3563 = ~pi0695 & pi0696;
assign w3564 = w3562 & w3563;
assign w3565 = ~w3561 & w12154;
assign w3566 = pi0382 & ~pi0647;
assign w3567 = w1229 & w3566;
assign w3568 = ~w3565 & ~w3567;
assign w3569 = ~pi0696 & w3562;
assign w3570 = pi0695 & ~w3559;
assign w3571 = w3569 & w3570;
assign w3572 = ~w1231 & ~w3564;
assign w3573 = (pi1626 & ~w3572) | (pi1626 & w12155) | (~w3572 & w12155);
assign w3574 = w3560 & w3567;
assign w3575 = pi1747 & ~w3571;
assign w3576 = ~w3574 & w3575;
assign w3577 = ~w3573 & w3576;
assign w3578 = ~w3568 & w3577;
assign w3579 = pi0413 & pi1272;
assign w3580 = ~pi0413 & ~pi1272;
assign w3581 = ~w3579 & ~w3580;
assign w3582 = ~pi0411 & ~pi1277;
assign w3583 = pi0411 & pi1277;
assign w3584 = pi0410 & pi1022;
assign w3585 = ~w3583 & ~w3584;
assign w3586 = (~pi1023 & w3585) | (~pi1023 & w12156) | (w3585 & w12156);
assign w3587 = ~w3585 & w12157;
assign w3588 = ~pi0412 & ~w3587;
assign w3589 = ~w3588 & w12158;
assign w3590 = ~pi1121 & ~w3579;
assign w3591 = ~w3589 & w3590;
assign w3592 = (pi0442 & w3589) | (pi0442 & w12159) | (w3589 & w12159);
assign w3593 = (~w3579 & w3588) | (~w3579 & w12160) | (w3588 & w12160);
assign w3594 = pi1121 & ~w3580;
assign w3595 = ~w3593 & w3594;
assign w3596 = (~pi1274 & w3593) | (~pi1274 & w12161) | (w3593 & w12161);
assign w3597 = ~w3592 & w3596;
assign w3598 = pi0510 & ~w3597;
assign w3599 = ~w3593 & w12162;
assign w3600 = pi0442 & pi1274;
assign w3601 = (w3600 & w3589) | (w3600 & w12163) | (w3589 & w12163);
assign w3602 = ~w3599 & ~w3601;
assign w3603 = ~pi1270 & w3602;
assign w3604 = ~w3598 & w3603;
assign w3605 = pi0388 & ~w3604;
assign w3606 = ~pi0510 & w3602;
assign w3607 = pi1270 & ~w3597;
assign w3608 = ~w3606 & w3607;
assign w3609 = ~pi1267 & ~w3608;
assign w3610 = ~w3605 & w3609;
assign w3611 = pi0482 & ~w3610;
assign w3612 = ~pi0388 & ~w3608;
assign w3613 = pi1267 & ~w3604;
assign w3614 = ~w3612 & w3613;
assign w3615 = ~pi1119 & ~w3614;
assign w3616 = ~w3611 & w3615;
assign w3617 = w3471 & ~w3616;
assign w3618 = pi0482 & pi1119;
assign w3619 = ~w3610 & w3618;
assign w3620 = pi1119 & pi1267;
assign w3621 = ~w3604 & w3620;
assign w3622 = ~w3612 & w3621;
assign w3623 = ~pi0441 & ~w3622;
assign w3624 = ~w3619 & w3623;
assign w3625 = ~pi0410 & ~pi0411;
assign w3626 = ~pi0412 & ~pi0413;
assign w3627 = ~pi0442 & ~pi0510;
assign w3628 = w3626 & w3627;
assign w3629 = ~pi0388 & ~pi0482;
assign w3630 = w3628 & w3629;
assign w3631 = w3628 & w12164;
assign w3632 = (w3631 & w12166) | (w3631 & w12167) | (w12166 & w12167);
assign w3633 = ~w3624 & w3632;
assign w3634 = w3617 & w3633;
assign w3635 = w3631 & w12168;
assign w3636 = w3631 & w12169;
assign w3637 = pi0481 & pi1690;
assign w3638 = ~pi0481 & ~pi1690;
assign w3639 = ~w3637 & ~w3638;
assign w3640 = pi0383 & ~w3639;
assign w3641 = (w3640 & w3634) | (w3640 & w12170) | (w3634 & w12170);
assign w3642 = (w3631 & w12171) | (w3631 & w12172) | (w12171 & w12172);
assign w3643 = ~w3624 & w3642;
assign w3644 = w3617 & w3643;
assign w3645 = ~pi0384 & ~pi0481;
assign w3646 = (~pi0383 & ~w3631) | (~pi0383 & w12174) | (~w3631 & w12174);
assign w3647 = (pi1122 & w3644) | (pi1122 & w12175) | (w3644 & w12175);
assign w3648 = ~w3641 & w3647;
assign w3649 = w3472 & ~w3616;
assign w3650 = (~w3635 & ~w3649) | (~w3635 & w12176) | (~w3649 & w12176);
assign w3651 = pi0384 & pi1122;
assign w3652 = w3650 & w3651;
assign w3653 = ~pi0384 & pi1122;
assign w3654 = ~w3650 & w3653;
assign w3655 = ~w3652 & ~w3654;
assign w3656 = pi0385 & w1860;
assign w3657 = w1829 & w12177;
assign w3658 = pi0897 & w1813;
assign w3659 = pi0898 & w1865;
assign w3660 = pi0896 & w1867;
assign w3661 = ~w3658 & ~w3660;
assign w3662 = ~w3657 & w3661;
assign w3663 = ~w3656 & w3662;
assign w3664 = ~w3659 & w3663;
assign w3665 = ~pi1690 & w3482;
assign w3666 = w3479 & w3665;
assign w3667 = (w3472 & w3460) | (w3472 & w12178) | (w3460 & w12178);
assign w3668 = ~w3466 & w3667;
assign w3669 = (pi0386 & w3668) | (pi0386 & w12179) | (w3668 & w12179);
assign w3670 = ~w3668 & w12180;
assign w3671 = pi1122 & ~w3669;
assign w3672 = ~w3670 & w3671;
assign w3673 = ~w3437 & ~w3461;
assign w3674 = (~w3457 & w12181) | (~w3457 & w12182) | (w12181 & w12182);
assign w3675 = pi1122 & pi1690;
assign w3676 = w3471 & w3675;
assign w3677 = (w3457 & w12183) | (w3457 & w12184) | (w12183 & w12184);
assign w3678 = ~w3674 & w3676;
assign w3679 = ~w3677 & w3678;
assign w3680 = (pi1122 & ~w3471) | (pi1122 & w3681) | (~w3471 & w3681);
assign w3681 = pi1122 & ~pi1690;
assign w3682 = w3482 & w12185;
assign w3683 = ~pi0387 & ~w3682;
assign w3684 = ~w3666 & w3680;
assign w3685 = ~w3683 & w3684;
assign w3686 = ~w3679 & ~w3685;
assign w3687 = ~pi0410 & ~pi1690;
assign w3688 = ~pi0411 & w3687;
assign w3689 = w3628 & w3688;
assign w3690 = ~w3604 & ~w3608;
assign w3691 = w3676 & w3690;
assign w3692 = (~pi0388 & ~w3689) | (~pi0388 & w12186) | (~w3689 & w12186);
assign w3693 = ~w3691 & w3692;
assign w3694 = w3680 & ~w3689;
assign w3695 = pi0388 & ~w3694;
assign w3696 = (w3695 & w3690) | (w3695 & w12187) | (w3690 & w12187);
assign w3697 = ~w3693 & ~w3696;
assign w3698 = w2868 & w12188;
assign w3699 = pi0064 & w2938;
assign w3700 = ~pi0389 & w2936;
assign w3701 = pi1747 & ~w3698;
assign w3702 = ~w3699 & w3701;
assign w3703 = ~w3700 & w3702;
assign w3704 = w2868 & w12189;
assign w3705 = pi0014 & w2938;
assign w3706 = ~pi0390 & w2936;
assign w3707 = pi1747 & ~w3704;
assign w3708 = ~w3705 & w3707;
assign w3709 = ~w3706 & w3708;
assign w3710 = w2868 & w12190;
assign w3711 = pi0015 & w2938;
assign w3712 = ~pi0391 & w2936;
assign w3713 = pi1747 & ~w3710;
assign w3714 = ~w3711 & w3713;
assign w3715 = ~w3712 & w3714;
assign w3716 = w2868 & w12191;
assign w3717 = pi0953 & w2938;
assign w3718 = ~pi0392 & w2936;
assign w3719 = pi1747 & ~w3716;
assign w3720 = ~w3717 & w3719;
assign w3721 = ~w3718 & w3720;
assign w3722 = w2868 & w12192;
assign w3723 = pi0332 & w2938;
assign w3724 = ~pi0393 & w2936;
assign w3725 = pi1747 & ~w3722;
assign w3726 = ~w3723 & w3725;
assign w3727 = ~w3724 & w3726;
assign w3728 = w2868 & w12193;
assign w3729 = pi0057 & w2938;
assign w3730 = ~pi0394 & w2936;
assign w3731 = pi1747 & ~w3728;
assign w3732 = ~w3729 & w3731;
assign w3733 = ~w3730 & w3732;
assign w3734 = w2868 & w12194;
assign w3735 = pi0299 & w2938;
assign w3736 = ~pi0395 & w2936;
assign w3737 = pi1747 & ~w3734;
assign w3738 = ~w3735 & w3737;
assign w3739 = ~w3736 & w3738;
assign w3740 = w2868 & w12195;
assign w3741 = ~pi0396 & w2936;
assign w3742 = pi1481 & w2938;
assign w3743 = pi1747 & ~w3740;
assign w3744 = ~w3741 & w3743;
assign w3745 = ~w3742 & w3744;
assign w3746 = w2868 & w12196;
assign w3747 = pi0223 & w2938;
assign w3748 = ~pi0397 & w2936;
assign w3749 = pi1747 & ~w3746;
assign w3750 = ~w3747 & w3749;
assign w3751 = ~w3748 & w3750;
assign w3752 = w2868 & w12197;
assign w3753 = ~pi0398 & w2936;
assign w3754 = pi0154 & w2938;
assign w3755 = pi1747 & ~w3752;
assign w3756 = ~w3753 & w3755;
assign w3757 = ~w3754 & w3756;
assign w3758 = w2868 & w12198;
assign w3759 = ~pi0399 & w2936;
assign w3760 = pi0254 & w2938;
assign w3761 = pi1747 & ~w3758;
assign w3762 = ~w3759 & w3761;
assign w3763 = ~w3760 & w3762;
assign w3764 = w2868 & w12199;
assign w3765 = ~pi0400 & w2936;
assign w3766 = pi0124 & w2938;
assign w3767 = pi1747 & ~w3764;
assign w3768 = ~w3765 & w3767;
assign w3769 = ~w3766 & w3768;
assign w3770 = w2868 & w12200;
assign w3771 = pi0155 & w2938;
assign w3772 = ~pi0401 & w2936;
assign w3773 = pi1747 & ~w3770;
assign w3774 = ~w3771 & w3773;
assign w3775 = ~w3772 & w3774;
assign w3776 = w2868 & w12201;
assign w3777 = pi0056 & w2938;
assign w3778 = ~pi0402 & w2936;
assign w3779 = pi1747 & ~w3776;
assign w3780 = ~w3777 & w3779;
assign w3781 = ~w3778 & w3780;
assign w3782 = w2868 & w12202;
assign w3783 = ~pi0403 & w2936;
assign w3784 = pi0063 & w2938;
assign w3785 = pi1747 & ~w3782;
assign w3786 = ~w3783 & w3785;
assign w3787 = ~w3784 & w3786;
assign w3788 = w2868 & w12203;
assign w3789 = pi0027 & w2938;
assign w3790 = ~pi0404 & w2936;
assign w3791 = pi1747 & ~w3788;
assign w3792 = ~w3789 & w3791;
assign w3793 = ~w3790 & w3792;
assign w3794 = w2868 & w12204;
assign w3795 = ~pi0405 & w2936;
assign w3796 = pi0022 & w2938;
assign w3797 = pi1747 & ~w3794;
assign w3798 = ~w3795 & w3797;
assign w3799 = ~w3796 & w3798;
assign w3800 = w2868 & w12205;
assign w3801 = ~pi1672 & w3191;
assign w3802 = ~pi0406 & w3193;
assign w3803 = pi1747 & ~w3800;
assign w3804 = ~w3801 & w3803;
assign w3805 = ~w3802 & w3804;
assign w3806 = w2868 & w12206;
assign w3807 = ~pi1666 & w3191;
assign w3808 = ~pi0407 & w3193;
assign w3809 = pi1747 & ~w3806;
assign w3810 = ~w3807 & w3809;
assign w3811 = ~w3808 & w3810;
assign w3812 = (pi1690 & ~w3471) | (pi1690 & w12207) | (~w3471 & w12207);
assign w3813 = (~w3471 & w12208) | (~w3471 & w12209) | (w12208 & w12209);
assign w3814 = (pi1122 & w3812) | (pi1122 & w12210) | (w3812 & w12210);
assign w3815 = ~w3813 & w3814;
assign w3816 = w2849 & w2850;
assign w3817 = pi0258 & w1755;
assign w3818 = w2555 & w12211;
assign w3819 = ~w3816 & ~w3818;
assign w3820 = (w3471 & w12212) | (w3471 & w12213) | (w12212 & w12213);
assign w3821 = (~w3471 & w12214) | (~w3471 & w12215) | (w12214 & w12215);
assign w3822 = pi1122 & ~w3820;
assign w3823 = ~w3821 & w3822;
assign w3824 = pi0411 & ~w3687;
assign w3825 = ~w3688 & ~w3824;
assign w3826 = w3680 & ~w3825;
assign w3827 = ~w3582 & ~w3583;
assign w3828 = ~w3584 & ~w3827;
assign w3829 = w3584 & w3827;
assign w3830 = ~w3828 & ~w3829;
assign w3831 = w3676 & w3830;
assign w3832 = ~w3826 & ~w3831;
assign w3833 = ~w3586 & ~w3587;
assign w3834 = (~w3688 & ~w3833) | (~w3688 & w12216) | (~w3833 & w12216);
assign w3835 = ~pi0412 & w3834;
assign w3836 = (pi1122 & w3834) | (pi1122 & w12217) | (w3834 & w12217);
assign w3837 = ~w3835 & w3836;
assign w3838 = ~pi0412 & w3625;
assign w3839 = (pi0413 & ~w3838) | (pi0413 & w12218) | (~w3838 & w12218);
assign w3840 = w3680 & w3839;
assign w3841 = w3626 & w3688;
assign w3842 = w3688 & w12219;
assign w3843 = (~w3581 & w3588) | (~w3581 & w12220) | (w3588 & w12220);
assign w3844 = ~w3589 & w3676;
assign w3845 = ~w3843 & w3844;
assign w3846 = ~w3840 & ~w3842;
assign w3847 = ~w3845 & w3846;
assign w3848 = w3152 & w12221;
assign w3849 = ~pi0414 & w3155;
assign w3850 = w2868 & w12222;
assign w3851 = pi1747 & ~w3850;
assign w3852 = w3152 & w12223;
assign w3853 = ~w3849 & w3851;
assign w3854 = ~w3848 & w3853;
assign w3855 = ~w3852 & w3854;
assign w3856 = w3152 & w11974;
assign w3857 = ~pi0415 & w3155;
assign w3858 = w2868 & w12224;
assign w3859 = pi1747 & ~w3858;
assign w3860 = w3152 & w12225;
assign w3861 = ~w3857 & w3859;
assign w3862 = ~w3856 & w3861;
assign w3863 = ~w3860 & w3862;
assign w3864 = w3152 & w12226;
assign w3865 = ~pi0416 & w3155;
assign w3866 = w2868 & w12227;
assign w3867 = pi1747 & ~w3866;
assign w3868 = w3152 & w11977;
assign w3869 = ~w3865 & w3867;
assign w3870 = ~w3864 & w3869;
assign w3871 = ~w3868 & w3870;
assign w3872 = w3152 & w12228;
assign w3873 = ~pi0417 & w3155;
assign w3874 = w2868 & w12229;
assign w3875 = pi1747 & ~w3874;
assign w3876 = w3152 & w11980;
assign w3877 = ~w3873 & w3875;
assign w3878 = ~w3872 & w3877;
assign w3879 = ~w3876 & w3878;
assign w3880 = w3152 & w11983;
assign w3881 = ~pi0418 & w3155;
assign w3882 = w2868 & w12230;
assign w3883 = pi1747 & ~w3882;
assign w3884 = w3152 & w12231;
assign w3885 = ~w3881 & w3883;
assign w3886 = ~w3880 & w3885;
assign w3887 = ~w3884 & w3886;
assign w3888 = w3152 & w11986;
assign w3889 = ~pi0419 & w3155;
assign w3890 = w2868 & w12232;
assign w3891 = pi1747 & ~w3890;
assign w3892 = w3152 & w12233;
assign w3893 = ~w3889 & w3891;
assign w3894 = ~w3888 & w3893;
assign w3895 = ~w3892 & w3894;
assign w3896 = w3152 & w12234;
assign w3897 = ~pi0420 & w3155;
assign w3898 = w2868 & w12235;
assign w3899 = pi1747 & ~w3898;
assign w3900 = w3152 & w11989;
assign w3901 = ~w3897 & w3899;
assign w3902 = ~w3896 & w3901;
assign w3903 = ~w3900 & w3902;
assign w3904 = w3152 & w12236;
assign w3905 = ~pi0421 & w3155;
assign w3906 = w2868 & w12237;
assign w3907 = pi1747 & ~w3906;
assign w3908 = w3152 & w11994;
assign w3909 = ~w3905 & w3907;
assign w3910 = ~w3904 & w3909;
assign w3911 = ~w3908 & w3910;
assign w3912 = w3152 & w11995;
assign w3913 = ~pi0422 & w3155;
assign w3914 = w2868 & w12238;
assign w3915 = pi1747 & ~w3914;
assign w3916 = w3152 & w12239;
assign w3917 = ~w3913 & w3915;
assign w3918 = ~w3912 & w3917;
assign w3919 = ~w3916 & w3918;
assign w3920 = w3152 & w12240;
assign w3921 = ~pi0423 & w3155;
assign w3922 = w2868 & w12241;
assign w3923 = pi1747 & ~w3922;
assign w3924 = w3152 & w11932;
assign w3925 = ~w3921 & w3923;
assign w3926 = ~w3920 & w3925;
assign w3927 = ~w3924 & w3926;
assign w3928 = w3152 & w12242;
assign w3929 = ~pi0424 & w3155;
assign w3930 = w2868 & w12243;
assign w3931 = pi1747 & ~w3930;
assign w3932 = w3152 & w12001;
assign w3933 = ~w3929 & w3931;
assign w3934 = ~w3928 & w3933;
assign w3935 = ~w3932 & w3934;
assign w3936 = w3152 & w12244;
assign w3937 = ~pi0425 & w3155;
assign w3938 = w2868 & w12245;
assign w3939 = pi1747 & ~w3938;
assign w3940 = w3152 & w12006;
assign w3941 = ~w3937 & w3939;
assign w3942 = ~w3936 & w3941;
assign w3943 = ~w3940 & w3942;
assign w3944 = w3152 & w12246;
assign w3945 = ~pi0426 & w3155;
assign w3946 = w2868 & w12247;
assign w3947 = pi1747 & ~w3946;
assign w3948 = w3152 & w11931;
assign w3949 = ~w3945 & w3947;
assign w3950 = ~w3944 & w3949;
assign w3951 = ~w3948 & w3950;
assign w3952 = pi1761 & w2863;
assign w3953 = w3952 & w11919;
assign w3954 = w2868 & w3953;
assign w3955 = (pi1459 & ~w2868) | (pi1459 & w12248) | (~w2868 & w12248);
assign w3956 = w3955 & w11922;
assign w3957 = pi1459 & ~w2873;
assign w3958 = (~w3957 & ~w2868) | (~w3957 & w12249) | (~w2868 & w12249);
assign w3959 = ~pi0427 & w3958;
assign w3960 = w2868 & w12250;
assign w3961 = pi1747 & ~w3960;
assign w3962 = w3955 & w12251;
assign w3963 = ~w3959 & w3961;
assign w3964 = ~w3956 & w3963;
assign w3965 = ~w3962 & w3964;
assign w3966 = w3955 & w12252;
assign w3967 = ~pi0428 & w3958;
assign w3968 = w2868 & w12253;
assign w3969 = pi1747 & ~w3968;
assign w3970 = w3955 & w11926;
assign w3971 = ~w3967 & w3969;
assign w3972 = ~w3966 & w3971;
assign w3973 = ~w3970 & w3972;
assign w3974 = ~pi0269 & pi1039;
assign w3975 = w357 & w1174;
assign w3976 = pi0251 & ~pi1042;
assign w3977 = ~pi0271 & pi1040;
assign w3978 = pi0253 & ~pi1313;
assign w3979 = pi0273 & ~pi1017;
assign w3980 = ~pi0252 & pi1044;
assign w3981 = pi0271 & ~pi1040;
assign w3982 = ~pi0270 & pi1041;
assign w3983 = pi0250 & ~pi1318;
assign w3984 = ~pi0263 & pi1043;
assign w3985 = ~pi0250 & pi1318;
assign w3986 = pi0263 & ~pi1043;
assign w3987 = ~pi0253 & pi1313;
assign w3988 = pi0272 & ~pi1049;
assign w3989 = pi0270 & ~pi1041;
assign w3990 = ~pi0251 & pi1042;
assign w3991 = pi0269 & ~pi1039;
assign w3992 = pi0255 & ~pi1317;
assign w3993 = ~pi0272 & pi1049;
assign w3994 = pi0252 & ~pi1044;
assign w3995 = ~pi0255 & pi1317;
assign w3996 = ~pi0273 & pi1017;
assign w3997 = ~w3974 & ~w3976;
assign w3998 = ~w3977 & ~w3978;
assign w3999 = ~w3979 & ~w3980;
assign w4000 = ~w3981 & ~w3982;
assign w4001 = ~w3983 & ~w3984;
assign w4002 = ~w3985 & ~w3986;
assign w4003 = ~w3987 & ~w3988;
assign w4004 = ~w3989 & ~w3990;
assign w4005 = ~w3991 & ~w3992;
assign w4006 = ~w3993 & ~w3994;
assign w4007 = ~w3995 & ~w3996;
assign w4008 = w4006 & w4007;
assign w4009 = w4004 & w4005;
assign w4010 = w4002 & w4003;
assign w4011 = w4000 & w4001;
assign w4012 = w3998 & w3999;
assign w4013 = w3997 & w4012;
assign w4014 = w4010 & w4011;
assign w4015 = w4008 & w4009;
assign w4016 = w4014 & w4015;
assign w4017 = w4013 & w4016;
assign w4018 = w3975 & w4017;
assign w4019 = w2868 & w12254;
assign w4020 = ~pi0430 & w2936;
assign w4021 = pi0310 & w2938;
assign w4022 = pi1747 & ~w4019;
assign w4023 = ~w4020 & w4022;
assign w4024 = ~w4021 & w4023;
assign w4025 = (~w1529 & w12255) | (~w1529 & w12256) | (w12255 & w12256);
assign w4026 = ~w3177 & ~w4025;
assign w4027 = w3152 & w11998;
assign w4028 = ~pi0432 & w3155;
assign w4029 = w2868 & w12257;
assign w4030 = pi1747 & ~w4029;
assign w4031 = w3152 & w12258;
assign w4032 = ~w4028 & w4030;
assign w4033 = ~w4027 & w4032;
assign w4034 = ~w4031 & w4033;
assign w4035 = pi0469 & pi1671;
assign w4036 = (~pi0433 & ~w4035) | (~pi0433 & w12259) | (~w4035 & w12259);
assign w4037 = w4035 & w12260;
assign w4038 = ~pi0705 & ~w4036;
assign w4039 = ~w4037 & w4038;
assign w4040 = w2870 & w12261;
assign w4041 = ~pi0435 & w2875;
assign w4042 = w2868 & w12262;
assign w4043 = pi1747 & ~w4042;
assign w4044 = w2870 & w12263;
assign w4045 = ~w4041 & w4043;
assign w4046 = ~w4040 & w4045;
assign w4047 = ~w4044 & w4046;
assign w4048 = w3955 & w12007;
assign w4049 = ~pi0436 & w3958;
assign w4050 = w2868 & w12264;
assign w4051 = pi1747 & ~w4050;
assign w4052 = w3955 & w12265;
assign w4053 = ~w4049 & w4051;
assign w4054 = ~w4048 & w4053;
assign w4055 = ~w4052 & w4054;
assign w4056 = w3952 & w12010;
assign w4057 = w2868 & w4056;
assign w4058 = (pi1480 & ~w2868) | (pi1480 & w12266) | (~w2868 & w12266);
assign w4059 = w4058 & w11926;
assign w4060 = pi1480 & ~w2873;
assign w4061 = (~w4060 & ~w2868) | (~w4060 & w12267) | (~w2868 & w12267);
assign w4062 = ~pi0437 & w4061;
assign w4063 = w2868 & w12268;
assign w4064 = pi1747 & ~w4063;
assign w4065 = w4058 & w12269;
assign w4066 = ~w4062 & w4064;
assign w4067 = ~w4059 & w4066;
assign w4068 = ~w4065 & w4067;
assign w4069 = w2870 & w12270;
assign w4070 = ~pi0438 & w2875;
assign w4071 = w2868 & w12271;
assign w4072 = pi1747 & ~w4071;
assign w4073 = w2870 & w12272;
assign w4074 = ~w4070 & w4072;
assign w4075 = ~w4069 & w4074;
assign w4076 = ~w4073 & w4075;
assign w4077 = w3955 & w12273;
assign w4078 = ~pi0439 & w3958;
assign w4079 = w2868 & w12274;
assign w4080 = pi1747 & ~w4079;
assign w4081 = w3955 & w12275;
assign w4082 = ~w4078 & w4080;
assign w4083 = ~w4077 & w4082;
assign w4084 = ~w4081 & w4083;
assign w4085 = w2868 & w12276;
assign w4086 = pi0057 & w3191;
assign w4087 = ~pi0440 & w3193;
assign w4088 = pi1747 & ~w4085;
assign w4089 = ~w4086 & w4088;
assign w4090 = ~w4087 & w4089;
assign w4091 = ~w3619 & ~w3622;
assign w4092 = (pi0441 & ~w3617) | (pi0441 & w12277) | (~w3617 & w12277);
assign w4093 = (pi1690 & ~w3617) | (pi1690 & w12278) | (~w3617 & w12278);
assign w4094 = ~w4092 & w4093;
assign w4095 = pi0441 & ~w3631;
assign w4096 = (~pi1690 & ~w3631) | (~pi1690 & w12279) | (~w3631 & w12279);
assign w4097 = ~w4095 & w4096;
assign w4098 = pi1122 & ~w4097;
assign w4099 = ~w4094 & w4098;
assign w4100 = w3680 & ~w3841;
assign w4101 = ~w3591 & ~w3595;
assign w4102 = pi0442 & ~w4100;
assign w4103 = (w4102 & w4101) | (w4102 & w12280) | (w4101 & w12280);
assign w4104 = ~pi0442 & ~w3842;
assign w4105 = (w4104 & ~w4101) | (w4104 & w12281) | (~w4101 & w12281);
assign w4106 = ~w4103 & ~w4105;
assign w4107 = w2868 & w12282;
assign w4108 = pi0022 & w3191;
assign w4109 = ~pi0443 & w3193;
assign w4110 = pi1747 & ~w4107;
assign w4111 = ~w4108 & w4110;
assign w4112 = ~w4109 & w4111;
assign w4113 = w3955 & w11977;
assign w4114 = ~pi0444 & w3958;
assign w4115 = w2868 & w12283;
assign w4116 = pi1747 & ~w4115;
assign w4117 = w3955 & w12284;
assign w4118 = ~w4114 & w4116;
assign w4119 = ~w4113 & w4118;
assign w4120 = ~w4117 & w4119;
assign w4121 = w2868 & w12285;
assign w4122 = pi0124 & w3191;
assign w4123 = ~pi0445 & w3193;
assign w4124 = pi1747 & ~w4121;
assign w4125 = ~w4122 & w4124;
assign w4126 = ~w4123 & w4125;
assign w4127 = w2868 & w12286;
assign w4128 = pi0254 & w3191;
assign w4129 = ~pi0446 & w3193;
assign w4130 = pi1747 & ~w4127;
assign w4131 = ~w4128 & w4130;
assign w4132 = ~w4129 & w4131;
assign w4133 = w2870 & w12287;
assign w4134 = ~pi0447 & w2875;
assign w4135 = w2868 & w12288;
assign w4136 = pi1747 & ~w4135;
assign w4137 = w2870 & w12289;
assign w4138 = ~w4134 & w4136;
assign w4139 = ~w4133 & w4138;
assign w4140 = ~w4137 & w4139;
assign w4141 = w4037 & w12290;
assign w4142 = w4037 & w12291;
assign w4143 = pi0448 & w4142;
assign w4144 = (~pi0705 & w4142) | (~pi0705 & w12292) | (w4142 & w12292);
assign w4145 = ~w4143 & w4144;
assign w4146 = w3955 & w12293;
assign w4147 = ~pi0449 & w3958;
assign w4148 = w2868 & w12294;
assign w4149 = pi1747 & ~w4148;
assign w4150 = w3955 & w11954;
assign w4151 = ~w4147 & w4149;
assign w4152 = ~w4146 & w4151;
assign w4153 = ~w4150 & w4152;
assign w4154 = w3955 & w12295;
assign w4155 = ~pi0450 & w3958;
assign w4156 = w2868 & w12296;
assign w4157 = pi1747 & ~w4156;
assign w4158 = w3955 & w11950;
assign w4159 = ~w4155 & w4157;
assign w4160 = ~w4154 & w4159;
assign w4161 = ~w4158 & w4160;
assign w4162 = w3955 & w12297;
assign w4163 = ~pi0451 & w3958;
assign w4164 = w2868 & w12298;
assign w4165 = pi1747 & ~w4164;
assign w4166 = w3955 & w11938;
assign w4167 = ~w4163 & w4165;
assign w4168 = ~w4162 & w4167;
assign w4169 = ~w4166 & w4168;
assign w4170 = w3955 & w11935;
assign w4171 = ~pi0452 & w3958;
assign w4172 = w2868 & w12299;
assign w4173 = pi1747 & ~w4172;
assign w4174 = w3955 & w12300;
assign w4175 = ~w4171 & w4173;
assign w4176 = ~w4170 & w4175;
assign w4177 = ~w4174 & w4176;
assign w4178 = w3955 & w12301;
assign w4179 = ~pi0453 & w3958;
assign w4180 = w2868 & w12302;
assign w4181 = pi1747 & ~w4180;
assign w4182 = w3955 & w11941;
assign w4183 = ~w4179 & w4181;
assign w4184 = ~w4178 & w4183;
assign w4185 = ~w4182 & w4184;
assign w4186 = w3952 & w11944;
assign w4187 = w2868 & w12303;
assign w4188 = pi1459 & ~w2934;
assign w4189 = (~w4188 & ~w2868) | (~w4188 & w12304) | (~w2868 & w12304);
assign w4190 = ~pi0454 & w4189;
assign w4191 = (w4188 & ~w2868) | (w4188 & w12305) | (~w2868 & w12305);
assign w4192 = pi0011 & w4191;
assign w4193 = pi1747 & ~w4187;
assign w4194 = ~w4190 & w4193;
assign w4195 = ~w4192 & w4194;
assign w4196 = w3955 & w11951;
assign w4197 = ~pi0455 & w3958;
assign w4198 = w2868 & w12306;
assign w4199 = pi1747 & ~w4198;
assign w4200 = w3955 & w12307;
assign w4201 = ~w4197 & w4199;
assign w4202 = ~w4196 & w4201;
assign w4203 = ~w4200 & w4202;
assign w4204 = w2868 & w12308;
assign w4205 = ~pi0456 & w4189;
assign w4206 = pi0016 & w4191;
assign w4207 = pi1747 & ~w4204;
assign w4208 = ~w4205 & w4207;
assign w4209 = ~w4206 & w4208;
assign w4210 = w2868 & w12309;
assign w4211 = pi0007 & w4191;
assign w4212 = ~pi0457 & w4189;
assign w4213 = pi1747 & ~w4210;
assign w4214 = ~w4211 & w4213;
assign w4215 = ~w4212 & w4214;
assign w4216 = w2870 & w12310;
assign w4217 = ~pi0458 & w2875;
assign w4218 = w2868 & w12311;
assign w4219 = pi1747 & ~w4218;
assign w4220 = w2870 & w12312;
assign w4221 = ~w4217 & w4219;
assign w4222 = ~w4216 & w4221;
assign w4223 = ~w4220 & w4222;
assign w4224 = w3955 & w12313;
assign w4225 = ~pi0459 & w3958;
assign w4226 = w2868 & w12314;
assign w4227 = pi1747 & ~w4226;
assign w4228 = w3955 & w11959;
assign w4229 = ~w4225 & w4227;
assign w4230 = ~w4224 & w4229;
assign w4231 = ~w4228 & w4230;
assign w4232 = w2868 & w12315;
assign w4233 = pi0019 & w4191;
assign w4234 = ~pi0460 & w4189;
assign w4235 = pi1747 & ~w4232;
assign w4236 = ~w4233 & w4235;
assign w4237 = ~w4234 & w4236;
assign w4238 = w2868 & w12316;
assign w4239 = pi0023 & w4191;
assign w4240 = ~pi0461 & w4189;
assign w4241 = pi1747 & ~w4238;
assign w4242 = ~w4239 & w4241;
assign w4243 = ~w4240 & w4242;
assign w4244 = w2868 & w12317;
assign w4245 = ~pi0462 & w4189;
assign w4246 = pi0046 & w4191;
assign w4247 = pi1747 & ~w4244;
assign w4248 = ~w4245 & w4247;
assign w4249 = ~w4246 & w4248;
assign w4250 = w2868 & w12318;
assign w4251 = pi0028 & w4191;
assign w4252 = ~pi0463 & w4189;
assign w4253 = pi1747 & ~w4250;
assign w4254 = ~w4251 & w4253;
assign w4255 = ~w4252 & w4254;
assign w4256 = w2868 & w12319;
assign w4257 = ~pi0464 & w4189;
assign w4258 = pi0030 & w4191;
assign w4259 = pi1747 & ~w4256;
assign w4260 = ~w4257 & w4259;
assign w4261 = ~w4258 & w4260;
assign w4262 = w4142 & w12321;
assign w4263 = w4142 & w12322;
assign w4264 = w4263 & w12324;
assign w4265 = (w4263 & w12325) | (w4263 & w12326) | (w12325 & w12326);
assign w4266 = ~w4264 & w4265;
assign w4267 = ~pi0466 & ~w3484;
assign w4268 = (w3681 & ~w3484) | (w3681 & w12327) | (~w3484 & w12327);
assign w4269 = ~w4267 & w4268;
assign w4270 = w3469 & ~w3475;
assign w4271 = w3471 & w12328;
assign w4272 = w4270 & w4271;
assign w4273 = pi0466 & w3675;
assign w4274 = (w4273 & ~w4270) | (w4273 & w12329) | (~w4270 & w12329);
assign w4275 = ~w4269 & ~w4272;
assign w4276 = ~w4274 & w4275;
assign w4277 = (~pi0467 & ~w4142) | (~pi0467 & w12330) | (~w4142 & w12330);
assign w4278 = (~pi0705 & ~w4142) | (~pi0705 & w12331) | (~w4142 & w12331);
assign w4279 = ~w4277 & w4278;
assign w4280 = (w3524 & w12334) | (w3524 & w12335) | (w12334 & w12335);
assign w4281 = (w3524 & w12336) | (w3524 & w12337) | (w12336 & w12337);
assign w4282 = w4280 & w4281;
assign w4283 = (~pi0468 & ~w3499) | (~pi0468 & w12338) | (~w3499 & w12338);
assign w4284 = ~w4282 & w4283;
assign w4285 = (w3492 & ~w3499) | (w3492 & w12339) | (~w3499 & w12339);
assign w4286 = pi0562 & w3491;
assign w4287 = (pi0468 & ~w3491) | (pi0468 & w12340) | (~w3491 & w12340);
assign w4288 = (w3499 & w12341) | (w3499 & w12342) | (w12341 & w12342);
assign w4289 = (w4288 & w3540) | (w4288 & w12343) | (w3540 & w12343);
assign w4290 = ~w4284 & ~w4289;
assign w4291 = ~pi0469 & ~pi1671;
assign w4292 = ~pi0705 & ~w4035;
assign w4293 = ~w4291 & w4292;
assign w4294 = (w3551 & w3550) | (w3551 & w12344) | (w3550 & w12344);
assign w4295 = w3546 & ~w3550;
assign w4296 = ~w4294 & ~w4295;
assign w4297 = pi0564 & pi1679;
assign w4298 = ~pi0564 & ~pi1679;
assign w4299 = ~w4297 & ~w4298;
assign w4300 = ~pi0514 & ~pi0541;
assign w4301 = ~pi0588 & w4300;
assign w4302 = ~pi0511 & ~pi0512;
assign w4303 = ~pi0513 & w4302;
assign w4304 = w4301 & w4303;
assign w4305 = ~pi0486 & ~pi0565;
assign w4306 = w4304 & w12345;
assign w4307 = w4304 & w12346;
assign w4308 = pi1679 & w3535;
assign w4309 = (pi0472 & ~w3535) | (pi0472 & w12347) | (~w3535 & w12347);
assign w4310 = (~w4309 & w4307) | (~w4309 & w12348) | (w4307 & w12348);
assign w4311 = pi0471 & pi1131;
assign w4312 = (w4311 & ~w4310) | (w4311 & w12349) | (~w4310 & w12349);
assign w4313 = pi0514 & pi1028;
assign w4314 = ~pi0514 & ~pi1028;
assign w4315 = ~w4313 & ~w4314;
assign w4316 = ~pi0512 & ~pi1310;
assign w4317 = pi0512 & pi1310;
assign w4318 = pi0511 & pi1027;
assign w4319 = ~w4317 & ~w4318;
assign w4320 = (~pi1129 & w4319) | (~pi1129 & w12350) | (w4319 & w12350);
assign w4321 = ~w4319 & w12351;
assign w4322 = ~pi0513 & ~w4321;
assign w4323 = ~w4322 & w12352;
assign w4324 = (pi1083 & w4323) | (pi1083 & w12353) | (w4323 & w12353);
assign w4325 = ~w4323 & w12354;
assign w4326 = pi0541 & ~w4325;
assign w4327 = (pi1130 & w4326) | (pi1130 & w12355) | (w4326 & w12355);
assign w4328 = ~pi0588 & ~w4327;
assign w4329 = ~w4326 & w12356;
assign w4330 = pi1076 & ~w4329;
assign w4331 = ~w4328 & w4330;
assign w4332 = ~pi0486 & ~w4331;
assign w4333 = pi0588 & ~w4329;
assign w4334 = ~pi1076 & ~w4327;
assign w4335 = ~w4333 & w4334;
assign w4336 = pi1029 & ~w4335;
assign w4337 = ~w4332 & w4336;
assign w4338 = ~pi0565 & ~w4337;
assign w4339 = pi0560 & pi1127;
assign w4340 = ~pi0560 & ~pi1127;
assign w4341 = ~w4339 & ~w4340;
assign w4342 = pi0486 & ~w4335;
assign w4343 = ~pi1029 & ~w4331;
assign w4344 = ~w4342 & w4343;
assign w4345 = w4341 & ~w4344;
assign w4346 = ~w4338 & w4345;
assign w4347 = pi0472 & ~w4339;
assign w4348 = w4311 & w4347;
assign w4349 = ~w4346 & w4347;
assign w4350 = ~pi0471 & pi1131;
assign w4351 = w4310 & w12357;
assign w4352 = ~w4349 & w4351;
assign w4353 = (~w4312 & w4346) | (~w4312 & w12358) | (w4346 & w12358);
assign w4354 = ~w4352 & w4353;
assign w4355 = ~w4307 & ~w4339;
assign w4356 = pi0472 & pi1131;
assign w4357 = ~w4346 & w12359;
assign w4358 = ~w4307 & w12360;
assign w4359 = (pi0472 & w4307) | (pi0472 & w12361) | (w4307 & w12361);
assign w4360 = pi1131 & ~w4358;
assign w4361 = ~w4359 & w4360;
assign w4362 = (~w4361 & w4346) | (~w4361 & w12362) | (w4346 & w12362);
assign w4363 = ~w4357 & ~w4362;
assign w4364 = ~pi0473 & ~w4263;
assign w4365 = (~pi0705 & ~w4263) | (~pi0705 & w12363) | (~w4263 & w12363);
assign w4366 = ~w4364 & w4365;
assign w4367 = ~pi0474 & ~w4035;
assign w4368 = (~pi0705 & ~w4035) | (~pi0705 & w12364) | (~w4035 & w12364);
assign w4369 = ~w4367 & w4368;
assign w4370 = ~pi0475 & ~w4037;
assign w4371 = (~pi0705 & ~w4037) | (~pi0705 & w12365) | (~w4037 & w12365);
assign w4372 = ~w4370 & w4371;
assign w4373 = (~pi0476 & ~w4037) | (~pi0476 & w12366) | (~w4037 & w12366);
assign w4374 = ~pi0705 & ~w4141;
assign w4375 = ~w4373 & w4374;
assign w4376 = (~pi0477 & ~w4037) | (~pi0477 & w12367) | (~w4037 & w12367);
assign w4377 = ~pi0705 & ~w4142;
assign w4378 = ~w4376 & w4377;
assign w4379 = (~pi0478 & ~w4142) | (~pi0478 & w12368) | (~w4142 & w12368);
assign w4380 = ~pi0705 & ~w4263;
assign w4381 = ~w4379 & w4380;
assign w4382 = (~pi0479 & ~w4142) | (~pi0479 & w12369) | (~w4142 & w12369);
assign w4383 = ~pi0705 & ~w4262;
assign w4384 = ~w4382 & w4383;
assign w4385 = (w3457 & w12370) | (w3457 & w12371) | (w12370 & w12371);
assign w4386 = ~w3459 & ~w4385;
assign w4387 = w3676 & ~w4386;
assign w4388 = ~w3665 & w3680;
assign w4389 = w3482 & w12372;
assign w4390 = (pi0480 & w4388) | (pi0480 & w12373) | (w4388 & w12373);
assign w4391 = ~pi0480 & pi0484;
assign w4392 = w3482 & w12374;
assign w4393 = ~w4390 & ~w4392;
assign w4394 = ~w4387 & w4393;
assign w4395 = ~pi0481 & pi1122;
assign w4396 = (w4395 & w3634) | (w4395 & w12375) | (w3634 & w12375);
assign w4397 = pi0481 & pi1122;
assign w4398 = ~w3634 & w12376;
assign w4399 = ~w4396 & ~w4398;
assign w4400 = ~pi0388 & w3689;
assign w4401 = w3472 & ~w3610;
assign w4402 = (~w4400 & ~w4401) | (~w4400 & w12377) | (~w4401 & w12377);
assign w4403 = pi0482 & ~w4402;
assign w4404 = (pi1122 & ~w4402) | (pi1122 & w12378) | (~w4402 & w12378);
assign w4405 = ~w4403 & w4404;
assign w4406 = w3491 & ~w3535;
assign w4407 = (w3492 & ~w3495) | (w3492 & w12379) | (~w3495 & w12379);
assign w4408 = ~w4406 & ~w4407;
assign w4409 = w3492 & ~w3493;
assign w4410 = w4408 & ~w4409;
assign w4411 = (pi0483 & ~w4408) | (pi0483 & w12380) | (~w4408 & w12380);
assign w4412 = (~w3528 & w3524) | (~w3528 & w12381) | (w3524 & w12381);
assign w4413 = ~w3527 & ~w4412;
assign w4414 = w3491 & w3535;
assign w4415 = (w4414 & w4413) | (w4414 & w12382) | (w4413 & w12382);
assign w4416 = ~pi0483 & w3493;
assign w4417 = w3497 & w12383;
assign w4418 = ~w4411 & ~w4417;
assign w4419 = ~w4415 & w4418;
assign w4420 = ~w3443 & w3457;
assign w4421 = ~w3458 & ~w4420;
assign w4422 = w3676 & ~w4421;
assign w4423 = (~w4389 & ~w4388) | (~w4389 & w12384) | (~w4388 & w12384);
assign w4424 = ~w4422 & w4423;
assign w4425 = pi0549 & w4408;
assign w4426 = (~pi0485 & ~w4408) | (~pi0485 & w12385) | (~w4408 & w12385);
assign w4427 = ~w4410 & ~w4426;
assign w4428 = ~w3505 & ~w3528;
assign w4429 = ~w3524 & w4428;
assign w4430 = (w4414 & ~w3524) | (w4414 & w12386) | (~w3524 & w12386);
assign w4431 = ~w4429 & w4430;
assign w4432 = ~w4427 & ~w4431;
assign w4433 = w3492 & ~w4304;
assign w4434 = ~w4331 & ~w4335;
assign w4435 = ~w4433 & w12387;
assign w4436 = (w4435 & w4434) | (w4435 & w12388) | (w4434 & w12388);
assign w4437 = (~pi0486 & ~w4304) | (~pi0486 & w12389) | (~w4304 & w12389);
assign w4438 = (w4437 & ~w4434) | (w4437 & w12390) | (~w4434 & w12390);
assign w4439 = ~w4436 & ~w4438;
assign w4440 = w2868 & w12391;
assign w4441 = pi0064 & w3191;
assign w4442 = ~pi0487 & w3193;
assign w4443 = pi1747 & ~w4440;
assign w4444 = ~w4441 & w4443;
assign w4445 = ~w4442 & w4444;
assign w4446 = w2868 & w12392;
assign w4447 = pi0014 & w3191;
assign w4448 = ~pi0488 & w3193;
assign w4449 = pi1747 & ~w4446;
assign w4450 = ~w4447 & w4449;
assign w4451 = ~w4448 & w4450;
assign w4452 = w2868 & w12393;
assign w4453 = pi0015 & w3191;
assign w4454 = ~pi0489 & w3193;
assign w4455 = pi1747 & ~w4452;
assign w4456 = ~w4453 & w4455;
assign w4457 = ~w4454 & w4456;
assign w4458 = w2868 & w12394;
assign w4459 = pi0953 & w3191;
assign w4460 = ~pi0490 & w3193;
assign w4461 = pi1747 & ~w4458;
assign w4462 = ~w4459 & w4461;
assign w4463 = ~w4460 & w4462;
assign w4464 = w2868 & w12395;
assign w4465 = pi0310 & w3191;
assign w4466 = ~pi0491 & w3193;
assign w4467 = pi1747 & ~w4464;
assign w4468 = ~w4465 & w4467;
assign w4469 = ~w4466 & w4468;
assign w4470 = w2868 & w12396;
assign w4471 = pi0332 & w3191;
assign w4472 = ~pi0492 & w3193;
assign w4473 = pi1747 & ~w4470;
assign w4474 = ~w4471 & w4473;
assign w4475 = ~w4472 & w4474;
assign w4476 = w2868 & w12397;
assign w4477 = pi0299 & w3191;
assign w4478 = ~pi0493 & w3193;
assign w4479 = pi1747 & ~w4476;
assign w4480 = ~w4477 & w4479;
assign w4481 = ~w4478 & w4480;
assign w4482 = w2868 & w12398;
assign w4483 = pi0286 & w3191;
assign w4484 = ~pi0494 & w3193;
assign w4485 = pi1747 & ~w4482;
assign w4486 = ~w4483 & w4485;
assign w4487 = ~w4484 & w4486;
assign w4488 = w2868 & w12399;
assign w4489 = pi1481 & w3191;
assign w4490 = ~pi0495 & w3193;
assign w4491 = pi1747 & ~w4488;
assign w4492 = ~w4489 & w4491;
assign w4493 = ~w4490 & w4492;
assign w4494 = w2868 & w12400;
assign w4495 = pi0223 & w3191;
assign w4496 = ~pi0496 & w3193;
assign w4497 = pi1747 & ~w4494;
assign w4498 = ~w4495 & w4497;
assign w4499 = ~w4496 & w4498;
assign w4500 = w2868 & w12401;
assign w4501 = pi0154 & w3191;
assign w4502 = ~pi0497 & w3193;
assign w4503 = pi1747 & ~w4500;
assign w4504 = ~w4501 & w4503;
assign w4505 = ~w4502 & w4504;
assign w4506 = w2868 & w12402;
assign w4507 = pi0155 & w3191;
assign w4508 = ~pi0498 & w3193;
assign w4509 = pi1747 & ~w4506;
assign w4510 = ~w4507 & w4509;
assign w4511 = ~w4508 & w4510;
assign w4512 = w2868 & w12403;
assign w4513 = pi0056 & w3191;
assign w4514 = ~pi0499 & w3193;
assign w4515 = pi1747 & ~w4512;
assign w4516 = ~w4513 & w4515;
assign w4517 = ~w4514 & w4516;
assign w4518 = w2868 & w12404;
assign w4519 = pi0063 & w3191;
assign w4520 = ~pi0500 & w3193;
assign w4521 = pi1747 & ~w4518;
assign w4522 = ~w4519 & w4521;
assign w4523 = ~w4520 & w4522;
assign w4524 = w2868 & w12405;
assign w4525 = pi0194 & w3191;
assign w4526 = ~pi0501 & w3193;
assign w4527 = pi1747 & ~w4524;
assign w4528 = ~w4525 & w4527;
assign w4529 = ~w4526 & w4528;
assign w4530 = w2868 & w12406;
assign w4531 = pi0049 & w3191;
assign w4532 = ~pi0502 & w3193;
assign w4533 = pi1747 & ~w4530;
assign w4534 = ~w4531 & w4533;
assign w4535 = ~w4532 & w4534;
assign w4536 = w2868 & w12407;
assign w4537 = pi0027 & w3191;
assign w4538 = ~pi0503 & w3193;
assign w4539 = pi1747 & ~w4536;
assign w4540 = ~w4537 & w4539;
assign w4541 = ~w4538 & w4540;
assign w4542 = w2868 & w12408;
assign w4543 = ~pi1672 & w4191;
assign w4544 = ~pi0504 & w4189;
assign w4545 = pi1747 & ~w4542;
assign w4546 = ~w4543 & w4545;
assign w4547 = ~w4544 & w4546;
assign w4548 = w2868 & w12409;
assign w4549 = ~pi0505 & w4189;
assign w4550 = ~pi1666 & w4191;
assign w4551 = pi1747 & ~w4548;
assign w4552 = ~w4549 & w4551;
assign w4553 = ~w4550 & w4552;
assign w4554 = (pi1679 & ~w3535) | (pi1679 & w12410) | (~w3535 & w12410);
assign w4555 = (~w3535 & w12411) | (~w3535 & w12412) | (w12411 & w12412);
assign w4556 = (pi1131 & w4554) | (pi1131 & w12413) | (w4554 & w12413);
assign w4557 = ~w4555 & w4556;
assign w4558 = ~pi1690 & w3480;
assign w4559 = w3680 & ~w4558;
assign w4560 = (~pi0507 & ~w3681) | (~pi0507 & w12414) | (~w3681 & w12414);
assign w4561 = w4559 & ~w4560;
assign w4562 = ~w3447 & ~w3448;
assign w4563 = w3449 & ~w4562;
assign w4564 = ~w3449 & w4562;
assign w4565 = ~w4563 & ~w4564;
assign w4566 = w3676 & w4565;
assign w4567 = ~w4561 & ~w4566;
assign w4568 = ~pi0508 & w3480;
assign w4569 = w3681 & w4568;
assign w4570 = w3680 & w12415;
assign w4571 = ~w3446 & ~w3451;
assign w4572 = ~w3452 & ~w4571;
assign w4573 = (~w4569 & w4572) | (~w4569 & w12416) | (w4572 & w12416);
assign w4574 = ~w4570 & w4573;
assign w4575 = ~w3454 & ~w3455;
assign w4576 = w3676 & w4575;
assign w4577 = (~pi0509 & ~w3481) | (~pi0509 & w12417) | (~w3481 & w12417);
assign w4578 = ~w4576 & w4577;
assign w4579 = pi0509 & ~w4388;
assign w4580 = (w4579 & w4575) | (w4579 & w12418) | (w4575 & w12418);
assign w4581 = ~w4578 & ~w4580;
assign w4582 = w3688 & w12419;
assign w4583 = w3472 & ~w3597;
assign w4584 = (~w4582 & ~w4583) | (~w4582 & w12420) | (~w4583 & w12420);
assign w4585 = pi0510 & ~w4584;
assign w4586 = (pi1122 & ~w4584) | (pi1122 & w12421) | (~w4584 & w12421);
assign w4587 = ~w4585 & w4586;
assign w4588 = (w3535 & w12422) | (w3535 & w12423) | (w12422 & w12423);
assign w4589 = (~w3535 & w12424) | (~w3535 & w12425) | (w12424 & w12425);
assign w4590 = pi1131 & ~w4588;
assign w4591 = ~w4589 & w4590;
assign w4592 = ~w3535 & w12426;
assign w4593 = pi0511 & pi0512;
assign w4594 = ~w4302 & ~w4593;
assign w4595 = w3492 & ~w4594;
assign w4596 = ~w4316 & ~w4317;
assign w4597 = ~w4318 & ~w4596;
assign w4598 = w4318 & w4596;
assign w4599 = ~w4597 & ~w4598;
assign w4600 = w4414 & w4599;
assign w4601 = ~w4592 & ~w4595;
assign w4602 = ~w4600 & w4601;
assign w4603 = ~pi1679 & w4302;
assign w4604 = w4308 & ~w4320;
assign w4605 = (~w4603 & ~w4604) | (~w4603 & w12427) | (~w4604 & w12427);
assign w4606 = pi0513 & ~w4605;
assign w4607 = (pi1131 & ~w4605) | (pi1131 & w12428) | (~w4605 & w12428);
assign w4608 = ~w4606 & w4607;
assign w4609 = w4302 & w12429;
assign w4610 = w3492 & w4609;
assign w4611 = w3492 & ~w4303;
assign w4612 = ~w4406 & ~w4611;
assign w4613 = (~w4315 & w4322) | (~w4315 & w12430) | (w4322 & w12430);
assign w4614 = ~w4323 & w4414;
assign w4615 = ~w4613 & w4614;
assign w4616 = (~w4610 & w4612) | (~w4610 & w12431) | (w4612 & w12431);
assign w4617 = ~w4615 & w4616;
assign w4618 = w4058 & w11922;
assign w4619 = ~pi0515 & w4061;
assign w4620 = w2868 & w12432;
assign w4621 = pi1747 & ~w4620;
assign w4622 = w4058 & w12433;
assign w4623 = ~w4619 & w4621;
assign w4624 = ~w4618 & w4623;
assign w4625 = ~w4622 & w4624;
assign w4626 = w2870 & w12275;
assign w4627 = ~pi0516 & w2875;
assign w4628 = w2868 & w12434;
assign w4629 = pi1747 & ~w4628;
assign w4630 = w2870 & w12435;
assign w4631 = ~w4627 & w4629;
assign w4632 = ~w4626 & w4631;
assign w4633 = ~w4630 & w4632;
assign w4634 = w2870 & w12221;
assign w4635 = ~pi0517 & w2875;
assign w4636 = w2868 & w12436;
assign w4637 = pi1747 & ~w4636;
assign w4638 = w2870 & w12437;
assign w4639 = ~w4635 & w4637;
assign w4640 = ~w4634 & w4639;
assign w4641 = ~w4638 & w4640;
assign w4642 = w2870 & w12438;
assign w4643 = ~pi0518 & w2875;
assign w4644 = w2868 & w12439;
assign w4645 = pi1747 & ~w4644;
assign w4646 = w2870 & w12440;
assign w4647 = ~w4643 & w4645;
assign w4648 = ~w4642 & w4647;
assign w4649 = ~w4646 & w4648;
assign w4650 = w2870 & w12441;
assign w4651 = ~pi0519 & w2875;
assign w4652 = w2868 & w12442;
assign w4653 = pi1747 & ~w4652;
assign w4654 = w2870 & w12443;
assign w4655 = ~w4651 & w4653;
assign w4656 = ~w4650 & w4655;
assign w4657 = ~w4654 & w4656;
assign w4658 = w3955 & w12444;
assign w4659 = ~pi0520 & w3958;
assign w4660 = w2868 & w12445;
assign w4661 = pi1747 & ~w4660;
assign w4662 = w3955 & w11971;
assign w4663 = ~w4659 & w4661;
assign w4664 = ~w4658 & w4663;
assign w4665 = ~w4662 & w4664;
assign w4666 = w3955 & w12446;
assign w4667 = ~pi0521 & w3958;
assign w4668 = w2868 & w12447;
assign w4669 = pi1747 & ~w4668;
assign w4670 = w3955 & w12221;
assign w4671 = ~w4667 & w4669;
assign w4672 = ~w4666 & w4671;
assign w4673 = ~w4670 & w4672;
assign w4674 = w3955 & w12448;
assign w4675 = ~pi0522 & w3958;
assign w4676 = w2868 & w12449;
assign w4677 = pi1747 & ~w4676;
assign w4678 = w3955 & w12438;
assign w4679 = ~w4675 & w4677;
assign w4680 = ~w4674 & w4679;
assign w4681 = ~w4678 & w4680;
assign w4682 = w3955 & w12450;
assign w4683 = ~pi0523 & w3958;
assign w4684 = w2868 & w12451;
assign w4685 = pi1747 & ~w4684;
assign w4686 = w3955 & w11974;
assign w4687 = ~w4683 & w4685;
assign w4688 = ~w4682 & w4687;
assign w4689 = ~w4686 & w4688;
assign w4690 = w3955 & w12452;
assign w4691 = ~pi0524 & w3958;
assign w4692 = w2868 & w12453;
assign w4693 = pi1747 & ~w4692;
assign w4694 = w3955 & w11983;
assign w4695 = ~w4691 & w4693;
assign w4696 = ~w4690 & w4695;
assign w4697 = ~w4694 & w4696;
assign w4698 = w3955 & w12454;
assign w4699 = ~pi0525 & w3958;
assign w4700 = w2868 & w12455;
assign w4701 = pi1747 & ~w4700;
assign w4702 = w3955 & w12270;
assign w4703 = ~w4699 & w4701;
assign w4704 = ~w4698 & w4703;
assign w4705 = ~w4702 & w4704;
assign w4706 = w3955 & w11994;
assign w4707 = ~pi0526 & w3958;
assign w4708 = w2868 & w12456;
assign w4709 = pi1747 & ~w4708;
assign w4710 = w3955 & w12457;
assign w4711 = ~w4707 & w4709;
assign w4712 = ~w4706 & w4711;
assign w4713 = ~w4710 & w4712;
assign w4714 = w3955 & w11995;
assign w4715 = ~pi0527 & w3958;
assign w4716 = w2868 & w12458;
assign w4717 = pi1747 & ~w4716;
assign w4718 = w3955 & w12459;
assign w4719 = ~w4715 & w4717;
assign w4720 = ~w4714 & w4719;
assign w4721 = ~w4718 & w4720;
assign w4722 = w3955 & w12443;
assign w4723 = ~pi0528 & w3958;
assign w4724 = w2868 & w12460;
assign w4725 = pi1747 & ~w4724;
assign w4726 = w3955 & w12461;
assign w4727 = ~w4723 & w4725;
assign w4728 = ~w4722 & w4727;
assign w4729 = ~w4726 & w4728;
assign w4730 = w3955 & w11980;
assign w4731 = ~pi0529 & w3958;
assign w4732 = w2868 & w12462;
assign w4733 = pi1747 & ~w4732;
assign w4734 = w3955 & w12463;
assign w4735 = ~w4731 & w4733;
assign w4736 = ~w4730 & w4735;
assign w4737 = ~w4734 & w4736;
assign w4738 = w3955 & w12001;
assign w4739 = ~pi0530 & w3958;
assign w4740 = w2868 & w12464;
assign w4741 = pi1747 & ~w4740;
assign w4742 = w3955 & w12465;
assign w4743 = ~w4739 & w4741;
assign w4744 = ~w4738 & w4743;
assign w4745 = ~w4742 & w4744;
assign w4746 = w3955 & w12466;
assign w4747 = ~pi0531 & w3958;
assign w4748 = w2868 & w12467;
assign w4749 = pi1747 & ~w4748;
assign w4750 = w3955 & w12006;
assign w4751 = ~w4747 & w4749;
assign w4752 = ~w4746 & w4751;
assign w4753 = ~w4750 & w4752;
assign w4754 = w2868 & w12468;
assign w4755 = ~pi0532 & w4189;
assign w4756 = pi0018 & w4191;
assign w4757 = pi1747 & ~w4754;
assign w4758 = ~w4755 & w4757;
assign w4759 = ~w4756 & w4758;
assign w4760 = ~pi0533 & pi1127;
assign w4761 = (w3524 & w12471) | (w3524 & w12472) | (w12471 & w12472);
assign w4762 = (~pi0533 & ~w3497) | (~pi0533 & w12473) | (~w3497 & w12473);
assign w4763 = pi1131 & ~w3499;
assign w4764 = ~w4762 & w4763;
assign w4765 = (~w4764 & w4761) | (~w4764 & w12474) | (w4761 & w12474);
assign w4766 = pi0533 & ~w3536;
assign w4767 = (pi1679 & ~w3536) | (pi1679 & w12475) | (~w3536 & w12475);
assign w4768 = ~w4766 & w4767;
assign w4769 = ~w4765 & ~w4768;
assign w4770 = w3152 & w12476;
assign w4771 = ~pi0534 & w3155;
assign w4772 = w2868 & w12477;
assign w4773 = pi1747 & ~w4772;
assign w4774 = w3152 & w12261;
assign w4775 = ~w4771 & w4773;
assign w4776 = ~w4770 & w4775;
assign w4777 = ~w4774 & w4776;
assign w4778 = (pi1480 & w1221) | (pi1480 & w12478) | (w1221 & w12478);
assign w4779 = ~pi0535 & ~w4778;
assign w4780 = w1773 & ~w4779;
assign w4781 = w3152 & w12270;
assign w4782 = ~pi0536 & w3155;
assign w4783 = w2868 & w12479;
assign w4784 = pi1747 & ~w4783;
assign w4785 = w3152 & w12480;
assign w4786 = ~w4782 & w4784;
assign w4787 = ~w4781 & w4786;
assign w4788 = ~w4785 & w4787;
assign w4789 = w2868 & w12481;
assign w4790 = pi0049 & w4191;
assign w4791 = ~pi0537 & w4189;
assign w4792 = pi1747 & ~w4789;
assign w4793 = ~w4790 & w4792;
assign w4794 = ~w4791 & w4793;
assign w4795 = w2868 & w12482;
assign w4796 = ~pi0538 & w4189;
assign w4797 = pi0299 & w4191;
assign w4798 = pi1747 & ~w4795;
assign w4799 = ~w4796 & w4798;
assign w4800 = ~w4797 & w4799;
assign w4801 = w2868 & w12483;
assign w4802 = pi0124 & w4191;
assign w4803 = ~pi0539 & w4189;
assign w4804 = pi1747 & ~w4801;
assign w4805 = ~w4802 & w4804;
assign w4806 = ~w4803 & w4805;
assign w4807 = w2868 & w12484;
assign w4808 = ~pi0540 & w4189;
assign w4809 = pi0223 & w4191;
assign w4810 = pi1747 & ~w4807;
assign w4811 = ~w4808 & w4810;
assign w4812 = ~w4809 & w4811;
assign w4813 = ~pi1679 & w4609;
assign w4814 = (~w4323 & w12485) | (~w4323 & w12486) | (w12485 & w12486);
assign w4815 = ~w4325 & w4814;
assign w4816 = ~w4815 & w12487;
assign w4817 = (pi0541 & w4815) | (pi0541 & w12488) | (w4815 & w12488);
assign w4818 = pi1131 & ~w4816;
assign w4819 = ~w4817 & w4818;
assign w4820 = w4058 & w12443;
assign w4821 = ~pi0542 & w4061;
assign w4822 = w2868 & w12489;
assign w4823 = pi1747 & ~w4822;
assign w4824 = w4058 & w12490;
assign w4825 = ~w4821 & w4823;
assign w4826 = ~w4820 & w4825;
assign w4827 = ~w4824 & w4826;
assign w4828 = w2868 & w12491;
assign w4829 = pi0953 & w4191;
assign w4830 = ~pi0543 & w4189;
assign w4831 = pi1747 & ~w4828;
assign w4832 = ~w4829 & w4831;
assign w4833 = ~w4830 & w4832;
assign w4834 = w4058 & w11995;
assign w4835 = ~pi0544 & w4061;
assign w4836 = w2868 & w12492;
assign w4837 = pi1747 & ~w4836;
assign w4838 = w4058 & w12493;
assign w4839 = ~w4835 & w4837;
assign w4840 = ~w4834 & w4839;
assign w4841 = ~w4838 & w4840;
assign w4842 = ~w1520 & ~w1525;
assign w4843 = ~w1359 & w4842;
assign w4844 = w1359 & ~w4842;
assign w4845 = ~w4843 & ~w4844;
assign w4846 = w4058 & w11986;
assign w4847 = ~pi0546 & w4061;
assign w4848 = w2868 & w12494;
assign w4849 = pi1747 & ~w4848;
assign w4850 = w4058 & w12495;
assign w4851 = ~w4847 & w4849;
assign w4852 = ~w4846 & w4851;
assign w4853 = ~w4850 & w4852;
assign w4854 = w4058 & w12289;
assign w4855 = ~pi0547 & w4061;
assign w4856 = w2868 & w12496;
assign w4857 = pi1747 & ~w4856;
assign w4858 = w4058 & w12497;
assign w4859 = ~w4855 & w4857;
assign w4860 = ~w4854 & w4859;
assign w4861 = ~w4858 & w4860;
assign w4862 = w3152 & w12498;
assign w4863 = ~pi0548 & w3155;
assign w4864 = w2868 & w12499;
assign w4865 = pi1747 & ~w4864;
assign w4866 = w3152 & w12289;
assign w4867 = ~w4863 & w4865;
assign w4868 = ~w4862 & w4867;
assign w4869 = ~w4866 & w4868;
assign w4870 = ~w3520 & ~w3522;
assign w4871 = (w4425 & w4870) | (w4425 & w12500) | (w4870 & w12500);
assign w4872 = w4414 & w4870;
assign w4873 = (~pi0549 & ~w3497) | (~pi0549 & w12501) | (~w3497 & w12501);
assign w4874 = ~w4872 & w4873;
assign w4875 = ~w4871 & ~w4874;
assign w4876 = w4058 & w11954;
assign w4877 = ~pi0550 & w4061;
assign w4878 = w2868 & w12502;
assign w4879 = pi1747 & ~w4878;
assign w4880 = w4058 & w12503;
assign w4881 = ~w4877 & w4879;
assign w4882 = ~w4876 & w4881;
assign w4883 = ~w4880 & w4882;
assign w4884 = w4058 & w11938;
assign w4885 = ~pi0551 & w4061;
assign w4886 = w2868 & w12504;
assign w4887 = pi1747 & ~w4886;
assign w4888 = w4058 & w12505;
assign w4889 = ~w4885 & w4887;
assign w4890 = ~w4884 & w4889;
assign w4891 = ~w4888 & w4890;
assign w4892 = pi0642 & pi1139;
assign w4893 = pi0591 & pi1258;
assign w4894 = ~pi0591 & ~pi1258;
assign w4895 = ~w4893 & ~w4894;
assign w4896 = ~pi0589 & ~pi1342;
assign w4897 = pi0589 & pi1342;
assign w4898 = pi0594 & pi1032;
assign w4899 = ~w4897 & ~w4898;
assign w4900 = (~pi1141 & w4899) | (~pi1141 & w12506) | (w4899 & w12506);
assign w4901 = ~w4899 & w12507;
assign w4902 = ~pi0590 & ~w4901;
assign w4903 = ~w4902 & w12508;
assign w4904 = (pi1033 & w4903) | (pi1033 & w12509) | (w4903 & w12509);
assign w4905 = ~w4903 & w12510;
assign w4906 = pi0627 & ~w4905;
assign w4907 = (pi1142 & w4906) | (pi1142 & w12511) | (w4906 & w12511);
assign w4908 = ~pi0655 & ~w4907;
assign w4909 = ~w4906 & w12512;
assign w4910 = pi1265 & ~w4909;
assign w4911 = ~w4908 & w4910;
assign w4912 = ~pi0568 & ~w4911;
assign w4913 = pi0655 & ~w4909;
assign w4914 = ~pi1265 & ~w4907;
assign w4915 = ~w4913 & w4914;
assign w4916 = pi1034 & ~w4915;
assign w4917 = ~w4912 & w4916;
assign w4918 = ~pi0631 & ~w4917;
assign w4919 = ~pi0642 & ~pi1139;
assign w4920 = ~w4892 & ~w4919;
assign w4921 = pi0568 & ~w4915;
assign w4922 = ~pi1034 & ~w4911;
assign w4923 = ~w4921 & w4922;
assign w4924 = w4920 & ~w4923;
assign w4925 = ~w4918 & w4924;
assign w4926 = w3241 & w12513;
assign w4927 = (w4926 & w4925) | (w4926 & w12514) | (w4925 & w12514);
assign w4928 = pi0552 & w3242;
assign w4929 = ~pi0594 & ~pi1697;
assign w4930 = ~pi0589 & w4929;
assign w4931 = w4929 & w12515;
assign w4932 = ~pi0591 & w4931;
assign w4933 = w4931 & w6235;
assign w4934 = w4931 & w12516;
assign w4935 = ~pi0568 & w4934;
assign w4936 = w4934 & w12518;
assign w4937 = w4934 & w12519;
assign w4938 = (pi0552 & ~w4934) | (pi0552 & w12520) | (~w4934 & w12520);
assign w4939 = ~w4937 & ~w4938;
assign w4940 = ~w4939 & w12521;
assign w4941 = ~w4939 & w12522;
assign w4942 = (~w4940 & w4925) | (~w4940 & w12523) | (w4925 & w12523);
assign w4943 = ~w4927 & w4942;
assign w4944 = w4058 & w11935;
assign w4945 = ~pi0553 & w4061;
assign w4946 = w2868 & w12524;
assign w4947 = pi1747 & ~w4946;
assign w4948 = w4058 & w12525;
assign w4949 = ~w4945 & w4947;
assign w4950 = ~w4944 & w4949;
assign w4951 = ~w4948 & w4950;
assign w4952 = w4058 & w11941;
assign w4953 = ~pi0554 & w4061;
assign w4954 = w2868 & w12526;
assign w4955 = pi1747 & ~w4954;
assign w4956 = w4058 & w12527;
assign w4957 = ~w4953 & w4955;
assign w4958 = ~w4952 & w4957;
assign w4959 = ~w4956 & w4958;
assign w4960 = w4058 & w11950;
assign w4961 = ~pi0555 & w4061;
assign w4962 = w2868 & w12528;
assign w4963 = pi1747 & ~w4962;
assign w4964 = w4058 & w12529;
assign w4965 = ~w4961 & w4963;
assign w4966 = ~w4960 & w4965;
assign w4967 = ~w4964 & w4966;
assign w4968 = w4058 & w11951;
assign w4969 = ~pi0556 & w4061;
assign w4970 = w2868 & w12530;
assign w4971 = pi1747 & ~w4970;
assign w4972 = w4058 & w12531;
assign w4973 = ~w4969 & w4971;
assign w4974 = ~w4968 & w4973;
assign w4975 = ~w4972 & w4974;
assign w4976 = w4058 & w12310;
assign w4977 = ~pi0557 & w4061;
assign w4978 = w2868 & w12532;
assign w4979 = pi1747 & ~w4978;
assign w4980 = w4058 & w12533;
assign w4981 = ~w4977 & w4979;
assign w4982 = ~w4976 & w4981;
assign w4983 = ~w4980 & w4982;
assign w4984 = w4058 & w11959;
assign w4985 = ~pi0558 & w4061;
assign w4986 = w2868 & w12534;
assign w4987 = pi1747 & ~w4986;
assign w4988 = w4058 & w12535;
assign w4989 = ~w4985 & w4987;
assign w4990 = ~w4984 & w4989;
assign w4991 = ~w4988 & w4990;
assign w4992 = w3152 & w12536;
assign w4993 = ~pi0559 & w3155;
assign w4994 = w2868 & w12537;
assign w4995 = pi1747 & ~w4994;
assign w4996 = w3152 & w12310;
assign w4997 = ~w4993 & w4995;
assign w4998 = ~w4992 & w4997;
assign w4999 = ~w4996 & w4998;
assign w5000 = (pi0560 & ~w4304) | (pi0560 & w12538) | (~w4304 & w12538);
assign w5001 = ~w4306 & ~w5000;
assign w5002 = ~w3535 & w12539;
assign w5003 = (~w5002 & w5001) | (~w5002 & w12540) | (w5001 & w12540);
assign w5004 = (w5003 & w4346) | (w5003 & w12541) | (w4346 & w12541);
assign w5005 = ~w4338 & ~w4344;
assign w5006 = w3535 & ~w4341;
assign w5007 = (w5006 & w5001) | (w5006 & w12542) | (w5001 & w12542);
assign w5008 = ~w5005 & w5007;
assign w5009 = ~w5004 & ~w5008;
assign w5010 = ~pi0753 & ~pi1773;
assign w5011 = pi1773 & ~pi1807;
assign w5012 = ~w5010 & ~w5011;
assign w5013 = (~pi0562 & ~w3499) | (~pi0562 & w12543) | (~w3499 & w12543);
assign w5014 = w4285 & ~w5013;
assign w5015 = ~w3540 & w4286;
assign w5016 = ~w4282 & ~w5014;
assign w5017 = ~w5015 & w5016;
assign w5018 = ~pi0649 & w4937;
assign w5019 = w3242 & w12544;
assign w5020 = pi0563 & pi1143;
assign w5021 = ~w5018 & w12545;
assign w5022 = (~w4892 & ~w4937) | (~w4892 & w12546) | (~w4937 & w12546);
assign w5023 = (~w4937 & w12547) | (~w4937 & w12548) | (w12547 & w12548);
assign w5024 = ~w4925 & w5022;
assign w5025 = ~pi0563 & pi1143;
assign w5026 = (w5025 & w5018) | (w5025 & w12549) | (w5018 & w12549);
assign w5027 = ~w5024 & w5026;
assign w5028 = (~w5021 & w4925) | (~w5021 & w12550) | (w4925 & w12550);
assign w5029 = ~w5027 & w5028;
assign w5030 = pi0564 & pi1131;
assign w5031 = ~w4310 & w5030;
assign w5032 = w4347 & w5030;
assign w5033 = ~pi0564 & pi1131;
assign w5034 = w4310 & w5033;
assign w5035 = (w5034 & w4346) | (w5034 & w12551) | (w4346 & w12551);
assign w5036 = (~w5031 & w4346) | (~w5031 & w12552) | (w4346 & w12552);
assign w5037 = ~w5035 & w5036;
assign w5038 = ~w4337 & ~w4344;
assign w5039 = w3491 & ~w5038;
assign w5040 = pi0486 & w3492;
assign w5041 = ~w4433 & w12553;
assign w5042 = (pi0565 & w5039) | (pi0565 & w12554) | (w5039 & w12554);
assign w5043 = ~pi0565 & w4414;
assign w5044 = w5038 & w5043;
assign w5045 = w4304 & w12555;
assign w5046 = ~w5044 & ~w5045;
assign w5047 = ~w5042 & w5046;
assign w5048 = ~w3212 & w3238;
assign w5049 = ~w3239 & ~w5048;
assign w5050 = w3251 & ~w5049;
assign w5051 = (~pi0566 & ~w3203) | (~pi0566 & w12556) | (~w3203 & w12556);
assign w5052 = ~w3205 & w3243;
assign w5053 = ~w5051 & w5052;
assign w5054 = ~w5050 & ~w5053;
assign w5055 = w3492 & ~w3495;
assign w5056 = ~w4406 & ~w5055;
assign w5057 = pi0622 & w5056;
assign w5058 = (~pi0567 & ~w5056) | (~pi0567 & w12557) | (~w5056 & w12557);
assign w5059 = ~w4408 & ~w5058;
assign w5060 = ~w3518 & w12558;
assign w5061 = ~w3519 & w4414;
assign w5062 = ~w5060 & w5061;
assign w5063 = ~w5059 & ~w5062;
assign w5064 = ~w4911 & ~w4915;
assign w5065 = ~w3242 & ~w4934;
assign w5066 = pi0568 & ~w5065;
assign w5067 = (w5066 & w5064) | (w5066 & w12559) | (w5064 & w12559);
assign w5068 = ~pi0568 & ~w4934;
assign w5069 = (w5068 & ~w5064) | (w5068 & w12560) | (~w5064 & w12560);
assign w5070 = pi1143 & ~w5067;
assign w5071 = ~w5069 & w5070;
assign w5072 = ~pi0569 & ~w3203;
assign w5073 = w3243 & ~w5072;
assign w5074 = (w3235 & w12561) | (w3235 & w12562) | (w12561 & w12562);
assign w5075 = ~w3237 & ~w5074;
assign w5076 = (~w5073 & w5075) | (~w5073 & w12563) | (w5075 & w12563);
assign w5077 = ~w3204 & ~w5076;
assign w5078 = w2868 & w12564;
assign w5079 = pi0064 & w4191;
assign w5080 = ~pi0570 & w4189;
assign w5081 = pi1747 & ~w5078;
assign w5082 = ~w5079 & w5081;
assign w5083 = ~w5080 & w5082;
assign w5084 = w2868 & w12565;
assign w5085 = pi0014 & w4191;
assign w5086 = ~pi0571 & w4189;
assign w5087 = pi1747 & ~w5084;
assign w5088 = ~w5085 & w5087;
assign w5089 = ~w5086 & w5088;
assign w5090 = w2868 & w12566;
assign w5091 = ~pi0572 & w4189;
assign w5092 = pi0015 & w4191;
assign w5093 = pi1747 & ~w5090;
assign w5094 = ~w5091 & w5093;
assign w5095 = ~w5092 & w5094;
assign w5096 = w2868 & w12567;
assign w5097 = ~pi0573 & w4189;
assign w5098 = pi0310 & w4191;
assign w5099 = pi1747 & ~w5096;
assign w5100 = ~w5097 & w5099;
assign w5101 = ~w5098 & w5100;
assign w5102 = w2868 & w12568;
assign w5103 = ~pi0574 & w4189;
assign w5104 = pi0332 & w4191;
assign w5105 = pi1747 & ~w5102;
assign w5106 = ~w5103 & w5105;
assign w5107 = ~w5104 & w5106;
assign w5108 = w2868 & w12569;
assign w5109 = pi0057 & w4191;
assign w5110 = ~pi0575 & w4189;
assign w5111 = pi1747 & ~w5108;
assign w5112 = ~w5109 & w5111;
assign w5113 = ~w5110 & w5112;
assign w5114 = w2868 & w12570;
assign w5115 = pi1481 & w4191;
assign w5116 = ~pi0576 & w4189;
assign w5117 = pi1747 & ~w5114;
assign w5118 = ~w5115 & w5117;
assign w5119 = ~w5116 & w5118;
assign w5120 = w2868 & w12571;
assign w5121 = ~pi0577 & w4189;
assign w5122 = pi0254 & w4191;
assign w5123 = pi1747 & ~w5120;
assign w5124 = ~w5121 & w5123;
assign w5125 = ~w5122 & w5124;
assign w5126 = w2868 & w12572;
assign w5127 = ~pi0578 & w4189;
assign w5128 = pi0286 & w4191;
assign w5129 = pi1747 & ~w5126;
assign w5130 = ~w5127 & w5129;
assign w5131 = ~w5128 & w5130;
assign w5132 = w2868 & w12573;
assign w5133 = pi0155 & w4191;
assign w5134 = ~pi0579 & w4189;
assign w5135 = pi1747 & ~w5132;
assign w5136 = ~w5133 & w5135;
assign w5137 = ~w5134 & w5136;
assign w5138 = w2868 & w12574;
assign w5139 = pi0154 & w4191;
assign w5140 = ~pi0580 & w4189;
assign w5141 = pi1747 & ~w5138;
assign w5142 = ~w5139 & w5141;
assign w5143 = ~w5140 & w5142;
assign w5144 = w2868 & w12575;
assign w5145 = pi0194 & w4191;
assign w5146 = ~pi0581 & w4189;
assign w5147 = pi1747 & ~w5144;
assign w5148 = ~w5145 & w5147;
assign w5149 = ~w5146 & w5148;
assign w5150 = w2868 & w12576;
assign w5151 = ~pi0582 & w4189;
assign w5152 = pi0056 & w4191;
assign w5153 = pi1747 & ~w5150;
assign w5154 = ~w5151 & w5153;
assign w5155 = ~w5152 & w5154;
assign w5156 = w2868 & w12577;
assign w5157 = pi0063 & w4191;
assign w5158 = ~pi0583 & w4189;
assign w5159 = pi1747 & ~w5156;
assign w5160 = ~w5157 & w5159;
assign w5161 = ~w5158 & w5160;
assign w5162 = w2868 & w12578;
assign w5163 = pi0027 & w4191;
assign w5164 = ~pi0584 & w4189;
assign w5165 = pi1747 & ~w5162;
assign w5166 = ~w5163 & w5165;
assign w5167 = ~w5164 & w5166;
assign w5168 = w2868 & w12579;
assign w5169 = pi0022 & w4191;
assign w5170 = ~pi0585 & w4189;
assign w5171 = pi1747 & ~w5168;
assign w5172 = ~w5169 & w5171;
assign w5173 = ~w5170 & w5172;
assign w5174 = (pi1697 & ~w3241) | (pi1697 & w12580) | (~w3241 & w12580);
assign w5175 = (~w3241 & w12581) | (~w3241 & w12582) | (w12581 & w12582);
assign w5176 = (pi1143 & w5174) | (pi1143 & w12583) | (w5174 & w12583);
assign w5177 = ~w5175 & w5176;
assign w5178 = ~w3495 & w12584;
assign w5179 = ~w3513 & ~w3514;
assign w5180 = w3491 & ~w5179;
assign w5181 = (pi0587 & w5180) | (pi0587 & w12585) | (w5180 & w12585);
assign w5182 = ~pi0587 & w4414;
assign w5183 = w5179 & w5182;
assign w5184 = ~w5178 & ~w5183;
assign w5185 = ~w5181 & w5184;
assign w5186 = w4609 & w12586;
assign w5187 = w4308 & ~w4327;
assign w5188 = (~w5186 & ~w5187) | (~w5186 & w12587) | (~w5187 & w12587);
assign w5189 = pi0588 & ~w5188;
assign w5190 = (pi1131 & ~w5188) | (pi1131 & w12588) | (~w5188 & w12588);
assign w5191 = ~w5189 & w5190;
assign w5192 = ~w4896 & ~w4897;
assign w5193 = w4898 & w5192;
assign w5194 = ~w4898 & ~w5192;
assign w5195 = ~w5193 & ~w5194;
assign w5196 = (~w4930 & ~w5195) | (~w4930 & w12589) | (~w5195 & w12589);
assign w5197 = pi1143 & ~w5196;
assign w5198 = pi0589 & ~w4929;
assign w5199 = w3243 & w5198;
assign w5200 = ~w5197 & ~w5199;
assign w5201 = w3242 & ~w4900;
assign w5202 = (~w4901 & w5201) | (~w4901 & w12590) | (w5201 & w12590);
assign w5203 = pi0590 & w5202;
assign w5204 = (pi1143 & w5202) | (pi1143 & w12591) | (w5202 & w12591);
assign w5205 = ~w5203 & w5204;
assign w5206 = pi0591 & ~w4931;
assign w5207 = ~w4932 & ~w5206;
assign w5208 = w3243 & ~w5207;
assign w5209 = (~w4895 & w4902) | (~w4895 & w12592) | (w4902 & w12592);
assign w5210 = w3251 & ~w4903;
assign w5211 = ~w5209 & w5210;
assign w5212 = ~w5208 & ~w5211;
assign w5213 = (pi1459 & w1221) | (pi1459 & w12593) | (w1221 & w12593);
assign w5214 = ~pi0592 & ~w5213;
assign w5215 = w1769 & ~w5214;
assign w5216 = w4058 & w11971;
assign w5217 = ~pi0593 & w4061;
assign w5218 = w2868 & w12594;
assign w5219 = pi1747 & ~w5218;
assign w5220 = w4058 & w12595;
assign w5221 = ~w5217 & w5219;
assign w5222 = ~w5216 & w5221;
assign w5223 = ~w5220 & w5222;
assign w5224 = (w3241 & w12596) | (w3241 & w12597) | (w12596 & w12597);
assign w5225 = (~w3241 & w12598) | (~w3241 & w12599) | (w12598 & w12599);
assign w5226 = pi1143 & ~w5224;
assign w5227 = ~w5225 & w5226;
assign w5228 = w4058 & w12221;
assign w5229 = ~pi0595 & w4061;
assign w5230 = w2868 & w12600;
assign w5231 = pi1747 & ~w5230;
assign w5232 = w4058 & w12601;
assign w5233 = ~w5229 & w5231;
assign w5234 = ~w5228 & w5233;
assign w5235 = ~w5232 & w5234;
assign w5236 = w4058 & w12438;
assign w5237 = ~pi0596 & w4061;
assign w5238 = w2868 & w12602;
assign w5239 = pi1747 & ~w5238;
assign w5240 = w4058 & w12603;
assign w5241 = ~w5237 & w5239;
assign w5242 = ~w5236 & w5241;
assign w5243 = ~w5240 & w5242;
assign w5244 = w4058 & w11974;
assign w5245 = ~pi0597 & w4061;
assign w5246 = w2868 & w12604;
assign w5247 = pi1747 & ~w5246;
assign w5248 = w4058 & w12605;
assign w5249 = ~w5245 & w5247;
assign w5250 = ~w5244 & w5249;
assign w5251 = ~w5248 & w5250;
assign w5252 = w4058 & w11977;
assign w5253 = ~pi0598 & w4061;
assign w5254 = w2868 & w12606;
assign w5255 = pi1747 & ~w5254;
assign w5256 = w4058 & w12607;
assign w5257 = ~w5253 & w5255;
assign w5258 = ~w5252 & w5257;
assign w5259 = ~w5256 & w5258;
assign w5260 = w4058 & w11980;
assign w5261 = ~pi0599 & w4061;
assign w5262 = w2868 & w12608;
assign w5263 = pi1747 & ~w5262;
assign w5264 = w4058 & w12609;
assign w5265 = ~w5261 & w5263;
assign w5266 = ~w5260 & w5265;
assign w5267 = ~w5264 & w5266;
assign w5268 = w4058 & w11983;
assign w5269 = ~pi0600 & w4061;
assign w5270 = w2868 & w12610;
assign w5271 = pi1747 & ~w5270;
assign w5272 = w4058 & w12611;
assign w5273 = ~w5269 & w5271;
assign w5274 = ~w5268 & w5273;
assign w5275 = ~w5272 & w5274;
assign w5276 = w4058 & w12275;
assign w5277 = ~pi0601 & w4061;
assign w5278 = w2868 & w12612;
assign w5279 = pi1747 & ~w5278;
assign w5280 = w4058 & w12613;
assign w5281 = ~w5277 & w5279;
assign w5282 = ~w5276 & w5281;
assign w5283 = ~w5280 & w5282;
assign w5284 = w4058 & w11989;
assign w5285 = ~pi0602 & w4061;
assign w5286 = w2868 & w12614;
assign w5287 = pi1747 & ~w5286;
assign w5288 = w4058 & w12615;
assign w5289 = ~w5285 & w5287;
assign w5290 = ~w5284 & w5289;
assign w5291 = ~w5288 & w5290;
assign w5292 = w4058 & w11994;
assign w5293 = ~pi0603 & w4061;
assign w5294 = w2868 & w12616;
assign w5295 = pi1747 & ~w5294;
assign w5296 = w4058 & w12617;
assign w5297 = ~w5293 & w5295;
assign w5298 = ~w5292 & w5297;
assign w5299 = ~w5296 & w5298;
assign w5300 = w4058 & w12270;
assign w5301 = ~pi0604 & w4061;
assign w5302 = w2868 & w12618;
assign w5303 = pi1747 & ~w5302;
assign w5304 = w4058 & w12619;
assign w5305 = ~w5301 & w5303;
assign w5306 = ~w5300 & w5305;
assign w5307 = ~w5304 & w5306;
assign w5308 = w4058 & w11932;
assign w5309 = ~pi0605 & w4061;
assign w5310 = w2868 & w12620;
assign w5311 = pi1747 & ~w5310;
assign w5312 = w4058 & w12621;
assign w5313 = ~w5309 & w5311;
assign w5314 = ~w5308 & w5313;
assign w5315 = ~w5312 & w5314;
assign w5316 = w4058 & w11998;
assign w5317 = ~pi0606 & w4061;
assign w5318 = w2868 & w12622;
assign w5319 = pi1747 & ~w5318;
assign w5320 = w4058 & w12623;
assign w5321 = ~w5317 & w5319;
assign w5322 = ~w5316 & w5321;
assign w5323 = ~w5320 & w5322;
assign w5324 = w4058 & w12261;
assign w5325 = ~pi0607 & w4061;
assign w5326 = w2868 & w12624;
assign w5327 = pi1747 & ~w5326;
assign w5328 = w4058 & w12625;
assign w5329 = ~w5325 & w5327;
assign w5330 = ~w5324 & w5329;
assign w5331 = ~w5328 & w5330;
assign w5332 = w4058 & w12001;
assign w5333 = ~pi0608 & w4061;
assign w5334 = w2868 & w12626;
assign w5335 = pi1747 & ~w5334;
assign w5336 = w4058 & w12627;
assign w5337 = ~w5333 & w5335;
assign w5338 = ~w5332 & w5337;
assign w5339 = ~w5336 & w5338;
assign w5340 = w4058 & w12006;
assign w5341 = ~pi0609 & w4061;
assign w5342 = w2868 & w12628;
assign w5343 = pi1747 & ~w5342;
assign w5344 = w4058 & w12629;
assign w5345 = ~w5341 & w5343;
assign w5346 = ~w5340 & w5345;
assign w5347 = ~w5344 & w5346;
assign w5348 = w4058 & w12007;
assign w5349 = ~pi0610 & w4061;
assign w5350 = w2868 & w12630;
assign w5351 = pi1747 & ~w5350;
assign w5352 = w4058 & w12631;
assign w5353 = ~w5349 & w5351;
assign w5354 = ~w5348 & w5353;
assign w5355 = ~w5352 & w5354;
assign w5356 = w4058 & w11931;
assign w5357 = ~pi0611 & w4061;
assign w5358 = w2868 & w12632;
assign w5359 = pi1747 & ~w5358;
assign w5360 = w4058 & w12633;
assign w5361 = ~w5357 & w5359;
assign w5362 = ~w5356 & w5361;
assign w5363 = ~w5360 & w5362;
assign w5364 = w3152 & w12634;
assign w5365 = ~pi0612 & w3155;
assign w5366 = w2868 & w12635;
assign w5367 = pi1747 & ~w5366;
assign w5368 = w3152 & w11971;
assign w5369 = ~w5365 & w5367;
assign w5370 = ~w5364 & w5369;
assign w5371 = ~w5368 & w5370;
assign w5372 = w3152 & w12636;
assign w5373 = ~pi0613 & w3155;
assign w5374 = w2868 & w12637;
assign w5375 = pi1747 & ~w5374;
assign w5376 = w3152 & w12275;
assign w5377 = ~w5373 & w5375;
assign w5378 = ~w5372 & w5377;
assign w5379 = ~w5376 & w5378;
assign w5380 = w3152 & w12638;
assign w5381 = ~pi0614 & w3155;
assign w5382 = w2868 & w12639;
assign w5383 = pi1747 & ~w5382;
assign w5384 = w3152 & w12438;
assign w5385 = ~w5381 & w5383;
assign w5386 = ~w5380 & w5385;
assign w5387 = ~w5384 & w5386;
assign w5388 = (pi1430 & w1221) | (pi1430 & w12640) | (w1221 & w12640);
assign w5389 = ~pi0615 & ~w5388;
assign w5390 = w1777 & ~w5389;
assign w5391 = w3152 & w12641;
assign w5392 = ~pi0616 & w3155;
assign w5393 = w2868 & w12642;
assign w5394 = pi1747 & ~w5393;
assign w5395 = w3152 & w12443;
assign w5396 = ~w5392 & w5394;
assign w5397 = ~w5391 & w5396;
assign w5398 = ~w5395 & w5397;
assign w5399 = (pi1447 & w1221) | (pi1447 & w12643) | (w1221 & w12643);
assign w5400 = ~pi0617 & ~w5399;
assign w5401 = w1783 & ~w5400;
assign w5402 = ~w3509 & ~w3510;
assign w5403 = ~w3511 & ~w5402;
assign w5404 = w3511 & w5402;
assign w5405 = ~w5403 & ~w5404;
assign w5406 = pi0506 & ~pi1679;
assign w5407 = pi0618 & ~w5406;
assign w5408 = ~pi0618 & w5406;
assign w5409 = ~w5407 & ~w5408;
assign w5410 = ~w4308 & w5409;
assign w5411 = (pi1131 & ~w5405) | (pi1131 & w12644) | (~w5405 & w12644);
assign w5412 = ~w5410 & w5411;
assign w5413 = pi0619 & pi0634;
assign w5414 = ~w19 & ~w25;
assign w5415 = ~w5413 & w5414;
assign w5416 = w22 & w5415;
assign w5417 = pi1747 & ~w5416;
assign w5418 = (~w1510 & w1517) | (~w1510 & w12645) | (w1517 & w12645);
assign w5419 = (w5418 & ~w4842) | (w5418 & w12646) | (~w4842 & w12646);
assign w5420 = w1528 & ~w5419;
assign w5421 = pi0645 & w3246;
assign w5422 = w3241 & w12647;
assign w5423 = (~w3238 & w12648) | (~w3238 & w12649) | (w12648 & w12649);
assign w5424 = pi0621 & pi1143;
assign w5425 = ~w5423 & w12650;
assign w5426 = ~pi0621 & pi1143;
assign w5427 = (w5426 & w5423) | (w5426 & w12651) | (w5423 & w12651);
assign w5428 = ~w5425 & ~w5427;
assign w5429 = ~w3516 & ~w3517;
assign w5430 = (w5057 & w5429) | (w5057 & w12652) | (w5429 & w12652);
assign w5431 = w4414 & w5429;
assign w5432 = (~pi0622 & ~w3495) | (~pi0622 & w12653) | (~w3495 & w12653);
assign w5433 = ~w5431 & w5432;
assign w5434 = ~w5430 & ~w5433;
assign w5435 = (~pi0623 & ~w3203) | (~pi0623 & w12654) | (~w3203 & w12654);
assign w5436 = ~w3206 & w3243;
assign w5437 = ~w5435 & w5436;
assign w5438 = (~w3238 & w12655) | (~w3238 & w12656) | (w12655 & w12656);
assign w5439 = ~w3240 & w3251;
assign w5440 = ~w5438 & w5439;
assign w5441 = ~w5437 & ~w5440;
assign w5442 = w3952 & w12029;
assign w5443 = w2868 & w12657;
assign w5444 = pi1480 & ~w2934;
assign w5445 = (~w5444 & ~w2868) | (~w5444 & w12658) | (~w2868 & w12658);
assign w5446 = ~pi0624 & w5445;
assign w5447 = (w5444 & ~w2868) | (w5444 & w12659) | (~w2868 & w12659);
assign w5448 = pi0030 & w5447;
assign w5449 = pi1747 & ~w5443;
assign w5450 = ~w5446 & w5449;
assign w5451 = ~w5448 & w5450;
assign w5452 = pi0982 & pi1236;
assign w5453 = ~pi0982 & ~pi1236;
assign w5454 = ~w5452 & ~w5453;
assign w5455 = pi1227 & pi1228;
assign w5456 = pi1016 & pi1229;
assign w5457 = ~pi1016 & ~pi1229;
assign w5458 = ~w5456 & ~w5457;
assign w5459 = ~w5454 & w5455;
assign w5460 = ~w5458 & w5459;
assign w5461 = w3955 & w12660;
assign w5462 = ~pi0626 & w3958;
assign w5463 = w2868 & w12661;
assign w5464 = pi1747 & ~w5463;
assign w5465 = w3955 & w12261;
assign w5466 = ~w5462 & w5464;
assign w5467 = ~w5461 & w5466;
assign w5468 = ~w5465 & w5467;
assign w5469 = (~w4903 & w12662) | (~w4903 & w12663) | (w12662 & w12663);
assign w5470 = ~w4905 & w5469;
assign w5471 = ~w5470 & w12664;
assign w5472 = (pi0627 & w5470) | (pi0627 & w12665) | (w5470 & w12665);
assign w5473 = pi1143 & ~w5471;
assign w5474 = ~w5472 & w5473;
assign w5475 = w2868 & w12666;
assign w5476 = ~pi0628 & w5445;
assign w5477 = pi0028 & w5447;
assign w5478 = pi1747 & ~w5475;
assign w5479 = ~w5476 & w5478;
assign w5480 = ~w5477 & w5479;
assign w5481 = w3955 & w12667;
assign w5482 = ~pi0629 & w3958;
assign w5483 = w2868 & w12668;
assign w5484 = pi1747 & ~w5483;
assign w5485 = w3955 & w11998;
assign w5486 = ~w5482 & w5484;
assign w5487 = ~w5481 & w5486;
assign w5488 = ~w5485 & w5487;
assign w5489 = pi1401 & w25;
assign w5490 = w21 & w5489;
assign w5491 = (~w5490 & ~w17) | (~w5490 & w12670) | (~w17 & w12670);
assign w5492 = w3242 & ~w4917;
assign w5493 = (~w4935 & ~w5492) | (~w4935 & w12671) | (~w5492 & w12671);
assign w5494 = pi0631 & pi1143;
assign w5495 = w5493 & w5494;
assign w5496 = ~pi0631 & pi1143;
assign w5497 = ~w5493 & w5496;
assign w5498 = ~w5495 & ~w5497;
assign w5499 = w3955 & w12310;
assign w5500 = ~pi0632 & w3958;
assign w5501 = w2868 & w12672;
assign w5502 = pi1747 & ~w5501;
assign w5503 = w3955 & w12673;
assign w5504 = ~w5500 & w5502;
assign w5505 = ~w5499 & w5504;
assign w5506 = ~w5503 & w5505;
assign w5507 = w2868 & w12674;
assign w5508 = pi0023 & w5447;
assign w5509 = ~pi0633 & w5445;
assign w5510 = pi1747 & ~w5507;
assign w5511 = ~w5508 & w5510;
assign w5512 = ~w5509 & w5511;
assign w5513 = pi0677 & pi1747;
assign w5514 = w20 & w5513;
assign w5515 = w26 & w5514;
assign w5516 = w2868 & w12675;
assign w5517 = pi0011 & w5447;
assign w5518 = ~pi0635 & w5445;
assign w5519 = pi1747 & ~w5516;
assign w5520 = ~w5517 & w5519;
assign w5521 = ~w5518 & w5520;
assign w5522 = w2868 & w12676;
assign w5523 = ~pi0636 & w5445;
assign w5524 = pi0016 & w5447;
assign w5525 = pi1747 & ~w5522;
assign w5526 = ~w5523 & w5525;
assign w5527 = ~w5524 & w5526;
assign w5528 = w2868 & w12677;
assign w5529 = ~pi0637 & w5445;
assign w5530 = pi0007 & w5447;
assign w5531 = pi1747 & ~w5528;
assign w5532 = ~w5529 & w5531;
assign w5533 = ~w5530 & w5532;
assign w5534 = w2868 & w12678;
assign w5535 = pi0019 & w5447;
assign w5536 = ~pi0638 & w5445;
assign w5537 = pi1747 & ~w5534;
assign w5538 = ~w5535 & w5537;
assign w5539 = ~w5536 & w5538;
assign w5540 = w2868 & w12679;
assign w5541 = ~pi0639 & w5445;
assign w5542 = pi0018 & w5447;
assign w5543 = pi1747 & ~w5540;
assign w5544 = ~w5541 & w5543;
assign w5545 = ~w5542 & w5544;
assign w5546 = w3955 & w12289;
assign w5547 = ~pi0640 & w3958;
assign w5548 = w2868 & w12680;
assign w5549 = pi1747 & ~w5548;
assign w5550 = w3955 & w12681;
assign w5551 = ~w5547 & w5549;
assign w5552 = ~w5546 & w5551;
assign w5553 = ~w5550 & w5552;
assign w5554 = w2868 & w12682;
assign w5555 = pi0046 & w5447;
assign w5556 = ~pi0641 & w5445;
assign w5557 = pi1747 & ~w5554;
assign w5558 = ~w5555 & w5557;
assign w5559 = ~w5556 & w5558;
assign w5560 = w3242 & ~w4920;
assign w5561 = (w5560 & w4918) | (w5560 & w12683) | (w4918 & w12683);
assign w5562 = w3242 & w4925;
assign w5563 = (pi0642 & ~w4934) | (pi0642 & w12684) | (~w4934 & w12684);
assign w5564 = ~w3242 & ~w4936;
assign w5565 = (pi1143 & ~w5564) | (pi1143 & w12685) | (~w5564 & w12685);
assign w5566 = ~w5561 & w5565;
assign w5567 = ~w5562 & w5566;
assign w5568 = ~pi0886 & ~pi1773;
assign w5569 = pi1773 & ~pi1809;
assign w5570 = ~w5568 & ~w5569;
assign w5571 = ~pi0644 & pi0893;
assign w5572 = w1885 & ~w5571;
assign w5573 = (w3243 & ~w3246) | (w3243 & w12686) | (~w3246 & w12686);
assign w5574 = pi1143 & pi1697;
assign w5575 = (w3238 & w12687) | (w3238 & w12688) | (w12687 & w12688);
assign w5576 = ~pi0645 & ~w3246;
assign w5577 = (~w5576 & w5575) | (~w5576 & w12689) | (w5575 & w12689);
assign w5578 = ~pi0645 & w3250;
assign w5579 = w3250 & w12690;
assign w5580 = ~w5577 & ~w5579;
assign w5581 = (pi1747 & ~w17) | (pi1747 & w12691) | (~w17 & w12691);
assign w5582 = w34 & w5581;
assign w5583 = ~w1231 & ~w5455;
assign w5584 = w3560 & ~w5583;
assign w5585 = ~w3572 & w5584;
assign w5586 = (~w1231 & ~w5584) | (~w1231 & w12692) | (~w5584 & w12692);
assign w5587 = w3577 & ~w5586;
assign w5588 = ~w3218 & w3235;
assign w5589 = ~w3236 & ~w5588;
assign w5590 = w3251 & ~w5589;
assign w5591 = (~pi0648 & ~w3200) | (~pi0648 & w12693) | (~w3200 & w12693);
assign w5592 = ~w3203 & w3243;
assign w5593 = ~w5591 & w5592;
assign w5594 = ~w5590 & ~w5593;
assign w5595 = pi0649 & w4937;
assign w5596 = ~w5019 & ~w5595;
assign w5597 = (~w4892 & ~w4937) | (~w4892 & w12694) | (~w4937 & w12694);
assign w5598 = (~w5596 & w4925) | (~w5596 & w12695) | (w4925 & w12695);
assign w5599 = ~pi0649 & ~w4937;
assign w5600 = (~w4937 & w12697) | (~w4937 & w12698) | (w12697 & w12698);
assign w5601 = ~w4925 & w5600;
assign w5602 = (pi1143 & ~w5599) | (pi1143 & w12699) | (~w5599 & w12699);
assign w5603 = ~w5601 & w5602;
assign w5604 = ~w5598 & w5603;
assign w5605 = ~w3233 & w12700;
assign w5606 = ~w3234 & ~w5605;
assign w5607 = w3251 & ~w5606;
assign w5608 = (~pi0650 & ~w3200) | (~pi0650 & w12701) | (~w3200 & w12701);
assign w5609 = ~w3202 & w3243;
assign w5610 = ~w5608 & w5609;
assign w5611 = ~w5607 & ~w5610;
assign w5612 = w2868 & w12702;
assign w5613 = ~pi0651 & w5445;
assign w5614 = ~pi1672 & w5447;
assign w5615 = pi1747 & ~w5612;
assign w5616 = ~w5613 & w5615;
assign w5617 = ~w5614 & w5616;
assign w5618 = w2868 & w12703;
assign w5619 = ~pi0652 & w5445;
assign w5620 = ~pi1666 & w5447;
assign w5621 = pi1747 & ~w5618;
assign w5622 = ~w5619 & w5621;
assign w5623 = ~w5620 & w5622;
assign w5624 = ~w3225 & ~w3226;
assign w5625 = w3231 & ~w5624;
assign w5626 = ~w3231 & w5624;
assign w5627 = ~w5625 & ~w5626;
assign w5628 = w3251 & w5627;
assign w5629 = (~pi0653 & ~w3198) | (~pi0653 & w12704) | (~w3198 & w12704);
assign w5630 = ~w3200 & ~w5629;
assign w5631 = w3243 & w5630;
assign w5632 = ~w5628 & ~w5631;
assign w5633 = (~w3224 & w3232) | (~w3224 & w12705) | (w3232 & w12705);
assign w5634 = ~w3233 & ~w5633;
assign w5635 = w3251 & ~w5634;
assign w5636 = ~pi0654 & ~w3200;
assign w5637 = ~w3201 & ~w5636;
assign w5638 = w3243 & w5637;
assign w5639 = ~w5635 & ~w5638;
assign w5640 = w3242 & ~w4907;
assign w5641 = (~w4933 & ~w5640) | (~w4933 & w12706) | (~w5640 & w12706);
assign w5642 = pi0655 & ~w5641;
assign w5643 = (pi1143 & ~w5641) | (pi1143 & w12707) | (~w5641 & w12707);
assign w5644 = ~w5642 & w5643;
assign w5645 = w3955 & w11986;
assign w5646 = ~pi0656 & w3958;
assign w5647 = w2868 & w12708;
assign w5648 = pi1747 & ~w5647;
assign w5649 = w3955 & w12709;
assign w5650 = ~w5646 & w5648;
assign w5651 = ~w5645 & w5650;
assign w5652 = ~w5649 & w5651;
assign w5653 = w3955 & w11989;
assign w5654 = ~pi0657 & w3958;
assign w5655 = w2868 & w12710;
assign w5656 = pi1747 & ~w5655;
assign w5657 = w3955 & w12711;
assign w5658 = ~w5654 & w5656;
assign w5659 = ~w5653 & w5658;
assign w5660 = ~w5657 & w5659;
assign w5661 = w3955 & w11932;
assign w5662 = ~pi0658 & w3958;
assign w5663 = w2868 & w12712;
assign w5664 = pi1747 & ~w5663;
assign w5665 = w3955 & w12713;
assign w5666 = ~w5662 & w5664;
assign w5667 = ~w5661 & w5666;
assign w5668 = ~w5665 & w5667;
assign w5669 = w3955 & w11931;
assign w5670 = ~pi0659 & w3958;
assign w5671 = w2868 & w12714;
assign w5672 = pi1747 & ~w5671;
assign w5673 = w3955 & w12715;
assign w5674 = ~w5670 & w5672;
assign w5675 = ~w5669 & w5674;
assign w5676 = ~w5673 & w5675;
assign w5677 = w2550 & w12716;
assign w5678 = w7 & w12717;
assign w5679 = ~w5677 & ~w5678;
assign w5680 = w1755 & ~w5679;
assign w5681 = ~pi0883 & ~pi1773;
assign w5682 = pi1773 & ~pi1806;
assign w5683 = ~w5681 & ~w5682;
assign w5684 = ~w3227 & ~w3228;
assign w5685 = ~w3229 & w5684;
assign w5686 = w3229 & ~w5684;
assign w5687 = ~w5685 & ~w5686;
assign w5688 = w3251 & w5687;
assign w5689 = ~pi0662 & ~w3198;
assign w5690 = ~w3199 & ~w5689;
assign w5691 = w3243 & w5690;
assign w5692 = ~w5688 & ~w5691;
assign w5693 = pi1102 & w3291;
assign w5694 = ~pi0698 & ~pi1338;
assign w5695 = pi0698 & pi1338;
assign w5696 = pi0700 & pi1105;
assign w5697 = ~w5695 & ~w5696;
assign w5698 = (~pi1106 & w5697) | (~pi1106 & w12718) | (w5697 & w12718);
assign w5699 = ~w5697 & w12719;
assign w5700 = ~pi0699 & ~w5699;
assign w5701 = ~w5700 & w12720;
assign w5702 = ~pi0669 & ~w5701;
assign w5703 = (~pi1107 & w5700) | (~pi1107 & w12721) | (w5700 & w12721);
assign w5704 = pi1108 & ~w5703;
assign w5705 = ~w5702 & w5704;
assign w5706 = ~pi0710 & ~w5705;
assign w5707 = pi0669 & ~w5703;
assign w5708 = ~pi1108 & ~w5701;
assign w5709 = ~w5707 & w5708;
assign w5710 = pi1081 & ~w5709;
assign w5711 = ~w5706 & w5710;
assign w5712 = ~pi0707 & ~w5711;
assign w5713 = ~pi1081 & w5709;
assign w5714 = ~pi0710 & ~pi1081;
assign w5715 = ~w5705 & w5714;
assign w5716 = ~w5713 & ~w5715;
assign w5717 = pi1109 & w5716;
assign w5718 = ~w5712 & w5717;
assign w5719 = ~pi0679 & ~pi1110;
assign w5720 = ~w5718 & w5719;
assign w5721 = pi0707 & w5716;
assign w5722 = ~pi1109 & ~pi1110;
assign w5723 = ~w5711 & w5722;
assign w5724 = ~w5721 & w5723;
assign w5725 = w3291 & ~w5724;
assign w5726 = ~w5720 & w5725;
assign w5727 = ~w5693 & ~w5726;
assign w5728 = ~pi0679 & ~w5718;
assign w5729 = ~pi1109 & ~w5711;
assign w5730 = ~w5721 & w5729;
assign w5731 = pi1110 & ~w5730;
assign w5732 = ~w5728 & w5731;
assign w5733 = (~pi0720 & ~w3291) | (~pi0720 & w12722) | (~w3291 & w12722);
assign w5734 = ~w5732 & w5733;
assign w5735 = ~w5727 & ~w5734;
assign w5736 = ~pi0709 & ~pi0720;
assign w5737 = ~w5732 & w5736;
assign w5738 = pi1102 & ~w5724;
assign w5739 = ~w5720 & w5738;
assign w5740 = ~pi0709 & ~w5739;
assign w5741 = ~w5737 & ~w5740;
assign w5742 = w5735 & w5741;
assign w5743 = ~pi0698 & ~pi0700;
assign w5744 = ~pi0669 & ~pi0699;
assign w5745 = ~pi0710 & w5744;
assign w5746 = ~pi0679 & ~pi0707;
assign w5747 = w5745 & w5746;
assign w5748 = w5745 & w12723;
assign w5749 = w5748 & w5736;
assign w5750 = ~pi0663 & pi1111;
assign w5751 = (w5748 & w12725) | (w5748 & w12726) | (w12725 & w12726);
assign w5752 = (w5751 & w5742) | (w5751 & w12993) | (w5742 & w12993);
assign w5753 = pi0663 & w3294;
assign w5754 = pi0663 & w3254;
assign w5755 = (w5754 & ~w5748) | (w5754 & w12727) | (~w5748 & w12727);
assign w5756 = (~w5755 & w5742) | (~w5755 & w12728) | (w5742 & w12728);
assign w5757 = ~w5752 & w5756;
assign w5758 = ~pi0359 & w3291;
assign w5759 = (w5758 & w3287) | (w5758 & w12729) | (w3287 & w12729);
assign w5760 = ~w3289 & w5759;
assign w5761 = pi0664 & pi1699;
assign w5762 = ~w5760 & w5761;
assign w5763 = pi1699 & w3291;
assign w5764 = ~pi0359 & ~pi0664;
assign w5765 = w3291 & w12730;
assign w5766 = (w5765 & w3287) | (w5765 & w12731) | (w3287 & w12731);
assign w5767 = ~w3289 & w5766;
assign w5768 = w3299 & w12732;
assign w5769 = pi0664 & w5768;
assign w5770 = (~pi1699 & w5768) | (~pi1699 & w12733) | (w5768 & w12733);
assign w5771 = ~w5769 & w5770;
assign w5772 = ~w5767 & ~w5771;
assign w5773 = ~w5762 & w5772;
assign w5774 = pi1111 & ~w5773;
assign w5775 = w5768 & w12733;
assign w5776 = pi0665 & pi1111;
assign w5777 = ~w5767 & w12734;
assign w5778 = ~pi0665 & pi1111;
assign w5779 = (w5778 & w5767) | (w5778 & w12735) | (w5767 & w12735);
assign w5780 = ~w5777 & ~w5779;
assign w5781 = ~pi0885 & ~pi1773;
assign w5782 = pi1773 & ~pi1808;
assign w5783 = ~w5781 & ~w5782;
assign w5784 = w2868 & w12736;
assign w5785 = pi0154 & w5447;
assign w5786 = ~pi0667 & w5445;
assign w5787 = pi1747 & ~w5784;
assign w5788 = ~w5785 & w5787;
assign w5789 = ~w5786 & w5788;
assign w5790 = w2868 & w12737;
assign w5791 = ~pi0668 & w5445;
assign w5792 = pi0286 & w5447;
assign w5793 = pi1747 & ~w5790;
assign w5794 = ~w5791 & w5793;
assign w5795 = ~w5792 & w5794;
assign w5796 = ~w5701 & w5763;
assign w5797 = ~w5703 & w5796;
assign w5798 = w5796 & w12738;
assign w5799 = ~pi1699 & w5743;
assign w5800 = w5744 & w5799;
assign w5801 = ~pi0699 & ~w3294;
assign w5802 = (pi0669 & ~w5801) | (pi0669 & w12739) | (~w5801 & w12739);
assign w5803 = ~w5797 & w5802;
assign w5804 = ~w5798 & ~w5800;
assign w5805 = ~w5803 & w5804;
assign w5806 = pi1111 & ~w5805;
assign w5807 = w2868 & w12740;
assign w5808 = pi0064 & w5447;
assign w5809 = ~pi0670 & w5445;
assign w5810 = pi1747 & ~w5807;
assign w5811 = ~w5808 & w5810;
assign w5812 = ~w5809 & w5811;
assign w5813 = w2868 & w12741;
assign w5814 = pi0310 & w5447;
assign w5815 = ~pi0671 & w5445;
assign w5816 = pi1747 & ~w5813;
assign w5817 = ~w5814 & w5816;
assign w5818 = ~w5815 & w5817;
assign w5819 = pi0759 & ~pi0848;
assign w5820 = ~pi0849 & pi0877;
assign w5821 = pi0748 & ~pi0810;
assign w5822 = ~pi0759 & pi0848;
assign w5823 = pi0809 & ~pi0847;
assign w5824 = ~pi0748 & pi0810;
assign w5825 = ~pi0808 & pi0846;
assign w5826 = ~pi0809 & pi0847;
assign w5827 = pi0808 & ~pi0846;
assign w5828 = pi0755 & ~pi0845;
assign w5829 = ~pi0755 & pi0845;
assign w5830 = pi0751 & ~pi0807;
assign w5831 = ~pi0751 & pi0807;
assign w5832 = pi0806 & ~pi0844;
assign w5833 = ~pi0806 & pi0844;
assign w5834 = ~pi0804 & pi0842;
assign w5835 = pi0750 & ~pi0754;
assign w5836 = pi0804 & ~pi0842;
assign w5837 = ~pi0750 & pi0754;
assign w5838 = ~pi0841 & pi0859;
assign w5839 = ~w5837 & w5838;
assign w5840 = ~w5835 & ~w5836;
assign w5841 = ~w5839 & w5840;
assign w5842 = ~w5833 & ~w5834;
assign w5843 = ~w5831 & ~w5832;
assign w5844 = (w5843 & w5841) | (w5843 & w12742) | (w5841 & w12742);
assign w5845 = ~w5829 & ~w5830;
assign w5846 = ~w5827 & ~w5828;
assign w5847 = ~w5825 & ~w5826;
assign w5848 = (~w5844 & w12744) | (~w5844 & w12745) | (w12744 & w12745);
assign w5849 = ~w5823 & ~w5824;
assign w5850 = ~w5821 & ~w5822;
assign w5851 = ~w5819 & ~w5820;
assign w5852 = (~w5848 & w12747) | (~w5848 & w12748) | (w12747 & w12748);
assign w5853 = pi0849 & ~pi0877;
assign w5854 = ~pi0749 & ~pi0850;
assign w5855 = ~pi0852 & w5854;
assign w5856 = ~w5853 & w5855;
assign w5857 = ~w5852 & w5856;
assign w5858 = w1516 & ~w1522;
assign w5859 = ~w1523 & ~w5858;
assign w5860 = pi0663 & pi0715;
assign w5861 = ~pi0674 & w3294;
assign w5862 = w5860 & w5861;
assign w5863 = ~pi0663 & w5736;
assign w5864 = w5747 & w5863;
assign w5865 = w5747 & w12749;
assign w5866 = ~pi0674 & w5865;
assign w5867 = w3254 & w5743;
assign w5868 = w5865 & w12750;
assign w5869 = pi1699 & w5860;
assign w5870 = pi0674 & pi1111;
assign w5871 = (w5870 & ~w5865) | (w5870 & w12751) | (~w5865 & w12751);
assign w5872 = (w5871 & ~w5742) | (w5871 & w12752) | (~w5742 & w12752);
assign w5873 = (~w5868 & ~w5742) | (~w5868 & w12753) | (~w5742 & w12753);
assign w5874 = ~w5872 & w5873;
assign w5875 = w3297 & w12754;
assign w5876 = pi0678 & w5875;
assign w5877 = (pi1111 & ~w3291) | (pi1111 & w3254) | (~w3291 & w3254);
assign w5878 = ~w5876 & w5877;
assign w5879 = ~w3283 & ~w3285;
assign w5880 = (pi0675 & w5876) | (pi0675 & w12755) | (w5876 & w12755);
assign w5881 = (w5880 & w5879) | (w5880 & w12756) | (w5879 & w12756);
assign w5882 = w3291 & w3294;
assign w5883 = (~pi0675 & ~w5875) | (~pi0675 & w12758) | (~w5875 & w12758);
assign w5884 = (w5883 & ~w5879) | (w5883 & w12759) | (~w5879 & w12759);
assign w5885 = ~w5881 & ~w5884;
assign w5886 = ~pi0387 & pi1175;
assign w5887 = ~pi0386 & pi1089;
assign w5888 = pi0387 & ~pi1175;
assign w5889 = pi0480 & ~pi1093;
assign w5890 = ~pi0480 & pi1093;
assign w5891 = ~pi0484 & pi1174;
assign w5892 = pi0484 & ~pi1174;
assign w5893 = pi0509 & ~pi1087;
assign w5894 = ~pi0509 & pi1087;
assign w5895 = ~pi0508 & pi1173;
assign w5896 = pi0508 & ~pi1173;
assign w5897 = ~pi0507 & pi1077;
assign w5898 = pi0507 & ~pi1077;
assign w5899 = ~pi0408 & pi1241;
assign w5900 = ~w5898 & w5899;
assign w5901 = (~w5896 & w5900) | (~w5896 & w12760) | (w5900 & w12760);
assign w5902 = ~w5894 & ~w5895;
assign w5903 = ~w5892 & ~w5893;
assign w5904 = (w5903 & w5901) | (w5903 & w12761) | (w5901 & w12761);
assign w5905 = ~w5890 & ~w5891;
assign w5906 = ~w5888 & ~w5889;
assign w5907 = ~w5886 & ~w5887;
assign w5908 = (~w5904 & w12763) | (~w5904 & w12764) | (w12763 & w12764);
assign w5909 = pi0466 & ~pi1176;
assign w5910 = pi0386 & ~pi1089;
assign w5911 = ~w5909 & ~w5910;
assign w5912 = ~pi0466 & pi1176;
assign w5913 = ~pi0379 & pi1082;
assign w5914 = ~w5912 & ~w5913;
assign w5915 = pi0470 & ~pi1177;
assign w5916 = pi0379 & ~pi1082;
assign w5917 = ~w5915 & ~w5916;
assign w5918 = ~pi0470 & pi1177;
assign w5919 = ~pi0381 & pi1179;
assign w5920 = ~w5918 & ~w5919;
assign w5921 = (w5908 & w12768) | (w5908 & w12769) | (w12768 & w12769);
assign w5922 = pi1256 & ~pi1257;
assign w5923 = pi0381 & ~pi1179;
assign w5924 = w5922 & ~w5923;
assign w5925 = ~pi0383 & ~pi0441;
assign w5926 = w3645 & w5925;
assign w5927 = w3630 & w5926;
assign w5928 = w3630 & w12770;
assign w5929 = w1501 & ~w5928;
assign w5930 = (~w5929 & w5921) | (~w5929 & w12771) | (w5921 & w12771);
assign w5931 = ~pi1607 & ~pi1734;
assign w5932 = w3675 & w5931;
assign w5933 = ~w5930 & w5932;
assign w5934 = ~w21 & ~w27;
assign w5935 = pi1747 & ~w5934;
assign w5936 = ~w5491 & w5935;
assign w5937 = ~pi0678 & ~w5875;
assign w5938 = w5878 & ~w5937;
assign w5939 = (~w3276 & w3274) | (~w3276 & w12772) | (w3274 & w12772);
assign w5940 = ~w3282 & w5882;
assign w5941 = ~w5939 & w5940;
assign w5942 = ~w5938 & ~w5941;
assign w5943 = ~w5730 & w5882;
assign w5944 = w5728 & w5943;
assign w5945 = ~w5718 & ~w5730;
assign w5946 = w5799 & w5745;
assign w5947 = ~pi0707 & w5946;
assign w5948 = w5877 & ~w5947;
assign w5949 = (~w5948 & w5945) | (~w5948 & w12773) | (w5945 & w12773);
assign w5950 = pi0679 & ~w5949;
assign w5951 = w3254 & w5748;
assign w5952 = ~w5944 & ~w5951;
assign w5953 = ~w5950 & w5952;
assign w5954 = w2868 & w12774;
assign w5955 = pi0014 & w5447;
assign w5956 = ~pi0680 & w5445;
assign w5957 = pi1747 & ~w5954;
assign w5958 = ~w5955 & w5957;
assign w5959 = ~w5956 & w5958;
assign w5960 = w2868 & w12775;
assign w5961 = ~pi0681 & w5445;
assign w5962 = pi0015 & w5447;
assign w5963 = pi1747 & ~w5960;
assign w5964 = ~w5961 & w5963;
assign w5965 = ~w5962 & w5964;
assign w5966 = w2868 & w12776;
assign w5967 = pi0953 & w5447;
assign w5968 = ~pi0682 & w5445;
assign w5969 = pi1747 & ~w5966;
assign w5970 = ~w5967 & w5969;
assign w5971 = ~w5968 & w5970;
assign w5972 = w2868 & w12777;
assign w5973 = pi0332 & w5447;
assign w5974 = ~pi0683 & w5445;
assign w5975 = pi1747 & ~w5972;
assign w5976 = ~w5973 & w5975;
assign w5977 = ~w5974 & w5976;
assign w5978 = w2868 & w12778;
assign w5979 = pi0057 & w5447;
assign w5980 = ~pi0684 & w5445;
assign w5981 = pi1747 & ~w5978;
assign w5982 = ~w5979 & w5981;
assign w5983 = ~w5980 & w5982;
assign w5984 = w2868 & w12779;
assign w5985 = pi0299 & w5447;
assign w5986 = ~pi0685 & w5445;
assign w5987 = pi1747 & ~w5984;
assign w5988 = ~w5985 & w5987;
assign w5989 = ~w5986 & w5988;
assign w5990 = w2868 & w12780;
assign w5991 = pi1481 & w5447;
assign w5992 = ~pi0686 & w5445;
assign w5993 = pi1747 & ~w5990;
assign w5994 = ~w5991 & w5993;
assign w5995 = ~w5992 & w5994;
assign w5996 = w2868 & w12781;
assign w5997 = ~pi0687 & w5445;
assign w5998 = pi0254 & w5447;
assign w5999 = pi1747 & ~w5996;
assign w6000 = ~w5997 & w5999;
assign w6001 = ~w5998 & w6000;
assign w6002 = w2868 & w12782;
assign w6003 = pi0223 & w5447;
assign w6004 = ~pi0688 & w5445;
assign w6005 = pi1747 & ~w6002;
assign w6006 = ~w6003 & w6005;
assign w6007 = ~w6004 & w6006;
assign w6008 = w2868 & w12783;
assign w6009 = ~pi0689 & w5445;
assign w6010 = pi0124 & w5447;
assign w6011 = pi1747 & ~w6008;
assign w6012 = ~w6009 & w6011;
assign w6013 = ~w6010 & w6012;
assign w6014 = w2868 & w12784;
assign w6015 = ~pi0690 & w5445;
assign w6016 = pi0155 & w5447;
assign w6017 = pi1747 & ~w6014;
assign w6018 = ~w6015 & w6017;
assign w6019 = ~w6016 & w6018;
assign w6020 = w2868 & w12785;
assign w6021 = pi0063 & w5447;
assign w6022 = ~pi0691 & w5445;
assign w6023 = pi1747 & ~w6020;
assign w6024 = ~w6021 & w6023;
assign w6025 = ~w6022 & w6024;
assign w6026 = w2868 & w12786;
assign w6027 = pi0056 & w5447;
assign w6028 = ~pi0692 & w5445;
assign w6029 = pi1747 & ~w6026;
assign w6030 = ~w6027 & w6029;
assign w6031 = ~w6028 & w6030;
assign w6032 = w2868 & w12787;
assign w6033 = ~pi0693 & w5445;
assign w6034 = pi0022 & w5447;
assign w6035 = pi1747 & ~w6032;
assign w6036 = ~w6033 & w6035;
assign w6037 = ~w6034 & w6036;
assign w6038 = w2868 & w12788;
assign w6039 = ~pi0694 & w5445;
assign w6040 = pi0027 & w5447;
assign w6041 = pi1747 & ~w6038;
assign w6042 = ~w6039 & w6041;
assign w6043 = ~w6040 & w6042;
assign w6044 = w3559 & w3569;
assign w6045 = w3569 & w12789;
assign w6046 = pi0695 & w6045;
assign w6047 = (w3564 & w3561) | (w3564 & w12790) | (w3561 & w12790);
assign w6048 = ~w5584 & w6047;
assign w6049 = w3577 & w6048;
assign w6050 = ~w6046 & ~w6049;
assign w6051 = (pi1699 & ~w3291) | (pi1699 & w12791) | (~w3291 & w12791);
assign w6052 = (~w3291 & w12792) | (~w3291 & w12793) | (w12792 & w12793);
assign w6053 = (pi1111 & w6051) | (pi1111 & w12794) | (w6051 & w12794);
assign w6054 = ~w6052 & w6053;
assign w6055 = ~pi0700 & ~pi1699;
assign w6056 = pi0698 & ~w6055;
assign w6057 = w5877 & w6056;
assign w6058 = ~w5694 & ~w5695;
assign w6059 = ~w5696 & ~w6058;
assign w6060 = w5696 & w6058;
assign w6061 = ~w6059 & ~w6060;
assign w6062 = (~w5867 & ~w6061) | (~w5867 & w12795) | (~w6061 & w12795);
assign w6063 = ~w6057 & w6062;
assign w6064 = ~w5698 & ~w5699;
assign w6065 = ~w5799 & w5877;
assign w6066 = (pi0699 & w6064) | (pi0699 & w12796) | (w6064 & w12796);
assign w6067 = ~w6065 & w6066;
assign w6068 = ~pi0699 & ~w5867;
assign w6069 = (w6068 & ~w6064) | (w6068 & w12797) | (~w6064 & w12797);
assign w6070 = ~w6067 & ~w6069;
assign w6071 = (w3291 & w12798) | (w3291 & w12799) | (w12798 & w12799);
assign w6072 = (~w3291 & w12800) | (~w3291 & w12801) | (w12800 & w12801);
assign w6073 = pi1111 & ~w6071;
assign w6074 = ~w6072 & w6073;
assign w6075 = ~pi0997 & w1345;
assign w6076 = ~w1609 & ~w6075;
assign w6077 = (~w17 & w12804) | (~w17 & w12805) | (w12804 & w12805);
assign w6078 = pi1747 & w24;
assign w6079 = w24 & w12806;
assign w6080 = ~w6077 & ~w6079;
assign w6081 = w2868 & w12807;
assign w6082 = pi0049 & w5447;
assign w6083 = ~pi0703 & w5445;
assign w6084 = pi1747 & ~w6081;
assign w6085 = ~w6082 & w6084;
assign w6086 = ~w6083 & w6085;
assign w6087 = w2868 & w12808;
assign w6088 = ~pi0704 & w5445;
assign w6089 = pi0194 & w5447;
assign w6090 = pi1747 & ~w6087;
assign w6091 = ~w6088 & w6090;
assign w6092 = ~w6089 & w6091;
assign w6093 = w5877 & ~w5946;
assign w6094 = ~w5711 & w5716;
assign w6095 = pi0707 & ~w6093;
assign w6096 = (w6095 & w6094) | (w6095 & w12809) | (w6094 & w12809);
assign w6097 = w5745 & w5867;
assign w6098 = ~pi0707 & ~w6097;
assign w6099 = (w6098 & ~w6094) | (w6098 & w12810) | (~w6094 & w12810);
assign w6100 = ~w6096 & ~w6099;
assign w6101 = w3254 & ~w3296;
assign w6102 = (~w3294 & w3296) | (~w3294 & w12811) | (w3296 & w12811);
assign w6103 = pi0708 & ~w6102;
assign w6104 = ~w5882 & ~w6103;
assign w6105 = (~w3258 & w3265) | (~w3258 & w12812) | (w3265 & w12812);
assign w6106 = ~w3266 & w5763;
assign w6107 = (~w6104 & ~w6106) | (~w6104 & w12813) | (~w6106 & w12813);
assign w6108 = ~pi0708 & w3254;
assign w6109 = w3296 & w6108;
assign w6110 = ~w6107 & ~w6109;
assign w6111 = ~pi0720 & ~w5732;
assign w6112 = w5739 & ~w6111;
assign w6113 = w5735 & ~w6112;
assign w6114 = pi0709 & w3294;
assign w6115 = (pi0709 & ~w5748) | (pi0709 & w12814) | (~w5748 & w12814);
assign w6116 = ~w5749 & ~w6115;
assign w6117 = w3254 & ~w6116;
assign w6118 = ~pi0709 & w3294;
assign w6119 = w6113 & w6118;
assign w6120 = (~w6117 & w6113) | (~w6117 & w12815) | (w6113 & w12815);
assign w6121 = ~w6119 & w6120;
assign w6122 = ~w5709 & w5882;
assign w6123 = w5706 & w6122;
assign w6124 = ~w5705 & ~w5709;
assign w6125 = ~w5800 & w5877;
assign w6126 = (~w6125 & w6124) | (~w6125 & w12816) | (w6124 & w12816);
assign w6127 = pi0710 & ~w6126;
assign w6128 = ~w6097 & ~w6123;
assign w6129 = ~w6127 & w6128;
assign w6130 = ~pi0471 & ~pi0472;
assign w6131 = ~pi0513 & ~pi0560;
assign w6132 = ~pi0564 & w6131;
assign w6133 = w4305 & w6130;
assign w6134 = w6132 & w6133;
assign w6135 = w4301 & w6134;
assign w6136 = w6134 & w12817;
assign w6137 = w1405 & ~w6136;
assign w6138 = ~pi0483 & pi1198;
assign w6139 = ~pi0485 & pi1197;
assign w6140 = pi0485 & ~pi1197;
assign w6141 = pi0549 & ~pi1264;
assign w6142 = ~pi0549 & pi1264;
assign w6143 = ~pi0567 & pi1196;
assign w6144 = pi0567 & ~pi1196;
assign w6145 = pi0622 & ~pi1195;
assign w6146 = ~pi0622 & pi1195;
assign w6147 = ~pi0587 & pi1194;
assign w6148 = pi0587 & ~pi1194;
assign w6149 = ~pi0618 & pi1276;
assign w6150 = pi0618 & ~pi1276;
assign w6151 = ~pi0506 & pi1192;
assign w6152 = ~w6150 & w6151;
assign w6153 = (~w6148 & w6152) | (~w6148 & w12818) | (w6152 & w12818);
assign w6154 = ~w6146 & ~w6147;
assign w6155 = ~w6144 & ~w6145;
assign w6156 = (w6155 & w6153) | (w6155 & w12819) | (w6153 & w12819);
assign w6157 = ~w6142 & ~w6143;
assign w6158 = ~w6140 & ~w6141;
assign w6159 = ~w6138 & ~w6139;
assign w6160 = (~w6156 & w12821) | (~w6156 & w12822) | (w12821 & w12822);
assign w6161 = pi0483 & ~pi1198;
assign w6162 = pi0533 & ~pi1199;
assign w6163 = ~w6161 & ~w6162;
assign w6164 = ~pi0380 & pi1249;
assign w6165 = ~pi0533 & pi1199;
assign w6166 = ~w6164 & ~w6165;
assign w6167 = pi0562 & ~pi1201;
assign w6168 = pi0380 & ~pi1249;
assign w6169 = ~w6167 & ~w6168;
assign w6170 = ~pi0468 & pi1036;
assign w6171 = ~pi0562 & pi1201;
assign w6172 = ~w6170 & ~w6171;
assign w6173 = (w6160 & w12826) | (w6160 & w12827) | (w12826 & w12827);
assign w6174 = pi1080 & ~pi1132;
assign w6175 = pi0468 & ~pi1036;
assign w6176 = w6174 & ~w6175;
assign w6177 = (~w6137 & w6173) | (~w6137 & w12828) | (w6173 & w12828);
assign w6178 = ~pi1608 & ~pi1730;
assign w6179 = w3491 & w6178;
assign w6180 = ~w6177 & w6179;
assign w6181 = w5875 & w3300;
assign w6182 = ~w3288 & ~w3290;
assign w6183 = w3294 & ~w6182;
assign w6184 = (pi0712 & w6181) | (pi0712 & w12829) | (w6181 & w12829);
assign w6185 = ~w6183 & w6184;
assign w6186 = w5882 & w6182;
assign w6187 = (~pi0712 & ~w5875) | (~pi0712 & w12831) | (~w5875 & w12831);
assign w6188 = ~w6186 & w6187;
assign w6189 = ~w6185 & ~w6188;
assign w6190 = ~pi0566 & pi1219;
assign w6191 = ~pi0623 & pi1056;
assign w6192 = pi0569 & ~pi1218;
assign w6193 = pi0566 & ~pi1219;
assign w6194 = ~pi0648 & pi1217;
assign w6195 = ~pi0569 & pi1218;
assign w6196 = pi0648 & ~pi1217;
assign w6197 = pi0650 & ~pi1066;
assign w6198 = ~pi0650 & pi1066;
assign w6199 = ~pi0654 & pi1216;
assign w6200 = pi0654 & ~pi1216;
assign w6201 = pi0653 & ~pi1215;
assign w6202 = ~pi0662 & pi1214;
assign w6203 = ~pi0653 & pi1215;
assign w6204 = pi0662 & ~pi1214;
assign w6205 = ~pi0586 & pi1213;
assign w6206 = ~w6204 & w6205;
assign w6207 = ~w6202 & ~w6203;
assign w6208 = ~w6206 & w6207;
assign w6209 = ~w6200 & ~w6201;
assign w6210 = ~w6198 & ~w6199;
assign w6211 = (w6210 & w6208) | (w6210 & w12832) | (w6208 & w12832);
assign w6212 = ~w6196 & ~w6197;
assign w6213 = ~w6194 & ~w6195;
assign w6214 = ~w6192 & ~w6193;
assign w6215 = (~w6211 & w12834) | (~w6211 & w12835) | (w12834 & w12835);
assign w6216 = ~w6190 & ~w6191;
assign w6217 = pi0358 & ~pi1057;
assign w6218 = pi0623 & ~pi1056;
assign w6219 = ~w6217 & ~w6218;
assign w6220 = ~pi0358 & pi1057;
assign w6221 = ~pi0645 & pi1232;
assign w6222 = ~w6220 & ~w6221;
assign w6223 = pi0621 & ~pi1266;
assign w6224 = pi0645 & ~pi1232;
assign w6225 = ~w6223 & ~w6224;
assign w6226 = (w6215 & w12839) | (w6215 & w12840) | (w12839 & w12840);
assign w6227 = ~pi0621 & pi1266;
assign w6228 = ~w1493 & ~w6227;
assign w6229 = ~w6226 & w6228;
assign w6230 = ~pi0589 & ~pi0594;
assign w6231 = w1493 & ~w6230;
assign w6232 = pi1144 & ~pi1259;
assign w6233 = ~pi0552 & ~pi0563;
assign w6234 = ~pi0568 & ~pi0590;
assign w6235 = ~pi0591 & ~pi0627;
assign w6236 = ~pi0631 & ~pi0642;
assign w6237 = ~pi0649 & ~pi0655;
assign w6238 = w6236 & w6237;
assign w6239 = w6234 & w6235;
assign w6240 = w6233 & w6239;
assign w6241 = (w1493 & ~w6240) | (w1493 & w12841) | (~w6240 & w12841);
assign w6242 = ~w6231 & ~w6232;
assign w6243 = ~pi1583 & ~pi1743;
assign w6244 = w5574 & w6243;
assign w6245 = (w6244 & w6241) | (w6244 & w12842) | (w6241 & w12842);
assign w6246 = ~w6229 & w6245;
assign w6247 = (w3291 & w12843) | (w3291 & w12844) | (w12843 & w12844);
assign w6248 = ~w5875 & ~w6247;
assign w6249 = ~w3273 & w3280;
assign w6250 = (~w6248 & w6249) | (~w6248 & w12845) | (w6249 & w12845);
assign w6251 = w5882 & w6249;
assign w6252 = (~pi0714 & ~w3298) | (~pi0714 & w12846) | (~w3298 & w12846);
assign w6253 = ~w6251 & w6252;
assign w6254 = ~w6250 & ~w6253;
assign w6255 = (~pi0715 & ~w5865) | (~pi0715 & w12847) | (~w5865 & w12847);
assign w6256 = pi1111 & ~w6255;
assign w6257 = (~w6256 & ~w5742) | (~w6256 & w12848) | (~w5742 & w12848);
assign w6258 = pi0715 & w5800;
assign w6259 = w5864 & w6258;
assign w6260 = (~w6259 & ~w5742) | (~w6259 & w12849) | (~w5742 & w12849);
assign w6261 = ~w6257 & w6260;
assign w6262 = (~w17 & w12850) | (~w17 & w12851) | (w12850 & w12851);
assign w6263 = ~pi1748 & w6078;
assign w6264 = ~w6262 & ~w6263;
assign w6265 = (w3291 & w3266) | (w3291 & w12852) | (w3266 & w12852);
assign w6266 = ~w3271 & w6265;
assign w6267 = ~pi0717 & ~w6266;
assign w6268 = (w3294 & ~w6266) | (w3294 & w12853) | (~w6266 & w12853);
assign w6269 = ~w6267 & w6268;
assign w6270 = ~pi0717 & ~w3297;
assign w6271 = (w3254 & ~w3297) | (w3254 & w12854) | (~w3297 & w12854);
assign w6272 = ~w6270 & w6271;
assign w6273 = ~w6269 & ~w6272;
assign w6274 = pi0697 & ~pi1699;
assign w6275 = ~pi0718 & ~w6274;
assign w6276 = pi0718 & w6274;
assign w6277 = ~w6275 & ~w6276;
assign w6278 = w5877 & w6277;
assign w6279 = ~w3259 & ~w3260;
assign w6280 = w3261 & ~w6279;
assign w6281 = ~w3261 & w6279;
assign w6282 = ~w6280 & ~w6281;
assign w6283 = w5882 & w6282;
assign w6284 = ~w6278 & ~w6283;
assign w6285 = ~pi0719 & ~w3295;
assign w6286 = w6101 & ~w6285;
assign w6287 = ~w3263 & w3291;
assign w6288 = w6287 & w3265;
assign w6289 = (~pi0719 & ~w6287) | (~pi0719 & w12855) | (~w6287 & w12855);
assign w6290 = w3294 & ~w6288;
assign w6291 = ~w6289 & w6290;
assign w6292 = ~w6286 & ~w6291;
assign w6293 = w5747 & w5799;
assign w6294 = ~w5720 & ~w5724;
assign w6295 = ~w5732 & w6294;
assign w6296 = w3294 & ~w6295;
assign w6297 = (pi0720 & w6293) | (pi0720 & w12856) | (w6293 & w12856);
assign w6298 = ~w6296 & w6297;
assign w6299 = (~pi0720 & ~w5748) | (~pi0720 & w12857) | (~w5748 & w12857);
assign w6300 = (w6299 & ~w6295) | (w6299 & w12858) | (~w6295 & w12858);
assign w6301 = ~w6298 & ~w6300;
assign w6302 = pi0712 & ~pi1346;
assign w6303 = pi0675 & ~pi1158;
assign w6304 = ~pi0675 & pi1158;
assign w6305 = ~pi0678 & pi1275;
assign w6306 = pi0678 & ~pi1275;
assign w6307 = pi0714 & ~pi1157;
assign w6308 = ~pi0714 & pi1157;
assign w6309 = ~pi0717 & pi1156;
assign w6310 = pi0717 & ~pi1156;
assign w6311 = pi0708 & ~pi1155;
assign w6312 = ~pi0708 & pi1155;
assign w6313 = ~pi0719 & pi1154;
assign w6314 = pi0718 & ~pi1283;
assign w6315 = ~pi0718 & pi1283;
assign w6316 = ~pi0697 & pi1331;
assign w6317 = ~w6315 & ~w6316;
assign w6318 = pi0719 & ~pi1154;
assign w6319 = ~w6314 & ~w6318;
assign w6320 = ~w6317 & w6319;
assign w6321 = ~w6312 & ~w6313;
assign w6322 = ~w6310 & ~w6311;
assign w6323 = (w6322 & w6320) | (w6322 & w12859) | (w6320 & w12859);
assign w6324 = ~w6308 & ~w6309;
assign w6325 = ~w6306 & ~w6307;
assign w6326 = ~w6304 & ~w6305;
assign w6327 = (~w6323 & w12861) | (~w6323 & w12862) | (w12861 & w12862);
assign w6328 = ~w6302 & ~w6303;
assign w6329 = ~pi0359 & pi1159;
assign w6330 = ~pi0712 & pi1346;
assign w6331 = ~w6329 & ~w6330;
assign w6332 = pi0359 & ~pi1159;
assign w6333 = pi0664 & ~pi1269;
assign w6334 = ~w6332 & ~w6333;
assign w6335 = ~pi0665 & pi1160;
assign w6336 = ~pi0664 & pi1269;
assign w6337 = ~w6335 & ~w6336;
assign w6338 = (w6327 & w12866) | (w6327 & w12867) | (w12866 & w12867);
assign w6339 = pi1112 & ~pi1113;
assign w6340 = pi0665 & ~pi1160;
assign w6341 = w6339 & ~w6340;
assign w6342 = ~w6338 & w6341;
assign w6343 = (w1586 & ~w5865) | (w1586 & w12869) | (~w5865 & w12869);
assign w6344 = ~w6342 & ~w6343;
assign w6345 = ~pi1604 & ~pi1728;
assign w6346 = w3294 & w6345;
assign w6347 = ~w6344 & w6346;
assign w6348 = (pi0722 & ~w5584) | (pi0722 & w12870) | (~w5584 & w12870);
assign w6349 = w5584 & w12871;
assign w6350 = ~pi0732 & ~pi1741;
assign w6351 = pi0732 & pi1741;
assign w6352 = ~w6350 & ~w6351;
assign w6353 = ~pi0744 & ~pi1722;
assign w6354 = pi0744 & pi1722;
assign w6355 = ~w6353 & ~w6354;
assign w6356 = w6352 & ~w6355;
assign w6357 = ~w6352 & w6355;
assign w6358 = ~w6356 & ~w6357;
assign w6359 = ~pi0727 & ~pi1733;
assign w6360 = pi0727 & pi1733;
assign w6361 = ~w6359 & ~w6360;
assign w6362 = w6358 & ~w6361;
assign w6363 = ~w6358 & w6361;
assign w6364 = ~w6362 & ~w6363;
assign w6365 = ~pi0730 & ~pi1735;
assign w6366 = pi0730 & pi1735;
assign w6367 = ~w6365 & ~w6366;
assign w6368 = pi0738 & ~w6367;
assign w6369 = ~pi0738 & w6367;
assign w6370 = ~w6368 & ~w6369;
assign w6371 = ~pi0723 & ~pi1740;
assign w6372 = pi0723 & pi1740;
assign w6373 = ~w6371 & ~w6372;
assign w6374 = ~pi0731 & ~pi1727;
assign w6375 = pi0731 & pi1727;
assign w6376 = ~w6374 & ~w6375;
assign w6377 = w6373 & ~w6376;
assign w6378 = ~w6373 & w6376;
assign w6379 = ~w6377 & ~w6378;
assign w6380 = w6370 & ~w6379;
assign w6381 = ~w6370 & w6379;
assign w6382 = ~w6380 & ~w6381;
assign w6383 = w6364 & w6382;
assign w6384 = ~w6364 & ~w6382;
assign w6385 = ~w6383 & ~w6384;
assign w6386 = w5584 & w12872;
assign w6387 = ~w6385 & w6386;
assign w6388 = pi1496 & ~pi1626;
assign w6389 = ~w6348 & ~w6388;
assign w6390 = (w6389 & ~w6385) | (w6389 & w12873) | (~w6385 & w12873);
assign w6391 = ~w6387 & w6390;
assign w6392 = w5584 & w12874;
assign w6393 = (pi0723 & ~w5584) | (pi0723 & w12875) | (~w5584 & w12875);
assign w6394 = ~w6388 & ~w6392;
assign w6395 = ~w6393 & w6394;
assign w6396 = pi1737 & pi1739;
assign w6397 = ~pi1668 & w6396;
assign w6398 = w2152 & w6397;
assign w6399 = pi0785 & ~pi1479;
assign w6400 = w2154 & w6399;
assign w6401 = ~w2156 & w6400;
assign w6402 = ~w6398 & ~w6401;
assign w6403 = w2150 & ~w6402;
assign w6404 = w2137 & w12876;
assign w6405 = w2167 & w6404;
assign w6406 = ~w6403 & ~w6405;
assign w6407 = ~pi0765 & pi0766;
assign w6408 = pi0761 & pi0787;
assign w6409 = ~pi0788 & ~w6408;
assign w6410 = (pi0783 & w6408) | (pi0783 & w12877) | (w6408 & w12877);
assign w6411 = pi0764 & pi0790;
assign w6412 = w6407 & w6411;
assign w6413 = ~w6410 & w6412;
assign w6414 = w6406 & ~w6413;
assign w6415 = ~pi0236 & pi0877;
assign w6416 = pi0243 & ~pi0759;
assign w6417 = pi0236 & ~pi0877;
assign w6418 = ~w6416 & ~w6417;
assign w6419 = ~pi0243 & pi0759;
assign w6420 = ~pi0224 & pi0810;
assign w6421 = ~w6419 & ~w6420;
assign w6422 = pi0224 & ~pi0810;
assign w6423 = pi0242 & ~pi0809;
assign w6424 = ~pi0241 & pi0808;
assign w6425 = ~pi0242 & pi0809;
assign w6426 = ~w6424 & ~w6425;
assign w6427 = pi0221 & ~pi0755;
assign w6428 = pi0241 & ~pi0808;
assign w6429 = ~pi0221 & pi0755;
assign w6430 = ~pi0240 & pi0807;
assign w6431 = ~w6429 & ~w6430;
assign w6432 = pi0239 & ~pi0806;
assign w6433 = ~pi0238 & pi0804;
assign w6434 = ~pi0239 & pi0806;
assign w6435 = ~w6433 & ~w6434;
assign w6436 = pi0237 & ~pi0750;
assign w6437 = pi0238 & ~pi0804;
assign w6438 = ~w6436 & ~w6437;
assign w6439 = w6435 & ~w6438;
assign w6440 = pi0240 & ~pi0807;
assign w6441 = ~w6432 & ~w6440;
assign w6442 = (w6431 & w6439) | (w6431 & w12878) | (w6439 & w12878);
assign w6443 = ~w6427 & ~w6428;
assign w6444 = ~w6422 & ~w6423;
assign w6445 = (~w6442 & w12880) | (~w6442 & w12881) | (w12880 & w12881);
assign w6446 = (w6418 & w6445) | (w6418 & w12882) | (w6445 & w12882);
assign w6447 = ~w6415 & ~w6446;
assign w6448 = pi0257 & ~pi0859;
assign w6449 = ~pi0237 & pi0750;
assign w6450 = ~w6415 & ~w6449;
assign w6451 = w6421 & w6450;
assign w6452 = w6426 & w6431;
assign w6453 = w6435 & w6452;
assign w6454 = w6453 & w12883;
assign w6455 = (~w6454 & w6446) | (~w6454 & w12884) | (w6446 & w12884);
assign w6456 = pi0797 & ~w6455;
assign w6457 = ~w1513 & ~w1514;
assign w6458 = w1339 & ~w6457;
assign w6459 = ~w1339 & w6457;
assign w6460 = ~w6458 & ~w6459;
assign w6461 = pi0737 & ~pi1738;
assign w6462 = ~pi0737 & pi1738;
assign w6463 = ~w6461 & ~w6462;
assign w6464 = pi1725 & ~w6463;
assign w6465 = ~pi1725 & w6463;
assign w6466 = ~w6464 & ~w6465;
assign w6467 = ~w6385 & ~w6466;
assign w6468 = w6385 & w6466;
assign w6469 = ~w6467 & ~w6468;
assign w6470 = pi0736 & w6469;
assign w6471 = ~pi0736 & ~w6469;
assign w6472 = ~w6470 & ~w6471;
assign w6473 = w5585 & ~w6472;
assign w6474 = (pi0727 & ~w5584) | (pi0727 & w12885) | (~w5584 & w12885);
assign w6475 = ~w6388 & ~w6474;
assign w6476 = ~w6473 & w6475;
assign w6477 = pi1676 & pi1726;
assign w6478 = ~pi0728 & ~w6477;
assign w6479 = w1885 & ~w6478;
assign w6480 = (pi0729 & ~w5584) | (pi0729 & w12886) | (~w5584 & w12886);
assign w6481 = w5585 & ~w6469;
assign w6482 = ~w6388 & ~w6480;
assign w6483 = ~w6481 & w6482;
assign w6484 = w5584 & w12887;
assign w6485 = (pi0730 & ~w5584) | (pi0730 & w12888) | (~w5584 & w12888);
assign w6486 = ~w6388 & ~w6484;
assign w6487 = ~w6485 & w6486;
assign w6488 = w5584 & w12889;
assign w6489 = (pi0731 & ~w5584) | (pi0731 & w12890) | (~w5584 & w12890);
assign w6490 = ~w6388 & ~w6488;
assign w6491 = ~w6489 & w6490;
assign w6492 = w5584 & w12891;
assign w6493 = (pi0732 & ~w5584) | (pi0732 & w12892) | (~w5584 & w12892);
assign w6494 = ~w6388 & ~w6492;
assign w6495 = ~w6493 & w6494;
assign w6496 = (pi0733 & ~w5584) | (pi0733 & w12893) | (~w5584 & w12893);
assign w6497 = w6349 & ~w6370;
assign w6498 = w6370 & w6386;
assign w6499 = ~w6388 & ~w6496;
assign w6500 = ~w6497 & w6499;
assign w6501 = ~w6498 & w6500;
assign w6502 = (pi0734 & ~w5584) | (pi0734 & w12894) | (~w5584 & w12894);
assign w6503 = w6367 & ~w6373;
assign w6504 = ~w6367 & w6373;
assign w6505 = ~w6503 & ~w6504;
assign w6506 = w5585 & ~w6505;
assign w6507 = ~w6388 & ~w6502;
assign w6508 = ~w6506 & w6507;
assign w6509 = (pi0735 & ~w5584) | (pi0735 & w12895) | (~w5584 & w12895);
assign w6510 = w5585 & ~w6379;
assign w6511 = ~w6388 & ~w6509;
assign w6512 = ~w6510 & w6511;
assign w6513 = (pi0736 & ~w5584) | (pi0736 & w12896) | (~w5584 & w12896);
assign w6514 = w5585 & ~w6358;
assign w6515 = ~w6388 & ~w6513;
assign w6516 = ~w6514 & w6515;
assign w6517 = (pi0737 & ~w5584) | (pi0737 & w12897) | (~w5584 & w12897);
assign w6518 = ~pi0729 & ~w6361;
assign w6519 = pi0729 & w6361;
assign w6520 = ~w6518 & ~w6519;
assign w6521 = w6352 & w6520;
assign w6522 = ~w6352 & ~w6520;
assign w6523 = w5585 & ~w6521;
assign w6524 = ~w6522 & w6523;
assign w6525 = ~w6388 & ~w6517;
assign w6526 = ~w6524 & w6525;
assign w6527 = (pi0738 & ~w5584) | (pi0738 & w12898) | (~w5584 & w12898);
assign w6528 = ~pi0722 & ~w6361;
assign w6529 = pi0722 & w6361;
assign w6530 = ~w6528 & ~w6529;
assign w6531 = w5585 & ~w6530;
assign w6532 = ~w6388 & ~w6527;
assign w6533 = ~w6531 & w6532;
assign w6534 = ~pi0257 & pi0859;
assign w6535 = w6453 & w12899;
assign w6536 = pi0873 & ~w6535;
assign w6537 = ~w6447 & w6536;
assign w6538 = w5584 & w12900;
assign w6539 = (pi0744 & ~w5584) | (pi0744 & w12901) | (~w5584 & w12901);
assign w6540 = ~w6388 & ~w6538;
assign w6541 = ~w6539 & w6540;
assign w6542 = (pi0745 & ~w5584) | (pi0745 & w12902) | (~w5584 & w12902);
assign w6543 = w6355 & ~w6376;
assign w6544 = ~w6355 & w6376;
assign w6545 = ~w6543 & ~w6544;
assign w6546 = w5585 & ~w6545;
assign w6547 = ~w6388 & ~w6542;
assign w6548 = ~w6546 & w6547;
assign w6549 = (pi0746 & ~w5584) | (pi0746 & w12903) | (~w5584 & w12903);
assign w6550 = pi0738 & ~w6466;
assign w6551 = ~pi0738 & w6466;
assign w6552 = ~w6550 & ~w6551;
assign w6553 = w5585 & ~w6552;
assign w6554 = ~w6388 & ~w6549;
assign w6555 = ~w6553 & w6554;
assign w6556 = (~w215 & w12906) | (~w215 & w12907) | (w12906 & w12907);
assign w6557 = (~w215 & w12908) | (~w215 & w12909) | (w12908 & w12909);
assign w6558 = ~w6556 & w6557;
assign w6559 = ~pi0497 & w1867;
assign w6560 = w1829 & w12910;
assign w6561 = ~pi0398 & w1813;
assign w6562 = pi0748 & w1860;
assign w6563 = ~pi0667 & w1865;
assign w6564 = ~w6559 & ~w6561;
assign w6565 = ~w6560 & w6564;
assign w6566 = ~w6562 & w6565;
assign w6567 = ~w6563 & w6566;
assign w6568 = ~pi0501 & w1867;
assign w6569 = w1829 & w12911;
assign w6570 = ~pi0377 & w1813;
assign w6571 = ~pi0704 & w1865;
assign w6572 = pi0749 & w1860;
assign w6573 = ~w6568 & ~w6570;
assign w6574 = ~w6569 & w6573;
assign w6575 = ~w6571 & w6574;
assign w6576 = ~w6572 & w6575;
assign w6577 = pi1092 & w1867;
assign w6578 = w1829 & w12912;
assign w6579 = pi1280 & w1813;
assign w6580 = pi1104 & w1865;
assign w6581 = pi0750 & w1860;
assign w6582 = ~w6577 & ~w6579;
assign w6583 = ~w6578 & w6582;
assign w6584 = ~w6580 & w6583;
assign w6585 = ~w6581 & w6584;
assign w6586 = ~pi0494 & w1867;
assign w6587 = w1829 & w12913;
assign w6588 = ~pi0378 & w1813;
assign w6589 = pi0751 & w1860;
assign w6590 = ~pi0668 & w1865;
assign w6591 = ~w6586 & ~w6588;
assign w6592 = ~w6587 & w6591;
assign w6593 = ~w6589 & w6592;
assign w6594 = ~w6590 & w6593;
assign w6595 = ~pi0366 & w1867;
assign w6596 = w1829 & w12914;
assign w6597 = ~pi0318 & w1813;
assign w6598 = ~pi0752 & w1860;
assign w6599 = ~pi0635 & w1865;
assign w6600 = ~w6595 & ~w6597;
assign w6601 = ~w6596 & w6600;
assign w6602 = ~w6598 & w6601;
assign w6603 = ~w6599 & w6602;
assign w6604 = w2863 & w12915;
assign w6605 = ~pi1759 & ~pi1760;
assign w6606 = w6604 & w12916;
assign w6607 = pi1479 & w6606;
assign w6608 = ~pi1759 & pi1760;
assign w6609 = w3952 & w12917;
assign w6610 = pi1165 & w6609;
assign w6611 = ~pi0684 & w5442;
assign w6612 = w3952 & w12918;
assign w6613 = pi1104 & w6612;
assign w6614 = ~pi0394 & w2932;
assign w6615 = w6604 & w12919;
assign w6616 = pi1319 & w6615;
assign w6617 = ~pi0529 & w3953;
assign w6618 = w2864 & w12917;
assign w6619 = pi1037 & w6618;
assign w6620 = w2864 & w12920;
assign w6621 = pi1280 & w6620;
assign w6622 = w3952 & w12920;
assign w6623 = pi1271 & w6622;
assign w6624 = w2864 & w12921;
assign w6625 = pi0991 & w6624;
assign w6626 = ~pi0440 & w3188;
assign w6627 = w2864 & w12918;
assign w6628 = pi1092 & w6627;
assign w6629 = w3952 & w12921;
assign w6630 = pi1035 & w6629;
assign w6631 = ~pi0417 & w3150;
assign w6632 = ~pi0575 & w4186;
assign w6633 = w6604 & w12922;
assign w6634 = pi0474 & w6633;
assign w6635 = ~pi0340 & w2866;
assign w6636 = ~pi0599 & w4056;
assign w6637 = w6604 & w12923;
assign w6638 = pi1487 & w6637;
assign w6639 = w6604 & w12924;
assign w6640 = pi1095 & w6639;
assign w6641 = w6604 & w12925;
assign w6642 = pi1684 & w6641;
assign w6643 = ~w6610 & ~w6611;
assign w6644 = ~w6613 & ~w6614;
assign w6645 = ~w6617 & ~w6619;
assign w6646 = ~w6621 & ~w6623;
assign w6647 = ~w6625 & ~w6626;
assign w6648 = ~w6628 & ~w6630;
assign w6649 = ~w6631 & ~w6632;
assign w6650 = ~w6635 & ~w6636;
assign w6651 = w6649 & w6650;
assign w6652 = w6647 & w6648;
assign w6653 = w6645 & w6646;
assign w6654 = w6643 & w6644;
assign w6655 = ~w6607 & ~w6616;
assign w6656 = ~w6634 & ~w6638;
assign w6657 = ~w6640 & ~w6642;
assign w6658 = w6656 & w6657;
assign w6659 = w6654 & w6655;
assign w6660 = w6652 & w6653;
assign w6661 = w6651 & w6660;
assign w6662 = w6658 & w6659;
assign w6663 = w6661 & w6662;
assign w6664 = ~pi0491 & w1867;
assign w6665 = w1829 & w12926;
assign w6666 = ~pi0430 & w1813;
assign w6667 = ~pi0671 & w1865;
assign w6668 = pi0754 & w1860;
assign w6669 = ~w6664 & ~w6666;
assign w6670 = ~w6665 & w6669;
assign w6671 = ~w6667 & w6670;
assign w6672 = ~w6668 & w6671;
assign w6673 = pi1028 & w1867;
assign w6674 = w1829 & w12927;
assign w6675 = pi1272 & w1813;
assign w6676 = pi0755 & w1860;
assign w6677 = pi1107 & w1865;
assign w6678 = ~w6673 & ~w6675;
assign w6679 = ~w6674 & w6678;
assign w6680 = ~w6676 & w6679;
assign w6681 = ~w6677 & w6680;
assign w6682 = ~pi0425 & w1867;
assign w6683 = w1829 & w12928;
assign w6684 = ~pi0348 & w1813;
assign w6685 = ~pi0756 & w1860;
assign w6686 = ~pi0609 & w1865;
assign w6687 = ~w6682 & ~w6684;
assign w6688 = ~w6683 & w6687;
assign w6689 = ~w6685 & w6688;
assign w6690 = ~w6686 & w6689;
assign w6691 = ~pi0371 & w1867;
assign w6692 = w1829 & w12929;
assign w6693 = ~pi0324 & w1813;
assign w6694 = ~pi0757 & w1860;
assign w6695 = ~pi0558 & w1865;
assign w6696 = ~w6691 & ~w6693;
assign w6697 = ~w6692 & w6696;
assign w6698 = ~w6694 & w6697;
assign w6699 = ~w6695 & w6698;
assign w6700 = ~pi0369 & w1867;
assign w6701 = w1829 & w12930;
assign w6702 = ~pi0322 & w1813;
assign w6703 = ~pi0758 & w1860;
assign w6704 = ~pi0636 & w1865;
assign w6705 = ~w6700 & ~w6702;
assign w6706 = ~w6701 & w6705;
assign w6707 = ~w6703 & w6706;
assign w6708 = ~w6704 & w6707;
assign w6709 = pi1029 & w1867;
assign w6710 = w1829 & w12931;
assign w6711 = pi1267 & w1813;
assign w6712 = pi0759 & w1860;
assign w6713 = pi1110 & w1865;
assign w6714 = ~w6709 & ~w6711;
assign w6715 = ~w6710 & w6714;
assign w6716 = ~w6712 & w6715;
assign w6717 = ~w6713 & w6716;
assign w6718 = pi1747 & ~pi1757;
assign w6719 = pi0760 & w2138;
assign w6720 = w2166 & w6719;
assign w6721 = w2166 & w12932;
assign w6722 = pi0773 & pi0937;
assign w6723 = ~w2136 & ~w6722;
assign w6724 = w2139 & w6723;
assign w6725 = w6724 & w12933;
assign w6726 = ~w6721 & ~w6725;
assign w6727 = w6718 & ~w6726;
assign w6728 = pi0872 & pi1665;
assign w6729 = w6406 & w12935;
assign w6730 = w6406 & w12936;
assign w6731 = w6406 & w12937;
assign w6732 = pi0761 & w6731;
assign w6733 = ~w6730 & ~w6732;
assign w6734 = ~pi0616 & w1867;
assign w6735 = w1829 & w12938;
assign w6736 = ~pi0519 & w1813;
assign w6737 = ~pi0542 & w1865;
assign w6738 = pi0762 & w1860;
assign w6739 = ~w6734 & ~w6736;
assign w6740 = ~w6735 & w6739;
assign w6741 = ~w6737 & w6740;
assign w6742 = ~w6738 & w6741;
assign w6743 = ~pi0791 & ~pi0792;
assign w6744 = pi0763 & ~w6743;
assign w6745 = w6406 & w12939;
assign w6746 = ~pi0763 & w6743;
assign w6747 = ~w6744 & ~w6746;
assign w6748 = w6745 & w6747;
assign w6749 = w6406 & w12940;
assign w6750 = w6406 & w12941;
assign w6751 = ~w6749 & ~w6750;
assign w6752 = w6406 & w12942;
assign w6753 = w6406 & w12943;
assign w6754 = ~w6752 & ~w6753;
assign w6755 = w6406 & w12944;
assign w6756 = w6406 & w12945;
assign w6757 = ~w6755 & ~w6756;
assign w6758 = pi0938 & w1867;
assign w6759 = w1829 & w12946;
assign w6760 = pi0861 & w1813;
assign w6761 = pi0767 & w1860;
assign w6762 = pi0992 & w1865;
assign w6763 = ~w6758 & ~w6760;
assign w6764 = ~w6759 & w6763;
assign w6765 = ~w6761 & w6764;
assign w6766 = ~w6762 & w6765;
assign w6767 = ~pi0424 & w1867;
assign w6768 = w1829 & w12947;
assign w6769 = ~pi0347 & w1813;
assign w6770 = ~pi0608 & w1865;
assign w6771 = pi0768 & w1860;
assign w6772 = ~w6767 & ~w6769;
assign w6773 = ~w6768 & w6772;
assign w6774 = ~w6770 & w6773;
assign w6775 = ~w6771 & w6774;
assign w6776 = ~pi1060 & ~pi1773;
assign w6777 = pi1773 & ~pi1829;
assign w6778 = ~w6776 & ~w6777;
assign w6779 = ~pi0419 & w1867;
assign w6780 = w1829 & w12948;
assign w6781 = ~pi0342 & w1813;
assign w6782 = ~pi0546 & w1865;
assign w6783 = pi0770 & w1860;
assign w6784 = ~w6779 & ~w6781;
assign w6785 = ~w6780 & w6784;
assign w6786 = ~w6782 & w6785;
assign w6787 = ~w6783 & w6786;
assign w6788 = pi1132 & w1867;
assign w6789 = w1829 & w12949;
assign w6790 = pi1257 & w1813;
assign w6791 = pi1113 & w1865;
assign w6792 = pi0771 & w1860;
assign w6793 = ~w6788 & ~w6790;
assign w6794 = ~w6789 & w6793;
assign w6795 = ~w6791 & w6794;
assign w6796 = ~w6792 & w6795;
assign w6797 = ~pi0422 & w1867;
assign w6798 = w1829 & w12950;
assign w6799 = ~pi0345 & w1813;
assign w6800 = ~pi0544 & w1865;
assign w6801 = pi0772 & w1860;
assign w6802 = ~w6797 & ~w6799;
assign w6803 = ~w6798 & w6802;
assign w6804 = ~w6800 & w6803;
assign w6805 = ~w6801 & w6804;
assign w6806 = ~pi1045 & w6718;
assign w6807 = ~pi1737 & ~pi1739;
assign w6808 = pi1674 & w6807;
assign w6809 = (~pi0937 & ~w6807) | (~pi0937 & w12951) | (~w6807 & w12951);
assign w6810 = ~w6397 & ~w6809;
assign w6811 = w6724 & w12952;
assign w6812 = ~w2133 & w6811;
assign w6813 = w6811 & w12953;
assign w6814 = w2140 & w12954;
assign w6815 = pi0984 & w6814;
assign w6816 = w6814 & w12955;
assign w6817 = ~w6813 & ~w6816;
assign w6818 = w6806 & ~w6817;
assign w6819 = pi0759 & ~pi0825;
assign w6820 = ~pi0826 & pi0877;
assign w6821 = pi0772 & ~pi0810;
assign w6822 = ~pi0759 & pi0825;
assign w6823 = pi0809 & ~pi0824;
assign w6824 = ~pi0772 & pi0810;
assign w6825 = ~pi0809 & pi0824;
assign w6826 = ~pi0808 & pi0823;
assign w6827 = pi0755 & ~pi0822;
assign w6828 = pi0808 & ~pi0823;
assign w6829 = ~pi0755 & pi0822;
assign w6830 = pi0770 & ~pi0807;
assign w6831 = ~pi0770 & pi0807;
assign w6832 = pi0806 & ~pi0821;
assign w6833 = ~pi0806 & pi0821;
assign w6834 = ~pi0804 & pi0819;
assign w6835 = pi0750 & ~pi0871;
assign w6836 = pi0804 & ~pi0819;
assign w6837 = ~pi0750 & pi0871;
assign w6838 = ~pi0818 & pi0859;
assign w6839 = ~w6837 & w6838;
assign w6840 = ~w6835 & ~w6836;
assign w6841 = ~w6839 & w6840;
assign w6842 = ~w6833 & ~w6834;
assign w6843 = ~w6831 & ~w6832;
assign w6844 = (w6843 & w6841) | (w6843 & w12956) | (w6841 & w12956);
assign w6845 = ~w6829 & ~w6830;
assign w6846 = ~w6827 & ~w6828;
assign w6847 = ~w6825 & ~w6826;
assign w6848 = (~w6844 & w12958) | (~w6844 & w12959) | (w12958 & w12959);
assign w6849 = ~w6823 & ~w6824;
assign w6850 = ~w6821 & ~w6822;
assign w6851 = ~w6819 & ~w6820;
assign w6852 = (~w6848 & w12961) | (~w6848 & w12962) | (w12961 & w12962);
assign w6853 = pi0826 & ~pi0877;
assign w6854 = ~pi0762 & ~pi0768;
assign w6855 = ~pi0827 & w6854;
assign w6856 = ~w6853 & w6855;
assign w6857 = ~w6852 & w6856;
assign w6858 = (w215 & w12963) | (w215 & w12964) | (w12963 & w12964);
assign w6859 = (~w215 & w12965) | (~w215 & w12966) | (w12965 & w12966);
assign w6860 = ~w634 & ~w6858;
assign w6861 = ~w6859 & w6860;
assign w6862 = ~pi0060 & ~w624;
assign w6863 = pi0778 & w624;
assign w6864 = ~w634 & ~w6862;
assign w6865 = ~w6863 & w6864;
assign w6866 = ~pi0052 & ~w624;
assign w6867 = pi0779 & w624;
assign w6868 = ~w634 & ~w6866;
assign w6869 = ~w6867 & w6868;
assign w6870 = ~pi1206 & w1867;
assign w6871 = ~pi1225 & w1862;
assign w6872 = ~pi1184 & w1813;
assign w6873 = ~pi1164 & w1865;
assign w6874 = pi0780 & w1860;
assign w6875 = ~w6870 & ~w6872;
assign w6876 = ~w6871 & w6875;
assign w6877 = ~w6873 & w6876;
assign w6878 = ~w6874 & w6877;
assign w6879 = ~pi1059 & ~pi1773;
assign w6880 = pi1773 & ~pi1828;
assign w6881 = ~w6879 & ~w6880;
assign w6882 = ~pi1061 & ~pi1773;
assign w6883 = pi1773 & ~pi1813;
assign w6884 = ~w6882 & ~w6883;
assign w6885 = pi1550 & w6729;
assign w6886 = pi0783 & w6731;
assign w6887 = ~w6885 & ~w6886;
assign w6888 = ~pi1072 & ~pi1773;
assign w6889 = pi1773 & ~pi1814;
assign w6890 = ~w6888 & ~w6889;
assign w6891 = ~pi0764 & ~pi0790;
assign w6892 = ~pi0761 & ~pi0787;
assign w6893 = ~pi0783 & ~pi0788;
assign w6894 = w6892 & w6893;
assign w6895 = w6891 & ~w6894;
assign w6896 = w6407 & ~w6895;
assign w6897 = w6406 & ~w6896;
assign w6898 = pi1675 & pi1680;
assign w6899 = ~pi0786 & ~w6898;
assign w6900 = w1885 & ~w6899;
assign w6901 = pi1705 & w6729;
assign w6902 = pi0787 & w6731;
assign w6903 = ~w6901 & ~w6902;
assign w6904 = pi1631 & w6729;
assign w6905 = pi0788 & w6731;
assign w6906 = ~w6904 & ~w6905;
assign w6907 = ~pi0917 & w5585;
assign w6908 = ~pi0789 & ~w1232;
assign w6909 = ~w6907 & ~w6908;
assign w6910 = pi1747 & ~w6909;
assign w6911 = pi1546 & w6729;
assign w6912 = ~pi0790 & w6731;
assign w6913 = ~w6911 & ~w6912;
assign w6914 = pi0791 & w6745;
assign w6915 = pi0791 & pi0792;
assign w6916 = ~w6743 & ~w6915;
assign w6917 = w6745 & w6916;
assign w6918 = pi0793 & ~w6746;
assign w6919 = ~pi0793 & w6746;
assign w6920 = ~w6918 & ~w6919;
assign w6921 = w6745 & w6920;
assign w6922 = ~pi0794 & ~pi1751;
assign w6923 = pi1315 & pi1747;
assign w6924 = ~w6922 & w6923;
assign w6925 = ~pi1084 & w1867;
assign w6926 = ~pi1140 & w1862;
assign w6927 = ~pi1120 & w1813;
assign w6928 = pi0795 & w1860;
assign w6929 = ~pi1103 & w1865;
assign w6930 = ~w6925 & ~w6927;
assign w6931 = ~w6926 & w6930;
assign w6932 = ~w6928 & w6931;
assign w6933 = ~w6929 & w6932;
assign w6934 = pi1131 & w1867;
assign w6935 = pi1143 & w1862;
assign w6936 = pi1122 & w1813;
assign w6937 = pi0796 & w1860;
assign w6938 = pi1111 & w1865;
assign w6939 = ~w6934 & ~w6936;
assign w6940 = ~w6935 & w6939;
assign w6941 = ~w6937 & w6940;
assign w6942 = ~w6938 & w6941;
assign w6943 = ~pi1133 & w1867;
assign w6944 = pi1255 & w1862;
assign w6945 = pi1025 & w1813;
assign w6946 = pi1051 & w1865;
assign w6947 = ~pi0797 & w1860;
assign w6948 = ~w6943 & ~w6945;
assign w6949 = ~w6944 & w6948;
assign w6950 = ~w6946 & w6949;
assign w6951 = ~w6947 & w6950;
assign w6952 = ~pi1369 & w1867;
assign w6953 = ~pi1413 & w1862;
assign w6954 = ~pi1360 & w1813;
assign w6955 = pi0798 & w1860;
assign w6956 = ~pi1361 & w1865;
assign w6957 = ~w6952 & ~w6954;
assign w6958 = ~w6953 & w6957;
assign w6959 = ~w6955 & w6958;
assign w6960 = ~w6956 & w6959;
assign w6961 = ~pi1137 & w1867;
assign w6962 = pi1242 & w1862;
assign w6963 = pi1124 & w1813;
assign w6964 = pi0799 & w1860;
assign w6965 = pi1118 & w1865;
assign w6966 = ~w6961 & ~w6963;
assign w6967 = ~w6962 & w6966;
assign w6968 = ~w6964 & w6967;
assign w6969 = ~w6965 & w6968;
assign w6970 = ~pi1030 & w1867;
assign w6971 = pi1261 & w1862;
assign w6972 = pi1252 & w1813;
assign w6973 = pi1074 & w1865;
assign w6974 = pi0800 & w1860;
assign w6975 = ~w6970 & ~w6972;
assign w6976 = ~w6971 & w6975;
assign w6977 = ~w6973 & w6976;
assign w6978 = ~w6974 & w6977;
assign w6979 = pi1080 & w1867;
assign w6980 = pi1144 & w1862;
assign w6981 = pi1256 & w1813;
assign w6982 = pi0801 & w1860;
assign w6983 = pi1112 & w1865;
assign w6984 = ~w6979 & ~w6981;
assign w6985 = ~w6980 & w6984;
assign w6986 = ~w6982 & w6985;
assign w6987 = ~w6983 & w6986;
assign w6988 = pi0939 & w1867;
assign w6989 = pi0969 & w1862;
assign w6990 = pi0863 & w1813;
assign w6991 = pi0802 & w1860;
assign w6992 = pi0994 & w1865;
assign w6993 = ~w6988 & ~w6990;
assign w6994 = ~w6989 & w6993;
assign w6995 = ~w6991 & w6994;
assign w6996 = ~w6992 & w6995;
assign w6997 = pi0942 & w1867;
assign w6998 = pi0973 & w1862;
assign w6999 = pi0876 & w1813;
assign w7000 = pi1014 & w1865;
assign w7001 = pi0803 & w1860;
assign w7002 = ~w6997 & ~w6999;
assign w7003 = ~w6998 & w7002;
assign w7004 = ~w7000 & w7003;
assign w7005 = ~w7001 & w7004;
assign w7006 = pi1027 & w1867;
assign w7007 = pi1032 & w1862;
assign w7008 = pi1022 & w1813;
assign w7009 = pi1105 & w1865;
assign w7010 = pi0804 & w1860;
assign w7011 = ~w7006 & ~w7008;
assign w7012 = ~w7007 & w7011;
assign w7013 = ~w7009 & w7012;
assign w7014 = ~w7010 & w7013;
assign w7015 = pi0941 & w1867;
assign w7016 = pi0968 & w1862;
assign w7017 = pi0862 & w1813;
assign w7018 = pi0993 & w1865;
assign w7019 = ~pi0805 & w1860;
assign w7020 = ~w7015 & ~w7017;
assign w7021 = ~w7016 & w7020;
assign w7022 = ~w7018 & w7021;
assign w7023 = ~w7019 & w7022;
assign w7024 = pi1310 & w1867;
assign w7025 = pi1342 & w1862;
assign w7026 = pi1277 & w1813;
assign w7027 = pi0806 & w1860;
assign w7028 = pi1338 & w1865;
assign w7029 = ~w7024 & ~w7026;
assign w7030 = ~w7025 & w7029;
assign w7031 = ~w7027 & w7030;
assign w7032 = ~w7028 & w7031;
assign w7033 = pi1129 & w1867;
assign w7034 = pi1141 & w1862;
assign w7035 = pi1023 & w1813;
assign w7036 = pi0807 & w1860;
assign w7037 = pi1106 & w1865;
assign w7038 = ~w7033 & ~w7035;
assign w7039 = ~w7034 & w7038;
assign w7040 = ~w7036 & w7039;
assign w7041 = ~w7037 & w7040;
assign w7042 = pi1083 & w1867;
assign w7043 = pi1033 & w1862;
assign w7044 = pi1121 & w1813;
assign w7045 = pi1108 & w1865;
assign w7046 = pi0808 & w1860;
assign w7047 = ~w7042 & ~w7044;
assign w7048 = ~w7043 & w7047;
assign w7049 = ~w7045 & w7048;
assign w7050 = ~w7046 & w7049;
assign w7051 = pi1130 & w1867;
assign w7052 = pi1142 & w1862;
assign w7053 = pi1274 & w1813;
assign w7054 = pi1081 & w1865;
assign w7055 = pi0809 & w1860;
assign w7056 = ~w7051 & ~w7053;
assign w7057 = ~w7052 & w7056;
assign w7058 = ~w7054 & w7057;
assign w7059 = ~w7055 & w7058;
assign w7060 = pi1076 & w1867;
assign w7061 = pi1265 & w1862;
assign w7062 = pi1270 & w1813;
assign w7063 = pi1109 & w1865;
assign w7064 = pi0810 & w1860;
assign w7065 = ~w7060 & ~w7062;
assign w7066 = ~w7061 & w7065;
assign w7067 = ~w7063 & w7066;
assign w7068 = ~w7064 & w7067;
assign w7069 = ~pi0612 & w1867;
assign w7070 = ~pi0520 & w1862;
assign w7071 = ~pi0337 & w1813;
assign w7072 = ~pi0593 & w1865;
assign w7073 = ~pi0811 & w1860;
assign w7074 = ~w7069 & ~w7071;
assign w7075 = ~w7070 & w7074;
assign w7076 = ~w7072 & w7075;
assign w7077 = ~w7073 & w7076;
assign w7078 = ~pi0364 & w1867;
assign w7079 = ~pi0451 & w1862;
assign w7080 = ~pi0316 & w1813;
assign w7081 = ~pi0812 & w1860;
assign w7082 = ~pi0551 & w1865;
assign w7083 = ~w7078 & ~w7080;
assign w7084 = ~w7079 & w7083;
assign w7085 = ~w7081 & w7084;
assign w7086 = ~w7082 & w7085;
assign w7087 = ~pi0367 & w1867;
assign w7088 = ~pi0450 & w1862;
assign w7089 = ~pi0319 & w1813;
assign w7090 = ~pi0813 & w1860;
assign w7091 = ~pi0555 & w1865;
assign w7092 = ~w7087 & ~w7089;
assign w7093 = ~w7088 & w7092;
assign w7094 = ~w7090 & w7093;
assign w7095 = ~w7091 & w7094;
assign w7096 = ~pi0613 & w1867;
assign w7097 = ~pi0439 & w1862;
assign w7098 = ~pi0516 & w1813;
assign w7099 = ~pi0601 & w1865;
assign w7100 = ~pi0814 & w1860;
assign w7101 = ~w7096 & ~w7098;
assign w7102 = ~w7097 & w7101;
assign w7103 = ~w7099 & w7102;
assign w7104 = ~w7100 & w7103;
assign w7105 = ~pi0365 & w1867;
assign w7106 = ~pi0453 & w1862;
assign w7107 = ~pi0317 & w1813;
assign w7108 = ~pi0815 & w1860;
assign w7109 = ~pi0554 & w1865;
assign w7110 = ~w7105 & ~w7107;
assign w7111 = ~w7106 & w7110;
assign w7112 = ~w7108 & w7111;
assign w7113 = ~w7109 & w7112;
assign w7114 = ~pi0368 & w1867;
assign w7115 = ~pi0455 & w1862;
assign w7116 = ~pi0320 & w1813;
assign w7117 = ~pi0556 & w1865;
assign w7118 = ~pi0816 & w1860;
assign w7119 = ~w7114 & ~w7116;
assign w7120 = ~w7115 & w7119;
assign w7121 = ~w7117 & w7120;
assign w7122 = ~w7118 & w7121;
assign w7123 = ~pi0414 & w1867;
assign w7124 = ~pi0521 & w1862;
assign w7125 = ~pi0517 & w1813;
assign w7126 = ~pi0817 & w1860;
assign w7127 = ~pi0595 & w1865;
assign w7128 = ~w7123 & ~w7125;
assign w7129 = ~w7124 & w7128;
assign w7130 = ~w7126 & w7129;
assign w7131 = ~w7127 & w7130;
assign w7132 = ~pi0614 & w1867;
assign w7133 = ~pi0522 & w1862;
assign w7134 = ~pi0518 & w1813;
assign w7135 = ~pi0596 & w1865;
assign w7136 = pi0818 & w1860;
assign w7137 = ~w7132 & ~w7134;
assign w7138 = ~w7133 & w7137;
assign w7139 = ~w7135 & w7138;
assign w7140 = ~w7136 & w7139;
assign w7141 = ~pi0416 & w1867;
assign w7142 = ~pi0444 & w1862;
assign w7143 = ~pi0339 & w1813;
assign w7144 = ~pi0598 & w1865;
assign w7145 = pi0819 & w1860;
assign w7146 = ~w7141 & ~w7143;
assign w7147 = ~w7142 & w7146;
assign w7148 = ~w7144 & w7147;
assign w7149 = ~w7145 & w7148;
assign w7150 = ~pi0417 & w1867;
assign w7151 = ~pi0529 & w1862;
assign w7152 = ~pi0340 & w1813;
assign w7153 = ~pi0820 & w1860;
assign w7154 = ~pi0599 & w1865;
assign w7155 = ~w7150 & ~w7152;
assign w7156 = ~w7151 & w7155;
assign w7157 = ~w7153 & w7156;
assign w7158 = ~w7154 & w7157;
assign w7159 = ~pi0418 & w1867;
assign w7160 = ~pi0524 & w1862;
assign w7161 = ~pi0341 & w1813;
assign w7162 = pi0821 & w1860;
assign w7163 = ~pi0600 & w1865;
assign w7164 = ~w7159 & ~w7161;
assign w7165 = ~w7160 & w7164;
assign w7166 = ~w7162 & w7165;
assign w7167 = ~w7163 & w7166;
assign w7168 = ~pi0536 & w1867;
assign w7169 = ~pi0525 & w1862;
assign w7170 = ~pi0438 & w1813;
assign w7171 = ~pi0604 & w1865;
assign w7172 = pi0822 & w1860;
assign w7173 = ~w7168 & ~w7170;
assign w7174 = ~w7169 & w7173;
assign w7175 = ~w7171 & w7174;
assign w7176 = ~w7172 & w7175;
assign w7177 = ~pi0420 & w1867;
assign w7178 = ~pi0657 & w1862;
assign w7179 = ~pi0343 & w1813;
assign w7180 = pi0823 & w1860;
assign w7181 = ~pi0602 & w1865;
assign w7182 = ~w7177 & ~w7179;
assign w7183 = ~w7178 & w7182;
assign w7184 = ~w7180 & w7183;
assign w7185 = ~w7181 & w7184;
assign w7186 = ~pi0421 & w1867;
assign w7187 = ~pi0526 & w1862;
assign w7188 = ~pi0344 & w1813;
assign w7189 = pi0824 & w1860;
assign w7190 = ~pi0603 & w1865;
assign w7191 = ~w7186 & ~w7188;
assign w7192 = ~w7187 & w7191;
assign w7193 = ~w7189 & w7192;
assign w7194 = ~w7190 & w7193;
assign w7195 = ~pi0432 & w1867;
assign w7196 = ~pi0629 & w1862;
assign w7197 = ~pi0346 & w1813;
assign w7198 = ~pi0606 & w1865;
assign w7199 = pi0825 & w1860;
assign w7200 = ~w7195 & ~w7197;
assign w7201 = ~w7196 & w7200;
assign w7202 = ~w7198 & w7201;
assign w7203 = ~w7199 & w7202;
assign w7204 = ~pi0423 & w1867;
assign w7205 = ~pi0658 & w1862;
assign w7206 = ~pi0314 & w1813;
assign w7207 = pi0826 & w1860;
assign w7208 = ~pi0605 & w1865;
assign w7209 = ~w7204 & ~w7206;
assign w7210 = ~w7205 & w7209;
assign w7211 = ~w7207 & w7210;
assign w7212 = ~w7208 & w7211;
assign w7213 = ~pi0350 & w1867;
assign w7214 = ~pi0427 & w1862;
assign w7215 = ~pi0311 & w1813;
assign w7216 = pi0827 & w1860;
assign w7217 = ~pi0515 & w1865;
assign w7218 = ~w7213 & ~w7215;
assign w7219 = ~w7214 & w7218;
assign w7220 = ~w7216 & w7219;
assign w7221 = ~w7217 & w7220;
assign w7222 = ~pi0534 & w1867;
assign w7223 = ~pi0626 & w1862;
assign w7224 = ~pi0435 & w1813;
assign w7225 = ~pi0828 & w1860;
assign w7226 = ~pi0607 & w1865;
assign w7227 = ~w7222 & ~w7224;
assign w7228 = ~w7223 & w7227;
assign w7229 = ~w7225 & w7228;
assign w7230 = ~w7226 & w7229;
assign w7231 = ~pi0351 & w1867;
assign w7232 = ~pi0428 & w1862;
assign w7233 = ~pi0312 & w1813;
assign w7234 = ~pi0829 & w1860;
assign w7235 = ~pi0437 & w1865;
assign w7236 = ~w7231 & ~w7233;
assign w7237 = ~w7232 & w7236;
assign w7238 = ~w7234 & w7237;
assign w7239 = ~w7235 & w7238;
assign w7240 = ~pi0559 & w1867;
assign w7241 = ~pi0632 & w1862;
assign w7242 = ~pi0458 & w1813;
assign w7243 = ~pi0830 & w1860;
assign w7244 = ~pi0557 & w1865;
assign w7245 = ~w7240 & ~w7242;
assign w7246 = ~w7241 & w7245;
assign w7247 = ~w7243 & w7246;
assign w7248 = ~w7244 & w7247;
assign w7249 = ~pi0548 & w1867;
assign w7250 = ~pi0640 & w1862;
assign w7251 = ~pi0447 & w1813;
assign w7252 = ~pi0831 & w1860;
assign w7253 = ~pi0547 & w1865;
assign w7254 = ~w7249 & ~w7251;
assign w7255 = ~w7250 & w7254;
assign w7256 = ~w7252 & w7255;
assign w7257 = ~w7253 & w7256;
assign w7258 = ~pi0362 & w1867;
assign w7259 = ~pi0449 & w1862;
assign w7260 = ~pi0321 & w1813;
assign w7261 = ~pi0550 & w1865;
assign w7262 = ~pi0832 & w1860;
assign w7263 = ~w7258 & ~w7260;
assign w7264 = ~w7259 & w7263;
assign w7265 = ~w7261 & w7264;
assign w7266 = ~w7262 & w7265;
assign w7267 = ~pi0356 & w1867;
assign w7268 = ~pi0436 & w1862;
assign w7269 = ~pi0349 & w1813;
assign w7270 = ~pi0833 & w1860;
assign w7271 = ~pi0610 & w1865;
assign w7272 = ~w7267 & ~w7269;
assign w7273 = ~w7268 & w7272;
assign w7274 = ~w7270 & w7273;
assign w7275 = ~w7271 & w7274;
assign w7276 = ~pi0426 & w1867;
assign w7277 = ~pi0659 & w1862;
assign w7278 = ~pi0313 & w1813;
assign w7279 = ~pi0611 & w1865;
assign w7280 = ~pi0834 & w1860;
assign w7281 = ~w7276 & ~w7278;
assign w7282 = ~w7277 & w7281;
assign w7283 = ~w7279 & w7282;
assign w7284 = ~w7280 & w7283;
assign w7285 = ~pi0487 & w1867;
assign w7286 = ~pi0570 & w1862;
assign w7287 = ~pi0389 & w1813;
assign w7288 = ~pi0670 & w1865;
assign w7289 = ~pi0835 & w1860;
assign w7290 = ~w7285 & ~w7287;
assign w7291 = ~w7286 & w7290;
assign w7292 = ~w7288 & w7291;
assign w7293 = ~w7289 & w7292;
assign w7294 = ~pi0372 & w1867;
assign w7295 = ~pi0460 & w1862;
assign w7296 = ~pi0325 & w1813;
assign w7297 = ~pi0836 & w1860;
assign w7298 = ~pi0638 & w1865;
assign w7299 = ~w7294 & ~w7296;
assign w7300 = ~w7295 & w7299;
assign w7301 = ~w7297 & w7300;
assign w7302 = ~w7298 & w7301;
assign w7303 = ~pi0488 & w1867;
assign w7304 = ~pi0571 & w1862;
assign w7305 = ~pi0390 & w1813;
assign w7306 = ~pi0837 & w1860;
assign w7307 = ~pi0680 & w1865;
assign w7308 = ~w7303 & ~w7305;
assign w7309 = ~w7304 & w7308;
assign w7310 = ~w7306 & w7309;
assign w7311 = ~w7307 & w7310;
assign w7312 = ~pi0370 & w1867;
assign w7313 = ~pi0457 & w1862;
assign w7314 = ~pi0323 & w1813;
assign w7315 = ~pi0838 & w1860;
assign w7316 = ~pi0637 & w1865;
assign w7317 = ~w7312 & ~w7314;
assign w7318 = ~w7313 & w7317;
assign w7319 = ~w7315 & w7318;
assign w7320 = ~w7316 & w7319;
assign w7321 = ~pi0373 & w1867;
assign w7322 = ~pi0532 & w1862;
assign w7323 = ~pi0326 & w1813;
assign w7324 = ~pi0639 & w1865;
assign w7325 = ~pi0839 & w1860;
assign w7326 = ~w7321 & ~w7323;
assign w7327 = ~w7322 & w7326;
assign w7328 = ~w7324 & w7327;
assign w7329 = ~w7325 & w7328;
assign w7330 = ~pi0489 & w1867;
assign w7331 = ~pi0572 & w1862;
assign w7332 = ~pi0391 & w1813;
assign w7333 = ~pi0681 & w1865;
assign w7334 = ~pi0840 & w1860;
assign w7335 = ~w7330 & ~w7332;
assign w7336 = ~w7331 & w7335;
assign w7337 = ~w7333 & w7336;
assign w7338 = ~w7334 & w7337;
assign w7339 = ~pi0490 & w1867;
assign w7340 = ~pi0543 & w1862;
assign w7341 = ~pi0392 & w1813;
assign w7342 = ~pi0682 & w1865;
assign w7343 = pi0841 & w1860;
assign w7344 = ~w7339 & ~w7341;
assign w7345 = ~w7340 & w7344;
assign w7346 = ~w7342 & w7345;
assign w7347 = ~w7343 & w7346;
assign w7348 = ~pi0492 & w1867;
assign w7349 = ~pi0574 & w1862;
assign w7350 = ~pi0393 & w1813;
assign w7351 = pi0842 & w1860;
assign w7352 = ~pi0683 & w1865;
assign w7353 = ~w7348 & ~w7350;
assign w7354 = ~w7349 & w7353;
assign w7355 = ~w7351 & w7354;
assign w7356 = ~w7352 & w7355;
assign w7357 = ~pi0440 & w1867;
assign w7358 = ~pi0575 & w1862;
assign w7359 = ~pi0394 & w1813;
assign w7360 = ~pi0684 & w1865;
assign w7361 = ~pi0843 & w1860;
assign w7362 = ~w7357 & ~w7359;
assign w7363 = ~w7358 & w7362;
assign w7364 = ~w7360 & w7363;
assign w7365 = ~w7361 & w7364;
assign w7366 = ~pi0493 & w1867;
assign w7367 = ~pi0538 & w1862;
assign w7368 = ~pi0395 & w1813;
assign w7369 = pi0844 & w1860;
assign w7370 = ~pi0685 & w1865;
assign w7371 = ~w7366 & ~w7368;
assign w7372 = ~w7367 & w7371;
assign w7373 = ~w7369 & w7372;
assign w7374 = ~w7370 & w7373;
assign w7375 = ~pi0495 & w1867;
assign w7376 = ~pi0576 & w1862;
assign w7377 = ~pi0396 & w1813;
assign w7378 = pi0845 & w1860;
assign w7379 = ~pi0686 & w1865;
assign w7380 = ~w7375 & ~w7377;
assign w7381 = ~w7376 & w7380;
assign w7382 = ~w7378 & w7381;
assign w7383 = ~w7379 & w7382;
assign w7384 = ~pi0446 & w1867;
assign w7385 = ~pi0577 & w1862;
assign w7386 = ~pi0399 & w1813;
assign w7387 = pi0846 & w1860;
assign w7388 = ~pi0687 & w1865;
assign w7389 = ~w7384 & ~w7386;
assign w7390 = ~w7385 & w7389;
assign w7391 = ~w7387 & w7390;
assign w7392 = ~w7388 & w7391;
assign w7393 = ~pi0496 & w1867;
assign w7394 = ~pi0540 & w1862;
assign w7395 = ~pi0397 & w1813;
assign w7396 = pi0847 & w1860;
assign w7397 = ~pi0688 & w1865;
assign w7398 = ~w7393 & ~w7395;
assign w7399 = ~w7394 & w7398;
assign w7400 = ~w7396 & w7399;
assign w7401 = ~w7397 & w7400;
assign w7402 = ~pi0498 & w1867;
assign w7403 = ~pi0579 & w1862;
assign w7404 = ~pi0401 & w1813;
assign w7405 = ~pi0690 & w1865;
assign w7406 = pi0848 & w1860;
assign w7407 = ~w7402 & ~w7404;
assign w7408 = ~w7403 & w7407;
assign w7409 = ~w7405 & w7408;
assign w7410 = ~w7406 & w7409;
assign w7411 = ~pi0445 & w1867;
assign w7412 = ~pi0539 & w1862;
assign w7413 = ~pi0400 & w1813;
assign w7414 = pi0849 & w1860;
assign w7415 = ~pi0689 & w1865;
assign w7416 = ~w7411 & ~w7413;
assign w7417 = ~w7412 & w7416;
assign w7418 = ~w7414 & w7417;
assign w7419 = ~w7415 & w7418;
assign w7420 = ~pi0406 & w1867;
assign w7421 = ~pi0504 & w1862;
assign w7422 = ~pi0334 & w1813;
assign w7423 = ~pi0651 & w1865;
assign w7424 = pi0850 & w1860;
assign w7425 = ~w7420 & ~w7422;
assign w7426 = ~w7421 & w7425;
assign w7427 = ~w7423 & w7426;
assign w7428 = ~w7424 & w7427;
assign w7429 = ~pi0499 & w1867;
assign w7430 = ~pi0582 & w1862;
assign w7431 = ~pi0402 & w1813;
assign w7432 = ~pi0692 & w1865;
assign w7433 = ~pi0851 & w1860;
assign w7434 = ~w7429 & ~w7431;
assign w7435 = ~w7430 & w7434;
assign w7436 = ~w7432 & w7435;
assign w7437 = ~w7433 & w7436;
assign w7438 = ~pi0500 & w1867;
assign w7439 = ~pi0583 & w1862;
assign w7440 = ~pi0403 & w1813;
assign w7441 = pi0852 & w1860;
assign w7442 = ~pi0691 & w1865;
assign w7443 = ~w7438 & ~w7440;
assign w7444 = ~w7439 & w7443;
assign w7445 = ~w7441 & w7444;
assign w7446 = ~w7442 & w7445;
assign w7447 = ~pi0407 & w1867;
assign w7448 = ~pi0505 & w1862;
assign w7449 = ~pi0335 & w1813;
assign w7450 = ~pi0853 & w1860;
assign w7451 = ~pi0652 & w1865;
assign w7452 = ~w7447 & ~w7449;
assign w7453 = ~w7448 & w7452;
assign w7454 = ~w7450 & w7453;
assign w7455 = ~w7451 & w7454;
assign w7456 = ~pi0374 & w1867;
assign w7457 = ~pi0462 & w1862;
assign w7458 = ~pi0328 & w1813;
assign w7459 = ~pi0854 & w1860;
assign w7460 = ~pi0641 & w1865;
assign w7461 = ~w7456 & ~w7458;
assign w7462 = ~w7457 & w7461;
assign w7463 = ~w7459 & w7462;
assign w7464 = ~w7460 & w7463;
assign w7465 = ~pi0376 & w1867;
assign w7466 = ~pi0463 & w1862;
assign w7467 = ~pi0329 & w1813;
assign w7468 = ~pi0628 & w1865;
assign w7469 = ~pi0855 & w1860;
assign w7470 = ~w7465 & ~w7467;
assign w7471 = ~w7466 & w7470;
assign w7472 = ~w7468 & w7471;
assign w7473 = ~w7469 & w7472;
assign w7474 = ~pi0357 & w1867;
assign w7475 = ~pi0461 & w1862;
assign w7476 = ~pi0327 & w1813;
assign w7477 = ~pi0633 & w1865;
assign w7478 = ~pi0856 & w1860;
assign w7479 = ~w7474 & ~w7476;
assign w7480 = ~w7475 & w7479;
assign w7481 = ~w7477 & w7480;
assign w7482 = ~w7478 & w7481;
assign w7483 = ~pi0503 & w1867;
assign w7484 = ~pi0584 & w1862;
assign w7485 = ~pi0404 & w1813;
assign w7486 = ~pi0694 & w1865;
assign w7487 = ~pi0857 & w1860;
assign w7488 = ~w7483 & ~w7485;
assign w7489 = ~w7484 & w7488;
assign w7490 = ~w7486 & w7489;
assign w7491 = ~w7487 & w7490;
assign w7492 = ~pi0443 & w1867;
assign w7493 = ~pi0585 & w1862;
assign w7494 = ~pi0405 & w1813;
assign w7495 = ~pi0693 & w1865;
assign w7496 = ~pi0858 & w1860;
assign w7497 = ~w7492 & ~w7494;
assign w7498 = ~w7493 & w7497;
assign w7499 = ~w7495 & w7498;
assign w7500 = ~w7496 & w7499;
assign w7501 = ~pi1126 & w1867;
assign w7502 = ~pi1031 & w1862;
assign w7503 = ~pi1235 & w1813;
assign w7504 = pi0859 & w1860;
assign w7505 = ~pi1237 & w1865;
assign w7506 = ~w7501 & ~w7503;
assign w7507 = ~w7502 & w7506;
assign w7508 = ~w7504 & w7507;
assign w7509 = ~w7505 & w7508;
assign w7510 = ~pi1128 & w1867;
assign w7511 = ~pi1273 & w1862;
assign w7512 = ~pi1268 & w1813;
assign w7513 = pi0860 & w1860;
assign w7514 = ~pi1243 & w1865;
assign w7515 = ~w7510 & ~w7512;
assign w7516 = ~w7511 & w7515;
assign w7517 = ~w7513 & w7516;
assign w7518 = ~w7514 & w7517;
assign w7519 = pi1430 & pi1698;
assign w7520 = pi1747 & ~w7519;
assign w7521 = pi0861 & w7520;
assign w7522 = pi1698 & pi1747;
assign w7523 = pi0064 & w7522;
assign w7524 = pi1430 & w7523;
assign w7525 = ~w7521 & ~w7524;
assign w7526 = pi0862 & w7520;
assign w7527 = pi0057 & w7522;
assign w7528 = pi1430 & w7527;
assign w7529 = ~w7526 & ~w7528;
assign w7530 = pi1430 & pi1695;
assign w7531 = pi1747 & ~w7530;
assign w7532 = pi0863 & w7531;
assign w7533 = pi0056 & pi1695;
assign w7534 = pi1747 & w7533;
assign w7535 = pi1430 & w7534;
assign w7536 = ~w7532 & ~w7535;
assign w7537 = ~pi0363 & w1867;
assign w7538 = ~pi0452 & w1862;
assign w7539 = ~pi0315 & w1813;
assign w7540 = ~pi0553 & w1865;
assign w7541 = ~pi0870 & w1860;
assign w7542 = ~w7537 & ~w7539;
assign w7543 = ~w7538 & w7542;
assign w7544 = ~w7540 & w7543;
assign w7545 = ~w7541 & w7544;
assign w7546 = ~pi0415 & w1867;
assign w7547 = ~pi0523 & w1862;
assign w7548 = ~pi0338 & w1813;
assign w7549 = pi0871 & w1860;
assign w7550 = ~pi0597 & w1865;
assign w7551 = ~w7546 & ~w7548;
assign w7552 = ~w7547 & w7551;
assign w7553 = ~w7549 & w7552;
assign w7554 = ~w7550 & w7553;
assign w7555 = ~pi0764 & ~w6894;
assign w7556 = pi0790 & ~w7555;
assign w7557 = pi0765 & ~w7556;
assign w7558 = pi0766 & ~w7557;
assign w7559 = w6406 & ~w7558;
assign w7560 = ~pi1078 & w1867;
assign w7561 = pi1145 & w1862;
assign w7562 = pi1024 & w1813;
assign w7563 = ~pi0873 & w1860;
assign w7564 = pi1114 & w1865;
assign w7565 = ~w7560 & ~w7562;
assign w7566 = ~w7561 & w7565;
assign w7567 = ~w7563 & w7566;
assign w7568 = ~w7564 & w7567;
assign w7569 = pi0876 & w7531;
assign w7570 = pi0049 & pi1695;
assign w7571 = pi1747 & w7570;
assign w7572 = pi1430 & w7571;
assign w7573 = ~w7569 & ~w7572;
assign w7574 = pi1127 & w1867;
assign w7575 = pi1139 & w1862;
assign w7576 = pi1119 & w1813;
assign w7577 = pi0877 & w1860;
assign w7578 = pi1102 & w1865;
assign w7579 = ~w7574 & ~w7576;
assign w7580 = ~w7575 & w7579;
assign w7581 = ~w7577 & w7580;
assign w7582 = ~w7578 & w7581;
assign w7583 = ~pi0051 & ~w624;
assign w7584 = pi0878 & w624;
assign w7585 = ~w634 & ~w7583;
assign w7586 = ~w7584 & w7585;
assign w7587 = ~pi0375 & w1867;
assign w7588 = ~pi0464 & w1862;
assign w7589 = ~pi0330 & w1813;
assign w7590 = ~pi0879 & w1860;
assign w7591 = ~pi0624 & w1865;
assign w7592 = ~w7587 & ~w7589;
assign w7593 = ~w7588 & w7592;
assign w7594 = ~w7590 & w7593;
assign w7595 = ~w7591 & w7594;
assign w7596 = ~pi0502 & w1867;
assign w7597 = ~pi0537 & w1862;
assign w7598 = ~pi0360 & w1813;
assign w7599 = ~pi0703 & w1865;
assign w7600 = ~pi0880 & w1860;
assign w7601 = ~w7596 & ~w7598;
assign w7602 = ~w7597 & w7601;
assign w7603 = ~w7599 & w7602;
assign w7604 = ~w7600 & w7603;
assign w7605 = pi0881 & ~w5585;
assign w7606 = pi0918 & w5585;
assign w7607 = ~w7605 & ~w7606;
assign w7608 = ~pi1300 & ~pi1773;
assign w7609 = pi1773 & ~pi1831;
assign w7610 = ~w7608 & ~w7609;
assign w7611 = pi0469 & w6633;
assign w7612 = ~pi0593 & w4056;
assign w7613 = ~pi0337 & w2866;
assign w7614 = pi0535 & w6609;
assign w7615 = ~pi1126 & w6627;
assign w7616 = pi1291 & w6615;
assign w7617 = ~pi0487 & w3188;
assign w7618 = ~pi0520 & w3953;
assign w7619 = ~pi1237 & w6612;
assign w7620 = ~pi0570 & w4186;
assign w7621 = ~pi0389 & w2932;
assign w7622 = pi0617 & w6618;
assign w7623 = ~pi0670 & w5442;
assign w7624 = pi0592 & w6629;
assign w7625 = ~pi0612 & w3150;
assign w7626 = pi0615 & w6624;
assign w7627 = pi1687 & w6641;
assign w7628 = ~pi1235 & w6620;
assign w7629 = ~pi1031 & w6622;
assign w7630 = pi1503 & w6637;
assign w7631 = pi1038 & w6606;
assign w7632 = pi1094 & w6639;
assign w7633 = ~w7612 & ~w7613;
assign w7634 = ~w7614 & ~w7615;
assign w7635 = ~w7617 & ~w7618;
assign w7636 = ~w7619 & ~w7620;
assign w7637 = ~w7621 & ~w7622;
assign w7638 = ~w7623 & ~w7624;
assign w7639 = ~w7625 & ~w7626;
assign w7640 = ~w7628 & ~w7629;
assign w7641 = w7639 & w7640;
assign w7642 = w7637 & w7638;
assign w7643 = w7635 & w7636;
assign w7644 = w7633 & w7634;
assign w7645 = ~w7611 & ~w7616;
assign w7646 = ~w7627 & ~w7630;
assign w7647 = ~w7631 & ~w7632;
assign w7648 = w7646 & w7647;
assign w7649 = w7644 & w7645;
assign w7650 = w7642 & w7643;
assign w7651 = w7641 & w7650;
assign w7652 = w7648 & w7649;
assign w7653 = w7651 & w7652;
assign w7654 = pi0884 & ~w5585;
assign w7655 = pi0887 & w5585;
assign w7656 = ~w7654 & ~w7655;
assign w7657 = pi0433 & w6633;
assign w7658 = pi1105 & w6612;
assign w7659 = ~pi0607 & w4056;
assign w7660 = ~pi0582 & w4186;
assign w7661 = pi0116 & w6624;
assign w7662 = pi1289 & w6615;
assign w7663 = pi1022 & w6620;
assign w7664 = ~pi0534 & w3150;
assign w7665 = ~pi0402 & w2932;
assign w7666 = pi1032 & w6622;
assign w7667 = pi1027 & w6627;
assign w7668 = ~pi0435 & w2866;
assign w7669 = ~pi0626 & w3953;
assign w7670 = ~pi0692 & w5442;
assign w7671 = ~pi0499 & w3188;
assign w7672 = pi0114 & w6629;
assign w7673 = pi1682 & w6641;
assign w7674 = pi0118 & w6618;
assign w7675 = pi0115 & w6609;
assign w7676 = pi1505 & w6637;
assign w7677 = pi1457 & w6606;
assign w7678 = pi1096 & w6639;
assign w7679 = ~w7658 & ~w7659;
assign w7680 = ~w7660 & ~w7661;
assign w7681 = ~w7663 & ~w7664;
assign w7682 = ~w7665 & ~w7666;
assign w7683 = ~w7667 & ~w7668;
assign w7684 = ~w7669 & ~w7670;
assign w7685 = ~w7671 & ~w7672;
assign w7686 = ~w7674 & ~w7675;
assign w7687 = w7685 & w7686;
assign w7688 = w7683 & w7684;
assign w7689 = w7681 & w7682;
assign w7690 = w7679 & w7680;
assign w7691 = ~w7657 & ~w7662;
assign w7692 = ~w7673 & ~w7676;
assign w7693 = ~w7677 & ~w7678;
assign w7694 = w7692 & w7693;
assign w7695 = w7690 & w7691;
assign w7696 = w7688 & w7689;
assign w7697 = w7687 & w7696;
assign w7698 = w7694 & w7695;
assign w7699 = w7697 & w7698;
assign w7700 = pi0475 & w6633;
assign w7701 = pi0958 & w6624;
assign w7702 = pi1310 & w6627;
assign w7703 = pi0959 & w6618;
assign w7704 = ~pi0502 & w3188;
assign w7705 = pi1069 & w6639;
assign w7706 = ~pi0425 & w3150;
assign w7707 = ~pi0609 & w4056;
assign w7708 = ~pi0531 & w3953;
assign w7709 = pi0970 & w6629;
assign w7710 = pi1277 & w6620;
assign w7711 = ~pi0537 & w4186;
assign w7712 = pi0957 & w6609;
assign w7713 = pi1342 & w6622;
assign w7714 = pi1338 & w6612;
assign w7715 = ~pi0348 & w2866;
assign w7716 = pi1504 & w6637;
assign w7717 = ~pi0703 & w5442;
assign w7718 = ~pi0360 & w2932;
assign w7719 = pi1700 & w6641;
assign w7720 = pi1320 & w6615;
assign w7721 = pi1731 & w6606;
assign w7722 = ~w7701 & ~w7702;
assign w7723 = ~w7703 & ~w7704;
assign w7724 = ~w7706 & ~w7707;
assign w7725 = ~w7708 & ~w7709;
assign w7726 = ~w7710 & ~w7711;
assign w7727 = ~w7712 & ~w7713;
assign w7728 = ~w7714 & ~w7715;
assign w7729 = ~w7717 & ~w7718;
assign w7730 = w7728 & w7729;
assign w7731 = w7726 & w7727;
assign w7732 = w7724 & w7725;
assign w7733 = w7722 & w7723;
assign w7734 = ~w7700 & ~w7705;
assign w7735 = ~w7716 & ~w7719;
assign w7736 = ~w7720 & ~w7721;
assign w7737 = w7735 & w7736;
assign w7738 = w7733 & w7734;
assign w7739 = w7731 & w7732;
assign w7740 = w7730 & w7739;
assign w7741 = w7737 & w7738;
assign w7742 = w7740 & w7741;
assign w7743 = pi0887 & ~w5585;
assign w7744 = pi1740 & w5585;
assign w7745 = ~w7743 & ~w7744;
assign w7746 = ~pi1301 & ~pi1773;
assign w7747 = pi1773 & ~pi1832;
assign w7748 = ~w7746 & ~w7747;
assign w7749 = pi0889 & ~w5585;
assign w7750 = pi1741 & w5585;
assign w7751 = ~w7749 & ~w7750;
assign w7752 = pi0890 & ~w5585;
assign w7753 = pi1727 & w5585;
assign w7754 = ~w7752 & ~w7753;
assign w7755 = pi0012 & pi0095;
assign w7756 = pi1510 & w7755;
assign w7757 = ~w397 & w7756;
assign w7758 = pi1447 & w7757;
assign w7759 = ~pi0891 & ~w7758;
assign w7760 = w1783 & ~w7759;
assign w7761 = pi1480 & w7757;
assign w7762 = ~pi0892 & ~w7761;
assign w7763 = w1773 & ~w7762;
assign w7764 = pi1233 & ~w1173;
assign w7765 = ~pi1494 & ~w406;
assign w7766 = pi0795 & pi1479;
assign w7767 = pi0771 & pi0799;
assign w7768 = w7766 & w7767;
assign w7769 = pi0803 & pi0860;
assign w7770 = pi0802 & w7769;
assign w7771 = w7768 & w7770;
assign w7772 = ~w370 & ~w7771;
assign w7773 = ~w7765 & ~w7772;
assign w7774 = pi0802 & pi0860;
assign w7775 = w1212 & w5455;
assign w7776 = w7768 & w7775;
assign w7777 = ~pi0803 & pi0860;
assign w7778 = pi0802 & ~w7777;
assign w7779 = ~pi0800 & w7766;
assign w7780 = ~w7769 & w7779;
assign w7781 = ~w7778 & w7780;
assign w7782 = pi0799 & ~w7781;
assign w7783 = w374 & ~w7782;
assign w7784 = pi0801 & ~w7783;
assign w7785 = ~pi0802 & ~w7767;
assign w7786 = ~w7784 & w7785;
assign w7787 = ~w7776 & ~w7786;
assign w7788 = ~w7774 & ~w7787;
assign w7789 = ~w7773 & ~w7788;
assign w7790 = ~pi1027 & ~pi1028;
assign w7791 = ~pi1029 & ~pi1076;
assign w7792 = ~pi1083 & ~pi1092;
assign w7793 = pi1126 & ~pi1127;
assign w7794 = ~pi1129 & ~pi1130;
assign w7795 = ~pi1310 & w7794;
assign w7796 = w7792 & w7793;
assign w7797 = w7790 & w7791;
assign w7798 = w7796 & w7797;
assign w7799 = w7795 & w7798;
assign w7800 = ~pi0380 & ~pi0468;
assign w7801 = ~w3534 & w7800;
assign w7802 = w4280 & w7801;
assign w7803 = ~w7799 & ~w7802;
assign w7804 = ~pi0379 & ~pi0381;
assign w7805 = ~pi0470 & w7804;
assign w7806 = ~w3475 & w7805;
assign w7807 = ~w3470 & w7806;
assign w7808 = ~pi1022 & ~pi1023;
assign w7809 = ~pi1119 & ~pi1121;
assign w7810 = pi1235 & ~pi1267;
assign w7811 = ~pi1270 & ~pi1272;
assign w7812 = ~pi1274 & ~pi1277;
assign w7813 = ~pi1280 & w7812;
assign w7814 = w7810 & w7811;
assign w7815 = w7808 & w7809;
assign w7816 = w7814 & w7815;
assign w7817 = w7813 & w7816;
assign w7818 = ~w7807 & ~w7817;
assign w7819 = ~pi1081 & ~pi1102;
assign w7820 = ~pi1104 & ~pi1105;
assign w7821 = ~pi1106 & ~pi1107;
assign w7822 = ~pi1108 & pi1237;
assign w7823 = ~pi1338 & w7822;
assign w7824 = w7820 & w7821;
assign w7825 = w5722 & w7819;
assign w7826 = w7824 & w7825;
assign w7827 = w7823 & w7826;
assign w7828 = ~pi0665 & w5764;
assign w7829 = ~w3290 & w7828;
assign w7830 = ~w3289 & w7829;
assign w7831 = ~w7827 & ~w7830;
assign w7832 = ~pi0621 & w5578;
assign w7833 = pi1031 & ~pi1032;
assign w7834 = ~pi1033 & ~pi1034;
assign w7835 = ~pi1139 & ~pi1141;
assign w7836 = ~pi1142 & ~pi1258;
assign w7837 = ~pi1265 & ~pi1271;
assign w7838 = ~pi1342 & w7837;
assign w7839 = w7835 & w7836;
assign w7840 = w7833 & w7834;
assign w7841 = w7839 & w7840;
assign w7842 = w7838 & w7841;
assign w7843 = ~w7832 & ~w7842;
assign w7844 = pi0966 & w2132;
assign w7845 = ~w6720 & ~w7844;
assign w7846 = ~pi1479 & ~w6720;
assign w7847 = ~w7845 & ~w7846;
assign w7848 = ~pi0954 & pi1021;
assign w7849 = w2169 & w7848;
assign w7850 = ~w2174 & ~w7849;
assign w7851 = ~pi1019 & w2179;
assign w7852 = pi0262 & pi1019;
assign w7853 = ~pi0916 & w7852;
assign w7854 = ~pi0900 & ~w7853;
assign w7855 = ~w7851 & w7854;
assign w7856 = ~w2171 & w7855;
assign w7857 = w7850 & w7856;
assign w7858 = ~w7847 & ~w7857;
assign w7859 = ~pi1676 & ~pi1726;
assign w7860 = ~pi0901 & ~w7859;
assign w7861 = w1885 & ~w7860;
assign w7862 = ~pi1286 & ~pi1773;
assign w7863 = pi1773 & ~pi1810;
assign w7864 = ~w7862 & ~w7863;
assign w7865 = pi1459 & w7757;
assign w7866 = ~pi0903 & ~w7865;
assign w7867 = w1769 & ~w7866;
assign w7868 = pi1430 & w7757;
assign w7869 = ~pi0904 & ~w7868;
assign w7870 = w1777 & ~w7869;
assign w7871 = ~pi1294 & ~pi1773;
assign w7872 = pi1773 & ~pi1822;
assign w7873 = ~w7871 & ~w7872;
assign w7874 = ~pi1299 & ~pi1773;
assign w7875 = pi1773 & ~pi1830;
assign w7876 = ~w7874 & ~w7875;
assign w7877 = ~pi1302 & ~pi1773;
assign w7878 = pi1773 & ~pi1834;
assign w7879 = ~w7877 & ~w7878;
assign w7880 = ~pi1298 & ~pi1773;
assign w7881 = pi1773 & ~pi1827;
assign w7882 = ~w7880 & ~w7881;
assign w7883 = ~pi1293 & ~pi1773;
assign w7884 = pi1773 & ~pi1826;
assign w7885 = ~w7883 & ~w7884;
assign w7886 = ~pi1297 & ~pi1773;
assign w7887 = pi1773 & ~pi1825;
assign w7888 = ~w7886 & ~w7887;
assign w7889 = ~pi1304 & ~pi1773;
assign w7890 = pi1773 & ~pi1812;
assign w7891 = ~w7889 & ~w7890;
assign w7892 = ~pi1303 & ~pi1773;
assign w7893 = pi1773 & ~pi1811;
assign w7894 = ~w7892 & ~w7893;
assign w7895 = ~pi1296 & ~pi1773;
assign w7896 = pi1773 & ~pi1824;
assign w7897 = ~w7895 & ~w7896;
assign w7898 = ~pi1295 & ~pi1773;
assign w7899 = pi1773 & ~pi1823;
assign w7900 = ~w7898 & ~w7899;
assign w7901 = ~pi1675 & ~pi1680;
assign w7902 = ~pi0915 & ~w7901;
assign w7903 = w1885 & ~w7902;
assign w7904 = w2147 & w6718;
assign w7905 = w2133 & w6720;
assign w7906 = ~pi0785 & w2154;
assign w7907 = ~w2157 & w7906;
assign w7908 = w2150 & w7907;
assign w7909 = pi0995 & w2143;
assign w7910 = pi0276 & w7909;
assign w7911 = ~pi0183 & w6405;
assign w7912 = ~w7905 & ~w7908;
assign w7913 = ~w7911 & w7912;
assign w7914 = ~w7849 & w7913;
assign w7915 = ~w7910 & w7914;
assign w7916 = w7904 & ~w7915;
assign w7917 = ~pi0917 & ~w1232;
assign w7918 = ~w5585 & ~w7917;
assign w7919 = pi1747 & ~w7918;
assign w7920 = pi0918 & ~w5585;
assign w7921 = pi1733 & w5585;
assign w7922 = ~w7920 & ~w7921;
assign w7923 = pi0937 & ~w6397;
assign w7924 = ~w6809 & ~w7923;
assign w7925 = w6811 & w7924;
assign w7926 = ~pi0963 & w7925;
assign w7927 = ~pi0919 & w7926;
assign w7928 = ~pi0919 & ~pi0984;
assign w7929 = ~w7926 & ~w7928;
assign w7930 = ~w7927 & ~w7929;
assign w7931 = pi0920 & ~w5585;
assign w7932 = pi1722 & w5585;
assign w7933 = ~w7931 & ~w7932;
assign w7934 = ~pi0921 & ~pi0984;
assign w7935 = ~w7927 & ~w7934;
assign w7936 = ~pi0921 & w7927;
assign w7937 = ~w7935 & ~w7936;
assign w7938 = pi0922 & ~w5585;
assign w7939 = pi1735 & w5585;
assign w7940 = ~w7938 & ~w7939;
assign w7941 = pi0923 & ~w5585;
assign w7942 = ~w6386 & ~w7941;
assign w7943 = pi0924 & ~w5585;
assign w7944 = pi1725 & w5585;
assign w7945 = ~w7943 & ~w7944;
assign w7946 = pi0925 & ~w5585;
assign w7947 = pi0889 & w5585;
assign w7948 = ~w7946 & ~w7947;
assign w7949 = pi0926 & ~w5585;
assign w7950 = pi0920 & w5585;
assign w7951 = ~w7949 & ~w7950;
assign w7952 = pi0927 & ~w5585;
assign w7953 = pi0890 & w5585;
assign w7954 = ~w7952 & ~w7953;
assign w7955 = pi0928 & ~w5585;
assign w7956 = pi0922 & w5585;
assign w7957 = ~w7955 & ~w7956;
assign w7958 = pi0929 & ~w5585;
assign w7959 = pi0923 & w5585;
assign w7960 = ~w7958 & ~w7959;
assign w7961 = pi0930 & ~w5585;
assign w7962 = pi0924 & w5585;
assign w7963 = ~w7961 & ~w7962;
assign w7964 = pi0931 & ~w5585;
assign w7965 = pi0925 & w5585;
assign w7966 = ~w7964 & ~w7965;
assign w7967 = pi0932 & ~w5585;
assign w7968 = pi0926 & w5585;
assign w7969 = ~w7967 & ~w7968;
assign w7970 = pi0933 & ~w5585;
assign w7971 = pi0927 & w5585;
assign w7972 = ~w7970 & ~w7971;
assign w7973 = pi0934 & ~w5585;
assign w7974 = pi0928 & w5585;
assign w7975 = ~w7973 & ~w7974;
assign w7976 = pi0935 & ~w5585;
assign w7977 = pi0929 & w5585;
assign w7978 = ~w7976 & ~w7977;
assign w7979 = pi0936 & ~w5585;
assign w7980 = pi0930 & w5585;
assign w7981 = ~w7979 & ~w7980;
assign w7982 = w6718 & w6810;
assign w7983 = w6812 & w7982;
assign w7984 = pi1447 & w7523;
assign w7985 = pi1447 & pi1698;
assign w7986 = pi1747 & ~w7985;
assign w7987 = pi0938 & w7986;
assign w7988 = ~w7984 & ~w7987;
assign w7989 = pi1447 & pi1695;
assign w7990 = pi1747 & ~w7989;
assign w7991 = pi0939 & w7990;
assign w7992 = pi1447 & w7534;
assign w7993 = ~w7991 & ~w7992;
assign w7994 = pi1447 & w7527;
assign w7995 = pi0941 & w7986;
assign w7996 = ~w7994 & ~w7995;
assign w7997 = pi0942 & w7990;
assign w7998 = pi1447 & w7571;
assign w7999 = ~w7997 & ~w7998;
assign w8000 = pi0943 & ~w5585;
assign w8001 = pi0881 & w5585;
assign w8002 = ~w8000 & ~w8001;
assign w8003 = pi0944 & ~w5585;
assign w8004 = pi0884 & w5585;
assign w8005 = ~w8003 & ~w8004;
assign w8006 = ~pi0715 & pi1269;
assign w8007 = pi0715 & ~pi1269;
assign w8008 = ~w8006 & ~w8007;
assign w8009 = ~pi0663 & pi1159;
assign w8010 = ~pi0709 & pi1346;
assign w8011 = pi0720 & ~pi1158;
assign w8012 = ~pi0720 & pi1158;
assign w8013 = ~w8011 & ~w8012;
assign w8014 = pi0679 & ~pi1275;
assign w8015 = ~pi0679 & pi1275;
assign w8016 = ~w8014 & ~w8015;
assign w8017 = pi0707 & ~pi1157;
assign w8018 = ~pi0707 & pi1157;
assign w8019 = ~w8017 & ~w8018;
assign w8020 = pi0710 & ~pi1156;
assign w8021 = ~pi0710 & pi1156;
assign w8022 = ~w8020 & ~w8021;
assign w8023 = ~pi0669 & pi1155;
assign w8024 = ~pi0698 & pi1283;
assign w8025 = pi0698 & ~pi1283;
assign w8026 = pi0700 & ~pi1331;
assign w8027 = ~w8025 & ~w8026;
assign w8028 = (~pi0699 & w8027) | (~pi0699 & w12978) | (w8027 & w12978);
assign w8029 = ~w8027 & w12967;
assign w8030 = pi1154 & ~w8029;
assign w8031 = ~w8028 & ~w8030;
assign w8032 = pi0669 & ~pi1155;
assign w8033 = ~w8023 & ~w8032;
assign w8034 = (w8033 & w8030) | (w8033 & w12979) | (w8030 & w12979);
assign w8035 = ~w8023 & ~w8034;
assign w8036 = ~w8034 & w12994;
assign w8037 = ~w8020 & ~w8036;
assign w8038 = w8019 & ~w8037;
assign w8039 = ~w8017 & ~w8038;
assign w8040 = w8016 & ~w8039;
assign w8041 = ~w8014 & ~w8040;
assign w8042 = w8013 & ~w8041;
assign w8043 = pi0709 & ~pi1346;
assign w8044 = ~w8011 & ~w8043;
assign w8045 = ~w8042 & w8044;
assign w8046 = ~w8010 & ~w8045;
assign w8047 = pi0663 & ~pi1159;
assign w8048 = ~w8009 & ~w8047;
assign w8049 = ~w8046 & w8048;
assign w8050 = ~w8009 & ~w8049;
assign w8051 = w8008 & w8050;
assign w8052 = ~w8008 & ~w8050;
assign w8053 = ~w8051 & ~w8052;
assign w8054 = ~pi0441 & pi1176;
assign w8055 = pi0482 & ~pi1089;
assign w8056 = ~pi0482 & pi1089;
assign w8057 = ~w8055 & ~w8056;
assign w8058 = pi0388 & ~pi1175;
assign w8059 = ~pi0388 & pi1175;
assign w8060 = ~w8058 & ~w8059;
assign w8061 = ~pi0510 & pi1093;
assign w8062 = pi0510 & ~pi1093;
assign w8063 = ~w8061 & ~w8062;
assign w8064 = ~pi0442 & pi1174;
assign w8065 = ~pi0413 & pi1087;
assign w8066 = pi0413 & ~pi1087;
assign w8067 = ~w8065 & ~w8066;
assign w8068 = ~pi0412 & pi1173;
assign w8069 = pi0412 & ~pi1173;
assign w8070 = ~pi0411 & pi1077;
assign w8071 = pi0411 & ~pi1077;
assign w8072 = pi0410 & ~pi1241;
assign w8073 = ~w8071 & ~w8072;
assign w8074 = ~w8070 & ~w8073;
assign w8075 = (~w8069 & w8073) | (~w8069 & w12968) | (w8073 & w12968);
assign w8076 = ~w8068 & ~w8075;
assign w8077 = w8067 & ~w8076;
assign w8078 = ~w8065 & ~w8077;
assign w8079 = pi0442 & ~pi1174;
assign w8080 = ~w8064 & ~w8079;
assign w8081 = ~w8078 & w8080;
assign w8082 = ~w8064 & ~w8081;
assign w8083 = w8063 & ~w8082;
assign w8084 = ~w8061 & ~w8083;
assign w8085 = w8060 & w8084;
assign w8086 = ~w8058 & ~w8085;
assign w8087 = w8057 & ~w8086;
assign w8088 = pi0441 & ~pi1176;
assign w8089 = ~w8055 & ~w8088;
assign w8090 = ~w8087 & w8089;
assign w8091 = ~w8054 & ~w8090;
assign w8092 = pi0384 & ~pi1082;
assign w8093 = ~w8091 & ~w8092;
assign w8094 = ~pi0384 & pi1082;
assign w8095 = ~pi0481 & pi1177;
assign w8096 = pi0481 & ~pi1177;
assign w8097 = ~w8095 & ~w8096;
assign w8098 = ~w8094 & w8097;
assign w8099 = ~w8093 & w8098;
assign w8100 = ~w8092 & ~w8094;
assign w8101 = w8091 & w8100;
assign w8102 = ~w8092 & ~w8097;
assign w8103 = ~w8101 & w8102;
assign w8104 = ~w8099 & ~w8103;
assign w8105 = pi0564 & ~pi1201;
assign w8106 = ~pi0564 & pi1201;
assign w8107 = ~w8105 & ~w8106;
assign w8108 = pi0472 & ~pi1249;
assign w8109 = pi0565 & ~pi1198;
assign w8110 = ~pi0565 & pi1198;
assign w8111 = ~w8109 & ~w8110;
assign w8112 = pi0486 & ~pi1197;
assign w8113 = ~pi0486 & pi1197;
assign w8114 = ~w8112 & ~w8113;
assign w8115 = ~pi0588 & pi1264;
assign w8116 = pi0588 & ~pi1264;
assign w8117 = ~w8115 & ~w8116;
assign w8118 = ~pi0541 & pi1196;
assign w8119 = ~pi0514 & pi1195;
assign w8120 = pi0514 & ~pi1195;
assign w8121 = ~w8119 & ~w8120;
assign w8122 = ~pi0513 & pi1194;
assign w8123 = pi0513 & ~pi1194;
assign w8124 = ~pi0512 & pi1276;
assign w8125 = pi0512 & ~pi1276;
assign w8126 = pi0511 & ~pi1192;
assign w8127 = ~w8125 & ~w8126;
assign w8128 = ~w8124 & ~w8127;
assign w8129 = (~w8123 & w8127) | (~w8123 & w12969) | (w8127 & w12969);
assign w8130 = ~w8122 & ~w8129;
assign w8131 = (w8121 & w8129) | (w8121 & w12980) | (w8129 & w12980);
assign w8132 = ~w8119 & ~w8131;
assign w8133 = pi0541 & ~pi1196;
assign w8134 = ~w8118 & ~w8133;
assign w8135 = (w8134 & w8131) | (w8134 & w12981) | (w8131 & w12981);
assign w8136 = ~w8118 & ~w8135;
assign w8137 = w8117 & ~w8136;
assign w8138 = ~w8115 & ~w8137;
assign w8139 = w8114 & w8138;
assign w8140 = ~w8112 & ~w8139;
assign w8141 = w8111 & ~w8140;
assign w8142 = ~w8109 & ~w8141;
assign w8143 = ~pi1199 & ~w8142;
assign w8144 = pi1199 & ~w8109;
assign w8145 = ~w8141 & w8144;
assign w8146 = pi0560 & ~w8145;
assign w8147 = ~w8143 & ~w8146;
assign w8148 = ~pi0472 & pi1249;
assign w8149 = ~w8108 & ~w8148;
assign w8150 = ~w8147 & w8149;
assign w8151 = ~w8108 & ~w8150;
assign w8152 = w8107 & w8151;
assign w8153 = ~w8107 & ~w8151;
assign w8154 = ~w8152 & ~w8153;
assign w8155 = ~pi0649 & pi1232;
assign w8156 = pi0649 & ~pi1232;
assign w8157 = ~w8155 & ~w8156;
assign w8158 = ~pi0552 & pi1057;
assign w8159 = ~pi0642 & pi1056;
assign w8160 = pi0631 & ~pi1219;
assign w8161 = ~pi0631 & pi1219;
assign w8162 = ~w8160 & ~w8161;
assign w8163 = ~pi0655 & pi1217;
assign w8164 = pi0655 & ~pi1217;
assign w8165 = ~w8163 & ~w8164;
assign w8166 = ~pi0627 & pi1066;
assign w8167 = ~pi0591 & pi1216;
assign w8168 = pi0591 & ~pi1216;
assign w8169 = ~w8167 & ~w8168;
assign w8170 = ~pi0590 & pi1215;
assign w8171 = pi0590 & ~pi1215;
assign w8172 = ~pi0589 & pi1214;
assign w8173 = pi0589 & ~pi1214;
assign w8174 = pi0594 & ~pi1213;
assign w8175 = ~w8173 & ~w8174;
assign w8176 = ~w8172 & ~w8175;
assign w8177 = (~w8171 & w8175) | (~w8171 & w12970) | (w8175 & w12970);
assign w8178 = ~w8170 & ~w8177;
assign w8179 = (w8169 & w8177) | (w8169 & w12971) | (w8177 & w12971);
assign w8180 = ~w8167 & ~w8179;
assign w8181 = pi0627 & ~pi1066;
assign w8182 = ~w8166 & ~w8181;
assign w8183 = (w8182 & w8179) | (w8182 & w12982) | (w8179 & w12982);
assign w8184 = ~w8166 & ~w8183;
assign w8185 = w8165 & ~w8184;
assign w8186 = ~w8163 & ~w8185;
assign w8187 = ~pi0568 & ~w8186;
assign w8188 = pi0568 & w8186;
assign w8189 = pi1218 & ~w8188;
assign w8190 = ~w8187 & ~w8189;
assign w8191 = w8162 & w8190;
assign w8192 = pi0642 & ~pi1056;
assign w8193 = ~w8160 & ~w8192;
assign w8194 = ~w8191 & w8193;
assign w8195 = ~w8159 & ~w8194;
assign w8196 = pi0552 & ~pi1057;
assign w8197 = ~w8158 & ~w8196;
assign w8198 = ~w8195 & w8197;
assign w8199 = ~w8158 & ~w8198;
assign w8200 = w8157 & w8199;
assign w8201 = ~w8157 & ~w8199;
assign w8202 = ~w8200 & ~w8201;
assign w8203 = ~pi1366 & ~pi1773;
assign w8204 = pi1773 & ~pi1836;
assign w8205 = ~w8203 & ~w8204;
assign w8206 = ~pi1367 & ~pi1773;
assign w8207 = pi1773 & ~pi1837;
assign w8208 = ~w8206 & ~w8207;
assign w8209 = ~pi1099 & ~pi1358;
assign w8210 = ~pi0257 & pi1099;
assign w8211 = ~w8209 & ~w8210;
assign w8212 = ~pi0277 & w2171;
assign w8213 = w2161 & ~w8212;
assign w8214 = w6718 & ~w8213;
assign w8215 = ~pi1368 & ~pi1773;
assign w8216 = pi1773 & ~pi1833;
assign w8217 = ~w8215 & ~w8216;
assign w8218 = ~pi1365 & ~pi1773;
assign w8219 = pi1773 & ~pi1835;
assign w8220 = ~w8218 & ~w8219;
assign w8221 = ~pi1511 & w7755;
assign w8222 = w397 & w8221;
assign w8223 = pi1480 & w8222;
assign w8224 = ~pi0957 & ~w8223;
assign w8225 = w1773 & ~w8224;
assign w8226 = pi1430 & w8222;
assign w8227 = ~pi0958 & ~w8226;
assign w8228 = w1777 & ~w8227;
assign w8229 = pi1447 & w8222;
assign w8230 = ~pi0959 & ~w8229;
assign w8231 = w1783 & ~w8230;
assign w8232 = w6407 & ~w6891;
assign w8233 = w6406 & w8232;
assign w8234 = ~pi1372 & ~pi1773;
assign w8235 = pi1773 & ~pi1817;
assign w8236 = ~w8234 & ~w8235;
assign w8237 = ~pi1373 & ~pi1773;
assign w8238 = pi1773 & ~pi1815;
assign w8239 = ~w8237 & ~w8238;
assign w8240 = pi0963 & ~w7925;
assign w8241 = ~pi0984 & ~w7926;
assign w8242 = ~w8240 & w8241;
assign w8243 = ~pi1392 & ~pi1773;
assign w8244 = pi1773 & ~pi1818;
assign w8245 = ~w8243 & ~w8244;
assign w8246 = pi1430 & pi1729;
assign w8247 = ~pi0965 & ~w8246;
assign w8248 = w1777 & ~w8247;
assign w8249 = ~pi0984 & w6718;
assign w8250 = ~w2132 & w2176;
assign w8251 = w2145 & w6808;
assign w8252 = pi1045 & w6814;
assign w8253 = pi0277 & w8252;
assign w8254 = ~w8250 & ~w8253;
assign w8255 = ~w8251 & w8254;
assign w8256 = w8249 & ~w8255;
assign w8257 = pi1459 & w7523;
assign w8258 = pi1459 & pi1698;
assign w8259 = pi1747 & ~w8258;
assign w8260 = pi0967 & w8259;
assign w8261 = ~w8257 & ~w8260;
assign w8262 = pi1459 & w7527;
assign w8263 = pi0968 & w8259;
assign w8264 = ~w8262 & ~w8263;
assign w8265 = pi1459 & pi1695;
assign w8266 = pi1747 & ~w8265;
assign w8267 = pi0969 & w8266;
assign w8268 = pi1459 & w7534;
assign w8269 = ~w8267 & ~w8268;
assign w8270 = pi1459 & w8222;
assign w8271 = ~pi0970 & ~w8270;
assign w8272 = w1769 & ~w8271;
assign w8273 = ~pi0872 & ~pi1683;
assign w8274 = w6718 & ~w6808;
assign w8275 = ~w2134 & w8274;
assign w8276 = w2145 & w8275;
assign w8277 = ~w8273 & w8276;
assign w8278 = w6403 & w6718;
assign w8279 = ~w8277 & ~w8278;
assign w8280 = ~pi1371 & ~pi1773;
assign w8281 = pi1773 & ~pi1816;
assign w8282 = ~w8280 & ~w8281;
assign w8283 = pi0973 & w8266;
assign w8284 = pi1459 & w7571;
assign w8285 = ~w8283 & ~w8284;
assign w8286 = ~pi0789 & w5585;
assign w8287 = pi0975 & ~w7847;
assign w8288 = ~w2179 & ~w8287;
assign w8289 = w7850 & w8288;
assign w8290 = ~w2171 & ~w8289;
assign w8291 = ~w2171 & ~w7852;
assign w8292 = w7845 & ~w7849;
assign w8293 = pi0976 & w8292;
assign w8294 = w8291 & ~w8293;
assign w8295 = ~pi0977 & pi1543;
assign w8296 = w1885 & ~w8295;
assign w8297 = w8046 & ~w8048;
assign w8298 = ~w8049 & ~w8297;
assign w8299 = ~w8091 & ~w8100;
assign w8300 = ~w8101 & ~w8299;
assign w8301 = w8147 & ~w8149;
assign w8302 = ~w8150 & ~w8301;
assign w8303 = w8195 & ~w8197;
assign w8304 = ~w8198 & ~w8303;
assign w8305 = pi0802 & w7765;
assign w8306 = pi0803 & ~pi1494;
assign w8307 = w406 & w8306;
assign w8308 = ~w8305 & ~w8307;
assign w8309 = w370 & ~w8308;
assign w8310 = ~pi0860 & w1705;
assign w8311 = ~pi0802 & ~w8310;
assign w8312 = w7783 & ~w8311;
assign w8313 = ~pi0795 & ~pi0860;
assign w8314 = pi1479 & ~w8313;
assign w8315 = w7767 & ~w8314;
assign w8316 = ~pi1236 & w5455;
assign w8317 = w8315 & ~w8316;
assign w8318 = ~pi0799 & pi0802;
assign w8319 = pi0795 & w1705;
assign w8320 = ~w7769 & w8319;
assign w8321 = ~w8318 & ~w8320;
assign w8322 = w376 & ~w8315;
assign w8323 = ~w8321 & w8322;
assign w8324 = ~w8317 & ~w8323;
assign w8325 = ~w8309 & w8324;
assign w8326 = ~w8312 & w8325;
assign w8327 = pi0802 & w7776;
assign w8328 = w1705 & w8312;
assign w8329 = ~w8327 & ~w8328;
assign w8330 = w7777 & ~w8329;
assign w8331 = w7772 & ~w8330;
assign w8332 = ~w8307 & ~w8331;
assign w8333 = ~pi0278 & w6815;
assign w8334 = ~w2172 & ~w8333;
assign w8335 = w6806 & ~w8334;
assign w8336 = pi0985 & w8291;
assign w8337 = w8292 & w8336;
assign w8338 = ~pi0986 & pi1548;
assign w8339 = w1885 & ~w8338;
assign w8340 = ~pi0987 & pi1523;
assign w8341 = w1885 & ~w8340;
assign w8342 = ~pi1414 & ~pi1773;
assign w8343 = pi1773 & ~pi1819;
assign w8344 = ~w8342 & ~w8343;
assign w8345 = ~pi1415 & ~pi1773;
assign w8346 = pi1773 & ~pi1821;
assign w8347 = ~w8345 & ~w8346;
assign w8348 = pi1447 & pi1729;
assign w8349 = ~pi0990 & ~w8348;
assign w8350 = w1783 & ~w8349;
assign w8351 = pi1430 & w1248;
assign w8352 = ~pi0991 & ~w8351;
assign w8353 = w1777 & ~w8352;
assign w8354 = pi1480 & w7523;
assign w8355 = pi1480 & pi1698;
assign w8356 = pi1747 & ~w8355;
assign w8357 = pi0992 & w8356;
assign w8358 = ~w8354 & ~w8357;
assign w8359 = pi1480 & w7527;
assign w8360 = pi0993 & w8356;
assign w8361 = ~w8359 & ~w8360;
assign w8362 = pi1480 & pi1695;
assign w8363 = pi1747 & ~w8362;
assign w8364 = pi0994 & w8363;
assign w8365 = pi1480 & w7534;
assign w8366 = ~w8364 & ~w8365;
assign w8367 = ~pi0276 & w7909;
assign w8368 = ~w2177 & ~w8367;
assign w8369 = w7904 & ~w8368;
assign w8370 = w397 & w1007;
assign w8371 = pi0811 & ~w397;
assign w8372 = pi0835 & w397;
assign w8373 = ~w8371 & ~w8372;
assign w8374 = pi0820 & ~w397;
assign w8375 = pi0843 & w397;
assign w8376 = ~w8374 & ~w8375;
assign w8377 = pi0828 & ~w397;
assign w8378 = pi0851 & w397;
assign w8379 = ~w8377 & ~w8378;
assign w8380 = pi0814 & ~w397;
assign w8381 = pi0837 & w397;
assign w8382 = ~w8380 & ~w8381;
assign w8383 = pi0815 & ~w397;
assign w8384 = pi0838 & w397;
assign w8385 = ~w8383 & ~w8384;
assign w8386 = pi0870 & ~w397;
assign w8387 = pi0752 & w397;
assign w8388 = ~w8386 & ~w8387;
assign w8389 = pi0816 & ~w397;
assign w8390 = pi0839 & w397;
assign w8391 = ~w8389 & ~w8390;
assign w8392 = pi0817 & ~w397;
assign w8393 = pi0840 & w397;
assign w8394 = ~w8392 & ~w8393;
assign w8395 = pi0756 & ~w397;
assign w8396 = pi0880 & w397;
assign w8397 = ~w8395 & ~w8396;
assign w8398 = pi0830 & ~w397;
assign w8399 = pi0854 & w397;
assign w8400 = ~w8398 & ~w8399;
assign w8401 = pi0831 & ~w397;
assign w8402 = pi0855 & w397;
assign w8403 = ~w8401 & ~w8402;
assign w8404 = pi0832 & ~w397;
assign w8405 = pi0856 & w397;
assign w8406 = ~w8404 & ~w8405;
assign w8407 = pi0757 & ~w397;
assign w8408 = pi0879 & w397;
assign w8409 = ~w8407 & ~w8408;
assign w8410 = pi0833 & ~w397;
assign w8411 = pi0857 & w397;
assign w8412 = ~w8410 & ~w8411;
assign w8413 = pi0834 & ~w397;
assign w8414 = pi0858 & w397;
assign w8415 = ~w8413 & ~w8414;
assign w8416 = pi0812 & ~w397;
assign w8417 = pi0758 & w397;
assign w8418 = ~w8416 & ~w8417;
assign w8419 = pi0813 & ~w397;
assign w8420 = pi0836 & w397;
assign w8421 = ~w8419 & ~w8420;
assign w8422 = pi1014 & w8363;
assign w8423 = pi1480 & w7571;
assign w8424 = ~w8422 & ~w8423;
assign w8425 = pi0728 & ~pi1329;
assign w8426 = pi0644 & ~pi1324;
assign w8427 = pi0987 & ~pi1325;
assign w8428 = pi0136 & ~pi1326;
assign w8429 = pi0986 & ~pi1339;
assign w8430 = pi0786 & ~pi1288;
assign w8431 = pi0915 & ~pi1327;
assign w8432 = pi0977 & ~pi1330;
assign w8433 = pi0901 & ~pi1328;
assign w8434 = ~pi1611 & pi1612;
assign w8435 = pi1613 & pi1620;
assign w8436 = w8434 & w8435;
assign w8437 = ~w8425 & ~w8426;
assign w8438 = ~w8427 & ~w8428;
assign w8439 = ~w8429 & ~w8430;
assign w8440 = ~w8431 & ~w8432;
assign w8441 = ~w8433 & w8440;
assign w8442 = w8438 & w8439;
assign w8443 = w8436 & w8437;
assign w8444 = w8442 & w8443;
assign w8445 = w8441 & w8444;
assign w8446 = ~pi1229 & w5455;
assign w8447 = w8315 & ~w8446;
assign w8448 = w376 & ~w7778;
assign w8449 = ~pi0802 & w374;
assign w8450 = w7777 & w8449;
assign w8451 = ~w8448 & ~w8450;
assign w8452 = w1705 & w7766;
assign w8453 = ~w8451 & w8452;
assign w8454 = ~w8447 & ~w8453;
assign w8455 = pi1017 & ~w3565;
assign w8456 = ~pi1738 & w3565;
assign w8457 = ~w8455 & ~w8456;
assign w8458 = w1298 & ~w1416;
assign w8459 = pi1018 & ~w8458;
assign w8460 = ~w1290 & ~w8459;
assign w8461 = pi1747 & ~w8460;
assign w8462 = w8273 & w8276;
assign w8463 = ~pi0262 & w6718;
assign w8464 = w2163 & w8463;
assign w8465 = ~w8462 & ~w8464;
assign w8466 = pi0986 & ~pi1323;
assign w8467 = pi0915 & pi1290;
assign w8468 = pi0136 & pi1289;
assign w8469 = pi0987 & pi1319;
assign w8470 = pi0786 & pi1320;
assign w8471 = pi0977 & ~pi1287;
assign w8472 = pi0728 & pi1322;
assign w8473 = pi0901 & pi1321;
assign w8474 = pi0644 & pi1291;
assign w8475 = pi1616 & ~pi1617;
assign w8476 = pi1618 & pi1619;
assign w8477 = w8475 & w8476;
assign w8478 = ~w8466 & ~w8467;
assign w8479 = ~w8468 & ~w8469;
assign w8480 = ~w8470 & ~w8471;
assign w8481 = ~w8472 & ~w8473;
assign w8482 = ~w8474 & w8481;
assign w8483 = w8479 & w8480;
assign w8484 = w8477 & w8478;
assign w8485 = w8483 & w8484;
assign w8486 = w8482 & w8485;
assign w8487 = w2133 & w6718;
assign w8488 = w6811 & w8487;
assign w8489 = w2868 & w6620;
assign w8490 = pi1747 & ~w8489;
assign w8491 = pi1022 & w8490;
assign w8492 = pi1747 & w8489;
assign w8493 = pi1776 & w8492;
assign w8494 = ~w8491 & ~w8493;
assign w8495 = pi1023 & w8490;
assign w8496 = pi1778 & w8492;
assign w8497 = ~w8495 & ~w8496;
assign w8498 = pi1024 & w8490;
assign w8499 = pi1790 & w8492;
assign w8500 = ~w8498 & ~w8499;
assign w8501 = pi1025 & w8490;
assign w8502 = pi1791 & w8492;
assign w8503 = ~w8501 & ~w8502;
assign w8504 = pi1026 & w8490;
assign w8505 = pi1792 & w8492;
assign w8506 = ~w8504 & ~w8505;
assign w8507 = w2868 & w6627;
assign w8508 = pi1747 & ~w8507;
assign w8509 = pi1027 & w8508;
assign w8510 = pi1747 & w8507;
assign w8511 = pi1776 & w8510;
assign w8512 = ~w8509 & ~w8511;
assign w8513 = pi1028 & w8508;
assign w8514 = pi1779 & w8510;
assign w8515 = ~w8513 & ~w8514;
assign w8516 = pi1029 & w8508;
assign w8517 = pi1783 & w8510;
assign w8518 = ~w8516 & ~w8517;
assign w8519 = ~pi1030 & w8508;
assign w8520 = pi1799 & w8510;
assign w8521 = ~w8519 & ~w8520;
assign w8522 = w2868 & w6622;
assign w8523 = pi1747 & w8522;
assign w8524 = pi1774 & w8523;
assign w8525 = pi1747 & ~w8522;
assign w8526 = ~pi1031 & w8525;
assign w8527 = ~w8524 & ~w8526;
assign w8528 = pi1776 & w8523;
assign w8529 = pi1032 & w8525;
assign w8530 = ~w8528 & ~w8529;
assign w8531 = pi1780 & w8523;
assign w8532 = pi1033 & w8525;
assign w8533 = ~w8531 & ~w8532;
assign w8534 = pi1783 & w8523;
assign w8535 = pi1034 & w8525;
assign w8536 = ~w8534 & ~w8535;
assign w8537 = pi1459 & w1248;
assign w8538 = ~pi1035 & ~w8537;
assign w8539 = w1769 & ~w8538;
assign w8540 = pi1036 & ~w3151;
assign w8541 = w3931 & ~w8540;
assign w8542 = pi1447 & w1248;
assign w8543 = ~pi1037 & ~w8542;
assign w8544 = w1783 & ~w8543;
assign w8545 = ~pi1038 & w6402;
assign w8546 = pi0971 & w2134;
assign w8547 = ~w2176 & ~w8546;
assign w8548 = ~w2163 & w8547;
assign w8549 = ~w2174 & w8548;
assign w8550 = ~w8545 & w8549;
assign w8551 = pi1039 & ~w3565;
assign w8552 = ~pi1733 & w3565;
assign w8553 = ~w8551 & ~w8552;
assign w8554 = pi1040 & ~w3565;
assign w8555 = ~pi1741 & w3565;
assign w8556 = ~w8554 & ~w8555;
assign w8557 = pi1041 & ~w3565;
assign w8558 = ~pi1727 & w3565;
assign w8559 = ~w8557 & ~w8558;
assign w8560 = pi1042 & ~w3565;
assign w8561 = ~pi1740 & w3565;
assign w8562 = ~w8560 & ~w8561;
assign w8563 = pi1043 & ~w3565;
assign w8564 = ~pi1735 & w3565;
assign w8565 = ~w8563 & ~w8564;
assign w8566 = pi1044 & ~w3565;
assign w8567 = ~pi1725 & w3565;
assign w8568 = ~w8566 & ~w8567;
assign w8569 = ~pi0277 & w8252;
assign w8570 = ~w2164 & ~w8569;
assign w8571 = w8249 & ~w8570;
assign w8572 = ~w2133 & ~w6397;
assign w8573 = pi0276 & ~w8572;
assign w8574 = w2151 & ~w8573;
assign w8575 = ~w2180 & ~w8574;
assign w8576 = w2150 & w6718;
assign w8577 = ~w8575 & w8576;
assign w8578 = ~w397 & w1007;
assign w8579 = pi1459 & pi1729;
assign w8580 = ~pi1048 & ~w8579;
assign w8581 = w1769 & ~w8580;
assign w8582 = pi1049 & ~w3565;
assign w8583 = ~pi1722 & w3565;
assign w8584 = ~w8582 & ~w8583;
assign w8585 = pi0183 & w6405;
assign w8586 = ~w2174 & ~w8585;
assign w8587 = w6718 & ~w8586;
assign w8588 = w2868 & w6612;
assign w8589 = pi1747 & ~w8588;
assign w8590 = pi1051 & w8589;
assign w8591 = pi1747 & w8588;
assign w8592 = pi1791 & w8591;
assign w8593 = ~w8590 & ~w8592;
assign w8594 = ~pi1052 & w8589;
assign w8595 = pi1787 & w8591;
assign w8596 = ~w8594 & ~w8595;
assign w8597 = ~pi1053 & ~w2869;
assign w8598 = w2982 & ~w8597;
assign w8599 = pi1054 & w8508;
assign w8600 = pi1792 & w8510;
assign w8601 = ~w8599 & ~w8600;
assign w8602 = ~pi1055 & ~w2869;
assign w8603 = w3144 & ~w8602;
assign w8604 = pi1056 & ~w3954;
assign w8605 = w5664 & ~w8604;
assign w8606 = pi1057 & ~w3954;
assign w8607 = w3961 & ~w8606;
assign w8608 = pi1738 & w6045;
assign w8609 = pi1747 & ~w6044;
assign w8610 = ~pi1058 & w8609;
assign w8611 = ~w8608 & ~w8610;
assign w8612 = ~pi1361 & w6612;
assign w8613 = ~pi0686 & w5442;
assign w8614 = ~pi0495 & w3188;
assign w8615 = pi0136 & w6637;
assign w8616 = ~pi0604 & w4056;
assign w8617 = pi0273 & w6633;
assign w8618 = ~pi1329 & w6615;
assign w8619 = ~pi0396 & w2932;
assign w8620 = ~pi0438 & w2866;
assign w8621 = ~pi1360 & w6620;
assign w8622 = ~pi0536 & w3150;
assign w8623 = ~pi1413 & w6622;
assign w8624 = ~pi0576 & w4186;
assign w8625 = ~pi0525 & w3953;
assign w8626 = ~pi1369 & w6627;
assign w8627 = ~w8612 & ~w8613;
assign w8628 = ~w8614 & ~w8616;
assign w8629 = ~w8619 & ~w8620;
assign w8630 = ~w8621 & ~w8622;
assign w8631 = ~w8623 & ~w8624;
assign w8632 = ~w8625 & ~w8626;
assign w8633 = w8631 & w8632;
assign w8634 = w8629 & w8630;
assign w8635 = w8627 & w8628;
assign w8636 = ~w8615 & ~w8617;
assign w8637 = ~w8618 & w8636;
assign w8638 = w8634 & w8635;
assign w8639 = w8633 & w8638;
assign w8640 = w8637 & w8639;
assign w8641 = ~pi0446 & w3188;
assign w8642 = ~pi0687 & w5442;
assign w8643 = ~pi0399 & w2932;
assign w8644 = pi0252 & w6633;
assign w8645 = ~pi0420 & w3150;
assign w8646 = ~pi1339 & w6615;
assign w8647 = pi0786 & w6637;
assign w8648 = ~pi1164 & w6612;
assign w8649 = ~pi0602 & w4056;
assign w8650 = ~pi0577 & w4186;
assign w8651 = ~pi0343 & w2866;
assign w8652 = ~pi1184 & w6620;
assign w8653 = ~pi1225 & w6622;
assign w8654 = ~pi1206 & w6627;
assign w8655 = ~pi0657 & w3953;
assign w8656 = ~w8641 & ~w8642;
assign w8657 = ~w8643 & ~w8645;
assign w8658 = ~w8648 & ~w8649;
assign w8659 = ~w8650 & ~w8651;
assign w8660 = ~w8652 & ~w8653;
assign w8661 = ~w8654 & ~w8655;
assign w8662 = w8660 & w8661;
assign w8663 = w8658 & w8659;
assign w8664 = w8656 & w8657;
assign w8665 = ~w8644 & ~w8646;
assign w8666 = ~w8647 & w8665;
assign w8667 = w8663 & w8664;
assign w8668 = w8662 & w8667;
assign w8669 = w8666 & w8668;
assign w8670 = pi1081 & w6612;
assign w8671 = ~pi0324 & w2866;
assign w8672 = pi1142 & w6622;
assign w8673 = pi0467 & w6633;
assign w8674 = ~pi0558 & w4056;
assign w8675 = pi1685 & w6641;
assign w8676 = ~pi1323 & w6615;
assign w8677 = ~pi0330 & w2932;
assign w8678 = ~pi0375 & w3188;
assign w8679 = ~pi0371 & w3150;
assign w8680 = ~pi0464 & w4186;
assign w8681 = pi1274 & w6620;
assign w8682 = ~pi0624 & w5442;
assign w8683 = ~pi0459 & w3953;
assign w8684 = pi1130 & w6627;
assign w8685 = ~w8670 & ~w8671;
assign w8686 = ~w8672 & ~w8674;
assign w8687 = ~w8677 & ~w8678;
assign w8688 = ~w8679 & ~w8680;
assign w8689 = ~w8681 & ~w8682;
assign w8690 = ~w8683 & ~w8684;
assign w8691 = w8689 & w8690;
assign w8692 = w8687 & w8688;
assign w8693 = w8685 & w8686;
assign w8694 = ~w8673 & ~w8675;
assign w8695 = ~w8676 & w8694;
assign w8696 = w8692 & w8693;
assign w8697 = w8691 & w8696;
assign w8698 = w8695 & w8697;
assign w8699 = ~pi1062 & ~w3954;
assign w8700 = w4173 & ~w8699;
assign w8701 = ~pi1063 & ~w3151;
assign w8702 = w3348 & ~w8701;
assign w8703 = ~pi1064 & ~w3954;
assign w8704 = w4733 & ~w8703;
assign w8705 = ~pi1065 & ~w3151;
assign w8706 = w5367 & ~w8705;
assign w8707 = pi1066 & ~w3954;
assign w8708 = w5656 & ~w8707;
assign w8709 = ~pi1067 & ~w2869;
assign w8710 = w4219 & ~w8709;
assign w8711 = w2868 & w6639;
assign w8712 = pi1747 & ~w8711;
assign w8713 = pi1068 & w8712;
assign w8714 = pi1747 & w8711;
assign w8715 = pi1779 & w8714;
assign w8716 = ~w8713 & ~w8715;
assign w8717 = pi1069 & w8712;
assign w8718 = pi1777 & w8714;
assign w8719 = ~w8717 & ~w8718;
assign w8720 = pi1070 & w8589;
assign w8721 = pi1795 & w8591;
assign w8722 = ~w8720 & ~w8721;
assign w8723 = ~pi1071 & ~w3954;
assign w8724 = w4669 & ~w8723;
assign w8725 = ~pi0404 & w2932;
assign w8726 = pi1076 & w6627;
assign w8727 = ~pi0694 & w5442;
assign w8728 = ~pi0584 & w4186;
assign w8729 = pi1270 & w6620;
assign w8730 = ~pi0610 & w4056;
assign w8731 = pi0479 & w6633;
assign w8732 = ~pi1287 & w6615;
assign w8733 = pi1265 & w6622;
assign w8734 = pi1109 & w6612;
assign w8735 = ~pi0356 & w3150;
assign w8736 = ~pi0349 & w2866;
assign w8737 = ~pi0436 & w3953;
assign w8738 = ~pi0503 & w3188;
assign w8739 = ~w8725 & ~w8726;
assign w8740 = ~w8727 & ~w8728;
assign w8741 = ~w8729 & ~w8730;
assign w8742 = ~w8733 & ~w8734;
assign w8743 = ~w8735 & ~w8736;
assign w8744 = ~w8737 & ~w8738;
assign w8745 = w8743 & w8744;
assign w8746 = w8741 & w8742;
assign w8747 = w8739 & w8740;
assign w8748 = ~w8731 & ~w8732;
assign w8749 = w8747 & w8748;
assign w8750 = w8745 & w8746;
assign w8751 = w8749 & w8750;
assign w8752 = ~pi1073 & ~w2869;
assign w8753 = w2962 & ~w8752;
assign w8754 = pi1074 & w8589;
assign w8755 = pi1799 & w8591;
assign w8756 = ~w8754 & ~w8755;
assign w8757 = ~pi1075 & ~w2869;
assign w8758 = w2886 & ~w8757;
assign w8759 = pi1076 & w8508;
assign w8760 = pi1782 & w8510;
assign w8761 = ~w8759 & ~w8760;
assign w8762 = pi1077 & ~w2869;
assign w8763 = w3080 & ~w8762;
assign w8764 = ~pi1078 & w8508;
assign w8765 = pi1790 & w8510;
assign w8766 = ~w8764 & ~w8765;
assign w8767 = pi1725 & w6045;
assign w8768 = ~pi1079 & w8609;
assign w8769 = ~w8767 & ~w8768;
assign w8770 = pi1080 & w8508;
assign w8771 = pi1800 & w8510;
assign w8772 = ~w8770 & ~w8771;
assign w8773 = pi1081 & w8589;
assign w8774 = pi1781 & w8591;
assign w8775 = ~w8773 & ~w8774;
assign w8776 = pi1082 & ~w2869;
assign w8777 = w2878 & ~w8776;
assign w8778 = pi1083 & w8508;
assign w8779 = pi1780 & w8510;
assign w8780 = ~w8778 & ~w8779;
assign w8781 = ~pi1084 & w8508;
assign w8782 = pi1786 & w8510;
assign w8783 = ~w8781 & ~w8782;
assign w8784 = ~pi1085 & ~w3954;
assign w8785 = w4165 & ~w8784;
assign w8786 = ~pi1086 & ~w3954;
assign w8787 = w4080 & ~w8786;
assign w8788 = pi1087 & ~w2869;
assign w8789 = w4072 & ~w8788;
assign w8790 = pi1088 & ~pi1101;
assign w8791 = ~w1290 & ~w8790;
assign w8792 = w13 & ~w8791;
assign w8793 = ~pi1547 & w2846;
assign w8794 = w224 & w226;
assign w8795 = w8793 & w8794;
assign w8796 = ~w8792 & ~w8795;
assign w8797 = w1755 & ~w8796;
assign w8798 = pi1089 & ~w2869;
assign w8799 = w3120 & ~w8798;
assign w8800 = w2841 & w2843;
assign w8801 = ~w8 & ~w8800;
assign w8802 = pi1747 & ~w8801;
assign w8803 = pi1091 & w15;
assign w8804 = w2838 & w2840;
assign w8805 = ~w8803 & ~w8804;
assign w8806 = w1755 & ~w8805;
assign w8807 = pi1092 & w8508;
assign w8808 = pi1775 & w8510;
assign w8809 = ~w8807 & ~w8808;
assign w8810 = pi1093 & ~w2869;
assign w8811 = w3104 & ~w8810;
assign w8812 = pi1094 & w8712;
assign w8813 = pi1774 & w8714;
assign w8814 = ~w8812 & ~w8813;
assign w8815 = pi1095 & w8712;
assign w8816 = pi1775 & w8714;
assign w8817 = ~w8815 & ~w8816;
assign w8818 = pi1096 & w8712;
assign w8819 = pi1776 & w8714;
assign w8820 = ~w8818 & ~w8819;
assign w8821 = pi1097 & w8712;
assign w8822 = pi1778 & w8714;
assign w8823 = ~w8821 & ~w8822;
assign w8824 = pi1098 & w8712;
assign w8825 = pi1780 & w8714;
assign w8826 = ~w8824 & ~w8825;
assign w8827 = w6418 & ~w6448;
assign w8828 = w6535 & w8827;
assign w8829 = w6445 & w8828;
assign w8830 = pi0112 & w404;
assign w8831 = ~w8829 & w8830;
assign w8832 = pi1787 & w8523;
assign w8833 = ~pi1100 & w8525;
assign w8834 = ~w8832 & ~w8833;
assign w8835 = pi1102 & w8589;
assign w8836 = pi1784 & w8591;
assign w8837 = ~w8835 & ~w8836;
assign w8838 = ~pi1103 & w8589;
assign w8839 = pi1786 & w8591;
assign w8840 = ~w8838 & ~w8839;
assign w8841 = pi1104 & w8589;
assign w8842 = pi1775 & w8591;
assign w8843 = ~w8841 & ~w8842;
assign w8844 = pi1105 & w8589;
assign w8845 = pi1776 & w8591;
assign w8846 = ~w8844 & ~w8845;
assign w8847 = pi1106 & w8589;
assign w8848 = pi1778 & w8591;
assign w8849 = ~w8847 & ~w8848;
assign w8850 = pi1107 & w8589;
assign w8851 = pi1779 & w8591;
assign w8852 = ~w8850 & ~w8851;
assign w8853 = pi1108 & w8589;
assign w8854 = pi1780 & w8591;
assign w8855 = ~w8853 & ~w8854;
assign w8856 = pi1109 & w8589;
assign w8857 = pi1782 & w8591;
assign w8858 = ~w8856 & ~w8857;
assign w8859 = pi1110 & w8589;
assign w8860 = pi1783 & w8591;
assign w8861 = ~w8859 & ~w8860;
assign w8862 = pi1111 & w8589;
assign w8863 = pi1789 & w8591;
assign w8864 = ~w8862 & ~w8863;
assign w8865 = pi1112 & w8589;
assign w8866 = pi1800 & w8591;
assign w8867 = ~w8865 & ~w8866;
assign w8868 = pi1113 & w8589;
assign w8869 = pi1801 & w8591;
assign w8870 = ~w8868 & ~w8869;
assign w8871 = pi1114 & w8589;
assign w8872 = pi1790 & w8591;
assign w8873 = ~w8871 & ~w8872;
assign w8874 = pi1115 & w8589;
assign w8875 = pi1792 & w8591;
assign w8876 = ~w8874 & ~w8875;
assign w8877 = pi1116 & w8589;
assign w8878 = pi1793 & w8591;
assign w8879 = ~w8877 & ~w8878;
assign w8880 = pi1117 & w8589;
assign w8881 = pi1794 & w8591;
assign w8882 = ~w8880 & ~w8881;
assign w8883 = pi1118 & w8589;
assign w8884 = pi1798 & w8591;
assign w8885 = ~w8883 & ~w8884;
assign w8886 = pi1119 & w8490;
assign w8887 = pi1784 & w8492;
assign w8888 = ~w8886 & ~w8887;
assign w8889 = ~pi1120 & w8490;
assign w8890 = pi1786 & w8492;
assign w8891 = ~w8889 & ~w8890;
assign w8892 = pi1121 & w8490;
assign w8893 = pi1780 & w8492;
assign w8894 = ~w8892 & ~w8893;
assign w8895 = pi1122 & w8490;
assign w8896 = pi1789 & w8492;
assign w8897 = ~w8895 & ~w8896;
assign w8898 = pi1123 & w8490;
assign w8899 = pi1794 & w8492;
assign w8900 = ~w8898 & ~w8899;
assign w8901 = pi1124 & w8490;
assign w8902 = pi1798 & w8492;
assign w8903 = ~w8901 & ~w8902;
assign w8904 = ~pi1125 & w8490;
assign w8905 = pi1787 & w8492;
assign w8906 = ~w8904 & ~w8905;
assign w8907 = ~pi1126 & w8508;
assign w8908 = pi1774 & w8510;
assign w8909 = ~w8907 & ~w8908;
assign w8910 = pi1127 & w8508;
assign w8911 = pi1784 & w8510;
assign w8912 = ~w8910 & ~w8911;
assign w8913 = ~pi1128 & w8508;
assign w8914 = pi1785 & w8510;
assign w8915 = ~w8913 & ~w8914;
assign w8916 = pi1129 & w8508;
assign w8917 = pi1778 & w8510;
assign w8918 = ~w8916 & ~w8917;
assign w8919 = pi1130 & w8508;
assign w8920 = pi1781 & w8510;
assign w8921 = ~w8919 & ~w8920;
assign w8922 = pi1131 & w8508;
assign w8923 = pi1789 & w8510;
assign w8924 = ~w8922 & ~w8923;
assign w8925 = pi1132 & w8508;
assign w8926 = pi1801 & w8510;
assign w8927 = ~w8925 & ~w8926;
assign w8928 = ~pi1133 & w8508;
assign w8929 = pi1791 & w8510;
assign w8930 = ~w8928 & ~w8929;
assign w8931 = pi1134 & w8508;
assign w8932 = pi1793 & w8510;
assign w8933 = ~w8931 & ~w8932;
assign w8934 = pi1135 & w8508;
assign w8935 = pi1794 & w8510;
assign w8936 = ~w8934 & ~w8935;
assign w8937 = pi1136 & w8508;
assign w8938 = pi1795 & w8510;
assign w8939 = ~w8937 & ~w8938;
assign w8940 = ~pi1137 & w8508;
assign w8941 = pi1798 & w8510;
assign w8942 = ~w8940 & ~w8941;
assign w8943 = ~pi1138 & w8508;
assign w8944 = pi1787 & w8510;
assign w8945 = ~w8943 & ~w8944;
assign w8946 = pi1784 & w8523;
assign w8947 = pi1139 & w8525;
assign w8948 = ~w8946 & ~w8947;
assign w8949 = pi1786 & w8523;
assign w8950 = ~pi1140 & w8525;
assign w8951 = ~w8949 & ~w8950;
assign w8952 = pi1778 & w8523;
assign w8953 = pi1141 & w8525;
assign w8954 = ~w8952 & ~w8953;
assign w8955 = pi1781 & w8523;
assign w8956 = pi1142 & w8525;
assign w8957 = ~w8955 & ~w8956;
assign w8958 = pi1789 & w8523;
assign w8959 = pi1143 & w8525;
assign w8960 = ~w8958 & ~w8959;
assign w8961 = pi1800 & w8523;
assign w8962 = pi1144 & w8525;
assign w8963 = ~w8961 & ~w8962;
assign w8964 = pi1790 & w8523;
assign w8965 = pi1145 & w8525;
assign w8966 = ~w8964 & ~w8965;
assign w8967 = pi1792 & w8523;
assign w8968 = pi1146 & w8525;
assign w8969 = ~w8967 & ~w8968;
assign w8970 = pi1795 & w8523;
assign w8971 = pi1147 & w8525;
assign w8972 = ~w8970 & ~w8971;
assign w8973 = pi1794 & w8523;
assign w8974 = pi1148 & w8525;
assign w8975 = ~w8973 & ~w8974;
assign w8976 = ~pi1149 & ~w4057;
assign w8977 = w5219 & ~w8976;
assign w8978 = ~pi1150 & ~w4057;
assign w8979 = w5279 & ~w8978;
assign w8980 = ~pi1151 & ~w4057;
assign w8981 = w4947 & ~w8980;
assign w8982 = ~pi1152 & ~w4057;
assign w8983 = w4971 & ~w8982;
assign w8984 = ~pi1153 & ~w4057;
assign w8985 = w5231 & ~w8984;
assign w8986 = pi1154 & ~w4057;
assign w8987 = w4849 & ~w8986;
assign w8988 = pi1155 & ~w4057;
assign w8989 = w5303 & ~w8988;
assign w8990 = pi1156 & ~w4057;
assign w8991 = w5287 & ~w8990;
assign w8992 = pi1157 & ~w4057;
assign w8993 = w5295 & ~w8992;
assign w8994 = pi1158 & ~w4057;
assign w8995 = w5319 & ~w8994;
assign w8996 = pi1159 & ~w4057;
assign w8997 = w4621 & ~w8996;
assign w8998 = pi1160 & ~w4057;
assign w8999 = w5335 & ~w8998;
assign w9000 = ~pi1161 & ~w4057;
assign w9001 = w4064 & ~w9000;
assign w9002 = ~pi1162 & ~w4057;
assign w9003 = w4857 & ~w9002;
assign w9004 = ~pi1163 & ~w4057;
assign w9005 = w5351 & ~w9004;
assign w9006 = pi1797 & w8591;
assign w9007 = ~pi1052 & pi1729;
assign w9008 = ~pi1164 & ~w9007;
assign w9009 = w8589 & w9008;
assign w9010 = ~w9006 & ~w9009;
assign w9011 = pi1480 & w1248;
assign w9012 = ~pi1165 & ~w9011;
assign w9013 = w1773 & ~w9012;
assign w9014 = ~pi1166 & ~w2869;
assign w9015 = w2918 & ~w9014;
assign w9016 = ~pi1167 & ~w2869;
assign w9017 = w2946 & ~w9016;
assign w9018 = ~pi1168 & ~w2869;
assign w9019 = w4629 & ~w9018;
assign w9020 = ~pi1169 & ~w2869;
assign w9021 = w2910 & ~w9020;
assign w9022 = ~pi1170 & ~w2869;
assign w9023 = w4637 & ~w9022;
assign w9024 = ~pi1171 & ~w2869;
assign w9025 = w3056 & ~w9024;
assign w9026 = ~pi1172 & ~w2869;
assign w9027 = w3072 & ~w9026;
assign w9028 = pi1173 & ~w2869;
assign w9029 = w3088 & ~w9028;
assign w9030 = pi1174 & ~w2869;
assign w9031 = w3096 & ~w9030;
assign w9032 = pi1175 & ~w2869;
assign w9033 = w3112 & ~w9032;
assign w9034 = pi1176 & ~w2869;
assign w9035 = w2902 & ~w9034;
assign w9036 = pi1177 & ~w2869;
assign w9037 = w4653 & ~w9036;
assign w9038 = ~pi1178 & ~w2869;
assign w9039 = w4043 & ~w9038;
assign w9040 = pi1179 & ~w2869;
assign w9041 = w3128 & ~w9040;
assign w9042 = ~pi1180 & ~w2869;
assign w9043 = w3136 & ~w9042;
assign w9044 = ~pi1181 & ~w2869;
assign w9045 = w4136 & ~w9044;
assign w9046 = ~pi1182 & ~w2869;
assign w9047 = w2894 & ~w9046;
assign w9048 = ~pi1183 & ~w4057;
assign w9049 = w5359 & ~w9048;
assign w9050 = pi1797 & w8492;
assign w9051 = ~pi1125 & pi1729;
assign w9052 = ~pi1184 & ~w9051;
assign w9053 = w8490 & w9052;
assign w9054 = ~w9050 & ~w9053;
assign w9055 = ~pi1185 & ~w3151;
assign w9056 = w3340 & ~w9055;
assign w9057 = ~pi1186 & ~w3151;
assign w9058 = w3362 & ~w9057;
assign w9059 = ~pi1187 & ~w3151;
assign w9060 = w5375 & ~w9059;
assign w9061 = ~pi1188 & ~w3151;
assign w9062 = w3332 & ~w9061;
assign w9063 = ~pi1189 & ~w3151;
assign w9064 = w3370 & ~w9063;
assign w9065 = ~pi1190 & ~w3151;
assign w9066 = w3851 & ~w9065;
assign w9067 = ~pi1191 & ~w3151;
assign w9068 = w3859 & ~w9067;
assign w9069 = pi1192 & ~w3151;
assign w9070 = w3867 & ~w9069;
assign w9071 = ~pi1193 & ~w3151;
assign w9072 = w3875 & ~w9071;
assign w9073 = pi1194 & ~w3151;
assign w9074 = w3891 & ~w9073;
assign w9075 = pi1195 & ~w3151;
assign w9076 = w4784 & ~w9075;
assign w9077 = pi1196 & ~w3151;
assign w9078 = w3899 & ~w9077;
assign w9079 = pi1197 & ~w3151;
assign w9080 = w3915 & ~w9079;
assign w9081 = pi1198 & ~w3151;
assign w9082 = w4030 & ~w9081;
assign w9083 = pi1199 & ~w3151;
assign w9084 = w3923 & ~w9083;
assign w9085 = ~pi1200 & ~w3151;
assign w9086 = w4773 & ~w9085;
assign w9087 = pi1201 & ~w3151;
assign w9088 = w5394 & ~w9087;
assign w9089 = ~pi1202 & ~w3151;
assign w9090 = w3939 & ~w9089;
assign w9091 = ~pi1203 & ~w3151;
assign w9092 = w4995 & ~w9091;
assign w9093 = ~pi1204 & ~w3151;
assign w9094 = w4865 & ~w9093;
assign w9095 = ~pi1205 & ~w3151;
assign w9096 = w3390 & ~w9095;
assign w9097 = pi1797 & w8510;
assign w9098 = ~pi1138 & pi1729;
assign w9099 = ~pi1206 & ~w9098;
assign w9100 = w8508 & w9099;
assign w9101 = ~w9097 & ~w9100;
assign w9102 = ~pi1207 & ~w3954;
assign w9103 = w4661 & ~w9102;
assign w9104 = ~pi1208 & ~w3954;
assign w9105 = w4157 & ~w9104;
assign w9106 = ~pi1209 & ~w3954;
assign w9107 = w4181 & ~w9106;
assign w9108 = ~pi1210 & ~w3954;
assign w9109 = w4199 & ~w9108;
assign w9110 = ~pi1211 & ~w3954;
assign w9111 = w4677 & ~w9110;
assign w9112 = ~pi1212 & ~w3954;
assign w9113 = w4685 & ~w9112;
assign w9114 = pi1213 & ~w3954;
assign w9115 = w4116 & ~w9114;
assign w9116 = pi1214 & ~w3954;
assign w9117 = w4693 & ~w9116;
assign w9118 = pi1215 & ~w3954;
assign w9119 = w5648 & ~w9118;
assign w9120 = pi1216 & ~w3954;
assign w9121 = w4701 & ~w9120;
assign w9122 = pi1217 & ~w3954;
assign w9123 = w4709 & ~w9122;
assign w9124 = pi1218 & ~w3954;
assign w9125 = w4717 & ~w9124;
assign w9126 = pi1219 & ~w3954;
assign w9127 = w5484 & ~w9126;
assign w9128 = ~pi1220 & ~w3954;
assign w9129 = w5464 & ~w9128;
assign w9130 = ~pi1221 & ~w3954;
assign w9131 = w3969 & ~w9130;
assign w9132 = ~pi1222 & ~w3954;
assign w9133 = w5502 & ~w9132;
assign w9134 = ~pi1223 & ~w3954;
assign w9135 = w4227 & ~w9134;
assign w9136 = ~pi1224 & ~w3954;
assign w9137 = w5672 & ~w9136;
assign w9138 = pi1797 & w8523;
assign w9139 = ~pi1100 & pi1729;
assign w9140 = ~pi1225 & ~w9139;
assign w9141 = w8525 & w9140;
assign w9142 = ~w9138 & ~w9141;
assign w9143 = ~pi1445 & ~pi1773;
assign w9144 = pi1773 & ~pi1820;
assign w9145 = ~w9143 & ~w9144;
assign w9146 = ~pi1733 & w6045;
assign w9147 = pi1227 & w8609;
assign w9148 = ~w9146 & ~w9147;
assign w9149 = ~pi1741 & w6045;
assign w9150 = pi1228 & w8609;
assign w9151 = ~w9149 & ~w9150;
assign w9152 = ~pi1722 & w6045;
assign w9153 = pi1229 & w8609;
assign w9154 = ~w9152 & ~w9153;
assign w9155 = pi1740 & w6045;
assign w9156 = ~pi1230 & w8609;
assign w9157 = ~w9155 & ~w9156;
assign w9158 = pi1735 & w6045;
assign w9159 = ~pi1231 & w8609;
assign w9160 = ~w9158 & ~w9159;
assign w9161 = pi1232 & ~w3954;
assign w9162 = w4725 & ~w9161;
assign w9163 = ~pi1627 & w1710;
assign w9164 = w3564 & w9163;
assign w9165 = ~pi1427 & ~w9164;
assign w9166 = ~pi1235 & w8490;
assign w9167 = pi1774 & w8492;
assign w9168 = ~w9166 & ~w9167;
assign w9169 = ~pi1727 & w6045;
assign w9170 = pi1236 & w8609;
assign w9171 = ~w9169 & ~w9170;
assign w9172 = ~pi1237 & w8589;
assign w9173 = pi1774 & w8591;
assign w9174 = ~w9172 & ~w9173;
assign w9175 = ~pi1238 & ~w3151;
assign w9176 = w3166 & ~w9175;
assign w9177 = ~pi1239 & ~w2869;
assign w9178 = w2926 & ~w9177;
assign w9179 = ~pi1240 & ~w3151;
assign w9180 = w3947 & ~w9179;
assign w9181 = pi1241 & ~w2869;
assign w9182 = w3064 & ~w9181;
assign w9183 = pi1798 & w8523;
assign w9184 = pi1242 & w8525;
assign w9185 = ~w9183 & ~w9184;
assign w9186 = ~pi1243 & w8589;
assign w9187 = pi1785 & w8591;
assign w9188 = ~w9186 & ~w9187;
assign w9189 = ~pi1244 & ~w3151;
assign w9190 = w3324 & ~w9189;
assign w9191 = ~pi1245 & ~w3151;
assign w9192 = w3183 & ~w9191;
assign w9193 = ~pi1246 & ~w2869;
assign w9194 = w2954 & ~w9193;
assign w9195 = ~pi1247 & ~w2869;
assign w9196 = w4645 & ~w9195;
assign w9197 = ~pi1248 & ~w3151;
assign w9198 = w5383 & ~w9197;
assign w9199 = pi1249 & ~w3151;
assign w9200 = w3158 & ~w9199;
assign w9201 = ~pi0073 & w1298;
assign w9202 = ~pi1418 & ~w9201;
assign w9203 = pi1252 & w8490;
assign w9204 = pi1799 & w8492;
assign w9205 = ~w9203 & ~w9204;
assign w9206 = pi1793 & w8523;
assign w9207 = pi1253 & w8525;
assign w9208 = ~w9206 & ~w9207;
assign w9209 = ~pi1254 & ~w2869;
assign w9210 = w3048 & ~w9209;
assign w9211 = pi1791 & w8523;
assign w9212 = pi1255 & w8525;
assign w9213 = ~w9211 & ~w9212;
assign w9214 = pi1256 & w8490;
assign w9215 = pi1800 & w8492;
assign w9216 = ~w9214 & ~w9215;
assign w9217 = pi1257 & w8490;
assign w9218 = pi1801 & w8492;
assign w9219 = ~w9217 & ~w9218;
assign w9220 = pi1779 & w8523;
assign w9221 = pi1258 & w8525;
assign w9222 = ~w9220 & ~w9221;
assign w9223 = pi1801 & w8523;
assign w9224 = pi1259 & w8525;
assign w9225 = ~w9223 & ~w9224;
assign w9226 = pi1260 & w8490;
assign w9227 = pi1793 & w8492;
assign w9228 = ~w9226 & ~w9227;
assign w9229 = pi1799 & w8523;
assign w9230 = pi1261 & w8525;
assign w9231 = ~w9229 & ~w9230;
assign w9232 = pi1262 & w8490;
assign w9233 = pi1795 & w8492;
assign w9234 = ~w9232 & ~w9233;
assign w9235 = ~pi1263 & ~w4057;
assign w9236 = w5343 & ~w9235;
assign w9237 = pi1264 & ~w3151;
assign w9238 = w3907 & ~w9237;
assign w9239 = pi1782 & w8523;
assign w9240 = pi1265 & w8525;
assign w9241 = ~w9239 & ~w9240;
assign w9242 = pi1266 & ~w3954;
assign w9243 = w4741 & ~w9242;
assign w9244 = pi1267 & w8490;
assign w9245 = pi1783 & w8492;
assign w9246 = ~w9244 & ~w9245;
assign w9247 = ~pi1268 & w8490;
assign w9248 = pi1785 & w8492;
assign w9249 = ~w9247 & ~w9248;
assign w9250 = pi1269 & ~w4057;
assign w9251 = w4823 & ~w9250;
assign w9252 = pi1270 & w8490;
assign w9253 = pi1782 & w8492;
assign w9254 = ~w9252 & ~w9253;
assign w9255 = pi1775 & w8523;
assign w9256 = pi1271 & w8525;
assign w9257 = ~w9255 & ~w9256;
assign w9258 = pi1272 & w8490;
assign w9259 = pi1779 & w8492;
assign w9260 = ~w9258 & ~w9259;
assign w9261 = pi1785 & w8523;
assign w9262 = ~pi1273 & w8525;
assign w9263 = ~w9261 & ~w9262;
assign w9264 = pi1274 & w8490;
assign w9265 = pi1781 & w8492;
assign w9266 = ~w9264 & ~w9265;
assign w9267 = pi1275 & ~w4057;
assign w9268 = w4837 & ~w9267;
assign w9269 = pi1276 & ~w3151;
assign w9270 = w3883 & ~w9269;
assign w9271 = pi1277 & w8490;
assign w9272 = pi1777 & w8492;
assign w9273 = ~w9271 & ~w9272;
assign w9274 = ~pi1278 & ~w3954;
assign w9275 = w4149 & ~w9274;
assign w9276 = ~pi1279 & ~w3954;
assign w9277 = w4051 & ~w9276;
assign w9278 = pi1280 & w8490;
assign w9279 = pi1775 & w8492;
assign w9280 = ~w9278 & ~w9279;
assign w9281 = ~pi1281 & ~w3954;
assign w9282 = w5549 & ~w9281;
assign w9283 = ~pi1282 & ~w3954;
assign w9284 = w4749 & ~w9283;
assign w9285 = pi1283 & ~w4057;
assign w9286 = w5271 & ~w9285;
assign w9287 = ~pi1284 & ~w4057;
assign w9288 = w5247 & ~w9287;
assign w9289 = pi1285 & ~w3574;
assign w9290 = ~pi1738 & w3574;
assign w9291 = ~w9289 & ~w9290;
assign w9292 = pi1129 & w6627;
assign w9293 = pi1097 & w6639;
assign w9294 = ~pi0374 & w3188;
assign w9295 = ~pi0641 & w5442;
assign w9296 = pi0476 & w6633;
assign w9297 = pi1686 & w6641;
assign w9298 = ~pi0557 & w4056;
assign w9299 = pi1290 & w6615;
assign w9300 = ~pi0328 & w2932;
assign w9301 = ~pi0458 & w2866;
assign w9302 = pi0903 & w6629;
assign w9303 = ~pi0462 & w4186;
assign w9304 = pi0892 & w6609;
assign w9305 = pi1023 & w6620;
assign w9306 = pi1141 & w6622;
assign w9307 = ~pi0632 & w3953;
assign w9308 = pi0904 & w6624;
assign w9309 = ~pi0559 & w3150;
assign w9310 = pi1106 & w6612;
assign w9311 = pi0891 & w6618;
assign w9312 = pi1742 & w6606;
assign w9313 = ~w9292 & ~w9294;
assign w9314 = ~w9295 & ~w9298;
assign w9315 = ~w9300 & ~w9301;
assign w9316 = ~w9302 & ~w9303;
assign w9317 = ~w9304 & ~w9305;
assign w9318 = ~w9306 & ~w9307;
assign w9319 = ~w9308 & ~w9309;
assign w9320 = ~w9310 & ~w9311;
assign w9321 = w9319 & w9320;
assign w9322 = w9317 & w9318;
assign w9323 = w9315 & w9316;
assign w9324 = w9313 & w9314;
assign w9325 = ~w9293 & ~w9296;
assign w9326 = ~w9297 & ~w9299;
assign w9327 = ~w9312 & w9326;
assign w9328 = w9324 & w9325;
assign w9329 = w9322 & w9323;
assign w9330 = w9321 & w9329;
assign w9331 = w9327 & w9328;
assign w9332 = w9330 & w9331;
assign w9333 = w2868 & w6615;
assign w9334 = pi1747 & w9333;
assign w9335 = pi1782 & w9334;
assign w9336 = pi1747 & ~w9333;
assign w9337 = ~pi1287 & w9336;
assign w9338 = ~w9335 & ~w9337;
assign w9339 = pi1793 & w9334;
assign w9340 = ~pi1288 & w9336;
assign w9341 = ~w9339 & ~w9340;
assign w9342 = pi1776 & w9334;
assign w9343 = pi1289 & w9336;
assign w9344 = ~w9342 & ~w9343;
assign w9345 = pi1778 & w9334;
assign w9346 = pi1290 & w9336;
assign w9347 = ~w9345 & ~w9346;
assign w9348 = pi1774 & w9334;
assign w9349 = pi1291 & w9336;
assign w9350 = ~w9348 & ~w9349;
assign w9351 = ~pi1292 & ~w4057;
assign w9352 = w5263 & ~w9351;
assign w9353 = pi1123 & w6620;
assign w9354 = ~pi0538 & w4186;
assign w9355 = ~pi0685 & w5442;
assign w9356 = pi1148 & w6622;
assign w9357 = pi1117 & w6612;
assign w9358 = pi0251 & w6633;
assign w9359 = pi0644 & w6637;
assign w9360 = ~pi1327 & w6615;
assign w9361 = ~pi0493 & w3188;
assign w9362 = ~pi0600 & w4056;
assign w9363 = ~pi1391 & w6618;
assign w9364 = ~pi1379 & w6629;
assign w9365 = ~pi0341 & w2866;
assign w9366 = ~pi1388 & w6624;
assign w9367 = ~pi0524 & w3953;
assign w9368 = pi1135 & w6627;
assign w9369 = ~pi1351 & w6609;
assign w9370 = ~pi0395 & w2932;
assign w9371 = ~pi0418 & w3150;
assign w9372 = ~w9353 & ~w9354;
assign w9373 = ~w9355 & ~w9356;
assign w9374 = ~w9357 & ~w9361;
assign w9375 = ~w9362 & ~w9363;
assign w9376 = ~w9364 & ~w9365;
assign w9377 = ~w9366 & ~w9367;
assign w9378 = ~w9368 & ~w9369;
assign w9379 = ~w9370 & ~w9371;
assign w9380 = w9378 & w9379;
assign w9381 = w9376 & w9377;
assign w9382 = w9374 & w9375;
assign w9383 = w9372 & w9373;
assign w9384 = ~w9358 & ~w9359;
assign w9385 = ~w9360 & w9384;
assign w9386 = w9382 & w9383;
assign w9387 = w9380 & w9381;
assign w9388 = w9386 & w9387;
assign w9389 = w9385 & w9388;
assign w9390 = ~pi1394 & w6618;
assign w9391 = ~pi1397 & w6624;
assign w9392 = ~pi0489 & w3188;
assign w9393 = ~pi0681 & w5442;
assign w9394 = ~pi0517 & w2866;
assign w9395 = ~pi0572 & w4186;
assign w9396 = pi1024 & w6620;
assign w9397 = pi1145 & w6622;
assign w9398 = ~pi0391 & w2932;
assign w9399 = ~pi0521 & w3953;
assign w9400 = pi1114 & w6612;
assign w9401 = ~pi0595 & w4056;
assign w9402 = ~pi0414 & w3150;
assign w9403 = pi0269 & w6633;
assign w9404 = ~pi1377 & w6629;
assign w9405 = ~pi1324 & w6615;
assign w9406 = ~pi1078 & w6627;
assign w9407 = ~pi1357 & w6609;
assign w9408 = ~w9390 & ~w9391;
assign w9409 = ~w9392 & ~w9393;
assign w9410 = ~w9394 & ~w9395;
assign w9411 = ~w9396 & ~w9397;
assign w9412 = ~w9398 & ~w9399;
assign w9413 = ~w9400 & ~w9401;
assign w9414 = ~w9402 & ~w9404;
assign w9415 = ~w9406 & ~w9407;
assign w9416 = w9414 & w9415;
assign w9417 = w9412 & w9413;
assign w9418 = w9410 & w9411;
assign w9419 = w9408 & w9409;
assign w9420 = ~w9403 & ~w9405;
assign w9421 = w9419 & w9420;
assign w9422 = w9417 & w9418;
assign w9423 = w9416 & w9422;
assign w9424 = w9421 & w9423;
assign w9425 = ~pi1387 & w6624;
assign w9426 = pi1025 & w6620;
assign w9427 = ~pi0490 & w3188;
assign w9428 = ~pi0596 & w4056;
assign w9429 = pi1051 & w6612;
assign w9430 = ~pi1378 & w6629;
assign w9431 = ~pi0614 & w3150;
assign w9432 = ~pi1402 & w6618;
assign w9433 = ~pi1133 & w6627;
assign w9434 = ~pi0682 & w5442;
assign w9435 = pi1255 & w6622;
assign w9436 = ~pi1355 & w6609;
assign w9437 = ~pi0522 & w3953;
assign w9438 = ~pi1325 & w6615;
assign w9439 = ~pi0392 & w2932;
assign w9440 = pi0271 & w6633;
assign w9441 = ~pi0543 & w4186;
assign w9442 = ~pi0518 & w2866;
assign w9443 = ~w9425 & ~w9426;
assign w9444 = ~w9427 & ~w9428;
assign w9445 = ~w9429 & ~w9430;
assign w9446 = ~w9431 & ~w9432;
assign w9447 = ~w9433 & ~w9434;
assign w9448 = ~w9435 & ~w9436;
assign w9449 = ~w9437 & ~w9439;
assign w9450 = ~w9441 & ~w9442;
assign w9451 = w9449 & w9450;
assign w9452 = w9447 & w9448;
assign w9453 = w9445 & w9446;
assign w9454 = w9443 & w9444;
assign w9455 = ~w9438 & ~w9440;
assign w9456 = w9454 & w9455;
assign w9457 = w9452 & w9453;
assign w9458 = w9451 & w9457;
assign w9459 = w9456 & w9458;
assign w9460 = ~pi1405 & w6629;
assign w9461 = pi1054 & w6627;
assign w9462 = pi1115 & w6612;
assign w9463 = ~pi0671 & w5442;
assign w9464 = ~pi0523 & w3953;
assign w9465 = ~pi0415 & w3150;
assign w9466 = ~pi0597 & w4056;
assign w9467 = ~pi0338 & w2866;
assign w9468 = ~pi0573 & w4186;
assign w9469 = ~pi0430 & w2932;
assign w9470 = ~pi0491 & w3188;
assign w9471 = ~pi1408 & w6618;
assign w9472 = ~pi1350 & w6609;
assign w9473 = ~pi1326 & w6615;
assign w9474 = ~pi1395 & w6624;
assign w9475 = pi0272 & w6633;
assign w9476 = pi1026 & w6620;
assign w9477 = pi1146 & w6622;
assign w9478 = ~w9460 & ~w9461;
assign w9479 = ~w9462 & ~w9463;
assign w9480 = ~w9464 & ~w9465;
assign w9481 = ~w9466 & ~w9467;
assign w9482 = ~w9468 & ~w9469;
assign w9483 = ~w9470 & ~w9471;
assign w9484 = ~w9472 & ~w9474;
assign w9485 = ~w9476 & ~w9477;
assign w9486 = w9484 & w9485;
assign w9487 = w9482 & w9483;
assign w9488 = w9480 & w9481;
assign w9489 = w9478 & w9479;
assign w9490 = ~w9473 & ~w9475;
assign w9491 = w9489 & w9490;
assign w9492 = w9487 & w9488;
assign w9493 = w9486 & w9492;
assign w9494 = w9491 & w9493;
assign w9495 = pi1253 & w6622;
assign w9496 = pi1260 & w6620;
assign w9497 = ~pi0416 & w3150;
assign w9498 = ~pi0598 & w4056;
assign w9499 = ~pi0444 & w3953;
assign w9500 = pi1134 & w6627;
assign w9501 = ~pi1380 & w6629;
assign w9502 = pi1116 & w6612;
assign w9503 = ~pi0492 & w3188;
assign w9504 = ~pi1389 & w6624;
assign w9505 = ~pi1411 & w6618;
assign w9506 = ~pi0393 & w2932;
assign w9507 = ~pi1354 & w6609;
assign w9508 = pi0270 & w6633;
assign w9509 = ~pi0574 & w4186;
assign w9510 = ~pi1288 & w6615;
assign w9511 = ~pi0339 & w2866;
assign w9512 = ~pi0683 & w5442;
assign w9513 = ~w9495 & ~w9496;
assign w9514 = ~w9497 & ~w9498;
assign w9515 = ~w9499 & ~w9500;
assign w9516 = ~w9501 & ~w9502;
assign w9517 = ~w9503 & ~w9504;
assign w9518 = ~w9505 & ~w9506;
assign w9519 = ~w9507 & ~w9509;
assign w9520 = ~w9511 & ~w9512;
assign w9521 = w9519 & w9520;
assign w9522 = w9517 & w9518;
assign w9523 = w9515 & w9516;
assign w9524 = w9513 & w9514;
assign w9525 = ~w9508 & ~w9510;
assign w9526 = w9524 & w9525;
assign w9527 = w9522 & w9523;
assign w9528 = w9521 & w9527;
assign w9529 = w9526 & w9528;
assign w9530 = ~pi1347 & w6609;
assign w9531 = ~pi1393 & w6624;
assign w9532 = ~pi0578 & w4186;
assign w9533 = ~pi0656 & w3953;
assign w9534 = ~pi0419 & w3150;
assign w9535 = pi0263 & w6633;
assign w9536 = pi0987 & w6637;
assign w9537 = ~pi1328 & w6615;
assign w9538 = ~pi0494 & w3188;
assign w9539 = ~pi0668 & w5442;
assign w9540 = pi1262 & w6620;
assign w9541 = pi1070 & w6612;
assign w9542 = pi1136 & w6627;
assign w9543 = ~pi0342 & w2866;
assign w9544 = pi1147 & w6622;
assign w9545 = ~pi1412 & w6618;
assign w9546 = ~pi0378 & w2932;
assign w9547 = ~pi0546 & w4056;
assign w9548 = ~pi1403 & w6629;
assign w9549 = ~w9530 & ~w9531;
assign w9550 = ~w9532 & ~w9533;
assign w9551 = ~w9534 & ~w9538;
assign w9552 = ~w9539 & ~w9540;
assign w9553 = ~w9541 & ~w9542;
assign w9554 = ~w9543 & ~w9544;
assign w9555 = ~w9545 & ~w9546;
assign w9556 = ~w9547 & ~w9548;
assign w9557 = w9555 & w9556;
assign w9558 = w9553 & w9554;
assign w9559 = w9551 & w9552;
assign w9560 = w9549 & w9550;
assign w9561 = ~w9535 & ~w9536;
assign w9562 = ~w9537 & w9561;
assign w9563 = w9559 & w9560;
assign w9564 = w9557 & w9558;
assign w9565 = w9563 & w9564;
assign w9566 = w9562 & w9565;
assign w9567 = ~pi0397 & w2932;
assign w9568 = ~pi1359 & w6618;
assign w9569 = pi1242 & w6622;
assign w9570 = ~pi1404 & w6624;
assign w9571 = ~pi0496 & w3188;
assign w9572 = pi0915 & w6637;
assign w9573 = pi0253 & w6633;
assign w9574 = ~pi1330 & w6615;
assign w9575 = pi1124 & w6620;
assign w9576 = ~pi1381 & w6609;
assign w9577 = ~pi0688 & w5442;
assign w9578 = ~pi0603 & w4056;
assign w9579 = ~pi0421 & w3150;
assign w9580 = ~pi1137 & w6627;
assign w9581 = ~pi1400 & w6629;
assign w9582 = pi1118 & w6612;
assign w9583 = ~pi0344 & w2866;
assign w9584 = ~pi0526 & w3953;
assign w9585 = ~pi0540 & w4186;
assign w9586 = ~w9567 & ~w9568;
assign w9587 = ~w9569 & ~w9570;
assign w9588 = ~w9571 & ~w9575;
assign w9589 = ~w9576 & ~w9577;
assign w9590 = ~w9578 & ~w9579;
assign w9591 = ~w9580 & ~w9581;
assign w9592 = ~w9582 & ~w9583;
assign w9593 = ~w9584 & ~w9585;
assign w9594 = w9592 & w9593;
assign w9595 = w9590 & w9591;
assign w9596 = w9588 & w9589;
assign w9597 = w9586 & w9587;
assign w9598 = ~w9572 & ~w9573;
assign w9599 = ~w9574 & w9598;
assign w9600 = w9596 & w9597;
assign w9601 = w9594 & w9595;
assign w9602 = w9600 & w9601;
assign w9603 = w9599 & w9602;
assign w9604 = ~pi0345 & w2866;
assign w9605 = ~pi1363 & w6609;
assign w9606 = pi1261 & w6622;
assign w9607 = ~pi0527 & w3953;
assign w9608 = pi1074 & w6612;
assign w9609 = ~pi0497 & w3188;
assign w9610 = ~pi0580 & w4186;
assign w9611 = ~pi1383 & w6624;
assign w9612 = ~pi0544 & w4056;
assign w9613 = ~pi0422 & w3150;
assign w9614 = ~pi0398 & w2932;
assign w9615 = ~pi0667 & w5442;
assign w9616 = ~pi1030 & w6627;
assign w9617 = pi0255 & w6633;
assign w9618 = ~pi1374 & w6629;
assign w9619 = pi0901 & w6637;
assign w9620 = ~pi1362 & w6618;
assign w9621 = pi1252 & w6620;
assign w9622 = ~w9604 & ~w9605;
assign w9623 = ~w9606 & ~w9607;
assign w9624 = ~w9608 & ~w9609;
assign w9625 = ~w9610 & ~w9611;
assign w9626 = ~w9612 & ~w9613;
assign w9627 = ~w9614 & ~w9615;
assign w9628 = ~w9616 & ~w9618;
assign w9629 = ~w9620 & ~w9621;
assign w9630 = w9628 & w9629;
assign w9631 = w9626 & w9627;
assign w9632 = w9624 & w9625;
assign w9633 = w9622 & w9623;
assign w9634 = ~w9617 & ~w9619;
assign w9635 = w9633 & w9634;
assign w9636 = w9631 & w9632;
assign w9637 = w9630 & w9636;
assign w9638 = w9635 & w9637;
assign w9639 = ~pi1390 & w6618;
assign w9640 = ~pi1406 & w6629;
assign w9641 = ~pi0401 & w2932;
assign w9642 = pi1144 & w6622;
assign w9643 = ~pi0579 & w4186;
assign w9644 = ~pi0498 & w3188;
assign w9645 = ~pi1384 & w6624;
assign w9646 = pi1112 & w6612;
assign w9647 = ~pi0690 & w5442;
assign w9648 = ~pi0346 & w2866;
assign w9649 = ~pi0432 & w3150;
assign w9650 = ~pi0606 & w4056;
assign w9651 = ~pi1382 & w6609;
assign w9652 = pi0728 & w6637;
assign w9653 = pi1080 & w6627;
assign w9654 = pi0250 & w6633;
assign w9655 = ~pi0629 & w3953;
assign w9656 = pi1256 & w6620;
assign w9657 = ~w9639 & ~w9640;
assign w9658 = ~w9641 & ~w9642;
assign w9659 = ~w9643 & ~w9644;
assign w9660 = ~w9645 & ~w9646;
assign w9661 = ~w9647 & ~w9648;
assign w9662 = ~w9649 & ~w9650;
assign w9663 = ~w9651 & ~w9653;
assign w9664 = ~w9655 & ~w9656;
assign w9665 = w9663 & w9664;
assign w9666 = w9661 & w9662;
assign w9667 = w9659 & w9660;
assign w9668 = w9657 & w9658;
assign w9669 = ~w9652 & ~w9654;
assign w9670 = w9668 & w9669;
assign w9671 = w9666 & w9667;
assign w9672 = w9665 & w9671;
assign w9673 = w9670 & w9672;
assign w9674 = ~pi0350 & w3150;
assign w9675 = ~pi0651 & w5442;
assign w9676 = ~pi0504 & w4186;
assign w9677 = pi0863 & w6620;
assign w9678 = ~pi1396 & w6624;
assign w9679 = ~pi1353 & w6609;
assign w9680 = pi0969 & w6622;
assign w9681 = ~pi0427 & w3953;
assign w9682 = ~pi0334 & w2932;
assign w9683 = pi0994 & w6612;
assign w9684 = ~pi0515 & w4056;
assign w9685 = ~pi0311 & w2866;
assign w9686 = ~pi0406 & w3188;
assign w9687 = pi0977 & w6637;
assign w9688 = pi0939 & w6627;
assign w9689 = pi0186 & w6633;
assign w9690 = ~pi1407 & w6629;
assign w9691 = ~pi1349 & w6618;
assign w9692 = ~w9674 & ~w9675;
assign w9693 = ~w9676 & ~w9677;
assign w9694 = ~w9678 & ~w9679;
assign w9695 = ~w9680 & ~w9681;
assign w9696 = ~w9682 & ~w9683;
assign w9697 = ~w9684 & ~w9685;
assign w9698 = ~w9686 & ~w9688;
assign w9699 = ~w9690 & ~w9691;
assign w9700 = w9698 & w9699;
assign w9701 = w9696 & w9697;
assign w9702 = w9694 & w9695;
assign w9703 = w9692 & w9693;
assign w9704 = ~w9687 & ~w9689;
assign w9705 = w9703 & w9704;
assign w9706 = w9701 & w9702;
assign w9707 = w9700 & w9706;
assign w9708 = w9705 & w9707;
assign w9709 = ~pi0548 & w3150;
assign w9710 = ~pi0376 & w3188;
assign w9711 = ~pi0463 & w4186;
assign w9712 = pi1028 & w6627;
assign w9713 = pi1107 & w6612;
assign w9714 = pi1321 & w6615;
assign w9715 = pi1068 & w6639;
assign w9716 = pi0477 & w6633;
assign w9717 = pi1681 & w6641;
assign w9718 = ~pi0447 & w2866;
assign w9719 = pi0131 & w6618;
assign w9720 = pi0130 & w6624;
assign w9721 = ~pi0329 & w2932;
assign w9722 = pi1272 & w6620;
assign w9723 = pi0128 & w6629;
assign w9724 = ~pi0547 & w4056;
assign w9725 = pi1258 & w6622;
assign w9726 = ~pi0628 & w5442;
assign w9727 = pi0129 & w6609;
assign w9728 = ~pi0640 & w3953;
assign w9729 = ~w9709 & ~w9710;
assign w9730 = ~w9711 & ~w9712;
assign w9731 = ~w9713 & ~w9718;
assign w9732 = ~w9719 & ~w9720;
assign w9733 = ~w9721 & ~w9722;
assign w9734 = ~w9723 & ~w9724;
assign w9735 = ~w9725 & ~w9726;
assign w9736 = ~w9727 & ~w9728;
assign w9737 = w9735 & w9736;
assign w9738 = w9733 & w9734;
assign w9739 = w9731 & w9732;
assign w9740 = w9729 & w9730;
assign w9741 = ~w9714 & ~w9715;
assign w9742 = ~w9716 & ~w9717;
assign w9743 = w9741 & w9742;
assign w9744 = w9739 & w9740;
assign w9745 = w9737 & w9738;
assign w9746 = w9744 & w9745;
assign w9747 = w9743 & w9746;
assign w9748 = pi1083 & w6627;
assign w9749 = pi1121 & w6620;
assign w9750 = pi1108 & w6612;
assign w9751 = pi0990 & w6618;
assign w9752 = ~pi0321 & w2866;
assign w9753 = pi1322 & w6615;
assign w9754 = pi0448 & w6633;
assign w9755 = pi1098 & w6639;
assign w9756 = pi1693 & w6641;
assign w9757 = pi1033 & w6622;
assign w9758 = ~pi0633 & w5442;
assign w9759 = ~pi0449 & w3953;
assign w9760 = pi1314 & w6609;
assign w9761 = ~pi0461 & w4186;
assign w9762 = ~pi0550 & w4056;
assign w9763 = pi0965 & w6624;
assign w9764 = ~pi0362 & w3150;
assign w9765 = pi1048 & w6629;
assign w9766 = ~pi0327 & w2932;
assign w9767 = ~pi0357 & w3188;
assign w9768 = ~w9748 & ~w9749;
assign w9769 = ~w9750 & ~w9751;
assign w9770 = ~w9752 & ~w9757;
assign w9771 = ~w9758 & ~w9759;
assign w9772 = ~w9760 & ~w9761;
assign w9773 = ~w9762 & ~w9763;
assign w9774 = ~w9764 & ~w9765;
assign w9775 = ~w9766 & ~w9767;
assign w9776 = w9774 & w9775;
assign w9777 = w9772 & w9773;
assign w9778 = w9770 & w9771;
assign w9779 = w9768 & w9769;
assign w9780 = ~w9753 & ~w9754;
assign w9781 = ~w9755 & ~w9756;
assign w9782 = w9780 & w9781;
assign w9783 = w9778 & w9779;
assign w9784 = w9776 & w9777;
assign w9785 = w9783 & w9784;
assign w9786 = w9782 & w9785;
assign w9787 = ~pi1305 & ~w4057;
assign w9788 = w5239 & ~w9787;
assign w9789 = ~w8010 & ~w8043;
assign w9790 = ~w8011 & ~w8042;
assign w9791 = w9789 & w9790;
assign w9792 = ~w9789 & ~w9790;
assign w9793 = ~w9791 & ~w9792;
assign w9794 = ~w8054 & ~w8088;
assign w9795 = ~w8055 & ~w8087;
assign w9796 = w9794 & w9795;
assign w9797 = ~w9794 & ~w9795;
assign w9798 = ~w9796 & ~w9797;
assign w9799 = ~pi0560 & w8145;
assign w9800 = pi0560 & w8143;
assign w9801 = ~w8147 & ~w9800;
assign w9802 = ~w9799 & ~w9801;
assign w9803 = ~w8159 & ~w8192;
assign w9804 = ~w8160 & ~w8191;
assign w9805 = w9803 & w9804;
assign w9806 = ~w9803 & ~w9804;
assign w9807 = ~w9805 & ~w9806;
assign w9808 = pi1310 & w8508;
assign w9809 = pi1777 & w8510;
assign w9810 = ~w9808 & ~w9809;
assign w9811 = ~pi1311 & ~w4057;
assign w9812 = w4963 & ~w9811;
assign w9813 = ~pi1312 & ~w4057;
assign w9814 = w4955 & ~w9813;
assign w9815 = pi1313 & ~w3574;
assign w9816 = ~pi1733 & w3574;
assign w9817 = ~w9815 & ~w9816;
assign w9818 = pi1480 & pi1729;
assign w9819 = ~pi1314 & ~w9818;
assign w9820 = w1773 & ~w9819;
assign w9821 = ~pi1316 & ~w4057;
assign w9822 = w4887 & ~w9821;
assign w9823 = pi1317 & ~w3574;
assign w9824 = ~pi1741 & w3574;
assign w9825 = ~w9823 & ~w9824;
assign w9826 = pi1318 & ~w3574;
assign w9827 = ~pi1722 & w3574;
assign w9828 = ~w9826 & ~w9827;
assign w9829 = pi1775 & w9334;
assign w9830 = pi1319 & w9336;
assign w9831 = ~w9829 & ~w9830;
assign w9832 = pi1777 & w9334;
assign w9833 = pi1320 & w9336;
assign w9834 = ~w9832 & ~w9833;
assign w9835 = pi1779 & w9334;
assign w9836 = pi1321 & w9336;
assign w9837 = ~w9835 & ~w9836;
assign w9838 = pi1780 & w9334;
assign w9839 = pi1322 & w9336;
assign w9840 = ~w9838 & ~w9839;
assign w9841 = pi1781 & w9334;
assign w9842 = ~pi1323 & w9336;
assign w9843 = ~w9841 & ~w9842;
assign w9844 = pi1790 & w9334;
assign w9845 = ~pi1324 & w9336;
assign w9846 = ~w9844 & ~w9845;
assign w9847 = pi1791 & w9334;
assign w9848 = ~pi1325 & w9336;
assign w9849 = ~w9847 & ~w9848;
assign w9850 = pi1792 & w9334;
assign w9851 = ~pi1326 & w9336;
assign w9852 = ~w9850 & ~w9851;
assign w9853 = pi1794 & w9334;
assign w9854 = ~pi1327 & w9336;
assign w9855 = ~w9853 & ~w9854;
assign w9856 = pi1795 & w9334;
assign w9857 = ~pi1328 & w9336;
assign w9858 = ~w9856 & ~w9857;
assign w9859 = pi1796 & w9334;
assign w9860 = ~pi1329 & w9336;
assign w9861 = ~w9859 & ~w9860;
assign w9862 = pi1798 & w9334;
assign w9863 = ~pi1330 & w9336;
assign w9864 = ~w9862 & ~w9863;
assign w9865 = pi1331 & ~w4057;
assign w9866 = w5255 & ~w9865;
assign w9867 = ~pi1332 & ~w4057;
assign w9868 = w4979 & ~w9867;
assign w9869 = ~pi1333 & ~w4057;
assign w9870 = w4987 & ~w9869;
assign w9871 = pi1334 & ~w3574;
assign w9872 = ~pi1727 & w3574;
assign w9873 = ~w9871 & ~w9872;
assign w9874 = pi1335 & ~w3574;
assign w9875 = ~pi1740 & w3574;
assign w9876 = ~w9874 & ~w9875;
assign w9877 = pi1336 & ~w3574;
assign w9878 = ~pi1735 & w3574;
assign w9879 = ~w9877 & ~w9878;
assign w9880 = pi1337 & ~w3574;
assign w9881 = ~pi1725 & w3574;
assign w9882 = ~w9880 & ~w9881;
assign w9883 = pi1338 & w8589;
assign w9884 = pi1777 & w8591;
assign w9885 = ~w9883 & ~w9884;
assign w9886 = pi1797 & w9334;
assign w9887 = ~pi1339 & w9336;
assign w9888 = ~w9886 & ~w9887;
assign w9889 = (~w8091 & w12983) | (~w8091 & w12984) | (w12983 & w12984);
assign w9890 = pi0383 & ~pi1179;
assign w9891 = ~pi0383 & pi1179;
assign w9892 = ~w9890 & ~w9891;
assign w9893 = w9889 & w9892;
assign w9894 = ~w9889 & ~w9892;
assign w9895 = ~w9893 & ~w9894;
assign w9896 = ~w8105 & ~w8108;
assign w9897 = ~w8105 & w8148;
assign w9898 = ~w8106 & ~w9897;
assign w9899 = (w9898 & ~w8147) | (w9898 & w12973) | (~w8147 & w12973);
assign w9900 = pi0471 & ~pi1036;
assign w9901 = ~pi0471 & pi1036;
assign w9902 = ~w9900 & ~w9901;
assign w9903 = w9899 & w9902;
assign w9904 = ~w9899 & ~w9902;
assign w9905 = ~w9903 & ~w9904;
assign w9906 = pi1777 & w8523;
assign w9907 = pi1342 & w8525;
assign w9908 = ~w9906 & ~w9907;
assign w9909 = ~pi1343 & ~w4057;
assign w9910 = w4879 & ~w9909;
assign w9911 = ~pi1344 & ~w4057;
assign w9912 = w5327 & ~w9911;
assign w9913 = ~pi1345 & ~pi1495;
assign w9914 = pi1345 & pi1495;
assign w9915 = pi1479 & ~w2132;
assign w9916 = ~pi1479 & ~w6396;
assign w9917 = ~w9915 & ~w9916;
assign w9918 = ~w9914 & ~w9917;
assign w9919 = pi1747 & ~w9913;
assign w9920 = ~w9918 & w9919;
assign w9921 = pi1346 & ~w4057;
assign w9922 = w5311 & ~w9921;
assign w9923 = w2868 & w6609;
assign w9924 = pi1747 & w9923;
assign w9925 = pi1795 & w9924;
assign w9926 = pi1747 & ~w9923;
assign w9927 = ~pi1347 & w9926;
assign w9928 = ~w9925 & ~w9927;
assign w9929 = pi1801 & w9924;
assign w9930 = ~pi1348 & w9926;
assign w9931 = ~w9929 & ~w9930;
assign w9932 = w2868 & w6618;
assign w9933 = pi1747 & w9932;
assign w9934 = pi1802 & w9933;
assign w9935 = pi1747 & ~w9932;
assign w9936 = ~pi1349 & w9935;
assign w9937 = ~w9934 & ~w9936;
assign w9938 = pi1792 & w9924;
assign w9939 = ~pi1350 & w9926;
assign w9940 = ~w9938 & ~w9939;
assign w9941 = pi1794 & w9924;
assign w9942 = ~pi1351 & w9926;
assign w9943 = ~w9941 & ~w9942;
assign w9944 = pi1803 & w9933;
assign w9945 = ~pi1352 & w9935;
assign w9946 = ~w9944 & ~w9945;
assign w9947 = pi1802 & w9924;
assign w9948 = ~pi1353 & w9926;
assign w9949 = ~w9947 & ~w9948;
assign w9950 = pi1793 & w9924;
assign w9951 = ~pi1354 & w9926;
assign w9952 = ~w9950 & ~w9951;
assign w9953 = pi1791 & w9924;
assign w9954 = ~pi1355 & w9926;
assign w9955 = ~w9953 & ~w9954;
assign w9956 = pi1803 & w9924;
assign w9957 = ~pi1356 & w9926;
assign w9958 = ~w9956 & ~w9957;
assign w9959 = pi1790 & w9924;
assign w9960 = ~pi1357 & w9926;
assign w9961 = ~w9959 & ~w9960;
assign w9962 = pi0103 & ~w1345;
assign w9963 = ~w1512 & ~w9962;
assign w9964 = pi1798 & w9933;
assign w9965 = ~pi1359 & w9935;
assign w9966 = ~w9964 & ~w9965;
assign w9967 = pi1360 & ~w9051;
assign w9968 = w8490 & ~w9967;
assign w9969 = pi1796 & w8492;
assign w9970 = ~w9968 & ~w9969;
assign w9971 = pi1361 & ~w9007;
assign w9972 = w8589 & ~w9971;
assign w9973 = pi1796 & w8591;
assign w9974 = ~w9972 & ~w9973;
assign w9975 = pi1799 & w9933;
assign w9976 = ~pi1362 & w9935;
assign w9977 = ~w9975 & ~w9976;
assign w9978 = pi1799 & w9924;
assign w9979 = ~pi1363 & w9926;
assign w9980 = ~w9978 & ~w9979;
assign w9981 = pi1801 & w9933;
assign w9982 = ~pi1364 & w9935;
assign w9983 = ~w9981 & ~w9982;
assign w9984 = ~pi1356 & w6609;
assign w9985 = pi0876 & w6620;
assign w9986 = pi1014 & w6612;
assign w9987 = ~pi1386 & w6624;
assign w9988 = ~pi0377 & w2932;
assign w9989 = ~pi0519 & w2866;
assign w9990 = ~pi0542 & w4056;
assign w9991 = pi0153 & w6633;
assign w9992 = ~pi1352 & w6618;
assign w9993 = ~pi1376 & w6629;
assign w9994 = ~pi0704 & w5442;
assign w9995 = pi0942 & w6627;
assign w9996 = ~pi0528 & w3953;
assign w9997 = pi0973 & w6622;
assign w9998 = ~pi0501 & w3188;
assign w9999 = ~pi0616 & w3150;
assign w10000 = ~pi0581 & w4186;
assign w10001 = ~w9984 & ~w9985;
assign w10002 = ~w9986 & ~w9987;
assign w10003 = ~w9988 & ~w9989;
assign w10004 = ~w9990 & ~w9992;
assign w10005 = ~w9993 & ~w9994;
assign w10006 = ~w9995 & ~w9996;
assign w10007 = ~w9997 & ~w9998;
assign w10008 = ~w9999 & ~w10000;
assign w10009 = w10007 & w10008;
assign w10010 = w10005 & w10006;
assign w10011 = w10003 & w10004;
assign w10012 = w10001 & w10002;
assign w10013 = ~w9991 & w10012;
assign w10014 = w10010 & w10011;
assign w10015 = w10009 & w10014;
assign w10016 = w10013 & w10015;
assign w10017 = ~pi0530 & w3953;
assign w10018 = ~pi0347 & w2866;
assign w10019 = pi0967 & w6622;
assign w10020 = pi0938 & w6627;
assign w10021 = ~pi0500 & w3188;
assign w10022 = ~pi0608 & w4056;
assign w10023 = ~pi0424 & w3150;
assign w10024 = ~pi0691 & w5442;
assign w10025 = pi0861 & w6620;
assign w10026 = pi0195 & w6633;
assign w10027 = ~pi0403 & w2932;
assign w10028 = ~pi0583 & w4186;
assign w10029 = pi0992 & w6612;
assign w10030 = ~w10017 & ~w10018;
assign w10031 = ~w10019 & ~w10020;
assign w10032 = ~w10021 & ~w10022;
assign w10033 = ~w10023 & ~w10024;
assign w10034 = ~w10025 & ~w10027;
assign w10035 = ~w10028 & ~w10029;
assign w10036 = w10034 & w10035;
assign w10037 = w10032 & w10033;
assign w10038 = w10030 & w10031;
assign w10039 = ~w10026 & w10038;
assign w10040 = w10036 & w10037;
assign w10041 = w10039 & w10040;
assign w10042 = ~pi0428 & w3953;
assign w10043 = pi0993 & w6612;
assign w10044 = pi0862 & w6620;
assign w10045 = ~pi0407 & w3188;
assign w10046 = ~pi0351 & w3150;
assign w10047 = ~pi0437 & w4056;
assign w10048 = ~pi0505 & w4186;
assign w10049 = ~pi0335 & w2932;
assign w10050 = ~pi0652 & w5442;
assign w10051 = pi0185 & w6633;
assign w10052 = pi0968 & w6622;
assign w10053 = pi0941 & w6627;
assign w10054 = ~pi0312 & w2866;
assign w10055 = ~w10042 & ~w10043;
assign w10056 = ~w10044 & ~w10045;
assign w10057 = ~w10046 & ~w10047;
assign w10058 = ~w10048 & ~w10049;
assign w10059 = ~w10050 & ~w10052;
assign w10060 = ~w10053 & ~w10054;
assign w10061 = w10059 & w10060;
assign w10062 = w10057 & w10058;
assign w10063 = w10055 & w10056;
assign w10064 = ~w10051 & w10063;
assign w10065 = w10061 & w10062;
assign w10066 = w10064 & w10065;
assign w10067 = ~pi0445 & w3188;
assign w10068 = ~pi0605 & w4056;
assign w10069 = ~pi0314 & w2866;
assign w10070 = ~pi0423 & w3150;
assign w10071 = ~pi1348 & w6609;
assign w10072 = ~pi1364 & w6618;
assign w10073 = pi1113 & w6612;
assign w10074 = pi0986 & w6637;
assign w10075 = ~pi0658 & w3953;
assign w10076 = pi1132 & w6627;
assign w10077 = ~pi1385 & w6624;
assign w10078 = pi1259 & w6622;
assign w10079 = ~pi0689 & w5442;
assign w10080 = ~pi0400 & w2932;
assign w10081 = ~pi1375 & w6629;
assign w10082 = pi1257 & w6620;
assign w10083 = ~pi0539 & w4186;
assign w10084 = ~w10067 & ~w10068;
assign w10085 = ~w10069 & ~w10070;
assign w10086 = ~w10071 & ~w10072;
assign w10087 = ~w10073 & ~w10075;
assign w10088 = ~w10076 & ~w10077;
assign w10089 = ~w10078 & ~w10079;
assign w10090 = ~w10080 & ~w10081;
assign w10091 = ~w10082 & ~w10083;
assign w10092 = w10090 & w10091;
assign w10093 = w10088 & w10089;
assign w10094 = w10086 & w10087;
assign w10095 = w10084 & w10085;
assign w10096 = ~w10074 & w10095;
assign w10097 = w10093 & w10094;
assign w10098 = w10092 & w10097;
assign w10099 = w10096 & w10098;
assign w10100 = pi1369 & ~w9098;
assign w10101 = w8508 & ~w10100;
assign w10102 = pi1796 & w8510;
assign w10103 = ~w10101 & ~w10102;
assign w10104 = w8793 & ~w8794;
assign w10105 = pi1088 & pi1101;
assign w10106 = w13 & w10105;
assign w10107 = ~w10104 & ~w10106;
assign w10108 = w1755 & ~w10107;
assign w10109 = pi1119 & w6620;
assign w10110 = pi1102 & w6612;
assign w10111 = pi1127 & w6627;
assign w10112 = ~pi0316 & w2866;
assign w10113 = ~pi0636 & w5442;
assign w10114 = pi1139 & w6622;
assign w10115 = ~pi0322 & w2932;
assign w10116 = ~pi0369 & w3188;
assign w10117 = ~pi0456 & w4186;
assign w10118 = pi0473 & w6633;
assign w10119 = ~pi0451 & w3953;
assign w10120 = ~pi0551 & w4056;
assign w10121 = ~pi0364 & w3150;
assign w10122 = ~w10109 & ~w10110;
assign w10123 = ~w10111 & ~w10112;
assign w10124 = ~w10113 & ~w10114;
assign w10125 = ~w10115 & ~w10116;
assign w10126 = ~w10117 & ~w10119;
assign w10127 = ~w10120 & ~w10121;
assign w10128 = w10126 & w10127;
assign w10129 = w10124 & w10125;
assign w10130 = w10122 & w10123;
assign w10131 = ~w10118 & w10130;
assign w10132 = w10128 & w10129;
assign w10133 = w10131 & w10132;
assign w10134 = ~pi1268 & w6620;
assign w10135 = ~pi0372 & w3188;
assign w10136 = ~pi1243 & w6612;
assign w10137 = ~pi0325 & w2932;
assign w10138 = ~pi1273 & w6622;
assign w10139 = ~pi0319 & w2866;
assign w10140 = ~pi0460 & w4186;
assign w10141 = ~pi0367 & w3150;
assign w10142 = ~pi0555 & w4056;
assign w10143 = ~pi0465 & w6633;
assign w10144 = ~pi0638 & w5442;
assign w10145 = ~pi1128 & w6627;
assign w10146 = ~pi0450 & w3953;
assign w10147 = ~w10134 & ~w10135;
assign w10148 = ~w10136 & ~w10137;
assign w10149 = ~w10138 & ~w10139;
assign w10150 = ~w10140 & ~w10141;
assign w10151 = ~w10142 & ~w10144;
assign w10152 = ~w10145 & ~w10146;
assign w10153 = w10151 & w10152;
assign w10154 = w10149 & w10150;
assign w10155 = w10147 & w10148;
assign w10156 = ~w10143 & w10155;
assign w10157 = w10153 & w10154;
assign w10158 = w10156 & w10157;
assign w10159 = ~pi0693 & w5442;
assign w10160 = pi1034 & w6622;
assign w10161 = pi1110 & w6612;
assign w10162 = ~pi0659 & w3953;
assign w10163 = ~pi0443 & w3188;
assign w10164 = ~pi0405 & w2932;
assign w10165 = ~pi0611 & w4056;
assign w10166 = pi1029 & w6627;
assign w10167 = ~pi0426 & w3150;
assign w10168 = pi0478 & w6633;
assign w10169 = ~pi0313 & w2866;
assign w10170 = pi1267 & w6620;
assign w10171 = ~pi0585 & w4186;
assign w10172 = ~w10159 & ~w10160;
assign w10173 = ~w10161 & ~w10162;
assign w10174 = ~w10163 & ~w10164;
assign w10175 = ~w10165 & ~w10166;
assign w10176 = ~w10167 & ~w10169;
assign w10177 = ~w10170 & ~w10171;
assign w10178 = w10176 & w10177;
assign w10179 = w10174 & w10175;
assign w10180 = w10172 & w10173;
assign w10181 = ~w10168 & w10180;
assign w10182 = w10178 & w10179;
assign w10183 = w10181 & w10182;
assign w10184 = w2868 & w6629;
assign w10185 = pi1747 & w10184;
assign w10186 = pi1799 & w10185;
assign w10187 = pi1747 & ~w10184;
assign w10188 = ~pi1374 & w10187;
assign w10189 = ~w10186 & ~w10188;
assign w10190 = pi1801 & w10185;
assign w10191 = ~pi1375 & w10187;
assign w10192 = ~w10190 & ~w10191;
assign w10193 = pi1803 & w10185;
assign w10194 = ~pi1376 & w10187;
assign w10195 = ~w10193 & ~w10194;
assign w10196 = pi1790 & w10185;
assign w10197 = ~pi1377 & w10187;
assign w10198 = ~w10196 & ~w10197;
assign w10199 = pi1791 & w10185;
assign w10200 = ~pi1378 & w10187;
assign w10201 = ~w10199 & ~w10200;
assign w10202 = pi1794 & w10185;
assign w10203 = ~pi1379 & w10187;
assign w10204 = ~w10202 & ~w10203;
assign w10205 = pi1793 & w10185;
assign w10206 = ~pi1380 & w10187;
assign w10207 = ~w10205 & ~w10206;
assign w10208 = pi1798 & w9924;
assign w10209 = ~pi1381 & w9926;
assign w10210 = ~w10208 & ~w10209;
assign w10211 = pi1800 & w9924;
assign w10212 = ~pi1382 & w9926;
assign w10213 = ~w10211 & ~w10212;
assign w10214 = w2868 & w6624;
assign w10215 = pi1747 & w10214;
assign w10216 = pi1799 & w10215;
assign w10217 = pi1747 & ~w10214;
assign w10218 = ~pi1383 & w10217;
assign w10219 = ~w10216 & ~w10218;
assign w10220 = pi1800 & w10215;
assign w10221 = ~pi1384 & w10217;
assign w10222 = ~w10220 & ~w10221;
assign w10223 = pi1801 & w10215;
assign w10224 = ~pi1385 & w10217;
assign w10225 = ~w10223 & ~w10224;
assign w10226 = pi1803 & w10215;
assign w10227 = ~pi1386 & w10217;
assign w10228 = ~w10226 & ~w10227;
assign w10229 = pi1791 & w10215;
assign w10230 = ~pi1387 & w10217;
assign w10231 = ~w10229 & ~w10230;
assign w10232 = pi1794 & w10215;
assign w10233 = ~pi1388 & w10217;
assign w10234 = ~w10232 & ~w10233;
assign w10235 = pi1793 & w10215;
assign w10236 = ~pi1389 & w10217;
assign w10237 = ~w10235 & ~w10236;
assign w10238 = pi1800 & w9933;
assign w10239 = ~pi1390 & w9935;
assign w10240 = ~w10238 & ~w10239;
assign w10241 = pi1794 & w9933;
assign w10242 = ~pi1391 & w9935;
assign w10243 = ~w10241 & ~w10242;
assign w10244 = ~pi0571 & w4186;
assign w10245 = ~pi0680 & w5442;
assign w10246 = ~pi1140 & w6622;
assign w10247 = ~pi0601 & w4056;
assign w10248 = ~pi1103 & w6612;
assign w10249 = ~pi0613 & w3150;
assign w10250 = ~pi1084 & w6627;
assign w10251 = ~pi0516 & w2866;
assign w10252 = ~pi0488 & w3188;
assign w10253 = ~pi0439 & w3953;
assign w10254 = ~pi0390 & w2932;
assign w10255 = ~pi1120 & w6620;
assign w10256 = ~w10244 & ~w10245;
assign w10257 = ~w10246 & ~w10247;
assign w10258 = ~w10248 & ~w10249;
assign w10259 = ~w10250 & ~w10251;
assign w10260 = ~w10252 & ~w10253;
assign w10261 = ~w10254 & ~w10255;
assign w10262 = w10260 & w10261;
assign w10263 = w10258 & w10259;
assign w10264 = w10256 & w10257;
assign w10265 = w10263 & w10264;
assign w10266 = w10262 & w10265;
assign w10267 = pi1795 & w10215;
assign w10268 = ~pi1393 & w10217;
assign w10269 = ~w10267 & ~w10268;
assign w10270 = pi1790 & w9933;
assign w10271 = ~pi1394 & w9935;
assign w10272 = ~w10270 & ~w10271;
assign w10273 = pi1792 & w10215;
assign w10274 = ~pi1395 & w10217;
assign w10275 = ~w10273 & ~w10274;
assign w10276 = pi1802 & w10215;
assign w10277 = ~pi1396 & w10217;
assign w10278 = ~w10276 & ~w10277;
assign w10279 = pi1790 & w10215;
assign w10280 = ~pi1397 & w10217;
assign w10281 = ~w10279 & ~w10280;
assign w10282 = ~w8007 & ~w8047;
assign w10283 = (w10282 & w8045) | (w10282 & w12974) | (w8045 & w12974);
assign w10284 = ~w8007 & w8009;
assign w10285 = ~w8006 & ~w10284;
assign w10286 = ~w10283 & w10285;
assign w10287 = pi0674 & ~pi1160;
assign w10288 = ~pi0674 & pi1160;
assign w10289 = ~w10287 & ~w10288;
assign w10290 = w10286 & w10289;
assign w10291 = ~w10286 & ~w10289;
assign w10292 = ~w10290 & ~w10291;
assign w10293 = ~w8156 & ~w8196;
assign w10294 = ~w8195 & w10293;
assign w10295 = ~w8156 & w8158;
assign w10296 = ~w8155 & ~w10295;
assign w10297 = ~w10294 & w10296;
assign w10298 = pi0563 & ~pi1266;
assign w10299 = ~pi0563 & pi1266;
assign w10300 = ~w10298 & ~w10299;
assign w10301 = w10297 & w10300;
assign w10302 = ~w10297 & ~w10300;
assign w10303 = ~w10301 & ~w10302;
assign w10304 = pi1798 & w10185;
assign w10305 = ~pi1400 & w10187;
assign w10306 = ~w10304 & ~w10305;
assign w10307 = pi0619 & pi1747;
assign w10308 = w2867 & w10307;
assign w10309 = pi1791 & w9933;
assign w10310 = ~pi1402 & w9935;
assign w10311 = ~w10309 & ~w10310;
assign w10312 = pi1795 & w10185;
assign w10313 = ~pi1403 & w10187;
assign w10314 = ~w10312 & ~w10313;
assign w10315 = pi1798 & w10215;
assign w10316 = ~pi1404 & w10217;
assign w10317 = ~w10315 & ~w10316;
assign w10318 = pi1792 & w10185;
assign w10319 = ~pi1405 & w10187;
assign w10320 = ~w10318 & ~w10319;
assign w10321 = pi1800 & w10185;
assign w10322 = ~pi1406 & w10187;
assign w10323 = ~w10321 & ~w10322;
assign w10324 = pi1802 & w10185;
assign w10325 = ~pi1407 & w10187;
assign w10326 = ~w10324 & ~w10325;
assign w10327 = pi1792 & w9933;
assign w10328 = ~pi1408 & w9935;
assign w10329 = ~w10327 & ~w10328;
assign w10330 = pi1793 & w9933;
assign w10331 = ~pi1411 & w9935;
assign w10332 = ~w10330 & ~w10331;
assign w10333 = pi1795 & w9933;
assign w10334 = ~pi1412 & w9935;
assign w10335 = ~w10333 & ~w10334;
assign w10336 = pi1413 & ~w9139;
assign w10337 = w8525 & ~w10336;
assign w10338 = pi1796 & w8523;
assign w10339 = ~w10337 & ~w10338;
assign w10340 = ~pi0370 & w3188;
assign w10341 = ~pi0453 & w3953;
assign w10342 = ~pi0637 & w5442;
assign w10343 = ~pi0457 & w4186;
assign w10344 = ~pi1138 & w6627;
assign w10345 = ~pi0317 & w2866;
assign w10346 = ~pi1052 & w6612;
assign w10347 = ~pi0554 & w4056;
assign w10348 = ~pi1125 & w6620;
assign w10349 = ~pi0365 & w3150;
assign w10350 = ~pi1100 & w6622;
assign w10351 = ~pi0323 & w2932;
assign w10352 = ~w10340 & ~w10341;
assign w10353 = ~w10342 & ~w10343;
assign w10354 = ~w10344 & ~w10345;
assign w10355 = ~w10346 & ~w10347;
assign w10356 = ~w10348 & ~w10349;
assign w10357 = ~w10350 & ~w10351;
assign w10358 = w10356 & w10357;
assign w10359 = w10354 & w10355;
assign w10360 = w10352 & w10353;
assign w10361 = w10359 & w10360;
assign w10362 = w10358 & w10361;
assign w10363 = ~pi0320 & w2866;
assign w10364 = ~pi0368 & w3150;
assign w10365 = pi1111 & w6612;
assign w10366 = pi1122 & w6620;
assign w10367 = ~pi0326 & w2932;
assign w10368 = pi1131 & w6627;
assign w10369 = ~pi0556 & w4056;
assign w10370 = ~pi0639 & w5442;
assign w10371 = ~pi0373 & w3188;
assign w10372 = ~pi0532 & w4186;
assign w10373 = pi1143 & w6622;
assign w10374 = ~pi0455 & w3953;
assign w10375 = ~w10363 & ~w10364;
assign w10376 = ~w10365 & ~w10366;
assign w10377 = ~w10367 & ~w10368;
assign w10378 = ~w10369 & ~w10370;
assign w10379 = ~w10371 & ~w10372;
assign w10380 = ~w10373 & ~w10374;
assign w10381 = w10379 & w10380;
assign w10382 = w10377 & w10378;
assign w10383 = w10375 & w10376;
assign w10384 = w10382 & w10383;
assign w10385 = w10381 & w10384;
assign w10386 = ~pi1460 & ~pi1465;
assign w10387 = pi1478 & ~pi1479;
assign w10388 = w10386 & w10387;
assign w10389 = pi1460 & pi1465;
assign w10390 = ~pi1478 & pi1479;
assign w10391 = w10389 & w10390;
assign w10392 = ~w10388 & ~w10391;
assign w10393 = ~pi1463 & pi1464;
assign w10394 = ~pi1466 & ~pi1472;
assign w10395 = ~pi1476 & w10394;
assign w10396 = w10393 & w10395;
assign w10397 = ~w10392 & w10396;
assign w10398 = pi1479 & pi1502;
assign w10399 = pi1518 & ~pi1521;
assign w10400 = w10398 & w10399;
assign w10401 = ~pi1479 & ~pi1502;
assign w10402 = ~pi1518 & pi1521;
assign w10403 = w10401 & w10402;
assign w10404 = ~w10400 & ~w10403;
assign w10405 = ~pi1506 & pi1508;
assign w10406 = ~pi1516 & ~pi1517;
assign w10407 = ~pi1519 & w10406;
assign w10408 = w10405 & w10407;
assign w10409 = ~w10404 & w10408;
assign w10410 = w2868 & w6641;
assign w10411 = pi1419 & ~w10410;
assign w10412 = ~pi1776 & w10410;
assign w10413 = ~w10411 & ~w10412;
assign w10414 = ~w8111 & w8140;
assign w10415 = ~w8141 & ~w10414;
assign w10416 = pi1192 & pi1276;
assign w10417 = ~pi1194 & ~w10416;
assign w10418 = ~pi1195 & w10417;
assign w10419 = ~pi1196 & w10418;
assign w10420 = ~pi1264 & w10419;
assign w10421 = ~pi1197 & w10420;
assign w10422 = ~pi1198 & w10421;
assign w10423 = ~pi1199 & w10422;
assign w10424 = ~pi1249 & w10423;
assign w10425 = ~pi1201 & w10424;
assign w10426 = pi1036 & ~w10425;
assign w10427 = ~pi1036 & w10425;
assign w10428 = ~w10426 & ~w10427;
assign w10429 = pi1747 & ~w215;
assign w10430 = pi1423 & ~w10410;
assign w10431 = ~pi1775 & w10410;
assign w10432 = ~w10430 & ~w10431;
assign w10433 = ~pi1748 & w2867;
assign w10434 = w6637 & w10433;
assign w10435 = pi1425 & ~w10410;
assign w10436 = ~pi1774 & w10410;
assign w10437 = ~w10435 & ~w10436;
assign w10438 = pi1426 & ~w10410;
assign w10439 = ~pi1777 & w10410;
assign w10440 = ~w10438 & ~w10439;
assign w10441 = ~pi1428 & ~pi1707;
assign w10442 = ~w10410 & ~w10441;
assign w10443 = pi1747 & ~w10442;
assign w10444 = pi1747 & ~w1092;
assign w10445 = ~w8013 & w8041;
assign w10446 = ~w8042 & ~w10445;
assign w10447 = ~w8057 & w8086;
assign w10448 = ~w8087 & ~w10447;
assign w10449 = ~w8162 & ~w8190;
assign w10450 = ~w8191 & ~w10449;
assign w10451 = pi1077 & pi1241;
assign w10452 = ~pi1173 & ~w10451;
assign w10453 = ~pi1087 & w10452;
assign w10454 = ~pi1174 & w10453;
assign w10455 = ~pi1093 & w10454;
assign w10456 = ~pi1175 & w10455;
assign w10457 = ~pi1089 & w10456;
assign w10458 = ~pi1082 & ~pi1176;
assign w10459 = w10457 & w10458;
assign w10460 = ~pi1177 & w10459;
assign w10461 = ~pi1179 & ~w10460;
assign w10462 = pi1179 & w10460;
assign w10463 = ~w10461 & ~w10462;
assign w10464 = ~pi1176 & w10457;
assign w10465 = pi1082 & ~w10464;
assign w10466 = ~w10459 & ~w10465;
assign w10467 = pi1213 & pi1214;
assign w10468 = ~pi1215 & ~w10467;
assign w10469 = ~pi1216 & w10468;
assign w10470 = ~pi1066 & w10469;
assign w10471 = ~pi1217 & w10470;
assign w10472 = ~pi1218 & w10471;
assign w10473 = ~pi1219 & w10472;
assign w10474 = ~pi1056 & w10473;
assign w10475 = pi1057 & ~w10474;
assign w10476 = ~pi1056 & ~pi1057;
assign w10477 = w10473 & w10476;
assign w10478 = ~w10475 & ~w10477;
assign w10479 = w6618 & w10433;
assign w10480 = pi1177 & ~w10459;
assign w10481 = ~w10460 & ~w10480;
assign w10482 = w6629 & w10433;
assign w10483 = w6624 & w10433;
assign w10484 = pi1232 & ~w10477;
assign w10485 = ~pi1232 & w10477;
assign w10486 = ~w10484 & ~w10485;
assign w10487 = ~w8016 & w8039;
assign w10488 = ~w8040 & ~w10487;
assign w10489 = ~w8060 & ~w8084;
assign w10490 = ~w8085 & ~w10489;
assign w10491 = ~w8114 & ~w8138;
assign w10492 = ~w8139 & ~w10491;
assign w10493 = ~pi0452 & w3953;
assign w10494 = ~pi0454 & w4186;
assign w10495 = ~pi0366 & w3188;
assign w10496 = ~pi0363 & w3150;
assign w10497 = ~pi0315 & w2866;
assign w10498 = ~pi0553 & w4056;
assign w10499 = ~pi0318 & w2932;
assign w10500 = ~pi0635 & w5442;
assign w10501 = ~w10493 & ~w10494;
assign w10502 = ~w10495 & ~w10496;
assign w10503 = ~w10497 & ~w10498;
assign w10504 = ~w10499 & ~w10500;
assign w10505 = w10503 & w10504;
assign w10506 = w10501 & w10502;
assign w10507 = w10505 & w10506;
assign w10508 = ~w8188 & w8190;
assign w10509 = ~pi1218 & ~w10508;
assign w10510 = ~w8187 & w8189;
assign w10511 = ~w10509 & ~w10510;
assign w10512 = pi1283 & pi1331;
assign w10513 = ~pi1154 & ~pi1155;
assign w10514 = ~pi1156 & w10513;
assign w10515 = ~pi1157 & w10514;
assign w10516 = ~w10512 & w10515;
assign w10517 = ~pi1275 & w10516;
assign w10518 = ~pi1158 & w10517;
assign w10519 = ~pi1346 & w10518;
assign w10520 = ~pi1159 & w10519;
assign w10521 = ~pi1269 & w10520;
assign w10522 = pi1160 & ~w10521;
assign w10523 = ~pi1160 & ~pi1269;
assign w10524 = w10520 & w10523;
assign w10525 = ~w10522 & ~w10524;
assign w10526 = pi1266 & ~w10485;
assign w10527 = ~pi1232 & ~pi1266;
assign w10528 = w10477 & w10527;
assign w10529 = ~w10526 & ~w10528;
assign w10530 = ~w8063 & w8082;
assign w10531 = ~w8083 & ~w10530;
assign w10532 = ~w8019 & w8037;
assign w10533 = ~w8038 & ~w10532;
assign w10534 = ~w8117 & w8136;
assign w10535 = ~w8137 & ~w10534;
assign w10536 = ~w8165 & w8184;
assign w10537 = ~w8185 & ~w10536;
assign w10538 = pi1198 & ~w10421;
assign w10539 = ~w10422 & ~w10538;
assign w10540 = pi1199 & ~w10422;
assign w10541 = ~w10423 & ~w10540;
assign w10542 = pi1201 & ~w10424;
assign w10543 = ~w10425 & ~w10542;
assign w10544 = ~pi0183 & pi1050;
assign w10545 = pi1457 & ~w2173;
assign w10546 = ~w10544 & ~w10545;
assign w10547 = pi1458 & ~w2677;
assign w10548 = ~w372 & ~w10547;
assign w10549 = pi1747 & ~w10548;
assign w10550 = pi1465 & pi1466;
assign w10551 = pi1464 & w10550;
assign w10552 = pi1472 & w10551;
assign w10553 = ~pi1460 & ~w10552;
assign w10554 = pi1460 & w10552;
assign w10555 = pi1626 & ~w10553;
assign w10556 = ~w10554 & w10555;
assign w10557 = pi1089 & ~w10456;
assign w10558 = ~w10457 & ~w10557;
assign w10559 = pi1176 & ~w10457;
assign w10560 = ~w10464 & ~w10559;
assign w10561 = pi1478 & w10554;
assign w10562 = ~pi1463 & ~w10561;
assign w10563 = pi1463 & w10561;
assign w10564 = pi1626 & ~w10562;
assign w10565 = ~w10563 & w10564;
assign w10566 = ~pi1464 & ~w10550;
assign w10567 = pi1626 & ~w10551;
assign w10568 = ~w10566 & w10567;
assign w10569 = ~pi1465 & ~pi1466;
assign w10570 = pi1626 & ~w10550;
assign w10571 = ~w10569 & w10570;
assign w10572 = ~pi1466 & pi1626;
assign w10573 = pi1159 & ~w10519;
assign w10574 = ~w10520 & ~w10573;
assign w10575 = pi1249 & ~w10423;
assign w10576 = ~w10424 & ~w10575;
assign w10577 = pi1269 & ~w10520;
assign w10578 = ~w10521 & ~w10577;
assign w10579 = ~pi0756 & ~pi0757;
assign w10580 = ~pi0811 & ~pi0812;
assign w10581 = ~pi0813 & ~pi0814;
assign w10582 = ~pi0815 & ~pi0816;
assign w10583 = ~pi0817 & ~pi0820;
assign w10584 = ~pi0828 & ~pi0830;
assign w10585 = ~pi0831 & ~pi0832;
assign w10586 = ~pi0833 & ~pi0834;
assign w10587 = ~pi0870 & w10586;
assign w10588 = w10584 & w10585;
assign w10589 = w10582 & w10583;
assign w10590 = w10580 & w10581;
assign w10591 = w10579 & w10590;
assign w10592 = w10588 & w10589;
assign w10593 = w10587 & w10592;
assign w10594 = w10591 & w10593;
assign w10595 = pi0829 & ~w10594;
assign w10596 = ~pi0752 & ~pi0758;
assign w10597 = ~pi0835 & ~pi0836;
assign w10598 = ~pi0837 & ~pi0838;
assign w10599 = ~pi0839 & ~pi0840;
assign w10600 = ~pi0843 & ~pi0851;
assign w10601 = ~pi0854 & ~pi0855;
assign w10602 = ~pi0856 & ~pi0857;
assign w10603 = ~pi0858 & ~pi0879;
assign w10604 = ~pi0880 & w10603;
assign w10605 = w10601 & w10602;
assign w10606 = w10599 & w10600;
assign w10607 = w10597 & w10598;
assign w10608 = w10596 & w10607;
assign w10609 = w10605 & w10606;
assign w10610 = w10604 & w10609;
assign w10611 = w10608 & w10610;
assign w10612 = pi0853 & ~w10611;
assign w10613 = ~pi1472 & ~w10551;
assign w10614 = pi1626 & ~w10552;
assign w10615 = ~w10613 & w10614;
assign w10616 = w6609 & w10433;
assign w10617 = pi1175 & ~w10455;
assign w10618 = ~w10456 & ~w10617;
assign w10619 = pi1218 & ~w10471;
assign w10620 = ~w10472 & ~w10619;
assign w10621 = ~pi1476 & ~w10563;
assign w10622 = pi1476 & w10563;
assign w10623 = pi1626 & ~w10621;
assign w10624 = ~w10622 & w10623;
assign w10625 = ~pi1087 & ~pi1089;
assign w10626 = ~pi1093 & ~pi1173;
assign w10627 = ~pi1174 & ~pi1175;
assign w10628 = ~pi1177 & ~pi1179;
assign w10629 = w10627 & w10628;
assign w10630 = w10625 & w10626;
assign w10631 = w10458 & w10630;
assign w10632 = w10629 & w10631;
assign w10633 = w5922 & ~w10632;
assign w10634 = ~pi1478 & ~w10554;
assign w10635 = pi1626 & ~w10561;
assign w10636 = ~w10634 & w10635;
assign w10637 = ~pi0760 & ~pi1479;
assign w10638 = ~w2168 & ~w10637;
assign w10639 = ~pi0333 & ~pi1099;
assign w10640 = ~pi0221 & pi1099;
assign w10641 = ~w10639 & ~w10640;
assign w10642 = pi1195 & ~w10417;
assign w10643 = ~w10418 & ~w10642;
assign w10644 = pi1158 & ~w10517;
assign w10645 = ~w10518 & ~w10644;
assign w10646 = pi1219 & ~w10472;
assign w10647 = ~w10473 & ~w10646;
assign w10648 = pi1346 & ~w10518;
assign w10649 = ~w10519 & ~w10648;
assign w10650 = pi1056 & ~w10473;
assign w10651 = ~w10474 & ~w10650;
assign w10652 = ~pi1611 & ~pi1617;
assign w10653 = pi1196 & ~w10418;
assign w10654 = ~w10419 & ~w10653;
assign w10655 = pi1194 & w10416;
assign w10656 = ~w10417 & ~w10655;
assign w10657 = pi1197 & ~w10420;
assign w10658 = ~w10421 & ~w10657;
assign w10659 = ~pi1066 & ~pi1215;
assign w10660 = ~pi1216 & ~pi1217;
assign w10661 = ~pi1218 & ~pi1219;
assign w10662 = w10660 & w10661;
assign w10663 = w10476 & w10659;
assign w10664 = w10527 & w10663;
assign w10665 = w10662 & w10664;
assign w10666 = w6232 & ~w10665;
assign w10667 = ~pi1036 & ~pi1194;
assign w10668 = ~pi1195 & ~pi1196;
assign w10669 = ~pi1197 & ~pi1198;
assign w10670 = ~pi1199 & ~pi1201;
assign w10671 = ~pi1249 & ~pi1264;
assign w10672 = w10670 & w10671;
assign w10673 = w10668 & w10669;
assign w10674 = w10667 & w10673;
assign w10675 = w10672 & w10674;
assign w10676 = w6174 & ~w10675;
assign w10677 = ~pi1493 & ~w2677;
assign w10678 = pi1747 & ~w372;
assign w10679 = ~w10677 & w10678;
assign w10680 = pi1494 & ~w371;
assign w10681 = ~w1213 & ~w10680;
assign w10682 = pi1747 & ~w10681;
assign w10683 = pi1087 & ~w10452;
assign w10684 = ~w10453 & ~w10683;
assign w10685 = ~w8022 & ~w8035;
assign w10686 = ~w8036 & ~w10685;
assign w10687 = w8078 & ~w8080;
assign w10688 = ~w8081 & ~w10687;
assign w10689 = w8132 & ~w8134;
assign w10690 = ~w8135 & ~w10689;
assign w10691 = w8180 & ~w8182;
assign w10692 = ~w8183 & ~w10691;
assign w10693 = pi1517 & pi1518;
assign w10694 = pi1508 & w10693;
assign w10695 = pi1506 & w10694;
assign w10696 = ~pi1502 & ~w10695;
assign w10697 = pi1502 & w10695;
assign w10698 = ~pi1581 & ~w10696;
assign w10699 = ~w10697 & w10698;
assign w10700 = pi1613 & pi1616;
assign w10701 = pi1619 & pi1620;
assign w10702 = pi1612 & pi1618;
assign w10703 = ~pi1506 & ~w10694;
assign w10704 = ~pi1581 & ~w10695;
assign w10705 = ~w10703 & w10704;
assign w10706 = pi1174 & ~w10453;
assign w10707 = ~w10454 & ~w10706;
assign w10708 = ~pi1508 & ~w10693;
assign w10709 = ~pi1581 & ~w10694;
assign w10710 = ~w10708 & w10709;
assign w10711 = pi1173 & w10451;
assign w10712 = ~w10452 & ~w10711;
assign w10713 = pi1093 & ~w10454;
assign w10714 = ~w10455 & ~w10713;
assign w10715 = pi1264 & ~w10419;
assign w10716 = ~w10420 & ~w10715;
assign w10717 = pi1275 & ~w10516;
assign w10718 = ~w10517 & ~w10717;
assign w10719 = pi1217 & ~w10470;
assign w10720 = ~w10471 & ~w10719;
assign w10721 = pi1521 & w10697;
assign w10722 = ~pi1516 & ~w10721;
assign w10723 = pi1516 & w10721;
assign w10724 = ~pi1581 & ~w10722;
assign w10725 = ~w10723 & w10724;
assign w10726 = ~pi1517 & ~pi1581;
assign w10727 = ~pi1517 & ~pi1518;
assign w10728 = ~pi1581 & ~w10693;
assign w10729 = ~w10727 & w10728;
assign w10730 = ~pi1519 & ~w10723;
assign w10731 = pi1519 & w10723;
assign w10732 = ~pi1581 & ~w10730;
assign w10733 = ~w10731 & w10732;
assign w10734 = ~pi1158 & ~pi1159;
assign w10735 = ~pi1275 & ~pi1346;
assign w10736 = w10734 & w10735;
assign w10737 = w10523 & w10736;
assign w10738 = w10515 & w10737;
assign w10739 = w6339 & ~w10738;
assign w10740 = ~pi1521 & ~w10697;
assign w10741 = ~pi1581 & ~w10721;
assign w10742 = ~w10740 & w10741;
assign w10743 = pi0788 & w6408;
assign w10744 = pi0783 & w10743;
assign w10745 = ~pi0764 & w10744;
assign w10746 = ~pi0790 & w10745;
assign w10747 = pi0765 & w10746;
assign w10748 = ~pi0766 & ~w10747;
assign w10749 = pi0766 & w10747;
assign w10750 = ~w10748 & ~w10749;
assign w10751 = pi1227 & ~pi1230;
assign w10752 = ~pi1227 & pi1230;
assign w10753 = ~w10751 & ~w10752;
assign w10754 = ~pi1079 & ~pi1236;
assign w10755 = pi1079 & pi1236;
assign w10756 = ~pi1058 & ~pi1229;
assign w10757 = pi1058 & pi1229;
assign w10758 = pi1228 & ~pi1231;
assign w10759 = ~pi1228 & pi1231;
assign w10760 = ~w10758 & ~w10759;
assign w10761 = ~w10754 & ~w10755;
assign w10762 = ~w10756 & ~w10757;
assign w10763 = w10761 & w10762;
assign w10764 = ~w10753 & ~w10760;
assign w10765 = w10763 & w10764;
assign w10766 = ~pi1154 & ~w10512;
assign w10767 = pi1155 & ~w10766;
assign w10768 = ~w10512 & w10513;
assign w10769 = ~w10767 & ~w10768;
assign w10770 = pi1216 & ~w10468;
assign w10771 = ~w10469 & ~w10770;
assign w10772 = w398 & w7755;
assign w10773 = ~pi0765 & ~w10746;
assign w10774 = ~w10747 & ~w10773;
assign w10775 = w8031 & ~w8033;
assign w10776 = ~w8034 & ~w10775;
assign w10777 = ~w8067 & w8076;
assign w10778 = ~w8077 & ~w10777;
assign w10779 = ~w8121 & w8130;
assign w10780 = ~w8131 & ~w10779;
assign w10781 = ~w8169 & w8178;
assign w10782 = ~w8179 & ~w10781;
assign w10783 = pi0764 & ~w10744;
assign w10784 = ~w10745 & ~w10783;
assign w10785 = pi1156 & ~w10768;
assign w10786 = ~w10512 & w10514;
assign w10787 = ~w10785 & ~w10786;
assign w10788 = pi0283 & pi0290;
assign w10789 = ~pi0292 & ~pi0293;
assign w10790 = ~pi1534 & w10789;
assign w10791 = w10788 & w10790;
assign w10792 = w2710 & w10791;
assign w10793 = pi1066 & ~w10469;
assign w10794 = ~w10470 & ~w10793;
assign w10795 = pi1215 & w10467;
assign w10796 = ~w10468 & ~w10795;
assign w10797 = pi1157 & ~w10786;
assign w10798 = ~w10516 & ~w10797;
assign w10799 = w1586 & ~w5866;
assign w10800 = w1501 & ~w5927;
assign w10801 = w1405 & ~w6135;
assign w10802 = pi0761 & pi0765;
assign w10803 = ~pi0766 & pi0783;
assign w10804 = ~pi0787 & ~pi0788;
assign w10805 = w10803 & w10804;
assign w10806 = w6891 & w10802;
assign w10807 = w10805 & w10806;
assign w10808 = pi1154 & w10512;
assign w10809 = ~w10766 & ~w10808;
assign w10810 = pi0790 & ~w10745;
assign w10811 = ~w10746 & ~w10810;
assign w10812 = ~pi0783 & ~w10743;
assign w10813 = ~w10744 & ~w10812;
assign w10814 = pi1551 & pi1694;
assign w10815 = ~pi1840 & ~w10814;
assign w10816 = pi1747 & ~w10815;
assign w10817 = ~w8122 & ~w8123;
assign w10818 = w8128 & ~w10817;
assign w10819 = ~w8128 & w10817;
assign w10820 = ~w10818 & ~w10819;
assign w10821 = ~w8068 & ~w8069;
assign w10822 = w8074 & ~w10821;
assign w10823 = ~w8074 & w10821;
assign w10824 = ~w10822 & ~w10823;
assign w10825 = ~w8029 & w8031;
assign w10826 = ~pi1154 & ~w10825;
assign w10827 = ~w8028 & w8030;
assign w10828 = ~w10826 & ~w10827;
assign w10829 = ~w8170 & ~w8171;
assign w10830 = w8176 & ~w10829;
assign w10831 = ~w8176 & w10829;
assign w10832 = ~w10830 & ~w10831;
assign w10833 = pi1556 & pi1689;
assign w10834 = ~pi1839 & ~w10833;
assign w10835 = pi1747 & ~w10834;
assign w10836 = ~w8172 & ~w8173;
assign w10837 = w8174 & ~w10836;
assign w10838 = ~w8174 & w10836;
assign w10839 = ~w10837 & ~w10838;
assign w10840 = ~w8124 & ~w8125;
assign w10841 = w8126 & ~w10840;
assign w10842 = ~w8126 & w10840;
assign w10843 = ~w10841 & ~w10842;
assign w10844 = ~w8070 & ~w8071;
assign w10845 = w8072 & ~w10844;
assign w10846 = ~w8072 & w10844;
assign w10847 = ~w10845 & ~w10846;
assign w10848 = ~w8024 & ~w8025;
assign w10849 = w8026 & ~w10848;
assign w10850 = ~w8026 & w10848;
assign w10851 = ~w10849 & ~w10850;
assign w10852 = pi1561 & pi1691;
assign w10853 = ~pi1838 & ~w10852;
assign w10854 = pi1747 & ~w10853;
assign w10855 = pi1562 & pi1696;
assign w10856 = ~pi1841 & ~w10855;
assign w10857 = pi1747 & ~w10856;
assign w10858 = pi1563 & ~w817;
assign w10859 = pi1825 & w817;
assign w10860 = ~w10858 & ~w10859;
assign w10861 = pi1564 & ~w817;
assign w10862 = pi1807 & w817;
assign w10863 = ~w10861 & ~w10862;
assign w10864 = ~pi1077 & ~pi1241;
assign w10865 = ~w10451 & ~w10864;
assign w10866 = ~pi1283 & ~pi1331;
assign w10867 = ~w10512 & ~w10866;
assign w10868 = ~pi1213 & ~pi1214;
assign w10869 = ~w10467 & ~w10868;
assign w10870 = ~pi1697 & ~w2873;
assign w10871 = ~pi1690 & ~w2873;
assign w10872 = ~pi1679 & ~w2873;
assign w10873 = pi1573 & ~w817;
assign w10874 = pi1837 & w817;
assign w10875 = ~w10873 & ~w10874;
assign w10876 = pi1574 & ~w817;
assign w10877 = pi1836 & w817;
assign w10878 = ~w10876 & ~w10877;
assign w10879 = pi1575 & ~w817;
assign w10880 = pi1813 & w817;
assign w10881 = ~w10879 & ~w10880;
assign w10882 = pi1576 & ~w817;
assign w10883 = pi1830 & w817;
assign w10884 = ~w10882 & ~w10883;
assign w10885 = pi1577 & ~w817;
assign w10886 = pi1827 & w817;
assign w10887 = ~w10885 & ~w10886;
assign w10888 = ~pi0047 & ~w361;
assign w10889 = pi1583 & ~pi1743;
assign w10890 = pi0713 & ~w10889;
assign w10891 = pi1747 & ~w10890;
assign w10892 = pi1584 & ~w817;
assign w10893 = pi1832 & w817;
assign w10894 = ~w10892 & ~w10893;
assign w10895 = pi1585 & ~w817;
assign w10896 = pi1833 & w817;
assign w10897 = ~w10895 & ~w10896;
assign w10898 = pi1586 & ~w817;
assign w10899 = pi1809 & w817;
assign w10900 = ~w10898 & ~w10899;
assign w10901 = pi1587 & ~w817;
assign w10902 = pi1806 & w817;
assign w10903 = ~w10901 & ~w10902;
assign w10904 = pi1588 & ~w817;
assign w10905 = pi1818 & w817;
assign w10906 = ~w10904 & ~w10905;
assign w10907 = pi1589 & ~w817;
assign w10908 = pi1808 & w817;
assign w10909 = ~w10907 & ~w10908;
assign w10910 = pi1590 & ~w817;
assign w10911 = pi1814 & w817;
assign w10912 = ~w10910 & ~w10911;
assign w10913 = pi1591 & ~w817;
assign w10914 = pi1824 & w817;
assign w10915 = ~w10913 & ~w10914;
assign w10916 = pi1592 & ~w817;
assign w10917 = pi1834 & w817;
assign w10918 = ~w10916 & ~w10917;
assign w10919 = pi1593 & ~w817;
assign w10920 = pi1820 & w817;
assign w10921 = ~w10919 & ~w10920;
assign w10922 = ~pi1699 & ~w2873;
assign w10923 = pi1595 & ~w817;
assign w10924 = pi1812 & w817;
assign w10925 = ~w10923 & ~w10924;
assign w10926 = pi1596 & ~w817;
assign w10927 = pi1811 & w817;
assign w10928 = ~w10926 & ~w10927;
assign w10929 = pi1597 & ~w817;
assign w10930 = pi1815 & w817;
assign w10931 = ~w10929 & ~w10930;
assign w10932 = pi1598 & ~w817;
assign w10933 = pi1826 & w817;
assign w10934 = ~w10932 & ~w10933;
assign w10935 = pi1599 & ~w817;
assign w10936 = pi1828 & w817;
assign w10937 = ~w10935 & ~w10936;
assign w10938 = pi1600 & ~w817;
assign w10939 = pi1821 & w817;
assign w10940 = ~w10938 & ~w10939;
assign w10941 = pi1601 & ~w817;
assign w10942 = pi1829 & w817;
assign w10943 = ~w10941 & ~w10942;
assign w10944 = pi1602 & ~w817;
assign w10945 = pi1831 & w817;
assign w10946 = ~w10944 & ~w10945;
assign w10947 = pi1603 & ~w817;
assign w10948 = pi1823 & w817;
assign w10949 = ~w10947 & ~w10948;
assign w10950 = pi1604 & ~pi1728;
assign w10951 = pi0721 & ~w10950;
assign w10952 = pi1747 & ~w10951;
assign w10953 = pi1605 & ~w817;
assign w10954 = pi1822 & w817;
assign w10955 = ~w10953 & ~w10954;
assign w10956 = pi1606 & ~w817;
assign w10957 = pi1810 & w817;
assign w10958 = ~w10956 & ~w10957;
assign w10959 = pi1607 & ~pi1734;
assign w10960 = pi0676 & ~w10959;
assign w10961 = pi1747 & ~w10960;
assign w10962 = pi1608 & ~pi1730;
assign w10963 = pi0711 & ~w10962;
assign w10964 = pi1747 & ~w10963;
assign w10965 = pi1609 & ~w817;
assign w10966 = pi1835 & w817;
assign w10967 = ~w10965 & ~w10966;
assign w10968 = pi1610 & ~w817;
assign w10969 = pi1816 & w817;
assign w10970 = ~w10968 & ~w10969;
assign w10971 = pi0990 & ~pi1412;
assign w10972 = ~pi0891 & ~pi0959;
assign w10973 = ~pi1411 & ~w10972;
assign w10974 = pi0118 & ~pi1408;
assign w10975 = pi0131 & ~pi1391;
assign w10976 = pi0617 & ~pi1394;
assign w10977 = pi1037 & ~pi1402;
assign w10978 = ~w10971 & ~w10974;
assign w10979 = ~w10975 & ~w10976;
assign w10980 = ~w10977 & w10979;
assign w10981 = ~w10973 & w10978;
assign w10982 = w10980 & w10981;
assign w10983 = pi0114 & ~pi1405;
assign w10984 = ~pi0903 & ~pi0970;
assign w10985 = ~pi1380 & ~w10984;
assign w10986 = pi0592 & ~pi1377;
assign w10987 = pi1035 & ~pi1378;
assign w10988 = pi0128 & ~pi1379;
assign w10989 = pi1048 & ~pi1403;
assign w10990 = ~w10983 & ~w10986;
assign w10991 = ~w10987 & ~w10988;
assign w10992 = ~w10989 & w10991;
assign w10993 = ~w10985 & w10990;
assign w10994 = w10992 & w10993;
assign w10995 = pi0116 & ~pi1395;
assign w10996 = ~pi0904 & ~pi0958;
assign w10997 = ~pi1389 & ~w10996;
assign w10998 = pi0130 & ~pi1388;
assign w10999 = pi0991 & ~pi1387;
assign w11000 = pi0965 & ~pi1393;
assign w11001 = pi0615 & ~pi1397;
assign w11002 = ~w10995 & ~w10998;
assign w11003 = ~w10999 & ~w11000;
assign w11004 = ~w11001 & w11003;
assign w11005 = ~w10997 & w11002;
assign w11006 = w11004 & w11005;
assign w11007 = pi1614 & ~w817;
assign w11008 = pi1817 & w817;
assign w11009 = ~w11007 & ~w11008;
assign w11010 = pi1615 & ~w817;
assign w11011 = pi1819 & w817;
assign w11012 = ~w11010 & ~w11011;
assign w11013 = pi0116 & ~pi1384;
assign w11014 = ~pi1385 & ~w10996;
assign w11015 = pi0965 & ~pi1386;
assign w11016 = pi0991 & ~pi1383;
assign w11017 = pi0130 & ~pi1396;
assign w11018 = pi0615 & ~pi1404;
assign w11019 = ~w11013 & ~w11015;
assign w11020 = ~w11016 & ~w11017;
assign w11021 = ~w11018 & w11020;
assign w11022 = ~w11014 & w11019;
assign w11023 = w11021 & w11022;
assign w11024 = pi0118 & ~pi1390;
assign w11025 = ~pi1364 & ~w10972;
assign w11026 = pi0131 & ~pi1349;
assign w11027 = pi1037 & ~pi1362;
assign w11028 = pi0617 & ~pi1359;
assign w11029 = pi0990 & ~pi1352;
assign w11030 = ~w11024 & ~w11026;
assign w11031 = ~w11027 & ~w11028;
assign w11032 = ~w11029 & w11031;
assign w11033 = ~w11025 & w11030;
assign w11034 = w11032 & w11033;
assign w11035 = pi0128 & ~pi1407;
assign w11036 = ~pi1375 & ~w10984;
assign w11037 = pi0592 & ~pi1400;
assign w11038 = pi0114 & ~pi1406;
assign w11039 = pi1048 & ~pi1376;
assign w11040 = pi1035 & ~pi1374;
assign w11041 = ~w11035 & ~w11037;
assign w11042 = ~w11038 & ~w11039;
assign w11043 = ~w11040 & w11042;
assign w11044 = ~w11036 & w11041;
assign w11045 = w11043 & w11044;
assign w11046 = pi0115 & ~pi1382;
assign w11047 = ~pi0892 & ~pi0957;
assign w11048 = ~pi1348 & ~w11047;
assign w11049 = pi0535 & ~pi1381;
assign w11050 = pi1314 & ~pi1356;
assign w11051 = pi0129 & ~pi1353;
assign w11052 = pi1165 & ~pi1363;
assign w11053 = ~w11046 & ~w11049;
assign w11054 = ~w11050 & ~w11051;
assign w11055 = ~w11052 & w11054;
assign w11056 = ~w11048 & w11053;
assign w11057 = w11055 & w11056;
assign w11058 = pi0535 & ~pi1357;
assign w11059 = ~pi1354 & ~w11047;
assign w11060 = pi0115 & ~pi1350;
assign w11061 = pi1165 & ~pi1355;
assign w11062 = pi0129 & ~pi1351;
assign w11063 = pi1314 & ~pi1347;
assign w11064 = ~w11058 & ~w11060;
assign w11065 = ~w11061 & ~w11062;
assign w11066 = ~w11063 & w11065;
assign w11067 = ~w11059 & w11064;
assign w11068 = w11066 & w11067;
assign w11069 = ~pi0295 & ~pi0296;
assign w11070 = pi0297 & pi0298;
assign w11071 = pi0307 & ~pi0308;
assign w11072 = w11070 & w11071;
assign w11073 = w2719 & w11069;
assign w11074 = w11072 & w11073;
assign w11075 = ~pi0700 & pi1331;
assign w11076 = ~w8026 & ~w11075;
assign w11077 = ~pi0594 & pi1213;
assign w11078 = ~w8174 & ~w11077;
assign w11079 = ~pi0410 & pi1241;
assign w11080 = ~w8072 & ~w11079;
assign w11081 = pi1747 & pi1755;
assign w11082 = pi1747 & pi1756;
assign w11083 = pi1747 & pi1754;
assign w11084 = ~pi0511 & pi1192;
assign w11085 = ~w8126 & ~w11084;
assign w11086 = ~w6409 & ~w10743;
assign w11087 = ~pi0038 & pi1101;
assign w11088 = pi1632 & ~w11087;
assign w11089 = pi1808 & w11087;
assign w11090 = ~w11088 & ~w11089;
assign w11091 = pi1633 & ~w11087;
assign w11092 = pi1837 & w11087;
assign w11093 = ~w11091 & ~w11092;
assign w11094 = pi1634 & ~w11087;
assign w11095 = pi1834 & w11087;
assign w11096 = ~w11094 & ~w11095;
assign w11097 = pi1635 & ~w11087;
assign w11098 = pi1812 & w11087;
assign w11099 = ~w11097 & ~w11098;
assign w11100 = pi1636 & ~w11087;
assign w11101 = pi1829 & w11087;
assign w11102 = ~w11100 & ~w11101;
assign w11103 = ~pi1192 & ~pi1276;
assign w11104 = ~w10416 & ~w11103;
assign w11105 = pi1638 & ~w11087;
assign w11106 = pi1825 & w11087;
assign w11107 = ~w11105 & ~w11106;
assign w11108 = pi1639 & ~w11087;
assign w11109 = pi1830 & w11087;
assign w11110 = ~w11108 & ~w11109;
assign w11111 = pi1640 & ~w11087;
assign w11112 = pi1824 & w11087;
assign w11113 = ~w11111 & ~w11112;
assign w11114 = pi1641 & ~w11087;
assign w11115 = pi1816 & w11087;
assign w11116 = ~w11114 & ~w11115;
assign w11117 = pi1642 & ~w11087;
assign w11118 = pi1810 & w11087;
assign w11119 = ~w11117 & ~w11118;
assign w11120 = pi1643 & ~w11087;
assign w11121 = pi1836 & w11087;
assign w11122 = ~w11120 & ~w11121;
assign w11123 = pi1644 & ~w11087;
assign w11124 = pi1833 & w11087;
assign w11125 = ~w11123 & ~w11124;
assign w11126 = pi1645 & ~w11087;
assign w11127 = pi1809 & w11087;
assign w11128 = ~w11126 & ~w11127;
assign w11129 = pi1646 & ~w11087;
assign w11130 = pi1811 & w11087;
assign w11131 = ~w11129 & ~w11130;
assign w11132 = pi1647 & ~w11087;
assign w11133 = pi1814 & w11087;
assign w11134 = ~w11132 & ~w11133;
assign w11135 = pi1648 & ~w11087;
assign w11136 = pi1832 & w11087;
assign w11137 = ~w11135 & ~w11136;
assign w11138 = pi1649 & ~w11087;
assign w11139 = pi1820 & w11087;
assign w11140 = ~w11138 & ~w11139;
assign w11141 = pi1650 & ~w11087;
assign w11142 = pi1806 & w11087;
assign w11143 = ~w11141 & ~w11142;
assign w11144 = pi1651 & ~w11087;
assign w11145 = pi1807 & w11087;
assign w11146 = ~w11144 & ~w11145;
assign w11147 = pi1652 & ~w11087;
assign w11148 = pi1835 & w11087;
assign w11149 = ~w11147 & ~w11148;
assign w11150 = pi1653 & ~w11087;
assign w11151 = pi1815 & w11087;
assign w11152 = ~w11150 & ~w11151;
assign w11153 = pi1654 & ~w11087;
assign w11154 = pi1827 & w11087;
assign w11155 = ~w11153 & ~w11154;
assign w11156 = pi1655 & ~w11087;
assign w11157 = pi1826 & w11087;
assign w11158 = ~w11156 & ~w11157;
assign w11159 = pi1656 & ~w11087;
assign w11160 = pi1822 & w11087;
assign w11161 = ~w11159 & ~w11160;
assign w11162 = pi1657 & ~w11087;
assign w11163 = pi1823 & w11087;
assign w11164 = ~w11162 & ~w11163;
assign w11165 = pi1658 & ~w11087;
assign w11166 = pi1813 & w11087;
assign w11167 = ~w11165 & ~w11166;
assign w11168 = pi1659 & ~w11087;
assign w11169 = pi1828 & w11087;
assign w11170 = ~w11168 & ~w11169;
assign w11171 = pi1660 & ~w11087;
assign w11172 = pi1819 & w11087;
assign w11173 = ~w11171 & ~w11172;
assign w11174 = pi1661 & ~w11087;
assign w11175 = pi1831 & w11087;
assign w11176 = ~w11174 & ~w11175;
assign w11177 = pi1662 & ~w11087;
assign w11178 = pi1818 & w11087;
assign w11179 = ~w11177 & ~w11178;
assign w11180 = pi1663 & ~w11087;
assign w11181 = pi1821 & w11087;
assign w11182 = ~w11180 & ~w11181;
assign w11183 = pi1664 & ~w11087;
assign w11184 = pi1817 & w11087;
assign w11185 = ~w11183 & ~w11184;
assign w11186 = ~pi0763 & ~pi0791;
assign w11187 = pi0792 & ~pi0793;
assign w11188 = w11186 & w11187;
assign w11189 = pi0012 & ~pi1099;
assign w11190 = ~pi0919 & ~pi0921;
assign w11191 = pi0963 & w11190;
assign w11192 = pi0274 & pi0275;
assign w11193 = pi0285 & w11192;
assign w11194 = w2680 & w11193;
assign w11195 = ~pi0200 & ~pi1099;
assign w11196 = ~w6408 & ~w6892;
assign w11197 = pi1749 & pi1750;
assign w11198 = w2 & ~pi1370;
assign w11199 = ~pi0309 & w1;
assign w11200 = w11 & ~w2;
assign w11201 = ~pi0677 & ~pi1401;
assign w11202 = w19 & w23;
assign w11203 = ~w33 & ~w137;
assign w11204 = ~pi0093 & pi0068;
assign w11205 = pi1753 & ~w189;
assign w11206 = ~pi0005 & pi0004;
assign w11207 = ~pi1753 & pi1667;
assign w11208 = w11207 & pi0000;
assign w11209 = pi0005 & ~pi0004;
assign w11210 = pi1753 & w189;
assign w11211 = w198 & pi1692;
assign w11212 = w198 & ~pi1692;
assign w11213 = ~w214 & ~w211;
assign w11214 = w216 & ~w185;
assign w11215 = w205 & ~w217;
assign w11216 = ~w219 & ~pi0199;
assign w11217 = ~pi0055 & ~pi0874;
assign w11218 = ~w228 & pi1586;
assign w11219 = ~w223 & pi1563;
assign w11220 = ~pi0193 & pi1638;
assign w11221 = ~w228 & pi1645;
assign w11222 = ~w228 & pi1614;
assign w11223 = ~w223 & pi1585;
assign w11224 = ~pi0193 & pi1644;
assign w11225 = ~w228 & pi1664;
assign w11226 = ~w203 & ~w257;
assign w11227 = w205 & ~w260;
assign w11228 = pi0779 & ~w259;
assign w11229 = ~w218 & w264;
assign w11230 = ~pi0005 & ~pi0004;
assign w11231 = ~w223 & pi1601;
assign w11232 = ~w228 & pi1658;
assign w11233 = ~pi0193 & pi1636;
assign w11234 = ~w228 & pi1575;
assign w11235 = ~w223 & pi1573;
assign w11236 = ~w228 & pi1663;
assign w11237 = ~pi0193 & pi1633;
assign w11238 = ~w228 & pi1600;
assign w11239 = pi0025 & ~w287;
assign w11240 = ~w218 & ~w289;
assign w11241 = w11207 & pi0001;
assign w11242 = pi0005 & pi0004;
assign w11243 = w11207 & pi0002;
assign w11244 = ~w223 & pi1591;
assign w11245 = ~w228 & pi1589;
assign w11246 = ~pi0193 & pi1640;
assign w11247 = ~w228 & pi1632;
assign w11248 = ~w223 & pi1584;
assign w11249 = ~w228 & pi1610;
assign w11250 = ~pi0193 & pi1648;
assign w11251 = ~w228 & pi1641;
assign w11252 = w205 & ~w315;
assign w11253 = pi0778 & ~w317;
assign w11254 = ~w218 & w320;
assign w11255 = w11207 & pi0003;
assign w11256 = ~w228 & pi1593;
assign w11257 = ~w223 & pi1574;
assign w11258 = ~pi0193 & pi1643;
assign w11259 = ~w228 & pi1649;
assign w11260 = ~w228 & pi1595;
assign w11261 = ~w223 & pi1599;
assign w11262 = ~pi0193 & pi1659;
assign w11263 = ~w228 & pi1635;
assign w11264 = ~pi0054 & ~w342;
assign w11265 = ~w218 & ~w344;
assign w11266 = ~w350 & w349;
assign w11267 = pi0352 & ~w359;
assign w11268 = ~pi0110 & ~pi0111;
assign w11269 = ~pi0095 & w361;
assign w11270 = ~pi0109 & ~pi0089;
assign w11271 = ~pi1229 & pi1236;
assign w11272 = ~pi0796 & ~pi1470;
assign w11273 = ~w369 & w368;
assign w11274 = w360 & w369;
assign w11275 = ~pi0796 & pi0024;
assign w11276 = w396 & w399;
assign w11277 = ~w396 & ~pi0776;
assign w11278 = pi0796 & pi0750;
assign w11279 = ~pi0771 & pi0148;
assign w11280 = ~w411 & pi0946;
assign w11281 = w411 & ~pi0946;
assign w11282 = pi0796 & pi0859;
assign w11283 = ~pi0771 & pi0187;
assign w11284 = ~w417 & ~pi0895;
assign w11285 = w412 & pi0940;
assign w11286 = pi0796 & pi0804;
assign w11287 = ~pi0238 & ~w424;
assign w11288 = pi0796 & pi0807;
assign w11289 = ~pi0240 & ~w429;
assign w11290 = w431 & pi0742;
assign w11291 = pi0796 & pi0806;
assign w11292 = ~pi0239 & ~w433;
assign w11293 = ~w435 & ~pi0741;
assign w11294 = w435 & pi0741;
assign w11295 = ~w421 & w439;
assign w11296 = ~w431 & ~pi0742;
assign w11297 = ~w443 & ~pi0945;
assign w11298 = pi0796 & pi0755;
assign w11299 = ~pi0221 & ~w445;
assign w11300 = ~w448 & pi0945;
assign w11301 = ~w448 & ~w11297;
assign w11302 = pi0796 & pi0808;
assign w11303 = ~pi0241 & ~w450;
assign w11304 = ~w452 & ~pi0867;
assign w11305 = w452 & pi0867;
assign w11306 = w443 & pi0945;
assign w11307 = pi0796 & pi0877;
assign w11308 = ~pi0236 & ~w458;
assign w11309 = ~w460 & ~pi0739;
assign w11310 = ~pi0771 & pi0190;
assign w11311 = pi0796 & pi0810;
assign w11312 = ~pi0224 & ~w465;
assign w11313 = ~w467 & ~pi0869;
assign w11314 = pi0796 & pi0809;
assign w11315 = ~pi0242 & ~w469;
assign w11316 = w471 & pi0868;
assign w11317 = ~w471 & ~pi0868;
assign w11318 = pi0796 & pi0759;
assign w11319 = ~pi0243 & ~w476;
assign w11320 = w478 & pi0875;
assign w11321 = ~w478 & ~pi0875;
assign w11322 = w449 & w484;
assign w11323 = w467 & pi0869;
assign w11324 = w481 & w464;
assign w11325 = w460 & pi0739;
assign w11326 = ~w490 & w495;
assign w11327 = ~pi0771 & pi0191;
assign w11328 = ~pi0774 & ~w498;
assign w11329 = ~w11326 & w499;
assign w11330 = ~pi0771 & pi0192;
assign w11331 = ~w500 & ~pi1099;
assign w11332 = ~w506 & ~w499;
assign w11333 = ~w506 & ~w11329;
assign w11334 = w11326 & w508;
assign w11335 = ~pi0774 & ~pi1099;
assign w11336 = ~w11334 & w510;
assign w11337 = ~w396 & pi0024;
assign w11338 = w396 & pi0672;
assign w11339 = ~w228 & pi1588;
assign w11340 = ~w223 & pi1592;
assign w11341 = ~pi0193 & pi1634;
assign w11342 = ~w228 & pi1662;
assign w11343 = ~w228 & pi1606;
assign w11344 = ~w223 & pi1598;
assign w11345 = ~pi0193 & pi1655;
assign w11346 = ~w228 & pi1642;
assign w11347 = ~w228 & pi1650;
assign w11348 = ~w223 & pi1605;
assign w11349 = ~w228 & pi1587;
assign w11350 = ~pi0193 & pi1656;
assign w11351 = ~w228 & pi1647;
assign w11352 = ~w223 & pi1576;
assign w11353 = ~w228 & pi1590;
assign w11354 = ~pi0193 & pi1639;
assign w11355 = ~w228 & pi1653;
assign w11356 = ~w223 & pi1602;
assign w11357 = ~w228 & pi1597;
assign w11358 = ~pi0193 & pi1661;
assign w11359 = ~w228 & pi1651;
assign w11360 = ~w223 & pi1603;
assign w11361 = ~w228 & pi1564;
assign w11362 = ~pi0193 & pi1657;
assign w11363 = ~w228 & pi1615;
assign w11364 = ~w223 & pi1609;
assign w11365 = ~pi0193 & pi1652;
assign w11366 = ~w228 & pi1660;
assign w11367 = ~w228 & pi1596;
assign w11368 = ~pi0193 & pi1654;
assign w11369 = ~pi1577 & ~w238;
assign w11370 = (~pi1646 & ~w228) | (~pi1646 & w12975) | (~w228 & w12975);
assign w11371 = ~w224 & ~w623;
assign w11372 = ~w624 & w631;
assign w11373 = pi0009 & ~w623;
assign w11374 = pi0009 & w11371;
assign w11375 = ~w634 & ~w11373;
assign w11376 = ~w634 & ~w11374;
assign w11377 = ~pi0010 & ~w623;
assign w11378 = ~pi0010 & w11371;
assign w11379 = ~w634 & ~w11377;
assign w11380 = ~w634 & ~w11378;
assign w11381 = w500 & ~w503;
assign w11382 = ~w490 & w641;
assign w11383 = ~w11382 & w644;
assign w11384 = w646 & ~w644;
assign w11385 = w646 & ~w11383;
assign w11386 = ~w490 & w648;
assign w11387 = ~pi0865 & ~pi1099;
assign w11388 = ~w645 & pi1099;
assign w11389 = ~w645 & ~w11387;
assign w11390 = pi0771 & pi0024;
assign w11391 = ~pi0771 & pi0029;
assign w11392 = ~w624 & w628;
assign w11393 = ~pi0013 & ~w623;
assign w11394 = ~pi0013 & w11371;
assign w11395 = ~w634 & ~w11393;
assign w11396 = ~w634 & ~w11394;
assign w11397 = ~w11326 & w663;
assign w11398 = w11326 & w665;
assign w11399 = pi0865 & pi0866;
assign w11400 = ~w11399 & ~pi1099;
assign w11401 = ~w669 & ~w672;
assign w11402 = w669 & pi0775;
assign w11403 = w449 & w483;
assign w11404 = ~w489 & ~w479;
assign w11405 = w11404 & w680;
assign w11406 = ~w11404 & w682;
assign w11407 = w11207 & pi0017;
assign w11408 = ~w218 & w689;
assign w11409 = ~w669 & ~w694;
assign w11410 = ~w650 & w696;
assign w11411 = ~w489 & w493;
assign w11412 = ~w11411 & ~w461;
assign w11413 = pi1099 & ~w701;
assign w11414 = w11207 & pi0020;
assign w11415 = pi0048 & ~w188;
assign w11416 = ~w218 & w710;
assign w11417 = w11207 & pi0021;
assign w11418 = ~pi0053 & w196;
assign w11419 = ~w218 & w717;
assign w11420 = w449 & w475;
assign w11421 = w468 & w722;
assign w11422 = w449 & ~pi1099;
assign w11423 = ~w756 & w757;
assign w11424 = ~w759 & w760;
assign w11425 = w761 & ~w760;
assign w11426 = w761 & ~w11424;
assign w11427 = ~w763 & w764;
assign w11428 = w765 & ~w764;
assign w11429 = w765 & ~w11427;
assign w11430 = ~pi0025 & ~w623;
assign w11431 = ~pi0025 & w11371;
assign w11432 = ~w634 & ~w11430;
assign w11433 = ~w634 & ~w11431;
assign w11434 = w11207 & pi0026;
assign w11435 = ~w218 & w781;
assign w11436 = ~w472 & w785;
assign w11437 = w472 & ~w785;
assign w11438 = w449 & ~w453;
assign w11439 = w721 & ~pi1099;
assign w11440 = pi1579 & pi0044;
assign w11441 = pi0040 & pi0039;
assign w11442 = w11441 & pi0041;
assign w11443 = pi0034 & pi0035;
assign w11444 = w11443 & pi0036;
assign w11445 = w11444 & pi0037;
assign w11446 = pi0045 & pi0042;
assign w11447 = w11446 & pi0031;
assign w11448 = ~w11446 & ~pi0031;
assign w11449 = ~pi1579 & ~pi0044;
assign w11450 = ~pi0040 & ~pi0039;
assign w11451 = ~w11441 & ~pi0041;
assign w11452 = ~pi0034 & ~pi0035;
assign w11453 = ~w11443 & ~pi0036;
assign w11454 = ~w11444 & ~pi0037;
assign w11455 = ~pi0045 & ~pi0042;
assign w11456 = ~w11447 & w893;
assign w11457 = w11447 & ~w893;
assign w11458 = w11446 & w897;
assign w11459 = w11458 & pi0032;
assign w11460 = w11459 & ~w901;
assign w11461 = ~w11459 & w901;
assign w11462 = ~w11458 & ~pi0032;
assign w11463 = ~w847 & ~w852;
assign w11464 = ~w857 & ~w862;
assign w11465 = ~w867 & ~w872;
assign w11466 = ~w877 & ~w882;
assign w11467 = ~w887 & ~w896;
assign w11468 = w11467 & w916;
assign w11469 = w909 & w918;
assign w11470 = w909 & w922;
assign w11471 = w11459 & pi0033;
assign w11472 = ~w11459 & ~pi0033;
assign w11473 = w909 & w929;
assign w11474 = w909 & w933;
assign w11475 = w909 & w937;
assign w11476 = w909 & w941;
assign w11477 = w909 & w945;
assign w11478 = w909 & w949;
assign w11479 = w909 & w953;
assign w11480 = w909 & w957;
assign w11481 = w909 & w961;
assign w11482 = w909 & w965;
assign w11483 = ~w11447 & ~pi0043;
assign w11484 = ~w11458 & w815;
assign w11485 = w909 & w971;
assign w11486 = w909 & w975;
assign w11487 = w909 & w979;
assign w11488 = ~w421 & w438;
assign w11489 = w436 & w982;
assign w11490 = ~w436 & ~w982;
assign w11491 = ~w214 & ~w217;
assign w11492 = ~pi0048 & ~w623;
assign w11493 = ~pi0048 & w11371;
assign w11494 = ~w634 & ~w11492;
assign w11495 = ~w634 & ~w11493;
assign w11496 = pi0796 & pi0012;
assign w11497 = ~pi0095 & pi1099;
assign w11498 = pi0756 & pi1099;
assign w11499 = pi0756 & w11497;
assign w11500 = ~pi0983 & ~pi1099;
assign w11501 = ~pi0983 & w1060;
assign w11502 = w421 & ~w438;
assign w11503 = ~pi0050 & ~w623;
assign w11504 = ~pi0050 & w11371;
assign w11505 = ~w634 & ~w11503;
assign w11506 = ~w634 & ~w11504;
assign w11507 = ~pi0051 & ~w623;
assign w11508 = ~pi0051 & w11371;
assign w11509 = ~w634 & ~w11507;
assign w11510 = ~w634 & ~w11508;
assign w11511 = ~pi0052 & ~w623;
assign w11512 = ~pi0052 & w11371;
assign w11513 = ~w634 & ~w11511;
assign w11514 = ~w634 & ~w11512;
assign w11515 = pi0053 & ~w623;
assign w11516 = pi0053 & w11371;
assign w11517 = ~w634 & ~w11515;
assign w11518 = ~w634 & ~w11516;
assign w11519 = pi0054 & ~w623;
assign w11520 = pi0054 & w11371;
assign w11521 = ~w634 & ~w11519;
assign w11522 = ~w634 & ~w11520;
assign w11523 = ~pi0828 & pi1099;
assign w11524 = ~pi0828 & w11497;
assign w11525 = pi0894 & ~pi1099;
assign w11526 = pi0894 & w1060;
assign w11527 = w421 & w1007;
assign w11528 = ~pi0820 & pi1099;
assign w11529 = ~pi0820 & w11497;
assign w11530 = w216 & w185;
assign w11531 = ~pi0060 & ~w623;
assign w11532 = ~pi0060 & w11371;
assign w11533 = ~w634 & ~w11531;
assign w11534 = ~w634 & ~w11532;
assign w11535 = ~pi0811 & pi1099;
assign w11536 = ~pi0811 & w11497;
assign w11537 = pi1625 & pi0094;
assign w11538 = ~pi1625 & ~pi0066;
assign w11539 = w1098 & pi0138;
assign w11540 = pi1049 & ~w1162;
assign w11541 = w1172 & pi1233;
assign w11542 = ~w1204 & pi1747;
assign w11543 = w11270 & pi0067;
assign w11544 = ~pi1479 & ~w369;
assign w11545 = ~w370 & ~w374;
assign w11546 = w381 & ~pi0801;
assign w11547 = w1210 & w1216;
assign w11548 = ~w360 & w1207;
assign w11549 = ~pi0109 & w1219;
assign w11550 = w1223 & w1225;
assign w11551 = ~w1232 & ~pi0138;
assign w11552 = pi0625 & ~pi0111;
assign w11553 = w1251 & w1252;
assign w11554 = w1210 & w368;
assign w11555 = w1211 & ~pi0121;
assign w11556 = pi1747 & pi0121;
assign w11557 = pi1747 & ~w11555;
assign w11558 = w396 & pi0762;
assign w11559 = ~w396 & pi0749;
assign w11560 = w396 & pi0768;
assign w11561 = ~w396 & pi0852;
assign w11562 = w396 & pi0827;
assign w11563 = ~w396 & pi0850;
assign w11564 = w396 & pi0826;
assign w11565 = ~w396 & pi0849;
assign w11566 = w1276 & w1281;
assign w11567 = pi1747 & ~pi0121;
assign w11568 = pi1747 & w11555;
assign w11569 = pi0075 & w224;
assign w11570 = ~w1290 & ~w224;
assign w11571 = ~w1290 & ~w11569;
assign w11572 = ~pi0073 & w1289;
assign w11573 = w11572 & ~pi0080;
assign w11574 = ~w1294 & pi0069;
assign w11575 = w1294 & ~pi0069;
assign w11576 = ~w1305 & ~w1306;
assign w11577 = w11575 & ~pi0074;
assign w11578 = ~w11577 & pi0070;
assign w11579 = ~pi0073 & w1297;
assign w11580 = pi1458 & pi0751;
assign w11581 = ~pi1458 & pi0770;
assign w11582 = w396 & pi0825;
assign w11583 = ~w396 & pi0848;
assign w11584 = w370 & w12985;
assign w11585 = (pi0748 & ~w370) | (pi0748 & w12986) | (~w370 & w12986);
assign w11586 = ~pi1458 & pi0871;
assign w11587 = pi1458 & pi0754;
assign w11588 = ~pi1458 & pi0818;
assign w11589 = pi1458 & pi0841;
assign w11590 = pi1458 & pi0842;
assign w11591 = ~pi1458 & pi0819;
assign w11592 = w396 & pi0821;
assign w11593 = ~w396 & pi0844;
assign w11594 = ~w1362 & w1365;
assign w11595 = w370 & w12987;
assign w11596 = (pi0845 & ~w370) | (pi0845 & w12988) | (~w370 & w12988);
assign w11597 = w370 & w12989;
assign w11598 = (pi0846 & ~w370) | (pi0846 & w12990) | (~w370 & w12990);
assign w11599 = ~w1372 & w1378;
assign w11600 = w370 & w12991;
assign w11601 = (pi0847 & ~w370) | (pi0847 & w12992) | (~w370 & w12992);
assign w11602 = w1384 & ~w1378;
assign w11603 = w1384 & ~w11599;
assign w11604 = ~w1388 & w1390;
assign w11605 = w1329 & ~w1320;
assign w11606 = ~w1329 & pi0807;
assign w11607 = ~pi0073 & ~pi0076;
assign w11608 = w11607 & ~pi0077;
assign w11609 = w11608 & ~pi0078;
assign w11610 = ~w11609 & pi0071;
assign w11611 = w11609 & ~pi0071;
assign w11612 = ~w1399 & w11567;
assign w11613 = ~w1399 & w11568;
assign w11614 = ~pi1541 & pi1839;
assign w11615 = ~pi0072 & ~w1404;
assign w11616 = w1329 & ~w1345;
assign w11617 = ~w1329 & pi0859;
assign w11618 = ~pi0055 & pi0073;
assign w11619 = pi0073 & ~w1417;
assign w11620 = w1418 & w11567;
assign w11621 = w1418 & w11568;
assign w11622 = ~w11575 & pi0074;
assign w11623 = w1329 & ~w1339;
assign w11624 = ~w1329 & pi0750;
assign w11625 = pi0073 & pi0076;
assign w11626 = w1329 & ~w1353;
assign w11627 = ~w1329 & pi0804;
assign w11628 = ~w11607 & pi0077;
assign w11629 = w1329 & ~w1359;
assign w11630 = ~w1329 & pi0806;
assign w11631 = ~w11608 & pi0078;
assign w11632 = w1329 & ~w1370;
assign w11633 = ~w1329 & pi0755;
assign w11634 = ~w11611 & pi0079;
assign w11635 = ~w1300 & w11567;
assign w11636 = ~w1300 & w11568;
assign w11637 = w1329 & ~w1376;
assign w11638 = ~w1329 & pi0808;
assign w11639 = ~w11572 & pi0080;
assign w11640 = w1329 & ~w1382;
assign w11641 = ~w1329 & pi0809;
assign w11642 = w1329 & ~w1332;
assign w11643 = ~w1329 & pi0810;
assign w11644 = pi0081 & pi0082;
assign w11645 = ~w1303 & ~w1482;
assign w11646 = w1321 & pi0759;
assign w11647 = ~w1328 & ~w1326;
assign w11648 = ~w1485 & w1267;
assign w11649 = ~w1293 & pi0083;
assign w11650 = ~w1304 & ~w1489;
assign w11651 = ~pi1538 & pi1840;
assign w11652 = ~pi0084 & ~w1492;
assign w11653 = ~pi1540 & pi1838;
assign w11654 = ~pi0085 & ~w1500;
assign w11655 = pi0103 & pi0104;
assign w11656 = ~pi0103 & ~pi0104;
assign w11657 = ~w1513 & ~w1511;
assign w11658 = pi0105 & pi0106;
assign w11659 = w1519 & w1510;
assign w11660 = ~pi0105 & ~pi0106;
assign w11661 = ~w1522 & w1524;
assign w11662 = ~w1521 & ~w1508;
assign w11663 = w1537 & ~w1541;
assign w11664 = w1545 & w1547;
assign w11665 = ~w1542 & w1549;
assign w11666 = w1537 & w1553;
assign w11667 = ~w1554 & ~w1552;
assign w11668 = pi0100 & pi0101;
assign w11669 = w1537 & w1558;
assign w11670 = ~w1559 & ~w1560;
assign w11671 = ~w1565 & ~w1569;
assign w11672 = w1572 & w1581;
assign w11673 = ~w1572 & ~w1581;
assign w11674 = ~pi1539 & pi1841;
assign w11675 = ~pi0087 & ~w1585;
assign w11676 = pi0067 & pi1747;
assign w11677 = pi0067 & w11542;
assign w11678 = ~w1210 & w368;
assign w11679 = w1596 & w11676;
assign w11680 = w1596 & w11677;
assign w11681 = w11549 & w1598;
assign w11682 = w1599 & pi1747;
assign w11683 = w1599 & w11542;
assign w11684 = ~w1232 & w11682;
assign w11685 = ~w1232 & w11683;
assign w11686 = ~pi0999 & ~pi1005;
assign w11687 = pi0999 & pi1005;
assign w11688 = ~pi1011 & pi1012;
assign w11689 = ~w1638 & ~w1634;
assign w11690 = w11689 & ~w1633;
assign w11691 = ~w1631 & w1641;
assign w11692 = w1644 & ~w1632;
assign w11693 = w1647 & ~w1641;
assign w11694 = w1647 & ~w11691;
assign w11695 = pi1012 & ~w1281;
assign w11696 = ~w1644 & ~w1281;
assign w11697 = ~w1653 & ~w1652;
assign w11698 = w1648 & ~pi1013;
assign w11699 = ~pi1000 & pi1001;
assign w11700 = ~w1648 & ~w1657;
assign w11701 = pi1000 & ~pi1001;
assign w11702 = w1648 & ~w1665;
assign w11703 = w1265 & w11676;
assign w11704 = w1265 & w11677;
assign w11705 = w1224 & pi1747;
assign w11706 = w1224 & w11542;
assign w11707 = w1690 & w11705;
assign w11708 = w1690 & w11706;
assign w11709 = w361 & w362;
assign w11710 = ~w1224 & ~w1716;
assign w11711 = w1485 & w406;
assign w11712 = ~w1631 & w1639;
assign w11713 = w1634 & w1645;
assign w11714 = ~w1649 & ~w1648;
assign w11715 = ~pi0257 & ~w415;
assign w11716 = ~pi0237 & ~w409;
assign w11717 = w1752 & w11682;
assign w11718 = w1752 & w11683;
assign w11719 = w1098 & w1755;
assign w11720 = w1276 & ~w1656;
assign w11721 = pi0877 & w406;
assign w11722 = w1789 & ~w1639;
assign w11723 = w1789 & ~w11712;
assign w11724 = ~w1844 & ~w1859;
assign w11725 = w1844 & ~pi0265;
assign w11726 = ~w1844 & w1859;
assign w11727 = ~w1912 & w1913;
assign w11728 = ~w1915 & w1916;
assign w11729 = w1917 & ~w1916;
assign w11730 = w1917 & ~w11728;
assign w11731 = ~w1919 & w1920;
assign w11732 = w1921 & ~w1920;
assign w11733 = w1921 & ~w11731;
assign w11734 = w1924 & ~w11732;
assign w11735 = w1924 & ~w11733;
assign w11736 = w1204 & ~w1207;
assign w11737 = ~w1789 & w1639;
assign w11738 = ~w1789 & w11712;
assign w11739 = ~w1630 & ~w1627;
assign w11740 = ~w1933 & ~w1627;
assign w11741 = ~w1933 & w11739;
assign w11742 = w1933 & w1627;
assign w11743 = w1933 & ~w11739;
assign w11744 = ~w1965 & w1966;
assign w11745 = ~w1968 & w1969;
assign w11746 = w1970 & ~w1969;
assign w11747 = w1970 & ~w11745;
assign w11748 = ~w1972 & w1973;
assign w11749 = w1943 & ~w1942;
assign w11750 = w1977 & w1942;
assign w11751 = w1977 & ~w11749;
assign w11752 = ~w2004 & w2005;
assign w11753 = ~w2007 & w2008;
assign w11754 = w2009 & ~w2008;
assign w11755 = w2009 & ~w11753;
assign w11756 = ~w2011 & w2012;
assign w11757 = w1982 & ~w1981;
assign w11758 = w2016 & w1981;
assign w11759 = w2016 & ~w11757;
assign w11760 = pi1747 & pi0997;
assign w11761 = pi1629 & pi0724;
assign w11762 = ~pi1677 & ~pi1050;
assign w11763 = ~pi0760 & w2136;
assign w11764 = w2141 & w2135;
assign w11765 = w11764 & ~pi0966;
assign w11766 = ~pi0995 & w2144;
assign w11767 = w11766 & w2134;
assign w11768 = ~pi0995 & ~pi0966;
assign w11769 = ~pi1345 & ~pi1479;
assign w11770 = ~pi0995 & w2162;
assign w11771 = w11763 & ~pi1050;
assign w11772 = ~pi1677 & w2170;
assign w11773 = w11772 & pi0277;
assign w11774 = w2137 & pi1677;
assign w11775 = ~pi0995 & pi0966;
assign w11776 = w2175 & w2132;
assign w11777 = pi1479 & ~pi1046;
assign w11778 = ~w2164 & ~w2172;
assign w11779 = ~w2216 & w2217;
assign w11780 = ~w2219 & w2220;
assign w11781 = w2221 & ~w2220;
assign w11782 = w2221 & ~w11780;
assign w11783 = ~w2223 & w2224;
assign w11784 = ~w2225 & ~w2224;
assign w11785 = ~w2225 & ~w11783;
assign w11786 = w2194 & w2229;
assign w11787 = pi0153 & pi0195;
assign w11788 = w234 & w2032;
assign w11789 = pi1747 & pi0999;
assign w11790 = ~pi0153 & ~pi0195;
assign w11791 = pi0199 & pi1579;
assign w11792 = ~pi0199 & pi1579;
assign w11793 = ~pi0197 & ~w2251;
assign w11794 = pi1747 & pi0998;
assign w11795 = w1564 & ~w1567;
assign w11796 = pi1713 & ~w2269;
assign w11797 = ~pi0202 & ~w2273;
assign w11798 = ~pi0203 & ~w2277;
assign w11799 = pi1718 & ~w2281;
assign w11800 = pi1711 & ~w2285;
assign w11801 = pi0874 & pi1579;
assign w11802 = ~pi0874 & pi1579;
assign w11803 = pi1716 & ~w2292;
assign w11804 = ~pi0207 & ~w2296;
assign w11805 = pi1716 & ~w2303;
assign w11806 = ~pi0209 & ~w2307;
assign w11807 = pi1713 & ~w2311;
assign w11808 = pi1714 & ~w2315;
assign w11809 = ~pi0212 & ~w2319;
assign w11810 = pi1718 & ~w2323;
assign w11811 = pi1711 & ~w2327;
assign w11812 = w1607 & ~w1602;
assign w11813 = w2331 & ~w1617;
assign w11814 = w1615 & ~w1629;
assign w11815 = pi1709 & ~w2337;
assign w11816 = w1561 & w2340;
assign w11817 = ~w1561 & ~w2340;
assign w11818 = ~pi0219 & ~w2345;
assign w11819 = pi1712 & ~w2349;
assign w11820 = pi0237 & pi0238;
assign w11821 = pi0239 & pi0240;
assign w11822 = ~w11821 & ~pi0221;
assign w11823 = w11821 & pi0221;
assign w11824 = pi0241 & pi0242;
assign w11825 = ~w11824 & ~pi0224;
assign w11826 = w11824 & pi0224;
assign w11827 = w2031 & pi0224;
assign w11828 = w2031 & ~w11825;
assign w11829 = pi1713 & ~w2368;
assign w11830 = ~pi0226 & ~w2372;
assign w11831 = ~pi0227 & ~w2376;
assign w11832 = pi1716 & ~w2380;
assign w11833 = pi1712 & ~w2387;
assign w11834 = ~pi0230 & ~w2391;
assign w11835 = ~pi0231 & ~w2395;
assign w11836 = ~pi0232 & ~w2399;
assign w11837 = pi1718 & ~w2403;
assign w11838 = ~pi0234 & ~w2407;
assign w11839 = pi1714 & ~w2411;
assign w11840 = w11826 & pi0243;
assign w11841 = pi0236 & w2031;
assign w11842 = ~pi0237 & ~pi0238;
assign w11843 = ~pi0239 & w2031;
assign w11844 = ~pi0239 & ~pi0240;
assign w11845 = ~pi0241 & w2031;
assign w11846 = ~pi0241 & ~pi0242;
assign w11847 = ~w11826 & ~pi0243;
assign w11848 = ~w2460 & w2461;
assign w11849 = ~w2463 & w2466;
assign w11850 = w2467 & ~w2466;
assign w11851 = w2467 & ~w11849;
assign w11852 = ~w2469 & w2470;
assign w11853 = w2471 & ~w2470;
assign w11854 = w2471 & ~w11852;
assign w11855 = pi0236 & pi0974;
assign w11856 = ~w1635 & ~w11742;
assign w11857 = ~w1635 & ~w11743;
assign w11858 = pi1718 & ~w2482;
assign w11859 = ~pi0247 & ~w2486;
assign w11860 = ~pi0248 & ~w2490;
assign w11861 = ~w2513 & w2514;
assign w11862 = ~w2516 & w2517;
assign w11863 = w2518 & ~w2517;
assign w11864 = w2518 & ~w11862;
assign w11865 = w2551 & pi1409;
assign w11866 = w2 & ~pi0660;
assign w11867 = pi0302 & pi0303;
assign w11868 = ~w2598 & w2599;
assign w11869 = ~w2601 & w2602;
assign w11870 = w2603 & ~w2602;
assign w11871 = w2603 & ~w11869;
assign w11872 = ~w2631 & w2632;
assign w11873 = ~w2634 & w2635;
assign w11874 = w2636 & ~w2635;
assign w11875 = w2636 & ~w11873;
assign w11876 = ~w2664 & w2665;
assign w11877 = ~w2667 & w2668;
assign w11878 = w2669 & ~w2668;
assign w11879 = w2669 & ~w11877;
assign w11880 = ~pi0274 & ~pi0275;
assign w11881 = ~pi0289 & pi0290;
assign w11882 = ~pi0291 & ~pi0283;
assign w11883 = w2711 & pi0283;
assign w11884 = w2711 & ~w11882;
assign w11885 = ~pi0302 & ~pi0303;
assign w11886 = w2161 & ~pi1621;
assign w11887 = w1538 & ~w1540;
assign w11888 = w1540 & ~pi0101;
assign w11889 = ~w1561 & w1326;
assign w11890 = ~w1568 & ~w2728;
assign w11891 = ~w1606 & w1603;
assign w11892 = ~pi0288 & ~pi0289;
assign w11893 = pi0290 & ~pi0291;
assign w11894 = w11893 & ~pi0283;
assign w11895 = w2161 & ~pi1534;
assign w11896 = ~w11893 & pi0283;
assign w11897 = w11867 & ~pi0284;
assign w11898 = ~w11867 & pi0284;
assign w11899 = pi0288 & pi0289;
assign w11900 = ~pi0290 & pi0291;
assign w11901 = ~pi0295 & ~pi0307;
assign w11902 = ~pi0296 & ~pi0297;
assign w11903 = pi0296 & pi0297;
assign w11904 = w11902 & ~pi0298;
assign w11905 = ~w11902 & pi0298;
assign w11906 = ~pi0306 & ~pi0304;
assign w11907 = pi0306 & pi0304;
assign w11908 = ~w11906 & pi0305;
assign w11909 = w11906 & ~pi0305;
assign w11910 = pi0295 & pi0307;
assign w11911 = w2556 & ~pi0258;
assign w11912 = w11911 & ~pi1250;
assign w11913 = w2839 & ~w2838;
assign w11914 = w11913 & ~pi0097;
assign w11915 = ~pi0138 & ~pi1547;
assign w11916 = w2848 & pi1101;
assign w11917 = ~w11916 & pi1747;
assign w11918 = w2851 & ~w2843;
assign w11919 = w2865 & w2862;
assign w11920 = w19 & ~pi1773;
assign w11921 = ~w2866 & pi1430;
assign w11922 = w2871 & ~pi1672;
assign w11923 = ~w2866 & ~w2874;
assign w11924 = w2866 & pi1802;
assign w11925 = pi1526 & pi1082;
assign w11926 = w2871 & ~pi1666;
assign w11927 = w2866 & pi1805;
assign w11928 = pi1526 & ~pi1075;
assign w11929 = pi1526 & ~pi1182;
assign w11930 = w2866 & pi1783;
assign w11931 = w2871 & pi0022;
assign w11932 = w2871 & pi0124;
assign w11933 = w2866 & pi1801;
assign w11934 = pi1526 & pi1176;
assign w11935 = w2871 & pi0011;
assign w11936 = w2866 & pi1788;
assign w11937 = pi1526 & ~pi1169;
assign w11938 = w2871 & pi0016;
assign w11939 = w2866 & pi1784;
assign w11940 = pi1526 & ~pi1166;
assign w11941 = w2871 & pi0007;
assign w11942 = w2866 & pi1787;
assign w11943 = pi1526 & ~pi1239;
assign w11944 = w2931 & w2862;
assign w11945 = w2932 & pi1788;
assign w11946 = ~w2932 & ~w2935;
assign w11947 = ~w2932 & w2935;
assign w11948 = pi1526 & ~pi1167;
assign w11949 = w2866 & pi1785;
assign w11950 = w2871 & pi0019;
assign w11951 = w2871 & pi0018;
assign w11952 = w2866 & pi1789;
assign w11953 = pi1526 & ~pi1246;
assign w11954 = w2871 & pi0023;
assign w11955 = w2866 & pi1780;
assign w11956 = pi1526 & ~pi1073;
assign w11957 = w2932 & pi1784;
assign w11958 = w2932 & pi1787;
assign w11959 = w2871 & pi0030;
assign w11960 = w2866 & pi1781;
assign w11961 = pi1526 & ~pi1053;
assign w11962 = w2932 & pi1785;
assign w11963 = w2932 & pi1789;
assign w11964 = w2932 & pi1780;
assign w11965 = w2932 & pi1778;
assign w11966 = w2932 & pi1779;
assign w11967 = w2932 & pi1781;
assign w11968 = w2932 & pi1802;
assign w11969 = w2932 & pi1805;
assign w11970 = w11911 & pi1250;
assign w11971 = w2871 & pi0064;
assign w11972 = w2866 & pi1774;
assign w11973 = pi1526 & ~pi1254;
assign w11974 = w2871 & pi0310;
assign w11975 = w2866 & pi1792;
assign w11976 = pi1526 & ~pi1171;
assign w11977 = w2871 & pi0332;
assign w11978 = w2866 & pi1793;
assign w11979 = pi1526 & pi1241;
assign w11980 = w2871 & pi0057;
assign w11981 = w2866 & pi1775;
assign w11982 = pi1526 & ~pi1172;
assign w11983 = w2871 & pi0299;
assign w11984 = w2866 & pi1794;
assign w11985 = pi1526 & pi1077;
assign w11986 = w2871 & pi0286;
assign w11987 = w2866 & pi1795;
assign w11988 = pi1526 & pi1173;
assign w11989 = w2871 & pi0254;
assign w11990 = w2866 & pi1797;
assign w11991 = pi1526 & pi1174;
assign w11992 = pi1526 & pi1093;
assign w11993 = w2866 & pi1798;
assign w11994 = w2871 & pi0223;
assign w11995 = w2871 & pi0154;
assign w11996 = w2866 & pi1799;
assign w11997 = pi1526 & pi1175;
assign w11998 = w2871 & pi0155;
assign w11999 = w2866 & pi1800;
assign w12000 = pi1526 & pi1089;
assign w12001 = w2871 & pi0063;
assign w12002 = w2866 & pi1804;
assign w12003 = pi1526 & pi1179;
assign w12004 = pi1526 & ~pi1180;
assign w12005 = w2866 & pi1777;
assign w12006 = w2871 & pi0049;
assign w12007 = w2871 & pi0027;
assign w12008 = w2866 & pi1782;
assign w12009 = pi1526 & ~pi1055;
assign w12010 = w2865 & w3149;
assign w12011 = ~w3150 & pi1447;
assign w12012 = ~w3150 & ~w3154;
assign w12013 = w3150 & pi1802;
assign w12014 = pi1526 & pi1249;
assign w12015 = w3150 & pi1805;
assign w12016 = pi1526 & ~pi1238;
assign w12017 = ~w1538 & ~w1546;
assign w12018 = w1531 & w3171;
assign w12019 = ~w1531 & ~w3171;
assign w12020 = ~w1537 & ~w1535;
assign w12021 = w3176 & ~w1535;
assign w12022 = w3176 & w12020;
assign w12023 = ~w1530 & ~w12021;
assign w12024 = ~w1530 & ~w12022;
assign w12025 = ~w1533 & ~w12023;
assign w12026 = ~w1533 & ~w12024;
assign w12027 = pi1526 & ~pi1245;
assign w12028 = w3150 & pi1782;
assign w12029 = w2931 & w3149;
assign w12030 = w3188 & pi1780;
assign w12031 = ~w3188 & w3190;
assign w12032 = ~w3188 & ~w3190;
assign w12033 = pi0662 & pi0653;
assign w12034 = pi0654 & pi0650;
assign w12035 = w12034 & pi0648;
assign w12036 = pi0569 & pi0566;
assign w12037 = w12036 & pi0623;
assign w12038 = w3227 & ~w3226;
assign w12039 = ~w3225 & w3224;
assign w12040 = w3222 & w3221;
assign w12041 = ~w3219 & ~w3221;
assign w12042 = ~w3219 & ~w12040;
assign w12043 = ~w3218 & ~w3216;
assign w12044 = w3215 & w3216;
assign w12045 = w3215 & ~w12043;
assign w12046 = ~w3213 & ~w12044;
assign w12047 = ~w3213 & ~w12045;
assign w12048 = ~w3212 & ~w3210;
assign w12049 = w3209 & ~w3210;
assign w12050 = w3209 & w12048;
assign w12051 = pi1569 & pi1459;
assign w12052 = ~pi1697 & pi1143;
assign w12053 = ~w3207 & ~pi1143;
assign w12054 = ~w3207 & ~w12052;
assign w12055 = w3244 & ~w12049;
assign w12056 = w3244 & ~w12050;
assign w12057 = pi0358 & ~w12055;
assign w12058 = pi0358 & ~w12056;
assign w12059 = w12037 & pi0358;
assign w12060 = w3206 & w3247;
assign w12061 = w3249 & ~w12049;
assign w12062 = w3249 & ~w12050;
assign w12063 = w3251 & w12061;
assign w12064 = w3251 & w12062;
assign w12065 = w3259 & ~pi1106;
assign w12066 = ~w3259 & pi1106;
assign w12067 = ~w3263 & w3258;
assign w12068 = ~w3267 & ~pi0717;
assign w12069 = w3263 & ~w3256;
assign w12070 = ~w3270 & ~pi1081;
assign w12071 = w3270 & pi1081;
assign w12072 = ~w3267 & w3278;
assign w12073 = w3255 & ~pi1110;
assign w12074 = ~w3284 & pi0675;
assign w12075 = ~pi1102 & pi0712;
assign w12076 = pi1594 & pi1480;
assign w12077 = w3289 & ~w3254;
assign w12078 = pi0719 & pi0708;
assign w12079 = pi0717 & pi0714;
assign w12080 = ~w3301 & ~w3294;
assign w12081 = ~w3289 & pi1699;
assign w12082 = pi1699 & w3307;
assign w12083 = w2932 & pi1777;
assign w12084 = pi1526 & ~pi1244;
assign w12085 = w3150 & pi1780;
assign w12086 = pi1526 & ~pi1188;
assign w12087 = w3150 & pi1788;
assign w12088 = pi1526 & ~pi1185;
assign w12089 = w3150 & pi1784;
assign w12090 = w3150 & pi1787;
assign w12091 = pi1526 & ~pi1063;
assign w12092 = w3188 & pi1788;
assign w12093 = pi1526 & ~pi1186;
assign w12094 = w3150 & pi1785;
assign w12095 = pi1526 & ~pi1189;
assign w12096 = w3150 & pi1789;
assign w12097 = w3188 & pi1784;
assign w12098 = w3188 & pi1787;
assign w12099 = pi1526 & ~pi1205;
assign w12100 = w3150 & pi1781;
assign w12101 = w3188 & pi1785;
assign w12102 = w3188 & pi1789;
assign w12103 = w3188 & pi1778;
assign w12104 = w3188 & pi1781;
assign w12105 = w3188 & pi1779;
assign w12106 = w2932 & pi1803;
assign w12107 = w2932 & pi1795;
assign w12108 = ~w3446 & ~w3444;
assign w12109 = pi1272 & ~pi0509;
assign w12110 = ~w3443 & ~w3441;
assign w12111 = w3440 & w3441;
assign w12112 = w3440 & ~w12110;
assign w12113 = ~w3438 & ~w12111;
assign w12114 = ~w3438 & ~w12112;
assign w12115 = ~w3437 & w12113;
assign w12116 = ~w3437 & w12114;
assign w12117 = w3462 & pi1119;
assign w12118 = ~w3461 & ~w12113;
assign w12119 = ~w3461 & ~w12114;
assign w12120 = ~w3465 & w3467;
assign w12121 = pi1571 & pi1430;
assign w12122 = ~w3465 & ~pi0386;
assign w12123 = ~w3462 & ~pi1119;
assign w12124 = pi0508 & pi0509;
assign w12125 = pi0387 & pi0386;
assign w12126 = pi0466 & ~pi1690;
assign w12127 = ~w3485 & w3486;
assign w12128 = w3485 & w3488;
assign w12129 = w3498 & pi0533;
assign w12130 = pi0380 & w3492;
assign w12131 = w3509 & ~pi1129;
assign w12132 = ~w3509 & pi1129;
assign w12133 = w3513 & ~pi1028;
assign w12134 = ~w3513 & pi1028;
assign w12135 = w3516 & w3508;
assign w12136 = w3506 & ~pi1130;
assign w12137 = ~w3521 & pi0549;
assign w12138 = w3505 & w3529;
assign w12139 = w3531 & ~w3529;
assign w12140 = w3531 & ~w12138;
assign w12141 = ~w3504 & ~w12139;
assign w12142 = ~w3504 & ~w12140;
assign w12143 = w3533 & ~w3529;
assign w12144 = w3533 & ~w12138;
assign w12145 = pi1572 & pi1447;
assign w12146 = ~w3532 & pi0380;
assign w12147 = w3538 & ~w12143;
assign w12148 = w3538 & ~w12144;
assign w12149 = w12126 & pi0379;
assign w12150 = ~w12149 & pi0470;
assign w12151 = pi1122 & pi0381;
assign w12152 = pi1690 & ~pi0379;
assign w12153 = pi0470 & w3555;
assign w12154 = w3560 & w3564;
assign w12155 = w3567 & pi1626;
assign w12156 = w3582 & ~pi1023;
assign w12157 = ~w3582 & pi1023;
assign w12158 = ~w3586 & w3581;
assign w12159 = ~w3590 & pi0442;
assign w12160 = w3586 & ~w3579;
assign w12161 = ~w3594 & ~pi1274;
assign w12162 = w3594 & pi1274;
assign w12163 = ~w3590 & w3600;
assign w12164 = w3629 & w3625;
assign w12165 = pi0441 & ~pi0384;
assign w12166 = pi1690 & pi0384;
assign w12167 = pi1690 & ~w12165;
assign w12168 = ~pi0441 & ~pi1690;
assign w12169 = w12168 & ~pi0384;
assign w12170 = w3636 & w3640;
assign w12171 = pi0481 & w12166;
assign w12172 = pi0481 & w12167;
assign w12173 = w12168 & w3645;
assign w12174 = ~w12173 & ~pi0383;
assign w12175 = ~w3646 & pi1122;
assign w12176 = w3624 & ~w3635;
assign w12177 = w1844 & ~pi0899;
assign w12178 = ~w3462 & w3472;
assign w12179 = w3666 & pi0386;
assign w12180 = ~w3666 & ~pi0386;
assign w12181 = ~w3673 & ~w12113;
assign w12182 = ~w3673 & ~w12114;
assign w12183 = w3673 & w12113;
assign w12184 = w3673 & w12114;
assign w12185 = w3681 & w3478;
assign w12186 = ~pi1122 & ~pi0388;
assign w12187 = ~w3675 & w3695;
assign w12188 = w2932 & pi1774;
assign w12189 = w2932 & pi1786;
assign w12190 = w2932 & pi1790;
assign w12191 = w2932 & pi1791;
assign w12192 = w2932 & pi1793;
assign w12193 = w2932 & pi1775;
assign w12194 = w2932 & pi1794;
assign w12195 = w2932 & pi1796;
assign w12196 = w2932 & pi1798;
assign w12197 = w2932 & pi1799;
assign w12198 = w2932 & pi1797;
assign w12199 = w2932 & pi1801;
assign w12200 = w2932 & pi1800;
assign w12201 = w2932 & pi1776;
assign w12202 = w2932 & pi1804;
assign w12203 = w2932 & pi1782;
assign w12204 = w2932 & pi1783;
assign w12205 = w3188 & pi1802;
assign w12206 = w3188 & pi1805;
assign w12207 = ~pi1022 & pi1690;
assign w12208 = ~pi0408 & pi1690;
assign w12209 = ~pi0408 & w12207;
assign w12210 = ~pi0408 & pi1122;
assign w12211 = w2556 & w3817;
assign w12212 = pi0410 & ~pi1690;
assign w12213 = pi0410 & ~w12207;
assign w12214 = ~pi0410 & pi1690;
assign w12215 = ~pi0410 & w12207;
assign w12216 = ~w3676 & ~w3688;
assign w12217 = ~pi0412 & pi1122;
assign w12218 = w3675 & pi0413;
assign w12219 = w3626 & pi1122;
assign w12220 = w3586 & ~w3581;
assign w12221 = w2871 & pi0015;
assign w12222 = w3150 & pi1790;
assign w12223 = pi1526 & ~pi1190;
assign w12224 = w3150 & pi1792;
assign w12225 = pi1526 & ~pi1191;
assign w12226 = pi1526 & pi1192;
assign w12227 = w3150 & pi1793;
assign w12228 = pi1526 & ~pi1193;
assign w12229 = w3150 & pi1775;
assign w12230 = w3150 & pi1794;
assign w12231 = pi1526 & pi1276;
assign w12232 = w3150 & pi1795;
assign w12233 = pi1526 & pi1194;
assign w12234 = pi1526 & pi1196;
assign w12235 = w3150 & pi1797;
assign w12236 = pi1526 & pi1264;
assign w12237 = w3150 & pi1798;
assign w12238 = w3150 & pi1799;
assign w12239 = pi1526 & pi1197;
assign w12240 = pi1526 & pi1199;
assign w12241 = w3150 & pi1801;
assign w12242 = pi1526 & pi1036;
assign w12243 = w3150 & pi1804;
assign w12244 = pi1526 & ~pi1202;
assign w12245 = w3150 & pi1777;
assign w12246 = pi1526 & ~pi1240;
assign w12247 = w3150 & pi1783;
assign w12248 = ~w3953 & pi1459;
assign w12249 = ~w3953 & ~w3957;
assign w12250 = w3953 & pi1802;
assign w12251 = pi1526 & pi1057;
assign w12252 = pi1526 & ~pi1221;
assign w12253 = w3953 & pi1805;
assign w12254 = w2932 & pi1792;
assign w12255 = ~w3176 & w1535;
assign w12256 = ~w3176 & ~w12020;
assign w12257 = w3150 & pi1800;
assign w12258 = pi1526 & pi1198;
assign w12259 = ~pi0474 & ~pi0433;
assign w12260 = pi0474 & pi0433;
assign w12261 = w2871 & pi0056;
assign w12262 = w2866 & pi1776;
assign w12263 = pi1526 & ~pi1178;
assign w12264 = w3953 & pi1782;
assign w12265 = pi1526 & ~pi1279;
assign w12266 = ~w4056 & pi1480;
assign w12267 = ~w4056 & ~w4060;
assign w12268 = w4056 & pi1805;
assign w12269 = pi1526 & ~pi1161;
assign w12270 = w2871 & pi1481;
assign w12271 = w2866 & pi1796;
assign w12272 = pi1526 & pi1087;
assign w12273 = pi1526 & ~pi1086;
assign w12274 = w3953 & pi1786;
assign w12275 = w2871 & pi0014;
assign w12276 = w3188 & pi1775;
assign w12277 = ~w4091 & pi0441;
assign w12278 = ~w3624 & pi1690;
assign w12279 = pi0441 & ~pi1690;
assign w12280 = ~w3675 & w4102;
assign w12281 = ~w3676 & w4104;
assign w12282 = w3188 & pi1783;
assign w12283 = w3953 & pi1793;
assign w12284 = pi1526 & pi1213;
assign w12285 = w3188 & pi1801;
assign w12286 = w3188 & pi1797;
assign w12287 = pi1526 & ~pi1181;
assign w12288 = w2866 & pi1779;
assign w12289 = w2871 & pi0028;
assign w12290 = pi0475 & pi0476;
assign w12291 = w12290 & pi0477;
assign w12292 = pi0448 & ~pi0705;
assign w12293 = pi1526 & ~pi1278;
assign w12294 = w3953 & pi1780;
assign w12295 = pi1526 & ~pi1208;
assign w12296 = w3953 & pi1785;
assign w12297 = pi1526 & ~pi1085;
assign w12298 = w3953 & pi1784;
assign w12299 = w3953 & pi1788;
assign w12300 = pi1526 & ~pi1062;
assign w12301 = pi1526 & ~pi1209;
assign w12302 = w3953 & pi1787;
assign w12303 = w4186 & pi1788;
assign w12304 = ~w4186 & ~w4188;
assign w12305 = ~w4186 & w4188;
assign w12306 = w3953 & pi1789;
assign w12307 = pi1526 & ~pi1210;
assign w12308 = w4186 & pi1784;
assign w12309 = w4186 & pi1787;
assign w12310 = w2871 & pi0046;
assign w12311 = w2866 & pi1778;
assign w12312 = pi1526 & ~pi1067;
assign w12313 = pi1526 & ~pi1223;
assign w12314 = w3953 & pi1781;
assign w12315 = w4186 & pi1785;
assign w12316 = w4186 & pi1780;
assign w12317 = w4186 & pi1778;
assign w12318 = w4186 & pi1779;
assign w12319 = w4186 & pi1781;
assign w12320 = pi0448 & pi0467;
assign w12321 = w12320 & pi0479;
assign w12322 = w12321 & pi0478;
assign w12323 = ~pi0473 & pi0465;
assign w12324 = pi0473 & ~pi0465;
assign w12325 = ~pi0705 & ~pi0465;
assign w12326 = ~pi0705 & ~w12323;
assign w12327 = ~pi0466 & w3681;
assign w12328 = w3675 & ~pi0466;
assign w12329 = ~w3471 & w4273;
assign w12330 = ~pi0448 & ~pi0467;
assign w12331 = ~w12320 & ~pi0705;
assign w12332 = pi0380 & pi0562;
assign w12333 = w12332 & w3492;
assign w12334 = ~pi0562 & w12141;
assign w12335 = ~pi0562 & w12142;
assign w12336 = w3491 & w12147;
assign w12337 = w3491 & w12148;
assign w12338 = ~w12333 & ~pi0468;
assign w12339 = ~w12332 & w3492;
assign w12340 = ~pi0562 & pi0468;
assign w12341 = w4287 & ~w3492;
assign w12342 = w4287 & ~w12339;
assign w12343 = ~w3491 & w4288;
assign w12344 = w3544 & w3551;
assign w12345 = w4305 & ~pi0560;
assign w12346 = w12345 & ~pi1679;
assign w12347 = ~pi1679 & pi0472;
assign w12348 = pi0472 & ~w4309;
assign w12349 = w4299 & w4311;
assign w12350 = w4316 & ~pi1129;
assign w12351 = ~w4316 & pi1129;
assign w12352 = ~w4320 & w4315;
assign w12353 = w4313 & pi1083;
assign w12354 = ~w4313 & ~pi1083;
assign w12355 = w4324 & pi1130;
assign w12356 = ~w4324 & ~pi1130;
assign w12357 = ~w4299 & w4350;
assign w12358 = ~w4348 & ~w4312;
assign w12359 = w4355 & ~w4356;
assign w12360 = ~w4308 & ~pi0472;
assign w12361 = w4308 & pi0472;
assign w12362 = ~w4355 & ~w4361;
assign w12363 = ~pi0473 & ~pi0705;
assign w12364 = ~pi0474 & ~pi0705;
assign w12365 = ~pi0475 & ~pi0705;
assign w12366 = ~pi0475 & ~pi0476;
assign w12367 = ~w12290 & ~pi0477;
assign w12368 = ~w12321 & ~pi0478;
assign w12369 = ~w12320 & ~pi0479;
assign w12370 = ~w3440 & ~w3441;
assign w12371 = ~w3440 & w12110;
assign w12372 = w3681 & ~pi0484;
assign w12373 = w4389 & pi0480;
assign w12374 = w3681 & w4391;
assign w12375 = w3636 & w4395;
assign w12376 = ~w3636 & w4397;
assign w12377 = w3614 & ~w4400;
assign w12378 = pi0482 & pi1122;
assign w12379 = ~w3496 & w3492;
assign w12380 = w4409 & pi0483;
assign w12381 = w3505 & ~w3528;
assign w12382 = w3530 & w4414;
assign w12383 = w3492 & w4416;
assign w12384 = ~pi0484 & ~w4389;
assign w12385 = ~pi0549 & ~pi0485;
assign w12386 = w4428 & w4414;
assign w12387 = ~w4406 & pi0486;
assign w12388 = ~w3491 & w4435;
assign w12389 = ~w3492 & ~pi0486;
assign w12390 = ~w4414 & w4437;
assign w12391 = w3188 & pi1774;
assign w12392 = w3188 & pi1786;
assign w12393 = w3188 & pi1790;
assign w12394 = w3188 & pi1791;
assign w12395 = w3188 & pi1792;
assign w12396 = w3188 & pi1793;
assign w12397 = w3188 & pi1794;
assign w12398 = w3188 & pi1795;
assign w12399 = w3188 & pi1796;
assign w12400 = w3188 & pi1798;
assign w12401 = w3188 & pi1799;
assign w12402 = w3188 & pi1800;
assign w12403 = w3188 & pi1776;
assign w12404 = w3188 & pi1804;
assign w12405 = w3188 & pi1803;
assign w12406 = w3188 & pi1777;
assign w12407 = w3188 & pi1782;
assign w12408 = w4186 & pi1802;
assign w12409 = w4186 & pi1805;
assign w12410 = ~pi1027 & pi1679;
assign w12411 = ~pi0506 & pi1679;
assign w12412 = ~pi0506 & w12410;
assign w12413 = ~pi0506 & pi1131;
assign w12414 = ~pi0408 & ~pi0507;
assign w12415 = ~w4558 & pi0508;
assign w12416 = ~w3676 & ~w4569;
assign w12417 = ~w3681 & ~pi0509;
assign w12418 = ~w3675 & w4579;
assign w12419 = w3626 & ~pi0442;
assign w12420 = ~w3602 & ~w4582;
assign w12421 = pi0510 & pi1122;
assign w12422 = pi0511 & ~pi1679;
assign w12423 = pi0511 & ~w12410;
assign w12424 = ~pi0511 & pi1679;
assign w12425 = ~pi0511 & w12410;
assign w12426 = w3491 & pi0512;
assign w12427 = w4321 & ~w4603;
assign w12428 = pi0513 & pi1131;
assign w12429 = ~pi0513 & ~pi0514;
assign w12430 = w4320 & ~w4315;
assign w12431 = ~pi0514 & ~w4610;
assign w12432 = w4056 & pi1802;
assign w12433 = pi1526 & pi1159;
assign w12434 = w2866 & pi1786;
assign w12435 = pi1526 & ~pi1168;
assign w12436 = w2866 & pi1790;
assign w12437 = pi1526 & ~pi1170;
assign w12438 = w2871 & pi0953;
assign w12439 = w2866 & pi1791;
assign w12440 = pi1526 & ~pi1247;
assign w12441 = pi1526 & pi1177;
assign w12442 = w2866 & pi1803;
assign w12443 = w2871 & pi0194;
assign w12444 = pi1526 & ~pi1207;
assign w12445 = w3953 & pi1774;
assign w12446 = pi1526 & ~pi1071;
assign w12447 = w3953 & pi1790;
assign w12448 = pi1526 & ~pi1211;
assign w12449 = w3953 & pi1791;
assign w12450 = pi1526 & ~pi1212;
assign w12451 = w3953 & pi1792;
assign w12452 = pi1526 & pi1214;
assign w12453 = w3953 & pi1794;
assign w12454 = pi1526 & pi1216;
assign w12455 = w3953 & pi1796;
assign w12456 = w3953 & pi1798;
assign w12457 = pi1526 & pi1217;
assign w12458 = w3953 & pi1799;
assign w12459 = pi1526 & pi1218;
assign w12460 = w3953 & pi1803;
assign w12461 = pi1526 & pi1232;
assign w12462 = w3953 & pi1775;
assign w12463 = pi1526 & ~pi1064;
assign w12464 = w3953 & pi1804;
assign w12465 = pi1526 & pi1266;
assign w12466 = pi1526 & ~pi1282;
assign w12467 = w3953 & pi1777;
assign w12468 = w4186 & pi1789;
assign w12469 = ~w3525 & ~w3529;
assign w12470 = ~w3525 & ~w12138;
assign w12471 = w4760 & ~w12469;
assign w12472 = w4760 & ~w12470;
assign w12473 = ~w3498 & ~pi0533;
assign w12474 = ~w3491 & ~w4764;
assign w12475 = ~w3532 & pi1679;
assign w12476 = pi1526 & ~pi1200;
assign w12477 = w3150 & pi1776;
assign w12478 = w1226 & pi1480;
assign w12479 = w3150 & pi1796;
assign w12480 = pi1526 & pi1195;
assign w12481 = w4186 & pi1777;
assign w12482 = w4186 & pi1794;
assign w12483 = w4186 & pi1801;
assign w12484 = w4186 & pi1798;
assign w12485 = w4308 & ~pi1083;
assign w12486 = w4308 & ~w12353;
assign w12487 = ~w4813 & ~pi0541;
assign w12488 = w4813 & pi0541;
assign w12489 = w4056 & pi1803;
assign w12490 = pi1526 & pi1269;
assign w12491 = w4186 & pi1791;
assign w12492 = w4056 & pi1799;
assign w12493 = pi1526 & pi1275;
assign w12494 = w4056 & pi1795;
assign w12495 = pi1526 & pi1154;
assign w12496 = w4056 & pi1779;
assign w12497 = pi1526 & ~pi1162;
assign w12498 = pi1526 & ~pi1204;
assign w12499 = w3150 & pi1779;
assign w12500 = ~w3491 & w4425;
assign w12501 = ~w3492 & ~pi0549;
assign w12502 = w4056 & pi1780;
assign w12503 = pi1526 & ~pi1343;
assign w12504 = w4056 & pi1784;
assign w12505 = pi1526 & ~pi1316;
assign w12506 = w4896 & ~pi1141;
assign w12507 = ~w4896 & pi1141;
assign w12508 = ~w4900 & w4895;
assign w12509 = w4893 & pi1033;
assign w12510 = ~w4893 & ~pi1033;
assign w12511 = w4904 & pi1142;
assign w12512 = ~w4904 & ~pi1142;
assign w12513 = w5574 & ~pi0552;
assign w12514 = w4892 & w4926;
assign w12515 = ~pi0589 & ~pi0590;
assign w12516 = w6235 & ~pi0655;
assign w12517 = ~pi0568 & ~pi0631;
assign w12518 = w12517 & ~pi0642;
assign w12519 = w12518 & ~pi0552;
assign w12520 = ~w12518 & pi0552;
assign w12521 = pi1143 & ~w4928;
assign w12522 = pi1143 & ~w4892;
assign w12523 = ~w4941 & ~w4940;
assign w12524 = w4056 & pi1788;
assign w12525 = pi1526 & ~pi1151;
assign w12526 = w4056 & pi1787;
assign w12527 = pi1526 & ~pi1312;
assign w12528 = w4056 & pi1785;
assign w12529 = pi1526 & ~pi1311;
assign w12530 = w4056 & pi1789;
assign w12531 = pi1526 & ~pi1152;
assign w12532 = w4056 & pi1778;
assign w12533 = pi1526 & ~pi1332;
assign w12534 = w4056 & pi1781;
assign w12535 = pi1526 & ~pi1333;
assign w12536 = pi1526 & ~pi1203;
assign w12537 = w3150 & pi1778;
assign w12538 = ~w4305 & pi0560;
assign w12539 = w3491 & pi0560;
assign w12540 = ~w3492 & ~w5002;
assign w12541 = ~w4414 & w5003;
assign w12542 = ~w3492 & w5006;
assign w12543 = ~pi0380 & ~pi0562;
assign w12544 = pi0552 & pi0649;
assign w12545 = ~w5019 & w5020;
assign w12546 = pi0649 & ~w4892;
assign w12547 = w5020 & ~w4892;
assign w12548 = w5020 & w12546;
assign w12549 = w5019 & w5025;
assign w12550 = ~w5023 & ~w5021;
assign w12551 = ~w4347 & w5034;
assign w12552 = ~w5032 & ~w5031;
assign w12553 = ~w4406 & ~w5040;
assign w12554 = ~w5041 & pi0565;
assign w12555 = w3492 & w4305;
assign w12556 = ~pi0569 & ~pi0566;
assign w12557 = ~pi0622 & ~pi0567;
assign w12558 = ~w3516 & ~w3508;
assign w12559 = ~pi1697 & w5066;
assign w12560 = ~w3242 & w5068;
assign w12561 = ~w3215 & ~w3216;
assign w12562 = ~w3215 & w12043;
assign w12563 = ~w3251 & ~w5073;
assign w12564 = w4186 & pi1774;
assign w12565 = w4186 & pi1786;
assign w12566 = w4186 & pi1790;
assign w12567 = w4186 & pi1792;
assign w12568 = w4186 & pi1793;
assign w12569 = w4186 & pi1775;
assign w12570 = w4186 & pi1796;
assign w12571 = w4186 & pi1797;
assign w12572 = w4186 & pi1795;
assign w12573 = w4186 & pi1800;
assign w12574 = w4186 & pi1799;
assign w12575 = w4186 & pi1803;
assign w12576 = w4186 & pi1776;
assign w12577 = w4186 & pi1804;
assign w12578 = w4186 & pi1782;
assign w12579 = w4186 & pi1783;
assign w12580 = ~pi1032 & pi1697;
assign w12581 = ~pi0586 & pi1697;
assign w12582 = ~pi0586 & w12580;
assign w12583 = ~pi0586 & pi1143;
assign w12584 = w3492 & w3494;
assign w12585 = ~w5056 & pi0587;
assign w12586 = ~pi1679 & ~pi0541;
assign w12587 = w4329 & ~w5186;
assign w12588 = pi0588 & pi1131;
assign w12589 = ~w3242 & ~w4930;
assign w12590 = w4930 & ~w4901;
assign w12591 = pi0590 & pi1143;
assign w12592 = w4900 & ~w4895;
assign w12593 = w1226 & pi1459;
assign w12594 = w4056 & pi1774;
assign w12595 = pi1526 & ~pi1149;
assign w12596 = pi0594 & ~pi1697;
assign w12597 = pi0594 & ~w12580;
assign w12598 = ~pi0594 & pi1697;
assign w12599 = ~pi0594 & w12580;
assign w12600 = w4056 & pi1790;
assign w12601 = pi1526 & ~pi1153;
assign w12602 = w4056 & pi1791;
assign w12603 = pi1526 & ~pi1305;
assign w12604 = w4056 & pi1792;
assign w12605 = pi1526 & ~pi1284;
assign w12606 = w4056 & pi1793;
assign w12607 = pi1526 & pi1331;
assign w12608 = w4056 & pi1775;
assign w12609 = pi1526 & ~pi1292;
assign w12610 = w4056 & pi1794;
assign w12611 = pi1526 & pi1283;
assign w12612 = w4056 & pi1786;
assign w12613 = pi1526 & ~pi1150;
assign w12614 = w4056 & pi1797;
assign w12615 = pi1526 & pi1156;
assign w12616 = w4056 & pi1798;
assign w12617 = pi1526 & pi1157;
assign w12618 = w4056 & pi1796;
assign w12619 = pi1526 & pi1155;
assign w12620 = w4056 & pi1801;
assign w12621 = pi1526 & pi1346;
assign w12622 = w4056 & pi1800;
assign w12623 = pi1526 & pi1158;
assign w12624 = w4056 & pi1776;
assign w12625 = pi1526 & ~pi1344;
assign w12626 = w4056 & pi1804;
assign w12627 = pi1526 & pi1160;
assign w12628 = w4056 & pi1777;
assign w12629 = pi1526 & ~pi1263;
assign w12630 = w4056 & pi1782;
assign w12631 = pi1526 & ~pi1163;
assign w12632 = w4056 & pi1783;
assign w12633 = pi1526 & ~pi1183;
assign w12634 = pi1526 & ~pi1065;
assign w12635 = w3150 & pi1774;
assign w12636 = pi1526 & ~pi1187;
assign w12637 = w3150 & pi1786;
assign w12638 = pi1526 & ~pi1248;
assign w12639 = w3150 & pi1791;
assign w12640 = w1226 & pi1430;
assign w12641 = pi1526 & pi1201;
assign w12642 = w3150 & pi1803;
assign w12643 = w1226 & pi1447;
assign w12644 = ~w4308 & pi1131;
assign w12645 = ~w1519 & ~w1510;
assign w12646 = w1359 & w5418;
assign w12647 = pi1697 & ~pi0645;
assign w12648 = w5422 & w12061;
assign w12649 = w5422 & w12062;
assign w12650 = ~w5421 & w5424;
assign w12651 = w5421 & w5426;
assign w12652 = ~w3491 & w5057;
assign w12653 = ~w3492 & ~pi0622;
assign w12654 = ~w12036 & ~pi0623;
assign w12655 = ~w3209 & w3210;
assign w12656 = ~w3209 & ~w12048;
assign w12657 = w5442 & pi1781;
assign w12658 = ~w5442 & ~w5444;
assign w12659 = ~w5442 & w5444;
assign w12660 = pi1526 & ~pi1220;
assign w12661 = w3953 & pi1776;
assign w12662 = w3242 & ~pi1033;
assign w12663 = w3242 & ~w12509;
assign w12664 = ~w4932 & ~pi0627;
assign w12665 = w4932 & pi0627;
assign w12666 = w5442 & pi1779;
assign w12667 = pi1526 & pi1219;
assign w12668 = w3953 & pi1800;
assign w12669 = pi0646 & ~w30;
assign w12670 = ~w12669 & ~w5490;
assign w12671 = w4923 & ~w4935;
assign w12672 = w3953 & pi1778;
assign w12673 = pi1526 & ~pi1222;
assign w12674 = w5442 & pi1780;
assign w12675 = w5442 & pi1788;
assign w12676 = w5442 & pi1784;
assign w12677 = w5442 & pi1787;
assign w12678 = w5442 & pi1785;
assign w12679 = w5442 & pi1789;
assign w12680 = w3953 & pi1779;
assign w12681 = pi1526 & ~pi1281;
assign w12682 = w5442 & pi1778;
assign w12683 = w4923 & w5560;
assign w12684 = ~w12517 & pi0642;
assign w12685 = w5563 & pi1143;
assign w12686 = ~pi0645 & w3243;
assign w12687 = w5574 & ~w12061;
assign w12688 = w5574 & ~w12062;
assign w12689 = w5573 & ~w5576;
assign w12690 = ~pi0645 & w3251;
assign w12691 = ~pi0646 & pi1747;
assign w12692 = w3572 & ~w1231;
assign w12693 = ~w12034 & ~pi0648;
assign w12694 = ~pi0649 & ~w4892;
assign w12695 = ~w5597 & ~w5596;
assign w12696 = pi0649 & pi1143;
assign w12697 = ~w4892 & ~pi1143;
assign w12698 = ~w4892 & ~w12696;
assign w12699 = w4928 & pi1143;
assign w12700 = ~w3222 & ~w3221;
assign w12701 = ~pi0654 & ~pi0650;
assign w12702 = w5442 & pi1802;
assign w12703 = w5442 & pi1805;
assign w12704 = ~pi0662 & ~pi0653;
assign w12705 = w3225 & ~w3224;
assign w12706 = w4909 & ~w4933;
assign w12707 = pi0655 & pi1143;
assign w12708 = w3953 & pi1795;
assign w12709 = pi1526 & pi1215;
assign w12710 = w3953 & pi1797;
assign w12711 = pi1526 & pi1066;
assign w12712 = w3953 & pi1801;
assign w12713 = pi1526 & pi1056;
assign w12714 = w3953 & pi1783;
assign w12715 = pi1526 & ~pi1224;
assign w12716 = w2551 & ~pi1409;
assign w12717 = pi1090 & pi1101;
assign w12718 = w5694 & ~pi1106;
assign w12719 = ~w5694 & pi1106;
assign w12720 = ~w5698 & pi1107;
assign w12721 = w5698 & ~pi1107;
assign w12722 = ~pi1102 & ~pi0720;
assign w12723 = w5746 & w5743;
assign w12724 = ~w5736 & ~pi1699;
assign w12725 = w5750 & pi1699;
assign w12726 = w5750 & ~w12724;
assign w12727 = ~w5736 & w5754;
assign w12728 = ~w5753 & ~w5755;
assign w12729 = pi1102 & w5758;
assign w12730 = pi1699 & w5764;
assign w12731 = pi1102 & w5765;
assign w12732 = w3301 & pi0359;
assign w12733 = pi0664 & ~pi1699;
assign w12734 = ~w5775 & w5776;
assign w12735 = w5775 & w5778;
assign w12736 = w5442 & pi1799;
assign w12737 = w5442 & pi1795;
assign w12738 = ~w5703 & ~pi0669;
assign w12739 = ~w5743 & pi0669;
assign w12740 = w5442 & pi1774;
assign w12741 = w5442 & pi1792;
assign w12742 = ~w5842 & w5843;
assign w12743 = ~w5845 & w5846;
assign w12744 = w5847 & ~w5846;
assign w12745 = w5847 & ~w12743;
assign w12746 = ~w5849 & w5850;
assign w12747 = w5851 & ~w5850;
assign w12748 = w5851 & ~w12746;
assign w12749 = w5863 & ~pi0715;
assign w12750 = ~pi0674 & w5867;
assign w12751 = ~w5799 & w5870;
assign w12752 = ~w5869 & w5871;
assign w12753 = ~w5862 & ~w5868;
assign w12754 = w12079 & ~pi1699;
assign w12755 = ~w5877 & pi0675;
assign w12756 = ~w3294 & w5880;
assign w12757 = pi0678 & pi1111;
assign w12758 = ~w12757 & ~pi0675;
assign w12759 = ~w5882 & w5883;
assign w12760 = w5897 & ~w5896;
assign w12761 = ~w5902 & w5903;
assign w12762 = ~w5905 & w5906;
assign w12763 = w5907 & ~w5906;
assign w12764 = w5907 & ~w12762;
assign w12765 = ~w5911 & w5914;
assign w12766 = w5917 & ~w5914;
assign w12767 = w5917 & ~w12765;
assign w12768 = w5920 & ~w12766;
assign w12769 = w5920 & ~w12767;
assign w12770 = w5926 & w3625;
assign w12771 = ~w5924 & ~w5929;
assign w12772 = ~w3280 & ~w3276;
assign w12773 = ~w3294 & ~w5948;
assign w12774 = w5442 & pi1786;
assign w12775 = w5442 & pi1790;
assign w12776 = w5442 & pi1791;
assign w12777 = w5442 & pi1793;
assign w12778 = w5442 & pi1775;
assign w12779 = w5442 & pi1794;
assign w12780 = w5442 & pi1796;
assign w12781 = w5442 & pi1797;
assign w12782 = w5442 & pi1798;
assign w12783 = w5442 & pi1801;
assign w12784 = w5442 & pi1800;
assign w12785 = w5442 & pi1804;
assign w12786 = w5442 & pi1776;
assign w12787 = w5442 & pi1783;
assign w12788 = w5442 & pi1782;
assign w12789 = w3559 & pi1747;
assign w12790 = ~w3560 & w3564;
assign w12791 = ~pi1105 & pi1699;
assign w12792 = ~pi0697 & pi1699;
assign w12793 = ~pi0697 & w12791;
assign w12794 = ~pi0697 & pi1111;
assign w12795 = ~w5882 & ~w5867;
assign w12796 = ~w3294 & pi0699;
assign w12797 = ~w5882 & w6068;
assign w12798 = pi0700 & ~pi1699;
assign w12799 = pi0700 & ~w12791;
assign w12800 = ~pi0700 & pi1699;
assign w12801 = ~pi0700 & w12791;
assign w12802 = w27 & pi1747;
assign w12803 = w27 & w12691;
assign w12804 = w28 & w12803;
assign w12805 = w28 & w12802;
assign w12806 = pi1747 & pi1748;
assign w12807 = w5442 & pi1777;
assign w12808 = w5442 & pi1803;
assign w12809 = ~w3294 & w6095;
assign w12810 = ~w5882 & w6098;
assign w12811 = ~w3254 & ~w3294;
assign w12812 = w3263 & ~w3258;
assign w12813 = w6105 & ~w6104;
assign w12814 = pi0720 & pi0709;
assign w12815 = ~w6114 & ~w6117;
assign w12816 = ~w3294 & ~w6125;
assign w12817 = w4301 & w4302;
assign w12818 = w6149 & ~w6148;
assign w12819 = ~w6154 & w6155;
assign w12820 = ~w6157 & w6158;
assign w12821 = w6159 & ~w6158;
assign w12822 = w6159 & ~w12820;
assign w12823 = ~w6163 & w6166;
assign w12824 = w6169 & ~w6166;
assign w12825 = w6169 & ~w12823;
assign w12826 = w6172 & ~w12824;
assign w12827 = w6172 & ~w12825;
assign w12828 = ~w6176 & ~w6137;
assign w12829 = ~w5877 & pi0712;
assign w12830 = w12757 & pi0675;
assign w12831 = ~w12830 & ~pi0712;
assign w12832 = ~w6209 & w6210;
assign w12833 = ~w6212 & w6213;
assign w12834 = w6214 & ~w6213;
assign w12835 = w6214 & ~w12833;
assign w12836 = ~w6216 & w6219;
assign w12837 = w6222 & ~w6219;
assign w12838 = w6222 & ~w12836;
assign w12839 = w6225 & ~w12837;
assign w12840 = w6225 & ~w12838;
assign w12841 = ~w6238 & w1493;
assign w12842 = ~w6242 & w6244;
assign w12843 = pi0714 & ~pi1111;
assign w12844 = pi0714 & ~w3254;
assign w12845 = ~w3294 & ~w6248;
assign w12846 = ~w3254 & ~pi0714;
assign w12847 = ~w5799 & ~pi0715;
assign w12848 = ~w5753 & ~w6256;
assign w12849 = ~w5869 & ~w6259;
assign w12850 = w29 & w12803;
assign w12851 = w29 & w12802;
assign w12852 = ~w3267 & w3291;
assign w12853 = ~pi0717 & w3294;
assign w12854 = ~pi0717 & w3254;
assign w12855 = w3264 & ~pi0719;
assign w12856 = ~w5877 & pi0720;
assign w12857 = ~w3254 & ~pi0720;
assign w12858 = ~w5882 & w6299;
assign w12859 = ~w6321 & w6322;
assign w12860 = ~w6324 & w6325;
assign w12861 = w6326 & ~w6325;
assign w12862 = w6326 & ~w12860;
assign w12863 = ~w6328 & w6331;
assign w12864 = w6334 & ~w6331;
assign w12865 = w6334 & ~w12863;
assign w12866 = w6337 & ~w12864;
assign w12867 = w6337 & ~w12865;
assign w12868 = ~pi0674 & w5743;
assign w12869 = ~w12868 & w1586;
assign w12870 = w3572 & pi0722;
assign w12871 = ~w3572 & ~pi1738;
assign w12872 = ~w3572 & pi1738;
assign w12873 = ~w6349 & w6389;
assign w12874 = ~w3572 & pi0733;
assign w12875 = w3572 & pi0723;
assign w12876 = ~pi1677 & pi1050;
assign w12877 = pi0788 & pi0783;
assign w12878 = ~w6441 & w6431;
assign w12879 = ~w6443 & w6426;
assign w12880 = w6444 & ~w6426;
assign w12881 = w6444 & ~w12879;
assign w12882 = ~w6421 & w6418;
assign w12883 = w6451 & w6448;
assign w12884 = w6415 & ~w6454;
assign w12885 = w3572 & pi0727;
assign w12886 = w3572 & pi0729;
assign w12887 = ~w3572 & pi0746;
assign w12888 = w3572 & pi0730;
assign w12889 = ~w3572 & pi0734;
assign w12890 = w3572 & pi0731;
assign w12891 = ~w3572 & pi0745;
assign w12892 = w3572 & pi0732;
assign w12893 = w3572 & pi0733;
assign w12894 = w3572 & pi0734;
assign w12895 = w3572 & pi0735;
assign w12896 = w3572 & pi0736;
assign w12897 = w3572 & pi0737;
assign w12898 = w3572 & pi0738;
assign w12899 = w6451 & ~w6534;
assign w12900 = ~w3572 & pi0735;
assign w12901 = w3572 & pi0744;
assign w12902 = w3572 & pi0745;
assign w12903 = w3572 & pi0746;
assign w12904 = ~pi0048 & w623;
assign w12905 = ~pi0048 & ~w11371;
assign w12906 = pi0747 & ~w623;
assign w12907 = pi0747 & w11371;
assign w12908 = ~w634 & ~w12904;
assign w12909 = ~w634 & ~w12905;
assign w12910 = w1844 & ~pi0580;
assign w12911 = w1844 & ~pi0581;
assign w12912 = w1844 & pi1271;
assign w12913 = w1844 & ~pi0578;
assign w12914 = w1844 & ~pi0454;
assign w12915 = ~pi1761 & ~pi1762;
assign w12916 = ~pi1758 & w6605;
assign w12917 = w2931 & w6608;
assign w12918 = w2865 & w6608;
assign w12919 = ~pi1758 & w2862;
assign w12920 = w2865 & w6605;
assign w12921 = w2931 & w6605;
assign w12922 = ~pi1758 & w6608;
assign w12923 = pi1758 & w2862;
assign w12924 = pi1758 & w6605;
assign w12925 = pi1758 & w6608;
assign w12926 = w1844 & ~pi0573;
assign w12927 = w1844 & pi1258;
assign w12928 = w1844 & ~pi0531;
assign w12929 = w1844 & ~pi0459;
assign w12930 = w1844 & ~pi0456;
assign w12931 = w1844 & pi1034;
assign w12932 = w6719 & ~w2133;
assign w12933 = w2165 & pi1670;
assign w12934 = pi1345 & ~pi1544;
assign w12935 = w12934 & w6728;
assign w12936 = w12935 & pi1673;
assign w12937 = w12934 & ~w6728;
assign w12938 = w1844 & ~pi0528;
assign w12939 = pi1345 & ~pi1665;
assign w12940 = w12935 & pi1532;
assign w12941 = w12937 & ~pi0764;
assign w12942 = w12935 & pi1527;
assign w12943 = w12937 & pi0765;
assign w12944 = w12935 & pi1522;
assign w12945 = w12937 & ~pi0766;
assign w12946 = w1844 & pi0967;
assign w12947 = w1844 & ~pi0530;
assign w12948 = w1844 & ~pi0656;
assign w12949 = w1844 & pi1259;
assign w12950 = w1844 & ~pi0527;
assign w12951 = ~pi1674 & ~pi0937;
assign w12952 = w2165 & ~pi1670;
assign w12953 = ~w2133 & ~w6810;
assign w12954 = w2141 & w2148;
assign w12955 = pi0984 & pi0278;
assign w12956 = ~w6842 & w6843;
assign w12957 = ~w6845 & w6846;
assign w12958 = w6847 & ~w6846;
assign w12959 = w6847 & ~w12957;
assign w12960 = ~w6849 & w6850;
assign w12961 = w6851 & ~w6850;
assign w12962 = w6851 & ~w12960;
assign w12963 = ~pi0050 & w623;
assign w12964 = ~pi0050 & ~w11371;
assign w12965 = pi0777 & ~w623;
assign w12966 = pi0777 & w11371;
assign w12967 = ~w8024 & pi0699;
assign w12968 = w8070 & ~w8069;
assign w12969 = w8124 & ~w8123;
assign w12970 = w8172 & ~w8171;
assign w12971 = w8170 & w8169;
assign w12972 = ~w8098 & ~w8096;
assign w12973 = ~w9896 & w9898;
assign w12974 = w8010 & w10282;
assign w12975 = ~w11368 & ~pi1646;
assign w12976 = ~w633 & w635;
assign w12977 = ~w658 & w659;
assign w12978 = w8024 & ~pi0699;
assign w12979 = w8028 & w8033;
assign w12980 = w8122 & w8121;
assign w12981 = w8119 & w8134;
assign w12982 = w8167 & w8182;
assign w12983 = w12972 & ~w8096;
assign w12984 = (~w8096 & w12972) | (~w8096 & ~w8092) | (w12972 & ~w8092);
assign w12985 = ~pi1458 & pi0772;
assign w12986 = pi1458 & pi0748;
assign w12987 = ~pi1458 & pi0822;
assign w12988 = pi1458 & pi0845;
assign w12989 = ~pi1458 & pi0823;
assign w12990 = pi1458 & pi0846;
assign w12991 = ~pi1458 & pi0824;
assign w12992 = pi1458 & pi0847;
assign w12993 = ~pi1699 & w5751;
assign w12994 = ~w8023 & w8022;
assign one = 1;
assign po0000 = pi0661;// level 0
assign po0001 = pi0561;// level 0
assign po0002 = pi0666;// level 0
assign po0003 = pi0643;// level 0
assign po0004 = pi0902;// level 0
assign po0005 = pi0912;// level 0
assign po0006 = pi0911;// level 0
assign po0007 = pi0782;// level 0
assign po0008 = pi0784;// level 0
assign po0009 = pi0962;// level 0
assign po0010 = pi0972;// level 0
assign po0011 = pi0961;// level 0
assign po0012 = pi0964;// level 0
assign po0013 = pi0988;// level 0
assign po0014 = pi1226;// level 0
assign po0015 = pi0989;// level 0
assign po0016 = pi0905;// level 0
assign po0017 = pi0914;// level 0
assign po0018 = pi0913;// level 0
assign po0019 = pi0910;// level 0
assign po0020 = pi0909;// level 0
assign po0021 = pi0908;// level 0
assign po0022 = pi0781;// level 0
assign po0023 = pi0769;// level 0
assign po0024 = pi0906;// level 0
assign po0025 = pi0882;// level 0
assign po0026 = pi0888;// level 0
assign po0027 = pi0955;// level 0
assign po0028 = pi0907;// level 0
assign po0029 = pi0956;// level 0
assign po0030 = pi0951;// level 0
assign po0031 = pi0952;// level 0
assign po0032 = ~w38;// level 10
assign po0033 = ~w41;// level 10
assign po0034 = ~w44;// level 10
assign po0035 = ~w47;// level 10
assign po0036 = ~w50;// level 10
assign po0037 = ~w53;// level 10
assign po0038 = ~w56;// level 10
assign po0039 = ~w59;// level 10
assign po0040 = ~w62;// level 10
assign po0041 = ~w65;// level 10
assign po0042 = ~w68;// level 10
assign po0043 = ~w71;// level 10
assign po0044 = ~w74;// level 10
assign po0045 = ~w77;// level 10
assign po0046 = ~w80;// level 10
assign po0047 = ~w83;// level 10
assign po0048 = ~w86;// level 10
assign po0049 = ~w89;// level 10
assign po0050 = ~w92;// level 10
assign po0051 = ~w95;// level 10
assign po0052 = ~w98;// level 10
assign po0053 = ~w101;// level 10
assign po0054 = ~w104;// level 10
assign po0055 = ~w107;// level 10
assign po0056 = ~w110;// level 10
assign po0057 = ~w113;// level 10
assign po0058 = ~w116;// level 10
assign po0059 = ~w119;// level 10
assign po0060 = ~w122;// level 10
assign po0061 = ~w125;// level 10
assign po0062 = ~w128;// level 10
assign po0063 = ~w131;// level 10
assign po0064 = pi0256;// level 0
assign po0065 = pi1020;// level 0
assign po0066 = pi1015;// level 0
assign po0067 = pi1701;// level 0
assign po0068 = pi1747;// level 0
assign po0069 = pi0047;// level 0
assign po0070 = pi0975;// level 0
assign po0071 = pi0900;// level 0
assign po0072 = ~w134;// level 2
assign po0073 = pi1707;// level 0
assign po0074 = one;// level 0
assign po0075 = ~w139;// level 8
assign po0076 = pi0085;// level 0
assign po0077 = pi0072;// level 0
assign po0078 = pi0084;// level 0
assign po0079 = pi0087;// level 0
assign po0080 = pi0021;// level 0
assign po0081 = pi0020;// level 0
assign po0082 = pi0002;// level 0
assign po0083 = pi0000;// level 0
assign po0084 = pi0017;// level 0
assign po0085 = pi0026;// level 0
assign po0086 = pi0003;// level 0
assign po0087 = pi0001;// level 0
assign po0088 = pi0985;// level 0
assign po0089 = pi0976;// level 0
assign po0090 = pi1708;// level 0
assign po0091 = pi1715;// level 0
assign po0092 = pi1710;// level 0
assign po0093 = pi1706;// level 0
assign po0094 = ~w142;// level 10
assign po0095 = ~w145;// level 10
assign po0096 = ~w148;// level 10
assign po0097 = ~w151;// level 10
assign po0098 = ~w154;// level 10
assign po0099 = ~w157;// level 10
assign po0100 = ~w160;// level 10
assign po0101 = ~w163;// level 10
assign po0102 = ~w166;// level 10
assign po0103 = ~w169;// level 10
assign po0104 = ~w172;// level 10
assign po0105 = ~w175;// level 10
assign po0106 = ~w178;// level 10
assign po0107 = ~w181;// level 10
assign po0108 = ~w184;// level 10
assign po0109 = pi1752;// level 0
assign po0110 = ~w268;// level 11
assign po0111 = ~w296;// level 12
assign po0112 = ~w323;// level 11
assign po0113 = ~w348;// level 12
assign po0114 = ~w387;// level 8
assign po0115 = ~w391;// level 6
assign po0116 = ~w403;// level 6
assign po0117 = ~w512;// level 14
assign po0118 = ~w516;// level 6
assign po0119 = ~w637;// level 19
assign po0120 = ~w639;// level 19
assign po0121 = w653;// level 15
assign po0122 = ~w656;// level 3
assign po0123 = ~w661;// level 19
assign po0124 = w668;// level 15
assign po0125 = w675;// level 15
assign po0126 = w685;// level 15
assign po0127 = ~w693;// level 12
assign po0128 = w698;// level 15
assign po0129 = ~w706;// level 15
assign po0130 = ~w713;// level 11
assign po0131 = ~w719;// level 11
assign po0132 = ~w726;// level 16
assign po0133 = w732;// level 14
assign po0134 = w771;// level 7
assign po0135 = ~w777;// level 17
assign po0136 = ~w784;// level 12
assign po0137 = ~w791;// level 16
assign po0138 = ~w798;// level 15
assign po0139 = w809;// level 4
assign po0140 = w814;// level 15
assign po0141 = ~w920;// level 14
assign po0142 = ~w924;// level 14
assign po0143 = ~w931;// level 14
assign po0144 = one;// level 0
assign po0145 = ~w935;// level 14
assign po0146 = ~w939;// level 14
assign po0147 = ~w943;// level 14
assign po0148 = ~w947;// level 14
assign po0149 = ~w951;// level 14
assign po0150 = ~w955;// level 14
assign po0151 = ~w959;// level 14
assign po0152 = ~w963;// level 14
assign po0153 = ~w967;// level 14
assign po0154 = ~w973;// level 14
assign po0155 = ~w977;// level 14
assign po0156 = ~w981;// level 14
assign po0157 = ~w989;// level 13
assign po0158 = w999;// level 7
assign po0159 = ~w1005;// level 15
assign po0160 = w1014;// level 12
assign po0161 = ~w1020;// level 15
assign po0162 = ~w1023;// level 15
assign po0163 = ~w1029;// level 15
assign po0164 = ~w1035;// level 15
assign po0165 = ~w1041;// level 15
assign po0166 = w1045;// level 6
assign po0167 = ~w1053;// level 11
assign po0168 = ~w1069;// level 9
assign po0169 = pi0062;// level 0
assign po0170 = ~w1073;// level 5
assign po0171 = ~w1076;// level 15
assign po0172 = w1078;// level 4
assign po0173 = ~w991;// level 5
assign po0174 = w1079;// level 1
assign po0175 = ~w1087;// level 8
assign po0176 = w1090;// level 3
assign po0177 = w1096;// level 6
assign po0178 = ~w1263;// level 13
assign po0179 = ~w186;// level 2
assign po0180 = w1308;// level 10
assign po0181 = ~w1314;// level 10
assign po0182 = w1403;// level 15
assign po0183 = pi1746;// level 0
assign po0184 = w1411;// level 5
assign po0185 = w1420;// level 15
assign po0186 = ~w1424;// level 10
assign po0187 = ~w1429;// level 10
assign po0188 = w1437;// level 15
assign po0189 = w1445;// level 15
assign po0190 = w1453;// level 15
assign po0191 = w1461;// level 15
assign po0192 = w1469;// level 15
assign po0193 = w1477;// level 15
assign po0194 = w1484;// level 15
assign po0195 = w1491;// level 11
assign po0196 = w1499;// level 5
assign po0197 = w1507;// level 5
assign po0198 = w1584;// level 16
assign po0199 = w1592;// level 5
assign po0200 = w1595;// level 13
assign po0201 = ~w1601;// level 13
assign po0202 = w1678;// level 19
assign po0203 = ~w1686;// level 19
assign po0204 = ~w1692;// level 13
assign po0205 = ~w1693;// level 8
assign po0206 = w1704;// level 9
assign po0207 = w1721;// level 13
assign po0208 = w1596;// level 8
assign po0209 = ~w1723;// level 15
assign po0210 = ~w1725;// level 15
assign po0211 = ~w1727;// level 15
assign po0212 = ~w1729;// level 11
assign po0213 = w1735;// level 16
assign po0214 = ~w1738;// level 15
assign po0215 = ~w1741;// level 15
assign po0216 = ~w1743;// level 15
assign po0217 = ~w1745;// level 15
assign po0218 = ~w1747;// level 15
assign po0219 = w1751;// level 13
assign po0220 = w1754;// level 13
assign po0221 = w1757;// level 13
assign po0222 = w1758;// level 13
assign po0223 = w1761;// level 13
assign po0224 = w1768;// level 18
assign po0225 = w1772;// level 3
assign po0226 = w1776;// level 3
assign po0227 = w1780;// level 3
assign po0228 = ~w1782;// level 15
assign po0229 = w1786;// level 3
assign po0230 = ~w1788;// level 9
assign po0231 = w1793;// level 14
assign po0232 = w1265;// level 8
assign po0233 = w1795;// level 17
assign po0234 = ~one;// level 0
assign po0235 = ~w1798;// level 2
assign po0236 = ~w1872;// level 10
assign po0237 = ~one;// level 0
assign po0238 = ~one;// level 0
assign po0239 = w1875;// level 3
assign po0240 = w1878;// level 3
assign po0241 = w1881;// level 3
assign po0242 = w1884;// level 3
assign po0243 = ~w1472;// level 13
assign po0244 = ~w1464;// level 13
assign po0245 = ~w1480;// level 13
assign po0246 = ~w1487;// level 10
assign po0247 = w1887;// level 2
assign po0248 = w1926;// level 7
assign po0249 = ~w1930;// level 13
assign po0250 = w1932;// level 13
assign po0251 = w1937;// level 13
assign po0252 = w1940;// level 2
assign po0253 = ~w1979;// level 8
assign po0254 = w2018;// level 8
assign po0255 = w2021;// level 2
assign po0256 = w2024;// level 2
assign po0257 = w2027;// level 2
assign po0258 = w2030;// level 2
assign po0259 = ~w1432;// level 13
assign po0260 = ~w1448;// level 13
assign po0261 = ~w1440;// level 13
assign po0262 = ~w1456;// level 13
assign po0263 = ~w2035;// level 6
assign po0264 = w2043;// level 4
assign po0265 = ~w2046;// level 2
assign po0266 = ~w2049;// level 2
assign po0267 = w2052;// level 2
assign po0268 = w2055;// level 2
assign po0269 = w2058;// level 2
assign po0270 = w2061;// level 2
assign po0271 = w2064;// level 2
assign po0272 = w2067;// level 2
assign po0273 = w2070;// level 2
assign po0274 = w2073;// level 2
assign po0275 = w2076;// level 2
assign po0276 = w2079;// level 2
assign po0277 = w2082;// level 2
assign po0278 = w2085;// level 2
assign po0279 = w2088;// level 2
assign po0280 = w2091;// level 2
assign po0281 = w2094;// level 2
assign po0282 = w2097;// level 2
assign po0283 = w2100;// level 2
assign po0284 = w2103;// level 2
assign po0285 = w2106;// level 2
assign po0286 = w2109;// level 2
assign po0287 = w2112;// level 2
assign po0288 = w2115;// level 2
assign po0289 = w2118;// level 2
assign po0290 = w2121;// level 2
assign po0291 = w2124;// level 2
assign po0292 = w2127;// level 2
assign po0293 = w2130;// level 2
assign po0294 = w2192;// level 10
assign po0295 = w2231;// level 8
assign po0296 = w2236;// level 5
assign po0297 = w2239;// level 4
assign po0298 = ~w1414;// level 13
assign po0299 = ~w1394;// level 13
assign po0300 = w1283;// level 8
assign po0301 = ~one;// level 0
assign po0302 = ~one;// level 0
assign po0303 = ~one;// level 0
assign po0304 = ~w2242;// level 6
assign po0305 = w2243;// level 1
assign po0306 = w2246;// level 4
assign po0307 = w2247;// level 1
assign po0308 = ~w2253;// level 4
assign po0309 = w2261;// level 5
assign po0310 = ~w2264;// level 6
assign po0311 = w2267;// level 16
assign po0312 = ~w2271;// level 4
assign po0313 = ~w2275;// level 4
assign po0314 = ~w2279;// level 4
assign po0315 = ~w2283;// level 4
assign po0316 = ~w2287;// level 4
assign po0317 = ~w2294;// level 4
assign po0318 = ~w2298;// level 4
assign po0319 = ~w2305;// level 4
assign po0320 = ~w2309;// level 4
assign po0321 = ~w2313;// level 4
assign po0322 = ~w2317;// level 4
assign po0323 = ~w2321;// level 4
assign po0324 = ~w2325;// level 4
assign po0325 = ~w2329;// level 4
assign po0326 = ~w2333;// level 12
assign po0327 = w2335;// level 13
assign po0328 = ~w2339;// level 4
assign po0329 = ~w2343;// level 15
assign po0330 = ~w2347;// level 4
assign po0331 = ~w2351;// level 4
assign po0332 = w2359;// level 5
assign po0333 = pi0267;// level 0
assign po0334 = ~w2362;// level 2
assign po0335 = w2366;// level 5
assign po0336 = ~w2370;// level 4
assign po0337 = ~w2374;// level 4
assign po0338 = ~w2378;// level 4
assign po0339 = ~w2382;// level 4
assign po0340 = ~w2389;// level 4
assign po0341 = ~w2393;// level 4
assign po0342 = ~w2397;// level 4
assign po0343 = ~w2401;// level 4
assign po0344 = ~w2405;// level 4
assign po0345 = ~w2409;// level 4
assign po0346 = ~w2413;// level 4
assign po0347 = w2417;// level 6
assign po0348 = w2420;// level 4
assign po0349 = w2423;// level 4
assign po0350 = w2426;// level 4
assign po0351 = w2429;// level 5
assign po0352 = w2432;// level 5
assign po0353 = w2435;// level 6
assign po0354 = w2438;// level 6
assign po0355 = w2475;// level 12
assign po0356 = w2480;// level 14
assign po0357 = ~w2484;// level 4
assign po0358 = ~w2488;// level 4
assign po0359 = ~w2492;// level 4
assign po0360 = ~w2525;// level 7
assign po0361 = ~w2529;// level 3
assign po0362 = ~w2532;// level 3
assign po0363 = ~w2535;// level 3
assign po0364 = ~w2538;// level 3
assign po0365 = ~w2541;// level 2
assign po0366 = ~w2544;// level 3
assign po0367 = w2546;// level 2
assign po0368 = w2549;// level 3
assign po0369 = w2560;// level 7
assign po0370 = w2564;// level 6
assign po0371 = w2567;// level 10
assign po0372 = ~w2568;// level 3
assign po0373 = w2574;// level 10
assign po0374 = ~w2577;// level 3
assign po0375 = ~w2610;// level 7
assign po0376 = ~w2643;// level 7
assign po0377 = ~w2676;// level 7
assign po0378 = w2679;// level 13
assign po0379 = w2684;// level 3
assign po0380 = ~w2687;// level 3
assign po0381 = ~w2690;// level 3
assign po0382 = ~w2693;// level 3
assign po0383 = ~w2696;// level 3
assign po0384 = ~w2699;// level 3
assign po0385 = w2703;// level 4
assign po0386 = w2707;// level 4
assign po0387 = w2713;// level 10
assign po0388 = w2716;// level 10
assign po0389 = w2721;// level 10
assign po0390 = w2726;// level 15
assign po0391 = w2730;// level 16
assign po0392 = w2735;// level 12
assign po0393 = w2745;// level 10
assign po0394 = w2754;// level 10
assign po0395 = w2758;// level 5
assign po0396 = w2761;// level 2
assign po0397 = w2764;// level 10
assign po0398 = w2767;// level 10
assign po0399 = w2770;// level 10
assign po0400 = w2773;// level 10
assign po0401 = w2776;// level 10
assign po0402 = w2780;// level 10
assign po0403 = w2784;// level 10
assign po0404 = w2785;// level 10
assign po0405 = w2789;// level 10
assign po0406 = w2794;// level 10
assign po0407 = w2798;// level 10
assign po0408 = w2802;// level 10
assign po0409 = ~w2805;// level 2
assign po0410 = w2808;// level 10
assign po0411 = w2811;// level 10
assign po0412 = w2814;// level 10
assign po0413 = w2817;// level 10
assign po0414 = w2822;// level 10
assign po0415 = w2826;// level 10
assign po0416 = w2829;// level 10
assign po0417 = w2832;// level 10
assign po0418 = w2836;// level 10
assign po0419 = ~w2858;// level 9
assign po0420 = ~w2861;// level 2
assign po0421 = ~w2882;// level 9
assign po0422 = ~w2890;// level 9
assign po0423 = ~w2898;// level 9
assign po0424 = ~w2906;// level 9
assign po0425 = ~w2914;// level 9
assign po0426 = ~w2922;// level 9
assign po0427 = ~w2930;// level 9
assign po0428 = ~w2942;// level 8
assign po0429 = ~w2950;// level 9
assign po0430 = ~w2958;// level 9
assign po0431 = ~w2966;// level 9
assign po0432 = ~w2972;// level 8
assign po0433 = ~w2978;// level 8
assign po0434 = ~w2986;// level 9
assign po0435 = ~w2992;// level 8
assign po0436 = ~w2998;// level 8
assign po0437 = ~w3004;// level 8
assign po0438 = ~w3010;// level 8
assign po0439 = ~w3016;// level 8
assign po0440 = ~w3022;// level 8
assign po0441 = w3023;// level 3
assign po0442 = ~w3026;// level 2
assign po0443 = w3029;// level 13
assign po0444 = ~w3035;// level 8
assign po0445 = ~w3041;// level 8
assign po0446 = w3044;// level 6
assign po0447 = ~w3052;// level 9
assign po0448 = ~w3060;// level 9
assign po0449 = ~w3068;// level 9
assign po0450 = ~w3076;// level 9
assign po0451 = ~w3084;// level 9
assign po0452 = ~w3092;// level 9
assign po0453 = ~w3100;// level 9
assign po0454 = ~w3108;// level 9
assign po0455 = ~w3116;// level 9
assign po0456 = ~w3124;// level 9
assign po0457 = ~w3132;// level 9
assign po0458 = ~w3140;// level 9
assign po0459 = ~w3148;// level 9
assign po0460 = ~w3162;// level 9
assign po0461 = ~w3170;// level 9
assign po0462 = w1205;// level 12
assign po0463 = w3175;// level 14
assign po0464 = pi0434;// level 0
assign po0465 = w3179;// level 13
assign po0466 = ~w3187;// level 9
assign po0467 = ~w3197;// level 8
assign po0468 = ~w3253;// level 9
assign po0469 = ~w3310;// level 16
assign po0470 = ~w3316;// level 8
assign po0471 = w3320;// level 9
assign po0472 = ~w3328;// level 9
assign po0473 = ~w3336;// level 9
assign po0474 = ~w3344;// level 9
assign po0475 = ~w3352;// level 9
assign po0476 = ~w3358;// level 8
assign po0477 = ~w3366;// level 9
assign po0478 = ~w3374;// level 9
assign po0479 = ~w3380;// level 8
assign po0480 = ~w3386;// level 8
assign po0481 = ~w3394;// level 9
assign po0482 = ~w3400;// level 8
assign po0483 = ~w3406;// level 8
assign po0484 = ~w3412;// level 8
assign po0485 = ~w3418;// level 8
assign po0486 = ~w3424;// level 8
assign po0487 = ~w3430;// level 8
assign po0488 = ~w3436;// level 8
assign po0489 = ~w3490;// level 13
assign po0490 = w3543;// level 14
assign po0491 = ~w3558;// level 14
assign po0492 = w3578;// level 7
assign po0493 = w3648;// level 17
assign po0494 = ~w3655;// level 17
assign po0495 = ~w3664;// level 10
assign po0496 = w3672;// level 12
assign po0497 = ~w3686;// level 10
assign po0498 = w3697;// level 13
assign po0499 = ~w3703;// level 8
assign po0500 = ~w3709;// level 8
assign po0501 = ~w3715;// level 8
assign po0502 = ~w3721;// level 8
assign po0503 = ~w3727;// level 8
assign po0504 = ~w3733;// level 8
assign po0505 = ~w3739;// level 8
assign po0506 = ~w3745;// level 8
assign po0507 = ~w3751;// level 8
assign po0508 = ~w3757;// level 8
assign po0509 = ~w3763;// level 8
assign po0510 = ~w3769;// level 8
assign po0511 = ~w3775;// level 8
assign po0512 = ~w3781;// level 8
assign po0513 = ~w3787;// level 8
assign po0514 = ~w3793;// level 8
assign po0515 = ~w3799;// level 8
assign po0516 = ~w3805;// level 8
assign po0517 = ~w3811;// level 8
assign po0518 = w3815;// level 5
assign po0519 = ~w3819;// level 6
assign po0520 = w3823;// level 5
assign po0521 = ~w3832;// level 6
assign po0522 = w3837;// level 7
assign po0523 = ~w3847;// level 8
assign po0524 = ~w3855;// level 9
assign po0525 = ~w3863;// level 9
assign po0526 = ~w3871;// level 9
assign po0527 = ~w3879;// level 9
assign po0528 = ~w3887;// level 9
assign po0529 = ~w3895;// level 9
assign po0530 = ~w3903;// level 9
assign po0531 = ~w3911;// level 9
assign po0532 = ~w3919;// level 9
assign po0533 = ~w3927;// level 9
assign po0534 = ~w3935;// level 9
assign po0535 = ~w3943;// level 9
assign po0536 = ~w3951;// level 9
assign po0537 = ~w3965;// level 9
assign po0538 = ~w3973;// level 9
assign po0539 = w4018;// level 13
assign po0540 = ~w4024;// level 8
assign po0541 = ~w4026;// level 13
assign po0542 = ~w4034;// level 9
assign po0543 = w4039;// level 4
assign po0544 = pi0630;// level 0
assign po0545 = ~w4047;// level 9
assign po0546 = ~w4055;// level 9
assign po0547 = ~w4068;// level 9
assign po0548 = ~w4076;// level 9
assign po0549 = ~w4084;// level 9
assign po0550 = ~w4090;// level 8
assign po0551 = w4099;// level 17
assign po0552 = w4106;// level 9
assign po0553 = ~w4112;// level 8
assign po0554 = ~w4120;// level 9
assign po0555 = ~w4126;// level 8
assign po0556 = ~w4132;// level 8
assign po0557 = ~w4140;// level 9
assign po0558 = w4145;// level 5
assign po0559 = ~w4153;// level 9
assign po0560 = ~w4161;// level 9
assign po0561 = ~w4169;// level 9
assign po0562 = ~w4177;// level 9
assign po0563 = ~w4185;// level 9
assign po0564 = ~w4195;// level 8
assign po0565 = ~w4203;// level 9
assign po0566 = ~w4209;// level 8
assign po0567 = ~w4215;// level 8
assign po0568 = ~w4223;// level 9
assign po0569 = ~w4231;// level 9
assign po0570 = ~w4237;// level 8
assign po0571 = ~w4243;// level 8
assign po0572 = ~w4249;// level 8
assign po0573 = ~w4255;// level 8
assign po0574 = ~w4261;// level 8
assign po0575 = w4266;// level 6
assign po0576 = ~w4276;// level 13
assign po0577 = w4279;// level 5
assign po0578 = w4290;// level 13
assign po0579 = w4293;// level 3
assign po0580 = ~w4296;// level 13
assign po0581 = ~w4354;// level 17
assign po0582 = w4363;// level 16
assign po0583 = w4366;// level 6
assign po0584 = w4369;// level 3
assign po0585 = w4372;// level 4
assign po0586 = w4375;// level 5
assign po0587 = w4378;// level 5
assign po0588 = w4381;// level 6
assign po0589 = w4384;// level 6
assign po0590 = ~w4394;// level 10
assign po0591 = ~w4399;// level 17
assign po0592 = w4405;// level 15
assign po0593 = ~w4419;// level 13
assign po0594 = ~w4424;// level 10
assign po0595 = ~w4432;// level 12
assign po0596 = w4439;// level 13
assign po0597 = ~w4445;// level 8
assign po0598 = ~w4451;// level 8
assign po0599 = ~w4457;// level 8
assign po0600 = ~w4463;// level 8
assign po0601 = ~w4469;// level 8
assign po0602 = ~w4475;// level 8
assign po0603 = ~w4481;// level 8
assign po0604 = ~w4487;// level 8
assign po0605 = ~w4493;// level 8
assign po0606 = ~w4499;// level 8
assign po0607 = ~w4505;// level 8
assign po0608 = ~w4511;// level 8
assign po0609 = ~w4517;// level 8
assign po0610 = ~w4523;// level 8
assign po0611 = ~w4529;// level 8
assign po0612 = ~w4535;// level 8
assign po0613 = ~w4541;// level 8
assign po0614 = ~w4547;// level 8
assign po0615 = ~w4553;// level 8
assign po0616 = w4557;// level 5
assign po0617 = ~w4567;// level 6
assign po0618 = ~w4574;// level 7
assign po0619 = w4581;// level 9
assign po0620 = w4587;// level 11
assign po0621 = w4591;// level 5
assign po0622 = ~w4602;// level 6
assign po0623 = w4608;// level 7
assign po0624 = ~w4617;// level 8
assign po0625 = ~w4625;// level 9
assign po0626 = ~w4633;// level 9
assign po0627 = ~w4641;// level 9
assign po0628 = ~w4649;// level 9
assign po0629 = ~w4657;// level 9
assign po0630 = ~w4665;// level 9
assign po0631 = ~w4673;// level 9
assign po0632 = ~w4681;// level 9
assign po0633 = ~w4689;// level 9
assign po0634 = ~w4697;// level 9
assign po0635 = ~w4705;// level 9
assign po0636 = ~w4713;// level 9
assign po0637 = ~w4721;// level 9
assign po0638 = ~w4729;// level 9
assign po0639 = ~w4737;// level 9
assign po0640 = ~w4745;// level 9
assign po0641 = ~w4753;// level 9
assign po0642 = ~w4759;// level 8
assign po0643 = w4769;// level 14
assign po0644 = ~w4777;// level 9
assign po0645 = w4780;// level 8
assign po0646 = ~w4788;// level 9
assign po0647 = ~w4794;// level 8
assign po0648 = ~w4800;// level 8
assign po0649 = ~w4806;// level 8
assign po0650 = ~w4812;// level 8
assign po0651 = w4819;// level 10
assign po0652 = ~w4827;// level 9
assign po0653 = ~w4833;// level 8
assign po0654 = ~w4841;// level 9
assign po0655 = w4845;// level 12
assign po0656 = ~w4853;// level 9
assign po0657 = ~w4861;// level 9
assign po0658 = ~w4869;// level 9
assign po0659 = w4875;// level 12
assign po0660 = ~w4883;// level 9
assign po0661 = ~w4891;// level 9
assign po0662 = ~w4943;// level 16
assign po0663 = ~w4951;// level 9
assign po0664 = ~w4959;// level 9
assign po0665 = ~w4967;// level 9
assign po0666 = ~w4975;// level 9
assign po0667 = ~w4983;// level 9
assign po0668 = ~w4991;// level 9
assign po0669 = ~w4999;// level 9
assign po0670 = w5009;// level 16
assign po0671 = w5012;// level 2
assign po0672 = ~w5017;// level 13
assign po0673 = ~w5029;// level 17
assign po0674 = ~w5037;// level 16
assign po0675 = ~w5047;// level 16
assign po0676 = ~w5054;// level 10
assign po0677 = ~w5063;// level 10
assign po0678 = w5071;// level 14
assign po0679 = w5077;// level 9
assign po0680 = ~w5083;// level 8
assign po0681 = ~w5089;// level 8
assign po0682 = ~w5095;// level 8
assign po0683 = ~w5101;// level 8
assign po0684 = ~w5107;// level 8
assign po0685 = ~w5113;// level 8
assign po0686 = ~w5119;// level 8
assign po0687 = ~w5125;// level 8
assign po0688 = ~w5131;// level 8
assign po0689 = ~w5137;// level 8
assign po0690 = ~w5143;// level 8
assign po0691 = ~w5149;// level 8
assign po0692 = ~w5155;// level 8
assign po0693 = ~w5161;// level 8
assign po0694 = ~w5167;// level 8
assign po0695 = ~w5173;// level 8
assign po0696 = w5177;// level 5
assign po0697 = ~w5185;// level 7
assign po0698 = w5191;// level 12
assign po0699 = ~w5200;// level 7
assign po0700 = w5205;// level 7
assign po0701 = ~w5212;// level 8
assign po0702 = w5215;// level 8
assign po0703 = ~w5223;// level 9
assign po0704 = w5227;// level 5
assign po0705 = ~w5235;// level 9
assign po0706 = ~w5243;// level 9
assign po0707 = ~w5251;// level 9
assign po0708 = ~w5259;// level 9
assign po0709 = ~w5267;// level 9
assign po0710 = ~w5275;// level 9
assign po0711 = ~w5283;// level 9
assign po0712 = ~w5291;// level 9
assign po0713 = ~w5299;// level 9
assign po0714 = ~w5307;// level 9
assign po0715 = ~w5315;// level 9
assign po0716 = ~w5323;// level 9
assign po0717 = ~w5331;// level 9
assign po0718 = ~w5339;// level 9
assign po0719 = ~w5347;// level 9
assign po0720 = ~w5355;// level 9
assign po0721 = ~w5363;// level 9
assign po0722 = ~w5371;// level 9
assign po0723 = ~w5379;// level 9
assign po0724 = ~w5387;// level 9
assign po0725 = w5390;// level 8
assign po0726 = ~w5398;// level 9
assign po0727 = w5401;// level 8
assign po0728 = w5412;// level 6
assign po0729 = ~w5417;// level 5
assign po0730 = w5420;// level 12
assign po0731 = ~w5428;// level 9
assign po0732 = w5434;// level 9
assign po0733 = ~w5441;// level 10
assign po0734 = ~w5451;// level 8
assign po0735 = ~w5460;// level 4
assign po0736 = ~w5468;// level 9
assign po0737 = w5474;// level 10
assign po0738 = ~w5480;// level 8
assign po0739 = ~w5488;// level 9
assign po0740 = ~w5491;// level 7
assign po0741 = ~w5498;// level 16
assign po0742 = ~w5506;// level 9
assign po0743 = ~w5512;// level 8
assign po0744 = w5515;// level 3
assign po0745 = ~w5521;// level 8
assign po0746 = ~w5527;// level 8
assign po0747 = ~w5533;// level 8
assign po0748 = ~w5539;// level 8
assign po0749 = ~w5545;// level 8
assign po0750 = ~w5553;// level 9
assign po0751 = ~w5559;// level 8
assign po0752 = w5567;// level 16
assign po0753 = w5570;// level 2
assign po0754 = w5572;// level 2
assign po0755 = ~w5580;// level 9
assign po0756 = w5582;// level 8
assign po0757 = w5587;// level 7
assign po0758 = ~w5594;// level 9
assign po0759 = w5604;// level 17
assign po0760 = ~w5611;// level 8
assign po0761 = ~w5617;// level 8
assign po0762 = ~w5623;// level 8
assign po0763 = ~w5632;// level 7
assign po0764 = ~w5639;// level 7
assign po0765 = w5644;// level 12
assign po0766 = ~w5652;// level 9
assign po0767 = ~w5660;// level 9
assign po0768 = ~w5668;// level 9
assign po0769 = ~w5676;// level 9
assign po0770 = w5680;// level 7
assign po0771 = w5683;// level 2
assign po0772 = ~w5692;// level 6
assign po0773 = ~w5757;// level 18
assign po0774 = w5774;// level 16
assign po0775 = ~w5780;// level 15
assign po0776 = w5783;// level 2
assign po0777 = ~w5789;// level 8
assign po0778 = ~w5795;// level 8
assign po0779 = w5806;// level 10
assign po0780 = ~w5812;// level 8
assign po0781 = ~w5818;// level 8
assign po0782 = w5857;// level 7
assign po0783 = w5859;// level 10
assign po0784 = ~w5874;// level 18
assign po0785 = w5885;// level 13
assign po0786 = w5933;// level 8
assign po0787 = w5936;// level 8
assign po0788 = ~w5942;// level 12
assign po0789 = ~w5953;// level 15
assign po0790 = ~w5959;// level 8
assign po0791 = ~w5965;// level 8
assign po0792 = ~w5971;// level 8
assign po0793 = ~w5977;// level 8
assign po0794 = ~w5983;// level 8
assign po0795 = ~w5989;// level 8
assign po0796 = ~w5995;// level 8
assign po0797 = ~w6001;// level 8
assign po0798 = ~w6007;// level 8
assign po0799 = ~w6013;// level 8
assign po0800 = ~w6019;// level 8
assign po0801 = ~w6025;// level 8
assign po0802 = ~w6031;// level 8
assign po0803 = ~w6037;// level 8
assign po0804 = ~w6043;// level 8
assign po0805 = ~w3577;// level 6
assign po0806 = ~w6050;// level 8
assign po0807 = w6054;// level 5
assign po0808 = ~w6063;// level 6
assign po0809 = w6070;// level 7
assign po0810 = w6074;// level 5
assign po0811 = w6076;// level 7
assign po0812 = ~w6080;// level 8
assign po0813 = ~w6086;// level 8
assign po0814 = ~w6092;// level 8
assign po0815 = w3975;// level 12
assign po0816 = w6100;// level 12
assign po0817 = ~w6110;// level 8
assign po0818 = ~w6121;// level 18
assign po0819 = ~w6129;// level 11
assign po0820 = w6180;// level 8
assign po0821 = w6189;// level 16
assign po0822 = w6246;// level 8
assign po0823 = w6254;// level 11
assign po0824 = w6261;// level 18
assign po0825 = ~w6264;// level 8
assign po0826 = ~w6273;// level 10
assign po0827 = ~w6284;// level 6
assign po0828 = ~w6292;// level 8
assign po0829 = w6301;// level 17
assign po0830 = w6347;// level 9
assign po0831 = ~w6391;// level 10
assign po0832 = ~w6395;// level 7
assign po0833 = w6414;// level 7
assign po0834 = w6456;// level 8
assign po0835 = w6460;// level 9
assign po0836 = ~w6476;// level 14
assign po0837 = w6479;// level 3
assign po0838 = ~w6483;// level 12
assign po0839 = ~w6487;// level 7
assign po0840 = ~w6491;// level 7
assign po0841 = ~w6495;// level 7
assign po0842 = ~w6501;// level 8
assign po0843 = ~w6508;// level 7
assign po0844 = ~w6512;// level 7
assign po0845 = ~w6516;// level 7
assign po0846 = ~w6526;// level 8
assign po0847 = ~w6533;// level 7
assign po0848 = pi1012;// level 0
assign po0849 = pi1001;// level 0
assign po0850 = pi1005;// level 0
assign po0851 = pi1006;// level 0
assign po0852 = w6537;// level 8
assign po0853 = ~w6541;// level 7
assign po0854 = ~w6548;// level 7
assign po0855 = ~w6555;// level 8
assign po0856 = ~w6558;// level 7
assign po0857 = ~w6567;// level 10
assign po0858 = ~w6576;// level 10
assign po0859 = ~w6585;// level 10
assign po0860 = ~w6594;// level 10
assign po0861 = ~w6603;// level 10
assign po0862 = ~w6663;// level 9
assign po0863 = ~w6672;// level 10
assign po0864 = ~w6681;// level 10
assign po0865 = ~w6690;// level 10
assign po0866 = ~w6699;// level 10
assign po0867 = ~w6708;// level 10
assign po0868 = ~w6717;// level 10
assign po0869 = w6727;// level 7
assign po0870 = ~w6733;// level 9
assign po0871 = ~w6742;// level 10
assign po0872 = w6748;// level 8
assign po0873 = ~w6751;// level 8
assign po0874 = ~w6754;// level 8
assign po0875 = ~w6757;// level 8
assign po0876 = ~w6766;// level 10
assign po0877 = ~w6775;// level 10
assign po0878 = w6778;// level 2
assign po0879 = ~w6787;// level 10
assign po0880 = ~w6796;// level 10
assign po0881 = ~w6805;// level 10
assign po0882 = w6818;// level 8
assign po0883 = ~pi1000;// level 0
assign po0884 = ~pi1004;// level 0
assign po0885 = w6857;// level 7
assign po0886 = ~w6861;// level 8
assign po0887 = ~w6865;// level 9
assign po0888 = ~w6869;// level 9
assign po0889 = ~w6878;// level 10
assign po0890 = w6881;// level 2
assign po0891 = w6884;// level 2
assign po0892 = ~w6887;// level 9
assign po0893 = w6890;// level 2
assign po0894 = w6897;// level 7
assign po0895 = w6900;// level 3
assign po0896 = ~w6903;// level 9
assign po0897 = ~w6906;// level 9
assign po0898 = w6910;// level 8
assign po0899 = ~w6913;// level 9
assign po0900 = w6914;// level 8
assign po0901 = w6917;// level 8
assign po0902 = w6921;// level 8
assign po0903 = w6924;// level 2
assign po0904 = ~w6933;// level 10
assign po0905 = ~w6942;// level 10
assign po0906 = ~w6951;// level 10
assign po0907 = ~w6960;// level 10
assign po0908 = ~w6969;// level 10
assign po0909 = ~w6978;// level 10
assign po0910 = ~w6987;// level 10
assign po0911 = ~w6996;// level 10
assign po0912 = ~w7005;// level 10
assign po0913 = ~w7014;// level 10
assign po0914 = ~w7023;// level 10
assign po0915 = ~w7032;// level 10
assign po0916 = ~w7041;// level 10
assign po0917 = ~w7050;// level 10
assign po0918 = ~w7059;// level 10
assign po0919 = ~w7068;// level 10
assign po0920 = ~w7077;// level 10
assign po0921 = ~w7086;// level 10
assign po0922 = ~w7095;// level 10
assign po0923 = ~w7104;// level 10
assign po0924 = ~w7113;// level 10
assign po0925 = ~w7122;// level 10
assign po0926 = ~w7131;// level 10
assign po0927 = ~w7140;// level 10
assign po0928 = ~w7149;// level 10
assign po0929 = ~w7158;// level 10
assign po0930 = ~w7167;// level 10
assign po0931 = ~w7176;// level 10
assign po0932 = ~w7185;// level 10
assign po0933 = ~w7194;// level 10
assign po0934 = ~w7203;// level 10
assign po0935 = ~w7212;// level 10
assign po0936 = ~w7221;// level 10
assign po0937 = ~w7230;// level 10
assign po0938 = ~w7239;// level 10
assign po0939 = ~w7248;// level 10
assign po0940 = ~w7257;// level 10
assign po0941 = ~w7266;// level 10
assign po0942 = ~w7275;// level 10
assign po0943 = ~w7284;// level 10
assign po0944 = ~w7293;// level 10
assign po0945 = ~w7302;// level 10
assign po0946 = ~w7311;// level 10
assign po0947 = ~w7320;// level 10
assign po0948 = ~w7329;// level 10
assign po0949 = ~w7338;// level 10
assign po0950 = ~w7347;// level 10
assign po0951 = ~w7356;// level 10
assign po0952 = ~w7365;// level 10
assign po0953 = ~w7374;// level 10
assign po0954 = ~w7383;// level 10
assign po0955 = ~w7392;// level 10
assign po0956 = ~w7401;// level 10
assign po0957 = ~w7410;// level 10
assign po0958 = ~w7419;// level 10
assign po0959 = ~w7428;// level 10
assign po0960 = ~w7437;// level 10
assign po0961 = ~w7446;// level 10
assign po0962 = ~w7455;// level 10
assign po0963 = ~w7464;// level 10
assign po0964 = ~w7473;// level 10
assign po0965 = ~w7482;// level 10
assign po0966 = ~w7491;// level 10
assign po0967 = ~w7500;// level 10
assign po0968 = ~w7509;// level 10
assign po0969 = ~w7518;// level 10
assign po0970 = ~w7525;// level 4
assign po0971 = ~w7529;// level 4
assign po0972 = ~w7536;// level 4
assign po0973 = ~pi1013;// level 0
assign po0974 = ~pi1002;// level 0
assign po0975 = ~pi1003;// level 0
assign po0976 = ~pi1008;// level 0
assign po0977 = ~pi1009;// level 0
assign po0978 = ~pi1010;// level 0
assign po0979 = ~w7545;// level 10
assign po0980 = ~w7554;// level 10
assign po0981 = w7559;// level 7
assign po0982 = ~w7568;// level 10
assign po0983 = pi0974;// level 0
assign po0984 = ~pi1011;// level 0
assign po0985 = ~w7573;// level 4
assign po0986 = ~w7582;// level 10
assign po0987 = ~w7586;// level 9
assign po0988 = ~w7595;// level 10
assign po0989 = ~w7604;// level 10
assign po0990 = w7607;// level 7
assign po0991 = w7610;// level 2
assign po0992 = ~w7653;// level 9
assign po0993 = w7656;// level 7
assign po0994 = ~w7699;// level 9
assign po0995 = ~w7742;// level 9
assign po0996 = w7745;// level 7
assign po0997 = w7748;// level 2
assign po0998 = w7751;// level 7
assign po0999 = w7754;// level 7
assign po1000 = w7760;// level 8
assign po1001 = w7763;// level 8
assign po1002 = w7764;// level 12
assign po1003 = ~w7789;// level 11
assign po1004 = pi0997;// level 0
assign po1005 = w7803;// level 13
assign po1006 = w7818;// level 12
assign po1007 = w7831;// level 15
assign po1008 = w7843;// level 10
assign po1009 = w7858;// level 9
assign po1010 = w7861;// level 3
assign po1011 = w7864;// level 2
assign po1012 = w7867;// level 8
assign po1013 = w7870;// level 8
assign po1014 = w7873;// level 2
assign po1015 = w7876;// level 2
assign po1016 = w7879;// level 2
assign po1017 = w7882;// level 2
assign po1018 = w7885;// level 2
assign po1019 = w7888;// level 2
assign po1020 = w7891;// level 2
assign po1021 = w7894;// level 2
assign po1022 = w7897;// level 2
assign po1023 = w7900;// level 2
assign po1024 = w7903;// level 3
assign po1025 = w7916;// level 11
assign po1026 = w7919;// level 7
assign po1027 = w7922;// level 7
assign po1028 = w7930;// level 9
assign po1029 = w7933;// level 7
assign po1030 = w7937;// level 10
assign po1031 = w7940;// level 7
assign po1032 = w7942;// level 7
assign po1033 = w7945;// level 7
assign po1034 = w7948;// level 7
assign po1035 = w7951;// level 7
assign po1036 = w7954;// level 7
assign po1037 = w7957;// level 7
assign po1038 = w7960;// level 7
assign po1039 = w7963;// level 7
assign po1040 = w7966;// level 7
assign po1041 = w7969;// level 7
assign po1042 = w7972;// level 7
assign po1043 = w7975;// level 7
assign po1044 = w7978;// level 7
assign po1045 = w7981;// level 7
assign po1046 = w7983;// level 7
assign po1047 = ~w7988;// level 4
assign po1048 = ~w7993;// level 4
assign po1049 = pi0999;// level 0
assign po1050 = ~w7996;// level 4
assign po1051 = ~w7999;// level 4
assign po1052 = w8002;// level 7
assign po1053 = w8005;// level 7
assign po1054 = pi1007;// level 0
assign po1055 = pi0998;// level 0
assign po1056 = ~w8053;// level 18
assign po1057 = ~w8104;// level 18
assign po1058 = w8154;// level 18
assign po1059 = ~w8202;// level 18
assign po1060 = w8205;// level 2
assign po1061 = w8208;// level 2
assign po1062 = w8211;// level 2
assign po1063 = w8214;// level 8
assign po1064 = w8217;// level 2
assign po1065 = w8220;// level 2
assign po1066 = w8225;// level 8
assign po1067 = w8228;// level 8
assign po1068 = w8231;// level 8
assign po1069 = w8233;// level 7
assign po1070 = w8236;// level 2
assign po1071 = w8239;// level 2
assign po1072 = w8242;// level 9
assign po1073 = w8245;// level 2
assign po1074 = w8248;// level 3
assign po1075 = w8256;// level 9
assign po1076 = ~w8261;// level 4
assign po1077 = ~w8264;// level 4
assign po1078 = ~w8269;// level 4
assign po1079 = w8272;// level 8
assign po1080 = ~w8279;// level 8
assign po1081 = w8282;// level 2
assign po1082 = ~w8285;// level 4
assign po1083 = w8286;// level 6
assign po1084 = w8290;// level 11
assign po1085 = ~w8294;// level 9
assign po1086 = w8296;// level 2
assign po1087 = w8298;// level 16
assign po1088 = ~w8300;// level 17
assign po1089 = ~w8302;// level 16
assign po1090 = w8304;// level 16
assign po1091 = ~w8326;// level 8
assign po1092 = w8332;// level 12
assign po1093 = w8335;// level 8
assign po1094 = w8337;// level 8
assign po1095 = w8339;// level 2
assign po1096 = w8341;// level 2
assign po1097 = w8344;// level 2
assign po1098 = w8347;// level 2
assign po1099 = w8350;// level 3
assign po1100 = w8353;// level 8
assign po1101 = ~w8358;// level 4
assign po1102 = ~w8361;// level 4
assign po1103 = ~w8366;// level 4
assign po1104 = w8369;// level 8
assign po1105 = w8370;// level 5
assign po1106 = w8373;// level 6
assign po1107 = w8376;// level 6
assign po1108 = w8379;// level 6
assign po1109 = w8382;// level 6
assign po1110 = w8385;// level 6
assign po1111 = w8388;// level 6
assign po1112 = w8391;// level 6
assign po1113 = w8394;// level 6
assign po1114 = w8397;// level 6
assign po1115 = w8400;// level 6
assign po1116 = w8403;// level 6
assign po1117 = w8406;// level 6
assign po1118 = w8409;// level 6
assign po1119 = w8412;// level 6
assign po1120 = w8415;// level 6
assign po1121 = w8418;// level 6
assign po1122 = w8421;// level 6
assign po1123 = ~w8424;// level 4
assign po1124 = ~w8445;// level 5
assign po1125 = ~w8454;// level 6
assign po1126 = ~w8457;// level 6
assign po1127 = w8461;// level 9
assign po1128 = ~w8465;// level 8
assign po1129 = ~w8486;// level 5
assign po1130 = w8488;// level 6
assign po1131 = ~w8494;// level 8
assign po1132 = ~w8497;// level 8
assign po1133 = ~w8500;// level 8
assign po1134 = ~w8503;// level 8
assign po1135 = ~w8506;// level 8
assign po1136 = ~w8512;// level 8
assign po1137 = ~w8515;// level 8
assign po1138 = ~w8518;// level 8
assign po1139 = ~w8521;// level 8
assign po1140 = ~w8527;// level 8
assign po1141 = ~w8530;// level 8
assign po1142 = ~w8533;// level 8
assign po1143 = ~w8536;// level 8
assign po1144 = w8539;// level 8
assign po1145 = ~w8541;// level 7
assign po1146 = w8544;// level 8
assign po1147 = w8550;// level 9
assign po1148 = ~w8553;// level 6
assign po1149 = ~w8556;// level 6
assign po1150 = ~w8559;// level 6
assign po1151 = ~w8562;// level 6
assign po1152 = ~w8565;// level 6
assign po1153 = ~w8568;// level 6
assign po1154 = w8571;// level 8
assign po1155 = w8577;// level 7
assign po1156 = w8578;// level 5
assign po1157 = w8581;// level 3
assign po1158 = ~w8584;// level 6
assign po1159 = w8587;// level 8
assign po1160 = ~w8593;// level 8
assign po1161 = ~w8596;// level 8
assign po1162 = ~w8598;// level 7
assign po1163 = ~w8601;// level 8
assign po1164 = ~w8603;// level 7
assign po1165 = ~w8605;// level 7
assign po1166 = ~w8607;// level 7
assign po1167 = w8611;// level 6
assign po1168 = ~w8640;// level 9
assign po1169 = ~w8669;// level 9
assign po1170 = ~w8698;// level 9
assign po1171 = ~w8700;// level 7
assign po1172 = ~w8702;// level 7
assign po1173 = ~w8704;// level 7
assign po1174 = ~w8706;// level 7
assign po1175 = ~w8708;// level 7
assign po1176 = ~w8710;// level 7
assign po1177 = ~w8716;// level 8
assign po1178 = ~w8719;// level 8
assign po1179 = ~w8722;// level 8
assign po1180 = ~w8724;// level 7
assign po1181 = ~w8751;// level 8
assign po1182 = ~w8753;// level 7
assign po1183 = ~w8756;// level 8
assign po1184 = ~w8758;// level 7
assign po1185 = ~w8761;// level 8
assign po1186 = ~w8763;// level 7
assign po1187 = ~w8766;// level 8
assign po1188 = w8769;// level 6
assign po1189 = ~w8772;// level 8
assign po1190 = ~w8775;// level 8
assign po1191 = ~w8777;// level 7
assign po1192 = ~w8780;// level 8
assign po1193 = ~w8783;// level 8
assign po1194 = ~w8785;// level 7
assign po1195 = ~w8787;// level 7
assign po1196 = ~w8789;// level 7
assign po1197 = w8797;// level 8
assign po1198 = ~w8799;// level 7
assign po1199 = w8802;// level 8
assign po1200 = w8806;// level 8
assign po1201 = ~w8809;// level 8
assign po1202 = ~w8811;// level 7
assign po1203 = ~w8814;// level 8
assign po1204 = ~w8817;// level 8
assign po1205 = ~w8820;// level 8
assign po1206 = ~w8823;// level 8
assign po1207 = ~w8826;// level 8
assign po1208 = w8831;// level 8
assign po1209 = ~w8834;// level 8
assign po1210 = ~w17;// level 6
assign po1211 = ~w8837;// level 8
assign po1212 = ~w8840;// level 8
assign po1213 = ~w8843;// level 8
assign po1214 = ~w8846;// level 8
assign po1215 = ~w8849;// level 8
assign po1216 = ~w8852;// level 8
assign po1217 = ~w8855;// level 8
assign po1218 = ~w8858;// level 8
assign po1219 = ~w8861;// level 8
assign po1220 = ~w8864;// level 8
assign po1221 = ~w8867;// level 8
assign po1222 = ~w8870;// level 8
assign po1223 = ~w8873;// level 8
assign po1224 = ~w8876;// level 8
assign po1225 = ~w8879;// level 8
assign po1226 = ~w8882;// level 8
assign po1227 = ~w8885;// level 8
assign po1228 = ~w8888;// level 8
assign po1229 = ~w8891;// level 8
assign po1230 = ~w8894;// level 8
assign po1231 = ~w8897;// level 8
assign po1232 = ~w8900;// level 8
assign po1233 = ~w8903;// level 8
assign po1234 = ~w8906;// level 8
assign po1235 = ~w8909;// level 8
assign po1236 = ~w8912;// level 8
assign po1237 = ~w8915;// level 8
assign po1238 = ~w8918;// level 8
assign po1239 = ~w8921;// level 8
assign po1240 = ~w8924;// level 8
assign po1241 = ~w8927;// level 8
assign po1242 = ~w8930;// level 8
assign po1243 = ~w8933;// level 8
assign po1244 = ~w8936;// level 8
assign po1245 = ~w8939;// level 8
assign po1246 = ~w8942;// level 8
assign po1247 = ~w8945;// level 8
assign po1248 = ~w8948;// level 8
assign po1249 = ~w8951;// level 8
assign po1250 = ~w8954;// level 8
assign po1251 = ~w8957;// level 8
assign po1252 = ~w8960;// level 8
assign po1253 = ~w8963;// level 8
assign po1254 = ~w8966;// level 8
assign po1255 = ~w8969;// level 8
assign po1256 = ~w8972;// level 8
assign po1257 = ~w8975;// level 8
assign po1258 = ~w8977;// level 7
assign po1259 = ~w8979;// level 7
assign po1260 = ~w8981;// level 7
assign po1261 = ~w8983;// level 7
assign po1262 = ~w8985;// level 7
assign po1263 = ~w8987;// level 7
assign po1264 = ~w8989;// level 7
assign po1265 = ~w8991;// level 7
assign po1266 = ~w8993;// level 7
assign po1267 = ~w8995;// level 7
assign po1268 = ~w8997;// level 7
assign po1269 = ~w8999;// level 7
assign po1270 = ~w9001;// level 7
assign po1271 = ~w9003;// level 7
assign po1272 = ~w9005;// level 7
assign po1273 = ~w9010;// level 8
assign po1274 = w9013;// level 8
assign po1275 = ~w9015;// level 7
assign po1276 = ~w9017;// level 7
assign po1277 = ~w9019;// level 7
assign po1278 = ~w9021;// level 7
assign po1279 = ~w9023;// level 7
assign po1280 = ~w9025;// level 7
assign po1281 = ~w9027;// level 7
assign po1282 = ~w9029;// level 7
assign po1283 = ~w9031;// level 7
assign po1284 = ~w9033;// level 7
assign po1285 = ~w9035;// level 7
assign po1286 = ~w9037;// level 7
assign po1287 = ~w9039;// level 7
assign po1288 = ~w9041;// level 7
assign po1289 = ~w9043;// level 7
assign po1290 = ~w9045;// level 7
assign po1291 = ~w9047;// level 7
assign po1292 = ~w9049;// level 7
assign po1293 = ~w9054;// level 8
assign po1294 = ~w9056;// level 7
assign po1295 = ~w9058;// level 7
assign po1296 = ~w9060;// level 7
assign po1297 = ~w9062;// level 7
assign po1298 = ~w9064;// level 7
assign po1299 = ~w9066;// level 7
assign po1300 = ~w9068;// level 7
assign po1301 = ~w9070;// level 7
assign po1302 = ~w9072;// level 7
assign po1303 = ~w9074;// level 7
assign po1304 = ~w9076;// level 7
assign po1305 = ~w9078;// level 7
assign po1306 = ~w9080;// level 7
assign po1307 = ~w9082;// level 7
assign po1308 = ~w9084;// level 7
assign po1309 = ~w9086;// level 7
assign po1310 = ~w9088;// level 7
assign po1311 = ~w9090;// level 7
assign po1312 = ~w9092;// level 7
assign po1313 = ~w9094;// level 7
assign po1314 = ~w9096;// level 7
assign po1315 = ~w9101;// level 8
assign po1316 = ~w9103;// level 7
assign po1317 = ~w9105;// level 7
assign po1318 = ~w9107;// level 7
assign po1319 = ~w9109;// level 7
assign po1320 = ~w9111;// level 7
assign po1321 = ~w9113;// level 7
assign po1322 = ~w9115;// level 7
assign po1323 = ~w9117;// level 7
assign po1324 = ~w9119;// level 7
assign po1325 = ~w9121;// level 7
assign po1326 = ~w9123;// level 7
assign po1327 = ~w9125;// level 7
assign po1328 = ~w9127;// level 7
assign po1329 = ~w9129;// level 7
assign po1330 = ~w9131;// level 7
assign po1331 = ~w9133;// level 7
assign po1332 = ~w9135;// level 7
assign po1333 = ~w9137;// level 7
assign po1334 = ~w9142;// level 8
assign po1335 = w9145;// level 2
assign po1336 = ~w9148;// level 6
assign po1337 = ~w9151;// level 6
assign po1338 = ~w9154;// level 6
assign po1339 = w9157;// level 6
assign po1340 = w9160;// level 6
assign po1341 = ~w9162;// level 7
assign po1342 = ~w9165;// level 5
assign po1343 = ~w1860;// level 6
assign po1344 = ~w9168;// level 8
assign po1345 = ~w9171;// level 6
assign po1346 = ~w9174;// level 8
assign po1347 = ~w9176;// level 7
assign po1348 = ~w9178;// level 7
assign po1349 = ~w9180;// level 7
assign po1350 = ~w9182;// level 7
assign po1351 = ~w9185;// level 8
assign po1352 = ~w9188;// level 8
assign po1353 = ~w9190;// level 7
assign po1354 = ~w9192;// level 7
assign po1355 = ~w9194;// level 7
assign po1356 = ~w9196;// level 7
assign po1357 = ~w9198;// level 7
assign po1358 = ~w9200;// level 7
assign po1359 = pi1410;// level 0
assign po1360 = ~w9202;// level 7
assign po1361 = ~w9205;// level 8
assign po1362 = ~w9208;// level 8
assign po1363 = ~w9210;// level 7
assign po1364 = ~w9213;// level 8
assign po1365 = ~w9216;// level 8
assign po1366 = ~w9219;// level 8
assign po1367 = ~w9222;// level 8
assign po1368 = ~w9225;// level 8
assign po1369 = ~w9228;// level 8
assign po1370 = ~w9231;// level 8
assign po1371 = ~w9234;// level 8
assign po1372 = ~w9236;// level 7
assign po1373 = ~w9238;// level 7
assign po1374 = ~w9241;// level 8
assign po1375 = ~w9243;// level 7
assign po1376 = ~w9246;// level 8
assign po1377 = ~w9249;// level 8
assign po1378 = ~w9251;// level 7
assign po1379 = ~w9254;// level 8
assign po1380 = ~w9257;// level 8
assign po1381 = ~w9260;// level 8
assign po1382 = ~w9263;// level 8
assign po1383 = ~w9266;// level 8
assign po1384 = ~w9268;// level 7
assign po1385 = ~w9270;// level 7
assign po1386 = ~w9273;// level 8
assign po1387 = ~w9275;// level 7
assign po1388 = ~w9277;// level 7
assign po1389 = ~w9280;// level 8
assign po1390 = ~w9282;// level 7
assign po1391 = ~w9284;// level 7
assign po1392 = ~w9286;// level 7
assign po1393 = ~w9288;// level 7
assign po1394 = ~w9291;// level 5
assign po1395 = ~w9332;// level 9
assign po1396 = ~w9338;// level 8
assign po1397 = ~w9341;// level 8
assign po1398 = ~w9344;// level 8
assign po1399 = ~w9347;// level 8
assign po1400 = ~w9350;// level 8
assign po1401 = ~w9352;// level 7
assign po1402 = ~w9389;// level 9
assign po1403 = ~w9424;// level 9
assign po1404 = ~w9459;// level 9
assign po1405 = ~w9494;// level 9
assign po1406 = ~w9529;// level 9
assign po1407 = ~w9566;// level 9
assign po1408 = ~w9603;// level 9
assign po1409 = ~w9638;// level 9
assign po1410 = ~w9673;// level 9
assign po1411 = ~w9708;// level 9
assign po1412 = ~w9747;// level 9
assign po1413 = ~w9786;// level 9
assign po1414 = ~w9788;// level 7
assign po1415 = w9793;// level 15
assign po1416 = w9798;// level 16
assign po1417 = ~w9802;// level 16
assign po1418 = w9807;// level 15
assign po1419 = ~w9810;// level 8
assign po1420 = ~w9812;// level 7
assign po1421 = ~w9814;// level 7
assign po1422 = ~w9817;// level 5
assign po1423 = w9820;// level 3
assign po1424 = ~w8549;// level 8
assign po1425 = ~w9822;// level 7
assign po1426 = ~w9825;// level 5
assign po1427 = ~w9828;// level 5
assign po1428 = ~w9831;// level 8
assign po1429 = ~w9834;// level 8
assign po1430 = ~w9837;// level 8
assign po1431 = ~w9840;// level 8
assign po1432 = ~w9843;// level 8
assign po1433 = ~w9846;// level 8
assign po1434 = ~w9849;// level 8
assign po1435 = ~w9852;// level 8
assign po1436 = ~w9855;// level 8
assign po1437 = ~w9858;// level 8
assign po1438 = ~w9861;// level 8
assign po1439 = ~w9864;// level 8
assign po1440 = ~w9866;// level 7
assign po1441 = ~w9868;// level 7
assign po1442 = ~w9870;// level 7
assign po1443 = ~w9873;// level 5
assign po1444 = ~w9876;// level 5
assign po1445 = ~w9879;// level 5
assign po1446 = ~w9882;// level 5
assign po1447 = ~w9885;// level 8
assign po1448 = ~w9888;// level 8
assign po1449 = w9895;// level 18
assign po1450 = ~w9905;// level 17
assign po1451 = ~w9908;// level 8
assign po1452 = ~w9910;// level 7
assign po1453 = ~w9912;// level 7
assign po1454 = w9920;// level 5
assign po1455 = ~w9922;// level 7
assign po1456 = ~w9928;// level 8
assign po1457 = ~w9931;// level 8
assign po1458 = ~w9937;// level 8
assign po1459 = ~w9940;// level 8
assign po1460 = ~w9943;// level 8
assign po1461 = ~w9946;// level 8
assign po1462 = ~w9949;// level 8
assign po1463 = ~w9952;// level 8
assign po1464 = ~w9955;// level 8
assign po1465 = ~w9958;// level 8
assign po1466 = ~w9961;// level 8
assign po1467 = ~w9963;// level 7
assign po1468 = ~w9966;// level 8
assign po1469 = ~w9970;// level 8
assign po1470 = ~w9974;// level 8
assign po1471 = ~w9977;// level 8
assign po1472 = ~w9980;// level 8
assign po1473 = ~w9983;// level 8
assign po1474 = ~w10016;// level 9
assign po1475 = ~w10041;// level 8
assign po1476 = ~w10066;// level 8
assign po1477 = ~w10099;// level 9
assign po1478 = ~w10103;// level 8
assign po1479 = w10108;// level 8
assign po1480 = ~w10133;// level 8
assign po1481 = ~w10158;// level 8
assign po1482 = ~w10183;// level 8
assign po1483 = ~w10189;// level 8
assign po1484 = ~w10192;// level 8
assign po1485 = ~w10195;// level 8
assign po1486 = ~w10198;// level 8
assign po1487 = ~w10201;// level 8
assign po1488 = ~w10204;// level 8
assign po1489 = ~w10207;// level 8
assign po1490 = ~w10210;// level 8
assign po1491 = ~w10213;// level 8
assign po1492 = ~w10219;// level 8
assign po1493 = ~w10222;// level 8
assign po1494 = ~w10225;// level 8
assign po1495 = ~w10228;// level 8
assign po1496 = ~w10231;// level 8
assign po1497 = ~w10234;// level 8
assign po1498 = ~w10237;// level 8
assign po1499 = ~w10240;// level 8
assign po1500 = ~w10243;// level 8
assign po1501 = ~w10266;// level 8
assign po1502 = ~w10269;// level 8
assign po1503 = ~w10272;// level 8
assign po1504 = ~w10275;// level 8
assign po1505 = ~w10278;// level 8
assign po1506 = ~w10281;// level 8
assign po1507 = ~w10292;// level 17
assign po1508 = ~w10303;// level 18
assign po1509 = ~w10306;// level 8
assign po1510 = w10308;// level 4
assign po1511 = ~w10311;// level 8
assign po1512 = ~w10314;// level 8
assign po1513 = ~w10317;// level 8
assign po1514 = ~w10320;// level 8
assign po1515 = ~w10323;// level 8
assign po1516 = ~w10326;// level 8
assign po1517 = ~w10329;// level 8
assign po1518 = pi1418;// level 0
assign po1519 = ~w10332;// level 8
assign po1520 = ~w10335;// level 8
assign po1521 = ~w10339;// level 8
assign po1522 = ~w10362;// level 8
assign po1523 = ~w10385;// level 8
assign po1524 = w10397;// level 4
assign po1525 = w10409;// level 4
assign po1526 = w1232;// level 3
assign po1527 = w10413;// level 7
assign po1528 = ~w10415;// level 12
assign po1529 = ~w10428;// level 12
assign po1530 = w10429;// level 6
assign po1531 = w10432;// level 7
assign po1532 = w10434;// level 5
assign po1533 = w10437;// level 7
assign po1534 = w10440;// level 7
assign po1535 = w3574;// level 3
assign po1536 = w10443;// level 7
assign po1537 = w10444;// level 6
assign po1538 = w1813;// level 4
assign po1539 = ~w10446;// level 13
assign po1540 = ~w10448;// level 14
assign po1541 = ~w10450;// level 13
assign po1542 = w10463;// level 11
assign po1543 = ~w10466;// level 10
assign po1544 = ~w10478;// level 10
assign po1545 = w10479;// level 5
assign po1546 = ~w10481;// level 10
assign po1547 = w10482;// level 5
assign po1548 = w10483;// level 5
assign po1549 = ~w10486;// level 10
assign po1550 = ~w10488;// level 11
assign po1551 = ~w10490;// level 12
assign po1552 = ~w10492;// level 10
assign po1553 = ~w10507;// level 7
assign po1554 = w10511;// level 14
assign po1555 = w1828;// level 4
assign po1556 = ~w10525;// level 11
assign po1557 = ~w10529;// level 11
assign po1558 = w10531;// level 10
assign po1559 = ~w10533;// level 9
assign po1560 = w10535;// level 8
assign po1561 = w10537;// level 8
assign po1562 = ~w10539;// level 8
assign po1563 = ~w10541;// level 9
assign po1564 = ~w10543;// level 11
assign po1565 = ~w10546;// level 7
assign po1566 = w10549;// level 5
assign po1567 = w1844;// level 4
assign po1568 = w10556;// level 6
assign po1569 = ~w10558;// level 8
assign po1570 = ~w10560;// level 9
assign po1571 = w10565;// level 8
assign po1572 = w10568;// level 4
assign po1573 = w10571;// level 3
assign po1574 = w10572;// level 1
assign po1575 = ~w10574;// level 9
assign po1576 = ~w10576;// level 10
assign po1577 = ~w10578;// level 10
assign po1578 = ~w10595;// level 6
assign po1579 = ~w10612;// level 6
assign po1580 = w10615;// level 5
assign po1581 = w10616;// level 5
assign po1582 = ~w10618;// level 7
assign po1583 = ~w10620;// level 7
assign po1584 = w10624;// level 9
assign po1585 = w10633;// level 5
assign po1586 = w10636;// level 7
assign po1587 = w10638;// level 5
assign po1588 = w1859;// level 4
assign po1589 = w10641;// level 2
assign po1590 = ~w10643;// level 4
assign po1591 = ~w10645;// level 7
assign po1592 = ~w10647;// level 8
assign po1593 = ~w10649;// level 8
assign po1594 = ~w10651;// level 9
assign po1595 = ~w10652;// level 1
assign po1596 = ~w10654;// level 5
assign po1597 = ~w10656;// level 3
assign po1598 = ~w10658;// level 7
assign po1599 = w10666;// level 5
assign po1600 = w10676;// level 5
assign po1601 = w10679;// level 4
assign po1602 = w10682;// level 5
assign po1603 = w9917;// level 3
assign po1604 = ~pi1626;// level 0
assign po1605 = ~w10684;// level 4
assign po1606 = ~w10686;// level 8
assign po1607 = w10688;// level 8
assign po1608 = w10690;// level 7
assign po1609 = w10692;// level 7
assign po1610 = w10699;// level 6
assign po1611 = ~w10700;// level 1
assign po1612 = ~w10701;// level 1
assign po1613 = ~w10702;// level 1
assign po1614 = w10705;// level 5
assign po1615 = ~w10707;// level 5
assign po1616 = w10710;// level 4
assign po1617 = ~w10712;// level 3
assign po1618 = w10611;// level 5
assign po1619 = w10594;// level 5
assign po1620 = ~w10714;// level 6
assign po1621 = ~w10716;// level 6
assign po1622 = ~w10718;// level 6
assign po1623 = ~w10720;// level 6
assign po1624 = w10725;// level 8
assign po1625 = w10726;// level 1
assign po1626 = w10729;// level 3
assign po1627 = w10733;// level 9
assign po1628 = w10739;// level 5
assign po1629 = w10742;// level 7
assign po1630 = ~w10750;// level 8
assign po1631 = ~w10765;// level 4
assign po1632 = ~w10769;// level 4
assign po1633 = ~w10771;// level 4
assign po1634 = w10772;// level 3
assign po1635 = w10774;// level 7
assign po1636 = w10776;// level 7
assign po1637 = w10778;// level 6
assign po1638 = w10780;// level 6
assign po1639 = w10782;// level 6
assign po1640 = w10784;// level 5
assign po1641 = ~w10787;// level 4
assign po1642 = w10792;// level 4
assign po1643 = ~w10794;// level 5
assign po1644 = ~w10796;// level 3
assign po1645 = ~w10798;// level 5
assign po1646 = w6241;// level 4
assign po1647 = w10799;// level 6
assign po1648 = w10800;// level 5
assign po1649 = w10801;// level 5
assign po1650 = ~pi1625;// level 0
assign po1651 = pi1578;// level 0
assign po1652 = w10807;// level 3
assign po1653 = ~w10809;// level 3
assign po1654 = w10811;// level 6
assign po1655 = w9201;// level 6
assign po1656 = pi1627;// level 0
assign po1657 = ~pi1667;// level 0
assign po1658 = w10813;// level 4
assign po1659 = w10816;// level 3
assign po1660 = w10820;// level 5
assign po1661 = w10824;// level 5
assign po1662 = w10828;// level 8
assign po1663 = w10832;// level 5
assign po1664 = w10835;// level 3
assign po1665 = w10839;// level 4
assign po1666 = w10843;// level 4
assign po1667 = w10847;// level 4
assign po1668 = w10851;// level 4
assign po1669 = w10854;// level 3
assign po1670 = w10857;// level 3
assign po1671 = ~w10860;// level 3
assign po1672 = ~w10863;// level 3
assign po1673 = w10865;// level 2
assign po1674 = w10867;// level 2
assign po1675 = w10869;// level 2
assign po1676 = w381;// level 2
assign po1677 = w10870;// level 2
assign po1678 = w372;// level 2
assign po1679 = w10871;// level 2
assign po1680 = w10872;// level 2
assign po1681 = ~w10875;// level 3
assign po1682 = ~w10878;// level 3
assign po1683 = ~w10881;// level 3
assign po1684 = ~w10884;// level 3
assign po1685 = ~w10887;// level 3
assign po1686 = pi0954;// level 0
assign po1687 = w1;// level 2
assign po1688 = w1213;// level 2
assign po1689 = ~w10888;// level 2
assign po1690 = w1209;// level 2
assign po1691 = w10891;// level 3
assign po1692 = ~w10894;// level 3
assign po1693 = ~w10897;// level 3
assign po1694 = ~w10900;// level 3
assign po1695 = ~w10903;// level 3
assign po1696 = ~w10906;// level 3
assign po1697 = ~w10909;// level 3
assign po1698 = ~w10912;// level 3
assign po1699 = ~w10915;// level 3
assign po1700 = ~w10918;// level 3
assign po1701 = ~w10921;// level 3
assign po1702 = w10922;// level 2
assign po1703 = ~w10925;// level 3
assign po1704 = ~w10928;// level 3
assign po1705 = ~w10931;// level 3
assign po1706 = ~w10934;// level 3
assign po1707 = ~w10937;// level 3
assign po1708 = ~w10940;// level 3
assign po1709 = ~w10943;// level 3
assign po1710 = ~w10946;// level 3
assign po1711 = ~w10949;// level 3
assign po1712 = w10952;// level 3
assign po1713 = ~w10955;// level 3
assign po1714 = ~w10958;// level 3
assign po1715 = w10961;// level 3
assign po1716 = w10964;// level 3
assign po1717 = ~w10967;// level 3
assign po1718 = ~w10970;// level 3
assign po1719 = ~w10982;// level 4
assign po1720 = ~w10994;// level 4
assign po1721 = ~w11006;// level 4
assign po1722 = ~w11009;// level 3
assign po1723 = ~w11012;// level 3
assign po1724 = ~w11023;// level 4
assign po1725 = ~w11034;// level 4
assign po1726 = ~w11045;// level 4
assign po1727 = ~w11057;// level 4
assign po1728 = ~w11068;// level 4
assign po1729 = w11074;// level 3
assign po1730 = ~w11076;// level 2
assign po1731 = ~w11078;// level 2
assign po1732 = ~w11080;// level 2
assign po1733 = ~w185;// level 1
assign po1734 = w11081;// level 1
assign po1735 = w11082;// level 1
assign po1736 = w11083;// level 1
assign po1737 = w2132;// level 1
assign po1738 = ~w11085;// level 2
assign po1739 = w11086;// level 3
assign po1740 = ~w11090;// level 3
assign po1741 = ~w11093;// level 3
assign po1742 = ~w11096;// level 3
assign po1743 = ~w11099;// level 3
assign po1744 = ~w11102;// level 3
assign po1745 = w11104;// level 2
assign po1746 = ~w11107;// level 3
assign po1747 = ~w11110;// level 3
assign po1748 = ~w11113;// level 3
assign po1749 = ~w11116;// level 3
assign po1750 = ~w11119;// level 3
assign po1751 = ~w11122;// level 3
assign po1752 = ~w11125;// level 3
assign po1753 = ~w11128;// level 3
assign po1754 = ~w11131;// level 3
assign po1755 = ~w11134;// level 3
assign po1756 = ~w11137;// level 3
assign po1757 = ~w11140;// level 3
assign po1758 = ~w11143;// level 3
assign po1759 = ~w11146;// level 3
assign po1760 = ~w11149;// level 3
assign po1761 = ~w11152;// level 3
assign po1762 = ~w11155;// level 3
assign po1763 = ~w11158;// level 3
assign po1764 = ~w11161;// level 3
assign po1765 = ~w11164;// level 3
assign po1766 = ~w11167;// level 3
assign po1767 = ~w11170;// level 3
assign po1768 = ~w11173;// level 3
assign po1769 = ~w11176;// level 3
assign po1770 = ~w11179;// level 3
assign po1771 = ~w11182;// level 3
assign po1772 = ~w11185;// level 3
assign po1773 = w11188;// level 2
assign po1774 = w11189;// level 1
assign po1775 = ~w2135;// level 1
assign po1776 = w6396;// level 1
assign po1777 = ~w4;// level 2
assign po1778 = w11191;// level 2
assign po1779 = w11194;// level 3
assign po1780 = w11195;// level 1
assign po1781 = w11196;// level 2
assign po1782 = w6807;// level 1
assign po1783 = pi1680;// level 0
assign po1784 = ~pi1726;// level 0
assign po1785 = ~w6718;// level 1
assign po1786 = ~pi1192;// level 0
assign po1787 = pi1730;// level 0
assign po1788 = pi1038;// level 0
assign po1789 = pi1719;// level 0
assign po1790 = pi1723;// level 0
assign po1791 = pi1724;// level 0
assign po1792 = pi1720;// level 0
assign po1793 = pi1736;// level 0
assign po1794 = pi1732;// level 0
assign po1795 = pi1745;// level 0
assign po1796 = w11197;// level 1
assign po1797 = pi1734;// level 0
assign po1798 = pi1753;// level 0
assign po1799 = pi1744;// level 0
assign po1800 = pi1743;// level 0
assign po1801 = pi0112;// level 0
assign po1802 = pi1728;// level 0
assign po1803 = pi1721;// level 0
assign po1804 = ~pi1241;// level 0
assign po1805 = ~pi1213;// level 0
assign po1806 = ~pi1331;// level 0
assign po1807 = ~pi0787;// level 0
assign po1808 = ~pi1426;// level 0
assign po1809 = ~pi1428;// level 0
assign po1810 = ~pi1425;// level 0
assign po1811 = ~pi0944;// level 0
assign po1812 = ~pi1419;// level 0
assign po1813 = ~pi0936;// level 0
assign po1814 = ~pi0943;// level 0
assign po1815 = ~pi0932;// level 0
assign po1816 = ~pi0933;// level 0
assign po1817 = ~pi1423;// level 0
assign po1818 = ~pi0931;// level 0
assign po1819 = ~pi0934;// level 0
assign po1820 = ~pi0935;// level 0
assign po1821 = pi1855;// level 0
assign po1822 = pi1851;// level 0
assign po1823 = pi1853;// level 0
assign po1824 = pi1844;// level 0
assign po1825 = pi1852;// level 0
assign po1826 = pi0794;// level 0
assign po1827 = pi1849;// level 0
assign po1828 = pi1457;// level 0
assign po1829 = pi1845;// level 0
assign po1830 = pi1562;// level 0
assign po1831 = pi1099;// level 0
assign po1832 = pi1556;// level 0
assign po1833 = pi1858;// level 0
assign po1834 = pi1854;// level 0
assign po1835 = pi1842;// level 0
assign po1836 = pi1561;// level 0
assign po1837 = pi1847;// level 0
assign po1838 = pi1857;// level 0
assign po1839 = pi1859;// level 0
assign po1840 = pi1848;// level 0
assign po1841 = pi1846;// level 0
assign po1842 = pi1843;// level 0
assign po1843 = pi1551;// level 0
assign po1844 = pi1856;// level 0
assign po1845 = pi1850;// level 0
endmodule
