//Written by the Majority Logic Package Thu Apr 30 13:27:53 2015
module top (
            pi000, pi001, pi002, pi003, pi004, pi005, pi006, pi007, pi008, pi009, pi010, pi011, pi012, pi013, pi014, pi015, pi016, pi017, pi018, pi019, pi020, pi021, pi022, pi023, pi024, pi025, pi026, pi027, pi028, pi029, pi030, pi031, pi032, pi033, pi034, pi035, pi036, pi037, pi038, pi039, pi040, pi041, pi042, pi043, pi044, pi045, pi046, pi047, pi048, pi049, pi050, pi051, pi052, pi053, pi054, pi055, pi056, pi057, pi058, pi059, pi060, pi061, pi062, pi063, pi064, pi065, pi066, pi067, pi068, pi069, pi070, pi071, pi072, pi073, pi074, pi075, pi076, pi077, pi078, pi079, pi080, pi081, pi082, pi083, pi084, pi085, pi086, pi087, pi088, pi089, pi090, pi091, pi092, pi093, pi094, pi095, pi096, pi097, pi098, pi099, pi100, pi101, pi102, pi103, pi104, pi105, pi106, pi107, pi108, pi109, pi110, pi111, pi112, pi113, pi114, pi115, pi116, pi117, pi118, pi119, pi120, pi121, pi122, pi123, pi124, pi125, pi126, pi127, pi128, pi129, pi130, pi131, pi132, pi133, pi134, pi135, pi136, pi137, pi138, pi139, pi140, pi141, pi142, pi143, pi144, pi145, pi146, pi147, 
            po000, po001, po002, po003, po004, po005, po006, po007, po008, po009, po010, po011, po012, po013, po014, po015, po016, po017, po018, po019, po020, po021, po022, po023, po024, po025, po026, po027, po028, po029, po030, po031, po032, po033, po034, po035, po036, po037, po038, po039, po040, po041, po042, po043, po044, po045, po046, po047, po048, po049, po050, po051, po052, po053, po054, po055, po056, po057, po058, po059, po060, po061, po062, po063, po064, po065, po066, po067, po068, po069, po070, po071, po072, po073, po074, po075, po076, po077, po078, po079, po080, po081, po082, po083, po084, po085, po086, po087, po088, po089, po090, po091, po092, po093, po094, po095, po096, po097, po098, po099, po100, po101, po102, po103, po104, po105, po106, po107, po108, po109, po110, po111, po112, po113, po114, po115, po116, po117, po118, po119, po120, po121, po122, po123, po124, po125, po126, po127, po128, po129, po130, po131, po132, po133, po134, po135, po136, po137, po138, po139, po140, po141, po142, po143, po144, po145, po146);
input pi000, pi001, pi002, pi003, pi004, pi005, pi006, pi007, pi008, pi009, pi010, pi011, pi012, pi013, pi014, pi015, pi016, pi017, pi018, pi019, pi020, pi021, pi022, pi023, pi024, pi025, pi026, pi027, pi028, pi029, pi030, pi031, pi032, pi033, pi034, pi035, pi036, pi037, pi038, pi039, pi040, pi041, pi042, pi043, pi044, pi045, pi046, pi047, pi048, pi049, pi050, pi051, pi052, pi053, pi054, pi055, pi056, pi057, pi058, pi059, pi060, pi061, pi062, pi063, pi064, pi065, pi066, pi067, pi068, pi069, pi070, pi071, pi072, pi073, pi074, pi075, pi076, pi077, pi078, pi079, pi080, pi081, pi082, pi083, pi084, pi085, pi086, pi087, pi088, pi089, pi090, pi091, pi092, pi093, pi094, pi095, pi096, pi097, pi098, pi099, pi100, pi101, pi102, pi103, pi104, pi105, pi106, pi107, pi108, pi109, pi110, pi111, pi112, pi113, pi114, pi115, pi116, pi117, pi118, pi119, pi120, pi121, pi122, pi123, pi124, pi125, pi126, pi127, pi128, pi129, pi130, pi131, pi132, pi133, pi134, pi135, pi136, pi137, pi138, pi139, pi140, pi141, pi142, pi143, pi144, pi145, pi146, pi147;
output po000, po001, po002, po003, po004, po005, po006, po007, po008, po009, po010, po011, po012, po013, po014, po015, po016, po017, po018, po019, po020, po021, po022, po023, po024, po025, po026, po027, po028, po029, po030, po031, po032, po033, po034, po035, po036, po037, po038, po039, po040, po041, po042, po043, po044, po045, po046, po047, po048, po049, po050, po051, po052, po053, po054, po055, po056, po057, po058, po059, po060, po061, po062, po063, po064, po065, po066, po067, po068, po069, po070, po071, po072, po073, po074, po075, po076, po077, po078, po079, po080, po081, po082, po083, po084, po085, po086, po087, po088, po089, po090, po091, po092, po093, po094, po095, po096, po097, po098, po099, po100, po101, po102, po103, po104, po105, po106, po107, po108, po109, po110, po111, po112, po113, po114, po115, po116, po117, po118, po119, po120, po121, po122, po123, po124, po125, po126, po127, po128, po129, po130, po131, po132, po133, po134, po135, po136, po137, po138, po139, po140, po141, po142, po143, po144, po145, po146;
wire one, w0, w1, w2, w3, w4, w5, w6, w7, w8, w9, w10, w11, w12, w13, w14, w15, w16, w17, w18, w19, w20, w21, w22, w23, w24, w25, w26, w27, w28, w29, w30, w31, w32, w33, w34, w35, w36, w37, w38, w39, w40, w41, w42, w43, w44, w45, w46, w47, w48, w49, w50, w51, w52, w53, w54, w55, w56, w57, w58, w59, w60, w61, w62, w63, w64, w65, w66, w67, w68, w69, w70, w71, w72, w73, w74, w75, w76, w77, w78, w79, w80, w81, w82, w83, w84, w85, w86, w87, w88, w89, w90, w91, w92, w93, w94, w95, w96, w97, w98, w99, w100, w101, w102, w103, w104, w105, w106, w107, w108, w109, w110, w111, w112, w113, w114, w115, w116, w117, w118, w119, w120, w121, w122, w123, w124, w125, w126, w127, w128, w129, w130, w131, w132, w133, w134, w135, w136, w137, w138, w139, w140, w141, w142, w143, w144, w145, w146, w147, w148, w149, w150, w151, w152, w153, w154, w155, w156, w157, w158, w159, w160, w161, w162, w163, w164, w165, w166, w167, w168, w169, w170, w171, w172, w173, w174, w175, w176, w177, w178, w179, w180, w181, w182, w183, w184, w185, w186, w187, w188, w189, w190, w191, w192, w193, w194, w195, w196, w197, w198, w199, w200, w201, w202, w203, w204, w205, w206, w207, w208, w209, w210, w211, w212, w213, w214, w215, w216, w217, w218, w219, w220, w221, w222, w223, w224, w225, w226, w227, w228, w229, w230, w231, w232, w233, w234, w235, w236, w237, w238, w239, w240, w241, w242, w243, w244, w245, w246, w247, w248, w249, w250, w251, w252, w253, w254, w255, w256, w257, w258, w259, w260, w261, w262, w263, w264, w265, w266, w267, w268, w269, w270, w271, w272, w273, w274, w275, w276, w277, w278, w279, w280, w281, w282, w283, w284, w285, w286, w287, w288, w289, w290, w291, w292, w293, w294, w295, w296, w297, w298, w299, w300, w301, w302, w303, w304, w305, w306, w307, w308, w309, w310, w311, w312, w313, w314, w315, w316, w317, w318, w319, w320, w321, w322, w323, w324, w325, w326, w327, w328, w329, w330, w331, w332, w333, w334, w335, w336, w337, w338, w339, w340, w341, w342, w343, w344, w345, w346, w347, w348, w349, w350, w351, w352, w353, w354, w355, w356, w357, w358, w359, w360, w361, w362, w363, w364, w365, w366, w367, w368, w369, w370, w371, w372, w373, w374, w375, w376, w377, w378, w379, w380, w381, w382, w383, w384, w385, w386, w387, w388, w389, w390, w391, w392, w393, w394, w395, w396, w397, w398, w399, w400, w401, w402, w403, w404, w405, w406, w407, w408, w409, w410, w411, w412, w413, w414, w415, w416, w417, w418, w419, w420, w421, w422, w423, w424, w425, w426, w427, w428, w429, w430, w431, w432, w433, w434, w435, w436, w437, w438, w439, w440, w441, w442, w443, w444, w445, w446, w447, w448, w449, w450, w451, w452, w453, w454, w455, w456, w457, w458, w459, w460, w461, w462, w463, w464, w465, w466, w467, w468, w469, w470, w471, w472, w473, w474, w475, w476, w477, w478, w479, w480, w481, w482, w483, w484, w485, w486, w487, w488, w489, w490, w491, w492, w493, w494, w495, w496, w497, w498, w499, w500, w501, w502, w503, w504, w505, w506, w507, w508, w509, w510, w511, w512, w513, w514, w515, w516, w517, w518, w519, w520, w521, w522, w523, w524, w525, w526, w527, w528, w529, w530, w531, w532, w533, w534, w535, w536, w537, w538, w539, w540, w541, w542, w543, w544, w545, w546, w547, w548, w549, w550, w551, w552, w553, w554, w555, w556, w557, w558, w559, w560, w561, w562, w563, w564, w565, w566, w567, w568, w569, w570, w571, w572, w573, w574, w575, w576, w577, w578, w579, w580, w581, w582, w583, w584, w585, w586, w587, w588, w589, w590, w591, w592, w593, w594, w595, w596, w597, w598, w599, w600, w601, w602, w603, w604, w605, w606, w607, w608, w609, w610, w611, w612, w613, w614, w615, w616, w617, w618, w619, w620, w621, w622, w623, w624, w625, w626, w627, w628, w629, w630, w631, w632, w633, w634, w635, w636, w637, w638, w639, w640, w641, w642, w643, w644, w645, w646, w647, w648, w649, w650, w651, w652, w653, w654, w655, w656, w657, w658, w659, w660, w661, w662, w663, w664, w665, w666, w667, w668, w669, w670, w671, w672, w673, w674, w675, w676, w677, w678, w679, w680, w681, w682, w683, w684, w685, w686, w687, w688, w689, w690, w691, w692, w693, w694, w695, w696, w697, w698, w699, w700, w701, w702, w703, w704, w705, w706, w707, w708, w709, w710, w711, w712, w713, w714, w715, w716, w717, w718, w719, w720, w721, w722, w723, w724, w725, w726, w727, w728, w729, w730, w731, w732, w733, w734, w735, w736, w737, w738, w739, w740, w741, w742, w743, w744, w745, w746, w747, w748, w749, w750, w751, w752, w753, w754, w755, w756, w757, w758, w759, w760, w761, w762, w763, w764, w765, w766, w767, w768, w769, w770, w771, w772, w773, w774, w775, w776, w777, w778, w779, w780, w781, w782, w783, w784, w785, w786, w787, w788, w789, w790, w791, w792, w793, w794, w795, w796, w797, w798, w799, w800, w801, w802, w803, w804, w805, w806, w807, w808, w809, w810, w811, w812, w813, w814, w815, w816, w817, w818, w819, w820, w821, w822, w823, w824, w825, w826, w827, w828, w829, w830, w831, w832, w833, w834, w835, w836;
assign w0 = ~pi000 & ~pi002;
assign w1 = (pi128 & ~w0) | (pi128 & w745) | (~w0 & w745);
assign w2 = pi120 & ~w1;
assign w3 = ~pi002 & ~pi063;
assign w4 = pi128 & ~w3;
assign w5 = ~w3 & w746;
assign w6 = ~w2 & ~w5;
assign w7 = pi128 & pi133;
assign w8 = ~pi138 & pi139;
assign w9 = pi134 & pi135;
assign w10 = pi130 & w9;
assign w11 = w10 & w722;
assign w12 = pi001 & ~w11;
assign w13 = pi004 & ~pi075;
assign w14 = ~pi004 & pi075;
assign w15 = ~w13 & ~w14;
assign w16 = ~pi005 & pi077;
assign w17 = w15 & ~w16;
assign w18 = pi005 & ~pi077;
assign w19 = (~pi063 & w15) | (~pi063 & w747) | (w15 & w747);
assign w20 = ~w17 & w19;
assign w21 = ~w12 & ~w20;
assign w22 = w7 & ~w21;
assign w23 = (~pi119 & w0) | (~pi119 & w748) | (w0 & w748);
assign w24 = pi002 & pi063;
assign w25 = w4 & ~w24;
assign w26 = ~w23 & ~w25;
assign w27 = pi136 & w9;
assign w28 = pi138 & ~pi139;
assign w29 = w27 & w28;
assign w30 = w27 & w749;
assign w31 = (~pi003 & ~w0) | (~pi003 & w750) | (~w0 & w750);
assign w32 = pi128 & ~w31;
assign w33 = ~w30 & w32;
assign w34 = pi005 & ~pi063;
assign w35 = pi004 & w34;
assign w36 = (pi128 & w34) | (pi128 & w751) | (w34 & w751);
assign w37 = ~w35 & w36;
assign w38 = ~pi005 & pi063;
assign w39 = pi128 & ~w34;
assign w40 = ~w38 & w39;
assign w41 = (pi006 & ~w34) | (pi006 & w752) | (~w34 & w752);
assign w42 = w34 & w753;
assign w43 = ~w41 & ~w42;
assign w44 = (pi007 & ~w34) | (pi007 & w754) | (~w34 & w754);
assign w45 = w34 & w755;
assign w46 = ~w44 & ~w45;
assign w47 = (pi008 & ~w34) | (pi008 & w756) | (~w34 & w756);
assign w48 = w34 & w757;
assign w49 = ~w47 & ~w48;
assign w50 = (pi009 & ~w34) | (pi009 & w758) | (~w34 & w758);
assign w51 = w34 & w759;
assign w52 = ~w50 & ~w51;
assign w53 = (pi010 & ~w34) | (pi010 & w760) | (~w34 & w760);
assign w54 = w34 & w761;
assign w55 = ~w53 & ~w54;
assign w56 = pi004 & ~pi005;
assign w57 = (pi011 & ~w56) | (pi011 & w762) | (~w56 & w762);
assign w58 = pi050 & ~pi063;
assign w59 = w56 & w58;
assign w60 = ~w57 & ~w59;
assign w61 = (pi012 & ~w56) | (pi012 & w763) | (~w56 & w763);
assign w62 = pi051 & ~pi063;
assign w63 = w56 & w62;
assign w64 = ~w61 & ~w63;
assign w65 = (pi013 & ~w56) | (pi013 & w764) | (~w56 & w764);
assign w66 = pi045 & ~pi063;
assign w67 = w56 & w66;
assign w68 = ~w65 & ~w67;
assign w69 = (pi014 & ~w56) | (pi014 & w765) | (~w56 & w765);
assign w70 = pi046 & ~pi063;
assign w71 = w56 & w70;
assign w72 = ~w69 & ~w71;
assign w73 = (pi015 & ~w56) | (pi015 & w766) | (~w56 & w766);
assign w74 = pi047 & ~pi063;
assign w75 = w56 & w74;
assign w76 = ~w73 & ~w75;
assign w77 = (pi016 & ~w56) | (pi016 & w767) | (~w56 & w767);
assign w78 = pi048 & ~pi063;
assign w79 = w56 & w78;
assign w80 = ~w77 & ~w79;
assign w81 = (pi017 & ~w56) | (pi017 & w768) | (~w56 & w768);
assign w82 = pi049 & ~pi063;
assign w83 = w56 & w82;
assign w84 = ~w81 & ~w83;
assign w85 = (pi018 & ~w56) | (pi018 & w769) | (~w56 & w769);
assign w86 = pi043 & ~pi063;
assign w87 = w56 & w86;
assign w88 = ~w85 & ~w87;
assign w89 = (pi019 & ~w34) | (pi019 & w770) | (~w34 & w770);
assign w90 = w34 & w771;
assign w91 = ~w89 & ~w90;
assign w92 = (pi020 & ~w34) | (pi020 & w772) | (~w34 & w772);
assign w93 = w34 & w773;
assign w94 = ~w92 & ~w93;
assign w95 = (pi021 & ~w34) | (pi021 & w774) | (~w34 & w774);
assign w96 = w34 & w775;
assign w97 = ~w95 & ~w96;
assign w98 = (pi022 & ~w34) | (pi022 & w776) | (~w34 & w776);
assign w99 = w34 & w777;
assign w100 = ~w98 & ~w99;
assign w101 = (pi023 & ~w34) | (pi023 & w778) | (~w34 & w778);
assign w102 = w34 & w779;
assign w103 = ~w101 & ~w102;
assign w104 = (pi024 & ~w34) | (pi024 & w780) | (~w34 & w780);
assign w105 = w34 & w781;
assign w106 = ~w104 & ~w105;
assign w107 = (pi025 & ~w34) | (pi025 & w782) | (~w34 & w782);
assign w108 = w34 & w783;
assign w109 = ~w107 & ~w108;
assign w110 = (pi026 & ~w34) | (pi026 & w784) | (~w34 & w784);
assign w111 = w34 & w785;
assign w112 = ~w110 & ~w111;
assign w113 = (pi027 & ~w34) | (pi027 & w786) | (~w34 & w786);
assign w114 = w34 & w787;
assign w115 = ~w113 & ~w114;
assign w116 = (pi028 & ~w34) | (pi028 & w788) | (~w34 & w788);
assign w117 = w34 & w789;
assign w118 = ~w116 & ~w117;
assign w119 = (pi029 & ~w34) | (pi029 & w790) | (~w34 & w790);
assign w120 = w34 & w791;
assign w121 = ~w119 & ~w120;
assign w122 = ~pi004 & ~pi005;
assign w123 = (pi030 & ~w122) | (pi030 & w792) | (~w122 & w792);
assign w124 = w58 & w122;
assign w125 = ~w123 & ~w124;
assign w126 = (pi031 & ~w122) | (pi031 & w793) | (~w122 & w793);
assign w127 = w62 & w122;
assign w128 = ~w126 & ~w127;
assign w129 = (pi032 & ~w122) | (pi032 & w794) | (~w122 & w794);
assign w130 = w70 & w122;
assign w131 = ~w129 & ~w130;
assign w132 = (pi033 & ~w122) | (pi033 & w795) | (~w122 & w795);
assign w133 = w74 & w122;
assign w134 = ~w132 & ~w133;
assign w135 = (pi034 & ~w122) | (pi034 & w796) | (~w122 & w796);
assign w136 = w78 & w122;
assign w137 = ~w135 & ~w136;
assign w138 = (pi035 & ~w122) | (pi035 & w797) | (~w122 & w797);
assign w139 = w86 & w122;
assign w140 = ~w138 & ~w139;
assign w141 = (pi036 & ~w122) | (pi036 & w798) | (~w122 & w798);
assign w142 = w66 & w122;
assign w143 = ~w141 & ~w142;
assign w144 = (pi037 & ~w122) | (pi037 & w799) | (~w122 & w799);
assign w145 = w82 & w122;
assign w146 = ~w144 & ~w145;
assign w147 = ~pi059 & ~pi060;
assign w148 = ~pi058 & w147;
assign w149 = w147 & w670;
assign w150 = ~pi054 & w149;
assign w151 = w149 & w671;
assign w152 = w149 & w672;
assign w153 = ~pi053 & w152;
assign w154 = w152 & w673;
assign w155 = w152 & w674;
assign w156 = w152 & w675;
assign w157 = w152 & w695;
assign w158 = pi039 & w157;
assign w159 = ~pi040 & ~pi044;
assign w160 = ~pi041 & w159;
assign w161 = (~pi038 & ~w159) | (~pi038 & w800) | (~w159 & w800);
assign w162 = w159 & w801;
assign w163 = ~w161 & ~w162;
assign w164 = w157 & w802;
assign w165 = pi083 & ~pi129;
assign w166 = ~pi083 & pi129;
assign w167 = pi076 & ~pi082;
assign w168 = ~pi076 & pi082;
assign w169 = ~w167 & ~w168;
assign w170 = ~w166 & w169;
assign w171 = w169 & w676;
assign w172 = ~pi039 & ~pi062;
assign w173 = w172 & w835;
assign w174 = (pi128 & w164) | (pi128 & w678) | (w164 & w678);
assign w175 = w157 & w723;
assign w176 = pi128 & ~w172;
assign w177 = ~pi062 & w157;
assign w178 = (w157 & w724) | (w157 & w725) | (w724 & w725);
assign w179 = ~w175 & w178;
assign w180 = ~w174 & ~w179;
assign w181 = pi039 & pi128;
assign w182 = pi128 & w172;
assign w183 = (w182 & ~w171) | (w182 & w803) | (~w171 & w803);
assign w184 = ~w181 & ~w183;
assign w185 = w157 & w804;
assign w186 = ~w184 & ~w185;
assign w187 = (pi040 & ~w157) | (pi040 & w726) | (~w157 & w726);
assign w188 = (~w172 & ~w157) | (~w172 & w727) | (~w157 & w727);
assign w189 = ~w187 & w188;
assign w190 = pi128 & ~w189;
assign w191 = w157 & w703;
assign w192 = ~pi041 & ~w172;
assign w193 = (w192 & ~w157) | (w192 & w805) | (~w157 & w805);
assign w194 = w157 & w728;
assign w195 = pi128 & ~w194;
assign w196 = ~w193 & w195;
assign w197 = (w374 & w176) | (w374 & ~w156) | (w176 & ~w156);
assign w198 = (w156 & w704) | (w156 & w705) | (w704 & w705);
assign w199 = (w156 & w806) | (w156 & w807) | (w806 & w807);
assign w200 = (w156 & w729) | (w156 & w730) | (w729 & w730);
assign w201 = (pi042 & ~w152) | (pi042 & w706) | (~w152 & w706);
assign w202 = ~w154 & ~w201;
assign w203 = w197 & ~w202;
assign w204 = ~w200 & ~w203;
assign w205 = ~w199 & w204;
assign w206 = pi043 & w836;
assign w207 = w157 & w709;
assign w208 = ~pi076 & ~pi129;
assign w209 = pi099 & w208;
assign w210 = pi076 & pi129;
assign w211 = pi111 & w210;
assign w212 = ~w209 & ~w211;
assign w213 = pi076 & ~pi129;
assign w214 = pi095 & w213;
assign w215 = ~pi076 & pi129;
assign w216 = pi089 & w215;
assign w217 = ~w214 & ~w216;
assign w218 = w212 & w217;
assign w219 = w172 & ~w218;
assign w220 = ~w207 & ~w219;
assign w221 = ~w206 & w220;
assign w222 = pi128 & ~w221;
assign w223 = ~pi044 & ~w172;
assign w224 = (~w223 & ~w157) | (~w223 & w731) | (~w157 & w731);
assign w225 = ~w191 & ~w224;
assign w226 = pi128 & ~w225;
assign w227 = pi045 & w836;
assign w228 = w157 & w710;
assign w229 = pi091 & w213;
assign w230 = pi086 & w215;
assign w231 = ~w229 & ~w230;
assign w232 = pi107 & w210;
assign w233 = pi102 & w208;
assign w234 = ~w232 & ~w233;
assign w235 = w231 & w234;
assign w236 = w172 & ~w235;
assign w237 = ~w228 & ~w236;
assign w238 = ~w227 & w237;
assign w239 = pi128 & ~w238;
assign w240 = pi046 & w836;
assign w241 = w157 & w711;
assign w242 = pi087 & w215;
assign w243 = pi092 & w213;
assign w244 = ~w242 & ~w243;
assign w245 = pi108 & w210;
assign w246 = pi103 & w208;
assign w247 = ~w245 & ~w246;
assign w248 = w244 & w247;
assign w249 = w172 & ~w248;
assign w250 = ~w241 & ~w249;
assign w251 = ~w240 & w250;
assign w252 = pi128 & ~w251;
assign w253 = pi047 & w836;
assign w254 = w157 & w712;
assign w255 = pi096 & w208;
assign w256 = pi097 & w210;
assign w257 = ~w255 & ~w256;
assign w258 = pi078 & w213;
assign w259 = pi081 & w215;
assign w260 = ~w258 & ~w259;
assign w261 = w257 & w260;
assign w262 = w172 & ~w261;
assign w263 = ~w254 & ~w262;
assign w264 = ~w253 & w263;
assign w265 = pi128 & ~w264;
assign w266 = pi048 & w836;
assign w267 = w157 & w713;
assign w268 = pi105 & w208;
assign w269 = pi109 & w210;
assign w270 = ~w268 & ~w269;
assign w271 = pi093 & w213;
assign w272 = pi088 & w215;
assign w273 = ~w271 & ~w272;
assign w274 = w270 & w273;
assign w275 = w172 & ~w274;
assign w276 = ~w267 & ~w275;
assign w277 = ~w266 & w276;
assign w278 = pi128 & ~w277;
assign w279 = pi049 & w836;
assign w280 = w157 & w714;
assign w281 = pi094 & w213;
assign w282 = pi079 & w215;
assign w283 = ~w281 & ~w282;
assign w284 = pi104 & w208;
assign w285 = pi110 & w210;
assign w286 = ~w284 & ~w285;
assign w287 = w283 & w286;
assign w288 = w172 & ~w287;
assign w289 = ~w280 & ~w288;
assign w290 = ~w279 & w289;
assign w291 = pi128 & ~w290;
assign w292 = pi050 & w836;
assign w293 = w157 & w715;
assign w294 = pi100 & w208;
assign w295 = pi098 & w210;
assign w296 = ~w294 & ~w295;
assign w297 = pi084 & w215;
assign w298 = pi080 & w213;
assign w299 = ~w297 & ~w298;
assign w300 = w296 & w299;
assign w301 = w172 & ~w300;
assign w302 = ~w293 & ~w301;
assign w303 = ~w292 & w302;
assign w304 = pi128 & ~w303;
assign w305 = pi051 & w836;
assign w306 = pi085 & w215;
assign w307 = pi090 & w213;
assign w308 = ~w306 & ~w307;
assign w309 = pi106 & w210;
assign w310 = pi101 & w208;
assign w311 = ~w309 & ~w310;
assign w312 = w308 & w311;
assign w313 = w172 & ~w312;
assign w314 = (~w313 & ~w158) | (~w313 & w690) | (~w158 & w690);
assign w315 = ~w305 & w314;
assign w316 = pi128 & ~w315;
assign w317 = (pi052 & ~w152) | (pi052 & w732) | (~w152 & w732);
assign w318 = ~w156 & ~w317;
assign w319 = w197 & ~w318;
assign w320 = pi123 & pi126;
assign w321 = (w156 & w808) | (w156 & w809) | (w808 & w809);
assign w322 = ~w319 & ~w321;
assign w323 = pi053 & ~w152;
assign w324 = ~w153 & ~w323;
assign w325 = w197 & ~w324;
assign w326 = ~w198 & ~w325;
assign w327 = (w156 & w733) | (w156 & w734) | (w733 & w734);
assign w328 = pi126 & w327;
assign w329 = pi114 & ~pi123;
assign w330 = (w156 & w735) | (w156 & w736) | (w735 & w736);
assign w331 = pi054 & ~w149;
assign w332 = ~w150 & ~w331;
assign w333 = w197 & w332;
assign w334 = ~w330 & ~w333;
assign w335 = ~w328 & ~w334;
assign w336 = (w156 & w737) | (w156 & w738) | (w737 & w738);
assign w337 = (pi055 & ~w147) | (pi055 & w810) | (~w147 & w810);
assign w338 = ~w149 & ~w337;
assign w339 = w338 & w197;
assign w340 = ~w336 & ~w339;
assign w341 = w320 & w327;
assign w342 = (pi056 & ~w149) | (pi056 & w739) | (~w149 & w739);
assign w343 = ~w152 & ~w342;
assign w344 = w197 & ~w343;
assign w345 = ~w198 & ~w344;
assign w346 = ~w341 & w345;
assign w347 = (pi057 & ~w152) | (pi057 & w740) | (~w152 & w740);
assign w348 = ~w155 & ~w347;
assign w349 = w197 & ~w348;
assign w350 = ~w200 & ~w349;
assign w351 = ~pi114 & w336;
assign w352 = pi058 & ~w147;
assign w353 = ~w148 & ~w352;
assign w354 = w353 & w197;
assign w355 = ~w351 & ~w354;
assign w356 = pi059 & w197;
assign w357 = ~pi114 & ~pi126;
assign w358 = (w156 & w741) | (w156 & w742) | (w741 & w742);
assign w359 = ~pi123 & w358;
assign w360 = ~w356 & ~w359;
assign w361 = pi059 & pi060;
assign w362 = ~w147 & ~w361;
assign w363 = w362 & w197;
assign w364 = ~w358 & ~w363;
assign w365 = (pi061 & ~w149) | (pi061 & w743) | (~w149 & w743);
assign w366 = ~w151 & ~w365;
assign w367 = w197 & ~w366;
assign w368 = ~w198 & ~w367;
assign w369 = ~w328 & w368;
assign w370 = pi062 & ~w157;
assign w371 = ~w177 & ~w370;
assign w372 = w181 & ~w371;
assign w373 = pi128 & w185;
assign w374 = ~w172 & w811;
assign w375 = ~w156 & w374;
assign w376 = ~pi075 & pi077;
assign w377 = pi009 & w376;
assign w378 = pi075 & pi077;
assign w379 = pi028 & w378;
assign w380 = ~w377 & ~w379;
assign w381 = pi075 & ~pi077;
assign w382 = pi017 & w381;
assign w383 = ~pi075 & ~pi077;
assign w384 = pi037 & w383;
assign w385 = ~w382 & ~w384;
assign w386 = w380 & w385;
assign w387 = w8 & ~w386;
assign w388 = pi138 & pi139;
assign w389 = pi119 & w388;
assign w390 = ~pi138 & ~pi139;
assign w391 = pi128 & w390;
assign w392 = ~pi072 & w28;
assign w393 = ~w391 & ~w392;
assign w394 = ~w389 & w393;
assign w395 = ~w387 & w394;
assign w396 = pi066 & ~pi113;
assign w397 = w10 & w744;
assign w398 = ~w165 & ~w169;
assign w399 = ~w170 & ~w398;
assign w400 = (~w396 & ~w399) | (~w396 & w812) | (~w399 & w812);
assign w401 = w7 & ~w400;
assign w402 = pi066 & w171;
assign w403 = w171 & w813;
assign w404 = pi025 & w378;
assign w405 = pi006 & w376;
assign w406 = ~w404 & ~w405;
assign w407 = pi032 & w383;
assign w408 = pi014 & w381;
assign w409 = ~w407 & ~w408;
assign w410 = w406 & w409;
assign w411 = pi117 & w388;
assign w412 = pi127 & w390;
assign w413 = ~w411 & ~w412;
assign w414 = (w413 & w410) | (w413 & w814) | (w410 & w814);
assign w415 = ~w403 & w414;
assign w416 = w171 & w815;
assign w417 = pi036 & w383;
assign w418 = pi013 & w381;
assign w419 = ~w417 & ~w418;
assign w420 = pi021 & w376;
assign w421 = pi024 & w378;
assign w422 = ~w420 & ~w421;
assign w423 = w419 & w422;
assign w424 = pi124 & w390;
assign w425 = pi116 & w388;
assign w426 = ~w424 & ~w425;
assign w427 = (w426 & w423) | (w426 & w816) | (w423 & w816);
assign w428 = ~w416 & w427;
assign w429 = w15 & w817;
assign w430 = pi001 & w28;
assign w431 = w429 & w430;
assign w432 = pi012 & w381;
assign w433 = pi020 & w376;
assign w434 = ~w432 & ~w433;
assign w435 = pi031 & w383;
assign w436 = pi023 & w378;
assign w437 = ~w435 & ~w436;
assign w438 = w434 & w437;
assign w439 = pi115 & w388;
assign w440 = pi126 & w390;
assign w441 = ~w439 & ~w440;
assign w442 = (w441 & w438) | (w441 & w818) | (w438 & w818);
assign w443 = ~w431 & w442;
assign w444 = pi008 & w376;
assign w445 = pi027 & w378;
assign w446 = ~w444 & ~w445;
assign w447 = pi016 & w381;
assign w448 = pi034 & w383;
assign w449 = ~w447 & ~w448;
assign w450 = w446 & w449;
assign w451 = w8 & ~w450;
assign w452 = pi122 & w390;
assign w453 = pi112 & w388;
assign w454 = ~w452 & ~w453;
assign w455 = ~w451 & w454;
assign w456 = ~pi001 & w28;
assign w457 = w429 & w456;
assign w458 = pi011 & w381;
assign w459 = pi019 & w376;
assign w460 = ~w458 & ~w459;
assign w461 = pi030 & w383;
assign w462 = pi022 & w378;
assign w463 = ~w461 & ~w462;
assign w464 = w460 & w463;
assign w465 = pi123 & w390;
assign w466 = pi114 & w388;
assign w467 = ~w465 & ~w466;
assign w468 = (w467 & w464) | (w467 & w819) | (w464 & w819);
assign w469 = ~w457 & w468;
assign w470 = (pi072 & ~w402) | (pi072 & w820) | (~w402 & w820);
assign w471 = (pi128 & ~w29) | (pi128 & w821) | (~w29 & w821);
assign w472 = ~w470 & w471;
assign w473 = pi018 & w381;
assign w474 = pi029 & w378;
assign w475 = ~w473 & ~w474;
assign w476 = pi010 & w376;
assign w477 = pi035 & w383;
assign w478 = ~w476 & ~w477;
assign w479 = w475 & w478;
assign w480 = w8 & ~w479;
assign w481 = pi120 & w388;
assign w482 = pi121 & w390;
assign w483 = pi003 & w28;
assign w484 = ~w482 & ~w483;
assign w485 = ~w481 & w484;
assign w486 = ~w480 & w485;
assign w487 = pi007 & w376;
assign w488 = pi026 & w378;
assign w489 = ~w487 & ~w488;
assign w490 = pi015 & w381;
assign w491 = pi033 & w383;
assign w492 = ~w490 & ~w491;
assign w493 = w489 & w492;
assign w494 = w8 & ~w493;
assign w495 = pi125 & w390;
assign w496 = pi118 & w388;
assign w497 = ~w495 & ~w496;
assign w498 = ~w494 & w497;
assign w499 = w11 & w378;
assign w500 = (w11 & w822) | (w11 & w823) | (w822 & w823);
assign w501 = ~w499 & w500;
assign w502 = pi113 & w210;
assign w503 = pi113 & pi129;
assign w504 = (pi128 & w503) | (pi128 & w824) | (w503 & w824);
assign w505 = ~w502 & w504;
assign w506 = ~pi077 & ~w11;
assign w507 = (pi128 & ~w11) | (pi128 & w825) | (~w11 & w825);
assign w508 = ~w506 & w507;
assign w509 = ~pi083 & w397;
assign w510 = w397 & w826;
assign w511 = (pi078 & ~w397) | (pi078 & w827) | (~w397 & w827);
assign w512 = w397 & w828;
assign w513 = ~w511 & ~w512;
assign w514 = pi083 & w397;
assign w515 = w397 & w829;
assign w516 = (pi079 & ~w397) | (pi079 & w830) | (~w397 & w830);
assign w517 = w397 & w831;
assign w518 = ~w516 & ~w517;
assign w519 = (pi080 & ~w397) | (pi080 & w832) | (~w397 & w832);
assign w520 = w397 & w833;
assign w521 = ~w519 & ~w520;
assign w522 = (pi081 & ~w397) | (pi081 & w834) | (~w397 & w834);
assign w523 = pi144 & w515;
assign w524 = ~w522 & ~w523;
assign w525 = pi082 & w514;
assign w526 = ~pi082 & ~w514;
assign w527 = pi128 & ~w526;
assign w528 = ~w525 & w527;
assign w529 = ~pi083 & ~w397;
assign w530 = pi128 & ~w514;
assign w531 = ~w529 & w530;
assign w532 = pi084 & ~w515;
assign w533 = pi140 & w515;
assign w534 = ~w532 & ~w533;
assign w535 = pi085 & ~w515;
assign w536 = pi141 & w515;
assign w537 = ~w535 & ~w536;
assign w538 = pi086 & ~w515;
assign w539 = pi142 & w515;
assign w540 = ~w538 & ~w539;
assign w541 = pi087 & ~w515;
assign w542 = pi143 & w515;
assign w543 = ~w541 & ~w542;
assign w544 = pi088 & ~w515;
assign w545 = pi145 & w515;
assign w546 = ~w544 & ~w545;
assign w547 = pi089 & ~w515;
assign w548 = pi147 & w515;
assign w549 = ~w547 & ~w548;
assign w550 = pi090 & ~w510;
assign w551 = pi141 & w510;
assign w552 = ~w550 & ~w551;
assign w553 = pi091 & ~w510;
assign w554 = pi142 & w510;
assign w555 = ~w553 & ~w554;
assign w556 = pi092 & ~w510;
assign w557 = pi143 & w510;
assign w558 = ~w556 & ~w557;
assign w559 = pi093 & ~w510;
assign w560 = pi145 & w510;
assign w561 = ~w559 & ~w560;
assign w562 = pi094 & ~w510;
assign w563 = pi146 & w510;
assign w564 = ~w562 & ~w563;
assign w565 = pi095 & ~w510;
assign w566 = pi147 & w510;
assign w567 = ~w565 & ~w566;
assign w568 = ~pi082 & w509;
assign w569 = pi096 & ~w568;
assign w570 = pi144 & w568;
assign w571 = ~w569 & ~w570;
assign w572 = pi097 & ~w525;
assign w573 = pi144 & w525;
assign w574 = ~w572 & ~w573;
assign w575 = pi098 & ~w525;
assign w576 = pi140 & w525;
assign w577 = ~w575 & ~w576;
assign w578 = pi099 & ~w568;
assign w579 = pi147 & w568;
assign w580 = ~w578 & ~w579;
assign w581 = pi100 & ~w568;
assign w582 = pi140 & w568;
assign w583 = ~w581 & ~w582;
assign w584 = pi101 & ~w568;
assign w585 = pi141 & w568;
assign w586 = ~w584 & ~w585;
assign w587 = pi102 & ~w568;
assign w588 = pi142 & w568;
assign w589 = ~w587 & ~w588;
assign w590 = pi103 & ~w568;
assign w591 = pi143 & w568;
assign w592 = ~w590 & ~w591;
assign w593 = pi104 & ~w568;
assign w594 = pi146 & w568;
assign w595 = ~w593 & ~w594;
assign w596 = pi105 & ~w568;
assign w597 = pi145 & w568;
assign w598 = ~w596 & ~w597;
assign w599 = pi106 & ~w525;
assign w600 = pi141 & w525;
assign w601 = ~w599 & ~w600;
assign w602 = pi107 & ~w525;
assign w603 = pi142 & w525;
assign w604 = ~w602 & ~w603;
assign w605 = pi108 & ~w525;
assign w606 = pi143 & w525;
assign w607 = ~w605 & ~w606;
assign w608 = pi109 & ~w525;
assign w609 = pi145 & w525;
assign w610 = ~w608 & ~w609;
assign w611 = pi110 & ~w525;
assign w612 = pi146 & w525;
assign w613 = ~w611 & ~w612;
assign w614 = pi111 & ~w525;
assign w615 = pi147 & w525;
assign w616 = ~w614 & ~w615;
assign w617 = w27 & w388;
assign w618 = pi112 & ~w617;
assign w619 = pi145 & w617;
assign w620 = ~w618 & ~w619;
assign w621 = pi114 & ~w617;
assign w622 = pi140 & w617;
assign w623 = ~w621 & ~w622;
assign w624 = pi115 & ~w617;
assign w625 = pi141 & w617;
assign w626 = ~w624 & ~w625;
assign w627 = pi116 & ~w617;
assign w628 = pi142 & w617;
assign w629 = ~w627 & ~w628;
assign w630 = pi117 & ~w617;
assign w631 = pi143 & w617;
assign w632 = ~w630 & ~w631;
assign w633 = pi118 & ~w617;
assign w634 = pi144 & w617;
assign w635 = ~w633 & ~w634;
assign w636 = pi119 & ~w617;
assign w637 = pi146 & w617;
assign w638 = ~w636 & ~w637;
assign w639 = pi120 & ~w617;
assign w640 = pi147 & w617;
assign w641 = ~w639 & ~w640;
assign w642 = w27 & w390;
assign w643 = pi121 & ~w642;
assign w644 = pi147 & w642;
assign w645 = ~w643 & ~w644;
assign w646 = pi122 & ~w642;
assign w647 = pi145 & w642;
assign w648 = ~w646 & ~w647;
assign w649 = pi123 & ~w642;
assign w650 = pi140 & w642;
assign w651 = ~w649 & ~w650;
assign w652 = pi124 & ~w642;
assign w653 = pi142 & w642;
assign w654 = ~w652 & ~w653;
assign w655 = ~pi125 & ~w642;
assign w656 = pi126 & ~w642;
assign w657 = pi141 & w642;
assign w658 = ~w656 & ~w657;
assign w659 = pi127 & ~w642;
assign w660 = pi143 & w642;
assign w661 = ~w659 & ~w660;
assign w662 = pi128 & ~w642;
assign w663 = pi146 & w642;
assign w664 = ~w662 & ~w663;
assign w665 = ~pi113 & ~pi129;
assign w666 = pi128 & ~w503;
assign w667 = ~w665 & w666;
assign w668 = ~pi130 & w9;
assign w669 = pi003 & pi121;
assign w670 = ~pi058 & ~pi055;
assign w671 = ~pi054 & ~pi061;
assign w672 = w671 & ~pi056;
assign w673 = ~pi053 & ~pi042;
assign w674 = w673 & ~pi057;
assign w675 = w673 & w693;
assign w676 = ~w166 & ~w165;
assign w677 = pi066 & pi124;
assign w678 = w173 & w694;
assign w679 = pi062 & ~pi040;
assign w680 = pi062 & w159;
assign w681 = ~pi062 & ~w172;
assign w682 = pi062 & pi049;
assign w683 = pi062 & pi051;
assign w684 = pi062 & pi045;
assign w685 = pi062 & pi046;
assign w686 = pi062 & pi047;
assign w687 = pi062 & pi048;
assign w688 = pi062 & pi137;
assign w689 = pi062 & pi050;
assign w690 = (~w689 & w312) | (~w689 & w717) | (w312 & w717);
assign w691 = ~pi115 & ~w176;
assign w692 = (~pi115 & ~w176) | (~pi115 & w718) | (~w176 & w718);
assign w693 = ~pi057 & ~pi052;
assign w694 = (w171 & w719) | (w171 & w720) | (w719 & w720);
assign w695 = w675 & ~pi064;
assign w696 = pi039 & pi062;
assign w697 = pi038 & pi124;
assign w698 = pi038 & w677;
assign w699 = ~pi127 & ~pi124;
assign w700 = ~pi127 & ~w677;
assign w701 = pi062 & ~pi038;
assign w702 = pi039 & w679;
assign w703 = pi039 & w680;
assign w704 = pi115 & ~w176;
assign w705 = (pi115 & ~w176) | (pi115 & w721) | (~w176 & w721);
assign w706 = pi053 & pi042;
assign w707 = w681 | ~w172;
assign w708 = (~w172 & w681) | (~w172 & ~pi039) | (w681 & ~pi039);
assign w709 = pi039 & w682;
assign w710 = pi039 & w683;
assign w711 = pi039 & w684;
assign w712 = pi039 & w685;
assign w713 = pi039 & w686;
assign w714 = pi039 & w687;
assign w715 = pi039 & w688;
assign w716 = ~w329 & ~w320;
assign w717 = ~w172 & ~w689;
assign w718 = ~pi064 & ~pi115;
assign w719 = pi128 & ~w697;
assign w720 = pi128 & ~w698;
assign w721 = ~pi064 & pi115;
assign w722 = w8 & ~pi136;
assign w723 = pi039 & pi038;
assign w724 = w176 & pi038;
assign w725 = w176 & ~w701;
assign w726 = ~w696 & pi040;
assign w727 = ~w702 & ~w172;
assign w728 = w703 & ~w192;
assign w729 = pi126 & w705;
assign w730 = pi126 & w704;
assign w731 = ~w702 & ~w223;
assign w732 = ~w674 & pi052;
assign w733 = pi114 & ~w176;
assign w734 = pi114 & ~w374;
assign w735 = ~w329 & w692;
assign w736 = ~w329 & w691;
assign w737 = w716 & w692;
assign w738 = w716 & w691;
assign w739 = ~w671 & pi056;
assign w740 = ~w673 & pi057;
assign w741 = w357 & w692;
assign w742 = w357 & w691;
assign w743 = pi054 & pi061;
assign w744 = w8 & pi136;
assign w745 = pi063 & pi128;
assign w746 = pi128 & pi000;
assign w747 = w18 & ~pi063;
assign w748 = ~pi128 & ~pi119;
assign w749 = w28 & pi147;
assign w750 = pi063 & ~pi003;
assign w751 = pi004 & pi128;
assign w752 = pi004 & pi006;
assign w753 = ~pi004 & pi046;
assign w754 = pi004 & pi007;
assign w755 = ~pi004 & pi047;
assign w756 = pi004 & pi008;
assign w757 = ~pi004 & pi048;
assign w758 = pi004 & pi009;
assign w759 = ~pi004 & pi049;
assign w760 = pi004 & pi010;
assign w761 = ~pi004 & pi043;
assign w762 = pi063 & pi011;
assign w763 = pi063 & pi012;
assign w764 = pi063 & pi013;
assign w765 = pi063 & pi014;
assign w766 = pi063 & pi015;
assign w767 = pi063 & pi016;
assign w768 = pi063 & pi017;
assign w769 = pi063 & pi018;
assign w770 = pi004 & pi019;
assign w771 = ~pi004 & pi050;
assign w772 = pi004 & pi020;
assign w773 = ~pi004 & pi051;
assign w774 = pi004 & pi021;
assign w775 = ~pi004 & pi045;
assign w776 = ~pi004 & pi022;
assign w777 = pi004 & pi050;
assign w778 = ~pi004 & pi023;
assign w779 = pi004 & pi051;
assign w780 = ~pi004 & pi024;
assign w781 = pi004 & pi045;
assign w782 = ~pi004 & pi025;
assign w783 = pi004 & pi046;
assign w784 = ~pi004 & pi026;
assign w785 = pi004 & pi047;
assign w786 = ~pi004 & pi027;
assign w787 = pi004 & pi048;
assign w788 = ~pi004 & pi028;
assign w789 = pi004 & pi049;
assign w790 = ~pi004 & pi029;
assign w791 = pi004 & pi043;
assign w792 = pi063 & pi030;
assign w793 = pi063 & pi031;
assign w794 = pi063 & pi032;
assign w795 = pi063 & pi033;
assign w796 = pi063 & pi034;
assign w797 = pi063 & pi035;
assign w798 = pi063 & pi036;
assign w799 = pi063 & pi037;
assign w800 = pi041 & ~pi038;
assign w801 = ~pi041 & pi127;
assign w802 = w696 & ~w163;
assign w803 = pi066 & w182;
assign w804 = w696 & w160;
assign w805 = ~w703 & w192;
assign w806 = pi123 & w705;
assign w807 = pi123 & w704;
assign w808 = w320 & w705;
assign w809 = w320 & w704;
assign w810 = pi058 & pi055;
assign w811 = pi128 & pi064;
assign w812 = ~w397 & ~w396;
assign w813 = pi066 & w28;
assign w814 = ~w8 & w413;
assign w815 = ~pi066 & w28;
assign w816 = ~w8 & w426;
assign w817 = ~w16 & ~w18;
assign w818 = ~w8 & w441;
assign w819 = ~w8 & w467;
assign w820 = ~w397 & pi072;
assign w821 = ~pi146 & pi128;
assign w822 = pi128 & pi075;
assign w823 = pi128 & ~w383;
assign w824 = pi076 & pi128;
assign w825 = ~pi077 & pi128;
assign w826 = ~pi083 & pi082;
assign w827 = ~w826 & pi078;
assign w828 = w826 & pi144;
assign w829 = pi083 & ~pi082;
assign w830 = ~w829 & pi079;
assign w831 = w829 & pi146;
assign w832 = ~w826 & pi080;
assign w833 = w826 & pi140;
assign w834 = ~w829 & pi081;
assign w835 = (~w699 & ~w700) | (~w699 & ~w171) | (~w700 & ~w171);
assign w836 = (w708 & w707) | (w708 & ~w157) | (w707 & ~w157);
assign one = 1;
assign po000 = pi071;// level 0
assign po001 = pi069;// level 0
assign po002 = pi068;// level 0
assign po003 = pi067;// level 0
assign po004 = pi074;// level 0
assign po005 = pi070;// level 0
assign po006 = pi065;// level 0
assign po007 = pi073;// level 0
assign po008 = pi130;// level 0
assign po009 = pi131;// level 0
assign po010 = pi038;// level 0
assign po011 = pi043;// level 0
assign po012 = one;// level 0
assign po013 = pi132;// level 0
assign po014 = ~w6;// level 4
assign po015 = w22;// level 6
assign po016 = w26;// level 4
assign po017 = w33;// level 4
assign po018 = pi133;// level 0
assign po019 = w37;// level 3
assign po020 = w40;// level 3
assign po021 = ~w43;// level 3
assign po022 = ~w46;// level 3
assign po023 = ~w49;// level 3
assign po024 = ~w52;// level 3
assign po025 = ~w55;// level 3
assign po026 = ~w60;// level 3
assign po027 = ~w64;// level 3
assign po028 = ~w68;// level 3
assign po029 = ~w72;// level 3
assign po030 = ~w76;// level 3
assign po031 = ~w80;// level 3
assign po032 = ~w84;// level 3
assign po033 = ~w88;// level 3
assign po034 = ~w91;// level 3
assign po035 = ~w94;// level 3
assign po036 = ~w97;// level 3
assign po037 = ~w100;// level 3
assign po038 = ~w103;// level 3
assign po039 = ~w106;// level 3
assign po040 = ~w109;// level 3
assign po041 = ~w112;// level 3
assign po042 = ~w115;// level 3
assign po043 = ~w118;// level 3
assign po044 = ~w121;// level 3
assign po045 = ~w125;// level 3
assign po046 = ~w128;// level 3
assign po047 = ~w131;// level 3
assign po048 = ~w134;// level 3
assign po049 = ~w137;// level 3
assign po050 = ~w140;// level 3
assign po051 = ~w143;// level 3
assign po052 = ~w146;// level 3
assign po053 = ~w180;// level 8
assign po054 = w186;// level 6
assign po055 = w190;// level 7
assign po056 = w196;// level 7
assign po057 = ~w205;// level 8
assign po058 = w222;// level 8
assign po059 = w226;// level 7
assign po060 = w239;// level 8
assign po061 = w252;// level 8
assign po062 = w265;// level 8
assign po063 = w278;// level 8
assign po064 = w291;// level 8
assign po065 = w304;// level 8
assign po066 = w316;// level 8
assign po067 = ~w322;// level 7
assign po068 = ~w326;// level 7
assign po069 = ~w335;// level 8
assign po070 = w340;// level 7
assign po071 = ~w346;// level 8
assign po072 = ~w350;// level 7
assign po073 = w355;// level 7
assign po074 = w360;// level 7
assign po075 = w364;// level 7
assign po076 = ~w369;// level 8
assign po077 = w372;// level 7
assign po078 = w373;// level 6
assign po079 = w375;// level 5
assign po080 = ~w395;// level 6
assign po081 = w401;// level 6
assign po082 = ~w415;// level 6
assign po083 = ~w428;// level 6
assign po084 = ~w443;// level 6
assign po085 = ~w455;// level 6
assign po086 = ~w469;// level 6
assign po087 = w472;// level 6
assign po088 = ~w486;// level 6
assign po089 = ~w498;// level 6
assign po090 = w501;// level 5
assign po091 = w505;// level 3
assign po092 = w508;// level 5
assign po093 = ~w513;// level 5
assign po094 = ~w518;// level 5
assign po095 = ~w521;// level 5
assign po096 = ~w524;// level 6
assign po097 = w528;// level 7
assign po098 = w531;// level 6
assign po099 = ~w534;// level 6
assign po100 = ~w537;// level 6
assign po101 = ~w540;// level 6
assign po102 = ~w543;// level 6
assign po103 = ~w546;// level 6
assign po104 = ~w549;// level 6
assign po105 = ~w552;// level 6
assign po106 = ~w555;// level 6
assign po107 = ~w558;// level 6
assign po108 = ~w561;// level 6
assign po109 = ~w564;// level 6
assign po110 = ~w567;// level 6
assign po111 = ~w571;// level 7
assign po112 = ~w574;// level 7
assign po113 = ~w577;// level 7
assign po114 = ~w580;// level 7
assign po115 = ~w583;// level 7
assign po116 = ~w586;// level 7
assign po117 = ~w589;// level 7
assign po118 = ~w592;// level 7
assign po119 = ~w595;// level 7
assign po120 = ~w598;// level 7
assign po121 = ~w601;// level 7
assign po122 = ~w604;// level 7
assign po123 = ~w607;// level 7
assign po124 = ~w610;// level 7
assign po125 = ~w613;// level 7
assign po126 = ~w616;// level 7
assign po127 = ~w620;// level 5
assign po128 = w183;// level 4
assign po129 = ~w623;// level 5
assign po130 = ~w626;// level 5
assign po131 = ~w629;// level 5
assign po132 = ~w632;// level 5
assign po133 = ~w635;// level 5
assign po134 = ~w638;// level 5
assign po135 = ~w641;// level 5
assign po136 = ~w645;// level 5
assign po137 = ~w648;// level 5
assign po138 = ~w651;// level 5
assign po139 = ~w654;// level 5
assign po140 = ~w655;// level 4
assign po141 = ~w658;// level 5
assign po142 = ~w661;// level 5
assign po143 = ~w664;// level 5
assign po144 = w667;// level 3
assign po145 = w668;// level 2
assign po146 = w669;// level 1
endmodule
