//Written by the Majority Logic Package Wed Apr 29 20:50:51 2015
module top (
            pi000, pi001, pi002, pi003, pi004, pi005, pi006, pi007, pi008, pi009, pi010, pi011, pi012, pi013, pi014, pi015, pi016, pi017, pi018, pi019, pi020, pi021, pi022, pi023, pi024, pi025, pi026, pi027, pi028, pi029, pi030, pi031, pi032, pi033, pi034, pi035, pi036, pi037, pi038, pi039, pi040, pi041, pi042, pi043, pi044, pi045, pi046, pi047, pi048, pi049, pi050, pi051, pi052, pi053, pi054, pi055, pi056, pi057, pi058, pi059, pi060, pi061, pi062, pi063, pi064, pi065, pi066, pi067, pi068, pi069, pi070, pi071, pi072, pi073, pi074, pi075, pi076, pi077, pi078, pi079, pi080, pi081, pi082, pi083, pi084, pi085, pi086, pi087, pi088, pi089, pi090, pi091, pi092, pi093, pi094, pi095, pi096, pi097, pi098, pi099, pi100, pi101, pi102, pi103, pi104, pi105, pi106, pi107, pi108, pi109, pi110, pi111, pi112, pi113, pi114, pi115, pi116, pi117, pi118, pi119, pi120, pi121, pi122, pi123, pi124, pi125, pi126, pi127, pi128, pi129, pi130, pi131, pi132, pi133, pi134, pi135, pi136, pi137, pi138, pi139, pi140, pi141, pi142, pi143, pi144, pi145, pi146, pi147, pi148, pi149, pi150, pi151, pi152, pi153, pi154, pi155, pi156, pi157, pi158, pi159, pi160, pi161, pi162, pi163, pi164, pi165, pi166, pi167, pi168, pi169, pi170, pi171, pi172, pi173, pi174, pi175, pi176, pi177, pi178, pi179, pi180, pi181, pi182, pi183, pi184, pi185, pi186, pi187, pi188, pi189, pi190, pi191, pi192, pi193, pi194, pi195, pi196, pi197, pi198, pi199, pi200, pi201, pi202, pi203, pi204, pi205, pi206, pi207, pi208, pi209, pi210, pi211, pi212, pi213, pi214, pi215, pi216, pi217, pi218, pi219, pi220, pi221, pi222, pi223, pi224, pi225, pi226, pi227, pi228, pi229, pi230, pi231, pi232, pi233, pi234, pi235, pi236, pi237, pi238, pi239, pi240, pi241, pi242, pi243, pi244, pi245, pi246, pi247, pi248, pi249, pi250, pi251, pi252, pi253, pi254, pi255, pi256, pi257, pi258, pi259, pi260, pi261, pi262, pi263, pi264, pi265, pi266, pi267, pi268, pi269, pi270, pi271, pi272, pi273, pi274, pi275, pi276, pi277, pi278, pi279, pi280, pi281, pi282, pi283, pi284, pi285, pi286, pi287, pi288, pi289, pi290, pi291, pi292, pi293, pi294, pi295, pi296, pi297, pi298, pi299, pi300, pi301, pi302, pi303, pi304, pi305, pi306, pi307, pi308, pi309, pi310, pi311, pi312, pi313, pi314, pi315, pi316, pi317, pi318, pi319, pi320, pi321, pi322, pi323, pi324, pi325, pi326, pi327, pi328, pi329, pi330, pi331, pi332, pi333, pi334, pi335, pi336, pi337, pi338, pi339, pi340, pi341, pi342, pi343, pi344, pi345, pi346, pi347, pi348, pi349, pi350, pi351, pi352, pi353, pi354, pi355, pi356, pi357, pi358, pi359, pi360, pi361, pi362, pi363, pi364, pi365, pi366, pi367, pi368, pi369, pi370, pi371, pi372, pi373, pi374, pi375, pi376, pi377, pi378, pi379, pi380, pi381, pi382, pi383, pi384, pi385, pi386, pi387, pi388, pi389, pi390, pi391, pi392, pi393, pi394, pi395, pi396, pi397, pi398, pi399, pi400, pi401, pi402, pi403, pi404, pi405, pi406, pi407, pi408, pi409, pi410, pi411, pi412, pi413, pi414, pi415, pi416, pi417, pi418, pi419, pi420, pi421, pi422, pi423, pi424, pi425, pi426, pi427, pi428, pi429, pi430, pi431, pi432, pi433, pi434, pi435, pi436, pi437, pi438, pi439, pi440, pi441, pi442, pi443, pi444, pi445, pi446, pi447, pi448, pi449, pi450, pi451, pi452, pi453, pi454, pi455, pi456, pi457, pi458, pi459, pi460, pi461, pi462, pi463, pi464, pi465, pi466, pi467, pi468, pi469, pi470, pi471, pi472, pi473, pi474, pi475, pi476, pi477, pi478, pi479, pi480, pi481, pi482, pi483, pi484, pi485, pi486, pi487, pi488, pi489, pi490, pi491, pi492, pi493, pi494, pi495, pi496, pi497, pi498, pi499, pi500, pi501, pi502, pi503, pi504, pi505, pi506, pi507, pi508, pi509, pi510, pi511, pi512, pi513, pi514, pi515, pi516, pi517, pi518, pi519, pi520, pi521, pi522, pi523, pi524, pi525, pi526, pi527, pi528, pi529, pi530, pi531, pi532, pi533, pi534, pi535, pi536, pi537, pi538, pi539, pi540, pi541, pi542, pi543, pi544, pi545, pi546, pi547, pi548, pi549, pi550, pi551, pi552, pi553, pi554, pi555, pi556, pi557, pi558, pi559, pi560, pi561, pi562, pi563, pi564, pi565, pi566, pi567, pi568, pi569, pi570, pi571, pi572, pi573, pi574, pi575, pi576, pi577, pi578, pi579, pi580, pi581, pi582, pi583, pi584, pi585, pi586, pi587, pi588, pi589, pi590, pi591, pi592, pi593, pi594, pi595, pi596, pi597, pi598, pi599, pi600, pi601, pi602, pi603, pi604, pi605, pi606, pi607, pi608, pi609, pi610, pi611, pi612, pi613, pi614, pi615, pi616, pi617, pi618, pi619, pi620, pi621, pi622, pi623, pi624, pi625, pi626, pi627, pi628, pi629, pi630, pi631, pi632, pi633, pi634, pi635, pi636, pi637, pi638, pi639, pi640, pi641, pi642, pi643, pi644, pi645, pi646, pi647, pi648, pi649, pi650, pi651, pi652, pi653, pi654, pi655, pi656, pi657, pi658, pi659, pi660, pi661, pi662, pi663, pi664, pi665, pi666, pi667, pi668, pi669, pi670, pi671, pi672, pi673, pi674, pi675, pi676, pi677, pi678, pi679, pi680, pi681, pi682, pi683, pi684, pi685, pi686, pi687, pi688, pi689, pi690, pi691, pi692, pi693, pi694, pi695, pi696, pi697, pi698, pi699, pi700, pi701, pi702, pi703, pi704, pi705, pi706, pi707, pi708, pi709, pi710, pi711, pi712, pi713, pi714, pi715, pi716, pi717, pi718, pi719, pi720, pi721, pi722, pi723, pi724, pi725, pi726, pi727, pi728, pi729, pi730, pi731, pi732, pi733, pi734, pi735, pi736, pi737, pi738, pi739, pi740, pi741, pi742, pi743, pi744, pi745, pi746, pi747, pi748, pi749, pi750, pi751, pi752, pi753, pi754, pi755, pi756, pi757, pi758, pi759, pi760, pi761, pi762, pi763, pi764, pi765, pi766, pi767, pi768, pi769, pi770, pi771, pi772, pi773, pi774, pi775, pi776, pi777, pi778, pi779, pi780, pi781, pi782, pi783, pi784, pi785, pi786, pi787, pi788, 
            po000, po001, po002, po003, po004, po005, po006, po007, po008, po009, po010, po011, po012, po013, po014, po015, po016, po017, po018, po019, po020, po021, po022, po023, po024, po025, po026, po027, po028, po029, po030, po031, po032, po033, po034, po035, po036, po037, po038, po039, po040, po041, po042, po043, po044, po045, po046, po047, po048, po049, po050, po051, po052, po053, po054, po055, po056, po057, po058, po059, po060, po061, po062, po063, po064, po065, po066, po067, po068, po069, po070, po071, po072, po073, po074, po075, po076, po077, po078, po079, po080, po081, po082, po083, po084, po085, po086, po087, po088, po089, po090, po091, po092, po093, po094, po095, po096, po097, po098, po099, po100, po101, po102, po103, po104, po105, po106, po107, po108, po109, po110, po111, po112, po113, po114, po115, po116, po117, po118, po119, po120, po121, po122, po123, po124, po125, po126, po127, po128, po129, po130, po131, po132, po133, po134, po135, po136, po137, po138, po139, po140, po141, po142, po143, po144, po145, po146, po147, po148, po149, po150, po151, po152, po153, po154, po155, po156, po157, po158, po159, po160, po161, po162, po163, po164, po165, po166, po167, po168, po169, po170, po171, po172, po173, po174, po175, po176, po177, po178, po179, po180, po181, po182, po183, po184, po185, po186, po187, po188, po189, po190, po191, po192, po193, po194, po195, po196, po197, po198, po199, po200, po201, po202, po203, po204, po205, po206, po207, po208, po209, po210, po211, po212, po213, po214, po215, po216, po217, po218, po219, po220, po221, po222, po223, po224, po225, po226, po227, po228, po229, po230, po231, po232, po233, po234, po235, po236, po237, po238, po239, po240, po241, po242, po243, po244, po245, po246, po247, po248, po249, po250, po251, po252, po253, po254, po255, po256, po257, po258, po259, po260, po261, po262, po263, po264, po265, po266, po267, po268, po269, po270, po271, po272, po273, po274, po275, po276, po277, po278, po279, po280, po281, po282, po283, po284, po285, po286, po287, po288, po289, po290, po291, po292, po293, po294, po295, po296, po297, po298, po299, po300, po301, po302, po303, po304, po305, po306, po307, po308, po309, po310, po311, po312, po313, po314, po315, po316, po317, po318, po319, po320, po321, po322, po323, po324, po325, po326, po327, po328, po329, po330, po331, po332, po333, po334, po335, po336, po337, po338, po339, po340, po341, po342, po343, po344, po345, po346, po347, po348, po349, po350, po351, po352, po353, po354, po355, po356, po357, po358, po359, po360, po361, po362, po363, po364, po365, po366, po367, po368, po369, po370, po371, po372, po373, po374, po375, po376, po377, po378, po379, po380, po381, po382, po383, po384, po385, po386, po387, po388, po389, po390, po391, po392, po393, po394, po395, po396, po397, po398, po399, po400, po401, po402, po403, po404, po405, po406, po407, po408, po409, po410, po411, po412, po413, po414, po415, po416, po417, po418, po419, po420, po421, po422, po423, po424, po425, po426, po427, po428, po429, po430, po431, po432, po433, po434, po435, po436, po437, po438, po439, po440, po441, po442, po443, po444, po445, po446, po447, po448, po449, po450, po451, po452, po453, po454, po455, po456, po457, po458, po459, po460, po461, po462, po463, po464, po465, po466, po467, po468, po469, po470, po471, po472, po473, po474, po475, po476, po477, po478, po479, po480, po481, po482, po483, po484, po485, po486, po487, po488, po489, po490, po491, po492, po493, po494, po495, po496, po497, po498, po499, po500, po501, po502, po503, po504, po505, po506, po507, po508, po509, po510, po511, po512, po513, po514, po515, po516, po517, po518, po519, po520, po521, po522, po523, po524, po525, po526, po527, po528, po529, po530, po531, po532, po533, po534, po535, po536, po537, po538, po539, po540, po541, po542, po543, po544, po545, po546, po547, po548, po549, po550, po551, po552, po553, po554, po555, po556, po557, po558, po559, po560, po561, po562, po563, po564, po565, po566, po567, po568, po569, po570, po571, po572, po573, po574, po575, po576, po577, po578, po579, po580, po581, po582, po583, po584, po585, po586, po587, po588, po589, po590, po591, po592, po593, po594, po595, po596, po597, po598, po599, po600, po601, po602, po603, po604, po605, po606, po607, po608, po609, po610, po611, po612, po613, po614, po615, po616, po617, po618, po619, po620, po621, po622, po623, po624, po625, po626, po627, po628, po629, po630, po631, po632, po633, po634, po635, po636, po637, po638, po639, po640, po641, po642, po643, po644, po645, po646, po647, po648, po649, po650, po651, po652, po653, po654, po655, po656, po657, po658, po659, po660, po661, po662, po663, po664, po665, po666, po667);
input pi000, pi001, pi002, pi003, pi004, pi005, pi006, pi007, pi008, pi009, pi010, pi011, pi012, pi013, pi014, pi015, pi016, pi017, pi018, pi019, pi020, pi021, pi022, pi023, pi024, pi025, pi026, pi027, pi028, pi029, pi030, pi031, pi032, pi033, pi034, pi035, pi036, pi037, pi038, pi039, pi040, pi041, pi042, pi043, pi044, pi045, pi046, pi047, pi048, pi049, pi050, pi051, pi052, pi053, pi054, pi055, pi056, pi057, pi058, pi059, pi060, pi061, pi062, pi063, pi064, pi065, pi066, pi067, pi068, pi069, pi070, pi071, pi072, pi073, pi074, pi075, pi076, pi077, pi078, pi079, pi080, pi081, pi082, pi083, pi084, pi085, pi086, pi087, pi088, pi089, pi090, pi091, pi092, pi093, pi094, pi095, pi096, pi097, pi098, pi099, pi100, pi101, pi102, pi103, pi104, pi105, pi106, pi107, pi108, pi109, pi110, pi111, pi112, pi113, pi114, pi115, pi116, pi117, pi118, pi119, pi120, pi121, pi122, pi123, pi124, pi125, pi126, pi127, pi128, pi129, pi130, pi131, pi132, pi133, pi134, pi135, pi136, pi137, pi138, pi139, pi140, pi141, pi142, pi143, pi144, pi145, pi146, pi147, pi148, pi149, pi150, pi151, pi152, pi153, pi154, pi155, pi156, pi157, pi158, pi159, pi160, pi161, pi162, pi163, pi164, pi165, pi166, pi167, pi168, pi169, pi170, pi171, pi172, pi173, pi174, pi175, pi176, pi177, pi178, pi179, pi180, pi181, pi182, pi183, pi184, pi185, pi186, pi187, pi188, pi189, pi190, pi191, pi192, pi193, pi194, pi195, pi196, pi197, pi198, pi199, pi200, pi201, pi202, pi203, pi204, pi205, pi206, pi207, pi208, pi209, pi210, pi211, pi212, pi213, pi214, pi215, pi216, pi217, pi218, pi219, pi220, pi221, pi222, pi223, pi224, pi225, pi226, pi227, pi228, pi229, pi230, pi231, pi232, pi233, pi234, pi235, pi236, pi237, pi238, pi239, pi240, pi241, pi242, pi243, pi244, pi245, pi246, pi247, pi248, pi249, pi250, pi251, pi252, pi253, pi254, pi255, pi256, pi257, pi258, pi259, pi260, pi261, pi262, pi263, pi264, pi265, pi266, pi267, pi268, pi269, pi270, pi271, pi272, pi273, pi274, pi275, pi276, pi277, pi278, pi279, pi280, pi281, pi282, pi283, pi284, pi285, pi286, pi287, pi288, pi289, pi290, pi291, pi292, pi293, pi294, pi295, pi296, pi297, pi298, pi299, pi300, pi301, pi302, pi303, pi304, pi305, pi306, pi307, pi308, pi309, pi310, pi311, pi312, pi313, pi314, pi315, pi316, pi317, pi318, pi319, pi320, pi321, pi322, pi323, pi324, pi325, pi326, pi327, pi328, pi329, pi330, pi331, pi332, pi333, pi334, pi335, pi336, pi337, pi338, pi339, pi340, pi341, pi342, pi343, pi344, pi345, pi346, pi347, pi348, pi349, pi350, pi351, pi352, pi353, pi354, pi355, pi356, pi357, pi358, pi359, pi360, pi361, pi362, pi363, pi364, pi365, pi366, pi367, pi368, pi369, pi370, pi371, pi372, pi373, pi374, pi375, pi376, pi377, pi378, pi379, pi380, pi381, pi382, pi383, pi384, pi385, pi386, pi387, pi388, pi389, pi390, pi391, pi392, pi393, pi394, pi395, pi396, pi397, pi398, pi399, pi400, pi401, pi402, pi403, pi404, pi405, pi406, pi407, pi408, pi409, pi410, pi411, pi412, pi413, pi414, pi415, pi416, pi417, pi418, pi419, pi420, pi421, pi422, pi423, pi424, pi425, pi426, pi427, pi428, pi429, pi430, pi431, pi432, pi433, pi434, pi435, pi436, pi437, pi438, pi439, pi440, pi441, pi442, pi443, pi444, pi445, pi446, pi447, pi448, pi449, pi450, pi451, pi452, pi453, pi454, pi455, pi456, pi457, pi458, pi459, pi460, pi461, pi462, pi463, pi464, pi465, pi466, pi467, pi468, pi469, pi470, pi471, pi472, pi473, pi474, pi475, pi476, pi477, pi478, pi479, pi480, pi481, pi482, pi483, pi484, pi485, pi486, pi487, pi488, pi489, pi490, pi491, pi492, pi493, pi494, pi495, pi496, pi497, pi498, pi499, pi500, pi501, pi502, pi503, pi504, pi505, pi506, pi507, pi508, pi509, pi510, pi511, pi512, pi513, pi514, pi515, pi516, pi517, pi518, pi519, pi520, pi521, pi522, pi523, pi524, pi525, pi526, pi527, pi528, pi529, pi530, pi531, pi532, pi533, pi534, pi535, pi536, pi537, pi538, pi539, pi540, pi541, pi542, pi543, pi544, pi545, pi546, pi547, pi548, pi549, pi550, pi551, pi552, pi553, pi554, pi555, pi556, pi557, pi558, pi559, pi560, pi561, pi562, pi563, pi564, pi565, pi566, pi567, pi568, pi569, pi570, pi571, pi572, pi573, pi574, pi575, pi576, pi577, pi578, pi579, pi580, pi581, pi582, pi583, pi584, pi585, pi586, pi587, pi588, pi589, pi590, pi591, pi592, pi593, pi594, pi595, pi596, pi597, pi598, pi599, pi600, pi601, pi602, pi603, pi604, pi605, pi606, pi607, pi608, pi609, pi610, pi611, pi612, pi613, pi614, pi615, pi616, pi617, pi618, pi619, pi620, pi621, pi622, pi623, pi624, pi625, pi626, pi627, pi628, pi629, pi630, pi631, pi632, pi633, pi634, pi635, pi636, pi637, pi638, pi639, pi640, pi641, pi642, pi643, pi644, pi645, pi646, pi647, pi648, pi649, pi650, pi651, pi652, pi653, pi654, pi655, pi656, pi657, pi658, pi659, pi660, pi661, pi662, pi663, pi664, pi665, pi666, pi667, pi668, pi669, pi670, pi671, pi672, pi673, pi674, pi675, pi676, pi677, pi678, pi679, pi680, pi681, pi682, pi683, pi684, pi685, pi686, pi687, pi688, pi689, pi690, pi691, pi692, pi693, pi694, pi695, pi696, pi697, pi698, pi699, pi700, pi701, pi702, pi703, pi704, pi705, pi706, pi707, pi708, pi709, pi710, pi711, pi712, pi713, pi714, pi715, pi716, pi717, pi718, pi719, pi720, pi721, pi722, pi723, pi724, pi725, pi726, pi727, pi728, pi729, pi730, pi731, pi732, pi733, pi734, pi735, pi736, pi737, pi738, pi739, pi740, pi741, pi742, pi743, pi744, pi745, pi746, pi747, pi748, pi749, pi750, pi751, pi752, pi753, pi754, pi755, pi756, pi757, pi758, pi759, pi760, pi761, pi762, pi763, pi764, pi765, pi766, pi767, pi768, pi769, pi770, pi771, pi772, pi773, pi774, pi775, pi776, pi777, pi778, pi779, pi780, pi781, pi782, pi783, pi784, pi785, pi786, pi787, pi788;
output po000, po001, po002, po003, po004, po005, po006, po007, po008, po009, po010, po011, po012, po013, po014, po015, po016, po017, po018, po019, po020, po021, po022, po023, po024, po025, po026, po027, po028, po029, po030, po031, po032, po033, po034, po035, po036, po037, po038, po039, po040, po041, po042, po043, po044, po045, po046, po047, po048, po049, po050, po051, po052, po053, po054, po055, po056, po057, po058, po059, po060, po061, po062, po063, po064, po065, po066, po067, po068, po069, po070, po071, po072, po073, po074, po075, po076, po077, po078, po079, po080, po081, po082, po083, po084, po085, po086, po087, po088, po089, po090, po091, po092, po093, po094, po095, po096, po097, po098, po099, po100, po101, po102, po103, po104, po105, po106, po107, po108, po109, po110, po111, po112, po113, po114, po115, po116, po117, po118, po119, po120, po121, po122, po123, po124, po125, po126, po127, po128, po129, po130, po131, po132, po133, po134, po135, po136, po137, po138, po139, po140, po141, po142, po143, po144, po145, po146, po147, po148, po149, po150, po151, po152, po153, po154, po155, po156, po157, po158, po159, po160, po161, po162, po163, po164, po165, po166, po167, po168, po169, po170, po171, po172, po173, po174, po175, po176, po177, po178, po179, po180, po181, po182, po183, po184, po185, po186, po187, po188, po189, po190, po191, po192, po193, po194, po195, po196, po197, po198, po199, po200, po201, po202, po203, po204, po205, po206, po207, po208, po209, po210, po211, po212, po213, po214, po215, po216, po217, po218, po219, po220, po221, po222, po223, po224, po225, po226, po227, po228, po229, po230, po231, po232, po233, po234, po235, po236, po237, po238, po239, po240, po241, po242, po243, po244, po245, po246, po247, po248, po249, po250, po251, po252, po253, po254, po255, po256, po257, po258, po259, po260, po261, po262, po263, po264, po265, po266, po267, po268, po269, po270, po271, po272, po273, po274, po275, po276, po277, po278, po279, po280, po281, po282, po283, po284, po285, po286, po287, po288, po289, po290, po291, po292, po293, po294, po295, po296, po297, po298, po299, po300, po301, po302, po303, po304, po305, po306, po307, po308, po309, po310, po311, po312, po313, po314, po315, po316, po317, po318, po319, po320, po321, po322, po323, po324, po325, po326, po327, po328, po329, po330, po331, po332, po333, po334, po335, po336, po337, po338, po339, po340, po341, po342, po343, po344, po345, po346, po347, po348, po349, po350, po351, po352, po353, po354, po355, po356, po357, po358, po359, po360, po361, po362, po363, po364, po365, po366, po367, po368, po369, po370, po371, po372, po373, po374, po375, po376, po377, po378, po379, po380, po381, po382, po383, po384, po385, po386, po387, po388, po389, po390, po391, po392, po393, po394, po395, po396, po397, po398, po399, po400, po401, po402, po403, po404, po405, po406, po407, po408, po409, po410, po411, po412, po413, po414, po415, po416, po417, po418, po419, po420, po421, po422, po423, po424, po425, po426, po427, po428, po429, po430, po431, po432, po433, po434, po435, po436, po437, po438, po439, po440, po441, po442, po443, po444, po445, po446, po447, po448, po449, po450, po451, po452, po453, po454, po455, po456, po457, po458, po459, po460, po461, po462, po463, po464, po465, po466, po467, po468, po469, po470, po471, po472, po473, po474, po475, po476, po477, po478, po479, po480, po481, po482, po483, po484, po485, po486, po487, po488, po489, po490, po491, po492, po493, po494, po495, po496, po497, po498, po499, po500, po501, po502, po503, po504, po505, po506, po507, po508, po509, po510, po511, po512, po513, po514, po515, po516, po517, po518, po519, po520, po521, po522, po523, po524, po525, po526, po527, po528, po529, po530, po531, po532, po533, po534, po535, po536, po537, po538, po539, po540, po541, po542, po543, po544, po545, po546, po547, po548, po549, po550, po551, po552, po553, po554, po555, po556, po557, po558, po559, po560, po561, po562, po563, po564, po565, po566, po567, po568, po569, po570, po571, po572, po573, po574, po575, po576, po577, po578, po579, po580, po581, po582, po583, po584, po585, po586, po587, po588, po589, po590, po591, po592, po593, po594, po595, po596, po597, po598, po599, po600, po601, po602, po603, po604, po605, po606, po607, po608, po609, po610, po611, po612, po613, po614, po615, po616, po617, po618, po619, po620, po621, po622, po623, po624, po625, po626, po627, po628, po629, po630, po631, po632, po633, po634, po635, po636, po637, po638, po639, po640, po641, po642, po643, po644, po645, po646, po647, po648, po649, po650, po651, po652, po653, po654, po655, po656, po657, po658, po659, po660, po661, po662, po663, po664, po665, po666, po667;
wire one, w0, w1, w2, w3, w4, w5, w6, w7, w8, w9, w10, w11, w12, w13, w14, w15, w16, w17, w18, w19, w20, w21, w22, w23, w24, w25, w26, w27, w28, w29, w30, w31, w32, w33, w34, w35, w36, w37, w38, w39, w40, w41, w42, w43, w44, w45, w46, w47, w48, w49, w50, w51, w52, w53, w54, w55, w56, w57, w58, w59, w60, w61, w62, w63, w64, w65, w66, w67, w68, w69, w70, w71, w72, w73, w74, w75, w76, w77, w78, w79, w80, w81, w82, w83, w84, w85, w86, w87, w88, w89, w90, w91, w92, w93, w94, w95, w96, w97, w98, w99, w100, w101, w102, w103, w104, w105, w106, w107, w108, w109, w110, w111, w112, w113, w114, w115, w116, w117, w118, w119, w120, w121, w122, w123, w124, w125, w126, w127, w128, w129, w130, w131, w132, w133, w134, w135, w136, w137, w138, w139, w140, w141, w142, w143, w144, w145, w146, w147, w148, w149, w150, w151, w152, w153, w154, w155, w156, w157, w158, w159, w160, w161, w162, w163, w164, w165, w166, w167, w168, w169, w170, w171, w172, w173, w174, w175, w176, w177, w178, w179, w180, w181, w182, w183, w184, w185, w186, w187, w188, w189, w190, w191, w192, w193, w194, w195, w196, w197, w198, w199, w200, w201, w202, w203, w204, w205, w206, w207, w208, w209, w210, w211, w212, w213, w214, w215, w216, w217, w218, w219, w220, w221, w222, w223, w224, w225, w226, w227, w228, w229, w230, w231, w232, w233, w234, w235, w236, w237, w238, w239, w240, w241, w242, w243, w244, w245, w246, w247, w248, w249, w250, w251, w252, w253, w254, w255, w256, w257, w258, w259, w260, w261, w262, w263, w264, w265, w266, w267, w268, w269, w270, w271, w272, w273, w274, w275, w276, w277, w278, w279, w280, w281, w282, w283, w284, w285, w286, w287, w288, w289, w290, w291, w292, w293, w294, w295, w296, w297, w298, w299, w300, w301, w302, w303, w304, w305, w306, w307, w308, w309, w310, w311, w312, w313, w314, w315, w316, w317, w318, w319, w320, w321, w322, w323, w324, w325, w326, w327, w328, w329, w330, w331, w332, w333, w334, w335, w336, w337, w338, w339, w340, w341, w342, w343, w344, w345, w346, w347, w348, w349, w350, w351, w352, w353, w354, w355, w356, w357, w358, w359, w360, w361, w362, w363, w364, w365, w366, w367, w368, w369, w370, w371, w372, w373, w374, w375, w376, w377, w378, w379, w380, w381, w382, w383, w384, w385, w386, w387, w388, w389, w390, w391, w392, w393, w394, w395, w396, w397, w398, w399, w400, w401, w402, w403, w404, w405, w406, w407, w408, w409, w410, w411, w412, w413, w414, w415, w416, w417, w418, w419, w420, w421, w422, w423, w424, w425, w426, w427, w428, w429, w430, w431, w432, w433, w434, w435, w436, w437, w438, w439, w440, w441, w442, w443, w444, w445, w446, w447, w448, w449, w450, w451, w452, w453, w454, w455, w456, w457, w458, w459, w460, w461, w462, w463, w464, w465, w466, w467, w468, w469, w470, w471, w472, w473, w474, w475, w476, w477, w478, w479, w480, w481, w482, w483, w484, w485, w486, w487, w488, w489, w490, w491, w492, w493, w494, w495, w496, w497, w498, w499, w500, w501, w502, w503, w504, w505, w506, w507, w508, w509, w510, w511, w512, w513, w514, w515, w516, w517, w518, w519, w520, w521, w522, w523, w524, w525, w526, w527, w528, w529, w530, w531, w532, w533, w534, w535, w536, w537, w538, w539, w540, w541, w542, w543, w544, w545, w546, w547, w548, w549, w550, w551, w552, w553, w554, w555, w556, w557, w558, w559, w560, w561, w562, w563, w564, w565, w566, w567, w568, w569, w570, w571, w572, w573, w574, w575, w576, w577, w578, w579, w580, w581, w582, w583, w584, w585, w586, w587, w588, w589, w590, w591, w592, w593, w594, w595, w596, w597, w598, w599, w600, w601, w602, w603, w604, w605, w606, w607, w608, w609, w610, w611, w612, w613, w614, w615, w616, w617, w618, w619, w620, w621, w622, w623, w624, w625, w626, w627, w628, w629, w630, w631, w632, w633, w634, w635, w636, w637, w638, w639, w640, w641, w642, w643, w644, w645, w646, w647, w648, w649, w650, w651, w652, w653, w654, w655, w656, w657, w658, w659, w660, w661, w662, w663, w664, w665, w666, w667, w668, w669, w670, w671, w672, w673, w674, w675, w676, w677, w678, w679, w680, w681, w682, w683, w684, w685, w686, w687, w688, w689, w690, w691, w692, w693, w694, w695, w696, w697, w698, w699, w700, w701, w702, w703, w704, w705, w706, w707, w708, w709, w710, w711, w712, w713, w714, w715, w716, w717, w718, w719, w720, w721, w722, w723, w724, w725, w726, w727, w728, w729, w730, w731, w732, w733, w734, w735, w736, w737, w738, w739, w740, w741, w742, w743, w744, w745, w746, w747, w748, w749, w750, w751, w752, w753, w754, w755, w756, w757, w758, w759, w760, w761, w762, w763, w764, w765, w766, w767, w768, w769, w770, w771, w772, w773, w774, w775, w776, w777, w778, w779, w780, w781, w782, w783, w784, w785, w786, w787, w788, w789, w790, w791, w792, w793, w794, w795, w796, w797, w798, w799, w800, w801, w802, w803, w804, w805, w806, w807, w808, w809, w810, w811, w812, w813, w814, w815, w816, w817, w818, w819, w820, w821, w822, w823, w824, w825, w826, w827, w828, w829, w830, w831, w832, w833, w834, w835, w836, w837, w838, w839, w840, w841, w842, w843, w844, w845, w846, w847, w848, w849, w850, w851, w852, w853, w854, w855, w856, w857, w858, w859, w860, w861, w862, w863, w864, w865, w866, w867, w868, w869, w870, w871, w872, w873, w874, w875, w876, w877, w878, w879, w880, w881, w882, w883, w884, w885, w886, w887, w888, w889, w890, w891, w892, w893, w894, w895, w896, w897, w898, w899, w900, w901, w902, w903, w904, w905, w906, w907, w908, w909, w910, w911, w912, w913, w914, w915, w916, w917, w918, w919, w920, w921, w922, w923, w924, w925, w926, w927, w928, w929, w930, w931, w932, w933, w934, w935, w936, w937, w938, w939, w940, w941, w942, w943, w944, w945, w946, w947, w948, w949, w950, w951, w952, w953, w954, w955, w956, w957, w958, w959, w960, w961, w962, w963, w964, w965, w966, w967, w968, w969, w970, w971, w972, w973, w974, w975, w976, w977, w978, w979, w980, w981, w982, w983, w984, w985, w986, w987, w988, w989, w990, w991, w992, w993, w994, w995, w996, w997, w998, w999, w1000, w1001, w1002, w1003, w1004, w1005, w1006, w1007, w1008, w1009, w1010, w1011, w1012, w1013, w1014, w1015, w1016, w1017, w1018, w1019, w1020, w1021, w1022, w1023, w1024, w1025, w1026, w1027, w1028, w1029, w1030, w1031, w1032, w1033, w1034, w1035, w1036, w1037, w1038, w1039, w1040, w1041, w1042, w1043, w1044, w1045, w1046, w1047, w1048, w1049, w1050, w1051, w1052, w1053, w1054, w1055, w1056, w1057, w1058, w1059, w1060, w1061, w1062, w1063, w1064, w1065, w1066, w1067, w1068, w1069, w1070, w1071, w1072, w1073, w1074, w1075, w1076, w1077, w1078, w1079, w1080, w1081, w1082, w1083, w1084, w1085, w1086, w1087, w1088, w1089, w1090, w1091, w1092, w1093, w1094, w1095, w1096, w1097, w1098, w1099, w1100, w1101, w1102, w1103, w1104, w1105, w1106, w1107, w1108, w1109, w1110, w1111, w1112, w1113, w1114, w1115, w1116, w1117, w1118, w1119, w1120, w1121, w1122, w1123, w1124, w1125, w1126, w1127, w1128, w1129, w1130, w1131, w1132, w1133, w1134, w1135, w1136, w1137, w1138, w1139, w1140, w1141, w1142, w1143, w1144, w1145, w1146, w1147, w1148, w1149, w1150, w1151, w1152, w1153, w1154, w1155, w1156, w1157, w1158, w1159, w1160, w1161, w1162, w1163, w1164, w1165, w1166, w1167, w1168, w1169, w1170, w1171, w1172, w1173, w1174, w1175, w1176, w1177, w1178, w1179, w1180, w1181, w1182, w1183, w1184, w1185, w1186, w1187, w1188, w1189, w1190, w1191, w1192, w1193, w1194, w1195, w1196, w1197, w1198, w1199, w1200, w1201, w1202, w1203, w1204, w1205, w1206, w1207, w1208, w1209, w1210, w1211, w1212, w1213, w1214, w1215, w1216, w1217, w1218, w1219, w1220, w1221, w1222, w1223, w1224, w1225, w1226, w1227, w1228, w1229, w1230, w1231, w1232, w1233, w1234, w1235, w1236, w1237, w1238, w1239, w1240, w1241, w1242, w1243, w1244, w1245, w1246, w1247, w1248, w1249, w1250, w1251, w1252, w1253, w1254, w1255, w1256, w1257, w1258, w1259, w1260, w1261, w1262, w1263, w1264, w1265, w1266, w1267, w1268, w1269, w1270, w1271, w1272, w1273, w1274, w1275, w1276, w1277, w1278, w1279, w1280, w1281, w1282, w1283, w1284, w1285, w1286, w1287, w1288, w1289, w1290, w1291, w1292, w1293, w1294, w1295, w1296, w1297, w1298, w1299, w1300, w1301, w1302, w1303, w1304, w1305, w1306, w1307, w1308, w1309, w1310, w1311, w1312, w1313, w1314, w1315, w1316, w1317, w1318, w1319, w1320, w1321, w1322, w1323, w1324, w1325, w1326, w1327, w1328, w1329, w1330, w1331, w1332, w1333, w1334, w1335, w1336, w1337, w1338, w1339, w1340, w1341, w1342, w1343, w1344, w1345, w1346, w1347, w1348, w1349, w1350, w1351, w1352, w1353, w1354, w1355, w1356, w1357, w1358, w1359, w1360, w1361, w1362, w1363, w1364, w1365, w1366, w1367, w1368, w1369, w1370, w1371, w1372, w1373, w1374, w1375, w1376, w1377, w1378, w1379, w1380, w1381, w1382, w1383, w1384, w1385, w1386, w1387, w1388, w1389, w1390, w1391, w1392, w1393, w1394, w1395, w1396, w1397, w1398, w1399, w1400, w1401, w1402, w1403, w1404, w1405, w1406, w1407, w1408, w1409, w1410, w1411, w1412, w1413, w1414, w1415, w1416, w1417, w1418, w1419, w1420, w1421, w1422, w1423, w1424, w1425, w1426, w1427, w1428, w1429, w1430, w1431, w1432, w1433, w1434, w1435, w1436, w1437, w1438, w1439, w1440, w1441, w1442, w1443, w1444, w1445, w1446, w1447, w1448, w1449, w1450, w1451, w1452, w1453, w1454, w1455, w1456, w1457, w1458, w1459, w1460, w1461, w1462, w1463, w1464, w1465, w1466, w1467, w1468, w1469, w1470, w1471, w1472, w1473, w1474, w1475, w1476, w1477, w1478, w1479, w1480, w1481, w1482, w1483, w1484, w1485, w1486, w1487, w1488, w1489, w1490, w1491, w1492, w1493, w1494, w1495, w1496, w1497, w1498, w1499, w1500, w1501, w1502, w1503, w1504, w1505, w1506, w1507, w1508, w1509, w1510, w1511, w1512, w1513, w1514, w1515, w1516, w1517, w1518, w1519, w1520, w1521, w1522, w1523, w1524, w1525, w1526, w1527, w1528, w1529, w1530, w1531, w1532, w1533, w1534, w1535, w1536, w1537, w1538, w1539, w1540, w1541, w1542, w1543, w1544, w1545, w1546, w1547, w1548, w1549, w1550, w1551, w1552, w1553, w1554, w1555, w1556, w1557, w1558, w1559, w1560, w1561, w1562, w1563, w1564, w1565, w1566, w1567, w1568, w1569, w1570, w1571, w1572, w1573, w1574, w1575, w1576, w1577, w1578, w1579, w1580, w1581, w1582, w1583, w1584, w1585, w1586, w1587, w1588, w1589, w1590, w1591, w1592, w1593, w1594, w1595, w1596, w1597, w1598, w1599, w1600, w1601, w1602, w1603, w1604, w1605, w1606, w1607, w1608, w1609, w1610, w1611, w1612, w1613, w1614, w1615, w1616, w1617, w1618, w1619, w1620, w1621, w1622, w1623, w1624, w1625, w1626, w1627, w1628, w1629, w1630, w1631, w1632, w1633, w1634, w1635, w1636, w1637, w1638, w1639, w1640, w1641, w1642, w1643, w1644, w1645, w1646, w1647, w1648, w1649, w1650, w1651, w1652, w1653, w1654, w1655, w1656, w1657, w1658, w1659, w1660, w1661, w1662, w1663, w1664, w1665, w1666, w1667, w1668, w1669, w1670, w1671, w1672, w1673, w1674, w1675, w1676, w1677, w1678, w1679, w1680, w1681, w1682, w1683, w1684, w1685, w1686, w1687, w1688, w1689, w1690, w1691, w1692, w1693, w1694, w1695, w1696, w1697, w1698, w1699, w1700, w1701, w1702, w1703, w1704, w1705, w1706, w1707, w1708, w1709, w1710, w1711, w1712, w1713, w1714, w1715, w1716, w1717, w1718, w1719, w1720, w1721, w1722, w1723, w1724, w1725, w1726, w1727, w1728, w1729, w1730, w1731, w1732, w1733, w1734, w1735, w1736, w1737, w1738, w1739, w1740, w1741, w1742, w1743, w1744, w1745, w1746, w1747, w1748, w1749, w1750, w1751, w1752, w1753, w1754, w1755, w1756, w1757, w1758, w1759, w1760, w1761, w1762, w1763, w1764, w1765, w1766, w1767, w1768, w1769, w1770, w1771, w1772, w1773, w1774, w1775, w1776, w1777, w1778, w1779, w1780, w1781, w1782, w1783, w1784, w1785, w1786, w1787, w1788, w1789, w1790, w1791, w1792, w1793, w1794, w1795, w1796, w1797, w1798, w1799, w1800, w1801, w1802, w1803, w1804, w1805, w1806, w1807, w1808, w1809, w1810, w1811, w1812, w1813, w1814, w1815, w1816, w1817, w1818, w1819, w1820, w1821, w1822, w1823, w1824, w1825, w1826, w1827, w1828, w1829, w1830, w1831, w1832, w1833, w1834, w1835, w1836, w1837, w1838, w1839, w1840, w1841, w1842, w1843, w1844, w1845, w1846, w1847, w1848, w1849, w1850, w1851, w1852, w1853, w1854, w1855, w1856, w1857, w1858, w1859, w1860, w1861, w1862, w1863, w1864, w1865, w1866, w1867, w1868, w1869, w1870, w1871, w1872, w1873, w1874, w1875, w1876, w1877, w1878, w1879, w1880, w1881, w1882, w1883, w1884, w1885, w1886, w1887, w1888, w1889, w1890, w1891, w1892, w1893, w1894, w1895, w1896, w1897, w1898, w1899, w1900, w1901, w1902, w1903, w1904, w1905, w1906, w1907, w1908, w1909, w1910, w1911, w1912, w1913, w1914, w1915, w1916, w1917, w1918, w1919, w1920, w1921, w1922, w1923, w1924, w1925, w1926, w1927, w1928, w1929, w1930, w1931, w1932, w1933, w1934, w1935, w1936, w1937, w1938, w1939, w1940, w1941, w1942, w1943, w1944, w1945, w1946, w1947, w1948, w1949, w1950, w1951, w1952, w1953, w1954, w1955, w1956, w1957, w1958, w1959, w1960, w1961, w1962, w1963, w1964, w1965, w1966, w1967, w1968, w1969, w1970, w1971, w1972, w1973, w1974, w1975, w1976, w1977, w1978, w1979, w1980, w1981, w1982, w1983, w1984, w1985, w1986, w1987, w1988, w1989, w1990, w1991, w1992, w1993, w1994, w1995, w1996, w1997, w1998, w1999, w2000, w2001, w2002, w2003, w2004, w2005, w2006, w2007, w2008, w2009, w2010, w2011, w2012, w2013, w2014, w2015, w2016, w2017, w2018, w2019, w2020, w2021, w2022, w2023, w2024, w2025, w2026, w2027, w2028, w2029, w2030, w2031, w2032, w2033, w2034, w2035, w2036, w2037, w2038, w2039, w2040, w2041, w2042, w2043, w2044, w2045, w2046, w2047, w2048, w2049, w2050, w2051, w2052, w2053, w2054, w2055, w2056, w2057, w2058, w2059, w2060, w2061, w2062, w2063, w2064, w2065, w2066, w2067, w2068, w2069, w2070, w2071, w2072, w2073, w2074, w2075, w2076, w2077, w2078, w2079, w2080, w2081, w2082, w2083, w2084, w2085, w2086, w2087, w2088, w2089, w2090, w2091, w2092, w2093, w2094, w2095, w2096, w2097, w2098, w2099, w2100, w2101, w2102, w2103, w2104, w2105, w2106, w2107, w2108, w2109, w2110, w2111, w2112, w2113, w2114, w2115, w2116, w2117, w2118, w2119, w2120, w2121, w2122, w2123, w2124, w2125, w2126, w2127, w2128, w2129, w2130, w2131, w2132, w2133, w2134, w2135, w2136, w2137, w2138, w2139, w2140, w2141, w2142, w2143, w2144, w2145, w2146, w2147, w2148, w2149, w2150, w2151, w2152, w2153, w2154, w2155, w2156, w2157, w2158, w2159, w2160, w2161, w2162, w2163, w2164, w2165, w2166, w2167, w2168, w2169, w2170, w2171, w2172, w2173, w2174, w2175, w2176, w2177, w2178, w2179, w2180, w2181, w2182, w2183, w2184, w2185, w2186, w2187, w2188, w2189, w2190, w2191, w2192, w2193, w2194, w2195, w2196, w2197, w2198, w2199, w2200, w2201, w2202, w2203, w2204, w2205, w2206, w2207, w2208, w2209, w2210, w2211, w2212, w2213, w2214, w2215, w2216, w2217, w2218, w2219, w2220, w2221, w2222, w2223, w2224, w2225, w2226, w2227, w2228, w2229, w2230, w2231, w2232, w2233, w2234, w2235, w2236, w2237, w2238, w2239, w2240, w2241, w2242, w2243, w2244, w2245, w2246, w2247, w2248, w2249, w2250, w2251, w2252, w2253, w2254, w2255, w2256, w2257, w2258, w2259, w2260, w2261, w2262, w2263, w2264, w2265, w2266, w2267, w2268, w2269, w2270, w2271, w2272, w2273, w2274, w2275, w2276, w2277, w2278, w2279, w2280, w2281, w2282, w2283, w2284, w2285, w2286, w2287, w2288, w2289, w2290, w2291, w2292, w2293, w2294, w2295, w2296, w2297, w2298, w2299, w2300, w2301, w2302, w2303, w2304, w2305, w2306, w2307, w2308, w2309, w2310, w2311, w2312, w2313, w2314, w2315, w2316, w2317, w2318, w2319, w2320, w2321, w2322, w2323, w2324, w2325, w2326, w2327, w2328, w2329, w2330, w2331, w2332, w2333, w2334, w2335, w2336, w2337, w2338, w2339, w2340, w2341, w2342, w2343, w2344, w2345, w2346, w2347, w2348, w2349, w2350, w2351, w2352, w2353, w2354, w2355, w2356, w2357, w2358, w2359, w2360, w2361, w2362, w2363, w2364, w2365, w2366, w2367, w2368, w2369, w2370, w2371, w2372, w2373, w2374, w2375, w2376, w2377, w2378, w2379, w2380, w2381, w2382, w2383, w2384, w2385, w2386, w2387, w2388, w2389, w2390, w2391, w2392, w2393, w2394, w2395, w2396, w2397, w2398, w2399, w2400, w2401, w2402, w2403, w2404, w2405, w2406, w2407, w2408, w2409, w2410, w2411, w2412, w2413, w2414, w2415, w2416, w2417, w2418, w2419, w2420, w2421, w2422, w2423, w2424, w2425, w2426, w2427, w2428, w2429, w2430, w2431, w2432, w2433, w2434, w2435, w2436, w2437, w2438, w2439, w2440, w2441, w2442, w2443, w2444, w2445, w2446, w2447, w2448, w2449, w2450, w2451, w2452, w2453, w2454, w2455, w2456, w2457, w2458, w2459, w2460, w2461, w2462, w2463, w2464, w2465, w2466, w2467, w2468, w2469, w2470, w2471, w2472, w2473, w2474, w2475, w2476, w2477, w2478, w2479, w2480, w2481, w2482, w2483, w2484, w2485, w2486, w2487, w2488, w2489, w2490, w2491, w2492, w2493, w2494, w2495, w2496, w2497, w2498, w2499, w2500, w2501, w2502, w2503, w2504, w2505, w2506, w2507, w2508, w2509, w2510, w2511, w2512, w2513, w2514, w2515, w2516, w2517, w2518, w2519, w2520, w2521, w2522, w2523, w2524, w2525, w2526, w2527, w2528, w2529, w2530, w2531, w2532, w2533, w2534, w2535, w2536, w2537, w2538, w2539, w2540, w2541, w2542, w2543, w2544, w2545, w2546, w2547, w2548, w2549, w2550, w2551, w2552, w2553, w2554, w2555, w2556, w2557, w2558, w2559, w2560, w2561, w2562, w2563, w2564, w2565, w2566, w2567, w2568, w2569, w2570, w2571, w2572, w2573, w2574, w2575, w2576, w2577, w2578, w2579, w2580, w2581, w2582, w2583, w2584, w2585, w2586, w2587, w2588, w2589, w2590, w2591, w2592, w2593, w2594, w2595, w2596, w2597, w2598, w2599, w2600, w2601, w2602, w2603, w2604, w2605, w2606, w2607, w2608, w2609, w2610, w2611, w2612, w2613, w2614, w2615, w2616, w2617, w2618, w2619, w2620, w2621, w2622, w2623, w2624, w2625, w2626, w2627, w2628, w2629, w2630, w2631, w2632, w2633, w2634, w2635, w2636, w2637, w2638, w2639, w2640, w2641, w2642, w2643, w2644, w2645, w2646, w2647, w2648, w2649, w2650, w2651, w2652, w2653, w2654, w2655, w2656, w2657, w2658, w2659, w2660, w2661, w2662, w2663, w2664, w2665, w2666, w2667, w2668, w2669, w2670, w2671, w2672, w2673, w2674, w2675, w2676, w2677, w2678, w2679, w2680, w2681, w2682, w2683, w2684, w2685, w2686, w2687, w2688, w2689, w2690, w2691, w2692, w2693, w2694, w2695, w2696, w2697, w2698, w2699, w2700, w2701, w2702, w2703, w2704, w2705, w2706, w2707, w2708, w2709, w2710, w2711, w2712, w2713, w2714, w2715, w2716, w2717, w2718, w2719, w2720, w2721, w2722, w2723, w2724, w2725, w2726, w2727, w2728, w2729, w2730, w2731, w2732, w2733, w2734, w2735, w2736, w2737, w2738, w2739, w2740, w2741, w2742, w2743, w2744, w2745, w2746, w2747, w2748, w2749, w2750, w2751, w2752, w2753, w2754, w2755, w2756, w2757, w2758, w2759, w2760, w2761, w2762, w2763, w2764, w2765, w2766, w2767, w2768, w2769, w2770, w2771, w2772, w2773, w2774, w2775, w2776, w2777, w2778, w2779, w2780, w2781, w2782, w2783, w2784, w2785, w2786, w2787, w2788, w2789, w2790, w2791, w2792, w2793, w2794, w2795, w2796, w2797, w2798, w2799, w2800, w2801, w2802, w2803, w2804, w2805, w2806, w2807, w2808, w2809, w2810, w2811, w2812, w2813, w2814, w2815, w2816, w2817, w2818, w2819, w2820, w2821, w2822, w2823, w2824, w2825, w2826, w2827, w2828, w2829, w2830, w2831, w2832, w2833, w2834, w2835, w2836, w2837, w2838, w2839, w2840, w2841, w2842, w2843, w2844, w2845, w2846, w2847, w2848, w2849, w2850, w2851, w2852, w2853, w2854, w2855, w2856, w2857, w2858, w2859, w2860, w2861, w2862, w2863, w2864, w2865, w2866, w2867, w2868, w2869, w2870, w2871, w2872, w2873, w2874, w2875, w2876, w2877, w2878, w2879, w2880, w2881, w2882, w2883, w2884, w2885, w2886, w2887, w2888, w2889, w2890, w2891, w2892, w2893, w2894, w2895, w2896, w2897, w2898, w2899, w2900, w2901, w2902, w2903, w2904, w2905, w2906, w2907, w2908, w2909, w2910, w2911, w2912, w2913, w2914, w2915, w2916, w2917, w2918, w2919, w2920, w2921, w2922, w2923, w2924, w2925, w2926, w2927, w2928, w2929, w2930, w2931, w2932, w2933, w2934, w2935, w2936, w2937, w2938, w2939, w2940, w2941, w2942, w2943, w2944, w2945, w2946, w2947, w2948, w2949, w2950, w2951, w2952, w2953, w2954, w2955, w2956, w2957, w2958, w2959, w2960, w2961, w2962, w2963, w2964, w2965, w2966, w2967, w2968, w2969, w2970, w2971, w2972, w2973, w2974, w2975, w2976, w2977, w2978, w2979, w2980, w2981, w2982, w2983, w2984, w2985, w2986, w2987, w2988, w2989, w2990, w2991, w2992, w2993, w2994, w2995, w2996, w2997, w2998, w2999, w3000, w3001, w3002, w3003, w3004, w3005, w3006, w3007, w3008, w3009, w3010, w3011, w3012, w3013, w3014, w3015, w3016, w3017, w3018, w3019, w3020, w3021, w3022, w3023, w3024, w3025, w3026, w3027, w3028, w3029, w3030, w3031, w3032, w3033, w3034, w3035, w3036, w3037, w3038, w3039, w3040, w3041, w3042, w3043, w3044, w3045, w3046, w3047, w3048, w3049, w3050, w3051, w3052, w3053, w3054, w3055, w3056, w3057, w3058, w3059, w3060, w3061, w3062, w3063, w3064, w3065, w3066, w3067, w3068, w3069, w3070, w3071, w3072, w3073, w3074, w3075, w3076, w3077, w3078, w3079, w3080, w3081, w3082, w3083, w3084, w3085, w3086, w3087, w3088, w3089, w3090, w3091, w3092, w3093, w3094, w3095, w3096, w3097, w3098, w3099, w3100, w3101, w3102, w3103, w3104, w3105, w3106, w3107, w3108, w3109, w3110, w3111, w3112, w3113, w3114, w3115, w3116, w3117, w3118, w3119, w3120, w3121, w3122, w3123, w3124, w3125, w3126, w3127, w3128, w3129, w3130, w3131, w3132, w3133, w3134, w3135, w3136, w3137, w3138, w3139, w3140, w3141, w3142, w3143, w3144, w3145, w3146, w3147, w3148, w3149, w3150, w3151, w3152, w3153, w3154, w3155, w3156, w3157, w3158, w3159, w3160, w3161, w3162, w3163, w3164, w3165, w3166, w3167, w3168, w3169, w3170, w3171, w3172, w3173, w3174, w3175, w3176, w3177, w3178, w3179, w3180, w3181, w3182, w3183, w3184, w3185, w3186, w3187, w3188, w3189, w3190, w3191, w3192, w3193, w3194, w3195, w3196, w3197, w3198, w3199, w3200, w3201, w3202, w3203, w3204, w3205, w3206, w3207, w3208, w3209, w3210, w3211, w3212, w3213, w3214, w3215, w3216, w3217, w3218, w3219, w3220, w3221, w3222, w3223, w3224, w3225, w3226, w3227, w3228, w3229, w3230, w3231, w3232, w3233, w3234, w3235, w3236, w3237, w3238, w3239, w3240, w3241, w3242, w3243, w3244, w3245, w3246, w3247, w3248, w3249, w3250, w3251, w3252, w3253, w3254, w3255, w3256, w3257, w3258, w3259, w3260, w3261, w3262, w3263, w3264, w3265, w3266, w3267, w3268, w3269, w3270, w3271, w3272, w3273, w3274, w3275, w3276, w3277, w3278, w3279, w3280, w3281, w3282, w3283, w3284, w3285, w3286, w3287, w3288, w3289, w3290, w3291, w3292, w3293, w3294, w3295, w3296, w3297, w3298, w3299, w3300, w3301, w3302, w3303, w3304, w3305, w3306, w3307, w3308, w3309, w3310, w3311, w3312, w3313, w3314, w3315, w3316, w3317, w3318, w3319, w3320, w3321, w3322, w3323, w3324, w3325, w3326, w3327, w3328, w3329, w3330, w3331, w3332, w3333, w3334, w3335, w3336, w3337, w3338, w3339, w3340, w3341, w3342, w3343, w3344, w3345, w3346, w3347, w3348, w3349, w3350, w3351, w3352, w3353, w3354, w3355, w3356, w3357, w3358, w3359, w3360, w3361, w3362, w3363, w3364, w3365, w3366, w3367, w3368, w3369, w3370, w3371, w3372, w3373, w3374, w3375, w3376, w3377, w3378, w3379, w3380, w3381, w3382, w3383, w3384, w3385, w3386, w3387, w3388, w3389, w3390, w3391, w3392, w3393, w3394, w3395, w3396, w3397, w3398, w3399, w3400, w3401, w3402, w3403, w3404, w3405, w3406, w3407, w3408, w3409, w3410, w3411, w3412, w3413, w3414, w3415, w3416, w3417, w3418, w3419, w3420, w3421, w3422, w3423, w3424, w3425, w3426, w3427, w3428, w3429, w3430, w3431, w3432, w3433, w3434, w3435, w3436, w3437, w3438, w3439, w3440, w3441, w3442, w3443, w3444, w3445, w3446, w3447, w3448, w3449, w3450, w3451, w3452, w3453, w3454, w3455, w3456, w3457, w3458, w3459, w3460, w3461, w3462, w3463, w3464, w3465, w3466, w3467, w3468, w3469, w3470, w3471, w3472, w3473, w3474, w3475, w3476, w3477, w3478, w3479, w3480, w3481, w3482, w3483, w3484, w3485, w3486, w3487, w3488, w3489, w3490, w3491, w3492, w3493, w3494, w3495, w3496, w3497, w3498, w3499, w3500, w3501, w3502, w3503, w3504, w3505, w3506, w3507, w3508, w3509, w3510, w3511, w3512, w3513, w3514, w3515, w3516, w3517, w3518, w3519, w3520, w3521, w3522, w3523, w3524, w3525, w3526, w3527, w3528, w3529, w3530, w3531, w3532, w3533, w3534, w3535, w3536, w3537, w3538, w3539, w3540, w3541, w3542, w3543, w3544, w3545, w3546, w3547, w3548, w3549, w3550, w3551, w3552, w3553, w3554, w3555, w3556, w3557, w3558, w3559, w3560, w3561, w3562, w3563, w3564, w3565, w3566, w3567, w3568, w3569, w3570, w3571, w3572, w3573, w3574, w3575, w3576, w3577, w3578, w3579, w3580, w3581, w3582, w3583, w3584, w3585, w3586, w3587, w3588, w3589, w3590, w3591, w3592, w3593, w3594, w3595, w3596, w3597, w3598, w3599, w3600, w3601, w3602, w3603, w3604, w3605, w3606, w3607, w3608, w3609, w3610, w3611, w3612, w3613, w3614, w3615, w3616, w3617, w3618, w3619, w3620, w3621, w3622, w3623, w3624, w3625, w3626, w3627, w3628, w3629, w3630, w3631, w3632, w3633, w3634, w3635, w3636, w3637, w3638, w3639, w3640, w3641, w3642, w3643, w3644, w3645, w3646, w3647, w3648, w3649, w3650, w3651, w3652, w3653, w3654, w3655, w3656, w3657, w3658, w3659, w3660, w3661, w3662, w3663, w3664, w3665, w3666, w3667, w3668, w3669, w3670, w3671, w3672, w3673, w3674, w3675, w3676, w3677, w3678, w3679, w3680, w3681, w3682, w3683, w3684, w3685, w3686, w3687, w3688, w3689, w3690, w3691, w3692, w3693, w3694, w3695, w3696, w3697, w3698, w3699, w3700, w3701, w3702, w3703, w3704, w3705, w3706, w3707, w3708, w3709, w3710, w3711, w3712, w3713, w3714, w3715, w3716, w3717, w3718, w3719, w3720, w3721, w3722, w3723, w3724, w3725, w3726, w3727, w3728, w3729, w3730, w3731, w3732, w3733, w3734, w3735, w3736, w3737, w3738, w3739, w3740, w3741, w3742, w3743, w3744, w3745, w3746, w3747, w3748, w3749, w3750, w3751, w3752, w3753, w3754, w3755, w3756, w3757, w3758, w3759, w3760, w3761, w3762, w3763, w3764, w3765, w3766, w3767, w3768, w3769, w3770, w3771, w3772, w3773, w3774, w3775, w3776, w3777, w3778, w3779, w3780, w3781, w3782, w3783, w3784, w3785, w3786, w3787, w3788, w3789, w3790, w3791, w3792, w3793, w3794, w3795, w3796, w3797, w3798, w3799, w3800, w3801, w3802, w3803, w3804, w3805, w3806, w3807, w3808, w3809, w3810, w3811, w3812, w3813, w3814, w3815, w3816, w3817, w3818, w3819, w3820, w3821, w3822, w3823, w3824, w3825, w3826, w3827, w3828, w3829, w3830, w3831, w3832, w3833, w3834, w3835, w3836, w3837, w3838, w3839, w3840, w3841, w3842, w3843, w3844, w3845, w3846, w3847, w3848, w3849, w3850, w3851, w3852, w3853, w3854, w3855, w3856, w3857, w3858, w3859, w3860, w3861, w3862, w3863, w3864, w3865, w3866, w3867, w3868, w3869, w3870, w3871, w3872, w3873, w3874, w3875, w3876, w3877, w3878, w3879, w3880, w3881, w3882, w3883, w3884, w3885, w3886, w3887, w3888, w3889, w3890, w3891, w3892, w3893, w3894, w3895, w3896, w3897, w3898, w3899, w3900, w3901, w3902, w3903, w3904, w3905, w3906, w3907, w3908, w3909, w3910, w3911, w3912, w3913, w3914, w3915, w3916, w3917, w3918, w3919, w3920, w3921, w3922, w3923, w3924, w3925, w3926, w3927, w3928, w3929, w3930, w3931, w3932, w3933, w3934, w3935, w3936, w3937, w3938, w3939, w3940, w3941, w3942, w3943, w3944, w3945, w3946, w3947, w3948, w3949, w3950, w3951, w3952, w3953, w3954, w3955, w3956, w3957, w3958, w3959, w3960, w3961, w3962, w3963, w3964, w3965, w3966, w3967, w3968, w3969, w3970, w3971, w3972, w3973, w3974, w3975, w3976, w3977, w3978, w3979, w3980, w3981, w3982, w3983, w3984, w3985, w3986, w3987, w3988, w3989, w3990, w3991, w3992, w3993, w3994, w3995, w3996, w3997, w3998, w3999, w4000, w4001, w4002, w4003, w4004, w4005, w4006, w4007, w4008, w4009, w4010, w4011, w4012, w4013, w4014, w4015, w4016, w4017, w4018, w4019, w4020, w4021, w4022, w4023, w4024, w4025, w4026, w4027, w4028, w4029, w4030, w4031, w4032, w4033, w4034, w4035, w4036, w4037, w4038, w4039, w4040, w4041, w4042, w4043, w4044, w4045, w4046, w4047, w4048, w4049, w4050, w4051, w4052, w4053, w4054, w4055, w4056, w4057, w4058, w4059, w4060, w4061, w4062, w4063, w4064, w4065, w4066, w4067, w4068, w4069, w4070, w4071, w4072, w4073, w4074, w4075, w4076, w4077, w4078, w4079, w4080, w4081, w4082, w4083, w4084, w4085, w4086, w4087, w4088, w4089, w4090, w4091, w4092, w4093, w4094, w4095, w4096, w4097, w4098, w4099, w4100, w4101, w4102, w4103, w4104, w4105, w4106, w4107, w4108, w4109, w4110, w4111, w4112, w4113, w4114, w4115, w4116, w4117, w4118, w4119, w4120, w4121, w4122, w4123, w4124, w4125, w4126, w4127, w4128, w4129, w4130, w4131, w4132, w4133, w4134, w4135, w4136, w4137, w4138, w4139, w4140, w4141, w4142, w4143, w4144, w4145, w4146, w4147, w4148, w4149, w4150, w4151, w4152, w4153, w4154, w4155, w4156, w4157, w4158, w4159, w4160, w4161, w4162, w4163, w4164, w4165, w4166, w4167, w4168, w4169, w4170, w4171, w4172, w4173, w4174, w4175, w4176, w4177, w4178, w4179, w4180, w4181, w4182, w4183, w4184, w4185, w4186, w4187, w4188, w4189, w4190, w4191, w4192, w4193, w4194, w4195, w4196, w4197, w4198, w4199, w4200, w4201, w4202, w4203, w4204, w4205, w4206, w4207, w4208, w4209, w4210, w4211, w4212, w4213, w4214, w4215, w4216, w4217, w4218, w4219, w4220, w4221, w4222, w4223, w4224, w4225, w4226, w4227, w4228, w4229, w4230, w4231, w4232, w4233, w4234, w4235, w4236, w4237, w4238, w4239, w4240, w4241, w4242, w4243, w4244, w4245, w4246, w4247, w4248, w4249, w4250, w4251, w4252, w4253, w4254, w4255, w4256, w4257, w4258, w4259, w4260, w4261, w4262, w4263, w4264, w4265, w4266, w4267, w4268, w4269, w4270, w4271, w4272, w4273, w4274, w4275, w4276, w4277, w4278, w4279, w4280, w4281, w4282, w4283, w4284, w4285, w4286, w4287, w4288, w4289, w4290, w4291, w4292, w4293, w4294, w4295, w4296, w4297, w4298, w4299, w4300, w4301, w4302, w4303, w4304, w4305, w4306, w4307, w4308, w4309, w4310, w4311, w4312, w4313, w4314, w4315, w4316, w4317, w4318, w4319, w4320, w4321, w4322, w4323, w4324, w4325, w4326, w4327, w4328, w4329, w4330, w4331, w4332, w4333, w4334, w4335, w4336, w4337, w4338, w4339, w4340, w4341, w4342, w4343, w4344, w4345, w4346, w4347, w4348, w4349, w4350, w4351, w4352, w4353, w4354, w4355, w4356, w4357, w4358, w4359, w4360, w4361, w4362, w4363, w4364, w4365, w4366, w4367, w4368, w4369, w4370, w4371, w4372, w4373, w4374, w4375, w4376, w4377, w4378, w4379, w4380, w4381, w4382, w4383, w4384, w4385, w4386, w4387, w4388, w4389, w4390, w4391, w4392, w4393, w4394, w4395, w4396, w4397, w4398, w4399, w4400, w4401, w4402, w4403, w4404, w4405, w4406, w4407, w4408, w4409, w4410, w4411, w4412, w4413, w4414, w4415, w4416, w4417, w4418, w4419, w4420, w4421, w4422, w4423, w4424, w4425, w4426, w4427, w4428, w4429, w4430, w4431, w4432, w4433, w4434, w4435, w4436, w4437, w4438, w4439, w4440, w4441, w4442, w4443, w4444, w4445, w4446, w4447, w4448, w4449, w4450, w4451, w4452, w4453, w4454, w4455, w4456, w4457, w4458, w4459, w4460, w4461, w4462, w4463, w4464, w4465, w4466, w4467, w4468, w4469, w4470, w4471, w4472, w4473, w4474, w4475, w4476, w4477, w4478, w4479, w4480, w4481, w4482, w4483, w4484, w4485, w4486, w4487, w4488, w4489, w4490, w4491, w4492, w4493, w4494, w4495, w4496, w4497, w4498, w4499, w4500, w4501, w4502, w4503, w4504, w4505, w4506, w4507, w4508, w4509, w4510, w4511, w4512, w4513, w4514, w4515, w4516, w4517, w4518, w4519, w4520, w4521, w4522, w4523, w4524, w4525, w4526, w4527, w4528, w4529, w4530, w4531, w4532, w4533, w4534, w4535, w4536, w4537, w4538, w4539, w4540, w4541, w4542, w4543, w4544, w4545, w4546, w4547, w4548, w4549, w4550, w4551, w4552, w4553, w4554, w4555, w4556, w4557, w4558, w4559, w4560, w4561, w4562, w4563, w4564, w4565, w4566, w4567, w4568, w4569, w4570, w4571, w4572, w4573, w4574, w4575, w4576, w4577, w4578, w4579, w4580, w4581, w4582, w4583, w4584, w4585, w4586, w4587, w4588, w4589, w4590, w4591, w4592, w4593, w4594, w4595, w4596, w4597, w4598, w4599, w4600, w4601, w4602, w4603, w4604, w4605, w4606, w4607, w4608, w4609, w4610, w4611, w4612, w4613, w4614, w4615, w4616, w4617, w4618, w4619, w4620, w4621, w4622, w4623, w4624, w4625, w4626, w4627, w4628, w4629, w4630, w4631, w4632, w4633, w4634, w4635, w4636, w4637, w4638, w4639, w4640, w4641, w4642, w4643, w4644, w4645, w4646, w4647, w4648, w4649, w4650, w4651, w4652, w4653, w4654, w4655, w4656, w4657, w4658, w4659, w4660, w4661, w4662, w4663, w4664, w4665, w4666, w4667, w4668, w4669, w4670, w4671, w4672, w4673, w4674, w4675, w4676, w4677, w4678, w4679, w4680, w4681, w4682, w4683, w4684, w4685, w4686, w4687, w4688, w4689, w4690, w4691, w4692, w4693, w4694, w4695, w4696, w4697, w4698, w4699, w4700, w4701, w4702, w4703, w4704, w4705, w4706, w4707, w4708, w4709, w4710, w4711, w4712, w4713, w4714, w4715, w4716, w4717, w4718, w4719, w4720, w4721, w4722, w4723, w4724, w4725, w4726, w4727, w4728, w4729, w4730, w4731, w4732, w4733, w4734, w4735, w4736, w4737, w4738, w4739, w4740, w4741, w4742, w4743, w4744, w4745, w4746, w4747, w4748, w4749, w4750, w4751, w4752, w4753, w4754, w4755, w4756, w4757, w4758, w4759, w4760, w4761, w4762, w4763, w4764, w4765, w4766, w4767, w4768, w4769, w4770, w4771, w4772, w4773, w4774, w4775, w4776, w4777, w4778, w4779, w4780, w4781, w4782, w4783, w4784, w4785, w4786, w4787, w4788, w4789, w4790, w4791, w4792, w4793, w4794, w4795, w4796, w4797, w4798, w4799, w4800, w4801, w4802, w4803, w4804, w4805, w4806, w4807, w4808, w4809, w4810, w4811, w4812, w4813, w4814, w4815, w4816, w4817, w4818, w4819, w4820, w4821, w4822, w4823, w4824, w4825, w4826, w4827, w4828, w4829, w4830, w4831, w4832, w4833, w4834, w4835, w4836, w4837, w4838, w4839, w4840, w4841, w4842, w4843, w4844, w4845, w4846, w4847, w4848, w4849, w4850, w4851, w4852, w4853, w4854, w4855, w4856, w4857, w4858, w4859, w4860, w4861, w4862, w4863, w4864, w4865, w4866, w4867, w4868, w4869, w4870, w4871, w4872, w4873, w4874, w4875, w4876, w4877, w4878, w4879, w4880, w4881, w4882, w4883, w4884, w4885, w4886, w4887, w4888, w4889, w4890, w4891, w4892, w4893, w4894, w4895, w4896, w4897, w4898, w4899, w4900, w4901, w4902, w4903, w4904, w4905, w4906, w4907, w4908, w4909, w4910, w4911, w4912, w4913, w4914, w4915, w4916, w4917, w4918, w4919, w4920, w4921, w4922, w4923, w4924, w4925, w4926, w4927, w4928, w4929, w4930, w4931, w4932, w4933, w4934, w4935, w4936, w4937, w4938, w4939, w4940, w4941, w4942, w4943, w4944, w4945, w4946, w4947, w4948, w4949, w4950, w4951, w4952, w4953, w4954, w4955, w4956, w4957, w4958, w4959, w4960, w4961, w4962, w4963, w4964, w4965, w4966, w4967, w4968, w4969, w4970, w4971, w4972, w4973, w4974, w4975, w4976, w4977, w4978, w4979, w4980, w4981, w4982, w4983, w4984, w4985, w4986, w4987, w4988, w4989, w4990, w4991, w4992, w4993, w4994, w4995, w4996, w4997, w4998, w4999, w5000, w5001, w5002, w5003, w5004, w5005, w5006, w5007, w5008, w5009, w5010, w5011, w5012, w5013, w5014, w5015, w5016, w5017, w5018, w5019, w5020, w5021, w5022, w5023, w5024, w5025, w5026, w5027, w5028, w5029, w5030, w5031, w5032, w5033, w5034, w5035, w5036, w5037, w5038, w5039, w5040, w5041, w5042, w5043, w5044, w5045, w5046, w5047, w5048, w5049, w5050, w5051, w5052, w5053, w5054, w5055, w5056, w5057, w5058, w5059, w5060, w5061, w5062, w5063, w5064, w5065, w5066, w5067, w5068, w5069, w5070, w5071, w5072, w5073, w5074, w5075, w5076, w5077, w5078, w5079, w5080, w5081, w5082, w5083, w5084, w5085, w5086, w5087, w5088, w5089, w5090, w5091, w5092, w5093, w5094, w5095, w5096, w5097, w5098, w5099, w5100, w5101, w5102, w5103, w5104, w5105, w5106, w5107, w5108, w5109, w5110, w5111, w5112, w5113, w5114, w5115, w5116, w5117, w5118, w5119, w5120, w5121, w5122, w5123, w5124, w5125, w5126, w5127, w5128, w5129, w5130, w5131, w5132, w5133, w5134, w5135, w5136, w5137, w5138, w5139, w5140, w5141, w5142, w5143, w5144, w5145, w5146, w5147, w5148, w5149, w5150, w5151, w5152, w5153, w5154, w5155, w5156, w5157, w5158, w5159, w5160, w5161, w5162, w5163, w5164, w5165, w5166, w5167, w5168, w5169, w5170, w5171, w5172, w5173, w5174, w5175, w5176, w5177, w5178, w5179, w5180, w5181, w5182, w5183, w5184, w5185, w5186, w5187, w5188, w5189, w5190, w5191, w5192, w5193, w5194, w5195, w5196, w5197, w5198, w5199, w5200, w5201, w5202, w5203, w5204, w5205, w5206, w5207, w5208, w5209, w5210, w5211, w5212, w5213, w5214, w5215, w5216, w5217, w5218, w5219, w5220, w5221, w5222, w5223, w5224, w5225, w5226, w5227, w5228, w5229, w5230, w5231, w5232, w5233, w5234, w5235, w5236, w5237, w5238, w5239, w5240, w5241, w5242, w5243, w5244, w5245, w5246, w5247, w5248, w5249, w5250, w5251, w5252, w5253, w5254, w5255, w5256, w5257, w5258, w5259, w5260, w5261, w5262, w5263, w5264, w5265, w5266, w5267, w5268, w5269, w5270, w5271, w5272, w5273, w5274, w5275, w5276, w5277, w5278, w5279, w5280, w5281, w5282, w5283, w5284, w5285, w5286, w5287, w5288, w5289, w5290, w5291, w5292, w5293, w5294, w5295, w5296, w5297, w5298, w5299, w5300, w5301, w5302, w5303, w5304, w5305, w5306, w5307, w5308, w5309, w5310, w5311, w5312, w5313, w5314, w5315, w5316, w5317, w5318, w5319, w5320, w5321, w5322, w5323, w5324, w5325, w5326, w5327, w5328, w5329, w5330, w5331, w5332, w5333, w5334, w5335, w5336, w5337, w5338, w5339, w5340, w5341, w5342, w5343, w5344, w5345, w5346, w5347, w5348, w5349, w5350, w5351, w5352, w5353, w5354, w5355, w5356, w5357, w5358, w5359, w5360, w5361, w5362, w5363, w5364, w5365, w5366, w5367, w5368, w5369, w5370, w5371, w5372, w5373, w5374, w5375, w5376, w5377, w5378, w5379, w5380, w5381, w5382, w5383, w5384, w5385, w5386, w5387, w5388, w5389, w5390, w5391, w5392, w5393, w5394, w5395, w5396, w5397, w5398, w5399, w5400, w5401, w5402, w5403, w5404, w5405, w5406, w5407, w5408, w5409, w5410, w5411, w5412, w5413, w5414, w5415, w5416, w5417, w5418, w5419, w5420, w5421, w5422, w5423, w5424, w5425, w5426, w5427, w5428, w5429, w5430, w5431, w5432, w5433, w5434, w5435, w5436, w5437, w5438, w5439, w5440, w5441, w5442, w5443, w5444, w5445, w5446, w5447, w5448, w5449, w5450, w5451, w5452, w5453, w5454, w5455, w5456, w5457, w5458, w5459, w5460, w5461, w5462, w5463, w5464, w5465, w5466, w5467, w5468, w5469, w5470, w5471, w5472, w5473, w5474, w5475, w5476, w5477, w5478, w5479, w5480, w5481, w5482, w5483, w5484, w5485, w5486, w5487, w5488, w5489, w5490, w5491, w5492, w5493, w5494, w5495, w5496, w5497, w5498, w5499, w5500, w5501, w5502, w5503, w5504, w5505, w5506, w5507, w5508, w5509, w5510, w5511, w5512, w5513, w5514, w5515, w5516, w5517, w5518, w5519, w5520, w5521, w5522, w5523, w5524, w5525, w5526, w5527, w5528, w5529, w5530, w5531, w5532, w5533, w5534, w5535, w5536, w5537, w5538, w5539, w5540, w5541, w5542, w5543, w5544, w5545, w5546, w5547, w5548, w5549, w5550, w5551, w5552, w5553, w5554, w5555, w5556, w5557, w5558, w5559, w5560, w5561, w5562, w5563, w5564, w5565, w5566, w5567, w5568, w5569, w5570, w5571, w5572, w5573, w5574, w5575, w5576, w5577, w5578, w5579, w5580, w5581, w5582, w5583, w5584, w5585, w5586, w5587, w5588, w5589, w5590, w5591, w5592, w5593, w5594, w5595, w5596, w5597, w5598, w5599, w5600, w5601, w5602, w5603, w5604, w5605, w5606, w5607, w5608, w5609, w5610, w5611, w5612, w5613, w5614, w5615, w5616, w5617, w5618, w5619, w5620, w5621, w5622, w5623, w5624, w5625, w5626, w5627, w5628, w5629, w5630, w5631, w5632, w5633, w5634, w5635, w5636, w5637, w5638, w5639, w5640, w5641, w5642, w5643, w5644, w5645, w5646, w5647, w5648, w5649, w5650, w5651, w5652, w5653, w5654, w5655, w5656, w5657, w5658, w5659, w5660, w5661, w5662, w5663, w5664, w5665, w5666, w5667, w5668, w5669, w5670, w5671, w5672, w5673, w5674, w5675, w5676, w5677, w5678, w5679, w5680, w5681, w5682, w5683, w5684, w5685, w5686, w5687, w5688, w5689, w5690, w5691, w5692, w5693, w5694, w5695, w5696, w5697, w5698, w5699, w5700, w5701, w5702, w5703, w5704, w5705, w5706, w5707, w5708, w5709, w5710, w5711, w5712, w5713, w5714, w5715, w5716, w5717, w5718, w5719, w5720, w5721, w5722, w5723, w5724, w5725, w5726, w5727, w5728, w5729, w5730, w5731, w5732, w5733, w5734, w5735, w5736, w5737, w5738, w5739, w5740, w5741, w5742, w5743, w5744, w5745, w5746, w5747, w5748, w5749, w5750, w5751, w5752, w5753, w5754, w5755, w5756, w5757, w5758, w5759, w5760, w5761, w5762, w5763, w5764, w5765, w5766, w5767, w5768, w5769, w5770, w5771, w5772, w5773, w5774, w5775, w5776, w5777, w5778, w5779, w5780, w5781, w5782, w5783, w5784, w5785, w5786, w5787, w5788, w5789, w5790, w5791, w5792, w5793, w5794, w5795, w5796, w5797, w5798, w5799, w5800, w5801, w5802, w5803, w5804, w5805, w5806, w5807, w5808, w5809, w5810, w5811, w5812, w5813, w5814, w5815, w5816, w5817, w5818, w5819, w5820, w5821, w5822, w5823, w5824, w5825, w5826, w5827, w5828, w5829, w5830, w5831, w5832, w5833, w5834, w5835, w5836, w5837, w5838, w5839, w5840, w5841, w5842, w5843, w5844, w5845, w5846, w5847, w5848, w5849, w5850, w5851, w5852, w5853, w5854, w5855, w5856, w5857, w5858, w5859, w5860, w5861, w5862, w5863, w5864, w5865, w5866, w5867, w5868, w5869, w5870, w5871, w5872, w5873, w5874, w5875, w5876, w5877, w5878, w5879, w5880, w5881, w5882, w5883, w5884, w5885, w5886, w5887, w5888, w5889, w5890, w5891, w5892, w5893, w5894, w5895, w5896, w5897, w5898, w5899, w5900, w5901, w5902, w5903, w5904, w5905, w5906, w5907, w5908, w5909, w5910, w5911, w5912, w5913, w5914, w5915, w5916, w5917, w5918, w5919, w5920, w5921, w5922, w5923, w5924, w5925, w5926, w5927, w5928, w5929, w5930, w5931, w5932, w5933, w5934, w5935, w5936, w5937, w5938, w5939, w5940, w5941, w5942, w5943, w5944, w5945, w5946, w5947, w5948, w5949, w5950, w5951, w5952, w5953, w5954, w5955, w5956, w5957, w5958, w5959, w5960, w5961, w5962, w5963, w5964, w5965, w5966, w5967, w5968, w5969, w5970, w5971, w5972, w5973, w5974, w5975, w5976, w5977, w5978, w5979, w5980, w5981, w5982, w5983, w5984, w5985, w5986, w5987, w5988, w5989, w5990, w5991, w5992, w5993, w5994, w5995, w5996, w5997, w5998, w5999, w6000, w6001, w6002, w6003, w6004, w6005, w6006, w6007, w6008, w6009, w6010, w6011, w6012, w6013, w6014, w6015, w6016, w6017, w6018, w6019, w6020, w6021, w6022, w6023, w6024, w6025, w6026, w6027, w6028, w6029, w6030, w6031, w6032, w6033, w6034, w6035, w6036, w6037, w6038, w6039, w6040, w6041, w6042, w6043, w6044, w6045, w6046, w6047, w6048, w6049, w6050, w6051, w6052, w6053, w6054, w6055, w6056, w6057, w6058, w6059, w6060, w6061, w6062, w6063, w6064, w6065, w6066, w6067, w6068, w6069, w6070, w6071, w6072, w6073, w6074, w6075, w6076, w6077, w6078, w6079, w6080, w6081, w6082, w6083, w6084, w6085, w6086, w6087, w6088, w6089, w6090, w6091, w6092, w6093, w6094, w6095, w6096, w6097, w6098, w6099, w6100, w6101, w6102, w6103, w6104, w6105, w6106, w6107, w6108, w6109, w6110, w6111, w6112, w6113, w6114, w6115, w6116, w6117, w6118, w6119, w6120, w6121, w6122, w6123, w6124, w6125, w6126, w6127, w6128, w6129, w6130, w6131, w6132, w6133, w6134, w6135, w6136, w6137, w6138, w6139, w6140, w6141, w6142, w6143, w6144, w6145, w6146, w6147, w6148, w6149, w6150, w6151, w6152, w6153, w6154, w6155, w6156, w6157, w6158, w6159, w6160, w6161, w6162, w6163, w6164, w6165, w6166, w6167, w6168, w6169, w6170, w6171, w6172, w6173, w6174, w6175, w6176, w6177, w6178, w6179, w6180, w6181, w6182, w6183, w6184, w6185, w6186, w6187, w6188, w6189, w6190, w6191, w6192, w6193, w6194, w6195, w6196, w6197, w6198, w6199, w6200, w6201, w6202, w6203, w6204, w6205, w6206, w6207, w6208, w6209, w6210, w6211, w6212, w6213, w6214, w6215, w6216, w6217, w6218, w6219, w6220, w6221, w6222, w6223, w6224, w6225, w6226, w6227, w6228, w6229, w6230, w6231, w6232, w6233, w6234, w6235, w6236, w6237, w6238, w6239, w6240, w6241, w6242, w6243, w6244, w6245, w6246, w6247, w6248, w6249, w6250, w6251, w6252, w6253, w6254, w6255, w6256, w6257, w6258, w6259, w6260, w6261, w6262, w6263, w6264, w6265, w6266, w6267, w6268, w6269, w6270, w6271, w6272, w6273, w6274, w6275, w6276, w6277, w6278, w6279, w6280, w6281, w6282, w6283, w6284, w6285, w6286, w6287, w6288, w6289, w6290, w6291, w6292, w6293, w6294, w6295, w6296, w6297, w6298, w6299, w6300, w6301, w6302, w6303, w6304, w6305, w6306, w6307, w6308, w6309, w6310, w6311, w6312, w6313, w6314, w6315, w6316, w6317, w6318, w6319, w6320, w6321, w6322, w6323, w6324, w6325, w6326, w6327, w6328, w6329, w6330, w6331, w6332, w6333, w6334, w6335, w6336, w6337, w6338, w6339, w6340, w6341, w6342, w6343, w6344, w6345, w6346, w6347, w6348, w6349, w6350, w6351, w6352, w6353, w6354, w6355, w6356, w6357, w6358, w6359, w6360, w6361, w6362, w6363, w6364, w6365, w6366, w6367, w6368, w6369, w6370, w6371, w6372, w6373, w6374, w6375, w6376, w6377, w6378, w6379, w6380, w6381, w6382, w6383, w6384, w6385, w6386, w6387, w6388, w6389, w6390, w6391, w6392, w6393, w6394, w6395, w6396, w6397, w6398, w6399, w6400, w6401, w6402, w6403, w6404, w6405, w6406, w6407, w6408, w6409, w6410, w6411, w6412, w6413, w6414, w6415, w6416, w6417, w6418, w6419, w6420, w6421, w6422, w6423, w6424, w6425, w6426, w6427, w6428, w6429, w6430, w6431, w6432, w6433, w6434, w6435, w6436, w6437, w6438, w6439, w6440, w6441, w6442, w6443, w6444, w6445, w6446, w6447, w6448, w6449, w6450, w6451, w6452, w6453, w6454, w6455, w6456, w6457, w6458, w6459, w6460, w6461, w6462, w6463, w6464, w6465, w6466, w6467, w6468, w6469, w6470, w6471, w6472, w6473, w6474, w6475, w6476, w6477, w6478, w6479, w6480, w6481, w6482, w6483, w6484, w6485, w6486, w6487, w6488, w6489, w6490, w6491, w6492, w6493, w6494, w6495, w6496, w6497, w6498, w6499, w6500, w6501, w6502, w6503, w6504, w6505, w6506, w6507, w6508, w6509, w6510, w6511, w6512, w6513, w6514, w6515, w6516, w6517, w6518, w6519, w6520, w6521, w6522, w6523, w6524, w6525, w6526, w6527, w6528, w6529, w6530, w6531, w6532, w6533, w6534, w6535, w6536, w6537, w6538, w6539, w6540, w6541, w6542, w6543, w6544, w6545, w6546, w6547, w6548, w6549, w6550, w6551, w6552, w6553, w6554, w6555, w6556, w6557, w6558, w6559, w6560, w6561, w6562, w6563, w6564, w6565, w6566, w6567, w6568, w6569, w6570, w6571, w6572, w6573, w6574, w6575, w6576, w6577, w6578, w6579, w6580, w6581, w6582, w6583, w6584, w6585, w6586, w6587, w6588, w6589, w6590, w6591, w6592, w6593, w6594, w6595, w6596, w6597, w6598, w6599, w6600, w6601, w6602, w6603, w6604, w6605, w6606, w6607, w6608, w6609, w6610, w6611, w6612, w6613, w6614, w6615, w6616, w6617, w6618, w6619, w6620, w6621, w6622, w6623, w6624, w6625, w6626, w6627, w6628, w6629, w6630, w6631, w6632, w6633, w6634, w6635, w6636, w6637, w6638, w6639, w6640, w6641, w6642, w6643, w6644, w6645, w6646, w6647, w6648, w6649, w6650, w6651, w6652, w6653, w6654, w6655, w6656, w6657, w6658, w6659, w6660, w6661, w6662, w6663, w6664, w6665, w6666, w6667, w6668, w6669, w6670, w6671, w6672, w6673, w6674, w6675, w6676, w6677, w6678, w6679, w6680, w6681, w6682, w6683, w6684, w6685, w6686, w6687, w6688, w6689, w6690, w6691, w6692, w6693, w6694, w6695, w6696, w6697, w6698, w6699, w6700, w6701, w6702, w6703, w6704, w6705, w6706, w6707, w6708, w6709, w6710, w6711, w6712, w6713, w6714, w6715, w6716, w6717, w6718, w6719, w6720, w6721, w6722, w6723, w6724, w6725, w6726, w6727, w6728, w6729, w6730, w6731, w6732, w6733, w6734, w6735, w6736, w6737, w6738, w6739, w6740, w6741, w6742, w6743, w6744, w6745, w6746, w6747, w6748, w6749, w6750, w6751, w6752, w6753, w6754, w6755, w6756, w6757, w6758, w6759, w6760, w6761, w6762, w6763, w6764, w6765, w6766, w6767, w6768, w6769, w6770, w6771, w6772, w6773, w6774, w6775, w6776, w6777, w6778, w6779, w6780, w6781, w6782, w6783, w6784, w6785, w6786, w6787, w6788, w6789, w6790, w6791, w6792, w6793, w6794, w6795, w6796, w6797, w6798, w6799, w6800, w6801, w6802, w6803, w6804, w6805, w6806, w6807, w6808, w6809, w6810, w6811, w6812, w6813, w6814, w6815, w6816, w6817, w6818, w6819, w6820, w6821, w6822, w6823, w6824, w6825, w6826, w6827, w6828, w6829, w6830, w6831, w6832, w6833, w6834, w6835, w6836, w6837, w6838, w6839, w6840, w6841, w6842, w6843, w6844, w6845, w6846, w6847, w6848, w6849, w6850, w6851, w6852, w6853, w6854, w6855, w6856, w6857, w6858, w6859, w6860, w6861, w6862, w6863, w6864, w6865, w6866, w6867, w6868, w6869, w6870, w6871, w6872, w6873, w6874, w6875, w6876, w6877, w6878, w6879, w6880, w6881, w6882, w6883, w6884, w6885, w6886, w6887, w6888, w6889, w6890, w6891, w6892, w6893, w6894, w6895, w6896, w6897, w6898, w6899, w6900, w6901, w6902, w6903, w6904, w6905, w6906, w6907, w6908, w6909, w6910, w6911, w6912, w6913, w6914, w6915, w6916, w6917, w6918, w6919, w6920, w6921, w6922, w6923, w6924, w6925, w6926, w6927, w6928, w6929, w6930, w6931, w6932, w6933, w6934, w6935, w6936, w6937, w6938, w6939, w6940, w6941, w6942, w6943, w6944, w6945, w6946, w6947, w6948, w6949, w6950, w6951, w6952, w6953, w6954, w6955, w6956, w6957, w6958, w6959, w6960, w6961, w6962, w6963, w6964, w6965, w6966, w6967, w6968, w6969, w6970, w6971, w6972, w6973, w6974, w6975, w6976, w6977, w6978, w6979, w6980, w6981, w6982, w6983, w6984, w6985, w6986, w6987, w6988, w6989, w6990, w6991, w6992, w6993, w6994, w6995, w6996, w6997, w6998, w6999, w7000, w7001, w7002, w7003, w7004, w7005, w7006, w7007, w7008, w7009, w7010, w7011, w7012, w7013, w7014, w7015, w7016, w7017, w7018, w7019, w7020, w7021, w7022, w7023, w7024, w7025, w7026, w7027, w7028, w7029, w7030, w7031, w7032, w7033, w7034, w7035, w7036, w7037, w7038, w7039, w7040, w7041, w7042, w7043, w7044, w7045, w7046, w7047, w7048, w7049, w7050, w7051, w7052, w7053, w7054, w7055, w7056, w7057, w7058, w7059, w7060, w7061, w7062, w7063, w7064, w7065, w7066, w7067, w7068, w7069, w7070, w7071, w7072, w7073, w7074, w7075, w7076, w7077, w7078, w7079, w7080, w7081, w7082, w7083, w7084, w7085, w7086, w7087, w7088, w7089, w7090, w7091, w7092, w7093, w7094, w7095, w7096, w7097, w7098, w7099, w7100, w7101, w7102, w7103, w7104, w7105, w7106, w7107, w7108, w7109, w7110, w7111, w7112, w7113, w7114, w7115, w7116, w7117, w7118, w7119, w7120, w7121, w7122, w7123, w7124, w7125, w7126, w7127, w7128, w7129, w7130, w7131, w7132, w7133, w7134, w7135, w7136, w7137, w7138, w7139, w7140, w7141, w7142, w7143, w7144, w7145, w7146, w7147, w7148, w7149, w7150, w7151, w7152, w7153, w7154, w7155, w7156, w7157, w7158, w7159, w7160, w7161, w7162, w7163, w7164, w7165, w7166, w7167, w7168, w7169, w7170, w7171, w7172, w7173, w7174, w7175, w7176, w7177, w7178, w7179, w7180, w7181, w7182, w7183, w7184, w7185, w7186, w7187, w7188, w7189, w7190, w7191, w7192, w7193, w7194, w7195, w7196, w7197, w7198, w7199, w7200, w7201, w7202, w7203, w7204, w7205, w7206, w7207, w7208, w7209, w7210, w7211, w7212, w7213, w7214, w7215, w7216, w7217, w7218, w7219, w7220, w7221, w7222, w7223, w7224, w7225, w7226, w7227, w7228, w7229, w7230, w7231, w7232, w7233, w7234, w7235, w7236, w7237, w7238, w7239, w7240, w7241, w7242, w7243, w7244, w7245, w7246, w7247, w7248, w7249, w7250, w7251, w7252, w7253, w7254, w7255, w7256, w7257, w7258, w7259, w7260, w7261, w7262, w7263, w7264, w7265, w7266, w7267, w7268, w7269, w7270, w7271, w7272, w7273, w7274, w7275, w7276, w7277, w7278, w7279, w7280, w7281, w7282, w7283, w7284, w7285, w7286, w7287, w7288, w7289, w7290, w7291, w7292, w7293, w7294, w7295, w7296, w7297, w7298, w7299, w7300, w7301, w7302, w7303, w7304, w7305, w7306, w7307, w7308, w7309, w7310, w7311, w7312, w7313, w7314, w7315, w7316, w7317, w7318, w7319, w7320, w7321, w7322, w7323, w7324, w7325, w7326, w7327, w7328, w7329, w7330, w7331, w7332, w7333, w7334, w7335, w7336, w7337, w7338, w7339, w7340, w7341, w7342, w7343, w7344, w7345, w7346, w7347, w7348, w7349, w7350, w7351, w7352, w7353, w7354, w7355, w7356, w7357, w7358, w7359, w7360, w7361, w7362, w7363, w7364, w7365, w7366, w7367, w7368, w7369, w7370, w7371, w7372, w7373, w7374, w7375, w7376, w7377, w7378, w7379, w7380, w7381, w7382, w7383, w7384, w7385, w7386, w7387, w7388, w7389, w7390, w7391, w7392, w7393, w7394, w7395, w7396, w7397, w7398, w7399, w7400, w7401, w7402, w7403, w7404, w7405, w7406, w7407, w7408, w7409, w7410, w7411, w7412, w7413, w7414, w7415, w7416, w7417, w7418, w7419, w7420, w7421, w7422, w7423, w7424, w7425, w7426, w7427, w7428, w7429, w7430, w7431, w7432, w7433, w7434, w7435, w7436, w7437, w7438, w7439, w7440, w7441, w7442, w7443, w7444, w7445, w7446, w7447, w7448, w7449, w7450, w7451, w7452, w7453, w7454, w7455, w7456, w7457, w7458, w7459, w7460, w7461, w7462, w7463, w7464, w7465, w7466, w7467, w7468, w7469, w7470, w7471, w7472, w7473, w7474, w7475, w7476, w7477, w7478, w7479, w7480, w7481, w7482, w7483, w7484, w7485, w7486, w7487, w7488, w7489, w7490, w7491, w7492, w7493, w7494, w7495, w7496, w7497, w7498, w7499, w7500, w7501, w7502, w7503, w7504, w7505, w7506, w7507, w7508, w7509, w7510, w7511, w7512, w7513, w7514, w7515, w7516, w7517, w7518, w7519, w7520, w7521, w7522, w7523, w7524, w7525, w7526, w7527, w7528, w7529, w7530, w7531, w7532, w7533, w7534, w7535, w7536, w7537, w7538, w7539, w7540, w7541, w7542, w7543, w7544, w7545, w7546, w7547, w7548, w7549, w7550, w7551, w7552, w7553, w7554, w7555, w7556, w7557, w7558, w7559, w7560, w7561, w7562, w7563, w7564, w7565, w7566, w7567, w7568, w7569, w7570, w7571, w7572, w7573, w7574, w7575, w7576, w7577, w7578, w7579, w7580, w7581, w7582, w7583, w7584, w7585, w7586, w7587, w7588, w7589, w7590, w7591, w7592, w7593, w7594, w7595, w7596, w7597, w7598, w7599, w7600, w7601, w7602, w7603, w7604, w7605, w7606, w7607, w7608, w7609, w7610, w7611, w7612, w7613, w7614, w7615, w7616, w7617, w7618, w7619, w7620, w7621, w7622, w7623, w7624, w7625, w7626, w7627, w7628, w7629, w7630, w7631, w7632, w7633, w7634, w7635, w7636, w7637, w7638, w7639, w7640, w7641, w7642, w7643, w7644, w7645, w7646, w7647, w7648, w7649, w7650, w7651, w7652, w7653, w7654, w7655, w7656, w7657, w7658, w7659, w7660, w7661, w7662, w7663, w7664, w7665, w7666, w7667, w7668, w7669, w7670, w7671, w7672, w7673, w7674, w7675, w7676, w7677, w7678, w7679, w7680, w7681, w7682, w7683, w7684, w7685, w7686, w7687, w7688, w7689, w7690, w7691, w7692, w7693, w7694, w7695, w7696, w7697, w7698, w7699, w7700, w7701, w7702, w7703, w7704, w7705, w7706, w7707, w7708, w7709, w7710, w7711, w7712, w7713, w7714, w7715, w7716, w7717, w7718, w7719, w7720, w7721, w7722, w7723, w7724, w7725, w7726, w7727, w7728, w7729, w7730, w7731, w7732, w7733, w7734, w7735, w7736, w7737, w7738, w7739, w7740, w7741, w7742, w7743, w7744, w7745, w7746, w7747, w7748, w7749, w7750, w7751, w7752, w7753, w7754, w7755, w7756, w7757, w7758, w7759, w7760, w7761, w7762, w7763, w7764, w7765, w7766, w7767, w7768, w7769, w7770, w7771, w7772, w7773, w7774, w7775, w7776, w7777, w7778, w7779, w7780, w7781, w7782, w7783, w7784, w7785, w7786, w7787, w7788, w7789, w7790, w7791, w7792, w7793, w7794, w7795, w7796, w7797, w7798, w7799, w7800, w7801, w7802, w7803, w7804, w7805, w7806, w7807, w7808, w7809, w7810, w7811, w7812, w7813, w7814, w7815, w7816, w7817, w7818, w7819, w7820, w7821, w7822, w7823, w7824, w7825, w7826, w7827, w7828, w7829, w7830, w7831, w7832, w7833, w7834, w7835, w7836, w7837, w7838, w7839, w7840, w7841, w7842, w7843, w7844, w7845, w7846, w7847, w7848, w7849, w7850, w7851, w7852, w7853, w7854, w7855, w7856, w7857, w7858, w7859, w7860, w7861, w7862, w7863, w7864, w7865, w7866, w7867, w7868, w7869, w7870, w7871, w7872, w7873, w7874, w7875, w7876, w7877, w7878, w7879, w7880, w7881, w7882, w7883, w7884, w7885, w7886, w7887, w7888, w7889, w7890, w7891, w7892, w7893, w7894, w7895, w7896, w7897, w7898, w7899, w7900, w7901, w7902, w7903, w7904, w7905, w7906, w7907, w7908, w7909, w7910, w7911, w7912, w7913, w7914, w7915, w7916, w7917, w7918, w7919, w7920, w7921, w7922, w7923, w7924, w7925, w7926, w7927, w7928, w7929, w7930, w7931, w7932, w7933, w7934, w7935, w7936, w7937, w7938, w7939, w7940, w7941, w7942, w7943, w7944, w7945, w7946, w7947, w7948, w7949, w7950, w7951, w7952, w7953, w7954, w7955, w7956, w7957, w7958, w7959, w7960, w7961, w7962, w7963, w7964, w7965, w7966, w7967, w7968, w7969, w7970, w7971, w7972, w7973, w7974, w7975, w7976, w7977, w7978, w7979, w7980, w7981, w7982, w7983, w7984, w7985, w7986, w7987, w7988, w7989, w7990, w7991, w7992, w7993, w7994, w7995, w7996, w7997, w7998, w7999, w8000, w8001, w8002, w8003, w8004, w8005, w8006, w8007, w8008, w8009, w8010, w8011, w8012, w8013, w8014, w8015, w8016, w8017, w8018, w8019, w8020, w8021, w8022, w8023, w8024, w8025, w8026, w8027, w8028, w8029, w8030, w8031, w8032, w8033, w8034, w8035, w8036, w8037, w8038, w8039, w8040, w8041, w8042, w8043, w8044, w8045, w8046, w8047, w8048, w8049, w8050, w8051, w8052, w8053, w8054, w8055, w8056, w8057, w8058, w8059, w8060, w8061, w8062, w8063, w8064, w8065, w8066, w8067, w8068, w8069, w8070, w8071, w8072, w8073, w8074, w8075, w8076, w8077, w8078, w8079, w8080, w8081, w8082, w8083, w8084, w8085, w8086, w8087, w8088, w8089, w8090, w8091, w8092, w8093, w8094, w8095, w8096, w8097, w8098, w8099, w8100, w8101, w8102, w8103, w8104, w8105, w8106, w8107, w8108, w8109, w8110, w8111, w8112, w8113, w8114, w8115, w8116, w8117, w8118, w8119, w8120, w8121, w8122, w8123, w8124, w8125, w8126, w8127, w8128, w8129, w8130, w8131, w8132, w8133, w8134, w8135, w8136, w8137, w8138, w8139, w8140, w8141, w8142, w8143, w8144, w8145, w8146, w8147, w8148, w8149, w8150, w8151, w8152, w8153, w8154, w8155, w8156, w8157, w8158, w8159, w8160, w8161, w8162, w8163, w8164, w8165, w8166, w8167, w8168, w8169, w8170, w8171, w8172, w8173, w8174, w8175, w8176, w8177, w8178, w8179, w8180, w8181, w8182, w8183, w8184, w8185, w8186, w8187, w8188, w8189, w8190, w8191, w8192, w8193, w8194, w8195, w8196, w8197, w8198, w8199, w8200, w8201, w8202, w8203, w8204, w8205, w8206, w8207, w8208, w8209, w8210, w8211, w8212, w8213, w8214, w8215, w8216, w8217, w8218, w8219, w8220, w8221, w8222, w8223, w8224, w8225, w8226, w8227, w8228, w8229, w8230, w8231, w8232, w8233, w8234, w8235, w8236, w8237, w8238, w8239, w8240, w8241, w8242, w8243, w8244, w8245, w8246, w8247, w8248, w8249, w8250, w8251, w8252, w8253, w8254, w8255, w8256, w8257, w8258, w8259, w8260, w8261, w8262, w8263, w8264, w8265, w8266, w8267, w8268, w8269, w8270, w8271, w8272, w8273, w8274, w8275, w8276, w8277, w8278, w8279, w8280, w8281, w8282, w8283, w8284, w8285, w8286, w8287, w8288, w8289, w8290, w8291, w8292, w8293, w8294, w8295, w8296, w8297, w8298, w8299, w8300, w8301, w8302, w8303, w8304, w8305, w8306, w8307, w8308, w8309, w8310, w8311, w8312, w8313, w8314, w8315, w8316, w8317, w8318, w8319, w8320, w8321, w8322, w8323, w8324, w8325, w8326, w8327, w8328, w8329, w8330, w8331, w8332, w8333, w8334, w8335, w8336, w8337, w8338, w8339, w8340, w8341, w8342, w8343, w8344, w8345, w8346, w8347, w8348, w8349, w8350, w8351, w8352, w8353, w8354, w8355, w8356, w8357, w8358, w8359, w8360, w8361, w8362, w8363, w8364, w8365, w8366, w8367, w8368, w8369, w8370, w8371, w8372, w8373, w8374, w8375, w8376, w8377, w8378, w8379, w8380, w8381, w8382, w8383, w8384, w8385, w8386, w8387, w8388, w8389, w8390, w8391, w8392, w8393, w8394, w8395, w8396, w8397, w8398, w8399, w8400, w8401, w8402, w8403, w8404, w8405, w8406, w8407, w8408, w8409, w8410, w8411, w8412, w8413, w8414, w8415, w8416, w8417, w8418, w8419, w8420, w8421, w8422, w8423, w8424, w8425, w8426, w8427, w8428, w8429, w8430, w8431, w8432, w8433, w8434, w8435, w8436, w8437, w8438, w8439, w8440, w8441, w8442, w8443, w8444, w8445, w8446, w8447, w8448, w8449, w8450, w8451, w8452, w8453, w8454, w8455, w8456, w8457, w8458, w8459, w8460, w8461, w8462, w8463, w8464, w8465, w8466, w8467, w8468, w8469, w8470, w8471, w8472, w8473, w8474, w8475, w8476, w8477, w8478, w8479, w8480, w8481, w8482, w8483, w8484, w8485, w8486, w8487, w8488, w8489, w8490, w8491, w8492, w8493, w8494, w8495, w8496, w8497, w8498, w8499, w8500, w8501, w8502, w8503, w8504, w8505, w8506, w8507, w8508, w8509, w8510, w8511, w8512, w8513, w8514, w8515, w8516, w8517, w8518, w8519, w8520, w8521, w8522, w8523, w8524, w8525, w8526, w8527, w8528, w8529, w8530, w8531, w8532, w8533, w8534, w8535, w8536, w8537, w8538, w8539, w8540, w8541, w8542, w8543, w8544, w8545, w8546, w8547, w8548, w8549, w8550, w8551, w8552, w8553, w8554, w8555, w8556, w8557, w8558, w8559, w8560, w8561, w8562, w8563, w8564, w8565, w8566, w8567, w8568, w8569, w8570, w8571, w8572, w8573, w8574, w8575, w8576, w8577, w8578, w8579, w8580, w8581, w8582, w8583, w8584, w8585, w8586, w8587, w8588, w8589, w8590, w8591, w8592, w8593, w8594, w8595, w8596, w8597, w8598, w8599, w8600, w8601, w8602, w8603, w8604, w8605, w8606, w8607, w8608, w8609, w8610, w8611, w8612, w8613, w8614, w8615, w8616, w8617, w8618, w8619, w8620, w8621, w8622, w8623, w8624, w8625, w8626, w8627, w8628, w8629, w8630, w8631, w8632, w8633, w8634, w8635, w8636, w8637, w8638, w8639, w8640, w8641, w8642, w8643, w8644, w8645, w8646, w8647, w8648, w8649, w8650, w8651, w8652, w8653, w8654, w8655, w8656, w8657, w8658, w8659, w8660, w8661, w8662, w8663, w8664, w8665, w8666, w8667, w8668, w8669, w8670, w8671, w8672, w8673, w8674, w8675, w8676, w8677, w8678, w8679, w8680, w8681, w8682, w8683, w8684, w8685, w8686, w8687, w8688, w8689, w8690, w8691, w8692, w8693, w8694, w8695, w8696, w8697, w8698, w8699, w8700, w8701, w8702, w8703, w8704, w8705, w8706, w8707, w8708, w8709, w8710, w8711, w8712, w8713, w8714, w8715, w8716, w8717, w8718, w8719, w8720, w8721, w8722, w8723, w8724, w8725, w8726, w8727, w8728, w8729, w8730, w8731, w8732, w8733, w8734, w8735, w8736, w8737, w8738, w8739, w8740, w8741, w8742, w8743, w8744, w8745, w8746, w8747, w8748, w8749, w8750, w8751, w8752, w8753, w8754, w8755, w8756, w8757, w8758, w8759, w8760, w8761, w8762, w8763, w8764, w8765, w8766, w8767, w8768, w8769, w8770, w8771, w8772, w8773, w8774, w8775, w8776, w8777, w8778, w8779, w8780, w8781, w8782, w8783, w8784, w8785, w8786, w8787, w8788, w8789, w8790, w8791, w8792, w8793, w8794, w8795, w8796, w8797, w8798, w8799, w8800, w8801, w8802, w8803, w8804, w8805, w8806, w8807, w8808, w8809, w8810, w8811, w8812, w8813, w8814, w8815, w8816, w8817, w8818, w8819, w8820, w8821, w8822, w8823, w8824, w8825, w8826, w8827, w8828, w8829, w8830, w8831, w8832, w8833, w8834, w8835, w8836, w8837, w8838, w8839, w8840, w8841, w8842, w8843, w8844, w8845, w8846, w8847, w8848, w8849, w8850, w8851, w8852, w8853, w8854, w8855, w8856, w8857, w8858, w8859, w8860, w8861, w8862, w8863, w8864, w8865, w8866, w8867, w8868, w8869, w8870, w8871, w8872, w8873, w8874, w8875, w8876, w8877, w8878, w8879, w8880, w8881, w8882, w8883, w8884, w8885, w8886, w8887, w8888, w8889, w8890, w8891, w8892, w8893, w8894, w8895, w8896, w8897, w8898, w8899, w8900, w8901, w8902, w8903, w8904, w8905, w8906, w8907, w8908, w8909, w8910, w8911, w8912, w8913, w8914, w8915, w8916, w8917, w8918, w8919, w8920, w8921, w8922, w8923, w8924, w8925, w8926, w8927, w8928, w8929, w8930, w8931, w8932, w8933, w8934, w8935, w8936, w8937, w8938, w8939, w8940, w8941, w8942, w8943, w8944, w8945, w8946, w8947, w8948, w8949, w8950, w8951, w8952, w8953, w8954, w8955, w8956, w8957, w8958, w8959, w8960, w8961, w8962, w8963, w8964, w8965, w8966, w8967, w8968, w8969, w8970, w8971, w8972, w8973, w8974, w8975, w8976, w8977, w8978, w8979, w8980, w8981, w8982, w8983, w8984, w8985, w8986, w8987, w8988, w8989, w8990, w8991, w8992, w8993, w8994, w8995, w8996, w8997, w8998, w8999, w9000, w9001, w9002, w9003, w9004, w9005, w9006, w9007, w9008, w9009, w9010, w9011, w9012, w9013, w9014, w9015, w9016, w9017, w9018, w9019, w9020, w9021, w9022, w9023, w9024, w9025, w9026, w9027, w9028, w9029, w9030, w9031, w9032, w9033, w9034, w9035, w9036, w9037, w9038, w9039, w9040, w9041, w9042, w9043, w9044, w9045, w9046, w9047, w9048, w9049, w9050, w9051, w9052, w9053, w9054, w9055, w9056, w9057, w9058, w9059, w9060, w9061, w9062, w9063, w9064, w9065, w9066, w9067, w9068, w9069, w9070, w9071, w9072, w9073, w9074, w9075, w9076, w9077, w9078, w9079, w9080, w9081, w9082, w9083, w9084, w9085, w9086, w9087, w9088, w9089, w9090, w9091, w9092, w9093, w9094, w9095, w9096, w9097, w9098, w9099, w9100, w9101, w9102, w9103, w9104, w9105, w9106, w9107, w9108, w9109, w9110, w9111, w9112, w9113, w9114, w9115, w9116, w9117, w9118, w9119, w9120, w9121, w9122, w9123, w9124, w9125, w9126, w9127, w9128, w9129, w9130, w9131, w9132, w9133, w9134, w9135, w9136, w9137, w9138, w9139, w9140, w9141, w9142, w9143, w9144, w9145, w9146, w9147, w9148, w9149, w9150, w9151, w9152, w9153, w9154, w9155, w9156, w9157, w9158, w9159, w9160, w9161, w9162, w9163, w9164, w9165, w9166, w9167, w9168, w9169, w9170, w9171, w9172, w9173, w9174, w9175, w9176, w9177, w9178, w9179, w9180, w9181, w9182, w9183, w9184, w9185, w9186, w9187, w9188, w9189, w9190, w9191, w9192, w9193, w9194, w9195, w9196, w9197, w9198, w9199, w9200, w9201, w9202, w9203, w9204, w9205, w9206, w9207, w9208, w9209, w9210, w9211, w9212, w9213, w9214, w9215, w9216, w9217, w9218, w9219, w9220, w9221, w9222, w9223, w9224, w9225, w9226, w9227, w9228, w9229, w9230, w9231, w9232, w9233, w9234, w9235, w9236, w9237, w9238, w9239, w9240, w9241, w9242, w9243, w9244, w9245, w9246, w9247, w9248, w9249, w9250, w9251, w9252, w9253, w9254, w9255, w9256, w9257, w9258, w9259, w9260, w9261, w9262, w9263, w9264, w9265, w9266, w9267, w9268, w9269, w9270, w9271, w9272, w9273, w9274, w9275, w9276, w9277, w9278, w9279, w9280, w9281, w9282, w9283, w9284, w9285, w9286, w9287, w9288, w9289, w9290, w9291, w9292, w9293, w9294, w9295, w9296, w9297, w9298, w9299, w9300, w9301, w9302, w9303, w9304, w9305, w9306, w9307, w9308, w9309, w9310, w9311, w9312, w9313, w9314, w9315, w9316, w9317, w9318, w9319, w9320, w9321, w9322, w9323, w9324, w9325, w9326, w9327, w9328, w9329, w9330, w9331, w9332, w9333, w9334, w9335, w9336, w9337, w9338, w9339, w9340, w9341, w9342, w9343, w9344, w9345, w9346, w9347, w9348, w9349, w9350, w9351, w9352, w9353, w9354, w9355, w9356, w9357, w9358, w9359, w9360, w9361, w9362, w9363, w9364, w9365, w9366, w9367, w9368, w9369, w9370, w9371, w9372, w9373, w9374, w9375, w9376, w9377, w9378, w9379, w9380, w9381, w9382, w9383, w9384, w9385, w9386, w9387, w9388, w9389, w9390, w9391, w9392, w9393, w9394, w9395, w9396, w9397, w9398, w9399, w9400, w9401, w9402, w9403, w9404, w9405, w9406, w9407, w9408, w9409, w9410, w9411, w9412, w9413, w9414, w9415, w9416, w9417, w9418, w9419, w9420, w9421, w9422, w9423, w9424, w9425, w9426, w9427, w9428, w9429, w9430, w9431, w9432, w9433, w9434, w9435, w9436, w9437, w9438, w9439, w9440, w9441, w9442, w9443, w9444, w9445, w9446, w9447, w9448, w9449, w9450, w9451, w9452, w9453, w9454, w9455, w9456, w9457, w9458, w9459, w9460, w9461, w9462, w9463, w9464, w9465, w9466, w9467, w9468, w9469, w9470, w9471, w9472, w9473, w9474, w9475, w9476, w9477, w9478, w9479, w9480, w9481, w9482, w9483, w9484, w9485, w9486, w9487, w9488, w9489, w9490, w9491, w9492, w9493, w9494, w9495, w9496, w9497, w9498, w9499, w9500, w9501, w9502, w9503, w9504, w9505, w9506, w9507, w9508, w9509, w9510, w9511, w9512, w9513, w9514, w9515, w9516, w9517, w9518, w9519, w9520, w9521, w9522, w9523, w9524, w9525, w9526, w9527, w9528, w9529, w9530, w9531, w9532, w9533, w9534, w9535, w9536, w9537, w9538, w9539, w9540, w9541, w9542, w9543, w9544, w9545, w9546, w9547, w9548, w9549, w9550, w9551, w9552, w9553, w9554, w9555, w9556, w9557, w9558, w9559, w9560, w9561, w9562, w9563, w9564, w9565, w9566, w9567, w9568, w9569, w9570, w9571, w9572, w9573, w9574, w9575, w9576, w9577, w9578, w9579, w9580, w9581, w9582, w9583, w9584, w9585, w9586, w9587, w9588, w9589, w9590, w9591, w9592, w9593, w9594, w9595, w9596, w9597, w9598, w9599, w9600, w9601, w9602, w9603, w9604, w9605, w9606, w9607, w9608, w9609, w9610, w9611, w9612, w9613, w9614, w9615, w9616, w9617, w9618, w9619, w9620, w9621, w9622, w9623, w9624, w9625, w9626, w9627, w9628, w9629, w9630, w9631, w9632, w9633, w9634, w9635, w9636, w9637, w9638, w9639, w9640, w9641, w9642, w9643, w9644, w9645, w9646, w9647, w9648, w9649, w9650, w9651, w9652, w9653, w9654, w9655, w9656, w9657, w9658, w9659, w9660, w9661, w9662, w9663, w9664, w9665, w9666, w9667, w9668, w9669, w9670, w9671, w9672, w9673, w9674, w9675, w9676, w9677, w9678, w9679, w9680, w9681, w9682, w9683, w9684, w9685, w9686, w9687, w9688, w9689, w9690, w9691, w9692, w9693, w9694, w9695, w9696, w9697, w9698, w9699, w9700, w9701, w9702, w9703, w9704, w9705, w9706, w9707, w9708, w9709, w9710, w9711, w9712, w9713, w9714, w9715, w9716, w9717, w9718, w9719, w9720, w9721, w9722, w9723, w9724, w9725, w9726, w9727, w9728, w9729, w9730, w9731, w9732, w9733, w9734, w9735, w9736, w9737, w9738, w9739, w9740, w9741, w9742, w9743, w9744, w9745, w9746, w9747, w9748, w9749, w9750, w9751, w9752, w9753, w9754, w9755, w9756, w9757, w9758, w9759, w9760, w9761, w9762, w9763, w9764, w9765, w9766, w9767, w9768, w9769, w9770, w9771, w9772, w9773, w9774, w9775, w9776, w9777, w9778, w9779, w9780, w9781, w9782, w9783, w9784, w9785, w9786, w9787, w9788, w9789, w9790, w9791, w9792, w9793, w9794, w9795, w9796, w9797, w9798, w9799, w9800, w9801, w9802, w9803, w9804, w9805, w9806, w9807, w9808, w9809, w9810, w9811, w9812, w9813, w9814, w9815, w9816, w9817, w9818, w9819, w9820, w9821, w9822, w9823, w9824, w9825, w9826, w9827, w9828, w9829, w9830, w9831, w9832, w9833, w9834, w9835, w9836, w9837, w9838, w9839, w9840, w9841, w9842, w9843, w9844, w9845, w9846, w9847, w9848, w9849, w9850, w9851, w9852, w9853, w9854, w9855, w9856, w9857, w9858, w9859, w9860, w9861, w9862, w9863, w9864, w9865, w9866, w9867, w9868, w9869, w9870, w9871, w9872, w9873, w9874, w9875, w9876, w9877, w9878, w9879, w9880, w9881, w9882, w9883, w9884, w9885, w9886, w9887, w9888, w9889, w9890, w9891, w9892, w9893, w9894, w9895, w9896, w9897, w9898, w9899, w9900, w9901, w9902, w9903, w9904, w9905, w9906, w9907, w9908, w9909, w9910, w9911, w9912, w9913, w9914, w9915, w9916, w9917, w9918, w9919, w9920, w9921, w9922, w9923, w9924, w9925, w9926, w9927, w9928, w9929, w9930, w9931, w9932, w9933, w9934, w9935, w9936, w9937, w9938, w9939, w9940, w9941, w9942, w9943, w9944, w9945, w9946, w9947, w9948, w9949, w9950, w9951, w9952, w9953, w9954, w9955, w9956, w9957, w9958, w9959, w9960, w9961, w9962, w9963, w9964, w9965, w9966, w9967, w9968, w9969, w9970, w9971, w9972, w9973, w9974, w9975, w9976, w9977, w9978, w9979, w9980, w9981, w9982, w9983, w9984, w9985, w9986, w9987, w9988, w9989, w9990, w9991, w9992, w9993, w9994, w9995, w9996, w9997, w9998, w9999, w10000, w10001, w10002, w10003, w10004, w10005, w10006, w10007, w10008, w10009, w10010, w10011, w10012, w10013, w10014, w10015, w10016, w10017, w10018, w10019, w10020, w10021, w10022, w10023, w10024, w10025, w10026, w10027, w10028, w10029, w10030, w10031, w10032, w10033, w10034, w10035, w10036, w10037, w10038, w10039, w10040, w10041, w10042, w10043, w10044, w10045, w10046, w10047, w10048, w10049, w10050, w10051, w10052, w10053, w10054, w10055, w10056, w10057, w10058, w10059, w10060, w10061, w10062, w10063, w10064, w10065, w10066, w10067, w10068, w10069, w10070, w10071, w10072, w10073, w10074, w10075, w10076, w10077, w10078, w10079, w10080, w10081, w10082, w10083, w10084, w10085, w10086, w10087, w10088, w10089, w10090, w10091, w10092, w10093, w10094, w10095, w10096, w10097, w10098, w10099, w10100, w10101, w10102, w10103, w10104, w10105, w10106, w10107, w10108, w10109, w10110, w10111, w10112, w10113, w10114, w10115, w10116, w10117, w10118, w10119, w10120, w10121, w10122, w10123, w10124, w10125, w10126, w10127, w10128, w10129, w10130, w10131, w10132, w10133, w10134, w10135, w10136, w10137, w10138, w10139, w10140, w10141, w10142, w10143, w10144, w10145, w10146, w10147, w10148, w10149, w10150, w10151, w10152, w10153, w10154, w10155, w10156, w10157, w10158, w10159, w10160, w10161, w10162, w10163, w10164, w10165, w10166, w10167, w10168, w10169, w10170, w10171, w10172, w10173, w10174, w10175, w10176, w10177, w10178, w10179, w10180, w10181, w10182, w10183, w10184, w10185, w10186, w10187, w10188, w10189, w10190, w10191, w10192, w10193, w10194, w10195, w10196, w10197, w10198, w10199, w10200, w10201, w10202, w10203, w10204, w10205, w10206, w10207, w10208, w10209, w10210, w10211, w10212, w10213, w10214, w10215, w10216, w10217, w10218, w10219, w10220, w10221, w10222, w10223, w10224, w10225, w10226, w10227, w10228, w10229, w10230, w10231, w10232, w10233, w10234, w10235, w10236, w10237, w10238, w10239, w10240, w10241, w10242, w10243, w10244, w10245, w10246, w10247, w10248, w10249, w10250, w10251, w10252, w10253, w10254, w10255, w10256, w10257, w10258, w10259, w10260, w10261, w10262, w10263, w10264, w10265, w10266, w10267, w10268, w10269, w10270, w10271, w10272, w10273, w10274, w10275, w10276, w10277, w10278, w10279, w10280, w10281, w10282, w10283, w10284, w10285, w10286, w10287, w10288, w10289, w10290, w10291, w10292, w10293, w10294, w10295, w10296, w10297, w10298, w10299, w10300, w10301, w10302, w10303, w10304, w10305, w10306, w10307, w10308, w10309, w10310, w10311, w10312, w10313, w10314, w10315, w10316, w10317, w10318, w10319, w10320, w10321, w10322, w10323, w10324, w10325, w10326, w10327, w10328, w10329, w10330, w10331, w10332, w10333, w10334, w10335, w10336, w10337, w10338, w10339, w10340, w10341, w10342, w10343, w10344, w10345, w10346, w10347, w10348, w10349, w10350, w10351, w10352, w10353, w10354, w10355, w10356, w10357, w10358, w10359, w10360, w10361, w10362, w10363, w10364, w10365, w10366, w10367, w10368, w10369, w10370, w10371, w10372, w10373, w10374, w10375, w10376, w10377, w10378, w10379, w10380, w10381, w10382, w10383, w10384, w10385, w10386, w10387, w10388, w10389, w10390, w10391, w10392, w10393, w10394, w10395, w10396, w10397, w10398, w10399, w10400, w10401, w10402, w10403, w10404, w10405, w10406, w10407, w10408, w10409, w10410, w10411, w10412, w10413, w10414, w10415, w10416, w10417, w10418, w10419, w10420, w10421, w10422, w10423, w10424, w10425, w10426, w10427, w10428, w10429, w10430, w10431, w10432, w10433, w10434, w10435, w10436, w10437, w10438, w10439, w10440, w10441, w10442, w10443, w10444, w10445, w10446, w10447, w10448, w10449, w10450, w10451, w10452, w10453, w10454, w10455, w10456, w10457, w10458, w10459, w10460, w10461, w10462, w10463, w10464, w10465, w10466, w10467, w10468, w10469, w10470, w10471, w10472, w10473, w10474, w10475, w10476, w10477, w10478, w10479, w10480, w10481, w10482, w10483, w10484, w10485, w10486, w10487, w10488, w10489, w10490, w10491, w10492, w10493, w10494, w10495, w10496, w10497, w10498, w10499, w10500, w10501, w10502, w10503, w10504, w10505, w10506, w10507, w10508, w10509, w10510, w10511, w10512, w10513, w10514, w10515, w10516, w10517, w10518, w10519, w10520, w10521, w10522, w10523, w10524, w10525, w10526, w10527, w10528, w10529, w10530, w10531, w10532, w10533, w10534, w10535, w10536, w10537, w10538, w10539, w10540, w10541, w10542, w10543, w10544, w10545, w10546, w10547, w10548, w10549, w10550, w10551, w10552, w10553, w10554, w10555, w10556, w10557, w10558, w10559, w10560, w10561, w10562, w10563, w10564, w10565, w10566, w10567, w10568, w10569, w10570, w10571, w10572, w10573, w10574, w10575, w10576, w10577, w10578, w10579, w10580, w10581, w10582, w10583, w10584, w10585, w10586, w10587, w10588, w10589, w10590, w10591, w10592, w10593, w10594, w10595, w10596, w10597, w10598, w10599, w10600, w10601, w10602, w10603, w10604, w10605, w10606, w10607, w10608, w10609, w10610, w10611, w10612, w10613, w10614, w10615, w10616, w10617, w10618, w10619, w10620, w10621, w10622, w10623, w10624, w10625, w10626, w10627, w10628, w10629, w10630, w10631, w10632, w10633, w10634, w10635, w10636, w10637, w10638, w10639, w10640, w10641, w10642, w10643, w10644, w10645, w10646, w10647, w10648, w10649, w10650, w10651, w10652, w10653, w10654, w10655, w10656, w10657, w10658, w10659, w10660, w10661, w10662, w10663, w10664, w10665, w10666, w10667, w10668, w10669, w10670, w10671, w10672, w10673, w10674, w10675, w10676, w10677, w10678, w10679, w10680, w10681, w10682, w10683, w10684, w10685, w10686, w10687, w10688, w10689, w10690, w10691, w10692, w10693, w10694, w10695, w10696, w10697, w10698, w10699, w10700, w10701, w10702, w10703, w10704, w10705, w10706, w10707, w10708, w10709, w10710, w10711, w10712, w10713, w10714, w10715, w10716, w10717, w10718, w10719, w10720, w10721, w10722, w10723, w10724, w10725, w10726, w10727, w10728, w10729, w10730, w10731, w10732, w10733, w10734, w10735, w10736, w10737, w10738, w10739, w10740, w10741, w10742, w10743, w10744, w10745, w10746, w10747, w10748, w10749, w10750, w10751, w10752, w10753, w10754, w10755, w10756, w10757, w10758, w10759, w10760, w10761, w10762, w10763, w10764, w10765, w10766, w10767, w10768, w10769, w10770, w10771, w10772, w10773, w10774, w10775, w10776, w10777, w10778, w10779, w10780, w10781, w10782, w10783, w10784, w10785, w10786, w10787, w10788, w10789, w10790, w10791, w10792, w10793, w10794, w10795, w10796, w10797, w10798, w10799, w10800, w10801, w10802, w10803, w10804, w10805, w10806, w10807, w10808, w10809, w10810, w10811, w10812, w10813, w10814, w10815, w10816, w10817, w10818, w10819, w10820, w10821, w10822, w10823, w10824, w10825, w10826, w10827, w10828, w10829, w10830, w10831, w10832, w10833, w10834, w10835, w10836, w10837, w10838, w10839, w10840, w10841, w10842, w10843, w10844, w10845, w10846, w10847, w10848, w10849, w10850, w10851, w10852, w10853, w10854, w10855, w10856, w10857, w10858, w10859, w10860, w10861, w10862, w10863, w10864, w10865, w10866, w10867, w10868, w10869, w10870, w10871, w10872, w10873, w10874, w10875, w10876, w10877, w10878, w10879, w10880, w10881, w10882, w10883, w10884, w10885, w10886, w10887, w10888, w10889, w10890, w10891, w10892, w10893, w10894, w10895, w10896, w10897, w10898, w10899, w10900, w10901, w10902, w10903, w10904, w10905, w10906, w10907, w10908, w10909, w10910, w10911, w10912, w10913, w10914, w10915, w10916, w10917, w10918, w10919, w10920, w10921, w10922, w10923, w10924, w10925, w10926, w10927, w10928, w10929, w10930, w10931, w10932, w10933, w10934, w10935, w10936, w10937, w10938, w10939, w10940, w10941, w10942, w10943, w10944, w10945, w10946, w10947, w10948, w10949, w10950, w10951, w10952, w10953, w10954, w10955, w10956, w10957, w10958, w10959, w10960, w10961, w10962, w10963, w10964, w10965, w10966, w10967, w10968, w10969, w10970, w10971, w10972, w10973, w10974, w10975, w10976, w10977, w10978, w10979, w10980, w10981, w10982, w10983, w10984, w10985, w10986, w10987, w10988, w10989, w10990, w10991, w10992, w10993, w10994, w10995, w10996, w10997, w10998, w10999, w11000, w11001, w11002, w11003, w11004, w11005, w11006, w11007, w11008, w11009, w11010, w11011, w11012, w11013, w11014, w11015, w11016, w11017, w11018, w11019, w11020, w11021, w11022, w11023, w11024, w11025, w11026, w11027, w11028, w11029, w11030, w11031, w11032, w11033, w11034, w11035, w11036, w11037, w11038, w11039, w11040, w11041, w11042, w11043, w11044, w11045, w11046, w11047, w11048, w11049, w11050, w11051, w11052, w11053, w11054, w11055, w11056, w11057, w11058, w11059, w11060, w11061, w11062, w11063, w11064, w11065, w11066, w11067, w11068, w11069, w11070, w11071, w11072, w11073, w11074, w11075, w11076, w11077, w11078, w11079, w11080, w11081, w11082, w11083, w11084, w11085, w11086, w11087, w11088, w11089, w11090, w11091, w11092, w11093, w11094, w11095, w11096, w11097, w11098, w11099, w11100, w11101, w11102, w11103, w11104, w11105, w11106, w11107, w11108, w11109, w11110, w11111, w11112, w11113, w11114, w11115, w11116, w11117, w11118, w11119, w11120, w11121, w11122, w11123, w11124, w11125, w11126, w11127, w11128, w11129, w11130, w11131, w11132, w11133, w11134, w11135, w11136, w11137, w11138, w11139, w11140, w11141, w11142, w11143, w11144, w11145, w11146, w11147, w11148, w11149, w11150, w11151, w11152, w11153, w11154, w11155, w11156, w11157, w11158, w11159, w11160, w11161, w11162, w11163, w11164, w11165, w11166, w11167, w11168, w11169, w11170, w11171, w11172, w11173, w11174, w11175, w11176, w11177, w11178, w11179, w11180, w11181, w11182, w11183, w11184, w11185, w11186, w11187, w11188, w11189, w11190, w11191, w11192, w11193, w11194, w11195, w11196, w11197, w11198, w11199, w11200, w11201, w11202, w11203, w11204, w11205, w11206, w11207, w11208, w11209, w11210, w11211, w11212, w11213, w11214, w11215, w11216, w11217, w11218, w11219, w11220, w11221, w11222, w11223, w11224, w11225, w11226, w11227, w11228, w11229, w11230, w11231, w11232, w11233, w11234, w11235, w11236, w11237, w11238, w11239, w11240, w11241, w11242, w11243, w11244, w11245, w11246, w11247, w11248, w11249, w11250, w11251, w11252, w11253, w11254, w11255, w11256, w11257, w11258, w11259, w11260, w11261, w11262, w11263, w11264, w11265, w11266, w11267, w11268, w11269, w11270, w11271, w11272, w11273, w11274, w11275, w11276, w11277, w11278, w11279, w11280, w11281, w11282, w11283, w11284, w11285, w11286, w11287, w11288, w11289, w11290, w11291, w11292, w11293, w11294, w11295, w11296, w11297, w11298, w11299, w11300, w11301, w11302, w11303, w11304, w11305, w11306, w11307, w11308, w11309, w11310, w11311, w11312, w11313, w11314, w11315, w11316, w11317, w11318, w11319, w11320, w11321, w11322, w11323, w11324, w11325, w11326, w11327, w11328, w11329, w11330, w11331, w11332, w11333, w11334, w11335, w11336, w11337, w11338, w11339, w11340, w11341, w11342, w11343, w11344, w11345, w11346, w11347, w11348, w11349, w11350, w11351, w11352, w11353, w11354, w11355, w11356, w11357, w11358, w11359, w11360, w11361, w11362, w11363, w11364, w11365, w11366, w11367, w11368, w11369, w11370, w11371, w11372, w11373, w11374, w11375, w11376, w11377, w11378, w11379, w11380, w11381, w11382, w11383, w11384, w11385, w11386, w11387, w11388, w11389, w11390, w11391, w11392, w11393, w11394, w11395, w11396, w11397, w11398, w11399, w11400, w11401, w11402, w11403, w11404, w11405, w11406, w11407, w11408, w11409, w11410, w11411, w11412, w11413, w11414, w11415, w11416, w11417, w11418, w11419, w11420, w11421, w11422, w11423, w11424, w11425, w11426, w11427, w11428, w11429, w11430, w11431, w11432, w11433, w11434, w11435, w11436, w11437, w11438, w11439, w11440, w11441, w11442, w11443, w11444, w11445, w11446, w11447, w11448, w11449, w11450, w11451, w11452, w11453, w11454, w11455, w11456, w11457, w11458, w11459, w11460, w11461, w11462, w11463, w11464, w11465, w11466, w11467, w11468, w11469, w11470, w11471, w11472, w11473, w11474, w11475, w11476, w11477, w11478, w11479, w11480, w11481, w11482, w11483, w11484, w11485, w11486, w11487, w11488, w11489, w11490, w11491, w11492, w11493, w11494, w11495, w11496, w11497, w11498, w11499, w11500, w11501, w11502, w11503, w11504, w11505, w11506, w11507, w11508, w11509, w11510, w11511, w11512, w11513, w11514, w11515, w11516, w11517, w11518, w11519, w11520, w11521, w11522, w11523, w11524, w11525, w11526, w11527, w11528, w11529, w11530, w11531, w11532, w11533, w11534, w11535, w11536, w11537, w11538, w11539, w11540, w11541, w11542, w11543, w11544, w11545, w11546, w11547, w11548, w11549, w11550, w11551, w11552, w11553, w11554, w11555, w11556, w11557, w11558, w11559, w11560, w11561, w11562, w11563, w11564, w11565, w11566, w11567, w11568, w11569, w11570, w11571, w11572, w11573, w11574, w11575, w11576, w11577, w11578, w11579, w11580, w11581, w11582, w11583, w11584, w11585, w11586, w11587, w11588, w11589, w11590, w11591, w11592, w11593, w11594, w11595, w11596, w11597, w11598, w11599, w11600, w11601, w11602, w11603, w11604, w11605, w11606, w11607, w11608, w11609, w11610, w11611, w11612, w11613, w11614, w11615, w11616, w11617, w11618, w11619, w11620, w11621, w11622, w11623, w11624, w11625, w11626, w11627, w11628, w11629, w11630, w11631, w11632, w11633, w11634, w11635, w11636, w11637, w11638, w11639, w11640, w11641, w11642, w11643, w11644, w11645, w11646, w11647, w11648, w11649, w11650, w11651, w11652, w11653, w11654, w11655, w11656, w11657, w11658, w11659, w11660, w11661, w11662, w11663, w11664, w11665, w11666, w11667, w11668, w11669, w11670, w11671, w11672, w11673, w11674, w11675, w11676, w11677, w11678, w11679, w11680, w11681, w11682, w11683, w11684, w11685, w11686, w11687, w11688, w11689, w11690, w11691, w11692, w11693, w11694, w11695, w11696, w11697, w11698, w11699, w11700, w11701, w11702, w11703, w11704, w11705, w11706, w11707, w11708, w11709, w11710, w11711, w11712, w11713, w11714, w11715, w11716, w11717, w11718, w11719, w11720, w11721, w11722, w11723, w11724, w11725, w11726, w11727, w11728, w11729, w11730, w11731, w11732, w11733, w11734, w11735, w11736, w11737, w11738, w11739, w11740, w11741, w11742, w11743, w11744, w11745, w11746, w11747, w11748, w11749, w11750, w11751, w11752, w11753, w11754, w11755, w11756, w11757, w11758, w11759, w11760, w11761, w11762, w11763, w11764, w11765, w11766, w11767, w11768, w11769, w11770, w11771, w11772, w11773, w11774, w11775, w11776, w11777, w11778, w11779, w11780, w11781, w11782, w11783, w11784, w11785, w11786, w11787, w11788, w11789, w11790, w11791, w11792, w11793, w11794, w11795, w11796, w11797, w11798, w11799, w11800, w11801, w11802, w11803, w11804, w11805, w11806, w11807, w11808, w11809, w11810, w11811, w11812, w11813, w11814, w11815, w11816, w11817, w11818, w11819, w11820, w11821, w11822, w11823, w11824, w11825, w11826, w11827, w11828, w11829, w11830, w11831, w11832, w11833, w11834, w11835, w11836, w11837, w11838, w11839, w11840, w11841, w11842, w11843, w11844, w11845, w11846, w11847, w11848, w11849, w11850, w11851, w11852, w11853, w11854, w11855, w11856, w11857, w11858, w11859, w11860, w11861, w11862, w11863, w11864, w11865, w11866, w11867, w11868, w11869, w11870, w11871, w11872, w11873, w11874, w11875, w11876, w11877, w11878, w11879, w11880, w11881, w11882, w11883, w11884, w11885, w11886, w11887, w11888, w11889, w11890, w11891, w11892, w11893, w11894, w11895, w11896, w11897, w11898, w11899, w11900, w11901, w11902, w11903, w11904, w11905, w11906, w11907, w11908, w11909, w11910, w11911, w11912, w11913, w11914, w11915, w11916, w11917, w11918, w11919, w11920, w11921, w11922, w11923, w11924, w11925, w11926, w11927, w11928, w11929, w11930, w11931, w11932, w11933, w11934, w11935, w11936, w11937, w11938, w11939, w11940, w11941, w11942, w11943, w11944, w11945, w11946, w11947, w11948, w11949, w11950, w11951, w11952, w11953, w11954, w11955, w11956, w11957, w11958, w11959, w11960, w11961, w11962, w11963, w11964, w11965, w11966, w11967, w11968, w11969, w11970, w11971, w11972, w11973, w11974, w11975, w11976, w11977, w11978, w11979, w11980, w11981, w11982, w11983, w11984, w11985, w11986, w11987, w11988, w11989, w11990, w11991, w11992, w11993, w11994, w11995, w11996, w11997, w11998, w11999, w12000, w12001, w12002, w12003, w12004, w12005, w12006, w12007, w12008, w12009, w12010, w12011, w12012, w12013, w12014, w12015, w12016, w12017, w12018, w12019, w12020, w12021, w12022, w12023, w12024, w12025, w12026, w12027, w12028, w12029, w12030, w12031, w12032, w12033, w12034, w12035, w12036, w12037, w12038, w12039, w12040, w12041, w12042, w12043, w12044, w12045, w12046, w12047, w12048, w12049, w12050, w12051, w12052, w12053, w12054, w12055, w12056, w12057, w12058, w12059, w12060, w12061, w12062, w12063, w12064, w12065, w12066, w12067, w12068, w12069, w12070, w12071, w12072, w12073, w12074, w12075, w12076, w12077, w12078, w12079, w12080, w12081, w12082, w12083, w12084, w12085, w12086, w12087, w12088, w12089, w12090, w12091, w12092, w12093, w12094, w12095, w12096, w12097, w12098, w12099, w12100, w12101, w12102, w12103, w12104, w12105, w12106, w12107, w12108, w12109, w12110, w12111, w12112, w12113, w12114, w12115, w12116, w12117, w12118, w12119, w12120, w12121, w12122, w12123, w12124, w12125, w12126, w12127, w12128, w12129, w12130, w12131, w12132, w12133, w12134, w12135, w12136, w12137, w12138, w12139, w12140, w12141, w12142, w12143, w12144, w12145, w12146, w12147, w12148, w12149, w12150, w12151, w12152, w12153, w12154, w12155, w12156, w12157, w12158, w12159, w12160, w12161, w12162, w12163, w12164, w12165, w12166, w12167, w12168, w12169, w12170, w12171, w12172, w12173, w12174, w12175, w12176, w12177, w12178, w12179, w12180, w12181, w12182, w12183, w12184, w12185, w12186, w12187, w12188, w12189, w12190, w12191, w12192, w12193, w12194, w12195, w12196, w12197, w12198, w12199, w12200, w12201, w12202, w12203, w12204, w12205, w12206, w12207, w12208, w12209, w12210, w12211, w12212, w12213, w12214, w12215, w12216, w12217, w12218, w12219, w12220, w12221, w12222, w12223, w12224, w12225, w12226, w12227, w12228, w12229, w12230, w12231, w12232, w12233, w12234, w12235, w12236, w12237, w12238, w12239, w12240, w12241, w12242, w12243, w12244, w12245, w12246, w12247, w12248, w12249, w12250, w12251, w12252, w12253, w12254, w12255, w12256, w12257, w12258, w12259, w12260, w12261, w12262, w12263, w12264, w12265, w12266, w12267, w12268, w12269, w12270, w12271, w12272, w12273, w12274, w12275, w12276, w12277, w12278, w12279, w12280, w12281, w12282, w12283, w12284, w12285, w12286, w12287, w12288, w12289, w12290, w12291, w12292, w12293, w12294, w12295, w12296, w12297, w12298, w12299, w12300, w12301, w12302, w12303, w12304, w12305, w12306, w12307, w12308, w12309, w12310, w12311, w12312, w12313, w12314, w12315, w12316, w12317, w12318, w12319, w12320, w12321, w12322, w12323, w12324, w12325, w12326, w12327, w12328, w12329, w12330, w12331, w12332, w12333, w12334, w12335, w12336, w12337, w12338, w12339, w12340, w12341, w12342, w12343, w12344, w12345, w12346, w12347, w12348, w12349, w12350, w12351, w12352, w12353, w12354, w12355, w12356, w12357, w12358, w12359, w12360, w12361, w12362, w12363, w12364, w12365, w12366, w12367, w12368, w12369, w12370, w12371, w12372, w12373, w12374, w12375, w12376, w12377, w12378, w12379, w12380, w12381, w12382, w12383, w12384, w12385, w12386, w12387, w12388, w12389, w12390, w12391, w12392, w12393, w12394, w12395, w12396, w12397, w12398, w12399, w12400, w12401, w12402, w12403, w12404, w12405, w12406, w12407, w12408, w12409, w12410, w12411, w12412, w12413, w12414, w12415, w12416, w12417, w12418, w12419, w12420, w12421, w12422, w12423, w12424, w12425, w12426, w12427, w12428, w12429, w12430, w12431, w12432, w12433, w12434, w12435, w12436, w12437, w12438, w12439, w12440, w12441, w12442, w12443, w12444, w12445, w12446, w12447, w12448, w12449, w12450, w12451, w12452, w12453, w12454, w12455, w12456, w12457, w12458, w12459, w12460, w12461, w12462, w12463, w12464, w12465, w12466, w12467, w12468, w12469, w12470, w12471, w12472, w12473, w12474, w12475, w12476, w12477, w12478, w12479, w12480, w12481, w12482, w12483, w12484, w12485, w12486, w12487, w12488, w12489, w12490, w12491, w12492, w12493, w12494, w12495, w12496, w12497, w12498, w12499, w12500, w12501, w12502, w12503, w12504, w12505, w12506, w12507, w12508, w12509, w12510, w12511, w12512, w12513, w12514, w12515, w12516, w12517, w12518, w12519, w12520, w12521, w12522, w12523, w12524, w12525, w12526, w12527, w12528, w12529, w12530, w12531, w12532, w12533, w12534, w12535, w12536, w12537, w12538, w12539, w12540, w12541, w12542, w12543, w12544, w12545, w12546, w12547, w12548, w12549, w12550, w12551, w12552, w12553, w12554, w12555, w12556, w12557, w12558, w12559, w12560, w12561, w12562, w12563, w12564, w12565, w12566, w12567, w12568, w12569, w12570, w12571, w12572, w12573, w12574, w12575, w12576, w12577, w12578, w12579, w12580, w12581, w12582, w12583, w12584, w12585, w12586, w12587, w12588, w12589, w12590, w12591, w12592, w12593, w12594, w12595, w12596, w12597, w12598, w12599, w12600, w12601, w12602, w12603, w12604, w12605, w12606, w12607, w12608, w12609, w12610, w12611, w12612, w12613, w12614, w12615, w12616, w12617, w12618, w12619, w12620, w12621, w12622, w12623, w12624, w12625, w12626, w12627, w12628, w12629, w12630, w12631, w12632, w12633, w12634, w12635, w12636, w12637, w12638, w12639, w12640, w12641, w12642, w12643, w12644, w12645, w12646, w12647, w12648, w12649, w12650, w12651, w12652, w12653, w12654, w12655, w12656, w12657, w12658, w12659, w12660, w12661, w12662, w12663, w12664, w12665, w12666, w12667, w12668, w12669, w12670, w12671, w12672, w12673, w12674, w12675, w12676, w12677, w12678, w12679, w12680, w12681, w12682, w12683, w12684, w12685, w12686, w12687, w12688, w12689, w12690, w12691, w12692, w12693, w12694, w12695, w12696, w12697, w12698, w12699, w12700, w12701, w12702, w12703, w12704, w12705, w12706, w12707, w12708, w12709, w12710, w12711, w12712, w12713, w12714, w12715, w12716, w12717, w12718, w12719, w12720, w12721, w12722, w12723, w12724, w12725, w12726, w12727, w12728, w12729, w12730, w12731, w12732, w12733, w12734, w12735, w12736, w12737, w12738, w12739, w12740, w12741, w12742, w12743, w12744, w12745, w12746, w12747, w12748, w12749, w12750, w12751, w12752, w12753, w12754, w12755, w12756, w12757, w12758, w12759, w12760, w12761, w12762, w12763, w12764, w12765, w12766, w12767, w12768, w12769, w12770, w12771, w12772, w12773, w12774, w12775, w12776, w12777, w12778, w12779, w12780, w12781, w12782, w12783, w12784, w12785, w12786, w12787, w12788, w12789, w12790, w12791, w12792, w12793, w12794, w12795, w12796, w12797, w12798, w12799, w12800, w12801, w12802, w12803, w12804, w12805, w12806, w12807, w12808, w12809, w12810, w12811, w12812, w12813, w12814, w12815, w12816, w12817, w12818, w12819, w12820, w12821, w12822, w12823, w12824, w12825, w12826, w12827, w12828, w12829, w12830, w12831, w12832, w12833, w12834, w12835, w12836, w12837, w12838, w12839, w12840, w12841, w12842, w12843, w12844, w12845, w12846, w12847, w12848, w12849, w12850, w12851, w12852, w12853, w12854, w12855, w12856, w12857, w12858, w12859, w12860, w12861, w12862, w12863, w12864, w12865, w12866, w12867, w12868, w12869, w12870, w12871, w12872, w12873, w12874, w12875, w12876, w12877, w12878, w12879, w12880, w12881, w12882, w12883, w12884, w12885, w12886, w12887, w12888, w12889, w12890, w12891, w12892, w12893, w12894, w12895, w12896, w12897, w12898, w12899, w12900, w12901, w12902, w12903, w12904, w12905, w12906, w12907, w12908, w12909, w12910, w12911, w12912, w12913, w12914, w12915, w12916, w12917, w12918, w12919, w12920, w12921, w12922, w12923, w12924, w12925, w12926, w12927, w12928, w12929, w12930, w12931, w12932, w12933, w12934, w12935, w12936, w12937, w12938, w12939, w12940, w12941, w12942, w12943, w12944, w12945, w12946, w12947, w12948, w12949, w12950, w12951, w12952, w12953, w12954, w12955, w12956, w12957, w12958, w12959, w12960, w12961, w12962, w12963, w12964, w12965, w12966, w12967, w12968, w12969, w12970, w12971, w12972, w12973, w12974, w12975, w12976, w12977, w12978, w12979, w12980, w12981, w12982, w12983, w12984, w12985, w12986, w12987, w12988, w12989, w12990, w12991, w12992, w12993, w12994, w12995, w12996, w12997, w12998, w12999, w13000, w13001, w13002, w13003, w13004, w13005, w13006, w13007, w13008, w13009, w13010, w13011, w13012, w13013, w13014, w13015, w13016, w13017, w13018, w13019, w13020, w13021, w13022, w13023, w13024, w13025, w13026, w13027, w13028, w13029, w13030, w13031, w13032, w13033, w13034, w13035, w13036, w13037, w13038, w13039, w13040, w13041, w13042, w13043, w13044, w13045, w13046, w13047, w13048, w13049, w13050, w13051, w13052, w13053, w13054, w13055, w13056, w13057, w13058, w13059, w13060, w13061, w13062, w13063, w13064, w13065, w13066, w13067, w13068, w13069, w13070, w13071, w13072, w13073, w13074, w13075, w13076, w13077, w13078, w13079, w13080, w13081, w13082, w13083, w13084, w13085, w13086, w13087, w13088, w13089, w13090, w13091, w13092, w13093, w13094, w13095, w13096, w13097, w13098, w13099, w13100, w13101, w13102, w13103, w13104, w13105, w13106, w13107, w13108, w13109, w13110, w13111, w13112, w13113, w13114, w13115, w13116, w13117, w13118, w13119, w13120, w13121, w13122, w13123, w13124, w13125, w13126, w13127, w13128, w13129, w13130, w13131, w13132, w13133, w13134, w13135, w13136, w13137, w13138, w13139, w13140, w13141, w13142, w13143, w13144, w13145, w13146, w13147, w13148, w13149, w13150, w13151, w13152, w13153, w13154, w13155, w13156, w13157, w13158, w13159, w13160, w13161, w13162, w13163, w13164, w13165, w13166, w13167, w13168, w13169, w13170, w13171, w13172, w13173, w13174, w13175, w13176, w13177, w13178, w13179, w13180, w13181, w13182, w13183, w13184, w13185, w13186, w13187, w13188, w13189, w13190, w13191, w13192, w13193, w13194, w13195, w13196, w13197, w13198, w13199, w13200, w13201, w13202, w13203, w13204, w13205, w13206, w13207, w13208, w13209, w13210, w13211, w13212, w13213, w13214, w13215, w13216, w13217, w13218, w13219, w13220, w13221, w13222, w13223, w13224, w13225, w13226, w13227, w13228, w13229, w13230, w13231, w13232, w13233, w13234, w13235, w13236, w13237, w13238, w13239, w13240, w13241, w13242, w13243, w13244, w13245, w13246, w13247, w13248, w13249, w13250, w13251, w13252, w13253, w13254, w13255, w13256, w13257, w13258, w13259, w13260, w13261, w13262, w13263, w13264, w13265, w13266, w13267, w13268, w13269, w13270, w13271, w13272, w13273, w13274, w13275, w13276, w13277, w13278, w13279, w13280, w13281, w13282, w13283, w13284, w13285, w13286, w13287, w13288, w13289, w13290, w13291, w13292, w13293, w13294, w13295, w13296, w13297, w13298, w13299, w13300, w13301, w13302, w13303, w13304, w13305, w13306, w13307, w13308, w13309, w13310, w13311, w13312, w13313, w13314, w13315, w13316, w13317, w13318, w13319, w13320, w13321, w13322, w13323, w13324, w13325, w13326, w13327, w13328, w13329, w13330, w13331, w13332, w13333, w13334, w13335, w13336, w13337, w13338, w13339, w13340, w13341, w13342, w13343, w13344, w13345, w13346, w13347, w13348, w13349, w13350, w13351, w13352, w13353, w13354, w13355, w13356, w13357, w13358, w13359, w13360, w13361, w13362, w13363, w13364, w13365, w13366, w13367, w13368, w13369, w13370, w13371, w13372, w13373, w13374, w13375, w13376, w13377, w13378, w13379, w13380, w13381, w13382, w13383, w13384, w13385, w13386, w13387, w13388, w13389, w13390, w13391, w13392, w13393, w13394, w13395, w13396, w13397, w13398, w13399, w13400, w13401, w13402, w13403, w13404, w13405, w13406, w13407, w13408, w13409, w13410, w13411, w13412, w13413, w13414, w13415, w13416, w13417, w13418, w13419, w13420, w13421, w13422, w13423, w13424, w13425, w13426, w13427, w13428, w13429, w13430, w13431, w13432, w13433, w13434, w13435, w13436, w13437, w13438, w13439, w13440, w13441, w13442, w13443, w13444, w13445, w13446, w13447, w13448, w13449, w13450, w13451, w13452, w13453, w13454, w13455, w13456, w13457, w13458, w13459, w13460, w13461, w13462, w13463, w13464, w13465, w13466, w13467, w13468, w13469, w13470, w13471, w13472, w13473, w13474, w13475, w13476, w13477, w13478, w13479, w13480, w13481, w13482, w13483, w13484, w13485, w13486, w13487, w13488, w13489, w13490, w13491, w13492, w13493, w13494, w13495, w13496, w13497, w13498, w13499, w13500, w13501, w13502, w13503, w13504, w13505, w13506, w13507, w13508, w13509, w13510, w13511, w13512, w13513, w13514, w13515, w13516, w13517, w13518, w13519, w13520, w13521, w13522, w13523, w13524, w13525, w13526, w13527, w13528, w13529, w13530, w13531, w13532, w13533, w13534, w13535, w13536, w13537, w13538, w13539, w13540, w13541, w13542, w13543, w13544, w13545, w13546, w13547, w13548, w13549, w13550, w13551, w13552, w13553, w13554, w13555, w13556, w13557, w13558, w13559, w13560, w13561, w13562, w13563, w13564, w13565, w13566, w13567, w13568, w13569, w13570, w13571, w13572, w13573, w13574, w13575, w13576, w13577, w13578, w13579, w13580, w13581, w13582, w13583, w13584, w13585, w13586, w13587, w13588, w13589, w13590, w13591, w13592, w13593, w13594, w13595, w13596, w13597, w13598, w13599, w13600, w13601, w13602, w13603, w13604, w13605, w13606, w13607, w13608, w13609, w13610, w13611, w13612, w13613, w13614, w13615, w13616, w13617, w13618, w13619, w13620, w13621, w13622, w13623, w13624, w13625, w13626, w13627, w13628, w13629, w13630, w13631, w13632, w13633, w13634, w13635, w13636, w13637, w13638, w13639, w13640, w13641, w13642, w13643, w13644, w13645, w13646, w13647, w13648, w13649, w13650, w13651, w13652, w13653, w13654, w13655, w13656, w13657, w13658, w13659, w13660, w13661, w13662, w13663, w13664, w13665, w13666, w13667, w13668, w13669, w13670, w13671, w13672, w13673, w13674, w13675, w13676, w13677, w13678, w13679, w13680, w13681, w13682, w13683, w13684, w13685, w13686, w13687, w13688, w13689, w13690, w13691, w13692, w13693, w13694, w13695, w13696, w13697, w13698, w13699, w13700, w13701, w13702, w13703, w13704, w13705, w13706, w13707, w13708, w13709, w13710, w13711, w13712, w13713, w13714, w13715, w13716, w13717, w13718, w13719, w13720, w13721, w13722, w13723, w13724, w13725, w13726, w13727, w13728, w13729, w13730, w13731, w13732, w13733, w13734, w13735, w13736, w13737, w13738, w13739, w13740, w13741, w13742, w13743, w13744, w13745, w13746, w13747, w13748, w13749, w13750, w13751, w13752, w13753, w13754, w13755, w13756, w13757, w13758, w13759, w13760, w13761, w13762, w13763, w13764, w13765, w13766, w13767, w13768, w13769, w13770, w13771, w13772, w13773, w13774, w13775, w13776, w13777, w13778, w13779, w13780, w13781, w13782, w13783, w13784, w13785, w13786, w13787, w13788, w13789, w13790, w13791, w13792, w13793, w13794, w13795, w13796, w13797, w13798, w13799, w13800, w13801, w13802, w13803, w13804, w13805, w13806, w13807, w13808, w13809, w13810, w13811, w13812, w13813, w13814, w13815, w13816, w13817, w13818, w13819, w13820, w13821, w13822, w13823, w13824, w13825, w13826, w13827, w13828, w13829, w13830, w13831, w13832, w13833, w13834, w13835, w13836, w13837, w13838, w13839, w13840, w13841, w13842, w13843, w13844, w13845, w13846, w13847, w13848, w13849, w13850, w13851, w13852, w13853, w13854, w13855, w13856, w13857, w13858, w13859, w13860, w13861, w13862, w13863, w13864, w13865, w13866, w13867, w13868, w13869, w13870, w13871, w13872, w13873, w13874, w13875, w13876, w13877, w13878, w13879, w13880, w13881, w13882, w13883, w13884, w13885, w13886, w13887, w13888, w13889, w13890, w13891, w13892, w13893, w13894, w13895, w13896, w13897, w13898, w13899, w13900, w13901, w13902, w13903, w13904, w13905, w13906, w13907, w13908, w13909, w13910, w13911, w13912, w13913, w13914, w13915, w13916, w13917, w13918, w13919, w13920, w13921, w13922, w13923, w13924, w13925, w13926, w13927, w13928, w13929, w13930, w13931, w13932, w13933, w13934, w13935, w13936, w13937, w13938, w13939, w13940, w13941, w13942, w13943, w13944, w13945, w13946, w13947, w13948, w13949, w13950, w13951, w13952, w13953, w13954, w13955, w13956, w13957, w13958, w13959, w13960, w13961, w13962, w13963, w13964, w13965, w13966, w13967, w13968, w13969, w13970, w13971, w13972, w13973, w13974, w13975, w13976, w13977, w13978, w13979, w13980, w13981, w13982, w13983, w13984, w13985, w13986, w13987, w13988, w13989, w13990, w13991, w13992, w13993, w13994, w13995, w13996, w13997, w13998, w13999, w14000, w14001, w14002, w14003, w14004, w14005, w14006, w14007, w14008, w14009, w14010, w14011, w14012, w14013, w14014, w14015, w14016, w14017, w14018, w14019, w14020, w14021, w14022, w14023, w14024, w14025, w14026, w14027, w14028, w14029, w14030, w14031, w14032, w14033, w14034, w14035, w14036, w14037, w14038, w14039, w14040, w14041, w14042, w14043, w14044, w14045, w14046, w14047, w14048, w14049, w14050, w14051, w14052, w14053, w14054, w14055, w14056, w14057, w14058, w14059, w14060, w14061, w14062, w14063, w14064, w14065, w14066, w14067, w14068, w14069, w14070, w14071, w14072, w14073, w14074, w14075, w14076, w14077, w14078, w14079, w14080, w14081, w14082, w14083, w14084, w14085, w14086, w14087, w14088, w14089, w14090, w14091, w14092, w14093, w14094, w14095, w14096, w14097, w14098, w14099, w14100, w14101, w14102, w14103, w14104, w14105, w14106, w14107, w14108, w14109, w14110, w14111, w14112, w14113, w14114, w14115, w14116, w14117, w14118, w14119, w14120, w14121, w14122, w14123, w14124, w14125, w14126, w14127, w14128, w14129, w14130, w14131, w14132, w14133, w14134, w14135, w14136, w14137, w14138, w14139, w14140, w14141, w14142, w14143, w14144, w14145, w14146, w14147, w14148, w14149, w14150, w14151, w14152, w14153, w14154, w14155, w14156, w14157, w14158, w14159, w14160, w14161, w14162, w14163, w14164, w14165, w14166, w14167, w14168, w14169, w14170, w14171, w14172, w14173, w14174, w14175, w14176, w14177, w14178, w14179, w14180, w14181, w14182, w14183, w14184, w14185, w14186, w14187, w14188, w14189, w14190, w14191, w14192, w14193, w14194, w14195, w14196, w14197, w14198, w14199, w14200, w14201, w14202, w14203, w14204, w14205, w14206, w14207, w14208, w14209, w14210, w14211, w14212, w14213, w14214, w14215, w14216, w14217, w14218, w14219, w14220, w14221, w14222, w14223, w14224, w14225, w14226, w14227, w14228, w14229, w14230, w14231, w14232, w14233, w14234, w14235, w14236, w14237, w14238, w14239, w14240, w14241, w14242, w14243, w14244, w14245, w14246, w14247, w14248, w14249, w14250, w14251, w14252, w14253, w14254, w14255, w14256, w14257, w14258, w14259, w14260, w14261, w14262, w14263, w14264, w14265, w14266, w14267, w14268, w14269, w14270, w14271, w14272, w14273, w14274, w14275, w14276, w14277, w14278, w14279, w14280, w14281, w14282, w14283, w14284, w14285, w14286, w14287, w14288, w14289, w14290, w14291, w14292, w14293, w14294, w14295, w14296, w14297, w14298, w14299, w14300, w14301, w14302, w14303, w14304, w14305, w14306, w14307, w14308, w14309, w14310, w14311, w14312, w14313, w14314, w14315, w14316, w14317, w14318, w14319, w14320, w14321, w14322, w14323, w14324, w14325, w14326, w14327, w14328, w14329, w14330, w14331, w14332, w14333, w14334, w14335, w14336, w14337, w14338, w14339, w14340, w14341, w14342, w14343, w14344, w14345, w14346, w14347, w14348, w14349, w14350, w14351, w14352, w14353, w14354, w14355, w14356, w14357, w14358, w14359, w14360, w14361, w14362, w14363, w14364, w14365, w14366, w14367, w14368, w14369, w14370, w14371, w14372, w14373, w14374, w14375, w14376, w14377, w14378, w14379, w14380, w14381, w14382, w14383, w14384, w14385, w14386, w14387, w14388, w14389, w14390, w14391, w14392, w14393, w14394, w14395, w14396, w14397, w14398, w14399, w14400, w14401, w14402, w14403, w14404, w14405, w14406, w14407, w14408, w14409, w14410, w14411, w14412, w14413, w14414, w14415, w14416, w14417, w14418, w14419, w14420, w14421, w14422, w14423, w14424, w14425, w14426, w14427, w14428, w14429, w14430, w14431, w14432, w14433, w14434, w14435, w14436, w14437, w14438, w14439, w14440, w14441, w14442, w14443, w14444, w14445, w14446, w14447, w14448, w14449, w14450, w14451, w14452, w14453, w14454, w14455, w14456, w14457, w14458, w14459, w14460, w14461, w14462, w14463, w14464, w14465, w14466, w14467, w14468, w14469, w14470, w14471, w14472, w14473, w14474, w14475, w14476, w14477, w14478, w14479, w14480, w14481, w14482, w14483, w14484, w14485, w14486, w14487, w14488, w14489, w14490, w14491, w14492, w14493, w14494, w14495, w14496, w14497, w14498, w14499, w14500, w14501, w14502, w14503, w14504, w14505, w14506, w14507, w14508, w14509, w14510, w14511, w14512, w14513, w14514, w14515, w14516, w14517, w14518, w14519, w14520, w14521, w14522, w14523, w14524, w14525, w14526, w14527, w14528, w14529, w14530, w14531, w14532, w14533, w14534, w14535, w14536, w14537, w14538, w14539, w14540, w14541, w14542, w14543, w14544, w14545, w14546, w14547, w14548, w14549, w14550, w14551, w14552, w14553, w14554, w14555, w14556, w14557, w14558, w14559, w14560, w14561, w14562, w14563, w14564, w14565, w14566, w14567, w14568, w14569, w14570, w14571, w14572, w14573, w14574, w14575, w14576, w14577, w14578, w14579, w14580, w14581, w14582, w14583, w14584, w14585, w14586, w14587, w14588, w14589, w14590, w14591, w14592, w14593, w14594, w14595, w14596, w14597, w14598, w14599, w14600, w14601, w14602, w14603, w14604, w14605, w14606, w14607, w14608, w14609, w14610, w14611, w14612, w14613, w14614, w14615, w14616, w14617, w14618, w14619, w14620, w14621, w14622, w14623, w14624, w14625, w14626, w14627, w14628, w14629, w14630, w14631, w14632, w14633, w14634, w14635, w14636, w14637, w14638, w14639, w14640, w14641, w14642, w14643, w14644, w14645, w14646, w14647, w14648, w14649, w14650, w14651, w14652, w14653, w14654, w14655, w14656, w14657, w14658, w14659, w14660, w14661, w14662, w14663, w14664, w14665, w14666, w14667, w14668, w14669, w14670, w14671, w14672, w14673, w14674, w14675, w14676, w14677, w14678, w14679, w14680, w14681, w14682, w14683, w14684, w14685, w14686, w14687, w14688, w14689, w14690, w14691, w14692, w14693, w14694, w14695, w14696, w14697, w14698, w14699, w14700, w14701, w14702, w14703, w14704, w14705, w14706, w14707, w14708, w14709, w14710, w14711, w14712, w14713, w14714, w14715, w14716, w14717, w14718, w14719, w14720, w14721, w14722, w14723, w14724, w14725, w14726, w14727, w14728, w14729, w14730, w14731, w14732, w14733, w14734, w14735, w14736, w14737, w14738, w14739, w14740, w14741, w14742, w14743, w14744, w14745, w14746, w14747, w14748, w14749, w14750, w14751, w14752, w14753, w14754, w14755, w14756, w14757, w14758, w14759, w14760, w14761, w14762, w14763, w14764, w14765, w14766, w14767, w14768, w14769, w14770, w14771, w14772, w14773, w14774, w14775, w14776, w14777, w14778, w14779, w14780, w14781, w14782, w14783, w14784, w14785, w14786, w14787, w14788, w14789, w14790, w14791, w14792, w14793, w14794, w14795, w14796, w14797, w14798, w14799, w14800, w14801, w14802, w14803, w14804, w14805, w14806, w14807, w14808, w14809, w14810, w14811, w14812, w14813, w14814, w14815, w14816, w14817, w14818, w14819, w14820, w14821, w14822, w14823, w14824, w14825, w14826, w14827, w14828, w14829, w14830, w14831, w14832, w14833, w14834, w14835, w14836, w14837, w14838, w14839, w14840, w14841, w14842, w14843, w14844, w14845, w14846, w14847, w14848, w14849, w14850, w14851, w14852, w14853, w14854, w14855, w14856, w14857, w14858, w14859, w14860, w14861, w14862, w14863, w14864, w14865, w14866, w14867, w14868, w14869, w14870, w14871, w14872, w14873, w14874, w14875, w14876, w14877, w14878, w14879, w14880, w14881, w14882, w14883, w14884, w14885, w14886, w14887, w14888, w14889, w14890, w14891, w14892, w14893, w14894, w14895, w14896, w14897, w14898, w14899, w14900, w14901, w14902, w14903, w14904, w14905, w14906, w14907, w14908, w14909, w14910, w14911, w14912, w14913, w14914, w14915, w14916, w14917, w14918, w14919, w14920, w14921, w14922, w14923, w14924, w14925, w14926, w14927, w14928, w14929, w14930, w14931, w14932, w14933, w14934, w14935, w14936, w14937, w14938, w14939, w14940, w14941, w14942, w14943, w14944, w14945, w14946, w14947, w14948, w14949, w14950, w14951, w14952, w14953, w14954, w14955, w14956, w14957, w14958, w14959, w14960, w14961, w14962, w14963, w14964, w14965, w14966, w14967, w14968, w14969, w14970, w14971, w14972, w14973, w14974, w14975, w14976, w14977, w14978, w14979, w14980, w14981, w14982, w14983, w14984, w14985, w14986, w14987, w14988, w14989, w14990, w14991, w14992, w14993, w14994, w14995, w14996, w14997, w14998, w14999, w15000, w15001, w15002, w15003, w15004, w15005, w15006, w15007, w15008, w15009, w15010, w15011, w15012, w15013, w15014, w15015, w15016, w15017, w15018, w15019, w15020, w15021, w15022, w15023, w15024, w15025, w15026, w15027, w15028, w15029, w15030, w15031, w15032, w15033, w15034, w15035, w15036, w15037, w15038, w15039, w15040, w15041, w15042, w15043, w15044, w15045, w15046, w15047, w15048, w15049, w15050, w15051, w15052, w15053, w15054, w15055, w15056, w15057, w15058, w15059, w15060, w15061, w15062, w15063, w15064, w15065, w15066, w15067, w15068, w15069, w15070, w15071, w15072, w15073, w15074, w15075, w15076, w15077, w15078, w15079, w15080, w15081, w15082, w15083, w15084, w15085, w15086, w15087, w15088, w15089, w15090, w15091, w15092, w15093, w15094, w15095, w15096, w15097, w15098, w15099, w15100, w15101, w15102, w15103, w15104, w15105, w15106, w15107, w15108, w15109, w15110, w15111, w15112, w15113, w15114, w15115, w15116, w15117, w15118, w15119, w15120, w15121, w15122, w15123, w15124, w15125, w15126, w15127, w15128, w15129, w15130, w15131, w15132, w15133, w15134, w15135, w15136, w15137, w15138, w15139, w15140, w15141, w15142, w15143, w15144, w15145, w15146, w15147, w15148, w15149, w15150, w15151, w15152, w15153, w15154, w15155, w15156, w15157, w15158, w15159, w15160, w15161, w15162, w15163, w15164, w15165, w15166, w15167, w15168, w15169, w15170, w15171, w15172, w15173, w15174, w15175, w15176, w15177, w15178, w15179, w15180, w15181, w15182, w15183, w15184, w15185, w15186, w15187, w15188, w15189, w15190, w15191, w15192, w15193, w15194, w15195, w15196, w15197, w15198, w15199, w15200, w15201, w15202, w15203, w15204, w15205, w15206, w15207, w15208, w15209, w15210, w15211, w15212, w15213, w15214, w15215, w15216, w15217, w15218, w15219, w15220, w15221, w15222, w15223, w15224, w15225, w15226, w15227, w15228, w15229, w15230, w15231, w15232, w15233, w15234, w15235, w15236, w15237, w15238, w15239, w15240, w15241, w15242, w15243, w15244, w15245, w15246, w15247, w15248, w15249, w15250, w15251, w15252, w15253, w15254, w15255, w15256, w15257, w15258, w15259, w15260, w15261, w15262, w15263, w15264, w15265, w15266, w15267, w15268, w15269, w15270, w15271, w15272, w15273, w15274, w15275, w15276, w15277, w15278, w15279, w15280, w15281, w15282, w15283, w15284, w15285, w15286, w15287, w15288, w15289, w15290, w15291, w15292, w15293, w15294, w15295, w15296, w15297, w15298, w15299, w15300, w15301, w15302, w15303, w15304, w15305, w15306, w15307, w15308, w15309, w15310, w15311, w15312, w15313, w15314, w15315, w15316, w15317, w15318, w15319, w15320, w15321, w15322, w15323, w15324, w15325, w15326, w15327, w15328, w15329, w15330, w15331, w15332, w15333, w15334, w15335, w15336, w15337, w15338, w15339, w15340, w15341, w15342, w15343, w15344, w15345, w15346, w15347, w15348, w15349, w15350, w15351, w15352, w15353, w15354, w15355, w15356, w15357, w15358, w15359, w15360, w15361, w15362, w15363, w15364, w15365, w15366, w15367, w15368, w15369, w15370, w15371, w15372, w15373, w15374, w15375, w15376, w15377, w15378, w15379, w15380, w15381, w15382, w15383, w15384, w15385, w15386, w15387, w15388, w15389, w15390, w15391, w15392, w15393, w15394, w15395, w15396, w15397, w15398, w15399, w15400, w15401, w15402, w15403, w15404, w15405, w15406, w15407, w15408, w15409, w15410, w15411, w15412, w15413, w15414, w15415, w15416, w15417, w15418, w15419, w15420, w15421, w15422, w15423, w15424, w15425, w15426, w15427, w15428, w15429, w15430, w15431, w15432, w15433, w15434, w15435, w15436, w15437, w15438, w15439, w15440, w15441, w15442, w15443, w15444, w15445, w15446, w15447, w15448, w15449, w15450, w15451, w15452, w15453, w15454, w15455, w15456, w15457, w15458, w15459, w15460, w15461, w15462, w15463, w15464, w15465, w15466, w15467, w15468, w15469, w15470, w15471, w15472, w15473, w15474, w15475, w15476, w15477, w15478, w15479, w15480, w15481, w15482, w15483, w15484, w15485, w15486, w15487, w15488, w15489, w15490, w15491, w15492, w15493, w15494, w15495, w15496, w15497, w15498, w15499, w15500, w15501, w15502, w15503, w15504, w15505, w15506, w15507, w15508, w15509, w15510, w15511, w15512, w15513, w15514, w15515, w15516, w15517, w15518, w15519, w15520, w15521, w15522, w15523, w15524, w15525, w15526, w15527, w15528, w15529, w15530, w15531, w15532, w15533, w15534, w15535, w15536, w15537, w15538, w15539, w15540, w15541, w15542, w15543, w15544, w15545, w15546, w15547, w15548, w15549, w15550, w15551, w15552, w15553, w15554, w15555, w15556, w15557, w15558, w15559, w15560, w15561, w15562, w15563, w15564, w15565, w15566, w15567, w15568, w15569, w15570, w15571, w15572, w15573, w15574, w15575, w15576, w15577, w15578, w15579, w15580, w15581, w15582, w15583, w15584, w15585, w15586, w15587, w15588, w15589, w15590, w15591, w15592, w15593, w15594, w15595, w15596, w15597, w15598, w15599, w15600, w15601, w15602, w15603, w15604, w15605, w15606, w15607, w15608, w15609, w15610, w15611, w15612, w15613, w15614, w15615, w15616, w15617, w15618, w15619, w15620, w15621, w15622, w15623, w15624, w15625, w15626, w15627, w15628, w15629, w15630, w15631, w15632, w15633, w15634, w15635, w15636, w15637, w15638, w15639, w15640, w15641, w15642, w15643, w15644, w15645, w15646, w15647, w15648, w15649, w15650, w15651, w15652, w15653, w15654, w15655, w15656, w15657, w15658, w15659, w15660, w15661, w15662, w15663, w15664, w15665, w15666, w15667, w15668, w15669, w15670, w15671, w15672, w15673, w15674, w15675, w15676, w15677, w15678, w15679, w15680, w15681, w15682, w15683, w15684, w15685, w15686, w15687, w15688, w15689, w15690, w15691, w15692, w15693, w15694, w15695, w15696, w15697, w15698, w15699, w15700, w15701, w15702, w15703, w15704, w15705, w15706, w15707, w15708, w15709, w15710, w15711, w15712, w15713, w15714, w15715, w15716, w15717, w15718, w15719, w15720, w15721, w15722, w15723, w15724, w15725, w15726, w15727, w15728, w15729, w15730, w15731, w15732, w15733, w15734, w15735, w15736, w15737, w15738, w15739, w15740, w15741, w15742, w15743, w15744, w15745, w15746, w15747, w15748, w15749, w15750, w15751, w15752, w15753, w15754, w15755, w15756, w15757, w15758, w15759, w15760, w15761, w15762, w15763, w15764, w15765, w15766, w15767, w15768, w15769, w15770, w15771, w15772, w15773, w15774, w15775, w15776, w15777, w15778, w15779, w15780, w15781, w15782, w15783, w15784, w15785, w15786, w15787, w15788, w15789, w15790, w15791, w15792, w15793, w15794, w15795, w15796, w15797, w15798, w15799, w15800, w15801, w15802, w15803, w15804, w15805, w15806, w15807, w15808, w15809, w15810, w15811, w15812, w15813, w15814, w15815, w15816, w15817, w15818, w15819, w15820, w15821, w15822, w15823, w15824, w15825, w15826, w15827, w15828, w15829, w15830, w15831, w15832, w15833, w15834, w15835, w15836, w15837, w15838, w15839, w15840, w15841, w15842, w15843, w15844, w15845, w15846, w15847, w15848, w15849, w15850, w15851, w15852, w15853, w15854, w15855, w15856, w15857, w15858, w15859, w15860, w15861, w15862, w15863, w15864, w15865, w15866, w15867, w15868, w15869, w15870, w15871, w15872, w15873, w15874, w15875, w15876, w15877, w15878, w15879, w15880, w15881, w15882, w15883, w15884, w15885, w15886, w15887, w15888, w15889, w15890, w15891, w15892, w15893, w15894, w15895, w15896, w15897, w15898, w15899, w15900, w15901, w15902, w15903, w15904, w15905, w15906, w15907, w15908, w15909, w15910, w15911, w15912, w15913, w15914, w15915, w15916, w15917, w15918, w15919, w15920, w15921, w15922, w15923, w15924, w15925, w15926, w15927, w15928, w15929, w15930, w15931, w15932, w15933, w15934, w15935, w15936, w15937, w15938, w15939, w15940, w15941, w15942, w15943, w15944, w15945, w15946, w15947, w15948, w15949, w15950, w15951, w15952, w15953, w15954, w15955, w15956, w15957, w15958, w15959, w15960, w15961, w15962, w15963, w15964, w15965, w15966, w15967, w15968, w15969, w15970, w15971, w15972, w15973, w15974, w15975, w15976, w15977, w15978, w15979, w15980, w15981, w15982, w15983, w15984, w15985, w15986, w15987, w15988, w15989, w15990, w15991, w15992, w15993, w15994, w15995, w15996, w15997, w15998, w15999, w16000, w16001, w16002, w16003, w16004, w16005, w16006, w16007, w16008, w16009, w16010, w16011, w16012, w16013, w16014, w16015, w16016, w16017, w16018, w16019, w16020, w16021, w16022, w16023, w16024, w16025, w16026, w16027, w16028, w16029, w16030, w16031, w16032, w16033, w16034, w16035, w16036, w16037, w16038, w16039, w16040, w16041, w16042, w16043, w16044, w16045, w16046, w16047, w16048, w16049, w16050, w16051, w16052, w16053, w16054, w16055, w16056, w16057, w16058, w16059, w16060, w16061, w16062, w16063, w16064, w16065, w16066, w16067, w16068, w16069, w16070, w16071, w16072, w16073, w16074, w16075, w16076, w16077, w16078, w16079, w16080, w16081, w16082, w16083, w16084, w16085, w16086, w16087, w16088, w16089, w16090, w16091, w16092, w16093, w16094, w16095, w16096, w16097, w16098, w16099, w16100, w16101, w16102, w16103, w16104, w16105, w16106, w16107, w16108, w16109, w16110, w16111, w16112, w16113, w16114, w16115, w16116, w16117, w16118, w16119, w16120, w16121, w16122, w16123, w16124, w16125, w16126, w16127, w16128, w16129, w16130, w16131, w16132, w16133, w16134, w16135, w16136, w16137, w16138, w16139, w16140, w16141, w16142, w16143, w16144, w16145, w16146, w16147, w16148, w16149, w16150, w16151, w16152, w16153, w16154, w16155, w16156, w16157, w16158, w16159, w16160, w16161, w16162, w16163, w16164, w16165, w16166, w16167, w16168, w16169, w16170, w16171, w16172, w16173, w16174, w16175, w16176, w16177, w16178, w16179, w16180, w16181, w16182, w16183, w16184, w16185, w16186, w16187, w16188, w16189, w16190, w16191, w16192, w16193, w16194, w16195, w16196, w16197, w16198, w16199, w16200, w16201, w16202, w16203, w16204, w16205, w16206, w16207, w16208, w16209, w16210, w16211, w16212, w16213, w16214, w16215, w16216, w16217, w16218, w16219, w16220, w16221, w16222, w16223, w16224, w16225, w16226, w16227, w16228, w16229, w16230, w16231, w16232, w16233, w16234, w16235, w16236, w16237, w16238, w16239, w16240, w16241, w16242, w16243, w16244, w16245, w16246, w16247, w16248, w16249, w16250, w16251, w16252, w16253, w16254, w16255, w16256, w16257, w16258, w16259, w16260, w16261, w16262, w16263, w16264, w16265, w16266, w16267, w16268, w16269, w16270, w16271, w16272, w16273, w16274, w16275, w16276, w16277, w16278, w16279, w16280, w16281, w16282, w16283, w16284, w16285, w16286, w16287, w16288, w16289, w16290, w16291, w16292, w16293, w16294, w16295, w16296, w16297, w16298, w16299, w16300, w16301, w16302, w16303, w16304, w16305, w16306, w16307, w16308, w16309, w16310, w16311, w16312, w16313, w16314, w16315, w16316, w16317, w16318, w16319, w16320, w16321, w16322, w16323, w16324, w16325, w16326, w16327, w16328, w16329, w16330, w16331, w16332, w16333, w16334, w16335, w16336, w16337, w16338, w16339, w16340, w16341, w16342, w16343, w16344, w16345, w16346, w16347, w16348, w16349, w16350, w16351, w16352, w16353, w16354, w16355, w16356, w16357, w16358, w16359, w16360, w16361, w16362, w16363, w16364, w16365, w16366, w16367, w16368, w16369, w16370, w16371, w16372, w16373, w16374, w16375, w16376, w16377, w16378, w16379, w16380, w16381, w16382, w16383, w16384, w16385, w16386, w16387, w16388, w16389, w16390, w16391, w16392, w16393, w16394, w16395, w16396, w16397, w16398, w16399, w16400, w16401, w16402, w16403, w16404, w16405, w16406, w16407, w16408, w16409, w16410, w16411, w16412, w16413, w16414, w16415, w16416, w16417, w16418, w16419, w16420, w16421, w16422, w16423, w16424, w16425, w16426, w16427, w16428, w16429, w16430, w16431, w16432, w16433, w16434, w16435, w16436, w16437, w16438, w16439, w16440, w16441, w16442, w16443, w16444, w16445, w16446, w16447, w16448, w16449, w16450, w16451, w16452, w16453, w16454, w16455, w16456, w16457, w16458, w16459, w16460, w16461, w16462, w16463, w16464, w16465, w16466, w16467, w16468, w16469, w16470, w16471, w16472, w16473, w16474, w16475, w16476, w16477, w16478, w16479, w16480, w16481, w16482, w16483, w16484, w16485, w16486, w16487, w16488, w16489, w16490, w16491, w16492, w16493, w16494, w16495, w16496, w16497, w16498, w16499, w16500, w16501, w16502, w16503, w16504, w16505, w16506, w16507, w16508, w16509, w16510, w16511, w16512, w16513, w16514, w16515, w16516, w16517, w16518, w16519, w16520, w16521, w16522, w16523, w16524, w16525, w16526, w16527, w16528, w16529, w16530, w16531, w16532, w16533, w16534, w16535, w16536, w16537, w16538, w16539, w16540, w16541, w16542, w16543, w16544, w16545, w16546, w16547, w16548, w16549, w16550, w16551, w16552, w16553, w16554, w16555, w16556, w16557, w16558, w16559, w16560, w16561, w16562, w16563, w16564, w16565, w16566, w16567, w16568, w16569, w16570, w16571, w16572, w16573, w16574, w16575, w16576, w16577, w16578, w16579, w16580, w16581, w16582, w16583, w16584, w16585, w16586, w16587, w16588, w16589, w16590, w16591, w16592, w16593, w16594, w16595, w16596, w16597, w16598, w16599, w16600, w16601, w16602, w16603, w16604, w16605, w16606, w16607, w16608, w16609, w16610, w16611, w16612, w16613, w16614, w16615, w16616, w16617, w16618, w16619, w16620, w16621, w16622, w16623, w16624, w16625, w16626, w16627, w16628, w16629, w16630, w16631, w16632, w16633, w16634, w16635, w16636, w16637, w16638, w16639, w16640, w16641, w16642, w16643, w16644, w16645, w16646, w16647, w16648, w16649, w16650, w16651, w16652, w16653, w16654, w16655, w16656, w16657, w16658, w16659, w16660, w16661, w16662, w16663, w16664, w16665, w16666, w16667, w16668, w16669, w16670, w16671, w16672, w16673, w16674, w16675, w16676, w16677, w16678, w16679, w16680, w16681, w16682, w16683, w16684, w16685, w16686, w16687, w16688, w16689, w16690, w16691, w16692, w16693, w16694, w16695, w16696, w16697, w16698, w16699, w16700, w16701, w16702, w16703, w16704, w16705, w16706, w16707, w16708, w16709, w16710, w16711, w16712, w16713, w16714, w16715, w16716, w16717, w16718, w16719, w16720, w16721, w16722, w16723, w16724, w16725, w16726, w16727, w16728, w16729, w16730, w16731, w16732, w16733, w16734, w16735, w16736, w16737, w16738, w16739, w16740, w16741, w16742, w16743, w16744, w16745, w16746, w16747, w16748, w16749, w16750, w16751, w16752, w16753, w16754, w16755, w16756, w16757, w16758, w16759, w16760, w16761, w16762, w16763, w16764, w16765, w16766, w16767, w16768, w16769, w16770, w16771, w16772, w16773, w16774, w16775, w16776, w16777, w16778, w16779, w16780, w16781, w16782, w16783, w16784, w16785, w16786, w16787, w16788, w16789, w16790, w16791, w16792, w16793, w16794, w16795, w16796, w16797, w16798, w16799, w16800, w16801, w16802, w16803, w16804, w16805, w16806, w16807, w16808, w16809, w16810, w16811, w16812, w16813, w16814, w16815, w16816, w16817, w16818, w16819, w16820, w16821, w16822, w16823, w16824, w16825, w16826, w16827, w16828, w16829, w16830, w16831, w16832, w16833, w16834, w16835, w16836, w16837, w16838, w16839, w16840, w16841, w16842, w16843, w16844, w16845, w16846, w16847, w16848, w16849, w16850, w16851, w16852, w16853, w16854, w16855, w16856, w16857, w16858, w16859, w16860, w16861, w16862, w16863, w16864, w16865, w16866, w16867, w16868, w16869, w16870, w16871, w16872, w16873, w16874, w16875, w16876, w16877, w16878, w16879, w16880, w16881, w16882, w16883, w16884, w16885, w16886, w16887, w16888, w16889, w16890, w16891, w16892, w16893, w16894, w16895, w16896, w16897, w16898, w16899, w16900, w16901, w16902, w16903, w16904, w16905, w16906, w16907, w16908, w16909, w16910, w16911, w16912, w16913, w16914, w16915, w16916, w16917, w16918, w16919, w16920, w16921, w16922, w16923, w16924, w16925, w16926, w16927, w16928, w16929, w16930, w16931, w16932, w16933, w16934, w16935, w16936, w16937, w16938, w16939, w16940, w16941, w16942, w16943, w16944, w16945, w16946, w16947, w16948, w16949, w16950, w16951, w16952, w16953, w16954, w16955, w16956, w16957, w16958, w16959, w16960, w16961, w16962, w16963, w16964, w16965, w16966, w16967, w16968, w16969, w16970, w16971, w16972, w16973, w16974, w16975, w16976, w16977, w16978, w16979, w16980, w16981, w16982, w16983, w16984, w16985, w16986, w16987, w16988, w16989, w16990, w16991, w16992, w16993, w16994, w16995, w16996, w16997, w16998, w16999, w17000, w17001, w17002, w17003, w17004, w17005, w17006, w17007, w17008, w17009, w17010, w17011, w17012, w17013, w17014, w17015, w17016, w17017, w17018, w17019, w17020, w17021, w17022, w17023, w17024, w17025, w17026, w17027, w17028, w17029, w17030, w17031, w17032, w17033, w17034, w17035, w17036, w17037, w17038, w17039, w17040, w17041, w17042, w17043, w17044, w17045, w17046, w17047, w17048, w17049, w17050, w17051, w17052, w17053, w17054, w17055, w17056, w17057, w17058, w17059, w17060, w17061, w17062, w17063, w17064, w17065, w17066, w17067, w17068, w17069, w17070, w17071, w17072, w17073, w17074, w17075, w17076, w17077, w17078, w17079, w17080, w17081, w17082, w17083, w17084, w17085, w17086, w17087, w17088, w17089, w17090, w17091, w17092, w17093, w17094, w17095, w17096, w17097, w17098, w17099, w17100, w17101, w17102, w17103, w17104, w17105, w17106, w17107, w17108, w17109, w17110, w17111, w17112, w17113, w17114, w17115, w17116, w17117, w17118, w17119, w17120, w17121, w17122, w17123, w17124, w17125, w17126, w17127, w17128, w17129, w17130, w17131, w17132, w17133, w17134, w17135, w17136, w17137, w17138, w17139, w17140, w17141, w17142, w17143, w17144, w17145, w17146, w17147, w17148, w17149, w17150, w17151, w17152, w17153, w17154, w17155, w17156, w17157, w17158, w17159, w17160, w17161, w17162, w17163, w17164, w17165, w17166, w17167, w17168, w17169, w17170, w17171, w17172, w17173, w17174, w17175, w17176, w17177, w17178, w17179, w17180, w17181, w17182, w17183, w17184, w17185, w17186, w17187, w17188, w17189, w17190, w17191, w17192, w17193, w17194, w17195, w17196, w17197, w17198, w17199, w17200, w17201, w17202, w17203, w17204, w17205, w17206, w17207, w17208, w17209, w17210, w17211, w17212, w17213, w17214, w17215, w17216, w17217, w17218, w17219, w17220, w17221, w17222, w17223, w17224, w17225, w17226, w17227, w17228, w17229, w17230, w17231, w17232, w17233, w17234, w17235, w17236, w17237, w17238, w17239, w17240, w17241, w17242, w17243, w17244, w17245, w17246, w17247, w17248, w17249, w17250, w17251, w17252, w17253, w17254, w17255, w17256, w17257, w17258, w17259, w17260, w17261, w17262, w17263, w17264, w17265, w17266, w17267, w17268, w17269, w17270, w17271, w17272, w17273, w17274, w17275, w17276, w17277, w17278, w17279, w17280, w17281, w17282, w17283, w17284, w17285, w17286, w17287, w17288, w17289, w17290, w17291, w17292, w17293, w17294, w17295, w17296, w17297, w17298, w17299, w17300, w17301, w17302, w17303, w17304, w17305, w17306, w17307, w17308, w17309, w17310, w17311, w17312, w17313, w17314, w17315, w17316, w17317, w17318, w17319, w17320, w17321, w17322, w17323, w17324, w17325, w17326, w17327, w17328, w17329, w17330, w17331, w17332, w17333, w17334, w17335, w17336, w17337, w17338, w17339, w17340, w17341, w17342, w17343, w17344, w17345, w17346, w17347, w17348, w17349, w17350, w17351, w17352, w17353, w17354, w17355, w17356, w17357, w17358, w17359, w17360, w17361, w17362, w17363, w17364, w17365, w17366, w17367, w17368, w17369, w17370, w17371, w17372, w17373, w17374, w17375, w17376, w17377, w17378, w17379, w17380, w17381, w17382, w17383, w17384, w17385, w17386, w17387, w17388, w17389, w17390, w17391, w17392, w17393, w17394, w17395, w17396, w17397, w17398, w17399, w17400, w17401, w17402, w17403, w17404, w17405, w17406, w17407, w17408, w17409, w17410, w17411, w17412, w17413, w17414, w17415, w17416, w17417, w17418, w17419, w17420, w17421, w17422, w17423, w17424, w17425, w17426, w17427, w17428, w17429, w17430, w17431, w17432, w17433, w17434, w17435, w17436, w17437, w17438, w17439, w17440, w17441, w17442, w17443, w17444, w17445, w17446, w17447, w17448, w17449, w17450, w17451, w17452, w17453, w17454, w17455, w17456, w17457, w17458, w17459, w17460, w17461, w17462, w17463, w17464, w17465, w17466, w17467, w17468, w17469, w17470, w17471, w17472, w17473, w17474, w17475, w17476, w17477, w17478, w17479, w17480, w17481, w17482, w17483, w17484, w17485, w17486, w17487, w17488, w17489, w17490, w17491, w17492, w17493, w17494, w17495, w17496, w17497, w17498, w17499, w17500, w17501, w17502, w17503, w17504, w17505, w17506, w17507, w17508, w17509, w17510, w17511, w17512, w17513, w17514, w17515, w17516, w17517, w17518, w17519, w17520, w17521, w17522, w17523, w17524, w17525, w17526, w17527, w17528, w17529, w17530, w17531, w17532, w17533, w17534, w17535, w17536, w17537, w17538, w17539, w17540, w17541, w17542, w17543, w17544, w17545, w17546, w17547, w17548, w17549, w17550, w17551, w17552, w17553, w17554, w17555, w17556, w17557, w17558, w17559, w17560, w17561, w17562, w17563, w17564, w17565, w17566, w17567, w17568, w17569, w17570, w17571, w17572, w17573, w17574, w17575, w17576, w17577, w17578, w17579, w17580, w17581, w17582, w17583, w17584, w17585, w17586, w17587, w17588, w17589, w17590, w17591, w17592, w17593, w17594, w17595, w17596, w17597, w17598, w17599, w17600, w17601, w17602, w17603, w17604, w17605, w17606, w17607, w17608, w17609, w17610, w17611, w17612, w17613, w17614, w17615, w17616, w17617, w17618, w17619, w17620, w17621, w17622, w17623, w17624, w17625, w17626, w17627, w17628, w17629, w17630, w17631, w17632, w17633, w17634, w17635, w17636, w17637, w17638, w17639, w17640, w17641, w17642, w17643, w17644, w17645, w17646, w17647, w17648, w17649, w17650, w17651, w17652, w17653, w17654, w17655, w17656, w17657, w17658, w17659, w17660, w17661, w17662, w17663, w17664, w17665, w17666, w17667, w17668, w17669, w17670, w17671, w17672, w17673, w17674, w17675, w17676, w17677, w17678, w17679, w17680, w17681, w17682, w17683, w17684, w17685, w17686, w17687, w17688, w17689, w17690, w17691, w17692, w17693, w17694, w17695, w17696, w17697, w17698, w17699, w17700, w17701, w17702, w17703, w17704, w17705, w17706, w17707, w17708, w17709, w17710, w17711, w17712, w17713, w17714, w17715, w17716, w17717, w17718, w17719, w17720, w17721, w17722, w17723, w17724, w17725, w17726, w17727, w17728, w17729, w17730, w17731, w17732, w17733, w17734, w17735, w17736, w17737, w17738, w17739, w17740, w17741, w17742, w17743, w17744, w17745, w17746, w17747, w17748, w17749, w17750, w17751, w17752, w17753, w17754, w17755, w17756, w17757, w17758, w17759, w17760, w17761, w17762, w17763, w17764, w17765, w17766, w17767, w17768, w17769, w17770, w17771, w17772, w17773, w17774, w17775, w17776, w17777, w17778, w17779, w17780, w17781, w17782, w17783, w17784, w17785, w17786, w17787, w17788, w17789, w17790, w17791, w17792, w17793, w17794, w17795, w17796, w17797, w17798, w17799, w17800, w17801, w17802, w17803, w17804, w17805, w17806, w17807, w17808, w17809, w17810, w17811, w17812, w17813, w17814, w17815, w17816, w17817, w17818, w17819, w17820, w17821, w17822, w17823, w17824, w17825, w17826, w17827, w17828, w17829, w17830, w17831, w17832, w17833, w17834, w17835, w17836, w17837, w17838, w17839, w17840, w17841, w17842, w17843, w17844, w17845, w17846, w17847, w17848, w17849, w17850, w17851, w17852, w17853, w17854, w17855, w17856, w17857, w17858, w17859, w17860, w17861, w17862, w17863, w17864, w17865, w17866, w17867, w17868, w17869, w17870, w17871, w17872, w17873, w17874, w17875, w17876, w17877, w17878, w17879, w17880, w17881, w17882, w17883, w17884, w17885, w17886, w17887, w17888, w17889, w17890, w17891, w17892, w17893, w17894, w17895, w17896, w17897, w17898, w17899, w17900, w17901, w17902, w17903, w17904, w17905, w17906, w17907, w17908, w17909, w17910, w17911, w17912, w17913, w17914, w17915, w17916, w17917, w17918, w17919, w17920, w17921, w17922, w17923, w17924, w17925, w17926, w17927, w17928, w17929, w17930, w17931, w17932, w17933, w17934, w17935, w17936, w17937, w17938, w17939, w17940, w17941, w17942, w17943, w17944, w17945, w17946, w17947, w17948, w17949, w17950, w17951, w17952, w17953, w17954, w17955, w17956, w17957, w17958, w17959, w17960, w17961, w17962, w17963, w17964, w17965, w17966, w17967, w17968, w17969, w17970, w17971, w17972, w17973, w17974, w17975, w17976, w17977, w17978, w17979, w17980, w17981, w17982, w17983, w17984, w17985, w17986, w17987, w17988, w17989, w17990, w17991, w17992, w17993, w17994, w17995, w17996, w17997, w17998, w17999, w18000, w18001, w18002, w18003, w18004, w18005, w18006, w18007, w18008, w18009, w18010, w18011, w18012, w18013, w18014, w18015, w18016, w18017, w18018, w18019, w18020, w18021, w18022, w18023, w18024, w18025, w18026, w18027, w18028, w18029, w18030, w18031, w18032, w18033, w18034, w18035, w18036, w18037, w18038, w18039, w18040, w18041, w18042, w18043, w18044, w18045, w18046, w18047, w18048, w18049, w18050, w18051, w18052, w18053, w18054, w18055, w18056, w18057, w18058, w18059, w18060, w18061, w18062, w18063, w18064, w18065, w18066, w18067, w18068, w18069, w18070, w18071, w18072, w18073, w18074, w18075, w18076, w18077, w18078, w18079, w18080, w18081, w18082, w18083, w18084, w18085, w18086, w18087, w18088, w18089, w18090, w18091, w18092, w18093, w18094, w18095, w18096, w18097, w18098, w18099, w18100, w18101, w18102, w18103, w18104, w18105, w18106, w18107, w18108, w18109, w18110, w18111, w18112, w18113, w18114, w18115, w18116, w18117, w18118, w18119, w18120, w18121, w18122, w18123, w18124, w18125, w18126, w18127, w18128, w18129, w18130, w18131, w18132, w18133, w18134, w18135, w18136, w18137, w18138, w18139, w18140, w18141, w18142, w18143, w18144, w18145, w18146, w18147, w18148, w18149, w18150, w18151, w18152, w18153, w18154, w18155, w18156, w18157, w18158, w18159, w18160, w18161, w18162, w18163, w18164, w18165, w18166, w18167, w18168, w18169, w18170, w18171, w18172, w18173, w18174, w18175, w18176, w18177, w18178, w18179, w18180, w18181, w18182, w18183, w18184, w18185, w18186, w18187, w18188, w18189, w18190, w18191, w18192, w18193, w18194, w18195, w18196, w18197, w18198, w18199, w18200, w18201, w18202, w18203, w18204, w18205, w18206, w18207, w18208, w18209, w18210, w18211, w18212, w18213, w18214, w18215, w18216, w18217, w18218, w18219, w18220, w18221, w18222, w18223, w18224, w18225, w18226, w18227, w18228, w18229, w18230, w18231, w18232, w18233, w18234, w18235, w18236, w18237, w18238, w18239, w18240, w18241, w18242, w18243, w18244, w18245, w18246, w18247, w18248, w18249, w18250, w18251, w18252, w18253, w18254, w18255, w18256, w18257, w18258, w18259, w18260, w18261, w18262, w18263, w18264, w18265, w18266, w18267, w18268, w18269, w18270, w18271, w18272, w18273, w18274, w18275, w18276, w18277, w18278, w18279, w18280, w18281, w18282, w18283, w18284, w18285, w18286, w18287, w18288, w18289, w18290, w18291, w18292, w18293, w18294, w18295, w18296, w18297, w18298, w18299, w18300, w18301, w18302, w18303, w18304, w18305, w18306, w18307, w18308, w18309, w18310, w18311, w18312, w18313, w18314, w18315, w18316, w18317, w18318, w18319, w18320, w18321, w18322, w18323, w18324, w18325, w18326, w18327, w18328, w18329, w18330, w18331, w18332, w18333, w18334, w18335, w18336, w18337, w18338, w18339, w18340, w18341, w18342, w18343, w18344, w18345, w18346, w18347, w18348, w18349, w18350, w18351, w18352, w18353, w18354, w18355, w18356, w18357, w18358, w18359, w18360, w18361, w18362, w18363, w18364, w18365, w18366, w18367, w18368, w18369, w18370, w18371, w18372, w18373, w18374, w18375, w18376, w18377, w18378, w18379, w18380, w18381, w18382, w18383, w18384, w18385, w18386, w18387, w18388, w18389, w18390, w18391, w18392, w18393, w18394, w18395, w18396, w18397, w18398, w18399, w18400, w18401, w18402, w18403, w18404, w18405, w18406, w18407, w18408, w18409, w18410, w18411, w18412, w18413, w18414, w18415, w18416, w18417, w18418, w18419, w18420, w18421, w18422, w18423, w18424, w18425, w18426, w18427, w18428, w18429, w18430, w18431, w18432, w18433, w18434, w18435, w18436, w18437, w18438, w18439, w18440, w18441, w18442, w18443, w18444, w18445, w18446, w18447, w18448, w18449, w18450, w18451, w18452, w18453, w18454, w18455, w18456, w18457, w18458, w18459, w18460, w18461, w18462, w18463, w18464, w18465, w18466, w18467, w18468, w18469, w18470, w18471, w18472, w18473, w18474, w18475, w18476, w18477, w18478, w18479, w18480, w18481, w18482, w18483, w18484, w18485, w18486, w18487, w18488, w18489, w18490, w18491, w18492, w18493, w18494, w18495, w18496, w18497, w18498, w18499, w18500, w18501, w18502, w18503, w18504, w18505, w18506, w18507, w18508, w18509, w18510, w18511, w18512, w18513, w18514, w18515, w18516, w18517, w18518, w18519, w18520, w18521, w18522, w18523, w18524, w18525, w18526, w18527, w18528, w18529, w18530, w18531, w18532, w18533, w18534, w18535, w18536, w18537, w18538, w18539, w18540, w18541, w18542, w18543, w18544, w18545, w18546, w18547, w18548, w18549, w18550, w18551, w18552, w18553, w18554, w18555, w18556, w18557, w18558, w18559, w18560, w18561, w18562, w18563, w18564, w18565, w18566, w18567, w18568, w18569, w18570, w18571, w18572, w18573, w18574, w18575, w18576, w18577, w18578, w18579, w18580, w18581, w18582, w18583, w18584, w18585, w18586, w18587, w18588, w18589, w18590, w18591, w18592, w18593, w18594, w18595, w18596, w18597, w18598, w18599, w18600, w18601, w18602, w18603, w18604, w18605, w18606, w18607, w18608, w18609, w18610, w18611, w18612, w18613, w18614, w18615, w18616, w18617, w18618, w18619, w18620, w18621, w18622, w18623, w18624, w18625, w18626, w18627, w18628, w18629, w18630, w18631, w18632, w18633, w18634, w18635, w18636, w18637, w18638, w18639, w18640, w18641, w18642, w18643, w18644, w18645, w18646, w18647, w18648, w18649, w18650, w18651, w18652, w18653, w18654, w18655, w18656, w18657, w18658, w18659, w18660, w18661, w18662, w18663, w18664, w18665, w18666, w18667, w18668, w18669, w18670, w18671, w18672, w18673, w18674, w18675, w18676, w18677, w18678, w18679, w18680, w18681, w18682, w18683, w18684, w18685, w18686, w18687, w18688, w18689, w18690, w18691, w18692, w18693, w18694, w18695, w18696, w18697, w18698, w18699, w18700, w18701, w18702, w18703, w18704, w18705, w18706, w18707, w18708, w18709, w18710, w18711, w18712, w18713, w18714, w18715, w18716, w18717, w18718, w18719, w18720, w18721, w18722, w18723, w18724, w18725, w18726, w18727, w18728, w18729, w18730, w18731, w18732, w18733, w18734, w18735, w18736, w18737, w18738, w18739, w18740, w18741, w18742, w18743, w18744, w18745, w18746, w18747, w18748, w18749, w18750, w18751, w18752, w18753, w18754, w18755, w18756, w18757, w18758, w18759, w18760, w18761, w18762, w18763, w18764, w18765, w18766, w18767, w18768, w18769, w18770, w18771, w18772, w18773, w18774, w18775, w18776, w18777, w18778, w18779, w18780, w18781, w18782, w18783, w18784, w18785, w18786, w18787, w18788, w18789, w18790, w18791, w18792, w18793, w18794, w18795, w18796, w18797, w18798, w18799, w18800, w18801, w18802, w18803, w18804, w18805, w18806, w18807, w18808, w18809, w18810, w18811, w18812, w18813, w18814, w18815, w18816, w18817, w18818, w18819, w18820, w18821, w18822, w18823, w18824, w18825, w18826, w18827, w18828, w18829, w18830, w18831, w18832, w18833, w18834, w18835, w18836, w18837, w18838, w18839, w18840, w18841, w18842, w18843, w18844, w18845, w18846, w18847, w18848, w18849, w18850, w18851, w18852, w18853, w18854, w18855, w18856, w18857, w18858, w18859, w18860, w18861, w18862, w18863, w18864, w18865, w18866, w18867, w18868, w18869, w18870, w18871, w18872, w18873, w18874, w18875, w18876, w18877, w18878, w18879, w18880, w18881, w18882, w18883, w18884, w18885, w18886, w18887, w18888, w18889, w18890, w18891, w18892, w18893, w18894, w18895, w18896, w18897, w18898, w18899, w18900, w18901, w18902, w18903, w18904, w18905, w18906, w18907, w18908, w18909, w18910, w18911, w18912, w18913, w18914, w18915, w18916, w18917, w18918, w18919, w18920, w18921, w18922, w18923, w18924, w18925, w18926, w18927, w18928, w18929, w18930, w18931, w18932, w18933, w18934, w18935, w18936, w18937, w18938, w18939, w18940, w18941, w18942, w18943, w18944, w18945, w18946, w18947, w18948, w18949, w18950, w18951, w18952, w18953, w18954, w18955, w18956, w18957, w18958, w18959, w18960, w18961, w18962, w18963, w18964, w18965, w18966, w18967, w18968, w18969, w18970, w18971, w18972, w18973, w18974, w18975, w18976, w18977, w18978, w18979, w18980, w18981, w18982, w18983, w18984, w18985, w18986, w18987, w18988, w18989, w18990, w18991, w18992, w18993, w18994, w18995, w18996, w18997, w18998, w18999, w19000, w19001, w19002, w19003, w19004, w19005, w19006, w19007, w19008, w19009, w19010, w19011, w19012, w19013, w19014, w19015, w19016, w19017, w19018, w19019, w19020, w19021, w19022, w19023, w19024, w19025, w19026, w19027, w19028, w19029, w19030, w19031, w19032, w19033, w19034, w19035, w19036, w19037, w19038, w19039, w19040, w19041, w19042, w19043, w19044, w19045, w19046, w19047, w19048, w19049, w19050, w19051, w19052, w19053, w19054, w19055, w19056, w19057, w19058, w19059, w19060, w19061, w19062, w19063, w19064, w19065, w19066, w19067, w19068, w19069, w19070, w19071, w19072, w19073, w19074, w19075, w19076, w19077, w19078, w19079, w19080, w19081, w19082, w19083, w19084, w19085, w19086, w19087, w19088, w19089, w19090, w19091, w19092, w19093, w19094, w19095, w19096, w19097, w19098, w19099, w19100, w19101, w19102, w19103, w19104, w19105, w19106, w19107, w19108, w19109, w19110, w19111, w19112, w19113, w19114, w19115, w19116, w19117, w19118, w19119, w19120, w19121, w19122, w19123, w19124, w19125, w19126, w19127, w19128, w19129, w19130, w19131, w19132, w19133, w19134, w19135, w19136, w19137, w19138, w19139, w19140, w19141, w19142, w19143, w19144, w19145, w19146, w19147, w19148, w19149, w19150, w19151, w19152, w19153, w19154, w19155, w19156, w19157, w19158, w19159, w19160, w19161, w19162, w19163, w19164, w19165, w19166, w19167, w19168, w19169, w19170, w19171, w19172, w19173, w19174, w19175, w19176, w19177, w19178, w19179, w19180, w19181, w19182, w19183, w19184, w19185, w19186, w19187, w19188, w19189, w19190, w19191, w19192, w19193, w19194, w19195, w19196, w19197, w19198, w19199, w19200, w19201, w19202, w19203, w19204, w19205, w19206, w19207, w19208, w19209, w19210, w19211, w19212, w19213, w19214, w19215, w19216, w19217, w19218, w19219, w19220, w19221, w19222, w19223, w19224, w19225, w19226, w19227, w19228, w19229, w19230, w19231, w19232, w19233, w19234, w19235, w19236, w19237, w19238, w19239, w19240, w19241, w19242, w19243, w19244, w19245, w19246, w19247, w19248, w19249, w19250, w19251, w19252, w19253, w19254, w19255, w19256, w19257, w19258, w19259, w19260, w19261, w19262, w19263, w19264, w19265, w19266, w19267, w19268, w19269, w19270, w19271, w19272, w19273, w19274, w19275, w19276, w19277, w19278, w19279, w19280, w19281, w19282, w19283, w19284, w19285, w19286, w19287, w19288, w19289, w19290, w19291, w19292, w19293, w19294, w19295, w19296, w19297, w19298, w19299, w19300, w19301, w19302, w19303, w19304, w19305, w19306, w19307, w19308, w19309, w19310, w19311, w19312, w19313, w19314, w19315, w19316, w19317, w19318, w19319, w19320, w19321, w19322, w19323, w19324, w19325, w19326, w19327, w19328, w19329, w19330, w19331, w19332, w19333, w19334, w19335, w19336, w19337, w19338, w19339, w19340, w19341, w19342, w19343, w19344, w19345, w19346, w19347, w19348, w19349, w19350, w19351, w19352, w19353, w19354, w19355, w19356, w19357, w19358, w19359, w19360, w19361, w19362, w19363, w19364, w19365, w19366, w19367, w19368, w19369, w19370, w19371, w19372, w19373, w19374, w19375, w19376, w19377, w19378, w19379, w19380, w19381, w19382, w19383, w19384, w19385, w19386, w19387, w19388, w19389, w19390, w19391, w19392, w19393, w19394, w19395, w19396, w19397, w19398, w19399, w19400, w19401, w19402, w19403, w19404, w19405, w19406, w19407, w19408, w19409, w19410, w19411, w19412, w19413, w19414, w19415, w19416, w19417, w19418, w19419, w19420, w19421, w19422, w19423, w19424, w19425, w19426, w19427, w19428, w19429, w19430, w19431, w19432, w19433, w19434, w19435, w19436, w19437, w19438, w19439, w19440, w19441, w19442, w19443, w19444, w19445, w19446, w19447, w19448, w19449, w19450, w19451, w19452, w19453, w19454, w19455, w19456, w19457, w19458, w19459, w19460, w19461, w19462, w19463, w19464, w19465, w19466, w19467, w19468, w19469, w19470, w19471, w19472, w19473, w19474, w19475, w19476, w19477, w19478, w19479, w19480, w19481, w19482, w19483, w19484, w19485, w19486, w19487, w19488, w19489, w19490, w19491, w19492, w19493, w19494, w19495, w19496, w19497, w19498, w19499, w19500, w19501, w19502, w19503, w19504, w19505, w19506, w19507, w19508, w19509, w19510, w19511, w19512, w19513, w19514, w19515, w19516, w19517, w19518, w19519, w19520, w19521, w19522, w19523, w19524, w19525, w19526, w19527, w19528, w19529, w19530, w19531, w19532, w19533, w19534, w19535, w19536, w19537, w19538, w19539, w19540, w19541, w19542, w19543, w19544, w19545, w19546, w19547, w19548, w19549, w19550, w19551, w19552, w19553, w19554, w19555, w19556, w19557, w19558, w19559, w19560, w19561, w19562, w19563, w19564, w19565, w19566, w19567, w19568, w19569, w19570, w19571, w19572, w19573, w19574, w19575, w19576, w19577, w19578, w19579, w19580, w19581, w19582, w19583, w19584, w19585, w19586, w19587, w19588, w19589, w19590, w19591, w19592, w19593, w19594, w19595, w19596, w19597, w19598, w19599, w19600, w19601, w19602, w19603, w19604, w19605, w19606, w19607, w19608, w19609, w19610, w19611, w19612, w19613, w19614, w19615, w19616, w19617, w19618, w19619, w19620, w19621, w19622, w19623, w19624, w19625, w19626, w19627, w19628, w19629, w19630, w19631, w19632, w19633, w19634, w19635, w19636, w19637, w19638, w19639, w19640, w19641, w19642, w19643, w19644, w19645, w19646, w19647, w19648, w19649, w19650, w19651, w19652, w19653, w19654, w19655, w19656, w19657, w19658, w19659, w19660, w19661, w19662, w19663, w19664, w19665, w19666, w19667, w19668, w19669, w19670, w19671, w19672, w19673, w19674, w19675, w19676, w19677, w19678, w19679, w19680, w19681, w19682, w19683, w19684, w19685, w19686, w19687, w19688, w19689, w19690, w19691, w19692, w19693, w19694, w19695, w19696, w19697, w19698, w19699, w19700, w19701, w19702, w19703, w19704, w19705, w19706, w19707, w19708, w19709, w19710, w19711, w19712, w19713, w19714, w19715, w19716, w19717, w19718, w19719, w19720, w19721, w19722, w19723, w19724, w19725, w19726, w19727, w19728, w19729, w19730, w19731, w19732, w19733, w19734, w19735, w19736, w19737, w19738, w19739, w19740, w19741, w19742, w19743, w19744, w19745, w19746, w19747, w19748, w19749, w19750, w19751, w19752, w19753, w19754, w19755, w19756, w19757, w19758, w19759, w19760, w19761, w19762, w19763, w19764, w19765, w19766, w19767, w19768, w19769, w19770, w19771, w19772, w19773, w19774, w19775, w19776, w19777, w19778, w19779, w19780, w19781, w19782, w19783, w19784, w19785, w19786, w19787, w19788, w19789, w19790, w19791, w19792, w19793, w19794, w19795, w19796, w19797, w19798, w19799, w19800, w19801, w19802, w19803, w19804, w19805, w19806, w19807, w19808, w19809, w19810, w19811, w19812, w19813, w19814, w19815, w19816, w19817, w19818, w19819, w19820, w19821, w19822, w19823, w19824, w19825, w19826, w19827, w19828, w19829, w19830, w19831, w19832, w19833, w19834, w19835, w19836, w19837, w19838, w19839, w19840, w19841, w19842, w19843, w19844, w19845, w19846, w19847, w19848, w19849, w19850, w19851, w19852, w19853, w19854, w19855, w19856, w19857, w19858, w19859, w19860, w19861, w19862, w19863, w19864, w19865, w19866, w19867, w19868, w19869, w19870, w19871, w19872, w19873, w19874, w19875, w19876, w19877, w19878, w19879, w19880, w19881, w19882, w19883, w19884, w19885, w19886, w19887, w19888, w19889, w19890, w19891, w19892, w19893, w19894, w19895, w19896, w19897, w19898, w19899, w19900, w19901, w19902, w19903, w19904, w19905, w19906, w19907, w19908, w19909, w19910, w19911, w19912, w19913, w19914, w19915, w19916, w19917, w19918, w19919, w19920, w19921, w19922, w19923, w19924, w19925, w19926, w19927, w19928, w19929, w19930, w19931, w19932, w19933, w19934, w19935, w19936, w19937, w19938, w19939, w19940, w19941, w19942, w19943, w19944, w19945, w19946, w19947, w19948, w19949, w19950, w19951, w19952, w19953, w19954, w19955, w19956, w19957, w19958, w19959, w19960, w19961, w19962, w19963, w19964, w19965, w19966, w19967, w19968, w19969, w19970, w19971, w19972, w19973, w19974, w19975, w19976, w19977, w19978, w19979, w19980, w19981, w19982, w19983, w19984, w19985, w19986, w19987, w19988, w19989, w19990, w19991, w19992, w19993, w19994, w19995, w19996, w19997, w19998, w19999, w20000, w20001, w20002, w20003, w20004, w20005, w20006, w20007, w20008, w20009, w20010, w20011, w20012, w20013, w20014, w20015, w20016, w20017, w20018, w20019, w20020, w20021, w20022, w20023, w20024, w20025, w20026, w20027, w20028, w20029, w20030, w20031, w20032, w20033, w20034, w20035, w20036, w20037, w20038, w20039, w20040, w20041, w20042, w20043, w20044, w20045, w20046, w20047, w20048, w20049, w20050, w20051, w20052, w20053, w20054, w20055, w20056, w20057, w20058, w20059, w20060, w20061, w20062, w20063, w20064, w20065, w20066, w20067, w20068, w20069, w20070, w20071, w20072, w20073, w20074, w20075, w20076, w20077, w20078, w20079, w20080, w20081, w20082, w20083, w20084, w20085, w20086, w20087, w20088, w20089, w20090, w20091, w20092, w20093, w20094, w20095, w20096, w20097, w20098, w20099, w20100, w20101, w20102, w20103, w20104, w20105, w20106, w20107, w20108, w20109, w20110, w20111, w20112, w20113, w20114, w20115, w20116, w20117, w20118, w20119, w20120, w20121, w20122, w20123, w20124, w20125, w20126, w20127, w20128, w20129, w20130, w20131, w20132, w20133, w20134, w20135, w20136, w20137, w20138, w20139, w20140, w20141, w20142, w20143, w20144, w20145, w20146, w20147, w20148, w20149, w20150, w20151, w20152, w20153, w20154, w20155, w20156, w20157, w20158, w20159, w20160, w20161, w20162, w20163, w20164, w20165, w20166, w20167, w20168, w20169, w20170, w20171, w20172, w20173, w20174, w20175, w20176, w20177, w20178, w20179, w20180, w20181, w20182, w20183, w20184, w20185, w20186, w20187, w20188, w20189, w20190, w20191, w20192, w20193, w20194, w20195, w20196, w20197, w20198, w20199, w20200, w20201, w20202, w20203, w20204, w20205, w20206, w20207, w20208, w20209, w20210, w20211, w20212, w20213, w20214, w20215, w20216, w20217, w20218, w20219, w20220, w20221, w20222, w20223, w20224, w20225, w20226, w20227, w20228, w20229, w20230, w20231, w20232, w20233, w20234, w20235, w20236, w20237, w20238, w20239, w20240, w20241, w20242, w20243, w20244, w20245, w20246, w20247, w20248, w20249, w20250, w20251, w20252, w20253, w20254, w20255, w20256, w20257, w20258, w20259, w20260, w20261, w20262, w20263, w20264, w20265, w20266, w20267, w20268, w20269, w20270, w20271, w20272, w20273, w20274, w20275, w20276, w20277, w20278, w20279, w20280, w20281, w20282, w20283, w20284, w20285, w20286, w20287, w20288, w20289, w20290, w20291, w20292, w20293, w20294, w20295, w20296, w20297, w20298, w20299, w20300, w20301, w20302, w20303, w20304, w20305, w20306, w20307, w20308, w20309, w20310, w20311, w20312, w20313, w20314, w20315, w20316, w20317, w20318, w20319, w20320, w20321, w20322, w20323, w20324, w20325, w20326, w20327, w20328, w20329, w20330, w20331, w20332, w20333, w20334, w20335, w20336, w20337, w20338, w20339, w20340, w20341, w20342, w20343, w20344, w20345, w20346, w20347, w20348, w20349, w20350, w20351, w20352, w20353, w20354, w20355, w20356, w20357, w20358, w20359, w20360, w20361, w20362, w20363, w20364, w20365, w20366, w20367, w20368, w20369, w20370, w20371, w20372, w20373, w20374, w20375, w20376, w20377, w20378, w20379, w20380, w20381, w20382, w20383, w20384, w20385, w20386, w20387, w20388, w20389, w20390, w20391, w20392, w20393, w20394, w20395, w20396, w20397, w20398, w20399, w20400, w20401, w20402, w20403, w20404, w20405, w20406, w20407, w20408, w20409, w20410, w20411, w20412, w20413, w20414, w20415, w20416, w20417, w20418, w20419, w20420, w20421, w20422, w20423, w20424, w20425, w20426, w20427, w20428, w20429, w20430, w20431, w20432, w20433, w20434, w20435, w20436, w20437, w20438, w20439, w20440, w20441, w20442, w20443, w20444, w20445, w20446, w20447, w20448, w20449, w20450, w20451, w20452, w20453, w20454, w20455, w20456, w20457, w20458, w20459, w20460, w20461, w20462, w20463, w20464, w20465, w20466, w20467, w20468, w20469, w20470, w20471, w20472, w20473, w20474, w20475, w20476, w20477, w20478, w20479, w20480, w20481, w20482, w20483, w20484, w20485, w20486, w20487, w20488, w20489, w20490, w20491, w20492, w20493, w20494, w20495, w20496, w20497, w20498, w20499, w20500, w20501, w20502, w20503, w20504, w20505, w20506, w20507, w20508, w20509, w20510, w20511, w20512, w20513, w20514, w20515, w20516, w20517, w20518, w20519, w20520, w20521, w20522, w20523, w20524, w20525, w20526, w20527, w20528, w20529, w20530, w20531, w20532, w20533, w20534, w20535, w20536, w20537, w20538, w20539, w20540, w20541, w20542, w20543, w20544, w20545, w20546, w20547, w20548, w20549, w20550, w20551, w20552, w20553, w20554, w20555, w20556, w20557, w20558, w20559, w20560, w20561, w20562, w20563, w20564, w20565, w20566, w20567, w20568, w20569, w20570, w20571, w20572, w20573, w20574, w20575, w20576, w20577, w20578, w20579, w20580, w20581, w20582, w20583, w20584, w20585, w20586, w20587, w20588, w20589, w20590, w20591, w20592, w20593, w20594, w20595, w20596, w20597, w20598, w20599, w20600, w20601, w20602, w20603, w20604, w20605, w20606, w20607, w20608, w20609, w20610, w20611, w20612, w20613, w20614, w20615, w20616, w20617, w20618, w20619, w20620, w20621, w20622, w20623, w20624, w20625, w20626, w20627, w20628, w20629, w20630, w20631, w20632, w20633, w20634, w20635, w20636, w20637, w20638, w20639, w20640, w20641, w20642, w20643, w20644, w20645, w20646, w20647, w20648, w20649, w20650, w20651, w20652, w20653, w20654, w20655, w20656, w20657, w20658, w20659, w20660, w20661, w20662, w20663, w20664, w20665, w20666, w20667, w20668, w20669, w20670, w20671, w20672, w20673, w20674, w20675, w20676, w20677, w20678, w20679, w20680, w20681, w20682, w20683, w20684, w20685, w20686, w20687, w20688, w20689, w20690, w20691, w20692, w20693, w20694, w20695, w20696, w20697, w20698, w20699, w20700, w20701, w20702, w20703, w20704, w20705, w20706, w20707, w20708, w20709, w20710, w20711, w20712, w20713, w20714, w20715, w20716, w20717, w20718, w20719, w20720, w20721, w20722, w20723, w20724, w20725, w20726, w20727, w20728, w20729, w20730, w20731, w20732, w20733, w20734, w20735, w20736, w20737, w20738, w20739, w20740, w20741, w20742, w20743, w20744, w20745, w20746, w20747, w20748, w20749, w20750, w20751, w20752, w20753, w20754, w20755, w20756, w20757, w20758, w20759, w20760, w20761, w20762, w20763, w20764, w20765, w20766, w20767, w20768, w20769, w20770, w20771, w20772, w20773, w20774, w20775, w20776, w20777, w20778, w20779, w20780, w20781, w20782, w20783, w20784, w20785, w20786, w20787, w20788, w20789, w20790, w20791, w20792, w20793, w20794, w20795, w20796, w20797, w20798, w20799, w20800, w20801, w20802, w20803, w20804, w20805, w20806, w20807, w20808, w20809, w20810, w20811, w20812, w20813, w20814, w20815, w20816, w20817, w20818, w20819, w20820, w20821, w20822, w20823, w20824, w20825, w20826, w20827, w20828, w20829, w20830, w20831, w20832, w20833, w20834, w20835, w20836, w20837, w20838, w20839, w20840, w20841, w20842, w20843, w20844, w20845, w20846, w20847, w20848, w20849, w20850, w20851, w20852, w20853, w20854, w20855, w20856, w20857, w20858, w20859, w20860, w20861, w20862, w20863, w20864, w20865, w20866, w20867, w20868, w20869, w20870, w20871, w20872, w20873, w20874, w20875, w20876, w20877, w20878, w20879, w20880, w20881, w20882, w20883, w20884, w20885, w20886, w20887, w20888, w20889, w20890, w20891, w20892, w20893, w20894, w20895, w20896, w20897, w20898, w20899, w20900, w20901, w20902, w20903, w20904, w20905, w20906, w20907, w20908, w20909, w20910, w20911, w20912, w20913, w20914, w20915, w20916, w20917, w20918, w20919, w20920, w20921, w20922, w20923, w20924, w20925, w20926, w20927, w20928, w20929, w20930, w20931, w20932, w20933, w20934, w20935, w20936, w20937, w20938, w20939, w20940, w20941, w20942, w20943, w20944, w20945, w20946;
assign w0 = pi014 & pi107;
assign w1 = ~pi082 & w0;
assign w2 = pi082 & ~pi108;
assign w3 = pi014 & ~pi072;
assign w4 = w2 & w3;
assign w5 = ~w1 & ~w4;
assign w6 = ~pi083 & ~w5;
assign w7 = ~pi072 & pi082;
assign w8 = ~pi014 & pi083;
assign w9 = pi107 & w8;
assign w10 = w7 & w9;
assign w11 = pi072 & pi108;
assign w12 = pi014 & ~pi082;
assign w13 = w11 & w12;
assign w14 = pi082 & pi108;
assign w15 = ~pi014 & ~pi072;
assign w16 = w14 & w15;
assign w17 = pi107 & w16;
assign w18 = ~w10 & ~w17;
assign w19 = ~w6 & w18;
assign w20 = ~pi072 & ~pi082;
assign w21 = pi107 & w20;
assign w22 = w20 & w17893;
assign w23 = ~pi014 & pi072;
assign w24 = w14 & w23;
assign w25 = pi072 & ~pi108;
assign w26 = ~pi014 & ~pi107;
assign w27 = w25 & w26;
assign w28 = ~w24 & ~w27;
assign w29 = pi072 & w2;
assign w30 = w0 & w29;
assign w31 = ~w22 & w28;
assign w32 = (~pi083 & ~w31) | (~pi083 & w17894) | (~w31 & w17894);
assign w33 = ~pi082 & ~pi108;
assign w34 = pi108 & w0;
assign w35 = ~w33 & ~w34;
assign w36 = ~pi072 & pi083;
assign w37 = (w36 & w34) | (w36 & w17895) | (w34 & w17895);
assign w38 = ~pi083 & pi108;
assign w39 = ~pi107 & w38;
assign w40 = pi014 & ~pi107;
assign w41 = pi072 & w40;
assign w42 = w40 & w11;
assign w43 = ~w39 & ~w42;
assign w44 = ~w37 & w43;
assign w45 = ~pi040 & ~w44;
assign w46 = pi014 & pi083;
assign w47 = pi072 & pi107;
assign w48 = w14 & w47;
assign w49 = w33 & w47;
assign w50 = ~pi107 & ~pi108;
assign w51 = w20 & w50;
assign w52 = ~w48 & ~w49;
assign w53 = (w46 & ~w52) | (w46 & w17896) | (~w52 & w17896);
assign w54 = ~w32 & ~w45;
assign w55 = ~w53 & w54;
assign w56 = pi072 & pi082;
assign w57 = pi107 & w56;
assign w58 = pi107 & w2;
assign w59 = ~w21 & ~w57;
assign w60 = ~pi107 & pi108;
assign w61 = ~pi072 & w60;
assign w62 = ~w58 & ~w61;
assign w63 = w8 & ~w62;
assign w64 = ~pi083 & w2;
assign w65 = w40 & w71;
assign w66 = ~w3 & w64;
assign w67 = ~w65 & ~w66;
assign w68 = ~w63 & w67;
assign w69 = w2 & w47;
assign w70 = ~pi014 & pi107;
assign w71 = pi072 & ~pi082;
assign w72 = w70 & w71;
assign w73 = w14 & w26;
assign w74 = ~w69 & ~w72;
assign w75 = (pi083 & ~w74) | (pi083 & w17899) | (~w74 & w17899);
assign w76 = (w70 & w64) | (w70 & w17900) | (w64 & w17900);
assign w77 = pi014 & w7;
assign w78 = pi083 & ~pi107;
assign w79 = w77 & w78;
assign w80 = ~pi072 & pi107;
assign w81 = w14 & w80;
assign w82 = pi014 & w81;
assign w83 = ~pi082 & pi108;
assign w84 = ~pi014 & ~pi083;
assign w85 = ~pi072 & w84;
assign w86 = w83 & w85;
assign w87 = ~w82 & ~w86;
assign w88 = pi040 & pi083;
assign w89 = pi082 & ~pi107;
assign w90 = ~w21 & ~w89;
assign w91 = pi014 & w2;
assign w92 = ~pi014 & w33;
assign w93 = ~w91 & ~w92;
assign w94 = w90 & w93;
assign w95 = w88 & ~w94;
assign w96 = pi040 & ~w87;
assign w97 = ~w95 & ~w96;
assign w98 = ~w76 & ~w79;
assign w99 = ~w75 & w98;
assign w100 = w97 & w99;
assign w101 = (pi078 & ~w100) | (pi078 & w17901) | (~w100 & w17901);
assign w102 = ~pi072 & pi108;
assign w103 = w89 & w102;
assign w104 = ~pi014 & w83;
assign w105 = w80 & w104;
assign w106 = w2 & w17902;
assign w107 = pi072 & w33;
assign w108 = w26 & w107;
assign w109 = ~w105 & ~w106;
assign w110 = ~w108 & w109;
assign w111 = ~w73 & ~w103;
assign w112 = pi083 & w111;
assign w113 = w110 & w112;
assign w114 = w7 & w50;
assign w115 = w56 & w60;
assign w116 = ~w114 & ~w115;
assign w117 = ~w60 & w71;
assign w118 = ~pi083 & ~w117;
assign w119 = w116 & w118;
assign w120 = pi040 & ~w84;
assign w121 = ~w119 & w120;
assign w122 = ~w113 & w121;
assign w123 = ~pi040 & pi083;
assign w124 = w56 & w70;
assign w125 = w3 & w33;
assign w126 = ~w82 & w17903;
assign w127 = w123 & ~w126;
assign w128 = w11 & w70;
assign w129 = w3 & w39;
assign w130 = ~w128 & ~w129;
assign w131 = ~pi083 & ~w28;
assign w132 = w130 & ~w131;
assign w133 = w26 & w56;
assign w134 = ~pi108 & w133;
assign w135 = ~pi072 & w33;
assign w136 = w0 & w135;
assign w137 = ~w134 & ~w136;
assign w138 = ~pi083 & ~w137;
assign w139 = ~pi040 & ~w132;
assign w140 = ~w138 & ~w139;
assign w141 = ~w122 & w140;
assign w142 = ~w127 & w141;
assign w143 = ~w101 & w142;
assign w144 = (~pi078 & ~w55) | (~pi078 & w17904) | (~w55 & w17904);
assign w145 = w142 & w20755;
assign w146 = ~pi082 & w23;
assign w147 = ~w71 & ~w80;
assign w148 = pi108 & ~w147;
assign w149 = (pi083 & w148) | (pi083 & w17905) | (w148 & w17905);
assign w150 = w47 & w83;
assign w151 = w3 & w14;
assign w152 = ~w150 & ~w151;
assign w153 = w33 & w17906;
assign w154 = w2 & w84;
assign w155 = ~w128 & ~w154;
assign w156 = w152 & ~w153;
assign w157 = w155 & w156;
assign w158 = ~pi083 & ~pi107;
assign w159 = pi072 & w50;
assign w160 = w3 & w83;
assign w161 = ~w159 & ~w160;
assign w162 = ~w4 & ~w16;
assign w163 = ~pi083 & ~w162;
assign w164 = pi072 & pi083;
assign w165 = w2 & w164;
assign w166 = w26 & w33;
assign w167 = ~w133 & ~w165;
assign w168 = ~w166 & w167;
assign w169 = ~w163 & w168;
assign w170 = (~pi040 & ~w169) | (~pi040 & w17907) | (~w169 & w17907);
assign w171 = w26 & w102;
assign w172 = ~pi082 & w128;
assign w173 = pi072 & w14;
assign w174 = w14 & w17902;
assign w175 = ~w172 & w17908;
assign w176 = ~pi083 & ~w175;
assign w177 = pi083 & pi107;
assign w178 = pi014 & w83;
assign w179 = ~w2 & ~w83;
assign w180 = ~pi072 & ~w179;
assign w181 = (w177 & w180) | (w177 & w17909) | (w180 & w17909);
assign w182 = w29 & w40;
assign w183 = ~w181 & ~w182;
assign w184 = ~w176 & w183;
assign w185 = ~w170 & w184;
assign w186 = (pi040 & ~w157) | (pi040 & w17910) | (~w157 & w17910);
assign w187 = ~pi072 & ~pi108;
assign w188 = ~pi107 & w187;
assign w189 = ~pi108 & w70;
assign w190 = w56 & w189;
assign w191 = w60 & w71;
assign w192 = ~pi083 & w191;
assign w193 = ~w160 & ~w192;
assign w194 = ~pi014 & w115;
assign w195 = w0 & w11;
assign w196 = pi082 & w195;
assign w197 = ~w194 & ~w196;
assign w198 = w193 & w197;
assign w199 = w8 & ~w20;
assign w200 = pi108 & w199;
assign w201 = ~w171 & ~w200;
assign w202 = pi014 & ~pi083;
assign w203 = w150 & w202;
assign w204 = pi072 & ~pi083;
assign w205 = w33 & ~w204;
assign w206 = pi107 & w205;
assign w207 = ~w203 & ~w206;
assign w208 = w201 & w207;
assign w209 = ~pi040 & ~w208;
assign w210 = pi082 & w70;
assign w211 = w11 & w210;
assign w212 = w2 & w0;
assign w213 = ~w211 & ~w212;
assign w214 = (~pi083 & w211) | (~pi083 & w17912) | (w211 & w17912);
assign w215 = w78 & w173;
assign w216 = ~pi014 & w114;
assign w217 = w46 & w188;
assign w218 = ~w216 & ~w217;
assign w219 = ~w215 & w218;
assign w220 = ~w214 & w219;
assign w221 = ~w209 & w220;
assign w222 = ~pi107 & w2;
assign w223 = ~w21 & ~w191;
assign w224 = (w84 & ~w223) | (w84 & w17914) | (~w223 & w17914);
assign w225 = pi082 & w41;
assign w226 = w152 & ~w225;
assign w227 = w20 & w60;
assign w228 = w202 & w227;
assign w229 = (~w228 & w226) | (~w228 & w17915) | (w226 & w17915);
assign w230 = (pi040 & ~w229) | (pi040 & w17916) | (~w229 & w17916);
assign w231 = w70 & w135;
assign w232 = ~w216 & ~w231;
assign w233 = w123 & ~w232;
assign w234 = ~pi040 & ~pi083;
assign w235 = pi014 & w14;
assign w236 = w14 & w40;
assign w237 = w80 & w91;
assign w238 = w160 & w177;
assign w239 = ~w237 & ~w238;
assign w240 = w234 & w236;
assign w241 = w77 & w17917;
assign w242 = w239 & w17918;
assign w243 = ~w233 & w242;
assign w244 = ~w230 & w243;
assign w245 = (~pi078 & ~w221) | (~pi078 & w17919) | (~w221 & w17919);
assign w246 = w244 & ~w245;
assign w247 = (pi078 & ~w185) | (pi078 & w17920) | (~w185 & w17920);
assign w248 = w246 & ~w247;
assign w249 = ~w145 & w248;
assign w250 = w145 & ~w248;
assign w251 = ~w249 & ~w250;
assign w252 = ~pi047 & ~pi093;
assign w253 = ~pi027 & w252;
assign w254 = pi047 & ~pi093;
assign w255 = pi027 & w254;
assign w256 = ~w253 & ~w255;
assign w257 = ~pi047 & ~pi111;
assign w258 = ~pi023 & ~pi027;
assign w259 = w257 & w258;
assign w260 = pi093 & w259;
assign w261 = ~pi023 & pi027;
assign w262 = pi111 & w261;
assign w263 = w261 & w282;
assign w264 = pi027 & ~pi047;
assign w265 = pi093 & ~pi111;
assign w266 = pi023 & w265;
assign w267 = w264 & w266;
assign w268 = ~w260 & ~w263;
assign w269 = ~w267 & w268;
assign w270 = pi023 & ~pi027;
assign w271 = ~pi093 & w270;
assign w272 = pi047 & ~pi111;
assign w273 = w271 & w272;
assign w274 = pi047 & pi093;
assign w275 = pi111 & w274;
assign w276 = w261 & w275;
assign w277 = ~pi027 & ~pi111;
assign w278 = w274 & w277;
assign w279 = ~w273 & ~w276;
assign w280 = (~pi123 & ~w279) | (~pi123 & w17921) | (~w279 & w17921);
assign w281 = ~pi023 & ~pi093;
assign w282 = ~pi047 & pi111;
assign w283 = w281 & w282;
assign w284 = ~pi027 & w283;
assign w285 = ~pi093 & pi111;
assign w286 = pi023 & pi027;
assign w287 = pi047 & w286;
assign w288 = w285 & w287;
assign w289 = ~w284 & ~w288;
assign w290 = ~w280 & w289;
assign w291 = (pi123 & ~w269) | (pi123 & w17922) | (~w269 & w17922);
assign w292 = w290 & ~w291;
assign w293 = ~pi023 & w254;
assign w294 = ~pi047 & pi093;
assign w295 = pi023 & ~pi111;
assign w296 = w294 & w295;
assign w297 = ~w293 & ~w296;
assign w298 = ~pi123 & ~w297;
assign w299 = ~pi111 & w252;
assign w300 = w270 & w299;
assign w301 = (pi048 & ~w299) | (pi048 & w17923) | (~w299 & w17923);
assign w302 = w252 & w261;
assign w303 = pi111 & w302;
assign w304 = ~pi023 & pi123;
assign w305 = w294 & w304;
assign w306 = ~w298 & w301;
assign w307 = ~w303 & ~w305;
assign w308 = w306 & w307;
assign w309 = w252 & w286;
assign w310 = (~pi048 & ~w309) | (~pi048 & w1118) | (~w309 & w1118);
assign w311 = pi023 & pi093;
assign w312 = w282 & w311;
assign w313 = pi123 & w312;
assign w314 = ~pi023 & pi093;
assign w315 = pi027 & pi047;
assign w316 = w314 & w315;
assign w317 = pi093 & pi111;
assign w318 = ~pi023 & ~pi123;
assign w319 = ~pi027 & ~w318;
assign w320 = w317 & ~w319;
assign w321 = ~w313 & ~w320;
assign w322 = w321 & w17924;
assign w323 = ~w308 & ~w322;
assign w324 = w264 & w265;
assign w325 = pi123 & ~w324;
assign w326 = pi047 & pi111;
assign w327 = w314 & w326;
assign w328 = ~w302 & ~w327;
assign w329 = w264 & w314;
assign w330 = w325 & w328;
assign w331 = ~w271 & ~w329;
assign w332 = w330 & w331;
assign w333 = ~pi093 & w259;
assign w334 = w265 & w315;
assign w335 = ~pi123 & ~w334;
assign w336 = w281 & w315;
assign w337 = ~w333 & w335;
assign w338 = ~w336 & w337;
assign w339 = ~w332 & ~w338;
assign w340 = w294 & ~w295;
assign w341 = ~w262 & w340;
assign w342 = ~pi123 & w341;
assign w343 = ~pi027 & pi123;
assign w344 = w266 & w343;
assign w345 = pi111 & w254;
assign w346 = w254 & w17925;
assign w347 = w254 & w286;
assign w348 = ~w344 & ~w346;
assign w349 = ~w342 & w348;
assign w350 = pi023 & w326;
assign w351 = ~w299 & ~w350;
assign w352 = pi123 & ~w351;
assign w353 = ~pi027 & ~pi123;
assign w354 = w254 & w353;
assign w355 = pi111 & w354;
assign w356 = ~w302 & ~w355;
assign w357 = ~w352 & w356;
assign w358 = ~pi048 & ~w357;
assign w359 = ~pi023 & w272;
assign w360 = ~w309 & ~w359;
assign w361 = pi123 & ~w360;
assign w362 = (pi027 & ~w252) | (pi027 & w17926) | (~w252 & w17926);
assign w363 = ~w360 & w17927;
assign w364 = w272 & w311;
assign w365 = ~pi027 & w364;
assign w366 = w364 & w353;
assign w367 = (~pi020 & ~w283) | (~pi020 & w17928) | (~w283 & w17928);
assign w368 = ~w366 & w367;
assign w369 = ~w363 & w368;
assign w370 = ~w358 & w369;
assign w371 = (pi048 & ~w349) | (pi048 & w17929) | (~w349 & w17929);
assign w372 = w370 & ~w371;
assign w373 = pi020 & ~w339;
assign w374 = ~w323 & w373;
assign w375 = ~w372 & ~w374;
assign w376 = ~pi027 & pi111;
assign w377 = ~pi023 & w274;
assign w378 = w376 & w377;
assign w379 = pi027 & ~pi111;
assign w380 = ~w252 & w379;
assign w381 = ~w333 & ~w378;
assign w382 = (~pi123 & ~w381) | (~pi123 & w17930) | (~w381 & w17930);
assign w383 = pi027 & pi123;
assign w384 = ~w345 & w383;
assign w385 = ~w345 & w17931;
assign w386 = pi123 & w270;
assign w387 = w254 & w386;
assign w388 = pi027 & w364;
assign w389 = ~pi111 & w294;
assign w390 = w261 & w389;
assign w391 = ~w387 & ~w388;
assign w392 = w391 & w17932;
assign w393 = ~w382 & w392;
assign w394 = pi027 & ~pi123;
assign w395 = ~pi023 & ~pi111;
assign w396 = w254 & w395;
assign w397 = w350 & w383;
assign w398 = w394 & w396;
assign w399 = ~w397 & ~w398;
assign w400 = (w399 & w393) | (w399 & w17933) | (w393 & w17933);
assign w401 = ~pi048 & ~w292;
assign w402 = ~w375 & w17934;
assign w403 = pi021 & ~pi098;
assign w404 = ~pi007 & w403;
assign w405 = ~pi021 & ~pi054;
assign w406 = pi007 & w405;
assign w407 = ~w404 & ~w406;
assign w408 = ~pi021 & ~pi098;
assign w409 = ~pi054 & w408;
assign w410 = (~pi114 & ~w408) | (~pi114 & w17935) | (~w408 & w17935);
assign w411 = pi007 & ~pi013;
assign w412 = w409 & w411;
assign w413 = ~pi007 & pi013;
assign w414 = ~pi021 & w413;
assign w415 = pi054 & ~pi098;
assign w416 = w414 & w415;
assign w417 = ~pi021 & pi098;
assign w418 = ~pi007 & pi114;
assign w419 = w417 & w418;
assign w420 = ~w412 & ~w416;
assign w421 = pi001 & ~w419;
assign w422 = w420 & w421;
assign w423 = ~w407 & w410;
assign w424 = w422 & ~w423;
assign w425 = pi007 & pi054;
assign w426 = w417 & w425;
assign w427 = pi114 & w426;
assign w428 = pi021 & pi098;
assign w429 = w413 & w428;
assign w430 = ~pi001 & ~w429;
assign w431 = ~w427 & w430;
assign w432 = pi007 & pi013;
assign w433 = w408 & w432;
assign w434 = ~pi114 & w433;
assign w435 = pi054 & pi098;
assign w436 = ~pi007 & ~pi114;
assign w437 = ~pi013 & ~w436;
assign w438 = w435 & ~w437;
assign w439 = ~w434 & ~w438;
assign w440 = w431 & w439;
assign w441 = ~w424 & ~w440;
assign w442 = ~pi007 & ~pi013;
assign w443 = w405 & w442;
assign w444 = ~pi098 & w443;
assign w445 = ~pi007 & ~pi098;
assign w446 = pi013 & pi021;
assign w447 = w445 & w446;
assign w448 = pi013 & ~pi054;
assign w449 = w428 & w448;
assign w450 = ~pi114 & ~w449;
assign w451 = ~pi098 & w411;
assign w452 = ~w414 & ~w451;
assign w453 = ~pi007 & pi021;
assign w454 = w435 & w453;
assign w455 = pi013 & ~pi021;
assign w456 = ~pi054 & pi098;
assign w457 = w455 & w456;
assign w458 = ~w454 & ~w457;
assign w459 = w452 & w458;
assign w460 = pi114 & w459;
assign w461 = ~w444 & w450;
assign w462 = ~w447 & w461;
assign w463 = ~w460 & ~w462;
assign w464 = pi029 & ~w463;
assign w465 = ~w441 & w464;
assign w466 = pi007 & ~pi054;
assign w467 = w428 & w466;
assign w468 = ~pi013 & w467;
assign w469 = pi054 & w413;
assign w470 = w417 & ~w466;
assign w471 = ~w469 & w470;
assign w472 = pi001 & w471;
assign w473 = (~pi114 & w472) | (~pi114 & w17936) | (w472 & w17936);
assign w474 = pi114 & w409;
assign w475 = pi021 & pi054;
assign w476 = pi007 & pi114;
assign w477 = w475 & w476;
assign w478 = pi054 & w403;
assign w479 = ~pi013 & ~pi114;
assign w480 = w413 & w408;
assign w481 = w478 & w479;
assign w482 = ~w480 & ~w481;
assign w483 = ~pi001 & ~w477;
assign w484 = ~w474 & w483;
assign w485 = w482 & w484;
assign w486 = pi114 & w411;
assign w487 = w403 & w17937;
assign w488 = w403 & w432;
assign w489 = pi001 & ~w488;
assign w490 = ~w487 & w489;
assign w491 = w456 & w486;
assign w492 = w490 & ~w491;
assign w493 = ~pi054 & w453;
assign w494 = ~w433 & ~w493;
assign w495 = pi114 & ~w494;
assign w496 = (pi013 & ~w408) | (pi013 & w17938) | (~w408 & w17938);
assign w497 = ~w494 & w17939;
assign w498 = w408 & w442;
assign w499 = pi054 & w498;
assign w500 = (~pi029 & ~w498) | (~pi029 & w17940) | (~w498 & w17940);
assign w501 = ~w497 & w500;
assign w502 = ~w485 & ~w492;
assign w503 = ~w502 & w17941;
assign w504 = ~w465 & ~w503;
assign w505 = w413 & w971;
assign w506 = w415 & w446;
assign w507 = ~pi054 & w417;
assign w508 = ~w411 & ~w413;
assign w509 = pi054 & w408;
assign w510 = w408 & w17942;
assign w511 = w507 & w508;
assign w512 = ~w510 & ~w511;
assign w513 = ~w505 & ~w506;
assign w514 = (pi114 & ~w512) | (pi114 & w17943) | (~w512 & w17943);
assign w515 = ~pi054 & ~pi098;
assign w516 = w453 & w515;
assign w517 = ~pi114 & w516;
assign w518 = (pi013 & w517) | (pi013 & w17944) | (w517 & w17944);
assign w519 = pi021 & ~pi054;
assign w520 = ~w445 & ~w446;
assign w521 = w428 & w469;
assign w522 = w519 & w520;
assign w523 = ~w521 & ~w522;
assign w524 = pi013 & w403;
assign w525 = w425 & w524;
assign w526 = ~w499 & ~w525;
assign w527 = ~pi001 & w526;
assign w528 = ~pi114 & ~w523;
assign w529 = w527 & ~w528;
assign w530 = w529 & w17945;
assign w531 = w442 & w475;
assign w532 = pi098 & w531;
assign w533 = ~w408 & w448;
assign w534 = ~w444 & ~w532;
assign w535 = (~pi114 & ~w534) | (~pi114 & w17946) | (~w534 & w17946);
assign w536 = pi013 & pi114;
assign w537 = w509 & w536;
assign w538 = ~pi013 & w403;
assign w539 = w446 & w466;
assign w540 = pi098 & w539;
assign w541 = ~pi007 & pi098;
assign w542 = ~pi054 & w541;
assign w543 = w455 & w542;
assign w544 = ~w540 & ~w543;
assign w545 = w476 & w538;
assign w546 = w544 & ~w545;
assign w547 = (pi001 & ~w509) | (pi001 & w17947) | (~w509 & w17947);
assign w548 = w546 & w17948;
assign w549 = ~w535 & w548;
assign w550 = ~w530 & ~w549;
assign w551 = ~w504 & ~w550;
assign w552 = ~w402 & w551;
assign w553 = w402 & ~w551;
assign w554 = ~w552 & ~w553;
assign w555 = w251 & ~w554;
assign w556 = ~w251 & w554;
assign w557 = ~w555 & ~w556;
assign w558 = pi069 & pi127;
assign w559 = ~pi063 & w558;
assign w560 = pi063 & ~pi126;
assign w561 = ~pi033 & pi069;
assign w562 = w560 & w561;
assign w563 = ~w559 & ~w562;
assign w564 = ~pi104 & ~w563;
assign w565 = pi063 & pi126;
assign w566 = ~pi033 & pi127;
assign w567 = w565 & w566;
assign w568 = ~pi069 & w567;
assign w569 = ~pi033 & pi063;
assign w570 = pi104 & pi127;
assign w571 = ~pi069 & w570;
assign w572 = ~pi063 & pi126;
assign w573 = pi033 & pi069;
assign w574 = w572 & w573;
assign w575 = w569 & w571;
assign w576 = ~w574 & ~w575;
assign w577 = ~w564 & w576;
assign w578 = (pi102 & ~w577) | (pi102 & w17949) | (~w577 & w17949);
assign w579 = pi033 & pi127;
assign w580 = pi069 & w560;
assign w581 = w579 & w580;
assign w582 = pi033 & ~pi069;
assign w583 = w565 & w582;
assign w584 = pi033 & ~pi126;
assign w585 = ~pi069 & ~pi127;
assign w586 = w584 & w585;
assign w587 = ~w583 & ~w586;
assign w588 = ~pi033 & ~pi063;
assign w589 = pi127 & w588;
assign w590 = w588 & w17950;
assign w591 = ~w581 & w587;
assign w592 = (~pi104 & ~w591) | (~pi104 & w17951) | (~w591 & w17951);
assign w593 = ~pi104 & pi126;
assign w594 = pi033 & pi126;
assign w595 = pi069 & w594;
assign w596 = (~pi127 & w595) | (~pi127 & w17952) | (w595 & w17952);
assign w597 = ~pi033 & pi104;
assign w598 = ~pi063 & ~pi126;
assign w599 = pi126 & w558;
assign w600 = ~w598 & ~w599;
assign w601 = (w597 & w599) | (w597 & w17953) | (w599 & w17953);
assign w602 = ~w596 & ~w601;
assign w603 = ~pi102 & ~w602;
assign w604 = pi069 & pi104;
assign w605 = w579 & w598;
assign w606 = w565 & w579;
assign w607 = ~pi033 & ~pi127;
assign w608 = w598 & w607;
assign w609 = ~w605 & ~w606;
assign w610 = (w604 & ~w609) | (w604 & w17954) | (~w609 & w17954);
assign w611 = ~w592 & ~w603;
assign w612 = ~w578 & w611;
assign w613 = pi127 & w560;
assign w614 = pi033 & pi063;
assign w615 = pi127 & w614;
assign w616 = ~w589 & ~w613;
assign w617 = ~pi069 & pi127;
assign w618 = w560 & w617;
assign w619 = pi033 & ~pi063;
assign w620 = pi069 & ~pi127;
assign w621 = w619 & w620;
assign w622 = ~pi069 & ~pi104;
assign w623 = w560 & w622;
assign w624 = ~pi033 & pi126;
assign w625 = w585 & w624;
assign w626 = ~pi126 & w614;
assign w627 = w614 & w17956;
assign w628 = pi104 & w625;
assign w629 = ~w627 & ~w628;
assign w630 = ~w618 & ~w621;
assign w631 = ~w623 & w630;
assign w632 = w629 & w631;
assign w633 = pi069 & w565;
assign w634 = w566 & w633;
assign w635 = ~pi033 & w622;
assign w636 = w572 & w635;
assign w637 = ~w634 & ~w636;
assign w638 = (w617 & w623) | (w617 & w17958) | (w623 & w17958);
assign w639 = pi104 & ~pi127;
assign w640 = pi069 & w639;
assign w641 = w569 & w640;
assign w642 = ~w638 & ~w641;
assign w643 = pi102 & ~w637;
assign w644 = w642 & ~w643;
assign w645 = pi102 & pi104;
assign w646 = pi063 & ~pi127;
assign w647 = ~w589 & ~w646;
assign w648 = ~pi069 & w598;
assign w649 = ~w580 & ~w648;
assign w650 = w647 & w649;
assign w651 = w645 & ~w650;
assign w652 = pi127 & w619;
assign w653 = w619 & w617;
assign w654 = w560 & w579;
assign w655 = w565 & w585;
assign w656 = ~w654 & ~w655;
assign w657 = (pi104 & ~w656) | (pi104 & w17959) | (~w656 & w17959);
assign w658 = ~w651 & ~w657;
assign w659 = w644 & w658;
assign w660 = pi033 & ~pi127;
assign w661 = w598 & w660;
assign w662 = (pi126 & w589) | (pi126 & w17960) | (w589 & w17960);
assign w663 = w565 & w607;
assign w664 = w560 & w573;
assign w665 = ~w663 & ~w664;
assign w666 = (~pi069 & w662) | (~pi069 & w17961) | (w662 & w17961);
assign w667 = w665 & ~w666;
assign w668 = ~pi102 & pi104;
assign w669 = w614 & w617;
assign w670 = ~pi063 & w561;
assign w671 = w561 & w598;
assign w672 = ~w634 & w17962;
assign w673 = w668 & ~w672;
assign w674 = ~pi127 & w624;
assign w675 = w624 & w620;
assign w676 = w594 & w617;
assign w677 = w587 & w17963;
assign w678 = pi104 & ~w676;
assign w679 = w585 & w626;
assign w680 = w558 & w588;
assign w681 = ~pi126 & w680;
assign w682 = ~w679 & ~w681;
assign w683 = ~pi033 & ~pi126;
assign w684 = ~w594 & ~w683;
assign w685 = w646 & ~w684;
assign w686 = pi033 & w598;
assign w687 = ~w652 & ~w686;
assign w688 = ~w685 & w687;
assign w689 = pi069 & ~pi104;
assign w690 = pi102 & w689;
assign w691 = ~w688 & w690;
assign w692 = ~pi104 & ~w682;
assign w693 = ~w691 & ~w692;
assign w694 = (~pi102 & w676) | (~pi102 & w17964) | (w676 & w17964);
assign w695 = ~w677 & w694;
assign w696 = w693 & w17965;
assign w697 = w645 & ~w667;
assign w698 = w696 & ~w697;
assign w699 = (pi012 & ~w659) | (pi012 & w17966) | (~w659 & w17966);
assign w700 = w698 & ~w699;
assign w701 = (~pi012 & ~w612) | (~pi012 & w17967) | (~w612 & w17967);
assign w702 = w700 & ~w701;
assign w703 = ~pi104 & ~pi127;
assign w704 = ~pi127 & w584;
assign w705 = w561 & w572;
assign w706 = ~w704 & ~w705;
assign w707 = ~pi033 & ~pi069;
assign w708 = w565 & w707;
assign w709 = ~w562 & ~w708;
assign w710 = ~pi104 & ~w709;
assign w711 = w614 & w17968;
assign w712 = w585 & w598;
assign w713 = w585 & w614;
assign w714 = ~w712 & ~w713;
assign w715 = ~w711 & w714;
assign w716 = ~w710 & w715;
assign w717 = pi127 & w624;
assign w718 = pi033 & w572;
assign w719 = w582 & w598;
assign w720 = ~w717 & ~w718;
assign w721 = (pi104 & ~w720) | (pi104 & w17969) | (~w720 & w17969);
assign w722 = w572 & w579;
assign w723 = w561 & w565;
assign w724 = ~w722 & ~w723;
assign w725 = ~pi033 & w598;
assign w726 = w598 & w17970;
assign w727 = ~w623 & ~w676;
assign w728 = w724 & w727;
assign w729 = ~w726 & w728;
assign w730 = (pi102 & ~w729) | (pi102 & w17971) | (~w729 & w17971);
assign w731 = w617 & w718;
assign w732 = w565 & w573;
assign w733 = ~w625 & ~w732;
assign w734 = ~w731 & w733;
assign w735 = ~pi104 & ~w734;
assign w736 = pi069 & w572;
assign w737 = ~pi033 & w572;
assign w738 = ~pi033 & w560;
assign w739 = ~w737 & ~w738;
assign w740 = (w570 & ~w739) | (w570 & w17972) | (~w739 & w17972);
assign w741 = w614 & w620;
assign w742 = ~pi126 & w741;
assign w743 = ~w735 & w17973;
assign w744 = ~w730 & w743;
assign w745 = (pi012 & ~w744) | (pi012 & w17974) | (~w744 & w17974);
assign w746 = ~pi127 & w683;
assign w747 = w582 & w613;
assign w748 = w703 & w718;
assign w749 = ~w705 & ~w748;
assign w750 = w558 & w594;
assign w751 = pi063 & w750;
assign w752 = pi126 & w713;
assign w753 = ~w751 & ~w752;
assign w754 = w749 & w753;
assign w755 = ~pi069 & pi104;
assign w756 = ~w588 & w755;
assign w757 = pi126 & w756;
assign w758 = ~w625 & ~w757;
assign w759 = w689 & w722;
assign w760 = ~w566 & ~w570;
assign w761 = w598 & ~w760;
assign w762 = ~w759 & ~w761;
assign w763 = w758 & w762;
assign w764 = ~pi102 & ~w763;
assign w765 = w560 & w558;
assign w766 = pi063 & w617;
assign w767 = w594 & w766;
assign w768 = ~w765 & ~w767;
assign w769 = (~pi104 & w767) | (~pi104 & w17976) | (w767 & w17976);
assign w770 = w620 & w683;
assign w771 = w565 & w660;
assign w772 = ~w770 & ~w771;
assign w773 = pi104 & ~w772;
assign w774 = w585 & w738;
assign w775 = ~w773 & ~w774;
assign w776 = ~w769 & w775;
assign w777 = ~w764 & w776;
assign w778 = (pi104 & ~w724) | (pi104 & w17978) | (~w724 & w17978);
assign w779 = w572 & w660;
assign w780 = ~pi127 & w560;
assign w781 = ~w589 & ~w780;
assign w782 = (w622 & ~w781) | (w622 & w17979) | (~w781 & w17979);
assign w783 = ~pi063 & w620;
assign w784 = w624 & w783;
assign w785 = w783 & w17980;
assign w786 = ~w778 & ~w782;
assign w787 = (pi102 & ~w786) | (pi102 & w17981) | (~w786 & w17981);
assign w788 = w560 & w755;
assign w789 = w607 & w788;
assign w790 = ~pi126 & w617;
assign w791 = w588 & w790;
assign w792 = ~w789 & ~w791;
assign w793 = w668 & ~w792;
assign w794 = w558 & w572;
assign w795 = w565 & w620;
assign w796 = ~w794 & ~w795;
assign w797 = w597 & ~w796;
assign w798 = ~pi104 & w565;
assign w799 = w558 & w738;
assign w800 = ~pi102 & w620;
assign w801 = w798 & w800;
assign w802 = ~w799 & ~w801;
assign w803 = ~w797 & w802;
assign w804 = ~w793 & w803;
assign w805 = ~w787 & w804;
assign w806 = (~pi012 & ~w777) | (~pi012 & w17982) | (~w777 & w17982);
assign w807 = w805 & ~w806;
assign w808 = ~w745 & w807;
assign w809 = ~w702 & w808;
assign w810 = w702 & ~w808;
assign w811 = ~w809 & ~w810;
assign w812 = w598 & w707;
assign w813 = ~pi127 & w812;
assign w814 = w561 & ~w598;
assign w815 = ~w752 & ~w814;
assign w816 = (~pi104 & ~w815) | (~pi104 & w17983) | (~w815 & w17983);
assign w817 = w604 & w686;
assign w818 = pi127 & w788;
assign w819 = ~w784 & ~w818;
assign w820 = w560 & w607;
assign w821 = w604 & w615;
assign w822 = w689 & w820;
assign w823 = ~w821 & ~w822;
assign w824 = (pi102 & ~w633) | (pi102 & w17984) | (~w633 & w17984);
assign w825 = w823 & w824;
assign w826 = ~w817 & w819;
assign w827 = w825 & w826;
assign w828 = ~w816 & w827;
assign w829 = ~w558 & ~w585;
assign w830 = w737 & ~w829;
assign w831 = ~w621 & ~w830;
assign w832 = pi033 & ~w649;
assign w833 = w831 & ~w832;
assign w834 = pi104 & ~w833;
assign w835 = w569 & w790;
assign w836 = w594 & w620;
assign w837 = pi063 & w836;
assign w838 = ~w835 & ~w837;
assign w839 = (~pi104 & ~w838) | (~pi104 & w17985) | (~w838 & w17985);
assign w840 = ~pi127 & w719;
assign w841 = ~w581 & ~w840;
assign w842 = w823 & w841;
assign w843 = ~pi102 & w842;
assign w844 = ~w834 & ~w839;
assign w845 = w843 & w844;
assign w846 = ~w828 & ~w845;
assign w847 = pi033 & w620;
assign w848 = ~pi063 & w593;
assign w849 = ~w711 & ~w765;
assign w850 = w717 & w755;
assign w851 = w849 & ~w850;
assign w852 = ~w847 & w848;
assign w853 = ~w566 & w852;
assign w854 = w851 & ~w853;
assign w855 = pi102 & ~w854;
assign w856 = w558 & w598;
assign w857 = pi063 & w607;
assign w858 = ~w856 & ~w857;
assign w859 = ~w601 & ~w755;
assign w860 = ~w858 & ~w859;
assign w861 = ~w615 & ~w725;
assign w862 = pi104 & ~w861;
assign w863 = ~pi126 & ~w707;
assign w864 = ~w623 & ~w783;
assign w865 = w863 & ~w864;
assign w866 = ~w862 & ~w865;
assign w867 = w567 & w622;
assign w868 = (~pi012 & ~w719) | (~pi012 & w17986) | (~w719 & w17986);
assign w869 = ~w867 & w868;
assign w870 = (w869 & w866) | (w869 & w17987) | (w866 & w17987);
assign w871 = pi104 & ~w705;
assign w872 = ~w771 & ~w783;
assign w873 = w871 & w872;
assign w874 = ~w790 & w873;
assign w875 = ~pi104 & ~w723;
assign w876 = w560 & w620;
assign w877 = w875 & ~w876;
assign w878 = ~w813 & w877;
assign w879 = ~w874 & ~w878;
assign w880 = (pi102 & ~w790) | (pi102 & w17988) | (~w790 & w17988);
assign w881 = ~pi104 & ~w598;
assign w882 = ~w781 & w881;
assign w883 = w572 & w639;
assign w884 = w584 & w783;
assign w885 = w880 & ~w882;
assign w886 = ~w883 & ~w884;
assign w887 = w885 & w886;
assign w888 = ~pi104 & w856;
assign w889 = ~pi069 & ~w703;
assign w890 = ~pi102 & ~w795;
assign w891 = pi104 & w722;
assign w892 = w890 & ~w891;
assign w893 = w594 & ~w889;
assign w894 = w892 & w17989;
assign w895 = ~w887 & ~w894;
assign w896 = pi012 & ~w879;
assign w897 = ~w895 & w896;
assign w898 = ~w855 & w870;
assign w899 = ~w860 & w898;
assign w900 = ~w897 & ~w899;
assign w901 = ~w846 & ~w900;
assign w902 = ~pi159 & w901;
assign w903 = pi159 & ~w901;
assign w904 = ~w902 & ~w903;
assign w905 = w811 & w904;
assign w906 = ~w811 & ~w904;
assign w907 = ~w905 & ~w906;
assign w908 = (~pi529 & w557) | (~pi529 & w17990) | (w557 & w17990);
assign w909 = w557 & ~w907;
assign w910 = w908 & ~w909;
assign w911 = ~pi159 & pi490;
assign w912 = pi529 & ~w911;
assign w913 = pi159 & ~pi490;
assign w914 = w912 & ~w913;
assign w915 = ~w910 & ~w914;
assign w916 = pi007 & w455;
assign w917 = w403 & w448;
assign w918 = ~w916 & ~w917;
assign w919 = ~pi114 & ~w918;
assign w920 = ~pi054 & w403;
assign w921 = w486 & w920;
assign w922 = w435 & w455;
assign w923 = ~w468 & ~w921;
assign w924 = ~w919 & w923;
assign w925 = (pi001 & ~w924) | (pi001 & w17991) | (~w924 & w17991);
assign w926 = ~pi114 & w541;
assign w927 = w413 & w435;
assign w928 = pi007 & w536;
assign w929 = w456 & w928;
assign w930 = ~w927 & ~w929;
assign w931 = ~w474 & ~w926;
assign w932 = w930 & w931;
assign w933 = ~pi001 & ~w932;
assign w934 = w415 & w442;
assign w935 = ~pi013 & pi021;
assign w936 = w435 & w935;
assign w937 = ~w934 & ~w936;
assign w938 = w408 & w466;
assign w939 = ~w525 & w937;
assign w940 = (~pi114 & ~w939) | (~pi114 & w17992) | (~w939 & w17992);
assign w941 = pi054 & w428;
assign w942 = w408 & w425;
assign w943 = ~w941 & ~w942;
assign w944 = w928 & ~w943;
assign w945 = w408 & w418;
assign w946 = w448 & w945;
assign w947 = (~pi029 & ~w945) | (~pi029 & w17993) | (~w945 & w17993);
assign w948 = ~w944 & w947;
assign w949 = ~w940 & w948;
assign w950 = ~pi013 & w408;
assign w951 = ~w453 & ~w950;
assign w952 = ~w406 & ~w524;
assign w953 = w951 & w952;
assign w954 = pi114 & ~w953;
assign w955 = w479 & w507;
assign w956 = ~w540 & ~w955;
assign w957 = (pi001 & w954) | (pi001 & w17994) | (w954 & w17994);
assign w958 = pi007 & ~pi114;
assign w959 = ~w475 & ~w507;
assign w960 = ~w507 & w17995;
assign w961 = w403 & w17935;
assign w962 = ~w505 & ~w961;
assign w963 = w442 & w456;
assign w964 = ~w418 & w538;
assign w965 = pi114 & w963;
assign w966 = ~w964 & ~w965;
assign w967 = w962 & w966;
assign w968 = (~pi001 & ~w967) | (~pi001 & w17996) | (~w967 & w17996);
assign w969 = pi098 & w442;
assign w970 = w442 & w428;
assign w971 = ~pi021 & pi054;
assign w972 = w411 & w971;
assign w973 = w403 & w425;
assign w974 = ~w972 & ~w973;
assign w975 = (pi114 & ~w974) | (pi114 & w17997) | (~w974 & w17997);
assign w976 = ~pi007 & w536;
assign w977 = w411 & w415;
assign w978 = pi029 & ~w977;
assign w979 = w519 & w976;
assign w980 = w978 & ~w979;
assign w981 = w538 & w958;
assign w982 = w980 & ~w981;
assign w983 = ~w957 & ~w968;
assign w984 = ~w975 & w982;
assign w985 = w983 & w984;
assign w986 = ~w925 & w949;
assign w987 = ~w933 & w986;
assign w988 = ~w985 & ~w987;
assign w989 = w519 & w541;
assign w990 = w417 & w466;
assign w991 = ~w454 & ~w990;
assign w992 = ~pi007 & ~pi021;
assign w993 = w415 & w992;
assign w994 = ~pi013 & ~w993;
assign w995 = w991 & w994;
assign w996 = ~w478 & w536;
assign w997 = ~w995 & ~w996;
assign w998 = ~w454 & ~w516;
assign w999 = ~w541 & w971;
assign w1000 = (pi013 & ~w998) | (pi013 & w17998) | (~w998 & w17998);
assign w1001 = (pi001 & w1000) | (pi001 & w5136) | (w1000 & w5136);
assign w1002 = ~w989 & ~w997;
assign w1003 = w1001 & ~w1002;
assign w1004 = w411 & w435;
assign w1005 = w413 & w456;
assign w1006 = (~pi114 & ~w937) | (~pi114 & w17999) | (~w937 & w17999);
assign w1007 = (~pi001 & w1006) | (~pi001 & w18000) | (w1006 & w18000);
assign w1008 = w442 & w478;
assign w1009 = ~pi054 & w433;
assign w1010 = ~w1008 & ~w1009;
assign w1011 = ~pi001 & pi114;
assign w1012 = w411 & w475;
assign w1013 = w408 & w448;
assign w1014 = ~w1012 & ~w1013;
assign w1015 = ~w540 & w1014;
assign w1016 = w1011 & ~w1015;
assign w1017 = ~pi114 & ~w1010;
assign w1018 = ~w1016 & ~w1017;
assign w1019 = ~w1007 & w1018;
assign w1020 = ~w1003 & w1019;
assign w1021 = ~w988 & w1020;
assign w1022 = ~pi023 & pi047;
assign w1023 = pi023 & w257;
assign w1024 = ~w1022 & ~w1023;
assign w1025 = w256 & w1024;
assign w1026 = pi123 & ~w1025;
assign w1027 = ~pi111 & w353;
assign w1028 = ~w287 & ~w1027;
assign w1029 = pi093 & ~w1028;
assign w1030 = ~pi027 & w294;
assign w1031 = pi047 & w295;
assign w1032 = w295 & w315;
assign w1033 = ~w1030 & ~w1032;
assign w1034 = w1029 & ~w1033;
assign w1035 = ~w1026 & ~w1034;
assign w1036 = w254 & ~w379;
assign w1037 = ~pi111 & w274;
assign w1038 = pi023 & ~w282;
assign w1039 = ~w1037 & w1038;
assign w1040 = w277 & w314;
assign w1041 = w270 & w254;
assign w1042 = ~w263 & ~w1041;
assign w1043 = pi123 & w1040;
assign w1044 = w1042 & ~w1043;
assign w1045 = (~pi123 & w1039) | (~pi123 & w18001) | (w1039 & w18001);
assign w1046 = w1044 & ~w1045;
assign w1047 = pi023 & w282;
assign w1048 = ~w377 & ~w1047;
assign w1049 = w326 & w18002;
assign w1050 = (~w1049 & w1048) | (~w1049 & w18003) | (w1048 & w18003);
assign w1051 = pi123 & ~w1050;
assign w1052 = w359 & w383;
assign w1053 = w270 & w285;
assign w1054 = ~w1052 & w18004;
assign w1055 = ~pi123 & w1041;
assign w1056 = w1054 & ~w1055;
assign w1057 = ~w1051 & w1056;
assign w1058 = ~pi048 & ~w1046;
assign w1059 = w1057 & ~w1058;
assign w1060 = pi048 & ~w1035;
assign w1061 = w1059 & ~w1060;
assign w1062 = ~pi047 & w286;
assign w1063 = ~pi093 & ~pi111;
assign w1064 = w315 & w1063;
assign w1065 = ~w1062 & ~w1064;
assign w1066 = ~pi123 & ~w1065;
assign w1067 = w272 & w386;
assign w1068 = w264 & w317;
assign w1069 = ~w365 & ~w1067;
assign w1070 = ~w1066 & w1069;
assign w1071 = ~pi123 & w314;
assign w1072 = w266 & w383;
assign w1073 = ~w1071 & ~w1072;
assign w1074 = w261 & w317;
assign w1075 = w252 & w18005;
assign w1076 = ~w1074 & ~w1075;
assign w1077 = (~pi048 & ~w1073) | (~pi048 & w18006) | (~w1073 & w18006);
assign w1078 = w252 & w295;
assign w1079 = (~pi123 & w288) | (~pi123 & w20756) | (w288 & w20756);
assign w1080 = pi023 & pi111;
assign w1081 = w252 & w1080;
assign w1082 = w311 & w326;
assign w1083 = ~w1081 & ~w1082;
assign w1084 = w383 & ~w1083;
assign w1085 = w274 & w376;
assign w1086 = w281 & w376;
assign w1087 = ~w1085 & ~w1086;
assign w1088 = ~pi123 & ~w1087;
assign w1089 = w257 & w281;
assign w1090 = w383 & w1089;
assign w1091 = ~w1084 & ~w1088;
assign w1092 = (~pi020 & ~w1089) | (~pi020 & w18007) | (~w1089 & w18007);
assign w1093 = w1091 & w1092;
assign w1094 = w1093 & w18008;
assign w1095 = (pi048 & ~w1070) | (pi048 & w20757) | (~w1070 & w20757);
assign w1096 = w1094 & ~w1095;
assign w1097 = w272 & w314;
assign w1098 = (pi093 & w1023) | (pi093 & w18009) | (w1023 & w18009);
assign w1099 = ~pi027 & ~w283;
assign w1100 = ~w1098 & w1099;
assign w1101 = ~w384 & ~w1100;
assign w1102 = ~w327 & ~w396;
assign w1103 = w282 & ~w314;
assign w1104 = (pi027 & ~w1102) | (pi027 & w18010) | (~w1102 & w18010);
assign w1105 = (pi048 & w1104) | (pi048 & w1416) | (w1104 & w1416);
assign w1106 = ~w1097 & ~w1101;
assign w1107 = w1105 & ~w1106;
assign w1108 = ~pi023 & w265;
assign w1109 = w311 & w376;
assign w1110 = w394 & w1108;
assign w1111 = ~w1109 & ~w1110;
assign w1112 = ~w1088 & w1111;
assign w1113 = ~pi048 & ~w1112;
assign w1114 = pi047 & w1086;
assign w1115 = w286 & w1063;
assign w1116 = ~pi047 & w1115;
assign w1117 = ~w1114 & ~w1116;
assign w1118 = ~pi048 & pi123;
assign w1119 = w326 & w270;
assign w1120 = w252 & w379;
assign w1121 = ~w388 & w18011;
assign w1122 = w1118 & ~w1121;
assign w1123 = ~pi123 & ~w1117;
assign w1124 = ~w1122 & ~w1123;
assign w1125 = ~w1113 & w1124;
assign w1126 = ~w1107 & w1125;
assign w1127 = ~w1061 & ~w1096;
assign w1128 = w1126 & ~w1127;
assign w1129 = ~w1021 & w1128;
assign w1130 = w1021 & ~w1128;
assign w1131 = ~w1129 & ~w1130;
assign w1132 = w408 & w5073;
assign w1133 = ~w467 & ~w1132;
assign w1134 = pi114 & ~w1133;
assign w1135 = (pi007 & w955) | (pi007 & w18012) | (w955 & w18012);
assign w1136 = pi054 & ~w417;
assign w1137 = w413 & ~w1136;
assign w1138 = ~w1134 & ~w1135;
assign w1139 = (pi001 & w409) | (pi001 & w18013) | (w409 & w18013);
assign w1140 = ~w445 & ~w519;
assign w1141 = pi013 & ~w1140;
assign w1142 = w425 & w428;
assign w1143 = ~w977 & ~w1142;
assign w1144 = ~w1141 & w1143;
assign w1145 = pi054 & w433;
assign w1146 = ~w927 & ~w1145;
assign w1147 = w541 & w405;
assign w1148 = ~pi013 & w426;
assign w1149 = ~w1147 & ~w1148;
assign w1150 = w1146 & w1149;
assign w1151 = pi114 & ~w1150;
assign w1152 = w403 & w466;
assign w1153 = pi001 & w1152;
assign w1154 = w403 & w17942;
assign w1155 = ~w543 & ~w1154;
assign w1156 = ~w1153 & w1155;
assign w1157 = (~pi114 & ~w1144) | (~pi114 & w18014) | (~w1144 & w18014);
assign w1158 = ~w1151 & w20758;
assign w1159 = (~pi001 & ~w1138) | (~pi001 & w18015) | (~w1138 & w18015);
assign w1160 = pi098 & w432;
assign w1161 = ~w487 & ~w1160;
assign w1162 = w446 & ~w1161;
assign w1163 = ~pi021 & w445;
assign w1164 = w456 & w479;
assign w1165 = ~w950 & ~w1164;
assign w1166 = ~w1163 & w1165;
assign w1167 = ~w1162 & w1166;
assign w1168 = ~pi013 & ~w998;
assign w1169 = (~pi001 & w1168) | (~pi001 & w18016) | (w1168 & w18016);
assign w1170 = pi013 & pi098;
assign w1171 = w475 & w1170;
assign w1172 = ~w443 & ~w1171;
assign w1173 = ~w1148 & w1172;
assign w1174 = ~pi114 & ~w1173;
assign w1175 = ~w509 & ~w519;
assign w1176 = w976 & ~w1175;
assign w1177 = w435 & ~w446;
assign w1178 = w1011 & w1177;
assign w1179 = ~w1176 & ~w1178;
assign w1180 = ~w1174 & w1179;
assign w1181 = ~w1169 & w1180;
assign w1182 = ~w498 & ~w531;
assign w1183 = w538 & w1182;
assign w1184 = w403 & w469;
assign w1185 = w469 & w18017;
assign w1186 = w509 & w928;
assign w1187 = pi114 & w442;
assign w1188 = ~w959 & w1187;
assign w1189 = ~w1188 & w18018;
assign w1190 = (~pi114 & w1183) | (~pi114 & w20759) | (w1183 & w20759);
assign w1191 = w507 & w536;
assign w1192 = ~pi114 & w1004;
assign w1193 = ~w921 & ~w1192;
assign w1194 = ~w416 & ~w444;
assign w1195 = w1193 & w1194;
assign w1196 = w958 & w1170;
assign w1197 = w418 & w1154;
assign w1198 = pi021 & w1196;
assign w1199 = ~w1197 & ~w1198;
assign w1200 = (w1195 & w20760) | (w1195 & w20761) | (w20760 & w20761);
assign w1201 = (~pi001 & w1190) | (~pi001 & w18020) | (w1190 & w18020);
assign w1202 = w1200 & ~w1201;
assign w1203 = (~pi029 & ~w1181) | (~pi029 & w18021) | (~w1181 & w18021);
assign w1204 = w1202 & ~w1203;
assign w1205 = (pi029 & ~w1158) | (pi029 & w18022) | (~w1158 & w18022);
assign w1206 = w1204 & ~w1205;
assign w1207 = (pi048 & w299) | (pi048 & w18023) | (w299 & w18023);
assign w1208 = ~w272 & ~w281;
assign w1209 = pi027 & ~w1208;
assign w1210 = ~w1053 & ~w1209;
assign w1211 = w1210 & w18024;
assign w1212 = ~pi123 & ~w1211;
assign w1213 = w252 & w277;
assign w1214 = ~w364 & ~w1213;
assign w1215 = (pi123 & ~w1214) | (pi123 & w18025) | (~w1214 & w18025);
assign w1216 = ~w329 & ~w1086;
assign w1217 = pi027 & w395;
assign w1218 = w1216 & ~w1217;
assign w1219 = w296 & w353;
assign w1220 = w1218 & ~w1219;
assign w1221 = (~pi048 & ~w1220) | (~pi048 & w18026) | (~w1220 & w18026);
assign w1222 = ~pi047 & w1109;
assign w1223 = w285 & w1062;
assign w1224 = ~w1222 & ~w1223;
assign w1225 = ~pi023 & w257;
assign w1226 = ~w262 & ~w1225;
assign w1227 = pi093 & ~w1226;
assign w1228 = w1224 & ~w1227;
assign w1229 = w254 & w295;
assign w1230 = w254 & w376;
assign w1231 = ~w390 & ~w1230;
assign w1232 = pi048 & w1229;
assign w1233 = w1231 & ~w1232;
assign w1234 = pi123 & ~w1228;
assign w1235 = w1233 & ~w1234;
assign w1236 = ~w1212 & ~w1221;
assign w1237 = w1235 & w1236;
assign w1238 = pi020 & ~w1237;
assign w1239 = pi027 & w274;
assign w1240 = w270 & w294;
assign w1241 = ~w1239 & ~w1240;
assign w1242 = (~w259 & w1241) | (~w259 & w18027) | (w1241 & w18027);
assign w1243 = ~pi123 & ~w1242;
assign w1244 = ~pi027 & ~w1102;
assign w1245 = w310 & ~w1244;
assign w1246 = w252 & ~w286;
assign w1247 = pi048 & ~w1246;
assign w1248 = w345 & w383;
assign w1249 = w1247 & ~w1248;
assign w1250 = ~w1029 & w1249;
assign w1251 = ~w1245 & ~w1250;
assign w1252 = ~w283 & ~w359;
assign w1253 = w383 & ~w1252;
assign w1254 = ~w315 & w317;
assign w1255 = w1118 & w1254;
assign w1256 = ~w1253 & ~w1255;
assign w1257 = ~w1251 & w18028;
assign w1258 = ~pi020 & ~w1257;
assign w1259 = ~pi111 & w254;
assign w1260 = w258 & w1259;
assign w1261 = ~w284 & ~w1041;
assign w1262 = (~pi123 & ~w1261) | (~pi123 & w18029) | (~w1261 & w18029);
assign w1263 = w383 & w1081;
assign w1264 = w285 & w394;
assign w1265 = w1022 & w1264;
assign w1266 = ~w1263 & ~w1265;
assign w1267 = (~pi048 & w1262) | (~pi048 & w18030) | (w1262 & w18030);
assign w1268 = (pi123 & w273) | (pi123 & w18031) | (w273 & w18031);
assign w1269 = ~pi123 & w1109;
assign w1270 = ~w303 & ~w333;
assign w1271 = ~w1269 & w1270;
assign w1272 = (pi048 & ~w1271) | (pi048 & w18032) | (~w1271 & w18032);
assign w1273 = w376 & w1022;
assign w1274 = (w1118 & w260) | (w1118 & w18033) | (w260 & w18033);
assign w1275 = ~pi123 & ~w315;
assign w1276 = w311 & w394;
assign w1277 = (~w1275 & w1114) | (~w1275 & w18034) | (w1114 & w18034);
assign w1278 = ~w1274 & ~w1277;
assign w1279 = ~w1272 & w1278;
assign w1280 = ~w1267 & w1279;
assign w1281 = ~w1258 & w1280;
assign w1282 = ~w1238 & w1281;
assign w1283 = ~w1206 & w1282;
assign w1284 = w1206 & ~w1282;
assign w1285 = ~w1283 & ~w1284;
assign w1286 = w1131 & ~w1285;
assign w1287 = ~w1131 & w1285;
assign w1288 = ~w1286 & ~w1287;
assign w1289 = w7 & w17893;
assign w1290 = ~pi107 & w16;
assign w1291 = (~pi083 & w1290) | (~pi083 & w18035) | (w1290 & w18035);
assign w1292 = w40 & w173;
assign w1293 = w8 & w29;
assign w1294 = pi083 & w151;
assign w1295 = ~w1293 & ~w1294;
assign w1296 = ~w237 & ~w1292;
assign w1297 = w1295 & w1296;
assign w1298 = w7 & w0;
assign w1299 = ~pi107 & w20;
assign w1300 = ~w104 & ~w1299;
assign w1301 = (~pi083 & ~w1300) | (~pi083 & w18036) | (~w1300 & w18036);
assign w1302 = pi107 & w11;
assign w1303 = ~w24 & ~w1302;
assign w1304 = pi083 & ~w1303;
assign w1305 = ~w80 & w91;
assign w1306 = ~w125 & ~w1305;
assign w1307 = ~w1304 & w1306;
assign w1308 = ~w172 & ~w1292;
assign w1309 = ~pi083 & ~w1308;
assign w1310 = (w8 & w135) | (w8 & w18037) | (w135 & w18037);
assign w1311 = w1 & w164;
assign w1312 = w1 & w18038;
assign w1313 = ~w1310 & ~w1312;
assign w1314 = ~w1309 & w18039;
assign w1315 = (pi040 & ~w1307) | (pi040 & w20762) | (~w1307 & w20762);
assign w1316 = w1314 & ~w1315;
assign w1317 = (~pi040 & ~w1297) | (~pi040 & w18040) | (~w1297 & w18040);
assign w1318 = ~w103 & ~w196;
assign w1319 = ~w61 & ~w235;
assign w1320 = (pi083 & ~w1319) | (pi083 & w18041) | (~w1319 & w18041);
assign w1321 = w1318 & ~w1320;
assign w1322 = w0 & w25;
assign w1323 = ~w114 & ~w1322;
assign w1324 = ~w78 & w178;
assign w1325 = w1323 & ~w1324;
assign w1326 = ~pi014 & w191;
assign w1327 = ~pi014 & ~w158;
assign w1328 = ~w16 & ~w49;
assign w1329 = w1327 & ~w1328;
assign w1330 = w2 & w23;
assign w1331 = ~w13 & ~w49;
assign w1332 = ~w114 & ~w1330;
assign w1333 = w1331 & w1332;
assign w1334 = ~pi083 & ~w1333;
assign w1335 = ~w1329 & ~w1334;
assign w1336 = (~pi040 & ~w1325) | (~pi040 & w18042) | (~w1325 & w18042);
assign w1337 = w1335 & ~w1336;
assign w1338 = (pi078 & ~w1337) | (pi078 & w18043) | (~w1337 & w18043);
assign w1339 = ~w231 & w18044;
assign w1340 = ~pi083 & ~w1339;
assign w1341 = ~pi082 & w1322;
assign w1342 = w20 & w34;
assign w1343 = ~w1341 & ~w1342;
assign w1344 = (~pi040 & w1340) | (~pi040 & w18045) | (w1340 & w18045);
assign w1345 = ~w57 & ~w103;
assign w1346 = pi014 & ~w1345;
assign w1347 = (w88 & w1346) | (w88 & w18046) | (w1346 & w18046);
assign w1348 = pi040 & ~pi083;
assign w1349 = w70 & ~w107;
assign w1350 = ~w135 & ~w146;
assign w1351 = ~w1349 & ~w1350;
assign w1352 = w50 & w56;
assign w1353 = (w1348 & w1351) | (w1348 & w18047) | (w1351 & w18047);
assign w1354 = w15 & w83;
assign w1355 = ~w166 & ~w1354;
assign w1356 = ~w211 & w1355;
assign w1357 = w123 & ~w1356;
assign w1358 = w40 & w135;
assign w1359 = w135 & w18048;
assign w1360 = ~w238 & ~w1359;
assign w1361 = ~w1347 & ~w1353;
assign w1362 = ~w1357 & w1360;
assign w1363 = w1361 & w1362;
assign w1364 = ~w1344 & w1363;
assign w1365 = ~w1338 & w1364;
assign w1366 = (~pi078 & ~w1316) | (~pi078 & w18049) | (~w1316 & w18049);
assign w1367 = w1365 & ~w1366;
assign w1368 = pi023 & w317;
assign w1369 = ~w1085 & ~w1368;
assign w1370 = pi123 & ~w1369;
assign w1371 = w255 & ~w295;
assign w1372 = ~w1120 & ~w1371;
assign w1373 = ~w1370 & w1372;
assign w1374 = w277 & w377;
assign w1375 = ~w1229 & ~w1374;
assign w1376 = ~w334 & ~w1230;
assign w1377 = pi123 & ~w1376;
assign w1378 = w287 & w1063;
assign w1379 = ~w276 & ~w1378;
assign w1380 = ~w1377 & w1379;
assign w1381 = (~pi123 & w1374) | (~pi123 & w18051) | (w1374 & w18051);
assign w1382 = ~w276 & ~w1222;
assign w1383 = ~pi123 & ~w1382;
assign w1384 = (w343 & w299) | (w343 & w18052) | (w299 & w18052);
assign w1385 = w252 & w258;
assign w1386 = ~w1263 & ~w1385;
assign w1387 = ~w1384 & w1386;
assign w1388 = ~w1383 & w1387;
assign w1389 = (~pi048 & ~w1380) | (~pi048 & w18053) | (~w1380 & w18053);
assign w1390 = w1388 & ~w1389;
assign w1391 = w315 & w1368;
assign w1392 = ~w1097 & ~w1391;
assign w1393 = ~w1031 & ~w1108;
assign w1394 = (pi123 & ~w1393) | (pi123 & w18055) | (~w1393 & w18055);
assign w1395 = w1392 & ~w1394;
assign w1396 = pi027 & w294;
assign w1397 = ~pi027 & w282;
assign w1398 = w285 & w286;
assign w1399 = ~w396 & ~w1398;
assign w1400 = w314 & w1397;
assign w1401 = w1399 & ~w1400;
assign w1402 = ~w396 & ~w1068;
assign w1403 = ~w1081 & ~w1230;
assign w1404 = w1402 & w1403;
assign w1405 = w1037 & ~w1071;
assign w1406 = ~pi123 & ~w1404;
assign w1407 = (~pi027 & w1405) | (~pi027 & w18056) | (w1405 & w18056);
assign w1408 = ~w1406 & ~w1407;
assign w1409 = (~pi048 & ~w1401) | (~pi048 & w18057) | (~w1401 & w18057);
assign w1410 = w1408 & ~w1409;
assign w1411 = (pi020 & ~w1410) | (pi020 & w18058) | (~w1410 & w18058);
assign w1412 = ~w300 & w18059;
assign w1413 = ~pi123 & ~w1412;
assign w1414 = ~w267 & ~w1223;
assign w1415 = (~pi048 & w1413) | (~pi048 & w18060) | (w1413 & w18060);
assign w1416 = pi048 & pi123;
assign w1417 = ~w350 & ~w1097;
assign w1418 = pi027 & ~w1417;
assign w1419 = (w1416 & w1418) | (w1416 & w18061) | (w1418 & w18061);
assign w1420 = pi048 & ~pi123;
assign w1421 = ~w1368 & w1397;
assign w1422 = w281 & w326;
assign w1423 = ~w1089 & ~w1422;
assign w1424 = ~w1421 & w1423;
assign w1425 = w1420 & ~w1424;
assign w1426 = ~pi048 & w343;
assign w1427 = ~pi023 & w252;
assign w1428 = ~w389 & ~w1082;
assign w1429 = (w1426 & ~w1428) | (w1426 & w18062) | (~w1428 & w18062);
assign w1430 = w1120 & w1420;
assign w1431 = pi023 & pi123;
assign w1432 = w324 & w1431;
assign w1433 = ~w1090 & ~w1430;
assign w1434 = ~w1432 & w1433;
assign w1435 = ~w1429 & w1434;
assign w1436 = w1435 & w18063;
assign w1437 = ~w1415 & w1436;
assign w1438 = ~w1411 & w1437;
assign w1439 = (~pi020 & ~w1390) | (~pi020 & w18064) | (~w1390 & w18064);
assign w1440 = w1438 & ~w1439;
assign w1441 = ~w1367 & w1440;
assign w1442 = w1367 & ~w1440;
assign w1443 = ~w1441 & ~w1442;
assign w1444 = w566 & w560;
assign w1445 = ~pi127 & w708;
assign w1446 = (~pi104 & w1445) | (~pi104 & w18065) | (w1445 & w18065);
assign w1447 = ~w597 & ~w660;
assign w1448 = w633 & ~w1447;
assign w1449 = w560 & w582;
assign w1450 = pi104 & w1449;
assign w1451 = ~w799 & ~w1448;
assign w1452 = ~w1450 & w1451;
assign w1453 = pi069 & w569;
assign w1454 = w569 & w558;
assign w1455 = ~pi127 & w588;
assign w1456 = ~pi069 & w572;
assign w1457 = ~w1455 & ~w1456;
assign w1458 = (~pi104 & ~w1457) | (~pi104 & w18066) | (~w1457 & w18066);
assign w1459 = pi127 & w594;
assign w1460 = ~w583 & ~w1459;
assign w1461 = pi104 & ~w1460;
assign w1462 = ~w566 & w580;
assign w1463 = ~w671 & ~w1462;
assign w1464 = ~w1461 & w1463;
assign w1465 = w559 & w584;
assign w1466 = ~pi126 & w585;
assign w1467 = ~w812 & ~w1466;
assign w1468 = ~w1465 & w1467;
assign w1469 = pi104 & ~w1468;
assign w1470 = w579 & w848;
assign w1471 = w848 & w18067;
assign w1472 = w689 & w771;
assign w1473 = ~w712 & ~w1472;
assign w1474 = ~w1471 & w1473;
assign w1475 = ~w1469 & w1474;
assign w1476 = (pi102 & ~w1464) | (pi102 & w18068) | (~w1464 & w18068);
assign w1477 = w1475 & ~w1476;
assign w1478 = (~pi102 & ~w1452) | (~pi102 & w18069) | (~w1452 & w18069);
assign w1479 = ~w663 & ~w751;
assign w1480 = ~w633 & ~w674;
assign w1481 = (pi104 & ~w1480) | (pi104 & w18070) | (~w1480 & w18070);
assign w1482 = w1479 & ~w1481;
assign w1483 = w558 & w584;
assign w1484 = ~w820 & ~w1483;
assign w1485 = ~w639 & w736;
assign w1486 = w1484 & ~w1485;
assign w1487 = w660 & w1456;
assign w1488 = ~w605 & ~w708;
assign w1489 = w889 & ~w1488;
assign w1490 = ~w574 & ~w605;
assign w1491 = ~w820 & ~w1449;
assign w1492 = w1490 & w1491;
assign w1493 = ~pi104 & ~w1492;
assign w1494 = ~w1489 & ~w1493;
assign w1495 = (~pi102 & ~w1486) | (~pi102 & w18071) | (~w1486 & w18071);
assign w1496 = w1494 & ~w1495;
assign w1497 = (pi012 & ~w1496) | (pi012 & w18072) | (~w1496 & w18072);
assign w1498 = w560 & w660;
assign w1499 = w585 & w619;
assign w1500 = ~w1498 & ~w1499;
assign w1501 = ~w608 & ~w719;
assign w1502 = w1500 & w1501;
assign w1503 = w689 & w725;
assign w1504 = (~w1503 & w1502) | (~w1503 & w18073) | (w1502 & w18073);
assign w1505 = ~w562 & ~w836;
assign w1506 = ~w791 & w1505;
assign w1507 = w559 & w684;
assign w1508 = (~w1507 & w1506) | (~w1507 & w18074) | (w1506 & w18074);
assign w1509 = ~w615 & ~w663;
assign w1510 = pi069 & ~w1509;
assign w1511 = (w645 & w1510) | (w645 & w18075) | (w1510 & w18075);
assign w1512 = w572 & w707;
assign w1513 = ~w712 & ~w1512;
assign w1514 = ~w767 & w1513;
assign w1515 = w668 & ~w1514;
assign w1516 = ~pi127 & w598;
assign w1517 = w604 & w1516;
assign w1518 = ~w794 & ~w1517;
assign w1519 = (w597 & w1517) | (w597 & w18076) | (w1517 & w18076);
assign w1520 = ~w1515 & ~w1519;
assign w1521 = ~w1511 & w1520;
assign w1522 = ~pi102 & ~w1508;
assign w1523 = pi102 & ~w1504;
assign w1524 = w1521 & w18077;
assign w1525 = ~w1497 & w1524;
assign w1526 = (~pi012 & ~w1477) | (~pi012 & w18078) | (~w1477 & w18078);
assign w1527 = w1525 & ~w1526;
assign w1528 = w1525 & w18079;
assign w1529 = (pi267 & ~w1525) | (pi267 & w18080) | (~w1525 & w18080);
assign w1530 = ~w1528 & ~w1529;
assign w1531 = w1443 & w1530;
assign w1532 = ~w1443 & ~w1530;
assign w1533 = ~w1531 & ~w1532;
assign w1534 = ~w1288 & ~w1533;
assign w1535 = ~pi529 & ~w1534;
assign w1536 = w1288 & w1533;
assign w1537 = w1535 & ~w1536;
assign w1538 = pi267 & pi503;
assign w1539 = pi529 & ~w1538;
assign w1540 = ~pi267 & ~pi503;
assign w1541 = w1539 & ~w1540;
assign w1542 = ~w1537 & ~w1541;
assign w1543 = pi061 & pi105;
assign w1544 = pi032 & ~pi064;
assign w1545 = w1543 & w1544;
assign w1546 = ~pi067 & w1545;
assign w1547 = (~pi117 & ~w1545) | (~pi117 & w1665) | (~w1545 & w1665);
assign w1548 = pi061 & ~pi064;
assign w1549 = pi032 & ~pi067;
assign w1550 = w1548 & w1549;
assign w1551 = ~w1547 & w1550;
assign w1552 = pi032 & pi067;
assign w1553 = ~pi061 & w1552;
assign w1554 = pi061 & ~pi105;
assign w1555 = ~pi064 & pi067;
assign w1556 = w1554 & w1555;
assign w1557 = ~w1553 & ~w1556;
assign w1558 = ~pi061 & pi067;
assign w1559 = pi064 & pi105;
assign w1560 = w1558 & w1559;
assign w1561 = (~w1560 & w1557) | (~w1560 & w18081) | (w1557 & w18081);
assign w1562 = ~w1551 & w1561;
assign w1563 = pi002 & ~w1562;
assign w1564 = ~pi061 & ~pi064;
assign w1565 = pi032 & w1564;
assign w1566 = w1564 & w18082;
assign w1567 = pi064 & ~pi067;
assign w1568 = w1543 & w1567;
assign w1569 = pi064 & ~pi105;
assign w1570 = ~pi032 & ~pi067;
assign w1571 = w1569 & w1570;
assign w1572 = ~w1568 & ~w1571;
assign w1573 = pi064 & w1554;
assign w1574 = w1552 & w1573;
assign w1575 = ~w1566 & w1572;
assign w1576 = (~pi117 & ~w1575) | (~pi117 & w18083) | (~w1575 & w18083);
assign w1577 = pi067 & pi117;
assign w1578 = pi032 & pi064;
assign w1579 = w1543 & w1578;
assign w1580 = ~pi032 & ~pi105;
assign w1581 = w1564 & w1580;
assign w1582 = ~pi061 & ~pi105;
assign w1583 = w1578 & w1582;
assign w1584 = ~w1579 & ~w1581;
assign w1585 = (w1577 & ~w1584) | (w1577 & w18084) | (~w1584 & w18084);
assign w1586 = pi105 & w1552;
assign w1587 = ~w1582 & ~w1586;
assign w1588 = ~pi002 & pi117;
assign w1589 = pi064 & pi067;
assign w1590 = pi117 & ~w1589;
assign w1591 = ~pi032 & pi105;
assign w1592 = ~pi002 & w1591;
assign w1593 = ~w1590 & w1592;
assign w1594 = ~pi036 & ~w1593;
assign w1595 = ~pi064 & w1588;
assign w1596 = ~w1587 & w1595;
assign w1597 = w1594 & ~w1596;
assign w1598 = ~w1585 & w1597;
assign w1599 = ~w1576 & w1598;
assign w1600 = ~w1563 & w1599;
assign w1601 = ~pi032 & pi061;
assign w1602 = pi067 & w1554;
assign w1603 = ~pi067 & w1582;
assign w1604 = ~w1601 & ~w1603;
assign w1605 = ~w1565 & ~w1602;
assign w1606 = w1604 & w1605;
assign w1607 = w1554 & w1578;
assign w1608 = ~pi061 & pi064;
assign w1609 = w1549 & w1608;
assign w1610 = ~w1607 & ~w1609;
assign w1611 = w1543 & w1570;
assign w1612 = pi002 & ~w1606;
assign w1613 = (pi117 & w1612) | (pi117 & w18085) | (w1612 & w18085);
assign w1614 = ~w1565 & ~w1573;
assign w1615 = pi061 & pi064;
assign w1616 = pi032 & w1615;
assign w1617 = pi032 & w1554;
assign w1618 = ~w1616 & ~w1617;
assign w1619 = w1614 & w1618;
assign w1620 = ~pi117 & ~w1619;
assign w1621 = ~pi064 & ~pi067;
assign w1622 = w1591 & w1621;
assign w1623 = ~pi032 & pi067;
assign w1624 = w1608 & w1623;
assign w1625 = ~pi032 & pi117;
assign w1626 = ~pi067 & w1554;
assign w1627 = ~w1625 & w1626;
assign w1628 = ~w1624 & ~w1627;
assign w1629 = pi117 & w1622;
assign w1630 = w1628 & ~w1629;
assign w1631 = ~w1620 & w1630;
assign w1632 = ~pi002 & ~w1631;
assign w1633 = pi067 & w1545;
assign w1634 = ~pi061 & pi105;
assign w1635 = ~pi117 & w1621;
assign w1636 = w1634 & w1635;
assign w1637 = ~w1633 & ~w1636;
assign w1638 = ~pi032 & w1577;
assign w1639 = ~pi067 & ~pi117;
assign w1640 = w1549 & w1569;
assign w1641 = pi036 & ~w1640;
assign w1642 = w1617 & w1639;
assign w1643 = w1641 & ~w1642;
assign w1644 = w1548 & w1638;
assign w1645 = w1643 & ~w1644;
assign w1646 = pi002 & ~w1637;
assign w1647 = w1645 & ~w1646;
assign w1648 = ~w1632 & w18086;
assign w1649 = ~w1600 & ~w1648;
assign w1650 = w1559 & w1601;
assign w1651 = ~pi064 & ~pi105;
assign w1652 = w1601 & w1651;
assign w1653 = ~w1650 & ~w1652;
assign w1654 = ~w1591 & w1608;
assign w1655 = (pi067 & ~w1653) | (pi067 & w18087) | (~w1653 & w18087);
assign w1656 = ~pi117 & ~w1655;
assign w1657 = ~pi067 & w1591;
assign w1658 = w1615 & w1657;
assign w1659 = ~pi067 & w1634;
assign w1660 = w1544 & w1659;
assign w1661 = ~w1658 & ~w1660;
assign w1662 = w1570 & w1582;
assign w1663 = pi064 & w1662;
assign w1664 = w1554 & w1589;
assign w1665 = pi067 & ~pi117;
assign w1666 = w1548 & w1591;
assign w1667 = ~w1664 & ~w1666;
assign w1668 = ~w1663 & w1667;
assign w1669 = ~w1665 & w1668;
assign w1670 = (pi002 & ~w1669) | (pi002 & w18088) | (~w1669 & w18088);
assign w1671 = ~w1656 & w1670;
assign w1672 = pi061 & w1549;
assign w1673 = w1549 & w1615;
assign w1674 = w1558 & w1651;
assign w1675 = ~w1633 & w18089;
assign w1676 = w1588 & ~w1675;
assign w1677 = ~pi032 & pi064;
assign w1678 = w1626 & w1677;
assign w1679 = ~pi064 & w1582;
assign w1680 = w1552 & w1679;
assign w1681 = ~w1678 & ~w1680;
assign w1682 = ~pi117 & ~w1572;
assign w1683 = w1549 & w1559;
assign w1684 = ~pi064 & w1591;
assign w1685 = w1665 & w1684;
assign w1686 = ~w1683 & ~w1685;
assign w1687 = ~w1682 & w1686;
assign w1688 = ~pi002 & ~w1687;
assign w1689 = ~pi117 & ~w1681;
assign w1690 = ~w1688 & w18090;
assign w1691 = ~w1671 & w1690;
assign w1692 = ~w1649 & w1691;
assign w1693 = pi008 & pi059;
assign w1694 = ~pi056 & w1693;
assign w1695 = pi056 & ~pi099;
assign w1696 = pi008 & ~pi095;
assign w1697 = w1695 & w1696;
assign w1698 = ~w1694 & ~w1697;
assign w1699 = ~pi115 & ~w1698;
assign w1700 = pi056 & ~pi095;
assign w1701 = ~pi008 & pi059;
assign w1702 = pi115 & w1701;
assign w1703 = w1700 & w1702;
assign w1704 = pi056 & pi099;
assign w1705 = pi059 & ~pi095;
assign w1706 = w1704 & w1705;
assign w1707 = ~pi008 & w1706;
assign w1708 = ~pi056 & pi099;
assign w1709 = pi008 & pi095;
assign w1710 = w1708 & w1709;
assign w1711 = ~w1703 & ~w1707;
assign w1712 = ~w1699 & w1711;
assign w1713 = (pi026 & ~w1712) | (pi026 & w18091) | (~w1712 & w18091);
assign w1714 = pi008 & w1695;
assign w1715 = pi059 & pi095;
assign w1716 = w1714 & w1715;
assign w1717 = ~pi008 & pi095;
assign w1718 = w1704 & w1717;
assign w1719 = ~pi008 & ~pi059;
assign w1720 = pi095 & ~pi099;
assign w1721 = w1719 & w1720;
assign w1722 = ~w1718 & ~w1721;
assign w1723 = ~pi056 & ~pi099;
assign w1724 = w1705 & w1723;
assign w1725 = ~w1716 & w1722;
assign w1726 = (~pi115 & ~w1725) | (~pi115 & w18092) | (~w1725 & w18092);
assign w1727 = ~pi056 & ~pi095;
assign w1728 = ~pi099 & pi115;
assign w1729 = w1727 & w1728;
assign w1730 = pi008 & pi115;
assign w1731 = pi059 & w1730;
assign w1732 = ~pi095 & pi099;
assign w1733 = w1731 & w1732;
assign w1734 = ~pi059 & ~pi115;
assign w1735 = pi099 & w1734;
assign w1736 = pi095 & pi099;
assign w1737 = pi008 & ~pi059;
assign w1738 = w1736 & w1737;
assign w1739 = ~w1729 & ~w1735;
assign w1740 = ~w1733 & w1739;
assign w1741 = pi095 & w1704;
assign w1742 = w1715 & w1723;
assign w1743 = ~w1741 & ~w1742;
assign w1744 = ~pi059 & ~pi099;
assign w1745 = w1727 & w1744;
assign w1746 = w1730 & w1745;
assign w1747 = (~pi030 & ~w1745) | (~pi030 & w18093) | (~w1745 & w18093);
assign w1748 = w1731 & ~w1743;
assign w1749 = w1747 & ~w1748;
assign w1750 = (~pi026 & ~w1740) | (~pi026 & w18094) | (~w1740 & w18094);
assign w1751 = w1749 & ~w1750;
assign w1752 = pi056 & ~pi059;
assign w1753 = pi059 & w1727;
assign w1754 = ~pi008 & w1723;
assign w1755 = ~w1752 & ~w1754;
assign w1756 = ~w1714 & ~w1753;
assign w1757 = w1755 & w1756;
assign w1758 = pi099 & w1719;
assign w1759 = w1695 & w1715;
assign w1760 = ~pi056 & pi095;
assign w1761 = w1701 & w1760;
assign w1762 = ~w1759 & ~w1761;
assign w1763 = w1719 & w1704;
assign w1764 = w1762 & ~w1763;
assign w1765 = pi026 & ~w1757;
assign w1766 = ~pi059 & pi099;
assign w1767 = pi056 & pi095;
assign w1768 = ~w1766 & w1767;
assign w1769 = pi059 & w1695;
assign w1770 = ~w1753 & ~w1768;
assign w1771 = ~pi059 & pi115;
assign w1772 = ~pi008 & w1695;
assign w1773 = ~pi008 & pi115;
assign w1774 = ~pi095 & w1766;
assign w1775 = w1737 & w1760;
assign w1776 = w1773 & w1774;
assign w1777 = ~w1775 & ~w1776;
assign w1778 = ~w1771 & w1772;
assign w1779 = w1777 & ~w1778;
assign w1780 = (~pi026 & ~w1779) | (~pi026 & w18096) | (~w1779 & w18096);
assign w1781 = pi008 & w1704;
assign w1782 = w1705 & w1781;
assign w1783 = ~pi008 & ~pi095;
assign w1784 = w1708 & w1783;
assign w1785 = ~pi115 & w1784;
assign w1786 = ~w1782 & ~w1785;
assign w1787 = pi056 & w1701;
assign w1788 = w1701 & w1695;
assign w1789 = ~pi059 & w1700;
assign w1790 = w1730 & w1789;
assign w1791 = w1701 & w1720;
assign w1792 = pi030 & ~w1791;
assign w1793 = ~w1790 & w1792;
assign w1794 = ~pi115 & w1788;
assign w1795 = w1793 & ~w1794;
assign w1796 = pi026 & ~w1786;
assign w1797 = w1795 & ~w1796;
assign w1798 = ~w1780 & w1797;
assign w1799 = (pi115 & w1765) | (pi115 & w18097) | (w1765 & w18097);
assign w1800 = w1798 & ~w1799;
assign w1801 = ~w1713 & w1751;
assign w1802 = ~w1726 & w1801;
assign w1803 = ~w1800 & ~w1802;
assign w1804 = ~pi095 & ~pi099;
assign w1805 = w1752 & w1804;
assign w1806 = w1766 & w1767;
assign w1807 = ~w1805 & ~w1806;
assign w1808 = w1760 & ~w1766;
assign w1809 = w1696 & w1723;
assign w1810 = ~pi059 & w1695;
assign w1811 = w1717 & w1810;
assign w1812 = (~pi115 & ~w1810) | (~pi115 & w18098) | (~w1810 & w18098);
assign w1813 = pi059 & w1809;
assign w1814 = w1812 & ~w1813;
assign w1815 = (pi008 & ~w1807) | (pi008 & w18099) | (~w1807 & w18099);
assign w1816 = w1814 & ~w1815;
assign w1817 = w1732 & w1752;
assign w1818 = ~pi059 & w1720;
assign w1819 = w1720 & w18100;
assign w1820 = w1705 & w1708;
assign w1821 = ~w1817 & ~w1820;
assign w1822 = w1821 & w18101;
assign w1823 = ~pi008 & ~w1822;
assign w1824 = w1695 & w1709;
assign w1825 = ~w1817 & ~w1824;
assign w1826 = pi115 & w1825;
assign w1827 = ~w1823 & w1826;
assign w1828 = (pi026 & w1827) | (pi026 & w18102) | (w1827 & w18102);
assign w1829 = (pi115 & ~w1781) | (pi115 & w20763) | (~w1781 & w20763);
assign w1830 = w1701 & w1767;
assign w1831 = ~w1809 & ~w1830;
assign w1832 = w1722 & w1814;
assign w1833 = w1829 & w1831;
assign w1834 = ~w1832 & ~w1833;
assign w1835 = w1696 & w1735;
assign w1836 = w1701 & w1736;
assign w1837 = ~pi026 & ~w1836;
assign w1838 = ~w1835 & w1837;
assign w1839 = ~w1834 & w1838;
assign w1840 = ~w1828 & ~w1839;
assign w1841 = ~w1803 & ~w1840;
assign w1842 = ~w1692 & w1841;
assign w1843 = w1692 & ~w1841;
assign w1844 = ~w1842 & ~w1843;
assign w1845 = w1582 & w1621;
assign w1846 = ~w1545 & ~w1607;
assign w1847 = (pi117 & ~w1846) | (pi117 & w18103) | (~w1846 & w18103);
assign w1848 = ~pi117 & w1660;
assign w1849 = pi064 & ~w1634;
assign w1850 = w1623 & ~w1849;
assign w1851 = ~w1571 & ~w1850;
assign w1852 = ~w1848 & w1851;
assign w1853 = (~pi002 & ~w1852) | (~pi002 & w18104) | (~w1852 & w18104);
assign w1854 = pi105 & w1609;
assign w1855 = w1552 & w1569;
assign w1856 = ~pi061 & w1855;
assign w1857 = ~w1854 & ~w1856;
assign w1858 = w1564 & w1591;
assign w1859 = w1559 & w1623;
assign w1860 = ~w1858 & ~w1859;
assign w1861 = (pi117 & ~w1857) | (pi117 & w18105) | (~w1857 & w18105);
assign w1862 = ~w1548 & ~w1580;
assign w1863 = pi067 & ~w1862;
assign w1864 = ~w1579 & ~w1640;
assign w1865 = ~w1863 & w1864;
assign w1866 = ~pi117 & ~w1865;
assign w1867 = w1582 & w18106;
assign w1868 = w1544 & w1554;
assign w1869 = ~pi117 & w1615;
assign w1870 = ~w1868 & ~w1869;
assign w1871 = (pi002 & ~w1870) | (pi002 & w18107) | (~w1870 & w18107);
assign w1872 = w1554 & w1567;
assign w1873 = w1558 & w1684;
assign w1874 = ~w1872 & ~w1873;
assign w1875 = ~w1866 & w18108;
assign w1876 = ~w1853 & w1875;
assign w1877 = (pi036 & ~w1876) | (pi036 & w18109) | (~w1876 & w18109);
assign w1878 = pi064 & pi117;
assign w1879 = w1621 & w18110;
assign w1880 = w1602 & w1878;
assign w1881 = ~w1879 & ~w1880;
assign w1882 = ~w1553 & ~w1587;
assign w1883 = w1881 & ~w1882;
assign w1884 = w1552 & w1582;
assign w1885 = ~pi117 & w1884;
assign w1886 = ~pi067 & ~w1653;
assign w1887 = w1564 & w1570;
assign w1888 = w1543 & w1589;
assign w1889 = ~w1887 & ~w1888;
assign w1890 = ~w1854 & w1889;
assign w1891 = ~pi117 & ~w1890;
assign w1892 = pi064 & w1582;
assign w1893 = ~w1548 & ~w1892;
assign w1894 = w1638 & ~w1893;
assign w1895 = pi064 & w1634;
assign w1896 = ~w1568 & ~w1895;
assign w1897 = w1588 & ~w1896;
assign w1898 = ~w1894 & ~w1897;
assign w1899 = ~w1891 & w1898;
assign w1900 = (~pi002 & w1886) | (~pi002 & w18111) | (w1886 & w18111);
assign w1901 = w1899 & ~w1900;
assign w1902 = w1570 & w1615;
assign w1903 = ~pi067 & w1858;
assign w1904 = (pi117 & w1903) | (pi117 & w18112) | (w1903 & w18112);
assign w1905 = w1878 & w1884;
assign w1906 = ~pi032 & w1664;
assign w1907 = w1626 & ~w1677;
assign w1908 = ~w1906 & ~w1907;
assign w1909 = (pi117 & ~w1884) | (pi117 & w18113) | (~w1884 & w18113);
assign w1910 = ~w1663 & ~w1905;
assign w1911 = w1908 & w1910;
assign w1912 = (~w1904 & w1911) | (~w1904 & w18114) | (w1911 & w18114);
assign w1913 = ~pi002 & ~w1912;
assign w1914 = ~pi064 & w1554;
assign w1915 = pi117 & w1549;
assign w1916 = w1914 & w1915;
assign w1917 = w1623 & w1892;
assign w1918 = ~pi067 & w1581;
assign w1919 = w1555 & w1634;
assign w1920 = pi117 & w1919;
assign w1921 = ~w1918 & ~w1920;
assign w1922 = ~pi117 & w1683;
assign w1923 = w1921 & ~w1922;
assign w1924 = ~w1916 & ~w1917;
assign w1925 = (pi002 & ~w1923) | (pi002 & w18115) | (~w1923 & w18115);
assign w1926 = w1552 & w18110;
assign w1927 = ~pi067 & pi117;
assign w1928 = w1573 & w1927;
assign w1929 = w1586 & w18116;
assign w1930 = w1573 & w18117;
assign w1931 = ~w1929 & ~w1930;
assign w1932 = ~w1925 & w1931;
assign w1933 = ~w1913 & w1932;
assign w1934 = (~pi036 & ~w1901) | (~pi036 & w18118) | (~w1901 & w18118);
assign w1935 = w1933 & ~w1934;
assign w1936 = ~w1877 & w1935;
assign w1937 = w1723 & w1783;
assign w1938 = ~w1706 & ~w1759;
assign w1939 = (pi115 & ~w1938) | (pi115 & w18119) | (~w1938 & w18119);
assign w1940 = ~pi095 & w1708;
assign w1941 = w1701 & w1940;
assign w1942 = ~pi059 & w1696;
assign w1943 = w1708 & w1737;
assign w1944 = ~w1721 & ~w1942;
assign w1945 = ~w1943 & w1944;
assign w1946 = w1940 & w18120;
assign w1947 = w1945 & ~w1946;
assign w1948 = (~pi026 & ~w1947) | (~pi026 & w18121) | (~w1947 & w18121);
assign w1949 = ~pi099 & w1727;
assign w1950 = (pi026 & w1949) | (pi026 & w18122) | (w1949 & w18122);
assign w1951 = ~w1700 & ~w1744;
assign w1952 = pi008 & ~w1951;
assign w1953 = w1704 & w1715;
assign w1954 = ~w1791 & ~w1953;
assign w1955 = ~w1952 & w1954;
assign w1956 = ~pi059 & w1727;
assign w1957 = ~w1761 & ~w1956;
assign w1958 = pi099 & ~w1957;
assign w1959 = w1693 & w1720;
assign w1960 = ~pi056 & w1959;
assign w1961 = ~w1738 & ~w1960;
assign w1962 = ~w1958 & w1961;
assign w1963 = pi115 & ~w1962;
assign w1964 = ~pi059 & w1708;
assign w1965 = w1696 & w1964;
assign w1966 = w1695 & w1705;
assign w1967 = w1695 & w1717;
assign w1968 = pi026 & w1966;
assign w1969 = ~w1967 & ~w1968;
assign w1970 = ~w1965 & w1969;
assign w1971 = ~w1963 & w1970;
assign w1972 = (~pi115 & ~w1955) | (~pi115 & w18123) | (~w1955 & w18123);
assign w1973 = w1971 & w18124;
assign w1974 = pi030 & ~w1973;
assign w1975 = ~pi099 & ~pi115;
assign w1976 = (~pi026 & ~w1694) | (~pi026 & w18125) | (~w1694 & w18125);
assign w1977 = ~pi008 & ~w1807;
assign w1978 = w1976 & ~w1977;
assign w1979 = pi099 & w1693;
assign w1980 = ~w1723 & ~w1979;
assign w1981 = ~w1694 & ~w1980;
assign w1982 = pi095 & w1695;
assign w1983 = w1695 & w18126;
assign w1984 = ~pi008 & ~pi115;
assign w1985 = w1732 & w1984;
assign w1986 = pi026 & ~w1985;
assign w1987 = pi008 & w1983;
assign w1988 = w1986 & ~w1987;
assign w1989 = ~w1981 & w1988;
assign w1990 = ~w1978 & ~w1989;
assign w1991 = pi099 & w1761;
assign w1992 = w1704 & w1709;
assign w1993 = w1727 & w1719;
assign w1994 = ~w1991 & w18127;
assign w1995 = ~pi115 & ~w1994;
assign w1996 = ~pi026 & pi115;
assign w1997 = pi095 & w1708;
assign w1998 = ~w1718 & ~w1997;
assign w1999 = w1996 & ~w1998;
assign w2000 = pi095 & w1737;
assign w2001 = w1723 & w2000;
assign w2002 = w2000 & w18128;
assign w2003 = ~w1790 & ~w2002;
assign w2004 = ~w1999 & w2003;
assign w2005 = ~w1995 & w2004;
assign w2006 = ~w1990 & w2005;
assign w2007 = ~pi095 & w1695;
assign w2008 = w1719 & w2007;
assign w2009 = pi095 & w1723;
assign w2010 = w1719 & w2009;
assign w2011 = ~w1788 & ~w2008;
assign w2012 = (~pi115 & ~w2011) | (~pi115 & w18129) | (~w2011 & w18129);
assign w2013 = w1709 & w1975;
assign w2014 = w1752 & w2013;
assign w2015 = w1731 & w2009;
assign w2016 = ~w2014 & ~w2015;
assign w2017 = (~pi026 & w2012) | (~pi026 & w18130) | (w2012 & w18130);
assign w2018 = w1719 & w1949;
assign w2019 = pi059 & w1736;
assign w2020 = w1696 & w1708;
assign w2021 = pi115 & w2020;
assign w2022 = w1702 & w2007;
assign w2023 = ~w2021 & ~w2022;
assign w2024 = w1984 & w2019;
assign w2025 = w2023 & ~w2024;
assign w2026 = ~w2001 & ~w2018;
assign w2027 = (pi026 & ~w2025) | (pi026 & w18131) | (~w2025 & w18131);
assign w2028 = w1719 & w1767;
assign w2029 = w1719 & w1940;
assign w2030 = (w1996 & w2029) | (w1996 & w18132) | (w2029 & w18132);
assign w2031 = pi115 & w1719;
assign w2032 = w1693 & w18133;
assign w2033 = w1982 & w2031;
assign w2034 = pi056 & w2032;
assign w2035 = ~w2033 & ~w2034;
assign w2036 = ~w2030 & w2035;
assign w2037 = ~w2027 & w2036;
assign w2038 = ~w2017 & w2037;
assign w2039 = ~pi030 & ~w2006;
assign w2040 = w2038 & ~w2039;
assign w2041 = ~w1974 & w2040;
assign w2042 = ~w1936 & w2041;
assign w2043 = w1936 & ~w2041;
assign w2044 = ~w2042 & ~w2043;
assign w2045 = w1844 & ~w2044;
assign w2046 = ~w1844 & w2044;
assign w2047 = ~w2045 & ~w2046;
assign w2048 = pi085 & ~pi087;
assign w2049 = pi046 & ~pi050;
assign w2050 = w2048 & w2049;
assign w2051 = ~pi028 & ~pi085;
assign w2052 = pi046 & pi050;
assign w2053 = ~pi087 & w2052;
assign w2054 = w2051 & w2053;
assign w2055 = (~pi092 & w2054) | (~pi092 & w18134) | (w2054 & w18134);
assign w2056 = pi028 & ~pi085;
assign w2057 = w2052 & w2056;
assign w2058 = pi087 & w2057;
assign w2059 = pi087 & w2049;
assign w2060 = ~pi028 & pi092;
assign w2061 = w2059 & w2060;
assign w2062 = pi028 & ~pi087;
assign w2063 = w2052 & w2062;
assign w2064 = pi092 & w2063;
assign w2065 = w2049 & w2062;
assign w2066 = pi085 & w2065;
assign w2067 = ~w2058 & ~w2061;
assign w2068 = ~w2064 & ~w2066;
assign w2069 = w2067 & w2068;
assign w2070 = (~pi089 & ~w2069) | (~pi089 & w18135) | (~w2069 & w18135);
assign w2071 = pi046 & pi085;
assign w2072 = w2062 & w2071;
assign w2073 = ~pi046 & ~pi087;
assign w2074 = ~pi085 & w2073;
assign w2075 = ~pi046 & pi050;
assign w2076 = ~w2072 & ~w2074;
assign w2077 = ~pi028 & pi087;
assign w2078 = w2052 & w2077;
assign w2079 = pi050 & pi087;
assign w2080 = pi085 & w2079;
assign w2081 = ~w2078 & ~w2080;
assign w2082 = pi092 & ~w2081;
assign w2083 = pi028 & w2049;
assign w2084 = ~w2048 & w2083;
assign w2085 = ~pi046 & ~pi050;
assign w2086 = w2062 & w2085;
assign w2087 = ~w2084 & ~w2086;
assign w2088 = ~w2082 & w2087;
assign w2089 = (pi089 & ~w2088) | (pi089 & w18137) | (~w2088 & w18137);
assign w2090 = w2051 & w2085;
assign w2091 = (~pi092 & ~w2057) | (~pi092 & w18138) | (~w2057 & w18138);
assign w2092 = ~pi028 & pi085;
assign w2093 = pi087 & w2075;
assign w2094 = w2092 & w2093;
assign w2095 = pi028 & pi085;
assign w2096 = pi087 & w2085;
assign w2097 = w2095 & w2096;
assign w2098 = ~pi028 & ~pi087;
assign w2099 = w2085 & w2098;
assign w2100 = ~pi050 & w2051;
assign w2101 = ~w2099 & ~w2100;
assign w2102 = ~w2097 & w2101;
assign w2103 = pi092 & w2102;
assign w2104 = w2091 & ~w2094;
assign w2105 = ~w2070 & ~w2089;
assign w2106 = (~w2090 & w2103) | (~w2090 & w18139) | (w2103 & w18139);
assign w2107 = pi050 & ~pi085;
assign w2108 = pi046 & ~pi087;
assign w2109 = w2107 & w2108;
assign w2110 = pi028 & w2052;
assign w2111 = pi085 & pi087;
assign w2112 = w2110 & w2111;
assign w2113 = ~w2109 & ~w2112;
assign w2114 = pi046 & w2048;
assign w2115 = ~pi087 & w2107;
assign w2116 = ~w2110 & ~w2114;
assign w2117 = (pi092 & ~w2116) | (pi092 & w18140) | (~w2116 & w18140);
assign w2118 = w2113 & ~w2117;
assign w2119 = ~pi046 & w2107;
assign w2120 = w2077 & w2119;
assign w2121 = ~pi050 & ~pi087;
assign w2122 = ~w2052 & w2095;
assign w2123 = ~w2121 & w2122;
assign w2124 = pi046 & ~pi085;
assign w2125 = w2121 & w2124;
assign w2126 = pi028 & ~pi092;
assign w2127 = w2075 & w2126;
assign w2128 = ~w2120 & ~w2123;
assign w2129 = ~w2125 & ~w2127;
assign w2130 = w2049 & w2077;
assign w2131 = w2085 & w2111;
assign w2132 = pi028 & pi087;
assign w2133 = w2075 & w2132;
assign w2134 = ~w2125 & ~w2130;
assign w2135 = ~w2131 & ~w2133;
assign w2136 = w2134 & w2135;
assign w2137 = ~w2096 & ~w2108;
assign w2138 = ~pi050 & pi087;
assign w2139 = w2092 & w2138;
assign w2140 = pi050 & w2060;
assign w2141 = ~w2139 & ~w2140;
assign w2142 = ~w2137 & ~w2141;
assign w2143 = w2048 & w2052;
assign w2144 = ~pi028 & w2143;
assign w2145 = ~w2142 & ~w2144;
assign w2146 = ~pi092 & ~w2136;
assign w2147 = w2145 & ~w2146;
assign w2148 = (~pi089 & ~w2128) | (~pi089 & w18141) | (~w2128 & w18141);
assign w2149 = w2147 & ~w2148;
assign w2150 = (pi053 & ~w2149) | (pi053 & w18142) | (~w2149 & w18142);
assign w2151 = w2073 & w2092;
assign w2152 = ~pi050 & w2151;
assign w2153 = w2056 & w2079;
assign w2154 = ~w2065 & ~w2153;
assign w2155 = ~w2152 & w2154;
assign w2156 = ~pi092 & ~w2155;
assign w2157 = pi028 & ~pi046;
assign w2158 = w2048 & w2157;
assign w2159 = pi050 & w2158;
assign w2160 = ~w2097 & ~w2159;
assign w2161 = (~pi089 & w2156) | (~pi089 & w18143) | (w2156 & w18143);
assign w2162 = pi089 & ~pi092;
assign w2163 = ~pi085 & pi087;
assign w2164 = w2049 & w2163;
assign w2165 = ~w2120 & ~w2164;
assign w2166 = w2077 & w2085;
assign w2167 = ~pi050 & ~pi085;
assign w2168 = w2073 & w2167;
assign w2169 = ~w2086 & ~w2166;
assign w2170 = ~w2168 & w2169;
assign w2171 = w2165 & w2170;
assign w2172 = pi089 & pi092;
assign w2173 = pi087 & w2071;
assign w2174 = ~w2109 & ~w2173;
assign w2175 = pi028 & ~w2174;
assign w2176 = (w2172 & w2175) | (w2172 & w18144) | (w2175 & w18144);
assign w2177 = ~pi089 & pi092;
assign w2178 = w2079 & w2092;
assign w2179 = pi046 & w2178;
assign w2180 = w2075 & w2098;
assign w2181 = ~w2090 & ~w2180;
assign w2182 = ~w2179 & w2181;
assign w2183 = w2177 & ~w2182;
assign w2184 = ~pi087 & w2085;
assign w2185 = pi092 & w2056;
assign w2186 = w2184 & w2185;
assign w2187 = pi028 & pi092;
assign w2188 = pi050 & w2048;
assign w2189 = w2187 & w2188;
assign w2190 = w2188 & w18145;
assign w2191 = ~w2186 & ~w2190;
assign w2192 = ~w2183 & w2191;
assign w2193 = ~w2176 & w2192;
assign w2194 = w2162 & ~w2171;
assign w2195 = w2193 & w18146;
assign w2196 = ~w2150 & w2195;
assign w2197 = (~pi053 & ~w2105) | (~pi053 & w18147) | (~w2105 & w18147);
assign w2198 = w2196 & ~w2197;
assign w2199 = ~pi008 & w1708;
assign w2200 = ~pi095 & ~w1752;
assign w2201 = ~w1753 & ~w1787;
assign w2202 = (~w2199 & ~w2201) | (~w2199 & w18148) | (~w2201 & w18148);
assign w2203 = ~w1718 & ~w2019;
assign w2204 = pi115 & ~w2203;
assign w2205 = ~w1705 & w1714;
assign w2206 = ~w1809 & ~w2205;
assign w2207 = ~w2204 & w2206;
assign w2208 = ~pi115 & ~w2202;
assign w2209 = w2207 & ~w2208;
assign w2210 = ~pi008 & w1817;
assign w2211 = (~pi115 & w2210) | (~pi115 & w18149) | (w2210 & w18149);
assign w2212 = w1696 & w1704;
assign w2213 = ~w1967 & ~w2212;
assign w2214 = pi115 & ~w2213;
assign w2215 = pi008 & w1806;
assign w2216 = pi059 & w1697;
assign w2217 = ~w2215 & ~w2216;
assign w2218 = ~w2214 & w2217;
assign w2219 = ~w1991 & ~w2215;
assign w2220 = ~pi115 & ~w2219;
assign w2221 = (w1773 & w1949) | (w1773 & w18150) | (w1949 & w18150);
assign w2222 = w1719 & w1723;
assign w2223 = ~w2015 & ~w2222;
assign w2224 = ~w2221 & w2223;
assign w2225 = ~w2220 & w2224;
assign w2226 = (~pi026 & ~w2218) | (~pi026 & w18151) | (~w2218 & w18151);
assign w2227 = w2225 & ~w2226;
assign w2228 = pi026 & ~w2209;
assign w2229 = w2227 & ~w2228;
assign w2230 = pi008 & w1953;
assign w2231 = ~w1817 & ~w2230;
assign w2232 = ~w1774 & ~w1781;
assign w2233 = (pi115 & ~w2232) | (pi115 & w18152) | (~w2232 & w18152);
assign w2234 = w2231 & ~w2233;
assign w2235 = w1717 & w1964;
assign w2236 = pi008 & w1708;
assign w2237 = ~w1771 & w2236;
assign w2238 = ~w1805 & ~w1959;
assign w2239 = ~w2235 & w2238;
assign w2240 = ~pi008 & ~w1734;
assign w2241 = w1704 & w1783;
assign w2242 = ~w1742 & ~w2241;
assign w2243 = w2240 & ~w2242;
assign w2244 = ~w1710 & ~w1742;
assign w2245 = ~w1805 & ~w1967;
assign w2246 = w2244 & w2245;
assign w2247 = ~pi115 & ~w2246;
assign w2248 = ~w2243 & ~w2247;
assign w2249 = (~pi026 & ~w2239) | (~pi026 & w18153) | (~w2239 & w18153);
assign w2250 = w2248 & ~w2249;
assign w2251 = (pi030 & ~w2250) | (pi030 & w18154) | (~w2250 & w18154);
assign w2252 = ~pi099 & w1701;
assign w2253 = w1727 & w2252;
assign w2254 = ~w1697 & ~w1738;
assign w2255 = ~w2253 & w2254;
assign w2256 = ~pi115 & ~w2255;
assign w2257 = w1727 & w1979;
assign w2258 = ~w1960 & ~w2257;
assign w2259 = (~pi026 & w2256) | (~pi026 & w18155) | (w2256 & w18155);
assign w2260 = pi026 & ~pi115;
assign w2261 = w1744 & w1767;
assign w2262 = w1717 & w1723;
assign w2263 = ~w1745 & ~w2261;
assign w2264 = ~w2235 & w2263;
assign w2265 = pi026 & pi115;
assign w2266 = pi059 & w1767;
assign w2267 = ~w1817 & ~w2266;
assign w2268 = pi008 & ~w2267;
assign w2269 = w1736 & w1787;
assign w2270 = ~w1784 & ~w2222;
assign w2271 = ~w2269 & w2270;
assign w2272 = w1996 & ~w2271;
assign w2273 = pi008 & pi026;
assign w2274 = w1727 & w1975;
assign w2275 = w2273 & w2274;
assign w2276 = ~w1746 & ~w2275;
assign w2277 = w2020 & w8537;
assign w2278 = w2276 & ~w2277;
assign w2279 = ~w2272 & w2278;
assign w2280 = (w2265 & w2268) | (w2265 & w18156) | (w2268 & w18156);
assign w2281 = w2279 & ~w2280;
assign w2282 = (w2260 & ~w2264) | (w2260 & w18157) | (~w2264 & w18157);
assign w2283 = w2281 & w18158;
assign w2284 = ~w2251 & w2283;
assign w2285 = ~pi030 & ~w2229;
assign w2286 = w2284 & ~w2285;
assign w2287 = ~w2198 & w2286;
assign w2288 = w2198 & ~w2286;
assign w2289 = ~w2287 & ~w2288;
assign w2290 = pi042 & ~pi071;
assign w2291 = pi075 & ~pi110;
assign w2292 = w2290 & w2291;
assign w2293 = pi042 & pi110;
assign w2294 = ~pi071 & ~pi079;
assign w2295 = w2293 & w2294;
assign w2296 = ~pi075 & w2295;
assign w2297 = (~pi080 & w2296) | (~pi080 & w18159) | (w2296 & w18159);
assign w2298 = pi071 & ~pi079;
assign w2299 = pi042 & ~pi110;
assign w2300 = w2298 & w2299;
assign w2301 = pi080 & w2300;
assign w2302 = pi075 & pi079;
assign w2303 = ~pi071 & w2299;
assign w2304 = w2302 & w2303;
assign w2305 = pi079 & w2293;
assign w2306 = pi071 & ~pi075;
assign w2307 = ~pi071 & pi080;
assign w2308 = ~w2306 & ~w2307;
assign w2309 = w2305 & ~w2308;
assign w2310 = ~w2301 & ~w2304;
assign w2311 = ~w2309 & w2310;
assign w2312 = pi075 & w2290;
assign w2313 = w2290 & w2302;
assign w2314 = ~pi042 & pi110;
assign w2315 = ~pi079 & w2314;
assign w2316 = ~pi042 & ~pi071;
assign w2317 = ~pi075 & w2316;
assign w2318 = ~w2315 & ~w2317;
assign w2319 = (~pi080 & ~w2318) | (~pi080 & w18160) | (~w2318 & w18160);
assign w2320 = w2293 & w2298;
assign w2321 = pi071 & pi110;
assign w2322 = pi075 & w2321;
assign w2323 = ~w2320 & ~w2322;
assign w2324 = pi080 & ~w2323;
assign w2325 = ~pi071 & pi075;
assign w2326 = pi079 & w2299;
assign w2327 = ~w2325 & w2326;
assign w2328 = ~pi071 & pi079;
assign w2329 = ~pi042 & ~pi110;
assign w2330 = w2328 & w2329;
assign w2331 = ~w2327 & ~w2330;
assign w2332 = ~w2324 & w2331;
assign w2333 = pi071 & ~pi110;
assign w2334 = ~pi042 & w2302;
assign w2335 = w2333 & w2334;
assign w2336 = w2294 & w2329;
assign w2337 = ~pi075 & ~pi079;
assign w2338 = ~pi110 & w2337;
assign w2339 = ~w2336 & ~w2338;
assign w2340 = ~w2335 & w2339;
assign w2341 = pi080 & ~w2340;
assign w2342 = pi079 & ~pi080;
assign w2343 = w2293 & w2306;
assign w2344 = w2342 & w2343;
assign w2345 = ~pi079 & ~pi080;
assign w2346 = ~pi042 & pi071;
assign w2347 = pi075 & pi110;
assign w2348 = w2346 & w2347;
assign w2349 = w2345 & w2348;
assign w2350 = w2329 & w2337;
assign w2351 = ~w2344 & ~w2349;
assign w2352 = ~w2350 & w2351;
assign w2353 = ~w2341 & w2352;
assign w2354 = (pi073 & ~w2332) | (pi073 & w18161) | (~w2332 & w18161);
assign w2355 = w2353 & ~w2354;
assign w2356 = (~pi073 & ~w2311) | (~pi073 & w18162) | (~w2311 & w18162);
assign w2357 = ~pi071 & ~pi075;
assign w2358 = w2293 & w2357;
assign w2359 = pi042 & pi071;
assign w2360 = pi110 & w2302;
assign w2361 = w2359 & w2360;
assign w2362 = ~w2358 & ~w2361;
assign w2363 = ~pi071 & pi110;
assign w2364 = ~w2305 & ~w2312;
assign w2365 = (pi080 & ~w2364) | (pi080 & w18163) | (~w2364 & w18163);
assign w2366 = w2362 & ~w2365;
assign w2367 = pi079 & w2314;
assign w2368 = ~pi075 & pi080;
assign w2369 = w2306 & w2314;
assign w2370 = w2299 & w2357;
assign w2371 = w2302 & w2333;
assign w2372 = ~w2370 & ~w2371;
assign w2373 = ~pi079 & w2369;
assign w2374 = w2372 & ~w2373;
assign w2375 = w2291 & w2346;
assign w2376 = pi071 & pi079;
assign w2377 = w2314 & w2376;
assign w2378 = ~w2300 & ~w2370;
assign w2379 = ~w2375 & ~w2377;
assign w2380 = w2378 & w2379;
assign w2381 = pi075 & ~pi079;
assign w2382 = pi042 & w2381;
assign w2383 = (~pi080 & ~w2381) | (~pi080 & w18164) | (~w2381 & w18164);
assign w2384 = w2346 & w2381;
assign w2385 = w2295 & ~w2383;
assign w2386 = ~pi110 & w2384;
assign w2387 = ~w2385 & ~w2386;
assign w2388 = ~pi080 & ~w2380;
assign w2389 = w2387 & ~w2388;
assign w2390 = (~pi073 & ~w2374) | (~pi073 & w18165) | (~w2374 & w18165);
assign w2391 = w2389 & ~w2390;
assign w2392 = (pi015 & ~w2391) | (pi015 & w18166) | (~w2391 & w18166);
assign w2393 = pi079 & w2321;
assign w2394 = w2321 & w5715;
assign w2395 = w2291 & w2316;
assign w2396 = ~pi079 & w2395;
assign w2397 = w2299 & w2328;
assign w2398 = ~w2396 & w18167;
assign w2399 = ~pi080 & ~w2398;
assign w2400 = w2316 & w2360;
assign w2401 = ~w2335 & ~w2400;
assign w2402 = (~pi073 & w2399) | (~pi073 & w18168) | (w2399 & w18168);
assign w2403 = pi073 & ~pi080;
assign w2404 = ~pi042 & w2298;
assign w2405 = w2316 & w18169;
assign w2406 = w2299 & w2306;
assign w2407 = ~w2330 & ~w2406;
assign w2408 = ~w2405 & w2407;
assign w2409 = pi073 & pi080;
assign w2410 = pi075 & w2359;
assign w2411 = ~w2358 & ~w2410;
assign w2412 = pi079 & ~w2411;
assign w2413 = pi075 & w2295;
assign w2414 = (w2409 & w2412) | (w2409 & w18170) | (w2412 & w18170);
assign w2415 = ~pi073 & pi080;
assign w2416 = w2321 & w2382;
assign w2417 = w2294 & w2314;
assign w2418 = ~w2350 & ~w2417;
assign w2419 = ~w2416 & w2418;
assign w2420 = w2415 & ~w2419;
assign w2421 = pi079 & pi080;
assign w2422 = w2316 & w2347;
assign w2423 = ~w2405 & ~w2422;
assign w2424 = w2421 & ~w2423;
assign w2425 = ~w2420 & ~w2424;
assign w2426 = ~w2414 & w2425;
assign w2427 = (w2403 & ~w2408) | (w2403 & w18171) | (~w2408 & w18171);
assign w2428 = w2426 & w18172;
assign w2429 = ~w2392 & w2428;
assign w2430 = (~pi015 & ~w2355) | (~pi015 & w18173) | (~w2355 & w18173);
assign w2431 = w2429 & ~w2430;
assign w2432 = w2429 & w18174;
assign w2433 = (pi268 & ~w2429) | (pi268 & w18175) | (~w2429 & w18175);
assign w2434 = ~w2432 & ~w2433;
assign w2435 = w2289 & w2434;
assign w2436 = ~w2289 & ~w2434;
assign w2437 = ~w2435 & ~w2436;
assign w2438 = ~w2047 & w2437;
assign w2439 = ~pi529 & ~w2438;
assign w2440 = w2047 & ~w2437;
assign w2441 = w2439 & ~w2440;
assign w2442 = ~pi268 & pi527;
assign w2443 = pi529 & ~w2442;
assign w2444 = pi268 & ~pi527;
assign w2445 = w2443 & ~w2444;
assign w2446 = ~w2441 & ~w2445;
assign w2447 = ~pi045 & pi081;
assign w2448 = ~pi041 & pi081;
assign w2449 = ~pi016 & ~pi045;
assign w2450 = ~w2448 & ~w2449;
assign w2451 = pi041 & ~pi081;
assign w2452 = pi016 & ~pi120;
assign w2453 = ~w2451 & w2452;
assign w2454 = ~w2447 & ~w2450;
assign w2455 = pi041 & ~pi045;
assign w2456 = ~pi120 & ~w2455;
assign w2457 = pi041 & pi081;
assign w2458 = ~pi120 & w2457;
assign w2459 = ~pi041 & pi045;
assign w2460 = ~pi016 & ~pi074;
assign w2461 = w2459 & w2460;
assign w2462 = ~w2458 & ~w2461;
assign w2463 = ~w2456 & ~w2462;
assign w2464 = ~pi016 & pi074;
assign w2465 = pi041 & w2464;
assign w2466 = w2464 & w2451;
assign w2467 = ~pi074 & ~pi120;
assign w2468 = w2447 & w2467;
assign w2469 = pi016 & ~pi074;
assign w2470 = w2447 & w2469;
assign w2471 = ~w2468 & ~w2470;
assign w2472 = ~w2466 & w2471;
assign w2473 = ~w2463 & w2472;
assign w2474 = (~pi003 & ~w2473) | (~pi003 & w18176) | (~w2473 & w18176);
assign w2475 = ~pi016 & pi081;
assign w2476 = pi016 & pi074;
assign w2477 = w2447 & w2476;
assign w2478 = ~pi045 & ~pi081;
assign w2479 = ~pi074 & w2478;
assign w2480 = ~pi041 & ~pi081;
assign w2481 = pi016 & w2480;
assign w2482 = ~w2477 & ~w2479;
assign w2483 = ~w2475 & ~w2481;
assign w2484 = w2482 & w2483;
assign w2485 = pi045 & w2476;
assign w2486 = w2448 & w2485;
assign w2487 = w2459 & w2467;
assign w2488 = ~pi081 & w2487;
assign w2489 = ~w2486 & ~w2488;
assign w2490 = pi120 & ~w2484;
assign w2491 = (pi003 & w2490) | (pi003 & w18177) | (w2490 & w18177);
assign w2492 = pi045 & w2460;
assign w2493 = w2460 & w2519;
assign w2494 = pi016 & w2447;
assign w2495 = w2447 & w18178;
assign w2496 = w2451 & w2469;
assign w2497 = ~w2493 & ~w2495;
assign w2498 = (pi120 & ~w2497) | (pi120 & w18179) | (~w2497 & w18179);
assign w2499 = pi074 & pi120;
assign w2500 = ~pi016 & w2448;
assign w2501 = w2455 & w2469;
assign w2502 = pi044 & ~w2501;
assign w2503 = w2499 & w2500;
assign w2504 = w2502 & ~w2503;
assign w2505 = pi016 & w2468;
assign w2506 = w2504 & ~w2505;
assign w2507 = ~w2474 & ~w2491;
assign w2508 = ~w2498 & w2506;
assign w2509 = w2507 & w2508;
assign w2510 = w2448 & w2469;
assign w2511 = ~pi045 & pi074;
assign w2512 = w2448 & w2511;
assign w2513 = ~pi081 & w2476;
assign w2514 = pi120 & ~w2510;
assign w2515 = ~w2512 & ~w2513;
assign w2516 = ~pi120 & w2515;
assign w2517 = ~w2514 & ~w2516;
assign w2518 = pi016 & ~pi041;
assign w2519 = pi045 & pi081;
assign w2520 = w2518 & w2519;
assign w2521 = ~pi074 & w2520;
assign w2522 = pi045 & ~pi081;
assign w2523 = pi074 & w2522;
assign w2524 = w2522 & w18180;
assign w2525 = (pi003 & w2517) | (pi003 & w18181) | (w2517 & w18181);
assign w2526 = pi041 & w2519;
assign w2527 = ~pi016 & w2455;
assign w2528 = ~w2526 & ~w2527;
assign w2529 = w2467 & ~w2528;
assign w2530 = ~pi016 & pi045;
assign w2531 = ~pi120 & w2530;
assign w2532 = pi041 & pi045;
assign w2533 = w2464 & w2532;
assign w2534 = ~w2531 & ~w2533;
assign w2535 = ~pi003 & ~w2534;
assign w2536 = ~pi041 & w2478;
assign w2537 = w2478 & w18182;
assign w2538 = pi016 & w2459;
assign w2539 = w2499 & w2538;
assign w2540 = w2478 & w2518;
assign w2541 = w2457 & w2476;
assign w2542 = ~pi045 & w2541;
assign w2543 = (~pi120 & w2542) | (~pi120 & w18183) | (w2542 & w18183);
assign w2544 = w2519 & w18178;
assign w2545 = pi016 & ~pi081;
assign w2546 = w2455 & w2545;
assign w2547 = w2449 & w2480;
assign w2548 = ~w2546 & ~w2547;
assign w2549 = (w2499 & ~w2548) | (w2499 & w20764) | (~w2548 & w20764);
assign w2550 = ~w2543 & ~w2549;
assign w2551 = (~pi003 & w2539) | (~pi003 & w18184) | (w2539 & w18184);
assign w2552 = w2550 & ~w2551;
assign w2553 = ~w2529 & ~w2535;
assign w2554 = ~pi044 & w2553;
assign w2555 = w2552 & w18185;
assign w2556 = ~w2509 & ~w2555;
assign w2557 = ~pi016 & w2519;
assign w2558 = w2449 & w2451;
assign w2559 = w2518 & w2522;
assign w2560 = ~w2557 & ~w2558;
assign w2561 = ~pi074 & ~w2559;
assign w2562 = w2560 & w2561;
assign w2563 = pi074 & pi081;
assign w2564 = w2455 & w2563;
assign w2565 = w2448 & w2530;
assign w2566 = ~w2564 & ~w2565;
assign w2567 = (w2566 & w2562) | (w2566 & w18186) | (w2562 & w18186);
assign w2568 = ~pi041 & ~pi045;
assign w2569 = w2475 & w2568;
assign w2570 = w2457 & w2530;
assign w2571 = ~w2569 & ~w2570;
assign w2572 = w2451 & ~w2530;
assign w2573 = (pi074 & ~w2571) | (pi074 & w18187) | (~w2571 & w18187);
assign w2574 = ~pi120 & ~w2573;
assign w2575 = ~w2567 & ~w2574;
assign w2576 = pi003 & w2575;
assign w2577 = w2449 & w2457;
assign w2578 = ~pi074 & w2577;
assign w2579 = w2511 & w2518;
assign w2580 = ~pi081 & w2579;
assign w2581 = ~w2578 & ~w2580;
assign w2582 = ~pi120 & ~w2581;
assign w2583 = w2457 & w2469;
assign w2584 = w2480 & w2511;
assign w2585 = ~w2583 & ~w2584;
assign w2586 = ~w2486 & w2585;
assign w2587 = pi120 & ~w2586;
assign w2588 = w2469 & w2532;
assign w2589 = w2459 & w2464;
assign w2590 = ~pi120 & w2589;
assign w2591 = ~w2588 & ~w2590;
assign w2592 = ~w2529 & w2591;
assign w2593 = ~w2587 & w2592;
assign w2594 = (~w2582 & w2593) | (~w2582 & w18188) | (w2593 & w18188);
assign w2595 = ~w2576 & w2594;
assign w2596 = ~w2556 & w2595;
assign w2597 = pi062 & pi101;
assign w2598 = pi103 & w2597;
assign w2599 = pi062 & ~pi119;
assign w2600 = pi103 & w2599;
assign w2601 = ~pi062 & ~pi101;
assign w2602 = pi103 & w2601;
assign w2603 = ~w2598 & ~w2600;
assign w2604 = (~pi118 & ~w2603) | (~pi118 & w18189) | (~w2603 & w18189);
assign w2605 = pi066 & ~pi101;
assign w2606 = w2599 & w2605;
assign w2607 = ~pi118 & ~w2606;
assign w2608 = ~w2606 & w18190;
assign w2609 = ~pi066 & pi118;
assign w2610 = w2600 & w2609;
assign w2611 = ~pi062 & pi101;
assign w2612 = pi066 & ~pi103;
assign w2613 = ~pi066 & pi119;
assign w2614 = ~pi101 & ~pi103;
assign w2615 = w2613 & w2614;
assign w2616 = w2611 & w2612;
assign w2617 = pi118 & w2615;
assign w2618 = ~w2616 & ~w2617;
assign w2619 = ~w2608 & w2618;
assign w2620 = w2619 & w18191;
assign w2621 = ~pi034 & ~w2620;
assign w2622 = pi062 & ~pi103;
assign w2623 = ~w2602 & ~w2622;
assign w2624 = pi066 & w2599;
assign w2625 = ~pi062 & ~pi119;
assign w2626 = ~pi066 & w2625;
assign w2627 = ~pi103 & w2613;
assign w2628 = w2613 & w2622;
assign w2629 = ~pi034 & ~w2628;
assign w2630 = ~w2624 & ~w2626;
assign w2631 = w2623 & w2630;
assign w2632 = ~pi066 & pi103;
assign w2633 = w2611 & w2632;
assign w2634 = pi103 & ~pi119;
assign w2635 = w2597 & w2634;
assign w2636 = ~w2633 & ~w2635;
assign w2637 = (w2636 & w2631) | (w2636 & w18192) | (w2631 & w18192);
assign w2638 = pi118 & ~w2637;
assign w2639 = pi062 & pi119;
assign w2640 = ~pi101 & pi103;
assign w2641 = w2639 & w2640;
assign w2642 = pi066 & w2641;
assign w2643 = ~pi066 & ~pi118;
assign w2644 = ~pi101 & pi119;
assign w2645 = w2643 & w2644;
assign w2646 = ~pi062 & w2645;
assign w2647 = ~w2642 & ~w2646;
assign w2648 = pi066 & pi118;
assign w2649 = pi062 & ~pi101;
assign w2650 = ~pi103 & w2649;
assign w2651 = w2648 & w2650;
assign w2652 = w2600 & w2643;
assign w2653 = pi101 & ~pi119;
assign w2654 = w2632 & w2653;
assign w2655 = ~w2651 & ~w2652;
assign w2656 = pi038 & ~w2654;
assign w2657 = w2655 & w2656;
assign w2658 = pi034 & ~w2647;
assign w2659 = w2657 & ~w2658;
assign w2660 = pi066 & pi103;
assign w2661 = ~pi062 & w2660;
assign w2662 = ~w2606 & ~w2661;
assign w2663 = ~pi118 & ~w2662;
assign w2664 = pi062 & w2640;
assign w2665 = w2613 & w2664;
assign w2666 = w2599 & w2640;
assign w2667 = w2609 & w2666;
assign w2668 = pi066 & pi101;
assign w2669 = ~pi062 & pi119;
assign w2670 = w2668 & w2669;
assign w2671 = ~w2665 & ~w2667;
assign w2672 = ~w2663 & w2671;
assign w2673 = pi101 & w2599;
assign w2674 = w2660 & w2673;
assign w2675 = w2597 & w2613;
assign w2676 = ~pi066 & pi101;
assign w2677 = ~pi103 & ~pi119;
assign w2678 = w2676 & w2677;
assign w2679 = ~w2675 & ~w2678;
assign w2680 = w2625 & w2640;
assign w2681 = ~w2674 & w2679;
assign w2682 = (~pi118 & ~w2681) | (~pi118 & w18193) | (~w2681 & w18193);
assign w2683 = pi103 & w2644;
assign w2684 = w2648 & w2683;
assign w2685 = ~pi103 & pi119;
assign w2686 = pi118 & ~w2668;
assign w2687 = w2685 & ~w2686;
assign w2688 = pi118 & ~pi119;
assign w2689 = w2601 & w2688;
assign w2690 = ~w2684 & ~w2687;
assign w2691 = (~pi034 & ~w2690) | (~pi034 & w18194) | (~w2690 & w18194);
assign w2692 = pi101 & pi103;
assign w2693 = w2625 & w2692;
assign w2694 = w2639 & w2692;
assign w2695 = ~w2693 & ~w2694;
assign w2696 = w2648 & ~w2695;
assign w2697 = ~pi103 & w2601;
assign w2698 = ~pi119 & w2648;
assign w2699 = w2697 & w2698;
assign w2700 = ~pi038 & ~w2699;
assign w2701 = ~w2696 & w2700;
assign w2702 = ~w2691 & w2701;
assign w2703 = ~w2682 & w2702;
assign w2704 = (pi034 & ~w2672) | (pi034 & w18195) | (~w2672 & w18195);
assign w2705 = w2703 & ~w2704;
assign w2706 = ~w2638 & w2659;
assign w2707 = ~w2621 & w2706;
assign w2708 = ~w2705 & ~w2707;
assign w2709 = ~w2625 & ~w2660;
assign w2710 = w2692 & w2709;
assign w2711 = w2605 & w2625;
assign w2712 = ~w2642 & ~w2710;
assign w2713 = pi101 & pi119;
assign w2714 = w2632 & w2713;
assign w2715 = ~pi118 & ~w2714;
assign w2716 = w2612 & w2644;
assign w2717 = w2679 & w2715;
assign w2718 = (~pi034 & ~w2717) | (~pi034 & w18196) | (~w2717 & w18196);
assign w2719 = ~pi101 & ~pi119;
assign w2720 = w2660 & w2719;
assign w2721 = ~pi066 & ~pi103;
assign w2722 = w2597 & w2721;
assign w2723 = ~pi119 & w2722;
assign w2724 = ~pi062 & w2720;
assign w2725 = ~w2723 & ~w2724;
assign w2726 = (w2712 & w3181) | (w2712 & w18197) | (w3181 & w18197);
assign w2727 = ~w2718 & w2725;
assign w2728 = ~w2726 & ~w2727;
assign w2729 = w2597 & w2688;
assign w2730 = w2599 & w2614;
assign w2731 = w2622 & w2713;
assign w2732 = ~w2730 & ~w2731;
assign w2733 = w2611 & ~w2685;
assign w2734 = (~pi118 & ~w2732) | (~pi118 & w18198) | (~w2732 & w18198);
assign w2735 = ~w2729 & ~w2734;
assign w2736 = w2649 & w2685;
assign w2737 = ~w2613 & ~w2736;
assign w2738 = ~w2623 & ~w2737;
assign w2739 = ~pi103 & w2625;
assign w2740 = w2676 & w2739;
assign w2741 = pi066 & ~w2735;
assign w2742 = (pi034 & w2741) | (pi034 & w18200) | (w2741 & w18200);
assign w2743 = ~w2728 & ~w2742;
assign w2744 = ~w2708 & w2743;
assign w2745 = ~w2596 & w2744;
assign w2746 = w2596 & ~w2744;
assign w2747 = ~w2745 & ~w2746;
assign w2748 = ~pi041 & ~pi074;
assign w2749 = w2478 & w2748;
assign w2750 = ~w2520 & ~w2749;
assign w2751 = (pi120 & ~w2750) | (pi120 & w18201) | (~w2750 & w18201);
assign w2752 = pi041 & ~w2522;
assign w2753 = w2455 & w2460;
assign w2754 = w2467 & w2559;
assign w2755 = ~w2753 & ~w2754;
assign w2756 = w2464 & ~w2752;
assign w2757 = w2755 & ~w2756;
assign w2758 = (~pi003 & ~w2757) | (~pi003 & w18202) | (~w2757 & w18202);
assign w2759 = pi074 & ~w2450;
assign w2760 = ~w2544 & ~w2759;
assign w2761 = (~pi120 & ~w2760) | (~pi120 & w18203) | (~w2760 & w18203);
assign w2762 = w2455 & w2476;
assign w2763 = ~pi081 & w2762;
assign w2764 = pi045 & w2496;
assign w2765 = ~w2763 & ~w2764;
assign w2766 = ~pi016 & w2480;
assign w2767 = ~w2465 & ~w2766;
assign w2768 = pi045 & ~w2767;
assign w2769 = w2765 & ~w2768;
assign w2770 = ~pi041 & ~pi120;
assign w2771 = w2478 & w2770;
assign w2772 = w2447 & w2518;
assign w2773 = ~w2458 & ~w2771;
assign w2774 = (pi003 & ~w2773) | (pi003 & w18204) | (~w2773 & w18204);
assign w2775 = pi041 & w2447;
assign w2776 = w2447 & w18205;
assign w2777 = ~pi081 & w2464;
assign w2778 = w2459 & w2777;
assign w2779 = ~w2776 & ~w2778;
assign w2780 = ~w2774 & w2779;
assign w2781 = pi120 & ~w2769;
assign w2782 = w2780 & ~w2781;
assign w2783 = w2782 & w18206;
assign w2784 = pi044 & ~w2783;
assign w2785 = ~w2478 & ~w2485;
assign w2786 = ~w2513 & ~w2785;
assign w2787 = w2499 & w2775;
assign w2788 = ~w2487 & ~w2787;
assign w2789 = ~w2786 & w2788;
assign w2790 = pi003 & ~w2789;
assign w2791 = w2476 & w2478;
assign w2792 = ~pi120 & w2791;
assign w2793 = ~pi074 & ~w2571;
assign w2794 = (~pi003 & w2793) | (~pi003 & w18207) | (w2793 & w18207);
assign w2795 = w2460 & w2480;
assign w2796 = pi045 & pi074;
assign w2797 = w2457 & w2796;
assign w2798 = ~w2795 & ~w2797;
assign w2799 = ~w2764 & w2798;
assign w2800 = ~pi120 & ~w2799;
assign w2801 = ~pi016 & w2499;
assign w2802 = pi041 & w2478;
assign w2803 = ~w2448 & ~w2802;
assign w2804 = w2801 & ~w2803;
assign w2805 = ~pi003 & pi120;
assign w2806 = w2532 & ~w2563;
assign w2807 = w2805 & w2806;
assign w2808 = ~w2804 & ~w2807;
assign w2809 = ~w2790 & ~w2794;
assign w2810 = ~w2800 & w2808;
assign w2811 = w2451 & w2460;
assign w2812 = ~pi045 & w2811;
assign w2813 = ~pi074 & w2569;
assign w2814 = ~w2812 & ~w2813;
assign w2815 = (~pi120 & ~w2814) | (~pi120 & w18208) | (~w2814 & w18208);
assign w2816 = w2457 & w2460;
assign w2817 = pi045 & w2795;
assign w2818 = (pi120 & w2817) | (pi120 & w18209) | (w2817 & w18209);
assign w2819 = w2447 & w2464;
assign w2820 = w2458 & w2819;
assign w2821 = pi041 & pi120;
assign w2822 = w2513 & w2821;
assign w2823 = w2513 & w18210;
assign w2824 = ~w2820 & ~w2823;
assign w2825 = ~w2818 & w2824;
assign w2826 = ~w2815 & w2825;
assign w2827 = w2476 & w18211;
assign w2828 = ~pi074 & pi120;
assign w2829 = w2527 & w2828;
assign w2830 = ~w2827 & ~w2829;
assign w2831 = ~pi041 & w2447;
assign w2832 = pi120 & w2469;
assign w2833 = w2831 & w2832;
assign w2834 = ~pi074 & w2547;
assign w2835 = ~pi041 & w2522;
assign w2836 = w2499 & w2835;
assign w2837 = w2465 & w2478;
assign w2838 = ~w2836 & ~w2837;
assign w2839 = ~pi120 & w2588;
assign w2840 = w2838 & ~w2839;
assign w2841 = ~w2833 & ~w2834;
assign w2842 = (pi003 & ~w2840) | (pi003 & w18212) | (~w2840 & w18212);
assign w2843 = pi081 & ~w2830;
assign w2844 = ~w2842 & ~w2843;
assign w2845 = ~pi003 & ~w2826;
assign w2846 = w2844 & ~w2845;
assign w2847 = (~pi044 & ~w2809) | (~pi044 & w18213) | (~w2809 & w18213);
assign w2848 = w2846 & ~w2847;
assign w2849 = ~w2784 & w2848;
assign w2850 = w2625 & w18214;
assign w2851 = ~w2635 & ~w2641;
assign w2852 = (pi118 & ~w2851) | (pi118 & w18215) | (~w2851 & w18215);
assign w2853 = ~pi118 & pi119;
assign w2854 = w2601 & w2632;
assign w2855 = pi066 & w2614;
assign w2856 = w2612 & w2669;
assign w2857 = ~w2678 & ~w2855;
assign w2858 = ~w2856 & w2857;
assign w2859 = w2853 & w2854;
assign w2860 = w2858 & ~w2859;
assign w2861 = (~pi034 & ~w2860) | (~pi034 & w18216) | (~w2860 & w18216);
assign w2862 = w2612 & w2713;
assign w2863 = pi066 & w2693;
assign w2864 = ~w2862 & ~w2863;
assign w2865 = w2669 & w2692;
assign w2866 = ~pi066 & w2865;
assign w2867 = w2614 & w2669;
assign w2868 = ~w2866 & ~w2867;
assign w2869 = w2864 & w2868;
assign w2870 = pi118 & ~w2869;
assign w2871 = ~w2649 & ~w2677;
assign w2872 = pi066 & ~w2871;
assign w2873 = ~w2654 & ~w2694;
assign w2874 = ~w2872 & w2873;
assign w2875 = ~pi118 & ~w2874;
assign w2876 = ~pi101 & ~pi118;
assign w2877 = w2625 & w2876;
assign w2878 = ~pi118 & w2597;
assign w2879 = ~w2666 & ~w2878;
assign w2880 = (pi034 & ~w2879) | (pi034 & w18217) | (~w2879 & w18217);
assign w2881 = w2599 & w2676;
assign w2882 = ~pi103 & w2669;
assign w2883 = w2605 & w2882;
assign w2884 = ~w2881 & ~w2883;
assign w2885 = ~w2875 & ~w2880;
assign w2886 = ~w2870 & w2885;
assign w2887 = w2886 & w18218;
assign w2888 = pi038 & ~w2887;
assign w2889 = pi066 & w2639;
assign w2890 = w2639 & w2668;
assign w2891 = ~w2866 & ~w2890;
assign w2892 = w2601 & w2721;
assign w2893 = ~w2866 & w18219;
assign w2894 = ~pi118 & ~w2893;
assign w2895 = ~pi034 & pi118;
assign w2896 = pi119 & w2611;
assign w2897 = ~w2675 & ~w2896;
assign w2898 = w2895 & ~w2897;
assign w2899 = w2668 & w2739;
assign w2900 = w2739 & w18220;
assign w2901 = ~w2651 & ~w2900;
assign w2902 = w2625 & w2660;
assign w2903 = ~pi118 & w2902;
assign w2904 = ~pi066 & ~w2732;
assign w2905 = ~w2639 & w2660;
assign w2906 = ~w2709 & ~w2905;
assign w2907 = ~w2645 & ~w2906;
assign w2908 = w2597 & w2698;
assign w2909 = ~w2904 & w18221;
assign w2910 = w2907 & w20765;
assign w2911 = ~w2909 & ~w2910;
assign w2912 = ~w2898 & w2901;
assign w2913 = ~w2894 & w2912;
assign w2914 = w2613 & w2697;
assign w2915 = pi118 & ~w2722;
assign w2916 = ~w2863 & ~w2914;
assign w2917 = w2915 & w2916;
assign w2918 = pi101 & w2612;
assign w2919 = w2599 & w2918;
assign w2920 = (~pi118 & ~w2918) | (~pi118 & w18222) | (~w2918 & w18222);
assign w2921 = ~pi066 & w2599;
assign w2922 = pi101 & ~pi103;
assign w2923 = w2921 & ~w2922;
assign w2924 = ~w2740 & ~w2923;
assign w2925 = (~pi034 & ~w2924) | (~pi034 & w18223) | (~w2924 & w18223);
assign w2926 = ~pi103 & w2653;
assign w2927 = w2660 & w2853;
assign w2928 = w2609 & w2926;
assign w2929 = ~pi103 & w2850;
assign w2930 = w2605 & w2669;
assign w2931 = pi118 & ~w2930;
assign w2932 = ~w2715 & ~w2931;
assign w2933 = ~w2667 & ~w2899;
assign w2934 = ~w2929 & w2933;
assign w2935 = ~w2932 & w2934;
assign w2936 = (pi062 & w2928) | (pi062 & w18224) | (w2928 & w18224);
assign w2937 = (~w2936 & w2935) | (~w2936 & w18225) | (w2935 & w18225);
assign w2938 = ~w2917 & w2925;
assign w2939 = w2937 & ~w2938;
assign w2940 = (~pi038 & w2911) | (~pi038 & w18226) | (w2911 & w18226);
assign w2941 = w2939 & ~w2940;
assign w2942 = ~w2888 & w2941;
assign w2943 = ~w2849 & w2942;
assign w2944 = w2849 & ~w2942;
assign w2945 = ~w2943 & ~w2944;
assign w2946 = w2747 & ~w2945;
assign w2947 = ~w2747 & w2945;
assign w2948 = ~w2946 & ~w2947;
assign w2949 = ~pi022 & pi057;
assign w2950 = pi000 & ~pi097;
assign w2951 = w2949 & w2950;
assign w2952 = ~pi022 & pi097;
assign w2953 = ~pi000 & pi057;
assign w2954 = w2952 & w2953;
assign w2955 = ~pi011 & w2954;
assign w2956 = (~pi116 & w2955) | (~pi116 & w18227) | (w2955 & w18227);
assign w2957 = pi022 & pi097;
assign w2958 = ~pi000 & pi011;
assign w2959 = w2957 & w2958;
assign w2960 = pi057 & w2959;
assign w2961 = pi000 & ~pi022;
assign w2962 = pi057 & ~pi097;
assign w2963 = pi011 & w2962;
assign w2964 = w2961 & w2963;
assign w2965 = ~pi011 & pi116;
assign w2966 = pi022 & w2962;
assign w2967 = w2965 & w2966;
assign w2968 = pi011 & ~pi022;
assign w2969 = pi057 & pi097;
assign w2970 = w2968 & w2969;
assign w2971 = pi116 & w2970;
assign w2972 = ~w2960 & ~w2964;
assign w2973 = ~w2967 & ~w2971;
assign w2974 = w2972 & w2973;
assign w2975 = (~pi058 & ~w2974) | (~pi058 & w18228) | (~w2974 & w18228);
assign w2976 = pi057 & w2957;
assign w2977 = w2957 & w18229;
assign w2978 = pi000 & pi022;
assign w2979 = (pi116 & ~w2978) | (pi116 & w18230) | (~w2978 & w18230);
assign w2980 = ~pi022 & ~pi057;
assign w2981 = ~pi000 & w2980;
assign w2982 = ~pi057 & pi097;
assign w2983 = ~pi011 & w2982;
assign w2984 = pi000 & pi011;
assign w2985 = w2949 & w2984;
assign w2986 = ~w2983 & ~w2985;
assign w2987 = (~pi116 & ~w2980) | (~pi116 & w18231) | (~w2980 & w18231);
assign w2988 = w2986 & w2987;
assign w2989 = ~w2977 & w2979;
assign w2990 = ~w2988 & ~w2989;
assign w2991 = ~w2961 & w2963;
assign w2992 = ~pi057 & ~pi097;
assign w2993 = w2968 & w2992;
assign w2994 = (pi058 & w2990) | (pi058 & w18232) | (w2990 & w18232);
assign w2995 = pi000 & ~pi011;
assign w2996 = w2957 & w2995;
assign w2997 = ~pi057 & w2996;
assign w2998 = ~w2960 & ~w2997;
assign w2999 = ~pi116 & ~w2998;
assign w3000 = ~pi000 & ~pi097;
assign w3001 = ~pi022 & w2992;
assign w3002 = (w2965 & w3001) | (w2965 & w18233) | (w3001 & w18233);
assign w3003 = pi022 & pi116;
assign w3004 = w2984 & w2992;
assign w3005 = w3003 & w3004;
assign w3006 = ~pi000 & ~pi011;
assign w3007 = w2992 & w3006;
assign w3008 = ~w3005 & ~w3007;
assign w3009 = ~w3002 & w3008;
assign w3010 = ~w2999 & w3009;
assign w3011 = ~w2975 & ~w2994;
assign w3012 = (~pi060 & ~w3011) | (~pi060 & w18234) | (~w3011 & w18234);
assign w3013 = w2976 & w2984;
assign w3014 = ~w2954 & ~w3013;
assign w3015 = pi000 & w2949;
assign w3016 = ~pi000 & w2952;
assign w3017 = pi011 & w2969;
assign w3018 = ~w3015 & ~w3016;
assign w3019 = (pi116 & ~w3018) | (pi116 & w18235) | (~w3018 & w18235);
assign w3020 = w3014 & ~w3019;
assign w3021 = pi022 & w2982;
assign w3022 = w3006 & w3021;
assign w3023 = ~pi022 & ~pi097;
assign w3024 = ~w2969 & w2984;
assign w3025 = ~w3023 & w3024;
assign w3026 = w2953 & w3023;
assign w3027 = pi011 & ~pi116;
assign w3028 = w2982 & w3027;
assign w3029 = ~w3022 & ~w3025;
assign w3030 = ~w3026 & ~w3028;
assign w3031 = ~pi011 & pi022;
assign w3032 = w2962 & w3031;
assign w3033 = pi011 & pi022;
assign w3034 = w2982 & w3033;
assign w3035 = w2978 & w2992;
assign w3036 = ~w3026 & ~w3032;
assign w3037 = ~w3034 & ~w3035;
assign w3038 = w3036 & w3037;
assign w3039 = ~pi011 & ~pi022;
assign w3040 = w2969 & w3039;
assign w3041 = ~pi000 & ~pi116;
assign w3042 = pi022 & ~pi057;
assign w3043 = w2995 & w3042;
assign w3044 = w3040 & ~w3041;
assign w3045 = ~pi097 & w3043;
assign w3046 = ~w3044 & ~w3045;
assign w3047 = ~pi116 & ~w3038;
assign w3048 = w3046 & ~w3047;
assign w3049 = (~pi058 & ~w3029) | (~pi058 & w18236) | (~w3029 & w18236);
assign w3050 = w3048 & ~w3049;
assign w3051 = (pi060 & ~w3050) | (pi060 & w18237) | (~w3050 & w18237);
assign w3052 = ~pi097 & w2995;
assign w3053 = w2980 & w3052;
assign w3054 = w2962 & w2968;
assign w3055 = ~w2959 & ~w3054;
assign w3056 = ~w3053 & w3055;
assign w3057 = ~pi116 & ~w3056;
assign w3058 = pi022 & w2992;
assign w3059 = w2984 & w3058;
assign w3060 = pi011 & ~pi057;
assign w3061 = pi000 & w3060;
assign w3062 = w2952 & w3061;
assign w3063 = ~w3059 & ~w3062;
assign w3064 = (~pi058 & w3057) | (~pi058 & w18238) | (w3057 & w18238);
assign w3065 = pi058 & ~pi116;
assign w3066 = pi022 & ~pi097;
assign w3067 = w2953 & w3066;
assign w3068 = w2992 & w3031;
assign w3069 = ~w2993 & ~w3067;
assign w3070 = ~w3068 & w3069;
assign w3071 = w2980 & w3000;
assign w3072 = ~w3022 & ~w3071;
assign w3073 = w3070 & w3072;
assign w3074 = w3065 & ~w3073;
assign w3075 = pi058 & pi116;
assign w3076 = pi022 & pi057;
assign w3077 = pi000 & w3076;
assign w3078 = ~w2954 & ~w3077;
assign w3079 = pi011 & ~w3078;
assign w3080 = pi000 & pi057;
assign w3081 = w2952 & w3080;
assign w3082 = (w3075 & w3079) | (w3075 & w18239) | (w3079 & w18239);
assign w3083 = ~pi058 & pi116;
assign w3084 = pi057 & w2995;
assign w3085 = w2957 & w3084;
assign w3086 = w2982 & w3039;
assign w3087 = ~w3007 & ~w3086;
assign w3088 = ~w3085 & w3087;
assign w3089 = w3083 & ~w3088;
assign w3090 = pi011 & pi116;
assign w3091 = ~pi000 & w3023;
assign w3092 = w3090 & w3091;
assign w3093 = w3091 & w18240;
assign w3094 = pi000 & pi116;
assign w3095 = w2968 & w2982;
assign w3096 = w3094 & w3095;
assign w3097 = ~w3093 & ~w3096;
assign w3098 = ~w3074 & ~w3082;
assign w3099 = ~w3089 & w3097;
assign w3100 = w3098 & w18241;
assign w3101 = ~w3051 & w3100;
assign w3102 = ~w3012 & w3101;
assign w3103 = ~pi066 & w2669;
assign w3104 = ~pi101 & ~w2622;
assign w3105 = pi062 & w2632;
assign w3106 = ~w2602 & ~w3105;
assign w3107 = (~w3103 & ~w3106) | (~w3103 & w18242) | (~w3106 & w18242);
assign w3108 = pi119 & w2692;
assign w3109 = ~w2675 & ~w3108;
assign w3110 = w2624 & ~w2640;
assign w3111 = ~w2711 & ~w3110;
assign w3112 = pi118 & ~w3109;
assign w3113 = w3111 & ~w3112;
assign w3114 = ~pi118 & ~w3107;
assign w3115 = w3113 & ~w3114;
assign w3116 = w2627 & w2649;
assign w3117 = (~pi118 & w3116) | (~pi118 & w18243) | (w3116 & w18243);
assign w3118 = w2605 & w2639;
assign w3119 = ~w2881 & ~w3118;
assign w3120 = pi118 & ~w3119;
assign w3121 = w2597 & w2612;
assign w3122 = pi119 & w3121;
assign w3123 = pi103 & w2606;
assign w3124 = ~w3122 & ~w3123;
assign w3125 = ~w3120 & w3124;
assign w3126 = ~w2866 & ~w3122;
assign w3127 = ~pi118 & ~w3126;
assign w3128 = w2648 & w2693;
assign w3129 = ~w2677 & ~w2689;
assign w3130 = w2599 & w2643;
assign w3131 = ~pi066 & ~w3130;
assign w3132 = ~w3129 & w3131;
assign w3133 = ~w3128 & ~w3132;
assign w3134 = ~w3127 & w3133;
assign w3135 = (~pi034 & ~w3125) | (~pi034 & w18244) | (~w3125 & w18244);
assign w3136 = w3134 & ~w3135;
assign w3137 = pi034 & ~w3115;
assign w3138 = w3136 & ~w3137;
assign w3139 = pi101 & w2639;
assign w3140 = w2660 & w3139;
assign w3141 = ~w2736 & ~w3140;
assign w3142 = ~w2664 & ~w2889;
assign w3143 = (pi118 & ~w3142) | (pi118 & w18245) | (~w3142 & w18245);
assign w3144 = w3141 & ~w3143;
assign w3145 = w2611 & w2627;
assign w3146 = ~w2719 & w2905;
assign w3147 = pi066 & ~pi118;
assign w3148 = w2669 & w3147;
assign w3149 = ~w3145 & ~w3146;
assign w3150 = ~w2730 & ~w3148;
assign w3151 = ~w2670 & ~w2693;
assign w3152 = ~w2730 & ~w2881;
assign w3153 = w3151 & w3152;
assign w3154 = w2613 & w2649;
assign w3155 = ~pi118 & ~w2640;
assign w3156 = ~pi066 & w2693;
assign w3157 = w3154 & ~w3155;
assign w3158 = ~w3156 & ~w3157;
assign w3159 = ~pi118 & ~w3153;
assign w3160 = w3158 & ~w3159;
assign w3161 = (~pi034 & ~w3149) | (~pi034 & w18246) | (~w3149 & w18246);
assign w3162 = w3160 & ~w3161;
assign w3163 = (pi038 & ~w3162) | (pi038 & w18247) | (~w3162 & w18247);
assign w3164 = w2626 & w2640;
assign w3165 = ~w2606 & ~w2862;
assign w3166 = ~w3164 & w3165;
assign w3167 = ~pi118 & ~w3166;
assign w3168 = pi066 & w2669;
assign w3169 = w2640 & w3168;
assign w3170 = ~w2863 & ~w3169;
assign w3171 = (~pi034 & w3167) | (~pi034 & w18248) | (w3167 & w18248);
assign w3172 = pi034 & ~pi118;
assign w3173 = w2599 & w2922;
assign w3174 = w2614 & w2625;
assign w3175 = ~w2711 & ~w3173;
assign w3176 = ~w3174 & w3175;
assign w3177 = w2625 & w2676;
assign w3178 = ~w3145 & ~w3177;
assign w3179 = w3176 & w3178;
assign w3180 = w3172 & ~w3179;
assign w3181 = pi034 & pi118;
assign w3182 = ~w2598 & ~w2736;
assign w3183 = pi066 & ~w3182;
assign w3184 = (w3181 & w3183) | (w3181 & w18249) | (w3183 & w18249);
assign w3185 = w2713 & w3105;
assign w3186 = w2625 & w2721;
assign w3187 = w2601 & w2613;
assign w3188 = ~w3186 & ~w3187;
assign w3189 = ~w3185 & w3188;
assign w3190 = w2895 & ~w3189;
assign w3191 = pi103 & pi118;
assign w3192 = w2930 & w3191;
assign w3193 = ~w2699 & ~w3192;
assign w3194 = ~w3190 & w3193;
assign w3195 = ~w3184 & w3194;
assign w3196 = w3195 & w18250;
assign w3197 = ~w3163 & w3196;
assign w3198 = ~pi038 & ~w3138;
assign w3199 = w3197 & ~w3198;
assign w3200 = ~w3102 & w3199;
assign w3201 = w3102 & ~w3199;
assign w3202 = ~w3200 & ~w3201;
assign w3203 = ~pi051 & pi112;
assign w3204 = pi049 & ~pi086;
assign w3205 = w3203 & w3204;
assign w3206 = ~pi049 & pi112;
assign w3207 = pi051 & ~pi086;
assign w3208 = w3206 & w3207;
assign w3209 = ~pi019 & w3208;
assign w3210 = (~pi090 & w3209) | (~pi090 & w18251) | (w3209 & w18251);
assign w3211 = ~pi051 & w3204;
assign w3212 = w3204 & w18252;
assign w3213 = pi112 & w3212;
assign w3214 = pi019 & ~pi049;
assign w3215 = pi051 & pi112;
assign w3216 = pi086 & w3215;
assign w3217 = w3214 & w3216;
assign w3218 = ~pi019 & pi086;
assign w3219 = w3203 & w3218;
assign w3220 = pi019 & ~pi086;
assign w3221 = w3215 & w3220;
assign w3222 = ~w3219 & ~w3221;
assign w3223 = pi090 & ~w3222;
assign w3224 = ~w3213 & ~w3223;
assign w3225 = w3224 & w18253;
assign w3226 = pi051 & ~pi112;
assign w3227 = ~pi019 & w3226;
assign w3228 = pi019 & pi112;
assign w3229 = ~pi049 & ~pi086;
assign w3230 = ~w3228 & ~w3229;
assign w3231 = ~pi086 & ~w3206;
assign w3232 = ~w3230 & w3231;
assign w3233 = pi049 & pi051;
assign w3234 = pi086 & w3233;
assign w3235 = w3215 & w3218;
assign w3236 = ~w3234 & ~w3235;
assign w3237 = pi090 & ~w3236;
assign w3238 = ~pi051 & ~pi112;
assign w3239 = w3220 & w3238;
assign w3240 = pi019 & w3203;
assign w3241 = ~w3204 & w3240;
assign w3242 = ~w3239 & ~w3241;
assign w3243 = ~w3237 & w3242;
assign w3244 = pi019 & ~pi090;
assign w3245 = ~pi049 & pi051;
assign w3246 = pi086 & pi112;
assign w3247 = w3245 & w3246;
assign w3248 = ~pi019 & ~pi049;
assign w3249 = w3238 & w3248;
assign w3250 = ~pi019 & ~pi090;
assign w3251 = pi049 & pi086;
assign w3252 = w3226 & w3251;
assign w3253 = w3250 & w3252;
assign w3254 = ~w3249 & ~w3253;
assign w3255 = w3244 & w3247;
assign w3256 = w3254 & ~w3255;
assign w3257 = ~pi051 & pi086;
assign w3258 = pi019 & pi049;
assign w3259 = ~pi112 & w3258;
assign w3260 = w3257 & w3259;
assign w3261 = w3259 & w18255;
assign w3262 = ~pi019 & pi090;
assign w3263 = ~pi086 & w3238;
assign w3264 = ~pi049 & ~pi051;
assign w3265 = (w3262 & w3263) | (w3262 & w18256) | (w3263 & w18256);
assign w3266 = ~w3261 & ~w3265;
assign w3267 = w3256 & w3266;
assign w3268 = (pi088 & ~w3243) | (pi088 & w18257) | (~w3243 & w18257);
assign w3269 = w3267 & ~w3268;
assign w3270 = ~pi088 & ~w3225;
assign w3271 = w3269 & ~w3270;
assign w3272 = pi086 & ~pi112;
assign w3273 = w3248 & w3272;
assign w3274 = (w3226 & w3273) | (w3226 & w18258) | (w3273 & w18258);
assign w3275 = w3203 & w3229;
assign w3276 = ~w3226 & ~w3257;
assign w3277 = w3258 & ~w3276;
assign w3278 = ~w3275 & ~w3277;
assign w3279 = (~pi088 & ~w3278) | (~pi088 & w18259) | (~w3278 & w18259);
assign w3280 = pi051 & pi086;
assign w3281 = w3228 & w3280;
assign w3282 = pi049 & w3281;
assign w3283 = ~w3208 & ~w3282;
assign w3284 = ~pi019 & ~pi086;
assign w3285 = w3215 & w3284;
assign w3286 = ~pi019 & pi049;
assign w3287 = pi112 & w3286;
assign w3288 = (~pi090 & ~w3286) | (~pi090 & w18260) | (~w3286 & w18260);
assign w3289 = w3272 & w3286;
assign w3290 = w3285 & ~w3288;
assign w3291 = ~pi051 & w3289;
assign w3292 = ~w3290 & ~w3291;
assign w3293 = (pi088 & w3282) | (pi088 & w18261) | (w3282 & w18261);
assign w3294 = w3292 & ~w3293;
assign w3295 = pi088 & pi090;
assign w3296 = ~pi086 & pi112;
assign w3297 = pi051 & ~w3230;
assign w3298 = pi049 & w3296;
assign w3299 = pi019 & ~pi112;
assign w3300 = w3280 & w3299;
assign w3301 = w3238 & w3251;
assign w3302 = ~w3219 & ~w3275;
assign w3303 = ~w3300 & ~w3301;
assign w3304 = w3302 & w3303;
assign w3305 = (w3295 & w3297) | (w3295 & w18262) | (w3297 & w18262);
assign w3306 = ~pi090 & ~w3304;
assign w3307 = ~w3305 & ~w3306;
assign w3308 = ~w3279 & w3294;
assign w3309 = w3307 & w3308;
assign w3310 = pi006 & ~w3309;
assign w3311 = w3263 & w3286;
assign w3312 = w3203 & w3220;
assign w3313 = w3214 & w3280;
assign w3314 = ~w3312 & ~w3313;
assign w3315 = ~w3311 & w3314;
assign w3316 = ~pi090 & ~w3315;
assign w3317 = pi019 & w3226;
assign w3318 = w3204 & w3317;
assign w3319 = ~w3260 & ~w3318;
assign w3320 = (~pi088 & w3316) | (~pi088 & w18263) | (w3316 & w18263);
assign w3321 = pi088 & ~pi090;
assign w3322 = w3246 & w3264;
assign w3323 = w3218 & w3238;
assign w3324 = w3229 & w3238;
assign w3325 = ~w3322 & ~w3323;
assign w3326 = ~w3324 & w3325;
assign w3327 = ~w3239 & ~w3273;
assign w3328 = (w3321 & ~w3326) | (w3321 & w18264) | (~w3326 & w18264);
assign w3329 = w3207 & w3287;
assign w3330 = pi049 & w3246;
assign w3331 = ~w3208 & ~w3330;
assign w3332 = pi019 & ~w3331;
assign w3333 = (w3295 & w3332) | (w3295 & w18265) | (w3332 & w18265);
assign w3334 = ~pi088 & pi090;
assign w3335 = w3280 & w3286;
assign w3336 = pi112 & w3335;
assign w3337 = w3226 & w3284;
assign w3338 = ~w3249 & ~w3337;
assign w3339 = ~w3336 & w3338;
assign w3340 = w3334 & ~w3339;
assign w3341 = pi090 & w3214;
assign w3342 = w3263 & w3341;
assign w3343 = w3220 & w3226;
assign w3344 = pi090 & w3343;
assign w3345 = w3343 & w6274;
assign w3346 = ~w3342 & ~w3345;
assign w3347 = ~w3328 & ~w3333;
assign w3348 = ~w3340 & w3346;
assign w3349 = w3347 & w3348;
assign w3350 = ~w3320 & w3349;
assign w3351 = ~w3310 & w3350;
assign w3352 = ~pi006 & ~w3271;
assign w3353 = w3351 & ~w3352;
assign w3354 = ~pi303 & w3353;
assign w3355 = pi303 & ~w3353;
assign w3356 = ~w3354 & ~w3355;
assign w3357 = w3202 & w3356;
assign w3358 = ~w3202 & ~w3356;
assign w3359 = ~w3357 & ~w3358;
assign w3360 = ~w2948 & ~w3359;
assign w3361 = ~pi529 & ~w3360;
assign w3362 = w2948 & w3359;
assign w3363 = w3361 & ~w3362;
assign w3364 = pi303 & pi478;
assign w3365 = pi529 & ~w3364;
assign w3366 = ~pi303 & ~pi478;
assign w3367 = w3365 & ~w3366;
assign w3368 = ~w3363 & ~w3367;
assign w3369 = ~pi077 & ~pi109;
assign w3370 = ~pi043 & w3369;
assign w3371 = pi076 & pi077;
assign w3372 = pi043 & ~pi109;
assign w3373 = w3371 & w3372;
assign w3374 = ~w3370 & ~w3373;
assign w3375 = ~pi070 & ~pi077;
assign w3376 = pi076 & w3375;
assign w3377 = ~pi076 & pi077;
assign w3378 = ~w3376 & ~w3377;
assign w3379 = w3374 & w3378;
assign w3380 = pi039 & ~w3379;
assign w3381 = pi077 & pi109;
assign w3382 = ~pi043 & ~pi076;
assign w3383 = w3381 & w3382;
assign w3384 = pi070 & ~pi109;
assign w3385 = w3371 & w3384;
assign w3386 = pi070 & ~pi077;
assign w3387 = ~pi043 & pi076;
assign w3388 = w3386 & w3387;
assign w3389 = ~w3383 & ~w3385;
assign w3390 = ~w3388 & w3389;
assign w3391 = ~pi070 & pi109;
assign w3392 = w3371 & ~w3391;
assign w3393 = ~w3376 & ~w3392;
assign w3394 = ~pi070 & pi122;
assign w3395 = ~pi076 & pi109;
assign w3396 = ~pi043 & w3395;
assign w3397 = pi043 & ~pi076;
assign w3398 = w3386 & w3397;
assign w3399 = w3394 & w3396;
assign w3400 = ~w3398 & ~w3399;
assign w3401 = pi077 & ~pi109;
assign w3402 = pi070 & w3401;
assign w3403 = w3401 & w18266;
assign w3404 = ~pi076 & pi122;
assign w3405 = ~pi043 & w3401;
assign w3406 = ~w3404 & w3405;
assign w3407 = ~w3403 & ~w3406;
assign w3408 = w3400 & w3407;
assign w3409 = ~pi077 & pi109;
assign w3410 = ~pi043 & ~pi070;
assign w3411 = w3409 & w3410;
assign w3412 = pi043 & pi076;
assign w3413 = w3381 & w3412;
assign w3414 = ~pi070 & w3413;
assign w3415 = ~pi122 & w3411;
assign w3416 = ~w3414 & ~w3415;
assign w3417 = pi076 & w3401;
assign w3418 = ~pi043 & ~pi122;
assign w3419 = ~pi070 & pi077;
assign w3420 = pi122 & w3397;
assign w3421 = w3384 & w3387;
assign w3422 = w3419 & w3420;
assign w3423 = ~w3421 & ~w3422;
assign w3424 = w3417 & w3418;
assign w3425 = w3423 & ~w3424;
assign w3426 = pi039 & ~w3416;
assign w3427 = w3425 & ~w3426;
assign w3428 = (~pi039 & ~w3408) | (~pi039 & w18267) | (~w3408 & w18267);
assign w3429 = w3427 & ~w3428;
assign w3430 = (pi122 & w3380) | (pi122 & w18268) | (w3380 & w18268);
assign w3431 = ~pi077 & w3412;
assign w3432 = w3372 & w3419;
assign w3433 = ~w3431 & ~w3432;
assign w3434 = ~pi122 & ~w3433;
assign w3435 = pi122 & w3387;
assign w3436 = w3419 & w3435;
assign w3437 = w3371 & w3391;
assign w3438 = ~pi043 & w3437;
assign w3439 = pi043 & pi070;
assign w3440 = w3409 & w3439;
assign w3441 = ~w3436 & ~w3438;
assign w3442 = ~w3434 & w3441;
assign w3443 = pi070 & w3381;
assign w3444 = pi070 & pi076;
assign w3445 = w3369 & w3444;
assign w3446 = ~w3443 & ~w3445;
assign w3447 = (pi122 & w3446) | (pi122 & w18269) | (w3446 & w18269);
assign w3448 = w3402 & w3412;
assign w3449 = ~pi043 & pi070;
assign w3450 = w3381 & w3449;
assign w3451 = w3382 & w3384;
assign w3452 = ~w3450 & ~w3451;
assign w3453 = ~pi070 & pi076;
assign w3454 = w3369 & w3453;
assign w3455 = ~w3448 & w3452;
assign w3456 = ~pi122 & ~w3454;
assign w3457 = w3455 & w3456;
assign w3458 = ~pi070 & w3369;
assign w3459 = ~pi039 & pi122;
assign w3460 = ~w3420 & ~w3459;
assign w3461 = w3458 & ~w3460;
assign w3462 = pi122 & ~w3439;
assign w3463 = w3395 & ~w3462;
assign w3464 = pi043 & pi122;
assign w3465 = pi076 & w3391;
assign w3466 = w3464 & w3465;
assign w3467 = ~w3463 & ~w3466;
assign w3468 = ~pi039 & ~w3467;
assign w3469 = ~w3461 & ~w3468;
assign w3470 = ~w3447 & ~w3457;
assign w3471 = w3469 & ~w3470;
assign w3472 = pi070 & pi077;
assign w3473 = w3395 & w3472;
assign w3474 = ~pi076 & ~pi109;
assign w3475 = w3419 & w3474;
assign w3476 = ~w3473 & ~w3475;
assign w3477 = w3386 & ~w3395;
assign w3478 = (pi043 & ~w3476) | (pi043 & w18270) | (~w3476 & w18270);
assign w3479 = ~pi122 & ~w3478;
assign w3480 = w3372 & w3472;
assign w3481 = w3395 & w3419;
assign w3482 = ~w3383 & ~w3480;
assign w3483 = pi122 & ~w3481;
assign w3484 = w3482 & w3483;
assign w3485 = pi076 & w3411;
assign w3486 = pi070 & w3369;
assign w3487 = w3382 & w3486;
assign w3488 = ~w3485 & ~w3487;
assign w3489 = w3484 & w3488;
assign w3490 = pi039 & ~w3489;
assign w3491 = pi070 & pi109;
assign w3492 = w3387 & w3491;
assign w3493 = w3391 & w3397;
assign w3494 = ~w3492 & ~w3493;
assign w3495 = w3452 & w3494;
assign w3496 = pi122 & ~w3492;
assign w3497 = (~pi039 & w3492) | (~pi039 & w3759) | (w3492 & w3759);
assign w3498 = ~w3495 & w3497;
assign w3499 = w3372 & w3453;
assign w3500 = ~pi077 & w3499;
assign w3501 = ~pi076 & w3401;
assign w3502 = w3449 & w3501;
assign w3503 = ~w3500 & ~w3502;
assign w3504 = ~pi122 & ~w3503;
assign w3505 = w3372 & w3375;
assign w3506 = w3371 & w3449;
assign w3507 = ~w3505 & ~w3506;
assign w3508 = ~w3414 & w3507;
assign w3509 = w3459 & ~w3508;
assign w3510 = ~w3498 & ~w3504;
assign w3511 = ~w3509 & w3510;
assign w3512 = ~w3479 & w3490;
assign w3513 = w3511 & ~w3512;
assign w3514 = (~pi017 & ~w3471) | (~pi017 & w18271) | (~w3471 & w18271);
assign w3515 = w3513 & ~w3514;
assign w3516 = (pi017 & ~w3429) | (pi017 & w18272) | (~w3429 & w18272);
assign w3517 = w3515 & ~w3516;
assign w3518 = ~pi052 & ~pi084;
assign w3519 = pi004 & w3518;
assign w3520 = ~pi004 & pi052;
assign w3521 = ~w3519 & ~w3520;
assign w3522 = pi052 & ~pi094;
assign w3523 = pi005 & w3522;
assign w3524 = ~pi052 & ~pi094;
assign w3525 = ~pi005 & w3524;
assign w3526 = ~w3523 & ~w3525;
assign w3527 = w3521 & w3526;
assign w3528 = pi091 & ~w3527;
assign w3529 = pi052 & pi094;
assign w3530 = pi004 & ~pi084;
assign w3531 = w3529 & w3530;
assign w3532 = pi005 & w3531;
assign w3533 = ~pi052 & pi094;
assign w3534 = ~pi005 & ~pi084;
assign w3535 = w3533 & w3534;
assign w3536 = ~pi091 & w3535;
assign w3537 = ~w3532 & ~w3536;
assign w3538 = (pi024 & w3528) | (pi024 & w18273) | (w3528 & w18273);
assign w3539 = pi052 & pi084;
assign w3540 = pi004 & w3539;
assign w3541 = pi004 & w3522;
assign w3542 = ~w3519 & ~w3540;
assign w3543 = pi004 & ~pi005;
assign w3544 = pi091 & ~w3543;
assign w3545 = pi005 & ~pi084;
assign w3546 = ~pi004 & ~pi084;
assign w3547 = ~pi005 & pi091;
assign w3548 = pi094 & w3547;
assign w3549 = ~pi052 & pi084;
assign w3550 = ~pi004 & pi005;
assign w3551 = w3549 & w3550;
assign w3552 = w3546 & w3548;
assign w3553 = ~w3551 & ~w3552;
assign w3554 = w3522 & ~w3545;
assign w3555 = ~w3544 & w3554;
assign w3556 = w3553 & ~w3555;
assign w3557 = (~pi024 & ~w3556) | (~pi024 & w18275) | (~w3556 & w18275);
assign w3558 = w3539 & w18279;
assign w3559 = w3543 & w3549;
assign w3560 = ~pi004 & ~pi005;
assign w3561 = w3529 & w3560;
assign w3562 = ~w3559 & ~w3561;
assign w3563 = ~w3558 & w3562;
assign w3564 = pi091 & ~w3563;
assign w3565 = pi052 & ~pi084;
assign w3566 = pi005 & pi091;
assign w3567 = ~pi004 & w3566;
assign w3568 = ~pi005 & ~pi091;
assign w3569 = w3522 & w3568;
assign w3570 = pi084 & ~pi094;
assign w3571 = w3543 & w3570;
assign w3572 = pi018 & ~w3571;
assign w3573 = pi004 & w3569;
assign w3574 = w3572 & ~w3573;
assign w3575 = w3565 & w3567;
assign w3576 = w3574 & ~w3575;
assign w3577 = ~w3538 & ~w3557;
assign w3578 = ~w3564 & w3576;
assign w3579 = w3577 & w3578;
assign w3580 = pi004 & pi005;
assign w3581 = ~pi052 & w3580;
assign w3582 = w3522 & w3545;
assign w3583 = ~w3581 & ~w3582;
assign w3584 = ~pi091 & ~w3583;
assign w3585 = ~pi005 & w3531;
assign w3586 = pi005 & pi084;
assign w3587 = w3533 & w3586;
assign w3588 = pi091 & w3543;
assign w3589 = w3565 & w3588;
assign w3590 = ~w3587 & ~w3589;
assign w3591 = ~w3584 & w3590;
assign w3592 = (pi024 & ~w3591) | (pi024 & w18276) | (~w3591 & w18276);
assign w3593 = ~pi004 & pi094;
assign w3594 = pi091 & ~w3586;
assign w3595 = ~pi084 & pi094;
assign w3596 = pi004 & w3595;
assign w3597 = ~pi094 & w3518;
assign w3598 = w3518 & w18277;
assign w3599 = w3566 & w3596;
assign w3600 = ~w3598 & ~w3599;
assign w3601 = (~pi024 & ~w3600) | (~pi024 & w18278) | (~w3600 & w18278);
assign w3602 = w3541 & w3586;
assign w3603 = w3518 & w18279;
assign w3604 = pi084 & w3529;
assign w3605 = ~pi004 & w3570;
assign w3606 = ~w3604 & ~w3605;
assign w3607 = w3568 & ~w3606;
assign w3608 = pi004 & pi084;
assign w3609 = ~pi004 & ~pi094;
assign w3610 = w3518 & w3609;
assign w3611 = ~w3524 & ~w3529;
assign w3612 = w3566 & ~w3611;
assign w3613 = ~w3608 & ~w3610;
assign w3614 = w3612 & ~w3613;
assign w3615 = ~w3607 & ~w3614;
assign w3616 = (~pi091 & w3602) | (~pi091 & w18280) | (w3602 & w18280);
assign w3617 = w3615 & w20766;
assign w3618 = w3617 & w18281;
assign w3619 = ~w3579 & ~w3618;
assign w3620 = ~pi004 & pi084;
assign w3621 = w3524 & w3620;
assign w3622 = (pi094 & w3519) | (pi094 & w18282) | (w3519 & w18282);
assign w3623 = pi005 & pi052;
assign w3624 = w3570 & w3623;
assign w3625 = w3520 & w3595;
assign w3626 = ~w3624 & ~w3625;
assign w3627 = pi091 & w3626;
assign w3628 = (~pi005 & w3622) | (~pi005 & w18283) | (w3622 & w18283);
assign w3629 = w3627 & ~w3628;
assign w3630 = w3522 & w3546;
assign w3631 = pi084 & pi094;
assign w3632 = w3520 & w3631;
assign w3633 = ~w3630 & ~w3632;
assign w3634 = w3549 & ~w3593;
assign w3635 = (pi005 & ~w3633) | (pi005 & w18284) | (~w3633 & w18284);
assign w3636 = (pi024 & w3635) | (pi024 & w3858) | (w3635 & w3858);
assign w3637 = ~w3629 & w3636;
assign w3638 = w3543 & w3631;
assign w3639 = ~pi084 & w3550;
assign w3640 = ~pi091 & pi094;
assign w3641 = w3639 & w3640;
assign w3642 = ~w3638 & ~w3641;
assign w3643 = ~w3607 & w3642;
assign w3644 = ~pi024 & ~w3643;
assign w3645 = pi084 & w3522;
assign w3646 = w3560 & w3645;
assign w3647 = pi005 & ~pi052;
assign w3648 = ~pi084 & ~pi094;
assign w3649 = w3647 & w3648;
assign w3650 = pi004 & w3649;
assign w3651 = ~w3646 & ~w3650;
assign w3652 = ~pi024 & pi091;
assign w3653 = w3539 & w3543;
assign w3654 = ~w3532 & w18285;
assign w3655 = w3652 & ~w3654;
assign w3656 = ~pi091 & ~w3651;
assign w3657 = ~w3655 & ~w3656;
assign w3658 = ~w3644 & w3657;
assign w3659 = ~w3637 & w3658;
assign w3660 = ~w3619 & w3659;
assign w3661 = ~w3517 & w3660;
assign w3662 = w3517 & ~w3660;
assign w3663 = ~w3661 & ~w3662;
assign w3664 = ~w3405 & ~w3458;
assign w3665 = ~w3372 & w3386;
assign w3666 = ~w3465 & ~w3665;
assign w3667 = pi043 & ~pi070;
assign w3668 = w3381 & w3667;
assign w3669 = w3409 & w3444;
assign w3670 = ~w3492 & ~w3668;
assign w3671 = ~w3669 & w3670;
assign w3672 = pi122 & ~w3666;
assign w3673 = w3671 & ~w3672;
assign w3674 = w3381 & w3410;
assign w3675 = ~w3432 & ~w3674;
assign w3676 = ~pi122 & ~w3675;
assign w3677 = ~pi076 & ~pi122;
assign w3678 = pi070 & w3474;
assign w3679 = w3409 & w3667;
assign w3680 = ~w3678 & ~w3679;
assign w3681 = ~w3677 & ~w3680;
assign w3682 = pi070 & pi122;
assign w3683 = w3401 & w3682;
assign w3684 = w3369 & w3382;
assign w3685 = w3382 & w3472;
assign w3686 = ~w3683 & ~w3684;
assign w3687 = ~w3685 & w3686;
assign w3688 = ~w3681 & w3687;
assign w3689 = (~pi039 & ~w3688) | (~pi039 & w18286) | (~w3688 & w18286);
assign w3690 = w3395 & w3410;
assign w3691 = ~pi043 & w3669;
assign w3692 = pi043 & pi077;
assign w3693 = w3692 & w3491;
assign w3694 = ~w3691 & w18287;
assign w3695 = ~pi122 & ~w3694;
assign w3696 = pi076 & pi122;
assign w3697 = pi043 & w3409;
assign w3698 = ~w3401 & ~w3409;
assign w3699 = ~pi070 & ~w3698;
assign w3700 = (w3696 & w3699) | (w3696 & w18288) | (w3699 & w18288);
assign w3701 = pi070 & ~pi076;
assign w3702 = w3692 & w3701;
assign w3703 = ~pi109 & w3702;
assign w3704 = ~w3700 & ~w3703;
assign w3705 = ~w3695 & w3704;
assign w3706 = ~w3689 & w3705;
assign w3707 = (pi017 & ~w3706) | (pi017 & w18289) | (~w3706 & w18289);
assign w3708 = ~pi070 & ~pi109;
assign w3709 = ~pi076 & w3708;
assign w3710 = w3417 & w3449;
assign w3711 = w3382 & w3443;
assign w3712 = w3412 & w3491;
assign w3713 = pi077 & w3712;
assign w3714 = w3409 & w3701;
assign w3715 = ~pi122 & w3714;
assign w3716 = ~w3713 & ~w3715;
assign w3717 = ~w3679 & ~w3711;
assign w3718 = w3716 & w3717;
assign w3719 = pi043 & ~pi122;
assign w3720 = w3669 & w3719;
assign w3721 = ~pi043 & pi122;
assign w3722 = ~w3453 & ~w3696;
assign w3723 = w3369 & ~w3722;
assign w3724 = ~w3375 & w3721;
assign w3725 = pi109 & w3724;
assign w3726 = ~w3723 & ~w3725;
assign w3727 = ~w3690 & ~w3720;
assign w3728 = w3726 & w3727;
assign w3729 = ~pi039 & ~w3728;
assign w3730 = pi076 & w3450;
assign w3731 = ~w3373 & ~w3730;
assign w3732 = pi077 & w3708;
assign w3733 = w3382 & w3732;
assign w3734 = pi122 & w3473;
assign w3735 = ~w3733 & ~w3734;
assign w3736 = w3464 & w3709;
assign w3737 = w3735 & ~w3736;
assign w3738 = (~pi122 & w3730) | (~pi122 & w18292) | (w3730 & w18292);
assign w3739 = w3737 & ~w3738;
assign w3740 = ~w3729 & w3739;
assign w3741 = (~pi017 & ~w3740) | (~pi017 & w18293) | (~w3740 & w18293);
assign w3742 = ~w3376 & ~w3501;
assign w3743 = (w3418 & ~w3742) | (w3418 & w18294) | (~w3742 & w18294);
assign w3744 = pi122 & w3669;
assign w3745 = w3375 & w3395;
assign w3746 = w3719 & w3745;
assign w3747 = ~w3744 & ~w3746;
assign w3748 = ~w3743 & w3747;
assign w3749 = pi039 & ~w3748;
assign w3750 = w3391 & w18295;
assign w3751 = ~w3481 & ~w3750;
assign w3752 = w3464 & ~w3751;
assign w3753 = w3387 & w3458;
assign w3754 = ~w3733 & ~w3753;
assign w3755 = w3459 & ~w3754;
assign w3756 = pi039 & pi122;
assign w3757 = ~w3668 & ~w3702;
assign w3758 = w3756 & ~w3757;
assign w3759 = ~pi039 & ~pi122;
assign w3760 = w3395 & w3692;
assign w3761 = w3371 & w3708;
assign w3762 = pi043 & w3761;
assign w3763 = w3759 & w3760;
assign w3764 = ~w3762 & ~w3763;
assign w3765 = ~w3752 & ~w3755;
assign w3766 = ~w3758 & w3764;
assign w3767 = w3765 & w3766;
assign w3768 = ~w3749 & w3767;
assign w3769 = ~w3741 & w3768;
assign w3770 = ~w3707 & w3769;
assign w3771 = w3529 & w3534;
assign w3772 = ~w3582 & ~w3771;
assign w3773 = ~pi004 & ~pi091;
assign w3774 = w3533 & w3545;
assign w3775 = ~w3605 & ~w3774;
assign w3776 = ~w3773 & ~w3775;
assign w3777 = w3522 & w18296;
assign w3778 = w3524 & w3560;
assign w3779 = w3539 & w3560;
assign w3780 = ~w3778 & ~w3779;
assign w3781 = ~w3777 & w3780;
assign w3782 = ~w3776 & w3781;
assign w3783 = ~pi005 & w3549;
assign w3784 = pi084 & w3533;
assign w3785 = ~w3596 & ~w3783;
assign w3786 = (pi091 & ~w3785) | (pi091 & w18297) | (~w3785 & w18297);
assign w3787 = ~pi091 & w3597;
assign w3788 = w3533 & w3608;
assign w3789 = w3529 & w3545;
assign w3790 = ~w3569 & ~w3638;
assign w3791 = ~w3788 & ~w3789;
assign w3792 = w3790 & w3791;
assign w3793 = ~w3787 & w3792;
assign w3794 = (pi024 & ~w3793) | (pi024 & w18298) | (~w3793 & w18298);
assign w3795 = ~pi052 & w3638;
assign w3796 = w3560 & w3595;
assign w3797 = w3529 & w3586;
assign w3798 = ~w3796 & ~w3797;
assign w3799 = ~w3795 & w3798;
assign w3800 = ~pi091 & ~w3799;
assign w3801 = pi004 & pi091;
assign w3802 = ~pi084 & w3533;
assign w3803 = ~pi084 & w3522;
assign w3804 = ~w3802 & ~w3803;
assign w3805 = pi005 & w3533;
assign w3806 = (w3801 & ~w3804) | (w3801 & w18299) | (~w3804 & w18299);
assign w3807 = w3550 & w3645;
assign w3808 = ~w3800 & w18300;
assign w3809 = ~w3794 & w3808;
assign w3810 = (pi018 & ~w3809) | (pi018 & w18301) | (~w3809 & w18301);
assign w3811 = ~pi004 & w3648;
assign w3812 = pi052 & w3543;
assign w3813 = w3570 & w3812;
assign w3814 = w3773 & w3784;
assign w3815 = ~w3774 & ~w3814;
assign w3816 = pi094 & w3779;
assign w3817 = w3580 & w3604;
assign w3818 = ~w3816 & ~w3817;
assign w3819 = w3815 & w3818;
assign w3820 = ~w3518 & w3548;
assign w3821 = ~w3796 & ~w3820;
assign w3822 = pi005 & ~pi091;
assign w3823 = w3788 & w3822;
assign w3824 = ~w3530 & ~w3801;
assign w3825 = w3524 & ~w3824;
assign w3826 = ~w3823 & ~w3825;
assign w3827 = w3821 & w3826;
assign w3828 = ~pi024 & ~w3827;
assign w3829 = w3631 & w3812;
assign w3830 = w3522 & w3580;
assign w3831 = (~pi091 & w3829) | (~pi091 & w18303) | (w3829 & w18303);
assign w3832 = w3566 & w3811;
assign w3833 = w3522 & w3560;
assign w3834 = pi091 & w3632;
assign w3835 = ~pi084 & w3833;
assign w3836 = ~w3834 & ~w3835;
assign w3837 = ~w3832 & w3836;
assign w3838 = ~w3831 & w3837;
assign w3839 = ~w3828 & w3838;
assign w3840 = ~pi004 & w3522;
assign w3841 = w3533 & w3620;
assign w3842 = ~w3519 & ~w3841;
assign w3843 = (w3568 & ~w3842) | (w3568 & w18305) | (~w3842 & w18305);
assign w3844 = w3802 & w3822;
assign w3845 = w3802 & w18306;
assign w3846 = pi091 & w3788;
assign w3847 = ~w3845 & ~w3846;
assign w3848 = ~w3843 & w3847;
assign w3849 = pi024 & ~w3848;
assign w3850 = w3547 & w3630;
assign w3851 = ~pi094 & w3543;
assign w3852 = w3518 & w3851;
assign w3853 = ~w3850 & ~w3852;
assign w3854 = w3652 & ~w3853;
assign w3855 = w3530 & w3533;
assign w3856 = ~w3625 & ~w3855;
assign w3857 = w3566 & ~w3856;
assign w3858 = pi024 & pi091;
assign w3859 = w3623 & w3858;
assign w3860 = w3529 & w3550;
assign w3861 = w3523 & w3530;
assign w3862 = ~pi024 & ~pi091;
assign w3863 = w3860 & w3862;
assign w3864 = ~w3861 & ~w3863;
assign w3865 = ~w3608 & ~w3648;
assign w3866 = w3859 & w3865;
assign w3867 = w3864 & ~w3866;
assign w3868 = ~w3854 & w3867;
assign w3869 = ~w3857 & w3868;
assign w3870 = ~w3849 & w3869;
assign w3871 = (~pi018 & ~w3839) | (~pi018 & w18307) | (~w3839 & w18307);
assign w3872 = w3870 & ~w3871;
assign w3873 = ~w3810 & w3872;
assign w3874 = ~w3770 & w3873;
assign w3875 = w3770 & ~w3873;
assign w3876 = ~w3874 & ~w3875;
assign w3877 = w3663 & ~w3876;
assign w3878 = ~w3663 & w3876;
assign w3879 = ~w3877 & ~w3878;
assign w3880 = ~pi077 & w3493;
assign w3881 = w3382 & w3409;
assign w3882 = ~w3669 & ~w3881;
assign w3883 = ~w3880 & w3882;
assign w3884 = ~pi122 & ~w3883;
assign w3885 = w3465 & w3721;
assign w3886 = ~w3373 & ~w3683;
assign w3887 = ~w3885 & w3886;
assign w3888 = (pi039 & w3884) | (pi039 & w18308) | (w3884 & w18308);
assign w3889 = ~w3394 & ~w3397;
assign w3890 = w3369 & ~w3889;
assign w3891 = w3472 & w3696;
assign w3892 = ~w3890 & ~w3891;
assign w3893 = (~pi039 & ~w3892) | (~pi039 & w18309) | (~w3892 & w18309);
assign w3894 = w3382 & w3419;
assign w3895 = w3437 & w3418;
assign w3896 = ~w3487 & ~w3895;
assign w3897 = (pi122 & w3500) | (pi122 & w18310) | (w3500 & w18310);
assign w3898 = w3896 & ~w3897;
assign w3899 = ~w3893 & w3898;
assign w3900 = ~w3888 & w3899;
assign w3901 = ~pi017 & ~w3900;
assign w3902 = ~w3501 & ~w3750;
assign w3903 = ~pi122 & ~w3902;
assign w3904 = ~pi109 & w3398;
assign w3905 = w3404 & w3409;
assign w3906 = ~w3753 & ~w3904;
assign w3907 = pi039 & ~w3905;
assign w3908 = w3906 & w3907;
assign w3909 = ~pi039 & ~w3760;
assign w3910 = ~w3744 & w3909;
assign w3911 = w3369 & w3412;
assign w3912 = ~pi122 & w3911;
assign w3913 = ~pi043 & ~w3677;
assign w3914 = w3491 & ~w3913;
assign w3915 = ~w3912 & ~w3914;
assign w3916 = w3910 & w3915;
assign w3917 = ~w3903 & w3908;
assign w3918 = ~w3916 & ~w3917;
assign w3919 = pi122 & ~w3679;
assign w3920 = ~pi077 & w3397;
assign w3921 = ~pi109 & w3387;
assign w3922 = ~w3473 & ~w3921;
assign w3923 = ~pi076 & w3369;
assign w3924 = w3410 & w3923;
assign w3925 = w3372 & w3377;
assign w3926 = ~w3668 & ~w3925;
assign w3927 = ~w3924 & w3926;
assign w3928 = ~pi122 & w3927;
assign w3929 = w3919 & w3922;
assign w3930 = ~w3920 & w3929;
assign w3931 = ~w3928 & ~w3930;
assign w3932 = (pi017 & w3918) | (pi017 & w18311) | (w3918 & w18311);
assign w3933 = ~pi122 & w3475;
assign w3934 = (pi043 & w3933) | (pi043 & w18312) | (w3933 & w18312);
assign w3935 = ~w3369 & w3667;
assign w3936 = ~w3711 & ~w3924;
assign w3937 = (~pi122 & ~w3936) | (~pi122 & w18313) | (~w3936 & w18313);
assign w3938 = ~w3414 & ~w3880;
assign w3939 = ~pi039 & ~w3934;
assign w3940 = ~w3934 & w3938;
assign w3941 = ~w3937 & w3940;
assign w3942 = ~w3939 & ~w3941;
assign w3943 = w3369 & w3449;
assign w3944 = ~w3398 & ~w3480;
assign w3945 = ~w3943 & w3944;
assign w3946 = w3375 & w3396;
assign w3947 = pi109 & w3412;
assign w3948 = w3375 & w3947;
assign w3949 = ~w3946 & ~w3948;
assign w3950 = w3945 & w3949;
assign w3951 = pi122 & ~w3950;
assign w3952 = ~w3474 & ~w3692;
assign w3953 = pi109 & w3702;
assign w3954 = w3419 & w3952;
assign w3955 = ~w3953 & ~w3954;
assign w3956 = ~w3448 & ~w3487;
assign w3957 = ~pi039 & w3956;
assign w3958 = ~pi122 & ~w3955;
assign w3959 = w3957 & ~w3958;
assign w3960 = w3464 & w3486;
assign w3961 = (pi039 & ~w3486) | (pi039 & w18314) | (~w3486 & w18314);
assign w3962 = w3417 & w3721;
assign w3963 = w3961 & ~w3962;
assign w3964 = ~w3951 & w3959;
assign w3965 = ~w3963 & ~w3964;
assign w3966 = ~w3901 & ~w3932;
assign w3967 = ~w3942 & ~w3965;
assign w3968 = w3966 & w3967;
assign w3969 = pi035 & ~pi100;
assign w3970 = ~pi031 & w3969;
assign w3971 = ~pi100 & ~pi128;
assign w3972 = ~pi035 & w3971;
assign w3973 = pi100 & ~pi128;
assign w3974 = pi035 & w3973;
assign w3975 = ~w3972 & ~w3974;
assign w3976 = (pi037 & ~w3975) | (pi037 & w18315) | (~w3975 & w18315);
assign w3977 = ~pi037 & ~pi100;
assign w3978 = ~pi031 & ~pi035;
assign w3979 = w3977 & w3978;
assign w3980 = pi128 & w3979;
assign w3981 = ~pi037 & pi128;
assign w3982 = pi031 & pi035;
assign w3983 = ~pi100 & w3982;
assign w3984 = w3981 & w3983;
assign w3985 = ~w3980 & ~w3984;
assign w3986 = ~w3976 & w3985;
assign w3987 = pi106 & ~w3986;
assign w3988 = pi031 & ~pi035;
assign w3989 = ~pi037 & pi100;
assign w3990 = ~pi128 & w3989;
assign w3991 = w3988 & w3990;
assign w3992 = pi100 & pi128;
assign w3993 = ~pi035 & ~pi037;
assign w3994 = w3992 & w3993;
assign w3995 = ~pi031 & pi035;
assign w3996 = pi037 & w3992;
assign w3997 = w3995 & w3996;
assign w3998 = ~w3991 & ~w3997;
assign w3999 = (~pi106 & ~w3998) | (~pi106 & w4112) | (~w3998 & w4112);
assign w4000 = pi037 & w3973;
assign w4001 = w3982 & w4000;
assign w4002 = ~pi031 & w3971;
assign w4003 = ~pi035 & pi037;
assign w4004 = w4002 & w4003;
assign w4005 = ~w4001 & ~w4004;
assign w4006 = ~pi065 & w4005;
assign w4007 = ~w3999 & w4006;
assign w4008 = w3978 & w3996;
assign w4009 = w3993 & w4002;
assign w4010 = pi035 & ~pi037;
assign w4011 = ~w3971 & w4010;
assign w4012 = ~w4008 & ~w4009;
assign w4013 = (~pi106 & ~w4012) | (~pi106 & w18316) | (~w4012 & w18316);
assign w4014 = w3970 & w3981;
assign w4015 = pi035 & pi106;
assign w4016 = pi037 & w3971;
assign w4017 = w4015 & w4016;
assign w4018 = pi031 & ~pi037;
assign w4019 = pi035 & w3992;
assign w4020 = w4018 & w4019;
assign w4021 = ~pi035 & pi106;
assign w4022 = pi031 & w3973;
assign w4023 = w4021 & w4022;
assign w4024 = ~w4020 & ~w4023;
assign w4025 = ~w4014 & ~w4017;
assign w4026 = w4024 & w4025;
assign w4027 = pi065 & w4026;
assign w4028 = ~w3987 & w4007;
assign w4029 = ~w4013 & w4027;
assign w4030 = ~w4028 & ~w4029;
assign w4031 = pi037 & pi100;
assign w4032 = pi031 & pi106;
assign w4033 = w4031 & w4032;
assign w4034 = ~pi031 & w3973;
assign w4035 = ~pi037 & ~pi106;
assign w4036 = w4034 & w4035;
assign w4037 = ~pi100 & pi128;
assign w4038 = w4018 & w4037;
assign w4039 = ~w4034 & ~w4038;
assign w4040 = ~pi106 & ~w4039;
assign w4041 = w3971 & w4018;
assign w4042 = ~pi035 & w4041;
assign w4043 = (pi065 & ~w4041) | (pi065 & w18317) | (~w4041 & w18317);
assign w4044 = ~pi031 & pi037;
assign w4045 = ~pi128 & w4044;
assign w4046 = w3969 & w4045;
assign w4047 = ~pi031 & pi106;
assign w4048 = w4037 & w4047;
assign w4049 = ~w4040 & w4043;
assign w4050 = ~w4046 & ~w4048;
assign w4051 = w4049 & w4050;
assign w4052 = pi031 & w3971;
assign w4053 = pi035 & ~pi106;
assign w4054 = (~pi065 & ~w4052) | (~pi065 & w18318) | (~w4052 & w18318);
assign w4055 = pi031 & pi037;
assign w4056 = w4037 & w4055;
assign w4057 = pi106 & w4056;
assign w4058 = w3992 & w3995;
assign w4059 = pi037 & pi128;
assign w4060 = ~pi031 & ~pi106;
assign w4061 = ~pi035 & ~w4060;
assign w4062 = w4059 & ~w4061;
assign w4063 = ~w4057 & ~w4058;
assign w4064 = w4063 & w18319;
assign w4065 = w4010 & w4037;
assign w4066 = pi106 & ~w4065;
assign w4067 = ~pi035 & ~pi128;
assign w4068 = pi031 & w4067;
assign w4069 = w3992 & w4044;
assign w4070 = ~w3970 & ~w4068;
assign w4071 = w4066 & w4070;
assign w4072 = ~w4069 & w4071;
assign w4073 = w3992 & w4010;
assign w4074 = w3973 & w3995;
assign w4075 = ~w4073 & ~w4074;
assign w4076 = ~w4009 & w4075;
assign w4077 = ~pi106 & w4076;
assign w4078 = ~w4072 & ~w4077;
assign w4079 = pi068 & ~w4078;
assign w4080 = ~w4051 & ~w4064;
assign w4081 = w4079 & ~w4080;
assign w4082 = pi037 & w3995;
assign w4083 = ~w4018 & w4037;
assign w4084 = ~w4082 & w4083;
assign w4085 = ~pi106 & w4084;
assign w4086 = pi037 & pi106;
assign w4087 = w3973 & w4086;
assign w4088 = pi128 & w4018;
assign w4089 = w4021 & w4088;
assign w4090 = w3973 & w3982;
assign w4091 = ~w4087 & ~w4090;
assign w4092 = ~w4089 & w4091;
assign w4093 = pi065 & w4092;
assign w4094 = pi106 & ~pi128;
assign w4095 = w3977 & w4094;
assign w4096 = ~pi128 & w3995;
assign w4097 = w3995 & w3971;
assign w4098 = ~pi035 & ~pi106;
assign w4099 = w3973 & w4098;
assign w4100 = pi037 & w4099;
assign w4101 = ~w4097 & ~w4100;
assign w4102 = ~w4033 & ~w4095;
assign w4103 = ~pi065 & w4102;
assign w4104 = w4101 & w4103;
assign w4105 = ~w4085 & w4093;
assign w4106 = ~pi031 & pi100;
assign w4107 = w3971 & w3982;
assign w4108 = ~pi037 & w4106;
assign w4109 = ~w4107 & ~w4108;
assign w4110 = ~w4021 & ~w4095;
assign w4111 = ~w4109 & ~w4110;
assign w4112 = ~pi106 & w3994;
assign w4113 = w3994 & w4838;
assign w4114 = (~pi068 & ~w4002) | (~pi068 & w18320) | (~w4002 & w18320);
assign w4115 = ~w4113 & w4114;
assign w4116 = ~w4111 & w4115;
assign w4117 = (w4116 & w4105) | (w4116 & w18321) | (w4105 & w18321);
assign w4118 = ~w4081 & ~w4117;
assign w4119 = (pi035 & w4036) | (pi035 & w18322) | (w4036 & w18322);
assign w4120 = ~w4118 & w18323;
assign w4121 = ~w3968 & w4120;
assign w4122 = w3968 & ~w4120;
assign w4123 = ~w4121 & ~w4122;
assign w4124 = ~pi025 & pi125;
assign w4125 = ~pi113 & ~w4124;
assign w4126 = ~pi055 & pi124;
assign w4127 = pi009 & ~pi125;
assign w4128 = pi025 & w4127;
assign w4129 = w4125 & ~w4128;
assign w4130 = w4126 & w4129;
assign w4131 = pi025 & pi055;
assign w4132 = ~pi124 & w4131;
assign w4133 = w4131 & w18324;
assign w4134 = ~pi025 & pi124;
assign w4135 = pi113 & pi125;
assign w4136 = ~pi009 & w4135;
assign w4137 = pi009 & pi125;
assign w4138 = pi055 & ~pi124;
assign w4139 = w4137 & w4138;
assign w4140 = w4134 & w4136;
assign w4141 = ~w4139 & ~w4140;
assign w4142 = ~w4130 & w4141;
assign w4143 = (pi096 & ~w4142) | (pi096 & w18325) | (~w4142 & w18325);
assign w4144 = ~pi055 & ~pi124;
assign w4145 = ~pi025 & w4144;
assign w4146 = pi125 & w4131;
assign w4147 = ~w4145 & ~w4146;
assign w4148 = pi113 & ~w4147;
assign w4149 = ~pi055 & w4127;
assign w4150 = ~pi009 & ~pi113;
assign w4151 = w4131 & w4150;
assign w4152 = ~w4149 & ~w4151;
assign w4153 = ~pi124 & ~w4152;
assign w4154 = ~w4148 & ~w4153;
assign w4155 = ~pi025 & ~pi124;
assign w4156 = ~pi055 & w4137;
assign w4157 = w4155 & w4156;
assign w4158 = ~pi009 & ~pi125;
assign w4159 = ~pi025 & pi055;
assign w4160 = w4158 & w4159;
assign w4161 = (pi113 & w4157) | (pi113 & w18326) | (w4157 & w18326);
assign w4162 = pi055 & pi124;
assign w4163 = w4124 & w4162;
assign w4164 = ~pi113 & w4163;
assign w4165 = w4163 & w4150;
assign w4166 = ~pi009 & pi025;
assign w4167 = w4144 & w4166;
assign w4168 = ~pi125 & w4167;
assign w4169 = (pi010 & ~w4167) | (pi010 & w18327) | (~w4167 & w18327);
assign w4170 = ~w4165 & w4169;
assign w4171 = ~w4161 & w4170;
assign w4172 = ~pi096 & ~w4154;
assign w4173 = w4171 & ~w4172;
assign w4174 = ~pi125 & w4138;
assign w4175 = w4124 & w4126;
assign w4176 = ~w4174 & ~w4175;
assign w4177 = ~pi113 & ~w4176;
assign w4178 = w4124 & w4144;
assign w4179 = ~pi009 & w4178;
assign w4180 = (pi096 & ~w4178) | (pi096 & w18328) | (~w4178 & w18328);
assign w4181 = pi113 & ~pi125;
assign w4182 = w4126 & w4181;
assign w4183 = pi025 & ~pi124;
assign w4184 = w4149 & w4183;
assign w4185 = ~w4177 & w4180;
assign w4186 = ~w4182 & ~w4184;
assign w4187 = w4185 & w4186;
assign w4188 = ~pi113 & pi124;
assign w4189 = pi025 & ~pi125;
assign w4190 = w4188 & w4189;
assign w4191 = ~pi096 & ~w4190;
assign w4192 = pi025 & pi124;
assign w4193 = pi009 & w4192;
assign w4194 = w4127 & w4162;
assign w4195 = w4137 & w4144;
assign w4196 = ~pi113 & w4195;
assign w4197 = pi025 & pi125;
assign w4198 = w4126 & w4197;
assign w4199 = pi113 & w4198;
assign w4200 = ~w4196 & ~w4199;
assign w4201 = ~w4193 & ~w4194;
assign w4202 = w4191 & w4201;
assign w4203 = w4200 & w4202;
assign w4204 = pi009 & ~pi025;
assign w4205 = w4126 & w4204;
assign w4206 = pi113 & ~w4205;
assign w4207 = ~pi009 & pi125;
assign w4208 = ~pi124 & w4207;
assign w4209 = w4162 & w4189;
assign w4210 = ~w4149 & ~w4208;
assign w4211 = w4206 & w4210;
assign w4212 = ~w4209 & w4211;
assign w4213 = pi009 & w4138;
assign w4214 = w4138 & w4127;
assign w4215 = w4162 & w4204;
assign w4216 = ~pi113 & ~w4215;
assign w4217 = w4145 & w4158;
assign w4218 = ~w4214 & w4216;
assign w4219 = ~w4217 & w4218;
assign w4220 = ~w4212 & ~w4219;
assign w4221 = ~pi010 & ~w4220;
assign w4222 = ~w4187 & ~w4203;
assign w4223 = w4221 & ~w4222;
assign w4224 = ~w4143 & w4173;
assign w4225 = ~w4223 & ~w4224;
assign w4226 = w4162 & w4166;
assign w4227 = ~pi125 & w4226;
assign w4228 = ~w4144 & w4204;
assign w4229 = ~w4217 & ~w4227;
assign w4230 = (~pi113 & ~w4229) | (~pi113 & w18329) | (~w4229 & w18329);
assign w4231 = pi009 & w4162;
assign w4232 = w4124 & w4231;
assign w4233 = ~pi025 & ~pi125;
assign w4234 = pi009 & w4126;
assign w4235 = w4233 & w4234;
assign w4236 = pi009 & pi113;
assign w4237 = pi025 & w4144;
assign w4238 = w4236 & w4237;
assign w4239 = ~w4232 & ~w4235;
assign w4240 = ~w4238 & w4239;
assign w4241 = pi009 & ~pi113;
assign w4242 = w4138 & w4233;
assign w4243 = w4146 & w4236;
assign w4244 = w4241 & w4242;
assign w4245 = ~w4243 & ~w4244;
assign w4246 = (pi096 & ~w4136) | (pi096 & w18330) | (~w4136 & w18330);
assign w4247 = w4245 & w4246;
assign w4248 = w4240 & w4247;
assign w4249 = ~w4230 & w4248;
assign w4250 = pi055 & w4155;
assign w4251 = w4207 & w4250;
assign w4252 = w4189 & w4231;
assign w4253 = ~pi009 & pi124;
assign w4254 = w4159 & w4253;
assign w4255 = ~w4251 & ~w4252;
assign w4256 = (~pi113 & ~w4255) | (~pi113 & w18331) | (~w4255 & w18331);
assign w4257 = pi009 & w4175;
assign w4258 = pi025 & ~pi055;
assign w4259 = w4127 & w4258;
assign w4260 = ~w4167 & ~w4259;
assign w4261 = ~w4257 & w4260;
assign w4262 = w4131 & w18332;
assign w4263 = ~pi025 & ~pi055;
assign w4264 = ~pi125 & w4263;
assign w4265 = w4253 & w4264;
assign w4266 = ~w4262 & ~w4265;
assign w4267 = w4261 & w4266;
assign w4268 = pi113 & ~w4267;
assign w4269 = w4197 & w4213;
assign w4270 = ~w4168 & ~w4269;
assign w4271 = w4245 & w4270;
assign w4272 = ~pi096 & w4271;
assign w4273 = ~w4256 & ~w4268;
assign w4274 = w4272 & w4273;
assign w4275 = ~w4249 & ~w4274;
assign w4276 = ~w4225 & ~w4275;
assign w4277 = ~pi185 & w4276;
assign w4278 = pi185 & ~w4276;
assign w4279 = ~w4277 & ~w4278;
assign w4280 = w4123 & w4279;
assign w4281 = ~w4123 & ~w4279;
assign w4282 = ~w4280 & ~w4281;
assign w4283 = ~w3879 & w4282;
assign w4284 = ~pi529 & ~w4283;
assign w4285 = w3879 & ~w4282;
assign w4286 = w4284 & ~w4285;
assign w4287 = ~pi185 & pi444;
assign w4288 = pi529 & ~w4287;
assign w4289 = pi185 & ~pi444;
assign w4290 = w4288 & ~w4289;
assign w4291 = ~w4286 & ~w4290;
assign w4292 = ~w3370 & ~w3925;
assign w4293 = pi122 & ~w4292;
assign w4294 = ~pi122 & ~w3384;
assign w4295 = ~w3952 & w4294;
assign w4296 = ~w3440 & ~w4295;
assign w4297 = ~w4293 & w4296;
assign w4298 = ~pi017 & ~w4297;
assign w4299 = ~w3481 & ~w3713;
assign w4300 = w3409 & w3387;
assign w4301 = ~w3713 & w18333;
assign w4302 = (pi039 & w4298) | (pi039 & w18334) | (w4298 & w18334);
assign w4303 = ~w3451 & ~w3760;
assign w4304 = ~w3905 & ~w3943;
assign w4305 = w4303 & w4304;
assign w4306 = pi122 & ~w3667;
assign w4307 = ~pi122 & w3437;
assign w4308 = w3370 & w3677;
assign w4309 = ~w4307 & ~w4308;
assign w4310 = w3401 & w4306;
assign w4311 = w4309 & ~w4310;
assign w4312 = (~pi039 & ~w4311) | (~pi039 & w18335) | (~w4311 & w18335);
assign w4313 = pi076 & ~w3692;
assign w4314 = ~w3386 & w4313;
assign w4315 = (pi122 & ~w3369) | (pi122 & w3696) | (~w3369 & w3696);
assign w4316 = pi039 & ~w4315;
assign w4317 = ~w3703 & ~w4314;
assign w4318 = (w4316 & ~w4317) | (w4316 & w18336) | (~w4317 & w18336);
assign w4319 = (w3464 & ~w3446) | (w3464 & w18337) | (~w3446 & w18337);
assign w4320 = ~pi043 & w3683;
assign w4321 = ~w3487 & ~w3946;
assign w4322 = ~w4320 & w4321;
assign w4323 = ~w4319 & w4322;
assign w4324 = ~w4318 & w4323;
assign w4325 = (pi017 & ~w4324) | (pi017 & w18338) | (~w4324 & w18338);
assign w4326 = ~w3678 & ~w3947;
assign w4327 = ~pi077 & ~w4326;
assign w4328 = ~pi122 & ~w3943;
assign w4329 = ~w3448 & w4328;
assign w4330 = ~w4327 & w4329;
assign w4331 = ~pi077 & w3667;
assign w4332 = w3496 & ~w4331;
assign w4333 = ~w3953 & w4332;
assign w4334 = ~w4330 & ~w4333;
assign w4335 = w3375 & ~w3387;
assign w4336 = w3384 & w3719;
assign w4337 = ~w3492 & ~w4336;
assign w4338 = ~pi039 & ~w4337;
assign w4339 = w3413 & w3394;
assign w4340 = ~pi076 & ~pi077;
assign w4341 = w4336 & w4340;
assign w4342 = ~w4338 & ~w4339;
assign w4343 = ~w3669 & ~w4341;
assign w4344 = ~w3396 & ~w3437;
assign w4345 = pi039 & ~w4344;
assign w4346 = ~w3487 & ~w3690;
assign w4347 = ~w4345 & w4346;
assign w4348 = pi039 & w3464;
assign w4349 = w3475 & w4348;
assign w4350 = ~w3746 & ~w4349;
assign w4351 = (w4350 & w4347) | (w4350 & w18339) | (w4347 & w18339);
assign w4352 = (~pi017 & ~w4342) | (~pi017 & w20767) | (~w4342 & w20767);
assign w4353 = w4351 & ~w4352;
assign w4354 = (~pi039 & w4334) | (~pi039 & w18340) | (w4334 & w18340);
assign w4355 = w4353 & ~w4354;
assign w4356 = ~w4302 & ~w4325;
assign w4357 = w4355 & w4356;
assign w4358 = ~w3519 & ~w3812;
assign w4359 = ~pi091 & w4358;
assign w4360 = pi005 & w3529;
assign w4361 = ~w3648 & ~w4360;
assign w4362 = w4359 & ~w4361;
assign w4363 = w3522 & w3550;
assign w4364 = ~w3525 & ~w4363;
assign w4365 = (~w3587 & w4364) | (~w3587 & w18341) | (w4364 & w18341);
assign w4366 = (pi024 & w4362) | (pi024 & w18342) | (w4362 & w18342);
assign w4367 = (~w3788 & ~w3532) | (~w3788 & w18343) | (~w3532 & w18343);
assign w4368 = w3570 & w3822;
assign w4369 = ~w3638 & ~w4368;
assign w4370 = pi084 & w3524;
assign w4371 = w3550 & w4370;
assign w4372 = ~pi024 & ~w4369;
assign w4373 = w4370 & w18344;
assign w4374 = ~w4372 & ~w4373;
assign w4375 = w4367 & w4374;
assign w4376 = ~w4366 & w4375;
assign w4377 = ~pi018 & ~w4376;
assign w4378 = ~pi005 & w3522;
assign w4379 = ~w3531 & ~w3778;
assign w4380 = (pi091 & ~w3522) | (pi091 & w3566) | (~w3522 & w3566);
assign w4381 = (~w4380 & ~w4379) | (~w4380 & w18345) | (~w4379 & w18345);
assign w4382 = w3560 & w3570;
assign w4383 = ~pi004 & pi091;
assign w4384 = w3533 & w4383;
assign w4385 = ~w3860 & ~w4382;
assign w4386 = ~w4384 & w4385;
assign w4387 = w3524 & w18346;
assign w4388 = ~w3777 & ~w4387;
assign w4389 = w4386 & w4388;
assign w4390 = (~pi024 & ~w4389) | (~pi024 & w18347) | (~w4389 & w18347);
assign w4391 = ~pi004 & w3524;
assign w4392 = (pi091 & ~w3524) | (pi091 & w3801) | (~w3524 & w3801);
assign w4393 = pi024 & ~w4392;
assign w4394 = (w4393 & ~w4359) | (w4393 & w18348) | (~w4359 & w18348);
assign w4395 = w3522 & w3530;
assign w4396 = w3524 & w3608;
assign w4397 = ~w3604 & ~w4395;
assign w4398 = (w3566 & ~w4397) | (w3566 & w18349) | (~w4397 & w18349);
assign w4399 = w3533 & w3546;
assign w4400 = ~pi005 & w4399;
assign w4401 = pi084 & w3778;
assign w4402 = w3547 & w3645;
assign w4403 = ~w4400 & ~w4401;
assign w4404 = ~w4402 & w4403;
assign w4405 = ~w4398 & w4404;
assign w4406 = ~w4394 & w4405;
assign w4407 = (pi018 & ~w4406) | (pi018 & w18350) | (~w4406 & w18350);
assign w4408 = w3533 & w3580;
assign w4409 = ~w3621 & ~w4408;
assign w4410 = ~w3602 & w4409;
assign w4411 = w3620 & w4360;
assign w4412 = ~pi052 & w3545;
assign w4413 = ~w3638 & ~w4412;
assign w4414 = ~w4411 & w4413;
assign w4415 = pi091 & ~w4414;
assign w4416 = w3518 & w3580;
assign w4417 = w3568 & w4370;
assign w4418 = ~w4417 & w18351;
assign w4419 = ~w4415 & w4418;
assign w4420 = (~pi024 & ~w4419) | (~pi024 & w18352) | (~w4419 & w18352);
assign w4421 = ~w3625 & ~w3817;
assign w4422 = ~pi005 & w3533;
assign w4423 = w3533 & w3543;
assign w4424 = ~w3771 & ~w4423;
assign w4425 = (pi024 & w3771) | (pi024 & w10858) | (w3771 & w10858);
assign w4426 = (w4425 & ~w4421) | (w4425 & w18353) | (~w4421 & w18353);
assign w4427 = w3630 & w3859;
assign w4428 = ~w3845 & ~w4427;
assign w4429 = pi091 & w3560;
assign w4430 = ~w3595 & ~w4370;
assign w4431 = w4429 & ~w4430;
assign w4432 = ~pi005 & w3593;
assign w4433 = ~w3531 & ~w4432;
assign w4434 = w3858 & ~w4433;
assign w4435 = ~w4431 & ~w4434;
assign w4436 = w4428 & w4435;
assign w4437 = ~w4426 & w4436;
assign w4438 = ~w4420 & w4437;
assign w4439 = ~w4377 & ~w4407;
assign w4440 = w4438 & w4439;
assign w4441 = ~w4357 & w4440;
assign w4442 = w4357 & ~w4440;
assign w4443 = ~w4441 & ~w4442;
assign w4444 = w3663 & ~w4443;
assign w4445 = ~w3663 & w4443;
assign w4446 = ~w4444 & ~w4445;
assign w4447 = w3971 & w4003;
assign w4448 = pi037 & w4037;
assign w4449 = ~w4088 & ~w4447;
assign w4450 = ~w4056 & ~w4073;
assign w4451 = w3971 & w4035;
assign w4452 = w3988 & w4059;
assign w4453 = ~w4099 & ~w4451;
assign w4454 = w4450 & w4453;
assign w4455 = ~w4452 & w4454;
assign w4456 = w3973 & w4010;
assign w4457 = ~w3994 & ~w4456;
assign w4458 = ~pi106 & w4457;
assign w4459 = ~w4000 & ~w4045;
assign w4460 = w4066 & w4459;
assign w4461 = ~w4458 & ~w4460;
assign w4462 = w3971 & w3978;
assign w4463 = w3978 & w4031;
assign w4464 = ~w4462 & ~w4463;
assign w4465 = ~w3984 & w4464;
assign w4466 = w3978 & w3981;
assign w4467 = pi037 & ~pi100;
assign w4468 = w3988 & w4467;
assign w4469 = pi128 & w4468;
assign w4470 = w3992 & w18356;
assign w4471 = ~w4469 & ~w4470;
assign w4472 = ~w4469 & w18357;
assign w4473 = ~pi106 & ~w4472;
assign w4474 = pi035 & w4037;
assign w4475 = ~w3973 & ~w4037;
assign w4476 = ~pi037 & ~w4475;
assign w4477 = (w4032 & w4476) | (w4032 & w18358) | (w4476 & w18358);
assign w4478 = w3973 & w4082;
assign w4479 = ~w4477 & ~w4478;
assign w4480 = ~w4473 & w4479;
assign w4481 = (~pi065 & w4461) | (~pi065 & w18359) | (w4461 & w18359);
assign w4482 = w4480 & ~w4481;
assign w4483 = (pi068 & ~w4482) | (pi068 & w18360) | (~w4482 & w18360);
assign w4484 = ~pi037 & ~pi128;
assign w4485 = ~pi031 & w4484;
assign w4486 = pi037 & ~pi128;
assign w4487 = pi100 & w3988;
assign w4488 = w4486 & w4487;
assign w4489 = w3982 & w4059;
assign w4490 = pi100 & w4489;
assign w4491 = w4060 & w4448;
assign w4492 = ~w4490 & ~w4491;
assign w4493 = ~w4008 & ~w4065;
assign w4494 = w4492 & w4493;
assign w4495 = ~w3977 & w4021;
assign w4496 = pi128 & w4495;
assign w4497 = ~w4466 & ~w4496;
assign w4498 = pi037 & ~pi106;
assign w4499 = w4053 & w4056;
assign w4500 = w4052 & ~w4498;
assign w4501 = ~w4499 & ~w4500;
assign w4502 = w4497 & w4501;
assign w4503 = ~pi065 & ~w4502;
assign w4504 = w4059 & w4487;
assign w4505 = ~w4090 & ~w4504;
assign w4506 = ~pi031 & w4015;
assign w4507 = pi106 & w4069;
assign w4508 = w3973 & w3978;
assign w4509 = ~pi037 & w4508;
assign w4510 = ~w4507 & ~w4509;
assign w4511 = w4484 & w4506;
assign w4512 = w4510 & ~w4511;
assign w4513 = (~pi106 & w4504) | (~pi106 & w18363) | (w4504 & w18363);
assign w4514 = w4512 & ~w4513;
assign w4515 = ~w4503 & w4514;
assign w4516 = (~pi068 & ~w4515) | (~pi068 & w18364) | (~w4515 & w18364);
assign w4517 = w3995 & w4031;
assign w4518 = (pi106 & ~w4450) | (pi106 & w20768) | (~w4450 & w20768);
assign w4519 = w4037 & w4044;
assign w4520 = pi031 & w3977;
assign w4521 = ~w4034 & ~w4519;
assign w4522 = (w4098 & ~w4521) | (w4098 & w18365) | (~w4521 & w18365);
assign w4523 = ~pi106 & w4065;
assign w4524 = w4065 & w4060;
assign w4525 = (pi065 & ~w18366) | (pi065 & w20769) | (~w18366 & w20769);
assign w4526 = ~pi065 & pi106;
assign w4527 = ~w4042 & ~w4509;
assign w4528 = w4526 & ~w4527;
assign w4529 = ~pi065 & ~pi106;
assign w4530 = w3973 & w4018;
assign w4531 = pi035 & w4530;
assign w4532 = ~w4106 & ~w4520;
assign w4533 = w3981 & w4015;
assign w4534 = ~w4532 & w4533;
assign w4535 = w4058 & w4529;
assign w4536 = ~w4534 & w18367;
assign w4537 = ~w4528 & w4536;
assign w4538 = ~w4525 & w4537;
assign w4539 = ~w4516 & w4538;
assign w4540 = ~w4483 & w4539;
assign w4541 = ~w3770 & w4540;
assign w4542 = w3770 & ~w4540;
assign w4543 = ~w4541 & ~w4542;
assign w4544 = pi125 & w4134;
assign w4545 = ~pi055 & w4166;
assign w4546 = pi025 & w4126;
assign w4547 = ~w4544 & ~w4545;
assign w4548 = ~pi009 & w4138;
assign w4549 = ~w4145 & ~w4548;
assign w4550 = ~pi113 & ~w4549;
assign w4551 = ~w4198 & ~w4215;
assign w4552 = w4192 & w4207;
assign w4553 = w4551 & ~w4552;
assign w4554 = ~w4550 & w4553;
assign w4555 = w4134 & w4150;
assign w4556 = pi055 & w4555;
assign w4557 = ~w4125 & w4205;
assign w4558 = ~w4133 & ~w4557;
assign w4559 = w4138 & w4204;
assign w4560 = w4131 & w4158;
assign w4561 = w4144 & w4158;
assign w4562 = ~w4560 & ~w4561;
assign w4563 = w4181 & w4183;
assign w4564 = w4562 & ~w4563;
assign w4565 = ~w4206 & w4559;
assign w4566 = w4564 & ~w4565;
assign w4567 = ~w4556 & w4558;
assign w4568 = w4566 & w4567;
assign w4569 = ~pi096 & ~w4568;
assign w4570 = pi125 & w4258;
assign w4571 = w4253 & w4570;
assign w4572 = pi009 & pi025;
assign w4573 = w4162 & w4572;
assign w4574 = w4134 & w4158;
assign w4575 = ~w4573 & ~w4574;
assign w4576 = ~w4571 & w4575;
assign w4577 = ~pi113 & ~w4576;
assign w4578 = w4189 & w4213;
assign w4579 = ~w4126 & ~w4138;
assign w4580 = ~pi025 & ~w4579;
assign w4581 = (w4135 & w4580) | (w4135 & w18369) | (w4580 & w18369);
assign w4582 = ~w4577 & w18370;
assign w4583 = ~pi125 & w4155;
assign w4584 = w4197 & w4548;
assign w4585 = (pi113 & w4584) | (pi113 & w18372) | (w4584 & w18372);
assign w4586 = pi055 & w4192;
assign w4587 = w4137 & w4586;
assign w4588 = w4126 & w4189;
assign w4589 = ~pi113 & w4588;
assign w4590 = ~w4587 & ~w4589;
assign w4591 = pi096 & ~w4205;
assign w4592 = ~w4227 & w4591;
assign w4593 = w4590 & w4592;
assign w4594 = ~pi009 & pi113;
assign w4595 = ~w4263 & w4594;
assign w4596 = pi124 & w4595;
assign w4597 = ~pi096 & ~w4574;
assign w4598 = ~w4596 & w4597;
assign w4599 = ~w4124 & ~w4135;
assign w4600 = w4144 & ~w4599;
assign w4601 = w4198 & w4241;
assign w4602 = ~w4600 & ~w4601;
assign w4603 = w4598 & w4602;
assign w4604 = ~w4585 & w4593;
assign w4605 = ~w4603 & ~w4604;
assign w4606 = pi055 & w4207;
assign w4607 = w4192 & w4606;
assign w4608 = ~w4139 & ~w4607;
assign w4609 = pi113 & w4209;
assign w4610 = ~pi124 & w4160;
assign w4611 = ~w4609 & ~w4610;
assign w4612 = w4236 & w4583;
assign w4613 = w4611 & ~w4612;
assign w4614 = (~pi113 & w4607) | (~pi113 & w18373) | (w4607 & w18373);
assign w4615 = (pi010 & w4605) | (pi010 & w18374) | (w4605 & w18374);
assign w4616 = w4127 & w4131;
assign w4617 = (pi113 & ~w4551) | (pi113 & w20770) | (~w4551 & w20770);
assign w4618 = pi125 & w4263;
assign w4619 = ~w4174 & ~w4588;
assign w4620 = (w4150 & ~w4619) | (w4150 & w18375) | (~w4619 & w18375);
assign w4621 = ~pi125 & w4134;
assign w4622 = w4241 & w4621;
assign w4623 = w4621 & w18376;
assign w4624 = (pi096 & ~w18377) | (pi096 & w20771) | (~w18377 & w20771);
assign w4625 = ~pi113 & w4162;
assign w4626 = ~pi096 & ~pi125;
assign w4627 = w4124 & w4138;
assign w4628 = pi113 & w4175;
assign w4629 = ~w4627 & ~w4628;
assign w4630 = w4625 & w4626;
assign w4631 = ~pi025 & pi113;
assign w4632 = ~pi096 & pi113;
assign w4633 = ~w4179 & ~w4610;
assign w4634 = w4194 & w4631;
assign w4635 = (~w4634 & w4633) | (~w4634 & w18378) | (w4633 & w18378);
assign w4636 = (pi009 & ~w4629) | (pi009 & w20772) | (~w4629 & w20772);
assign w4637 = w4635 & ~w4636;
assign w4638 = ~w4624 & w4637;
assign w4639 = ~w4615 & w4638;
assign w4640 = (w4569 & w20773) | (w4569 & w20774) | (w20773 & w20774);
assign w4641 = w4639 & ~w4640;
assign w4642 = w4639 & w20775;
assign w4643 = (pi138 & ~w4639) | (pi138 & w20776) | (~w4639 & w20776);
assign w4644 = ~w4642 & ~w4643;
assign w4645 = w4543 & w4644;
assign w4646 = ~w4543 & ~w4644;
assign w4647 = ~w4645 & ~w4646;
assign w4648 = ~w4446 & w4647;
assign w4649 = ~pi529 & ~w4648;
assign w4650 = w4446 & ~w4647;
assign w4651 = w4649 & ~w4650;
assign w4652 = ~pi138 & pi517;
assign w4653 = pi529 & ~w4652;
assign w4654 = pi138 & ~pi517;
assign w4655 = w4653 & ~w4654;
assign w4656 = ~w4651 & ~w4655;
assign w4657 = pi055 & ~pi125;
assign w4658 = ~pi009 & w4144;
assign w4659 = ~w4213 & ~w4618;
assign w4660 = ~w4657 & ~w4658;
assign w4661 = w4659 & w4660;
assign w4662 = ~pi125 & w4253;
assign w4663 = w4207 & w4258;
assign w4664 = w4138 & w4197;
assign w4665 = ~w4663 & ~w4664;
assign w4666 = w4253 & w4657;
assign w4667 = pi096 & ~w4661;
assign w4668 = pi009 & w4233;
assign w4669 = w4138 & ~w4668;
assign w4670 = ~w4146 & ~w4618;
assign w4671 = ~w4669 & w4670;
assign w4672 = ~pi113 & ~w4671;
assign w4673 = w4594 & w4621;
assign w4674 = w4138 & w4207;
assign w4675 = ~w4259 & ~w4674;
assign w4676 = ~w4673 & w4675;
assign w4677 = ~pi025 & w4150;
assign w4678 = w4126 & w4677;
assign w4679 = ~w4232 & ~w4678;
assign w4680 = pi009 & w4159;
assign w4681 = w4183 & w4207;
assign w4682 = w4181 & w4680;
assign w4683 = ~w4681 & ~w4682;
assign w4684 = ~pi113 & w4674;
assign w4685 = w4683 & ~w4684;
assign w4686 = pi096 & ~w4679;
assign w4687 = w4685 & ~w4686;
assign w4688 = (~pi096 & w4672) | (~pi096 & w18380) | (w4672 & w18380);
assign w4689 = w4687 & ~w4688;
assign w4690 = ~w4156 & ~w4559;
assign w4691 = ~pi113 & ~w4690;
assign w4692 = w4126 & w4572;
assign w4693 = pi055 & w4124;
assign w4694 = ~w4253 & ~w4594;
assign w4695 = w4693 & ~w4694;
assign w4696 = ~w4692 & ~w4695;
assign w4697 = ~w4691 & w4696;
assign w4698 = pi096 & ~w4697;
assign w4699 = (w4626 & w4193) | (w4626 & w18382) | (w4193 & w18382);
assign w4700 = w4162 & w4197;
assign w4701 = w4144 & w4197;
assign w4702 = ~w4700 & ~w4701;
assign w4703 = w4236 & ~w4702;
assign w4704 = pi124 & w4137;
assign w4705 = ~w4144 & ~w4704;
assign w4706 = pi009 & w4181;
assign w4707 = w4144 & w4706;
assign w4708 = (w4632 & w4704) | (w4632 & w18383) | (w4704 & w18383);
assign w4709 = ~w4707 & ~w4708;
assign w4710 = w4158 & w4183;
assign w4711 = ~w4226 & ~w4710;
assign w4712 = ~w4269 & w4711;
assign w4713 = (~pi113 & ~w4712) | (~pi113 & w18384) | (~w4712 & w18384);
assign w4714 = ~pi025 & ~w4709;
assign w4715 = ~w4713 & ~w4714;
assign w4716 = ~w4699 & ~w4703;
assign w4717 = ~w4698 & w4716;
assign w4718 = w4131 & w4207;
assign w4719 = w4144 & w4204;
assign w4720 = ~w4232 & w18385;
assign w4721 = pi113 & ~w4720;
assign w4722 = ~pi113 & ~w4711;
assign w4723 = ~w4552 & ~w4622;
assign w4724 = ~w4722 & w4723;
assign w4725 = ~w4721 & w4724;
assign w4726 = pi096 & pi113;
assign w4727 = ~w4175 & ~w4209;
assign w4728 = ~pi009 & ~w4727;
assign w4729 = w4162 & w4233;
assign w4730 = ~w4168 & ~w4262;
assign w4731 = ~w4728 & w4730;
assign w4732 = w4132 & w4158;
assign w4733 = ~w4157 & ~w4732;
assign w4734 = ~pi113 & ~w4733;
assign w4735 = ~w4209 & ~w4242;
assign w4736 = ~w4237 & ~w4570;
assign w4737 = w4735 & w4736;
assign w4738 = pi096 & ~pi113;
assign w4739 = pi009 & w4738;
assign w4740 = ~w4737 & w4739;
assign w4741 = ~w4734 & ~w4740;
assign w4742 = (w4726 & ~w4731) | (w4726 & w18386) | (~w4731 & w18386);
assign w4743 = w4741 & ~w4742;
assign w4744 = ~pi096 & ~w4725;
assign w4745 = w4743 & ~w4744;
assign w4746 = (pi010 & ~w4717) | (pi010 & w18387) | (~w4717 & w18387);
assign w4747 = w4745 & ~w4746;
assign w4748 = (~pi010 & ~w4689) | (~pi010 & w18388) | (~w4689 & w18388);
assign w4749 = w4747 & ~w4748;
assign w4750 = w4747 & w18389;
assign w4751 = (pi191 & ~w4747) | (pi191 & w18390) | (~w4747 & w18390);
assign w4752 = ~w4750 & ~w4751;
assign w4753 = w3524 & w3534;
assign w4754 = (pi091 & ~w18391) | (pi091 & w20777) | (~w18391 & w20777);
assign w4755 = w3593 & w3647;
assign w4756 = ~w3639 & ~w4382;
assign w4757 = ~w4755 & w4756;
assign w4758 = w3535 & w18392;
assign w4759 = w4757 & ~w4758;
assign w4760 = (~pi024 & ~w4759) | (~pi024 & w20778) | (~w4759 & w20778);
assign w4761 = (pi024 & w3597) | (pi024 & w18393) | (w3597 & w18393);
assign w4762 = ~w3565 & ~w3609;
assign w4763 = w3529 & w3608;
assign w4764 = ~w3571 & ~w4763;
assign w4765 = ~w4761 & w4764;
assign w4766 = (~pi091 & ~w4765) | (~pi091 & w18394) | (~w4765 & w18394);
assign w4767 = w3550 & w3631;
assign w4768 = w3570 & w3581;
assign w4769 = ~w4767 & ~w4768;
assign w4770 = ~w3795 & ~w4399;
assign w4771 = w4769 & w4770;
assign w4772 = pi091 & ~w4771;
assign w4773 = pi024 & w4395;
assign w4774 = w3522 & w18346;
assign w4775 = w3550 & w3802;
assign w4776 = ~w4773 & ~w4774;
assign w4777 = ~w4775 & w4776;
assign w4778 = ~w4772 & w18395;
assign w4779 = (pi018 & ~w4778) | (pi018 & w20779) | (~w4778 & w20779);
assign w4780 = pi094 & w3580;
assign w4781 = ~w3777 & ~w4780;
assign w4782 = w3623 & ~w4781;
assign w4783 = w3568 & w3595;
assign w4784 = ~w3525 & ~w4391;
assign w4785 = ~w4783 & w4784;
assign w4786 = ~w4782 & w4785;
assign w4787 = w3524 & w3580;
assign w4788 = ~pi091 & w4787;
assign w4789 = ~pi005 & ~w3633;
assign w4790 = w3518 & w3560;
assign w4791 = ~w3797 & ~w4790;
assign w4792 = ~w3795 & w4791;
assign w4793 = ~pi091 & ~w4792;
assign w4794 = ~w3565 & ~w4370;
assign w4795 = w3567 & ~w4794;
assign w4796 = ~w3623 & w3631;
assign w4797 = w3652 & w4796;
assign w4798 = ~w4795 & ~w4797;
assign w4799 = ~w4793 & w4798;
assign w4800 = (~pi024 & w4789) | (~pi024 & w18396) | (w4789 & w18396);
assign w4801 = w4799 & ~w4800;
assign w4802 = ~w3807 & ~w4401;
assign w4803 = (~pi091 & ~w4802) | (~pi091 & w18397) | (~w4802 & w18397);
assign w4804 = ~w3535 & ~w3539;
assign w4805 = w4429 & ~w4804;
assign w4806 = ~pi052 & w3566;
assign w4807 = w3570 & w4806;
assign w4808 = w4806 & w18398;
assign w4809 = ~w4805 & ~w4808;
assign w4810 = ~w4803 & w4809;
assign w4811 = ~pi024 & ~w4810;
assign w4812 = w3588 & w3803;
assign w4813 = w3566 & w3802;
assign w4814 = w3560 & w3597;
assign w4815 = ~w4813 & ~w4814;
assign w4816 = ~pi091 & w3638;
assign w4817 = w4815 & ~w4816;
assign w4818 = ~w4371 & ~w4812;
assign w4819 = (pi024 & ~w4817) | (pi024 & w18399) | (~w4817 & w18399);
assign w4820 = w3580 & w3640;
assign w4821 = w3645 & w18400;
assign w4822 = pi052 & w4820;
assign w4823 = ~w4821 & ~w4822;
assign w4824 = ~w4819 & w4823;
assign w4825 = ~w4811 & w4824;
assign w4826 = (~pi018 & ~w4801) | (~pi018 & w18401) | (~w4801 & w18401);
assign w4827 = w4825 & ~w4826;
assign w4828 = ~w4779 & w4827;
assign w4829 = ~w3660 & w4828;
assign w4830 = w3660 & ~w4828;
assign w4831 = ~w4829 & ~w4830;
assign w4832 = w3977 & w4067;
assign w4833 = w3973 & w4055;
assign w4834 = w3992 & w4018;
assign w4835 = ~w4832 & ~w4833;
assign w4836 = (pi106 & ~w4835) | (pi106 & w18402) | (~w4835 & w18402);
assign w4837 = w3993 & w4037;
assign w4838 = pi031 & ~pi106;
assign w4839 = w3978 & w4486;
assign w4840 = ~pi031 & ~pi037;
assign w4841 = pi035 & w4840;
assign w4842 = w3995 & w4037;
assign w4843 = ~w4839 & ~w4841;
assign w4844 = ~w4842 & w4843;
assign w4845 = w4837 & w4838;
assign w4846 = w4844 & ~w4845;
assign w4847 = (~pi065 & ~w4846) | (~pi065 & w18403) | (~w4846 & w18403);
assign w4848 = w3983 & w4486;
assign w4849 = ~w4469 & ~w4848;
assign w4850 = ~pi031 & w3981;
assign w4851 = w3981 & w18404;
assign w4852 = w3995 & w4059;
assign w4853 = ~w4851 & ~w4852;
assign w4854 = (pi106 & ~w4849) | (pi106 & w18405) | (~w4849 & w18405);
assign w4855 = w3992 & w4055;
assign w4856 = pi035 & w3989;
assign w4857 = w3988 & w4486;
assign w4858 = ~w4096 & ~w4855;
assign w4859 = ~w4856 & ~w4857;
assign w4860 = w4858 & w4859;
assign w4861 = ~pi106 & w4031;
assign w4862 = ~w4530 & ~w4861;
assign w4863 = (pi065 & ~w4862) | (pi065 & w18406) | (~w4862 & w18406);
assign w4864 = w3973 & w4003;
assign w4865 = ~w4014 & ~w4864;
assign w4866 = ~w4863 & w4865;
assign w4867 = ~pi106 & ~w4860;
assign w4868 = w4866 & ~w4867;
assign w4869 = ~w4847 & w4868;
assign w4870 = (pi068 & ~w4869) | (pi068 & w18407) | (~w4869 & w18407);
assign w4871 = (~pi106 & ~w4471) | (~pi106 & w18408) | (~w4471 & w18408);
assign w4872 = w3973 & w4840;
assign w4873 = ~w4069 & ~w4872;
assign w4874 = ~pi035 & ~w4873;
assign w4875 = w4054 & ~w4874;
assign w4876 = w3981 & w4098;
assign w4877 = w3982 & w3992;
assign w4878 = (pi065 & ~w3971) | (pi065 & w18409) | (~w3971 & w18409);
assign w4879 = w4000 & w4015;
assign w4880 = w4878 & ~w4879;
assign w4881 = ~w3972 & ~w4876;
assign w4882 = ~w4877 & w4881;
assign w4883 = w4880 & w4882;
assign w4884 = ~w4875 & ~w4883;
assign w4885 = w3992 & w4003;
assign w4886 = ~w4448 & ~w4885;
assign w4887 = w4526 & ~w4886;
assign w4888 = ~w3989 & ~w4016;
assign w4889 = w4506 & ~w4888;
assign w4890 = ~w4887 & ~w4889;
assign w4891 = ~w4884 & w18410;
assign w4892 = ~w4044 & w4067;
assign w4893 = pi100 & w4892;
assign w4894 = ~w4004 & ~w4893;
assign w4895 = (pi106 & w3980) | (pi106 & w18411) | (w3980 & w18411);
assign w4896 = w3973 & w4044;
assign w4897 = w4053 & w4896;
assign w4898 = w3971 & w4055;
assign w4899 = w4015 & w4898;
assign w4900 = ~w4897 & ~w4899;
assign w4901 = ~w4895 & w4900;
assign w4902 = ~pi106 & ~w4894;
assign w4903 = w4901 & ~w4902;
assign w4904 = pi100 & w4839;
assign w4905 = w3990 & w18412;
assign w4906 = ~w4904 & ~w4905;
assign w4907 = ~pi037 & w3969;
assign w4908 = ~w4452 & ~w4907;
assign w4909 = ~w4498 & ~w4533;
assign w4910 = ~w4908 & ~w4909;
assign w4911 = ~w4009 & ~w4046;
assign w4912 = ~w4910 & w4911;
assign w4913 = ~pi106 & w4877;
assign w4914 = (~w4913 & w4912) | (~w4913 & w18413) | (w4912 & w18413);
assign w4915 = pi106 & ~w4906;
assign w4916 = w4914 & ~w4915;
assign w4917 = ~pi065 & ~w4903;
assign w4918 = w4916 & ~w4917;
assign w4919 = ~pi068 & ~w4891;
assign w4920 = w4918 & ~w4919;
assign w4921 = ~w4870 & w4920;
assign w4922 = w3369 & w3410;
assign w4923 = ~w3385 & ~w3437;
assign w4924 = (pi122 & ~w4923) | (pi122 & w18414) | (~w4923 & w18414);
assign w4925 = ~pi122 & w3485;
assign w4926 = pi070 & ~w3409;
assign w4927 = w3397 & ~w4926;
assign w4928 = ~w3451 & ~w4927;
assign w4929 = ~w4925 & w4928;
assign w4930 = (~pi039 & ~w4929) | (~pi039 & w18415) | (~w4929 & w18415);
assign w4931 = w3397 & w3491;
assign w4932 = w3384 & w3431;
assign w4933 = ~w4931 & ~w4932;
assign w4934 = ~w3691 & ~w3745;
assign w4935 = w4933 & w4934;
assign w4936 = (~pi122 & w3458) | (~pi122 & w18416) | (w3458 & w18416);
assign w4937 = (pi039 & w4936) | (pi039 & w18417) | (w4936 & w18417);
assign w4938 = ~w3419 & ~w3474;
assign w4939 = pi043 & ~w4938;
assign w4940 = w3371 & w3491;
assign w4941 = ~w3421 & ~w4940;
assign w4942 = ~w4939 & w4941;
assign w4943 = ~pi122 & ~w4942;
assign w4944 = w3401 & w3449;
assign w4945 = ~w3880 & ~w4944;
assign w4946 = ~w4943 & w18418;
assign w4947 = ~w4930 & w4946;
assign w4948 = (pi017 & ~w4947) | (pi017 & w18419) | (~w4947 & w18419);
assign w4949 = ~pi043 & ~w3476;
assign w4950 = ~w3419 & ~w3486;
assign w4951 = w3420 & ~w4950;
assign w4952 = w3459 & w3491;
assign w4953 = ~w3692 & w4952;
assign w4954 = ~w4951 & ~w4953;
assign w4955 = (~pi039 & w4949) | (~pi039 & w18420) | (w4949 & w18420);
assign w4956 = w4954 & ~w4955;
assign w4957 = w3410 & w4340;
assign w4958 = ~w3691 & w18421;
assign w4959 = ~pi122 & ~w4958;
assign w4960 = w3391 & w3418;
assign w4961 = ~w3923 & ~w4960;
assign w4962 = ~w3370 & ~w3413;
assign w4963 = w4961 & w4962;
assign w4964 = (pi039 & ~w4963) | (pi039 & w18422) | (~w4963 & w18422);
assign w4965 = ~w4959 & ~w4964;
assign w4966 = w4956 & w4965;
assign w4967 = ~pi017 & ~w4966;
assign w4968 = w3486 & w18423;
assign w4969 = ~w3487 & ~w3703;
assign w4970 = (~pi122 & ~w4969) | (~pi122 & w18424) | (~w4969 & w18424);
assign w4971 = (~pi039 & w4970) | (~pi039 & w18425) | (w4970 & w18425);
assign w4972 = (w3394 & w3406) | (w3394 & w18426) | (w3406 & w18426);
assign w4973 = ~pi122 & w3492;
assign w4974 = ~w3904 & ~w3924;
assign w4975 = ~w4973 & w4974;
assign w4976 = (pi039 & ~w4975) | (pi039 & w18427) | (~w4975 & w18427);
assign w4977 = (w3459 & w3946) | (w3459 & w18428) | (w3946 & w18428);
assign w4978 = ~pi122 & w3413;
assign w4979 = w3404 & w4944;
assign w4980 = ~w4978 & ~w4979;
assign w4981 = ~w4977 & w4980;
assign w4982 = ~w4976 & w4981;
assign w4983 = ~w4971 & w4982;
assign w4984 = ~w4967 & w4983;
assign w4985 = ~w4948 & w4984;
assign w4986 = ~w4921 & w4985;
assign w4987 = w4921 & ~w4985;
assign w4988 = ~w4986 & ~w4987;
assign w4989 = w4831 & ~w4988;
assign w4990 = ~w4831 & w4988;
assign w4991 = ~w4989 & ~w4990;
assign w4992 = (~pi529 & w4991) | (~pi529 & w18429) | (w4991 & w18429);
assign w4993 = ~w4752 & w4991;
assign w4994 = w4992 & ~w4993;
assign w4995 = pi191 & pi405;
assign w4996 = pi529 & ~w4995;
assign w4997 = ~pi191 & ~pi405;
assign w4998 = w4996 & ~w4997;
assign w4999 = ~w4994 & ~w4998;
assign w5000 = pi111 & w294;
assign w5001 = ~w266 & ~w1397;
assign w5002 = ~pi123 & w299;
assign w5003 = ~w312 & ~w334;
assign w5004 = ~w354 & ~w1109;
assign w5005 = w5003 & w5004;
assign w5006 = ~w5002 & w5005;
assign w5007 = ~pi023 & w285;
assign w5008 = ~w345 & ~w5007;
assign w5009 = pi123 & w5008;
assign w5010 = ~w278 & ~w1064;
assign w5011 = ~pi123 & w5010;
assign w5012 = ~w5009 & ~w5011;
assign w5013 = ~w318 & w324;
assign w5014 = ~w1273 & ~w1385;
assign w5015 = ~w5013 & w5014;
assign w5016 = (~w1040 & w1241) | (~w1040 & w18432) | (w1241 & w18432);
assign w5017 = ~pi123 & ~w5016;
assign w5018 = ~w389 & ~w1259;
assign w5019 = (w1431 & ~w5018) | (w1431 & w18433) | (~w5018 & w18433);
assign w5020 = w261 & w345;
assign w5021 = ~w5019 & ~w5020;
assign w5022 = ~w5017 & w5021;
assign w5023 = (~pi048 & w5012) | (~pi048 & w18434) | (w5012 & w18434);
assign w5024 = w5022 & ~w5023;
assign w5025 = (pi020 & ~w5024) | (pi020 & w18435) | (~w5024 & w18435);
assign w5026 = w270 & w345;
assign w5027 = ~pi111 & w281;
assign w5028 = w282 & w314;
assign w5029 = ~pi123 & w5028;
assign w5030 = ~w1391 & ~w5029;
assign w5031 = ~w324 & ~w378;
assign w5032 = w5030 & w5031;
assign w5033 = ~w295 & ~w1431;
assign w5034 = w252 & ~w5033;
assign w5035 = w312 & w394;
assign w5036 = ~w257 & w343;
assign w5037 = pi093 & w5036;
assign w5038 = ~w5035 & ~w5037;
assign w5039 = ~w1040 & ~w5034;
assign w5040 = w5038 & w5039;
assign w5041 = ~pi048 & ~w5040;
assign w5042 = pi023 & w1085;
assign w5043 = ~w347 & ~w5042;
assign w5044 = (~pi123 & w5042) | (~pi123 & w18437) | (w5042 & w18437);
assign w5045 = w261 & w1063;
assign w5046 = ~w327 & ~w5045;
assign w5047 = pi123 & ~w5046;
assign w5048 = ~w1260 & ~w5047;
assign w5049 = ~w5044 & w5048;
assign w5050 = ~w5041 & w5049;
assign w5051 = ~w293 & ~w1023;
assign w5052 = (w353 & ~w5051) | (w353 & w18439) | (~w5051 & w18439);
assign w5053 = ~pi047 & w379;
assign w5054 = w1071 & w5053;
assign w5055 = ~w313 & ~w5054;
assign w5056 = ~w5052 & w5055;
assign w5057 = pi048 & ~w5056;
assign w5058 = ~pi048 & ~pi123;
assign w5059 = ~w1378 & ~w1432;
assign w5060 = w316 & w5058;
assign w5061 = w359 & w18440;
assign w5062 = w5059 & w18441;
assign w5063 = w261 & w326;
assign w5064 = ~w334 & ~w5063;
assign w5065 = (w1426 & w1078) | (w1426 & w18442) | (w1078 & w18442);
assign w5066 = w1416 & ~w5064;
assign w5067 = ~w5065 & ~w5066;
assign w5068 = w5062 & w5067;
assign w5069 = ~w5057 & w5068;
assign w5070 = (~pi020 & ~w5050) | (~pi020 & w18443) | (~w5050 & w18443);
assign w5071 = w5069 & ~w5070;
assign w5072 = ~w5025 & w5071;
assign w5073 = ~pi013 & ~pi054;
assign w5074 = w428 & w5073;
assign w5075 = ~w917 & ~w5074;
assign w5076 = ~pi114 & ~w5075;
assign w5077 = ~pi007 & w415;
assign w5078 = ~w457 & ~w5077;
assign w5079 = ~w487 & w1182;
assign w5080 = ~w5076 & w5079;
assign w5081 = ~pi013 & w971;
assign w5082 = ~w466 & ~w971;
assign w5083 = pi098 & ~w5082;
assign w5084 = ~w446 & ~w971;
assign w5085 = ~w426 & ~w449;
assign w5086 = ~w1004 & w5085;
assign w5087 = ~pi098 & ~pi114;
assign w5088 = w5084 & w5087;
assign w5089 = w5086 & ~w5088;
assign w5090 = (pi001 & ~w5089) | (pi001 & w18445) | (~w5089 & w18445);
assign w5091 = ~w963 & ~w1171;
assign w5092 = ~w1148 & w5091;
assign w5093 = ~pi114 & ~w5092;
assign w5094 = ~w507 & ~w920;
assign w5095 = pi013 & w417;
assign w5096 = (w476 & ~w5094) | (w476 & w18446) | (~w5094 & w18446);
assign w5097 = ~w5093 & w18447;
assign w5098 = ~w5090 & w5097;
assign w5099 = ~pi054 & w445;
assign w5100 = w451 & w475;
assign w5101 = w541 & w971;
assign w5102 = w475 & w1160;
assign w5103 = ~pi114 & w5101;
assign w5104 = ~w5102 & ~w5103;
assign w5105 = ~w457 & ~w532;
assign w5106 = w5104 & w5105;
assign w5107 = ~w466 & ~w476;
assign w5108 = w408 & ~w5107;
assign w5109 = ~pi013 & pi114;
assign w5110 = pi013 & ~pi114;
assign w5111 = w426 & w5110;
assign w5112 = ~w405 & w5109;
assign w5113 = pi098 & w5112;
assign w5114 = ~w5111 & ~w5113;
assign w5115 = ~w963 & ~w5108;
assign w5116 = w5114 & w5115;
assign w5117 = ~pi001 & ~w5116;
assign w5118 = pi098 & w1012;
assign w5119 = pi114 & w454;
assign w5120 = w404 & w5073;
assign w5121 = ~w5119 & ~w5120;
assign w5122 = w536 & w5099;
assign w5123 = w5121 & ~w5122;
assign w5124 = (~pi114 & w5118) | (~pi114 & w18450) | (w5118 & w18450);
assign w5125 = w5123 & ~w5124;
assign w5126 = ~w5117 & w5125;
assign w5127 = (~pi029 & ~w5126) | (~pi029 & w18451) | (~w5126 & w18451);
assign w5128 = (w479 & ~w407) | (w479 & w18452) | (~w407 & w18452);
assign w5129 = w436 & w457;
assign w5130 = ~w427 & ~w5129;
assign w5131 = ~w5128 & w5130;
assign w5132 = pi001 & ~w5131;
assign w5133 = w516 & w5109;
assign w5134 = ~w412 & ~w5133;
assign w5135 = w1011 & ~w5134;
assign w5136 = pi001 & pi114;
assign w5137 = w413 & w475;
assign w5138 = ~w449 & ~w5137;
assign w5139 = w5136 & ~w5138;
assign w5140 = ~w989 & ~w990;
assign w5141 = w536 & ~w5140;
assign w5142 = w466 & w524;
assign w5143 = ~pi001 & w446;
assign w5144 = w926 & w5143;
assign w5145 = ~w5142 & ~w5144;
assign w5146 = ~w5135 & ~w5139;
assign w5147 = ~w5141 & w5145;
assign w5148 = w5146 & w5147;
assign w5149 = ~w5132 & w5148;
assign w5150 = ~w5127 & w5149;
assign w5151 = (pi029 & ~w5098) | (pi029 & w18453) | (~w5098 & w18453);
assign w5152 = w5150 & ~w5151;
assign w5153 = ~w5072 & w5152;
assign w5154 = w5072 & ~w5152;
assign w5155 = ~w5153 & ~w5154;
assign w5156 = w1131 & ~w5155;
assign w5157 = ~w1131 & w5155;
assign w5158 = ~w5156 & ~w5157;
assign w5159 = w23 & w33;
assign w5160 = ~pi014 & w60;
assign w5161 = w20 & w5160;
assign w5162 = ~w106 & ~w1342;
assign w5163 = ~w65 & ~w5159;
assign w5164 = w5162 & w18454;
assign w5165 = pi083 & ~w5164;
assign w5166 = ~w77 & ~w188;
assign w5167 = ~pi083 & w5166;
assign w5168 = ~w7 & ~w236;
assign w5169 = w5167 & ~w5168;
assign w5170 = ~w30 & ~w108;
assign w5171 = ~pi040 & w5170;
assign w5172 = ~w5169 & w5171;
assign w5173 = ~pi014 & w51;
assign w5174 = w3 & ~w33;
assign w5175 = ~w194 & ~w5173;
assign w5176 = (~pi083 & ~w5175) | (~pi083 & w18455) | (~w5175 & w18455);
assign w5177 = pi014 & w20;
assign w5178 = w60 & w5177;
assign w5179 = w46 & w107;
assign w5180 = w8 & w58;
assign w5181 = ~w5179 & ~w5180;
assign w5182 = ~w82 & ~w5178;
assign w5183 = w5181 & w5182;
assign w5184 = pi040 & w5183;
assign w5185 = ~w5165 & w5172;
assign w5186 = ~w5176 & w5184;
assign w5187 = ~w5185 & ~w5186;
assign w5188 = w40 & w107;
assign w5189 = w78 & w83;
assign w5190 = ~w231 & ~w5188;
assign w5191 = pi040 & ~w5189;
assign w5192 = w5190 & w5191;
assign w5193 = ~pi083 & ~w179;
assign w5194 = ~w90 & w5193;
assign w5195 = w5192 & ~w5194;
assign w5196 = w0 & w33;
assign w5197 = (~pi040 & ~w5196) | (~pi040 & w123) | (~w5196 & w123);
assign w5198 = pi083 & w150;
assign w5199 = w11 & ~w1327;
assign w5200 = ~w236 & ~w5198;
assign w5201 = w5200 & w18456;
assign w5202 = pi083 & ~w160;
assign w5203 = ~pi082 & w40;
assign w5204 = ~w115 & ~w189;
assign w5205 = w5202 & w5204;
assign w5206 = ~w5203 & w5205;
assign w5207 = w2 & w40;
assign w5208 = ~pi083 & ~w151;
assign w5209 = ~w5173 & ~w5207;
assign w5210 = w5208 & w5209;
assign w5211 = ~w5206 & ~w5210;
assign w5212 = pi078 & ~w5211;
assign w5213 = ~w5195 & ~w5201;
assign w5214 = w5212 & ~w5213;
assign w5215 = ~w36 & ~w40;
assign w5216 = w33 & ~w5215;
assign w5217 = w23 & w64;
assign w5218 = w56 & w177;
assign w5219 = ~w5216 & ~w5217;
assign w5220 = ~pi040 & ~w5218;
assign w5221 = w5219 & w5220;
assign w5222 = ~w80 & w83;
assign w5223 = ~w41 & w5222;
assign w5224 = ~pi083 & w5223;
assign w5225 = pi040 & ~w165;
assign w5226 = ~w212 & w5225;
assign w5227 = w9 & w102;
assign w5228 = w5226 & ~w5227;
assign w5229 = ~w5224 & w5228;
assign w5230 = ~pi072 & w89;
assign w5231 = ~w5196 & ~w5230;
assign w5232 = pi083 & ~w5231;
assign w5233 = (pi014 & ~w33) | (pi014 & w17902) | (~w33 & w17902);
assign w5234 = ~w5231 & w18457;
assign w5235 = w16 & w18458;
assign w5236 = (~pi078 & ~w107) | (~pi078 & w18459) | (~w107 & w18459);
assign w5237 = ~w5235 & w5236;
assign w5238 = ~w5234 & w5237;
assign w5239 = (w5238 & w5229) | (w5238 & w18460) | (w5229 & w18460);
assign w5240 = ~w5214 & ~w5239;
assign w5241 = ~pi083 & w114;
assign w5242 = (pi014 & w5241) | (pi014 & w18461) | (w5241 & w18461);
assign w5243 = ~w5240 & w18462;
assign w5244 = ~w402 & w5243;
assign w5245 = w402 & ~w5243;
assign w5246 = ~w5244 & ~w5245;
assign w5247 = ~pi221 & w901;
assign w5248 = pi221 & ~w901;
assign w5249 = ~w5247 & ~w5248;
assign w5250 = w5246 & w5249;
assign w5251 = ~w5246 & ~w5249;
assign w5252 = ~w5250 & ~w5251;
assign w5253 = ~w5158 & w5252;
assign w5254 = ~pi529 & ~w5253;
assign w5255 = w5158 & ~w5252;
assign w5256 = w5254 & ~w5255;
assign w5257 = ~pi221 & pi432;
assign w5258 = pi529 & ~w5257;
assign w5259 = pi221 & ~pi432;
assign w5260 = w5258 & ~w5259;
assign w5261 = ~w5256 & ~w5260;
assign w5262 = (pi083 & ~w33) | (pi083 & w46) | (~w33 & w46);
assign w5263 = ~w5207 & w5262;
assign w5264 = w5166 & w18463;
assign w5265 = (~w13 & w5264) | (~w13 & w18464) | (w5264 & w18464);
assign w5266 = pi040 & ~w5265;
assign w5267 = w81 & w46;
assign w5268 = ~w150 & ~w5267;
assign w5269 = w25 & w202;
assign w5270 = ~w128 & ~w5269;
assign w5271 = w107 & w18465;
assign w5272 = ~pi040 & ~w5270;
assign w5273 = ~w5271 & ~w5272;
assign w5274 = w5268 & w5273;
assign w5275 = ~w5266 & w5274;
assign w5276 = ~pi078 & ~w5275;
assign w5277 = w2 & w8;
assign w5278 = ~pi083 & w81;
assign w5279 = ~pi107 & w33;
assign w5280 = w84 & w5279;
assign w5281 = ~w5278 & ~w5280;
assign w5282 = ~w27 & ~w165;
assign w5283 = ~w236 & w5282;
assign w5284 = w5281 & w5283;
assign w5285 = ~w5159 & ~w5189;
assign w5286 = ~w21 & ~w210;
assign w5287 = ~pi083 & ~w5286;
assign w5288 = w33 & w78;
assign w5289 = w41 & w64;
assign w5290 = ~w5288 & ~w5289;
assign w5291 = ~w5287 & w5290;
assign w5292 = pi040 & ~w5291;
assign w5293 = ~w49 & ~w173;
assign w5294 = (w46 & ~w5293) | (w46 & w18467) | (~w5293 & w18467);
assign w5295 = ~w108 & ~w1293;
assign w5296 = ~w5161 & w5295;
assign w5297 = ~w5294 & w5296;
assign w5298 = ~w5292 & w5297;
assign w5299 = (pi078 & ~w5298) | (pi078 & w18468) | (~w5298 & w18468);
assign w5300 = ~w128 & ~w5177;
assign w5301 = ~w1292 & w5300;
assign w5302 = pi083 & ~w5301;
assign w5303 = w50 & w71;
assign w5304 = w0 & w83;
assign w5305 = ~w5303 & ~w5304;
assign w5306 = ~w30 & w5305;
assign w5307 = ~pi083 & ~w5306;
assign w5308 = w84 & w107;
assign w5309 = w20 & ~w50;
assign w5310 = ~w70 & w5309;
assign w5311 = ~w5308 & ~w5310;
assign w5312 = ~w5302 & ~w5307;
assign w5313 = (~pi040 & ~w5312) | (~pi040 & w18469) | (~w5312 & w18469);
assign w5314 = w83 & w70;
assign w5315 = ~w16 & ~w5314;
assign w5316 = (pi040 & w16) | (pi040 & w1348) | (w16 & w1348);
assign w5317 = (w5316 & ~w1318) | (w5316 & w20780) | (~w1318 & w20780);
assign w5318 = w3 & w222;
assign w5319 = ~w81 & ~w5160;
assign w5320 = ~w5318 & w5319;
assign w5321 = w88 & ~w5320;
assign w5322 = ~w171 & ~w5303;
assign w5323 = w8 & ~w5322;
assign w5324 = ~w228 & ~w5323;
assign w5325 = ~w5321 & w5324;
assign w5326 = ~w5317 & w5325;
assign w5327 = ~w5313 & w5326;
assign w5328 = ~w5299 & w5327;
assign w5329 = ~w5276 & w5328;
assign w5330 = ~w364 & ~w1385;
assign w5331 = w252 & w376;
assign w5332 = ~w305 & ~w316;
assign w5333 = ~w1086 & ~w5331;
assign w5334 = w5332 & w5333;
assign w5335 = pi123 & w1036;
assign w5336 = w5334 & ~w5335;
assign w5337 = w252 & w304;
assign w5338 = ~w1265 & ~w5337;
assign w5339 = w1038 & w1275;
assign w5340 = ~w275 & ~w1081;
assign w5341 = (w383 & ~w5340) | (w383 & w18470) | (~w5340 & w18470);
assign w5342 = ~pi027 & w346;
assign w5343 = ~w260 & ~w284;
assign w5344 = ~w5342 & w5343;
assign w5345 = ~w5341 & w5344;
assign w5346 = (pi048 & ~w5338) | (pi048 & w18471) | (~w5338 & w18471);
assign w5347 = w5345 & ~w5346;
assign w5348 = (pi020 & ~w5347) | (pi020 & w18472) | (~w5347 & w18472);
assign w5349 = w286 & w294;
assign w5350 = ~w283 & ~w5331;
assign w5351 = ~pi123 & ~w5349;
assign w5352 = w5350 & w5351;
assign w5353 = ~w1109 & ~w5053;
assign w5354 = ~w276 & w5353;
assign w5355 = pi123 & w5354;
assign w5356 = ~w288 & w5352;
assign w5357 = ~w5355 & ~w5356;
assign w5358 = w257 & ~w270;
assign w5359 = ~w281 & w5358;
assign w5360 = (~pi048 & w5357) | (~pi048 & w18473) | (w5357 & w18473);
assign w5361 = ~w253 & ~w336;
assign w5362 = pi123 & ~w5361;
assign w5363 = ~w281 & ~w315;
assign w5364 = ~pi123 & ~w285;
assign w5365 = ~w5363 & w5364;
assign w5366 = ~w1068 & ~w5365;
assign w5367 = ~w5362 & w5366;
assign w5368 = pi048 & ~w5367;
assign w5369 = ~w1109 & ~w1264;
assign w5370 = ~pi048 & ~w5369;
assign w5371 = w364 & w383;
assign w5372 = w283 & w394;
assign w5373 = ~w5371 & ~w5372;
assign w5374 = ~w5370 & w5373;
assign w5375 = ~w312 & w5374;
assign w5376 = ~w5368 & w5375;
assign w5377 = ~pi020 & ~w5376;
assign w5378 = (pi048 & w278) | (pi048 & w1420) | (w278 & w1420);
assign w5379 = ~w278 & ~w1240;
assign w5380 = (w5378 & ~w1392) | (w5378 & w18474) | (~w1392 & w18474);
assign w5381 = pi093 & w258;
assign w5382 = ~w364 & ~w5381;
assign w5383 = w1416 & ~w5382;
assign w5384 = ~w283 & ~w1108;
assign w5385 = w343 & ~w5384;
assign w5386 = w261 & w1416;
assign w5387 = w1259 & w5386;
assign w5388 = ~w5054 & ~w5387;
assign w5389 = ~w5383 & ~w5385;
assign w5390 = w5388 & w5389;
assign w5391 = ~w5380 & w5390;
assign w5392 = ~w5360 & ~w5377;
assign w5393 = w5392 & w18475;
assign w5394 = ~w5329 & w5393;
assign w5395 = w5329 & ~w5393;
assign w5396 = ~w5394 & ~w5395;
assign w5397 = ~w1128 & w5152;
assign w5398 = w1128 & ~w5152;
assign w5399 = ~w5397 & ~w5398;
assign w5400 = w5396 & w5399;
assign w5401 = ~w5396 & ~w5399;
assign w5402 = ~w5400 & ~w5401;
assign w5403 = w807 & w18476;
assign w5404 = (pi121 & ~w807) | (pi121 & w18477) | (~w807 & w18477);
assign w5405 = ~w5403 & ~w5404;
assign w5406 = w251 & w5405;
assign w5407 = ~w251 & ~w5405;
assign w5408 = ~w5406 & ~w5407;
assign w5409 = (~pi529 & ~w5408) | (~pi529 & w18478) | (~w5408 & w18478);
assign w5410 = ~w5402 & ~w5408;
assign w5411 = w5409 & ~w5410;
assign w5412 = ~pi121 & pi441;
assign w5413 = pi529 & ~w5412;
assign w5414 = pi121 & ~pi441;
assign w5415 = w5413 & ~w5414;
assign w5416 = ~w5411 & ~w5415;
assign w5417 = ~w478 & ~w538;
assign w5418 = pi114 & w5417;
assign w5419 = ~w467 & ~w498;
assign w5420 = ~pi114 & w5419;
assign w5421 = ~w5418 & ~w5420;
assign w5422 = ~w419 & ~w429;
assign w5423 = w5422 & w18479;
assign w5424 = (~pi001 & w5421) | (~pi001 & w18480) | (w5421 & w18480);
assign w5425 = w958 & w5084;
assign w5426 = ~w945 & ~w5425;
assign w5427 = (pi001 & ~w5426) | (pi001 & w18481) | (~w5426 & w18481);
assign w5428 = (w536 & ~w943) | (w536 & w18482) | (~w943 & w18482);
assign w5429 = ~w487 & ~w1147;
assign w5430 = (~pi013 & ~w5429) | (~pi013 & w18483) | (~w5429 & w18483);
assign w5431 = ~w5427 & ~w5430;
assign w5432 = ~w5424 & w5431;
assign w5433 = w417 & w432;
assign w5434 = ~w993 & ~w5433;
assign w5435 = ~w525 & w5434;
assign w5436 = ~pi114 & ~w5435;
assign w5437 = pi013 & w405;
assign w5438 = ~w1004 & ~w5437;
assign w5439 = ~w521 & w5438;
assign w5440 = pi114 & ~w5439;
assign w5441 = w479 & w509;
assign w5442 = w405 & ~w411;
assign w5443 = ~w445 & w5442;
assign w5444 = ~w5441 & ~w5443;
assign w5445 = ~w5436 & ~w5440;
assign w5446 = (~pi001 & ~w5445) | (~pi001 & w18484) | (~w5445 & w18484);
assign w5447 = ~w447 & ~w950;
assign w5448 = pi114 & ~w5447;
assign w5449 = ~pi114 & ~w415;
assign w5450 = ~w520 & w5449;
assign w5451 = ~w922 & ~w5450;
assign w5452 = ~w5448 & w5451;
assign w5453 = pi001 & ~w5452;
assign w5454 = w414 & w18485;
assign w5455 = ~w426 & ~w5454;
assign w5456 = w415 & w5110;
assign w5457 = ~w1004 & ~w5456;
assign w5458 = w539 & w18486;
assign w5459 = ~pi001 & ~w5457;
assign w5460 = ~w5458 & ~w5459;
assign w5461 = w5455 & w5460;
assign w5462 = ~w5453 & w5461;
assign w5463 = ~pi029 & ~w5462;
assign w5464 = ~w989 & ~w5102;
assign w5465 = ~pi013 & w417;
assign w5466 = w417 & w411;
assign w5467 = ~w5074 & ~w5466;
assign w5468 = (pi001 & w5074) | (pi001 & w7311) | (w5074 & w7311);
assign w5469 = (w5468 & ~w5464) | (w5468 & w18487) | (~w5464 & w18487);
assign w5470 = ~w456 & ~w509;
assign w5471 = w1187 & ~w5470;
assign w5472 = ~w467 & ~w969;
assign w5473 = w5136 & ~w5472;
assign w5474 = pi001 & w536;
assign w5475 = w516 & w5474;
assign w5476 = ~w5129 & ~w5475;
assign w5477 = ~w5471 & ~w5473;
assign w5478 = w5476 & w5477;
assign w5479 = ~w5469 & w5478;
assign w5480 = ~w5463 & w18488;
assign w5481 = (pi029 & ~w5432) | (pi029 & w20781) | (~w5432 & w20781);
assign w5482 = w5480 & ~w5481;
assign w5483 = ~w1021 & w5482;
assign w5484 = w1021 & ~w5482;
assign w5485 = ~w5483 & ~w5484;
assign w5486 = w5155 & w5485;
assign w5487 = ~w5155 & ~w5485;
assign w5488 = ~w5486 & ~w5487;
assign w5489 = ~w567 & ~w712;
assign w5490 = ~w586 & ~w719;
assign w5491 = ~w711 & w5490;
assign w5492 = ~w788 & ~w795;
assign w5493 = ~w883 & w5492;
assign w5494 = w5491 & w5493;
assign w5495 = (~pi102 & ~w5494) | (~pi102 & w18489) | (~w5494 & w18489);
assign w5496 = ~w589 & ~w766;
assign w5497 = ~w742 & w5496;
assign w5498 = (pi104 & ~w598) | (pi104 & w570) | (~w598 & w570);
assign w5499 = pi102 & ~w5498;
assign w5500 = (w5499 & ~w5497) | (w5499 & w18490) | (~w5497 & w18490);
assign w5501 = pi033 & w565;
assign w5502 = ~w605 & ~w5501;
assign w5503 = (w604 & ~w5502) | (w604 & w18491) | (~w5502 & w18491);
assign w5504 = w607 & w1456;
assign w5505 = ~w840 & ~w1450;
assign w5506 = (pi012 & ~w1456) | (pi012 & w18492) | (~w1456 & w18492);
assign w5507 = w5505 & w5506;
assign w5508 = ~w5503 & w5507;
assign w5509 = ~w5500 & w5508;
assign w5510 = ~w5495 & w5509;
assign w5511 = ~w633 & ~w746;
assign w5512 = (~pi104 & ~w569) | (~pi104 & w622) | (~w569 & w622);
assign w5513 = w5511 & w5512;
assign w5514 = (pi104 & ~w598) | (pi104 & w604) | (~w598 & w604);
assign w5515 = ~w876 & w5514;
assign w5516 = (~w574 & w5513) | (~w574 & w18493) | (w5513 & w18493);
assign w5517 = pi102 & ~w5516;
assign w5518 = w783 & w18494;
assign w5519 = w584 & w689;
assign w5520 = ~w676 & ~w5519;
assign w5521 = ~pi012 & ~w722;
assign w5522 = w567 & w604;
assign w5523 = w5521 & ~w5522;
assign w5524 = ~pi102 & ~w5520;
assign w5525 = w5523 & ~w5524;
assign w5526 = ~w5518 & w5525;
assign w5527 = ~w5517 & w5526;
assign w5528 = ~w5510 & ~w5527;
assign w5529 = ~w661 & ~w719;
assign w5530 = ~pi104 & ~w794;
assign w5531 = w5529 & w5530;
assign w5532 = w678 & ~w837;
assign w5533 = ~w670 & w5532;
assign w5534 = ~w581 & w5531;
assign w5535 = ~w5533 & ~w5534;
assign w5536 = w572 & w607;
assign w5537 = ~w680 & ~w5536;
assign w5538 = (~pi102 & w5535) | (~pi102 & w18495) | (w5535 & w18495);
assign w5539 = (~pi104 & ~w1456) | (~pi104 & w703) | (~w1456 & w703);
assign w5540 = ~pi127 & w561;
assign w5541 = pi126 & w585;
assign w5542 = ~w567 & ~w5541;
assign w5543 = pi104 & w5542;
assign w5544 = w560 & w5540;
assign w5545 = w5543 & ~w5544;
assign w5546 = w1479 & w5539;
assign w5547 = ~w5545 & ~w5546;
assign w5548 = (pi102 & w5547) | (pi102 & w18496) | (w5547 & w18496);
assign w5549 = ~w661 & ~w674;
assign w5550 = w755 & ~w5549;
assign w5551 = ~w5538 & ~w5548;
assign w5552 = ~w785 & ~w5550;
assign w5553 = w5551 & w5552;
assign w5554 = ~w5528 & w5553;
assign w5555 = ~pi143 & w5554;
assign w5556 = pi143 & ~w5554;
assign w5557 = ~w5555 & ~w5556;
assign w5558 = ~w248 & w702;
assign w5559 = w248 & ~w702;
assign w5560 = ~w5558 & ~w5559;
assign w5561 = w5557 & w5560;
assign w5562 = ~w5557 & ~w5560;
assign w5563 = ~w5561 & ~w5562;
assign w5564 = w5488 & w5563;
assign w5565 = ~pi529 & ~w5564;
assign w5566 = ~w5488 & ~w5563;
assign w5567 = w5565 & ~w5566;
assign w5568 = ~pi143 & pi412;
assign w5569 = pi529 & ~w5568;
assign w5570 = pi143 & ~pi412;
assign w5571 = w5569 & ~w5570;
assign w5572 = ~w5567 & ~w5571;
assign w5573 = w700 & w18497;
assign w5574 = (pi150 & ~w700) | (pi150 & w18498) | (~w700 & w18498);
assign w5575 = ~w5573 & ~w5574;
assign w5576 = ~w1021 & w1206;
assign w5577 = w1021 & ~w1206;
assign w5578 = ~w5576 & ~w5577;
assign w5579 = w15 & w33;
assign w5580 = ~w69 & ~w81;
assign w5581 = (pi083 & ~w5580) | (pi083 & w18499) | (~w5580 & w18499);
assign w5582 = ~pi072 & w40;
assign w5583 = w12 & w60;
assign w5584 = ~w27 & ~w5582;
assign w5585 = ~w5583 & w5584;
assign w5586 = w104 & w18500;
assign w5587 = w5585 & ~w5586;
assign w5588 = (~pi040 & ~w5587) | (~pi040 & w18501) | (~w5587 & w18501);
assign w5589 = ~w42 & ~w1341;
assign w5590 = ~w172 & ~w227;
assign w5591 = w5589 & w5590;
assign w5592 = (~pi083 & w135) | (~pi083 & w18502) | (w135 & w18502);
assign w5593 = (pi040 & w5592) | (pi040 & w18503) | (w5592 & w18503);
assign w5594 = ~w48 & ~w189;
assign w5595 = w204 & ~w5594;
assign w5596 = ~w7 & ~w50;
assign w5597 = w202 & ~w5596;
assign w5598 = ~w5178 & ~w5597;
assign w5599 = ~w5595 & w5598;
assign w5600 = (~w5593 & w5591) | (~w5593 & w18504) | (w5591 & w18504);
assign w5601 = ~w5588 & w5600;
assign w5602 = ~pi014 & ~w116;
assign w5603 = w5197 & ~w5602;
assign w5604 = w15 & w38;
assign w5605 = pi040 & ~w5604;
assign w5606 = pi083 & w106;
assign w5607 = w5605 & ~w5606;
assign w5608 = ~w1 & ~w35;
assign w5609 = w5607 & ~w5608;
assign w5610 = w20 & w26;
assign w5611 = ~w172 & w18505;
assign w5612 = ~pi083 & ~w5611;
assign w5613 = pi014 & w5288;
assign w5614 = w5288 & w17902;
assign w5615 = pi072 & w83;
assign w5616 = pi108 & w23;
assign w5617 = ~w5615 & ~w5616;
assign w5618 = w123 & ~w5617;
assign w5619 = ~w5618 & w18506;
assign w5620 = ~w5612 & w5619;
assign w5621 = ~w5603 & ~w5609;
assign w5622 = w5620 & ~w5621;
assign w5623 = ~w15 & ~w70;
assign w5624 = ~w41 & w5623;
assign w5625 = w2 & ~w5624;
assign w5626 = (~pi083 & ~w107) | (~pi083 & w18507) | (~w107 & w18507);
assign w5627 = ~w5625 & w5626;
assign w5628 = pi083 & ~w133;
assign w5629 = ~w1341 & ~w5161;
assign w5630 = w5628 & w5629;
assign w5631 = w187 & w210;
assign w5632 = (pi083 & w5631) | (pi083 & w18508) | (w5631 & w18508);
assign w5633 = ~pi083 & w128;
assign w5634 = ~w5173 & ~w5188;
assign w5635 = ~w5633 & w5634;
assign w5636 = w0 & w38;
assign w5637 = w78 & w1330;
assign w5638 = pi082 & w5636;
assign w5639 = ~w5637 & ~w5638;
assign w5640 = (pi040 & ~w5635) | (pi040 & w18509) | (~w5635 & w18509);
assign w5641 = w5639 & ~w5640;
assign w5642 = ~w5627 & ~w5630;
assign w5643 = ~pi040 & w5642;
assign w5644 = w5641 & ~w5643;
assign w5645 = ~pi078 & ~w5622;
assign w5646 = w5644 & ~w5645;
assign w5647 = (pi078 & ~w5601) | (pi078 & w18510) | (~w5601 & w18510);
assign w5648 = w5646 & ~w5647;
assign w5649 = ~w1282 & w5648;
assign w5650 = w1282 & ~w5648;
assign w5651 = ~w5649 & ~w5650;
assign w5652 = w5578 & ~w5651;
assign w5653 = ~w5578 & w5651;
assign w5654 = ~w5652 & ~w5653;
assign w5655 = ~w5575 & w5654;
assign w5656 = w5575 & ~w5654;
assign w5657 = ~w5655 & ~w5656;
assign w5658 = ~pi150 & pi483;
assign w5659 = pi150 & ~pi483;
assign w5660 = ~w5658 & ~w5659;
assign w5661 = ~w145 & w5329;
assign w5662 = w145 & ~w5329;
assign w5663 = ~w5661 & ~w5662;
assign w5664 = w5155 & w5663;
assign w5665 = ~w5155 & ~w5663;
assign w5666 = ~w5664 & ~w5665;
assign w5667 = ~pi137 & w5554;
assign w5668 = pi137 & ~w5554;
assign w5669 = ~w5667 & ~w5668;
assign w5670 = w811 & w5669;
assign w5671 = ~w811 & ~w5669;
assign w5672 = ~w5670 & ~w5671;
assign w5673 = (~pi529 & ~w5666) | (~pi529 & w18511) | (~w5666 & w18511);
assign w5674 = ~w5666 & ~w5672;
assign w5675 = w5673 & ~w5674;
assign w5676 = ~pi137 & pi495;
assign w5677 = pi529 & ~w5676;
assign w5678 = pi137 & ~pi495;
assign w5679 = w5677 & ~w5678;
assign w5680 = ~w5675 & ~w5679;
assign w5681 = ~w2334 & ~w2397;
assign w5682 = ~pi080 & ~w5681;
assign w5683 = ~pi079 & pi080;
assign w5684 = w2292 & w5683;
assign w5685 = ~w2413 & ~w5684;
assign w5686 = ~w5682 & w5685;
assign w5687 = w2299 & w2376;
assign w5688 = pi075 & w5687;
assign w5689 = w2333 & w2337;
assign w5690 = ~w2320 & ~w5689;
assign w5691 = ~w5688 & w5690;
assign w5692 = (~pi080 & ~w5691) | (~pi080 & w18512) | (~w5691 & w18512);
assign w5693 = ~pi080 & pi110;
assign w5694 = (~pi075 & w2393) | (~pi075 & w18513) | (w2393 & w18513);
assign w5695 = pi075 & w2363;
assign w5696 = ~pi071 & w2329;
assign w5697 = w2421 & w5695;
assign w5698 = w2329 & w2307;
assign w5699 = ~w5697 & ~w5698;
assign w5700 = (~pi073 & ~w5699) | (~pi073 & w18514) | (~w5699 & w18514);
assign w5701 = w2347 & w2359;
assign w5702 = ~w2375 & ~w5701;
assign w5703 = (w2421 & ~w5702) | (w2421 & w18515) | (~w5702 & w18515);
assign w5704 = ~w5692 & ~w5700;
assign w5705 = ~w5703 & w5704;
assign w5706 = pi075 & w2316;
assign w5707 = pi075 & w2299;
assign w5708 = ~w2410 & ~w5706;
assign w5709 = ~pi079 & w2299;
assign w5710 = w2337 & w2363;
assign w5711 = pi080 & w5710;
assign w5712 = ~w2368 & w5709;
assign w5713 = ~w5711 & ~w5712;
assign w5714 = ~pi110 & w2359;
assign w5715 = ~pi075 & pi079;
assign w5716 = ~pi042 & w5715;
assign w5717 = w2359 & w18518;
assign w5718 = w5715 & w2346;
assign w5719 = ~w5717 & ~w5718;
assign w5720 = w5713 & w5719;
assign w5721 = (~pi073 & ~w5720) | (~pi073 & w18519) | (~w5720 & w18519);
assign w5722 = w2291 & w2359;
assign w5723 = w2293 & w2337;
assign w5724 = ~w2384 & ~w5723;
assign w5725 = (pi080 & ~w5724) | (pi080 & w18520) | (~w5724 & w18520);
assign w5726 = pi079 & w2290;
assign w5727 = w2333 & w2381;
assign w5728 = w2345 & w5707;
assign w5729 = ~w5727 & ~w5728;
assign w5730 = w2368 & w5726;
assign w5731 = w5729 & ~w5730;
assign w5732 = w2347 & w5726;
assign w5733 = ~pi071 & w2314;
assign w5734 = w2345 & w5733;
assign w5735 = ~w5732 & ~w5734;
assign w5736 = ~pi079 & w2329;
assign w5737 = ~w2326 & ~w5736;
assign w5738 = pi042 & ~pi075;
assign w5739 = ~w5706 & ~w5738;
assign w5740 = w5737 & w5739;
assign w5741 = w2409 & ~w5740;
assign w5742 = pi073 & ~w5735;
assign w5743 = ~w5741 & ~w5742;
assign w5744 = ~w5725 & w5731;
assign w5745 = w5743 & w5744;
assign w5746 = w2363 & w5715;
assign w5747 = (~pi080 & ~w5690) | (~pi080 & w18521) | (~w5690 & w18521);
assign w5748 = w2298 & w2347;
assign w5749 = (~pi073 & w5747) | (~pi073 & w18522) | (w5747 & w18522);
assign w5750 = ~pi079 & w2410;
assign w5751 = ~w5732 & ~w5750;
assign w5752 = (w2415 & ~w5751) | (w2415 & w18523) | (~w5751 & w18523);
assign w5753 = pi071 & w2293;
assign w5754 = w2337 & w5753;
assign w5755 = w2381 & w5733;
assign w5756 = ~w5754 & ~w5755;
assign w5757 = w2306 & w5736;
assign w5758 = ~w2358 & ~w5687;
assign w5759 = ~w5757 & w5758;
assign w5760 = w5756 & w5759;
assign w5761 = w2337 & w5714;
assign w5762 = w2302 & w5696;
assign w5763 = ~w5761 & ~w5762;
assign w5764 = ~w2343 & ~w2370;
assign w5765 = pi075 & w2346;
assign w5766 = pi071 & w2329;
assign w5767 = ~w5765 & ~w5766;
assign w5768 = w5764 & w5767;
assign w5769 = pi079 & w2403;
assign w5770 = ~w5768 & w5769;
assign w5771 = ~pi080 & ~w5763;
assign w5772 = ~w5770 & ~w5771;
assign w5773 = w2409 & ~w5760;
assign w5774 = w5772 & ~w5773;
assign w5775 = w5774 & w18524;
assign w5776 = (pi015 & ~w5745) | (pi015 & w20782) | (~w5745 & w20782);
assign w5777 = w5775 & ~w5776;
assign w5778 = (~pi015 & ~w5705) | (~pi015 & w18525) | (~w5705 & w18525);
assign w5779 = w5777 & ~w5778;
assign w5780 = w5777 & w18526;
assign w5781 = (pi190 & ~w5777) | (pi190 & w18527) | (~w5777 & w18527);
assign w5782 = ~w5780 & ~w5781;
assign w5783 = ~w1692 & w1936;
assign w5784 = w1692 & ~w1936;
assign w5785 = ~w5783 & ~w5784;
assign w5786 = w2071 & w2138;
assign w5787 = ~w2099 & ~w2143;
assign w5788 = (pi092 & ~w5787) | (pi092 & w18528) | (~w5787 & w18528);
assign w5789 = pi050 & w2151;
assign w5790 = ~pi085 & w2062;
assign w5791 = w2107 & w2157;
assign w5792 = w2051 & w2138;
assign w5793 = ~w5790 & ~w5791;
assign w5794 = ~w5792 & w5793;
assign w5795 = w2151 & w18529;
assign w5796 = w5794 & ~w5795;
assign w5797 = (~pi089 & ~w5796) | (~pi089 & w18530) | (~w5796 & w18530);
assign w5798 = ~w2097 & ~w2153;
assign w5799 = w2073 & w2107;
assign w5800 = ~w2094 & ~w5799;
assign w5801 = w5798 & w5800;
assign w5802 = pi087 & ~pi092;
assign w5803 = pi085 & w2121;
assign w5804 = (pi046 & w5803) | (pi046 & w18531) | (w5803 & w18531);
assign w5805 = ~pi050 & ~pi092;
assign w5806 = w2073 & w5805;
assign w5807 = (pi089 & w5804) | (pi089 & w18532) | (w5804 & w18532);
assign w5808 = ~w2108 & ~w2167;
assign w5809 = pi028 & ~w5808;
assign w5810 = w2052 & w2111;
assign w5811 = ~w2139 & ~w5810;
assign w5812 = ~w5809 & w5811;
assign w5813 = ~pi092 & ~w5812;
assign w5814 = w2062 & w2075;
assign w5815 = ~pi085 & w5814;
assign w5816 = ~w2130 & ~w5815;
assign w5817 = ~w5813 & w18533;
assign w5818 = ~w5797 & w5817;
assign w5819 = (pi053 & ~w5818) | (pi053 & w18534) | (~w5818 & w18534);
assign w5820 = w2049 & w18979;
assign w5821 = ~w2085 & ~w2095;
assign w5822 = ~w2122 & ~w5821;
assign w5823 = ~pi028 & ~pi092;
assign w5824 = ~pi087 & w5823;
assign w5825 = w5823 & w18535;
assign w5826 = ~w5822 & ~w5825;
assign w5827 = w2052 & w2132;
assign w5828 = w2051 & w2073;
assign w5829 = ~w2094 & w18536;
assign w5830 = ~w2078 & ~w2093;
assign w5831 = pi092 & w5830;
assign w5832 = w2085 & w2095;
assign w5833 = ~pi092 & ~w5832;
assign w5834 = w2052 & w2163;
assign w5835 = ~w2125 & ~w5834;
assign w5836 = ~pi028 & ~pi089;
assign w5837 = ~w5835 & w5836;
assign w5838 = ~w2137 & w2185;
assign w5839 = ~w5837 & ~w5838;
assign w5840 = (~pi089 & w5832) | (~pi089 & w2177) | (w5832 & w2177);
assign w5841 = ~w5831 & w5840;
assign w5842 = w5839 & ~w5841;
assign w5843 = ~pi092 & ~w5829;
assign w5844 = w2077 & w2124;
assign w5845 = w2098 & w2119;
assign w5846 = (pi092 & w5845) | (pi092 & w18538) | (w5845 & w18538);
assign w5847 = ~pi028 & w2049;
assign w5848 = ~pi046 & pi087;
assign w5849 = w2100 & w5848;
assign w5850 = ~w2163 & w5847;
assign w5851 = ~w5849 & ~w5850;
assign w5852 = ~pi092 & ~w5851;
assign w5853 = w2131 & w2187;
assign w5854 = ~pi092 & w2049;
assign w5855 = pi087 & w2056;
assign w5856 = w5854 & w5855;
assign w5857 = ~w5853 & ~w5856;
assign w5858 = ~w5852 & w18539;
assign w5859 = pi085 & w2049;
assign w5860 = w2098 & w5859;
assign w5861 = (pi092 & w5860) | (pi092 & w18540) | (w5860 & w18540);
assign w5862 = w2080 & w5823;
assign w5863 = w2073 & w2100;
assign w5864 = ~pi085 & w2138;
assign w5865 = w2157 & w5864;
assign w5866 = ~w5862 & ~w5863;
assign w5867 = ~w5865 & w5866;
assign w5868 = pi085 & ~pi092;
assign w5869 = w2059 & w18541;
assign w5870 = w2110 & w5868;
assign w5871 = ~w5869 & ~w5870;
assign w5872 = (pi089 & ~w5867) | (pi089 & w18542) | (~w5867 & w18542);
assign w5873 = w5871 & ~w5872;
assign w5874 = ~pi089 & ~w5858;
assign w5875 = w5873 & ~w5874;
assign w5876 = (~w5842 & w20783) | (~w5842 & w20784) | (w20783 & w20784);
assign w5877 = w5875 & ~w5876;
assign w5878 = ~w5819 & w5877;
assign w5879 = ~w2041 & w5878;
assign w5880 = w2041 & ~w5878;
assign w5881 = ~w5879 & ~w5880;
assign w5882 = w5785 & ~w5881;
assign w5883 = ~w5785 & w5881;
assign w5884 = ~w5882 & ~w5883;
assign w5885 = ~w5782 & w5884;
assign w5886 = w5782 & ~w5884;
assign w5887 = ~w5885 & ~w5886;
assign w5888 = ~pi190 & pi410;
assign w5889 = pi190 & ~pi410;
assign w5890 = ~w5888 & ~w5889;
assign w5891 = ~w5393 & w5482;
assign w5892 = w5393 & ~w5482;
assign w5893 = ~w5891 & ~w5892;
assign w5894 = w1131 & ~w5893;
assign w5895 = ~w1131 & w5893;
assign w5896 = ~w5894 & ~w5895;
assign w5897 = ~w248 & w5072;
assign w5898 = w248 & ~w5072;
assign w5899 = ~w5897 & ~w5898;
assign w5900 = w807 & w18544;
assign w5901 = (pi136 & ~w807) | (pi136 & w18545) | (~w807 & w18545);
assign w5902 = ~w5900 & ~w5901;
assign w5903 = w5899 & w5902;
assign w5904 = ~w5899 & ~w5902;
assign w5905 = ~w5903 & ~w5904;
assign w5906 = ~w5896 & w5905;
assign w5907 = ~pi529 & ~w5906;
assign w5908 = w5896 & ~w5905;
assign w5909 = w5907 & ~w5908;
assign w5910 = ~pi136 & pi438;
assign w5911 = pi529 & ~w5910;
assign w5912 = pi136 & ~pi438;
assign w5913 = w5911 & ~w5912;
assign w5914 = ~w5909 & ~w5913;
assign w5915 = w2451 & ~w2511;
assign w5916 = ~w2538 & ~w5915;
assign w5917 = pi016 & w2532;
assign w5918 = w2448 & w2796;
assign w5919 = ~w2468 & ~w2771;
assign w5920 = ~w5918 & w5919;
assign w5921 = ~w2563 & w5917;
assign w5922 = w5920 & ~w5921;
assign w5923 = w2519 & w2748;
assign w5924 = ~w2512 & ~w5923;
assign w5925 = w2460 & w2478;
assign w5926 = w2480 & w2485;
assign w5927 = ~pi045 & ~w2545;
assign w5928 = w2821 & w5927;
assign w5929 = ~w5926 & ~w5928;
assign w5930 = ~w2816 & ~w5925;
assign w5931 = ~w2836 & w5930;
assign w5932 = w5929 & w5931;
assign w5933 = (~pi003 & ~w5932) | (~pi003 & w18546) | (~w5932 & w18546);
assign w5934 = ~w2461 & ~w2797;
assign w5935 = ~w2764 & w5934;
assign w5936 = ~pi120 & ~w5935;
assign w5937 = w2464 & w2775;
assign w5938 = pi016 & pi120;
assign w5939 = ~w2831 & ~w2835;
assign w5940 = (w5938 & ~w5939) | (w5938 & w18547) | (~w5939 & w18547);
assign w5941 = ~w5936 & w18548;
assign w5942 = ~w5933 & w5941;
assign w5943 = ~pi016 & w2568;
assign w5944 = ~pi045 & w2583;
assign w5945 = ~pi041 & pi074;
assign w5946 = ~pi081 & w5945;
assign w5947 = ~w2541 & ~w5946;
assign w5948 = pi045 & ~w5947;
assign w5949 = ~pi074 & w2570;
assign w5950 = w2451 & w2530;
assign w5951 = ~pi120 & w5950;
assign w5952 = ~w5949 & ~w5951;
assign w5953 = ~w5948 & w5952;
assign w5954 = w2532 & w2545;
assign w5955 = pi074 & ~pi120;
assign w5956 = w5954 & w5955;
assign w5957 = ~w2518 & ~w5938;
assign w5958 = w2478 & ~w5957;
assign w5959 = ~w2480 & w2828;
assign w5960 = pi045 & w5959;
assign w5961 = ~w5958 & ~w5960;
assign w5962 = ~w2461 & ~w5956;
assign w5963 = w5961 & w5962;
assign w5964 = ~pi003 & ~w5963;
assign w5965 = pi081 & w2588;
assign w5966 = w2557 & w2821;
assign w5967 = ~w2813 & ~w5966;
assign w5968 = w2499 & w5943;
assign w5969 = w5967 & ~w5968;
assign w5970 = (~pi120 & w5965) | (~pi120 & w18551) | (w5965 & w18551);
assign w5971 = w5969 & ~w5970;
assign w5972 = ~w5964 & w5971;
assign w5973 = (~pi044 & ~w5972) | (~pi044 & w18552) | (~w5972 & w18552);
assign w5974 = ~pi016 & w2447;
assign w5975 = ~w2481 & ~w5950;
assign w5976 = (w2467 & ~w5975) | (w2467 & w18553) | (~w5975 & w18553);
assign w5977 = pi120 & w5954;
assign w5978 = w2835 & w5955;
assign w5979 = w2835 & w18554;
assign w5980 = ~w5977 & ~w5979;
assign w5981 = ~w5976 & w5980;
assign w5982 = pi003 & ~w5981;
assign w5983 = pi081 & w2589;
assign w5984 = ~pi003 & w2563;
assign w5985 = w2531 & w5984;
assign w5986 = pi016 & w2512;
assign w5987 = w2499 & w2559;
assign w5988 = ~w5985 & ~w5986;
assign w5989 = w2589 & w18555;
assign w5990 = w5988 & w18556;
assign w5991 = w2569 & w2828;
assign w5992 = w2545 & w2748;
assign w5993 = ~pi045 & w5992;
assign w5994 = ~w5991 & ~w5993;
assign w5995 = w2805 & ~w5994;
assign w5996 = pi003 & pi120;
assign w5997 = w2464 & w2457;
assign w5998 = ~w5918 & ~w5997;
assign w5999 = w5996 & ~w5998;
assign w6000 = ~w5995 & ~w5999;
assign w6001 = w5990 & w6000;
assign w6002 = ~w5982 & w6001;
assign w6003 = ~w5973 & w6002;
assign w6004 = (pi044 & ~w5942) | (pi044 & w18557) | (~w5942 & w18557);
assign w6005 = w6003 & ~w6004;
assign w6006 = ~pi097 & ~pi116;
assign w6007 = w3076 & w6006;
assign w6008 = w2958 & w6007;
assign w6009 = ~pi000 & w2992;
assign w6010 = pi000 & w2980;
assign w6011 = ~w3084 & ~w6010;
assign w6012 = (pi116 & ~w2992) | (pi116 & w3094) | (~w2992 & w3094);
assign w6013 = (~w6012 & ~w6011) | (~w6012 & w18558) | (~w6011 & w18558);
assign w6014 = (pi058 & w6013) | (pi058 & w18559) | (w6013 & w18559);
assign w6015 = ~pi011 & ~pi116;
assign w6016 = ~pi000 & w2982;
assign w6017 = w2982 & w18560;
assign w6018 = w6009 & w6015;
assign w6019 = ~w6017 & ~w6018;
assign w6020 = w2962 & w3003;
assign w6021 = w2969 & w2958;
assign w6022 = ~pi116 & w3081;
assign w6023 = w3006 & w3066;
assign w6024 = w2962 & w2965;
assign w6025 = ~w3068 & ~w6024;
assign w6026 = ~w6022 & w6025;
assign w6027 = ~w6023 & w6026;
assign w6028 = ~w6020 & ~w6021;
assign w6029 = w6019 & w6028;
assign w6030 = w6027 & w6029;
assign w6031 = ~w2951 & ~w2976;
assign w6032 = (w3090 & ~w6031) | (w3090 & w18561) | (~w6031 & w18561);
assign w6033 = ~pi022 & w2982;
assign w6034 = w3006 & w6033;
assign w6035 = w3031 & w6009;
assign w6036 = ~w2967 & ~w6034;
assign w6037 = ~w6035 & w6036;
assign w6038 = ~w6032 & w6037;
assign w6039 = ~pi058 & ~w6030;
assign w6040 = ~w6039 & w18562;
assign w6041 = pi060 & ~w6040;
assign w6042 = ~w3017 & ~w3054;
assign w6043 = (~pi116 & ~w3023) | (~pi116 & w18231) | (~w3023 & w18231);
assign w6044 = w6042 & w6043;
assign w6045 = w2958 & w2962;
assign w6046 = ~pi011 & w2992;
assign w6047 = ~w6045 & ~w6046;
assign w6048 = pi116 & w6047;
assign w6049 = ~w6044 & ~w6048;
assign w6050 = (pi058 & w6049) | (pi058 & w18563) | (w6049 & w18563);
assign w6051 = w2978 & w2982;
assign w6052 = w2970 & w3094;
assign w6053 = ~w6051 & ~w6052;
assign w6054 = w3027 & w3066;
assign w6055 = ~w2996 & ~w6054;
assign w6056 = ~pi000 & w3066;
assign w6057 = w3060 & w6056;
assign w6058 = w6056 & w18564;
assign w6059 = ~pi058 & ~w6055;
assign w6060 = ~w6058 & ~w6059;
assign w6061 = w6053 & w6060;
assign w6062 = ~w6050 & w6061;
assign w6063 = ~pi060 & ~w6062;
assign w6064 = pi097 & w2984;
assign w6065 = ~w6056 & ~w6064;
assign w6066 = ~pi057 & ~w6065;
assign w6067 = w2963 & w2978;
assign w6068 = ~pi022 & w3060;
assign w6069 = ~w2996 & ~w6068;
assign w6070 = ~w2960 & w6069;
assign w6071 = pi116 & ~w6070;
assign w6072 = w3060 & w2961;
assign w6073 = w2952 & w18566;
assign w6074 = ~pi116 & w3068;
assign w6075 = ~w6072 & ~w6073;
assign w6076 = ~w6074 & w6075;
assign w6077 = ~w6071 & w6076;
assign w6078 = (~pi058 & ~w6077) | (~pi058 & w18567) | (~w6077 & w18567);
assign w6079 = w2982 & w2995;
assign w6080 = ~w3040 & ~w6079;
assign w6081 = (pi058 & w3040) | (pi058 & w3065) | (w3040 & w3065);
assign w6082 = (w6081 & ~w3014) | (w6081 & w20785) | (~w3014 & w20785);
assign w6083 = ~pi000 & w3054;
assign w6084 = ~pi000 & pi097;
assign w6085 = ~pi011 & w6084;
assign w6086 = ~w3081 & ~w6085;
assign w6087 = ~w6083 & w6086;
assign w6088 = w3075 & ~w6087;
assign w6089 = pi116 & w3006;
assign w6090 = ~w2952 & ~w3058;
assign w6091 = w6089 & ~w6090;
assign w6092 = w3041 & w3095;
assign w6093 = ~w6091 & ~w6092;
assign w6094 = ~w6088 & w6093;
assign w6095 = ~w6082 & w6094;
assign w6096 = ~w6078 & w6095;
assign w6097 = ~w6063 & w6096;
assign w6098 = ~w6041 & w6097;
assign w6099 = ~w6005 & w6098;
assign w6100 = w6005 & ~w6098;
assign w6101 = ~w6099 & ~w6100;
assign w6102 = ~w2683 & ~w2896;
assign w6103 = (pi118 & ~w6102) | (pi118 & w18568) | (~w6102 & w18568);
assign w6104 = ~w2865 & ~w3118;
assign w6105 = ~w3130 & w6104;
assign w6106 = ~w2714 & ~w2877;
assign w6107 = w6105 & w6106;
assign w6108 = ~w2673 & ~w2930;
assign w6109 = ~w2606 & ~w3154;
assign w6110 = ~pi118 & ~w6109;
assign w6111 = ~w2722 & ~w3186;
assign w6112 = ~w3169 & w6111;
assign w6113 = ~w6110 & w6112;
assign w6114 = (~pi034 & ~w6113) | (~pi034 & w18570) | (~w6113 & w18570);
assign w6115 = (~pi118 & ~w2891) | (~pi118 & w18571) | (~w2891 & w18571);
assign w6116 = ~w2599 & ~w2669;
assign w6117 = ~pi101 & ~w6116;
assign w6118 = (w3191 & w6117) | (w3191 & w18572) | (w6117 & w18572);
assign w6119 = ~w2919 & ~w6118;
assign w6120 = ~w6115 & w6119;
assign w6121 = ~w6114 & w6120;
assign w6122 = (pi034 & ~w6107) | (pi034 & w18573) | (~w6107 & w18573);
assign w6123 = ~pi103 & w2719;
assign w6124 = w2600 & w2676;
assign w6125 = ~pi103 & w2675;
assign w6126 = w2611 & w2685;
assign w6127 = ~pi118 & w6126;
assign w6128 = ~w6125 & ~w6127;
assign w6129 = ~w2930 & ~w3140;
assign w6130 = w6128 & w6129;
assign w6131 = pi118 & ~w2601;
assign w6132 = (w2613 & w6131) | (w2613 & w2615) | (w6131 & w2615);
assign w6133 = ~w2640 & ~w3191;
assign w6134 = w2625 & ~w6133;
assign w6135 = w2865 & w3147;
assign w6136 = ~w6134 & ~w6135;
assign w6137 = (~pi034 & ~w6136) | (~pi034 & w18576) | (~w6136 & w18576);
assign w6138 = w2599 & w2660;
assign w6139 = ~w3185 & ~w6138;
assign w6140 = ~pi066 & w2649;
assign w6141 = w2688 & w2855;
assign w6142 = w2677 & w6140;
assign w6143 = ~w6141 & ~w6142;
assign w6144 = pi118 & w2731;
assign w6145 = w6143 & ~w6144;
assign w6146 = (~pi118 & w3185) | (~pi118 & w20786) | (w3185 & w20786);
assign w6147 = w6145 & ~w6146;
assign w6148 = ~w6137 & w6147;
assign w6149 = (~pi038 & ~w6148) | (~pi038 & w18577) | (~w6148 & w18577);
assign w6150 = ~pi103 & w2599;
assign w6151 = ~w2602 & ~w6150;
assign w6152 = (w2643 & ~w6151) | (w2643 & w18578) | (~w6151 & w18578);
assign w6153 = pi118 & w2865;
assign w6154 = w2614 & w3148;
assign w6155 = ~w6153 & ~w6154;
assign w6156 = ~w6152 & w6155;
assign w6157 = pi034 & ~w6156;
assign w6158 = w2609 & w2730;
assign w6159 = ~w3164 & ~w6158;
assign w6160 = w2895 & ~w6159;
assign w6161 = w2650 & w18579;
assign w6162 = ~w3118 & ~w3121;
assign w6163 = w3181 & ~w6162;
assign w6164 = ~pi034 & ~pi118;
assign w6165 = w2639 & w2612;
assign w6166 = w6164 & w6165;
assign w6167 = ~w6163 & ~w6166;
assign w6168 = ~w3123 & ~w3192;
assign w6169 = ~w6161 & w6168;
assign w6170 = w6167 & w6169;
assign w6171 = ~w6160 & w6170;
assign w6172 = ~w6157 & w6171;
assign w6173 = ~w6149 & w6172;
assign w6174 = (pi038 & ~w6121) | (pi038 & w18580) | (~w6121 & w18580);
assign w6175 = w6173 & ~w6174;
assign w6176 = ~w3054 & ~w3061;
assign w6177 = ~pi116 & ~w6176;
assign w6178 = pi116 & w2995;
assign w6179 = w2949 & w6178;
assign w6180 = ~w3034 & ~w6179;
assign w6181 = ~w6177 & w6180;
assign w6182 = (pi058 & ~w6181) | (pi058 & w18581) | (~w6181 & w18581);
assign w6183 = ~w2977 & ~w6023;
assign w6184 = w2961 & w2992;
assign w6185 = ~w6067 & ~w6184;
assign w6186 = (~pi116 & ~w6185) | (~pi116 & w18582) | (~w6185 & w18582);
assign w6187 = pi000 & w2952;
assign w6188 = w2952 & w18583;
assign w6189 = w2969 & w2978;
assign w6190 = ~w3035 & ~w6189;
assign w6191 = (w3090 & ~w6190) | (w3090 & w18584) | (~w6190 & w18584);
assign w6192 = ~pi022 & pi116;
assign w6193 = w2992 & w6192;
assign w6194 = ~w2959 & ~w6193;
assign w6195 = (~pi058 & ~w6194) | (~pi058 & w18585) | (~w6194 & w18585);
assign w6196 = ~pi060 & ~w3093;
assign w6197 = ~w6191 & ~w6195;
assign w6198 = w6196 & w6197;
assign w6199 = ~w2963 & ~w6046;
assign w6200 = ~w2953 & ~w6010;
assign w6201 = w6199 & w6200;
assign w6202 = pi058 & ~w6201;
assign w6203 = w2950 & w3076;
assign w6204 = w2969 & w3006;
assign w6205 = ~w3043 & ~w6203;
assign w6206 = pi000 & w2962;
assign w6207 = ~w3077 & ~w6010;
assign w6208 = w2958 & w3042;
assign w6209 = w2962 & w6015;
assign w6210 = w2965 & w6206;
assign w6211 = w2952 & w3006;
assign w6212 = pi116 & w6211;
assign w6213 = ~w6210 & ~w6212;
assign w6214 = ~w6007 & ~w6208;
assign w6215 = ~w6209 & w6214;
assign w6216 = w6213 & w6215;
assign w6217 = (~pi058 & ~w6216) | (~pi058 & w18587) | (~w6216 & w18587);
assign w6218 = pi000 & w2970;
assign w6219 = w6015 & w6033;
assign w6220 = ~w6218 & ~w6219;
assign w6221 = ~pi000 & w2949;
assign w6222 = w3090 & w6221;
assign w6223 = w6015 & w6206;
assign w6224 = w2995 & w3066;
assign w6225 = ~w6222 & ~w6223;
assign w6226 = pi060 & ~w6224;
assign w6227 = w6225 & w6226;
assign w6228 = pi058 & ~w6220;
assign w6229 = w6227 & ~w6228;
assign w6230 = ~w6217 & w6229;
assign w6231 = (pi116 & w6202) | (pi116 & w18588) | (w6202 & w18588);
assign w6232 = w6230 & ~w6231;
assign w6233 = ~w6182 & w6198;
assign w6234 = ~w6186 & w6233;
assign w6235 = ~w6232 & ~w6234;
assign w6236 = w2953 & w2957;
assign w6237 = ~w3026 & ~w6236;
assign w6238 = w3042 & ~w6084;
assign w6239 = w2953 & w3031;
assign w6240 = ~pi097 & w6239;
assign w6241 = (~pi116 & ~w6068) | (~pi116 & w18589) | (~w6068 & w18589);
assign w6242 = ~w6240 & w6241;
assign w6243 = (pi011 & ~w6237) | (pi011 & w18590) | (~w6237 & w18590);
assign w6244 = w6242 & ~w6243;
assign w6245 = w2952 & w18591;
assign w6246 = ~pi011 & w6245;
assign w6247 = w2962 & w3033;
assign w6248 = ~w6035 & ~w6247;
assign w6249 = ~w2954 & ~w6204;
assign w6250 = pi116 & w6249;
assign w6251 = w6248 & w6250;
assign w6252 = ~w6246 & w6251;
assign w6253 = w2952 & w2958;
assign w6254 = w2995 & w3076;
assign w6255 = ~w2993 & ~w6254;
assign w6256 = ~w6218 & w6255;
assign w6257 = pi116 & w6256;
assign w6258 = w6183 & ~w6253;
assign w6259 = w6242 & w6258;
assign w6260 = ~w6257 & ~w6259;
assign w6261 = ~pi058 & ~w2996;
assign w6262 = ~w6260 & w6261;
assign w6263 = (pi058 & w6252) | (pi058 & w18592) | (w6252 & w18592);
assign w6264 = ~w6262 & ~w6263;
assign w6265 = ~w6235 & ~w6264;
assign w6266 = ~w6175 & w6265;
assign w6267 = w6175 & ~w6265;
assign w6268 = ~w6266 & ~w6267;
assign w6269 = w6101 & w6268;
assign w6270 = ~w6101 & ~w6268;
assign w6271 = ~w6269 & ~w6270;
assign w6272 = ~w3259 & ~w3312;
assign w6273 = ~pi090 & ~w6272;
assign w6274 = pi049 & pi090;
assign w6275 = w3203 & w3284;
assign w6276 = w6274 & w6275;
assign w6277 = ~w3329 & ~w6276;
assign w6278 = ~w6273 & w6277;
assign w6279 = (pi088 & ~w6278) | (pi088 & w18593) | (~w6278 & w18593);
assign w6280 = pi049 & w3263;
assign w6281 = w3248 & w3257;
assign w6282 = ~w3235 & ~w6281;
assign w6283 = pi086 & w3203;
assign w6284 = w3258 & w6283;
assign w6285 = ~w6280 & w6282;
assign w6286 = (~pi090 & ~w6285) | (~pi090 & w18594) | (~w6285 & w18594);
assign w6287 = pi019 & pi090;
assign w6288 = pi049 & w6287;
assign w6289 = ~pi090 & w3245;
assign w6290 = ~w3313 & ~w6289;
assign w6291 = w3238 & w18595;
assign w6292 = w6290 & ~w6291;
assign w6293 = ~w3216 & ~w3301;
assign w6294 = w6288 & ~w6293;
assign w6295 = ~w3342 & ~w6294;
assign w6296 = (~pi088 & ~w6292) | (~pi088 & w18596) | (~w6292 & w18596);
assign w6297 = w6295 & ~w6296;
assign w6298 = ~w6279 & w6297;
assign w6299 = (~pi006 & ~w6298) | (~pi006 & w18597) | (~w6298 & w18597);
assign w6300 = ~pi086 & ~pi112;
assign w6301 = pi049 & w6300;
assign w6302 = pi049 & ~w3207;
assign w6303 = ~w3207 & w18598;
assign w6304 = ~w6301 & ~w6303;
assign w6305 = ~pi090 & ~w3257;
assign w6306 = ~pi090 & w3246;
assign w6307 = w3207 & w3248;
assign w6308 = ~w6306 & ~w6307;
assign w6309 = ~w6305 & ~w6308;
assign w6310 = w3203 & w3250;
assign w6311 = w3214 & w3272;
assign w6312 = w3203 & w3286;
assign w6313 = ~w6310 & ~w6311;
assign w6314 = ~w6312 & w6313;
assign w6315 = ~w6309 & w6314;
assign w6316 = w3203 & w3251;
assign w6317 = w3215 & w3248;
assign w6318 = ~w3289 & ~w6317;
assign w6319 = (pi090 & ~w6318) | (pi090 & w18599) | (~w6318 & w18599);
assign w6320 = w3257 & w3286;
assign w6321 = w3296 & w3341;
assign w6322 = ~w6320 & ~w6321;
assign w6323 = pi049 & w6310;
assign w6324 = w6322 & ~w6323;
assign w6325 = pi049 & w3221;
assign w6326 = w3207 & w3250;
assign w6327 = ~pi112 & w6326;
assign w6328 = ~w6325 & ~w6327;
assign w6329 = ~w3206 & ~w6301;
assign w6330 = ~pi019 & w3238;
assign w6331 = ~w3240 & ~w6330;
assign w6332 = w6329 & w6331;
assign w6333 = w3295 & ~w6332;
assign w6334 = pi088 & ~w6328;
assign w6335 = ~w6333 & ~w6334;
assign w6336 = ~w6319 & w6324;
assign w6337 = w6335 & w6336;
assign w6338 = w3264 & w3272;
assign w6339 = (pi051 & w6301) | (pi051 & w18600) | (w6301 & w18600);
assign w6340 = w3228 & w3257;
assign w6341 = ~w3208 & ~w6340;
assign w6342 = (~pi019 & w6339) | (~pi019 & w18601) | (w6339 & w18601);
assign w6343 = w6341 & ~w6342;
assign w6344 = w3286 & w3246;
assign w6345 = ~w6325 & w18602;
assign w6346 = w3334 & ~w6345;
assign w6347 = w3207 & w3214;
assign w6348 = ~w3335 & ~w6347;
assign w6349 = w6282 & w6348;
assign w6350 = pi090 & ~w3335;
assign w6351 = ~pi019 & w3322;
assign w6352 = w3258 & w3263;
assign w6353 = ~w6351 & ~w6352;
assign w6354 = ~pi090 & ~w6353;
assign w6355 = ~w3247 & ~w3275;
assign w6356 = ~w3245 & w3272;
assign w6357 = pi088 & w3244;
assign w6358 = (w6357 & ~w6355) | (w6357 & w18603) | (~w6355 & w18603);
assign w6359 = ~w6354 & ~w6358;
assign w6360 = (~pi088 & w3335) | (~pi088 & w18604) | (w3335 & w18604);
assign w6361 = ~w6349 & w6360;
assign w6362 = w6359 & w18605;
assign w6363 = w3295 & ~w6343;
assign w6364 = w6362 & ~w6363;
assign w6365 = (pi006 & ~w6337) | (pi006 & w18606) | (~w6337 & w18606);
assign w6366 = w6364 & ~w6365;
assign w6367 = ~w6299 & w6366;
assign w6368 = ~w3229 & ~w3246;
assign w6369 = pi051 & w6368;
assign w6370 = (pi090 & w6369) | (pi090 & w18607) | (w6369 & w18607);
assign w6371 = w3238 & w20787;
assign w6372 = ~w3221 & ~w3252;
assign w6373 = ~w3335 & ~w6310;
assign w6374 = w6372 & w6373;
assign w6375 = ~w6371 & w6374;
assign w6376 = (pi088 & ~w6375) | (pi088 & w18608) | (~w6375 & w18608);
assign w6377 = ~w3285 & ~w3312;
assign w6378 = ~pi090 & ~w6377;
assign w6379 = w3246 & w3248;
assign w6380 = ~w3249 & ~w6379;
assign w6381 = ~w3318 & w6380;
assign w6382 = pi086 & pi090;
assign w6383 = ~w3203 & ~w3264;
assign w6384 = w6382 & ~w6383;
assign w6385 = ~w6378 & w6381;
assign w6386 = ~w3344 & ~w6384;
assign w6387 = w3227 & w3251;
assign w6388 = ~w3281 & ~w6307;
assign w6389 = ~w6387 & w6388;
assign w6390 = ~pi090 & ~w6389;
assign w6391 = ~w3203 & ~w3226;
assign w6392 = ~pi086 & ~w6391;
assign w6393 = (w6274 & w6392) | (w6274 & w18609) | (w6392 & w18609);
assign w6394 = w3214 & w6283;
assign w6395 = ~w6390 & w18610;
assign w6396 = (~pi088 & ~w6385) | (~pi088 & w20788) | (~w6385 & w20788);
assign w6397 = (pi006 & ~w18611) | (pi006 & w20789) | (~w18611 & w20789);
assign w6398 = ~pi051 & w3229;
assign w6399 = ~pi051 & w3286;
assign w6400 = w3246 & w6399;
assign w6401 = w3245 & w3272;
assign w6402 = pi051 & w3248;
assign w6403 = w3246 & w6402;
assign w6404 = ~pi090 & w6401;
assign w6405 = ~w6403 & ~w6404;
assign w6406 = ~w3282 & ~w3343;
assign w6407 = w6405 & w6406;
assign w6408 = ~w3204 & ~w6274;
assign w6409 = w3238 & ~w6408;
assign w6410 = w3244 & w3252;
assign w6411 = w3262 & ~w6300;
assign w6412 = pi051 & w6411;
assign w6413 = ~w6410 & ~w6412;
assign w6414 = ~w6307 & ~w6409;
assign w6415 = w6413 & w6414;
assign w6416 = ~pi088 & ~w6415;
assign w6417 = w3203 & w3258;
assign w6418 = ~w3336 & ~w6417;
assign w6419 = pi090 & w3247;
assign w6420 = w3206 & w3284;
assign w6421 = w3229 & w6287;
assign w6422 = ~w6420 & ~w6421;
assign w6423 = ~pi051 & ~w6422;
assign w6424 = ~w6419 & ~w6423;
assign w6425 = (~pi090 & w3336) | (~pi090 & w18614) | (w3336 & w18614);
assign w6426 = w6424 & ~w6425;
assign w6427 = ~w6416 & w6426;
assign w6428 = (~pi006 & ~w6427) | (~pi006 & w18615) | (~w6427 & w18615);
assign w6429 = ~pi049 & w3203;
assign w6430 = ~w6301 & ~w6401;
assign w6431 = (w3250 & ~w6430) | (w3250 & w18616) | (~w6430 & w18616);
assign w6432 = pi086 & w3214;
assign w6433 = w3214 & w3246;
assign w6434 = ~w3221 & ~w6433;
assign w6435 = pi090 & ~w6434;
assign w6436 = pi090 & w3252;
assign w6437 = w3226 & w3229;
assign w6438 = w3244 & w6437;
assign w6439 = ~w6431 & ~w6435;
assign w6440 = ~w6436 & ~w6438;
assign w6441 = (pi088 & ~w6439) | (pi088 & w18617) | (~w6439 & w18617);
assign w6442 = ~w3228 & w3334;
assign w6443 = (w6442 & w3311) | (w6442 & w18618) | (w3311 & w18618);
assign w6444 = ~pi088 & w6289;
assign w6445 = w3204 & w3226;
assign w6446 = ~w3208 & ~w6445;
assign w6447 = w6287 & ~w6446;
assign w6448 = (w3228 & w6444) | (w3228 & w18619) | (w6444 & w18619);
assign w6449 = ~w6447 & ~w6448;
assign w6450 = ~w6443 & w6449;
assign w6451 = ~w6441 & w6450;
assign w6452 = ~w6428 & w6451;
assign w6453 = ~w6397 & w6452;
assign w6454 = ~w6367 & w6453;
assign w6455 = w6367 & ~w6453;
assign w6456 = ~w6454 & ~w6455;
assign w6457 = w3204 & w3215;
assign w6458 = ~w3249 & ~w6457;
assign w6459 = pi090 & ~pi112;
assign w6460 = w3245 & w6459;
assign w6461 = w3203 & w3262;
assign w6462 = w3228 & w3245;
assign w6463 = w3203 & w6382;
assign w6464 = ~w3323 & ~w6281;
assign w6465 = ~w6463 & w6464;
assign w6466 = ~w6460 & ~w6461;
assign w6467 = ~w6462 & w6466;
assign w6468 = w6465 & w6467;
assign w6469 = (~pi088 & ~w6468) | (~pi088 & w18620) | (~w6468 & w18620);
assign w6470 = ~pi049 & w3238;
assign w6471 = (pi090 & ~w3238) | (pi090 & w6274) | (~w3238 & w6274);
assign w6472 = pi088 & ~w6471;
assign w6473 = ~w6394 & w18621;
assign w6474 = w6472 & ~w6473;
assign w6475 = (w6287 & ~w6293) | (w6287 & w18622) | (~w6293 & w18622);
assign w6476 = ~w3249 & ~w6461;
assign w6477 = pi086 & ~w6476;
assign w6478 = w3227 & w3229;
assign w6479 = (pi006 & ~w3227) | (pi006 & w18623) | (~w3227 & w18623);
assign w6480 = ~w6477 & w6479;
assign w6481 = ~w6475 & w6480;
assign w6482 = ~w6474 & w6481;
assign w6483 = ~w6469 & w6482;
assign w6484 = w3203 & w3214;
assign w6485 = ~w6330 & ~w6484;
assign w6486 = pi090 & ~w6485;
assign w6487 = ~w3228 & ~w3264;
assign w6488 = w6305 & ~w6487;
assign w6489 = ~w3300 & ~w6488;
assign w6490 = ~w6486 & w6489;
assign w6491 = pi088 & ~w6490;
assign w6492 = w3244 & w3257;
assign w6493 = ~w3335 & ~w6492;
assign w6494 = w3244 & w6338;
assign w6495 = w6287 & w6457;
assign w6496 = ~pi006 & ~w3252;
assign w6497 = ~w6494 & ~w6495;
assign w6498 = w6496 & w6497;
assign w6499 = ~pi088 & ~w6493;
assign w6500 = w6498 & ~w6499;
assign w6501 = ~w6491 & w6500;
assign w6502 = ~w6483 & ~w6501;
assign w6503 = ~pi090 & ~w6338;
assign w6504 = w3226 & w3258;
assign w6505 = ~w6284 & w6503;
assign w6506 = ~w3323 & ~w6504;
assign w6507 = w6505 & w6506;
assign w6508 = ~pi086 & w3299;
assign w6509 = ~w3217 & w6350;
assign w6510 = ~w6508 & w6509;
assign w6511 = ~w6507 & ~w6510;
assign w6512 = w3299 & w3204;
assign w6513 = ~w6437 & ~w6512;
assign w6514 = (~pi088 & w6511) | (~pi088 & w18624) | (w6511 & w18624);
assign w6515 = w3226 & w3286;
assign w6516 = ~pi049 & w3220;
assign w6517 = w3203 & w6516;
assign w6518 = ~w6402 & ~w6457;
assign w6519 = ~w6517 & w6518;
assign w6520 = pi090 & w6519;
assign w6521 = ~pi090 & ~w6515;
assign w6522 = w3283 & w6521;
assign w6523 = ~w6520 & ~w6522;
assign w6524 = (pi088 & w6523) | (pi088 & w18625) | (w6523 & w18625);
assign w6525 = ~pi051 & w3273;
assign w6526 = (pi090 & w6525) | (pi090 & w18626) | (w6525 & w18626);
assign w6527 = ~w6514 & ~w6524;
assign w6528 = ~w6438 & ~w6526;
assign w6529 = w6527 & w6528;
assign w6530 = ~w6502 & w6529;
assign w6531 = ~pi171 & w6530;
assign w6532 = pi171 & ~w6530;
assign w6533 = ~w6531 & ~w6532;
assign w6534 = w6456 & w6533;
assign w6535 = ~w6456 & ~w6533;
assign w6536 = ~w6534 & ~w6535;
assign w6537 = w6271 & w6536;
assign w6538 = ~pi529 & ~w6537;
assign w6539 = ~w6271 & ~w6536;
assign w6540 = w6538 & ~w6539;
assign w6541 = ~pi171 & pi443;
assign w6542 = pi529 & ~w6541;
assign w6543 = pi171 & ~pi443;
assign w6544 = w6542 & ~w6543;
assign w6545 = ~w6540 & ~w6544;
assign w6546 = w6366 & w18627;
assign w6547 = (pi187 & ~w6366) | (pi187 & w18628) | (~w6366 & w18628);
assign w6548 = ~w6546 & ~w6547;
assign w6549 = ~w2596 & w2849;
assign w6550 = w2596 & ~w2849;
assign w6551 = ~w6549 & ~w6550;
assign w6552 = w2992 & w3039;
assign w6553 = ~w3081 & ~w6203;
assign w6554 = (pi116 & ~w6553) | (pi116 & w18629) | (~w6553 & w18629);
assign w6555 = pi022 & ~w2982;
assign w6556 = w2958 & ~w6555;
assign w6557 = ~w6023 & ~w6556;
assign w6558 = ~w6554 & w6557;
assign w6559 = ~w2959 & ~w3059;
assign w6560 = ~w2997 & ~w6073;
assign w6561 = w6559 & w6560;
assign w6562 = (~pi116 & w3001) | (~pi116 & w18630) | (w3001 & w18630);
assign w6563 = (pi058 & w6562) | (pi058 & w18631) | (w6562 & w18631);
assign w6564 = ~w6189 & ~w6224;
assign w6565 = ~pi116 & ~w6564;
assign w6566 = ~w2949 & ~w3000;
assign w6567 = w3027 & ~w6566;
assign w6568 = ~pi000 & w3060;
assign w6569 = w2952 & w6568;
assign w6570 = ~w6567 & ~w6569;
assign w6571 = ~w6565 & w6570;
assign w6572 = ~w3032 & w6571;
assign w6573 = (~w6563 & w6561) | (~w6563 & w18632) | (w6561 & w18632);
assign w6574 = w6572 & w6573;
assign w6575 = w2969 & w3033;
assign w6576 = w2980 & w3006;
assign w6577 = ~w2997 & w18634;
assign w6578 = ~pi116 & ~w6577;
assign w6579 = ~w2977 & ~w3021;
assign w6580 = w3083 & ~w6579;
assign w6581 = w3090 & w6009;
assign w6582 = w6009 & w18635;
assign w6583 = ~w6222 & ~w6582;
assign w6584 = ~pi116 & w3004;
assign w6585 = ~pi011 & ~w6237;
assign w6586 = ~w2984 & ~w2992;
assign w6587 = ~w3024 & ~w6586;
assign w6588 = w2963 & w3003;
assign w6589 = w2952 & w6015;
assign w6590 = ~w6588 & ~w6589;
assign w6591 = ~w6585 & w18636;
assign w6592 = pi058 & ~w6587;
assign w6593 = w6590 & w6592;
assign w6594 = ~w6591 & ~w6593;
assign w6595 = ~w6580 & w6583;
assign w6596 = ~w6578 & w6595;
assign w6597 = ~w6594 & w6596;
assign w6598 = pi116 & ~w3095;
assign w6599 = w2949 & w3052;
assign w6600 = ~pi116 & ~w2996;
assign w6601 = w6598 & ~w6599;
assign w6602 = ~w6600 & ~w6601;
assign w6603 = ~pi011 & w3071;
assign w6604 = ~w6057 & ~w6603;
assign w6605 = (pi058 & w6602) | (pi058 & w18637) | (w6602 & w18637);
assign w6606 = ~w2995 & ~w3039;
assign w6607 = w2962 & ~w6606;
assign w6608 = ~w6035 & ~w6607;
assign w6609 = ~pi116 & ~w6608;
assign w6610 = ~w3076 & ~w6033;
assign w6611 = w6089 & ~w6610;
assign w6612 = ~w3005 & ~w6008;
assign w6613 = ~w6611 & w6612;
assign w6614 = ~w6609 & w6613;
assign w6615 = w2984 & w18638;
assign w6616 = w2966 & w6089;
assign w6617 = pi057 & w6615;
assign w6618 = ~w6616 & ~w6617;
assign w6619 = (w6618 & w6614) | (w6618 & w18639) | (w6614 & w18639);
assign w6620 = ~w6605 & w6619;
assign w6621 = ~pi060 & ~w6597;
assign w6622 = w6620 & ~w6621;
assign w6623 = (pi060 & ~w6574) | (pi060 & w18640) | (~w6574 & w18640);
assign w6624 = w6622 & ~w6623;
assign w6625 = ~w2942 & w6624;
assign w6626 = w2942 & ~w6624;
assign w6627 = ~w6625 & ~w6626;
assign w6628 = w6551 & ~w6627;
assign w6629 = ~w6551 & w6627;
assign w6630 = ~w6628 & ~w6629;
assign w6631 = ~w6548 & w6630;
assign w6632 = w6548 & ~w6630;
assign w6633 = ~w6631 & ~w6632;
assign w6634 = ~pi187 & pi439;
assign w6635 = pi187 & ~pi439;
assign w6636 = ~w6634 & ~w6635;
assign w6637 = ~w6005 & w6175;
assign w6638 = w6005 & ~w6175;
assign w6639 = ~w6637 & ~w6638;
assign w6640 = w2747 & ~w6639;
assign w6641 = ~w2747 & w6639;
assign w6642 = ~w6640 & ~w6641;
assign w6643 = ~w2729 & ~w6138;
assign w6644 = w2609 & w2683;
assign w6645 = w6643 & ~w6644;
assign w6646 = ~w2918 & w3155;
assign w6647 = w2597 & w3191;
assign w6648 = w2612 & w2625;
assign w6649 = ~w2689 & ~w6647;
assign w6650 = ~w6648 & w6649;
assign w6651 = w2643 & w2673;
assign w6652 = ~w2650 & ~w2902;
assign w6653 = ~w2609 & ~w2689;
assign w6654 = ~w6652 & ~w6653;
assign w6655 = w2664 & w18641;
assign w6656 = (~pi038 & ~w2739) | (~pi038 & w18642) | (~w2739 & w18642);
assign w6657 = ~w6654 & w18643;
assign w6658 = (~pi034 & ~w6650) | (~pi034 & w20790) | (~w6650 & w20790);
assign w6659 = w6657 & ~w6658;
assign w6660 = (pi034 & ~w6645) | (pi034 & w18644) | (~w6645 & w18644);
assign w6661 = w6659 & ~w6660;
assign w6662 = ~pi118 & ~w2625;
assign w6663 = ~w2899 & ~w3164;
assign w6664 = w2669 & w18645;
assign w6665 = w6663 & ~w6664;
assign w6666 = (pi034 & ~w6665) | (pi034 & w18646) | (~w6665 & w18646);
assign w6667 = ~pi062 & w2612;
assign w6668 = ~pi119 & w2632;
assign w6669 = ~w2731 & ~w6668;
assign w6670 = w2599 & w2612;
assign w6671 = ~w3118 & ~w6670;
assign w6672 = ~pi118 & w6671;
assign w6673 = ~w2929 & w6672;
assign w6674 = w2931 & w6669;
assign w6675 = ~w6667 & w6674;
assign w6676 = ~w6673 & ~w6675;
assign w6677 = pi066 & w2713;
assign w6678 = w2853 & w2922;
assign w6679 = ~w6677 & ~w6678;
assign w6680 = ~w2903 & ~w6153;
assign w6681 = ~w6165 & w6679;
assign w6682 = w6680 & w6681;
assign w6683 = (pi038 & w6682) | (pi038 & w18647) | (w6682 & w18647);
assign w6684 = ~w6666 & w6683;
assign w6685 = ~w6676 & w6684;
assign w6686 = ~w6661 & ~w6685;
assign w6687 = ~w2624 & ~w6667;
assign w6688 = pi101 & ~w6687;
assign w6689 = ~w2914 & ~w3169;
assign w6690 = ~w6688 & w6689;
assign w6691 = ~w2677 & w6140;
assign w6692 = ~w3122 & ~w6691;
assign w6693 = ~w2674 & ~w2740;
assign w6694 = ~pi118 & ~w6692;
assign w6695 = w6693 & ~w6694;
assign w6696 = (pi118 & ~w6690) | (pi118 & w18568) | (~w6690 & w18568);
assign w6697 = w6695 & ~w6696;
assign w6698 = ~w2929 & ~w6125;
assign w6699 = ~pi118 & ~w6698;
assign w6700 = ~w2882 & ~w6662;
assign w6701 = w2605 & ~w6700;
assign w6702 = w2611 & w2698;
assign w6703 = ~w2610 & ~w2642;
assign w6704 = ~w6701 & w6703;
assign w6705 = ~w6702 & w6704;
assign w6706 = ~pi118 & w2730;
assign w6707 = (pi066 & w6706) | (pi066 & w18648) | (w6706 & w18648);
assign w6708 = (w6705 & w20791) | (w6705 & w20792) | (w20791 & w20792);
assign w6709 = ~pi034 & ~w6697;
assign w6710 = w6708 & ~w6709;
assign w6711 = ~w6686 & w6710;
assign w6712 = w2968 & ~w2992;
assign w6713 = pi097 & w6239;
assign w6714 = ~w6712 & ~w6713;
assign w6715 = (~pi116 & ~w6714) | (~pi116 & w18650) | (~w6714 & w18650);
assign w6716 = w3077 & w3090;
assign w6717 = w3054 & w3041;
assign w6718 = ~w6716 & ~w6717;
assign w6719 = w3058 & w3090;
assign w6720 = ~w6218 & ~w6569;
assign w6721 = ~w6719 & w6720;
assign w6722 = (pi058 & ~w6206) | (pi058 & w18651) | (~w6206 & w18651);
assign w6723 = w6721 & w18652;
assign w6724 = (pi022 & ~w6199) | (pi022 & w18653) | (~w6199 & w18653);
assign w6725 = ~w3062 & ~w6034;
assign w6726 = ~w6724 & w6725;
assign w6727 = pi116 & ~w6726;
assign w6728 = ~w2960 & ~w6599;
assign w6729 = (~pi116 & ~w6728) | (~pi116 & w18654) | (~w6728 & w18654);
assign w6730 = ~w6035 & ~w6067;
assign w6731 = ~pi058 & w6730;
assign w6732 = w6718 & w6731;
assign w6733 = ~w6729 & w6732;
assign w6734 = ~w6727 & w6733;
assign w6735 = ~w6715 & w6723;
assign w6736 = ~w6734 & ~w6735;
assign w6737 = pi011 & w2957;
assign w6738 = w3041 & w2957;
assign w6739 = ~w6584 & ~w6738;
assign w6740 = w3021 & w3094;
assign w6741 = (~pi058 & ~w2957) | (~pi058 & w18655) | (~w2957 & w18655);
assign w6742 = ~w6021 & w6741;
assign w6743 = w6739 & w18656;
assign w6744 = ~pi000 & w2962;
assign w6745 = ~w6245 & ~w6744;
assign w6746 = ~pi116 & ~w6745;
assign w6747 = ~w3053 & ~w6017;
assign w6748 = (pi058 & ~w6056) | (pi058 & w18657) | (~w6056 & w18657);
assign w6749 = w6747 & w6748;
assign w6750 = ~w6746 & w6749;
assign w6751 = ~w6743 & ~w6750;
assign w6752 = ~w3052 & ~w6236;
assign w6753 = w6598 & w6752;
assign w6754 = ~w6568 & w6753;
assign w6755 = ~w2970 & ~w6045;
assign w6756 = ~pi116 & w6755;
assign w6757 = ~w6603 & w6756;
assign w6758 = ~w6754 & ~w6757;
assign w6759 = pi060 & ~w6758;
assign w6760 = (w3076 & w6209) | (w3076 & w18658) | (w6209 & w18658);
assign w6761 = ~pi097 & w6568;
assign w6762 = ~pi058 & ~w6193;
assign w6763 = ~w6761 & w6762;
assign w6764 = ~w6760 & w6763;
assign w6765 = pi022 & w2958;
assign w6766 = ~w2961 & w2982;
assign w6767 = ~w6765 & w6766;
assign w6768 = ~pi116 & w6767;
assign w6769 = w2962 & w2984;
assign w6770 = pi058 & ~w6769;
assign w6771 = ~w6020 & w6770;
assign w6772 = w2965 & w6187;
assign w6773 = w6771 & ~w6772;
assign w6774 = ~w6768 & w6773;
assign w6775 = ~w3004 & ~w6221;
assign w6776 = pi116 & ~w6775;
assign w6777 = (pi011 & ~w2992) | (pi011 & w3033) | (~w2992 & w3033);
assign w6778 = ~w6775 & w18659;
assign w6779 = w3081 & w6015;
assign w6780 = (~pi060 & ~w6009) | (~pi060 & w18660) | (~w6009 & w18660);
assign w6781 = ~w6779 & w6780;
assign w6782 = ~w6778 & w6781;
assign w6783 = ~w6751 & w6759;
assign w6784 = (w6782 & w6774) | (w6782 & w18661) | (w6774 & w18661);
assign w6785 = ~w6783 & ~w6784;
assign w6786 = ~w6736 & ~w6785;
assign w6787 = ~w6711 & w6786;
assign w6788 = w6711 & ~w6786;
assign w6789 = ~w6787 & ~w6788;
assign w6790 = ~w6429 & ~w6445;
assign w6791 = ~pi090 & ~w6790;
assign w6792 = w3214 & w3238;
assign w6793 = pi086 & w6792;
assign w6794 = ~w3311 & ~w6793;
assign w6795 = ~w6791 & w6794;
assign w6796 = (pi088 & ~w6795) | (pi088 & w18662) | (~w6795 & w18662);
assign w6797 = ~w3247 & ~w6399;
assign w6798 = pi090 & w6797;
assign w6799 = w3299 & ~w6302;
assign w6800 = w6798 & ~w6799;
assign w6801 = w3238 & w3284;
assign w6802 = ~pi049 & w6801;
assign w6803 = ~pi090 & ~w3221;
assign w6804 = ~w6802 & w6803;
assign w6805 = ~w6484 & w6804;
assign w6806 = ~w6800 & ~w6805;
assign w6807 = pi019 & w3280;
assign w6808 = w3238 & w3258;
assign w6809 = ~pi090 & w6808;
assign w6810 = w3245 & w18663;
assign w6811 = ~w6809 & ~w6810;
assign w6812 = ~w6462 & ~w6807;
assign w6813 = ~w6436 & w6812;
assign w6814 = w6811 & w6813;
assign w6815 = (pi006 & w6814) | (pi006 & w18664) | (w6814 & w18664);
assign w6816 = ~pi090 & w3226;
assign w6817 = pi090 & w3286;
assign w6818 = ~w6417 & ~w6463;
assign w6819 = w3207 & w6817;
assign w6820 = w6818 & ~w6819;
assign w6821 = ~w6432 & w6816;
assign w6822 = ~w3204 & w6821;
assign w6823 = w6820 & ~w6822;
assign w6824 = ~w3263 & ~w3330;
assign w6825 = pi090 & ~w6824;
assign w6826 = pi086 & w6310;
assign w6827 = ~w6792 & ~w6826;
assign w6828 = ~w6825 & w6827;
assign w6829 = ~pi088 & ~w6828;
assign w6830 = (pi090 & w6352) | (pi090 & w18665) | (w6352 & w18665);
assign w6831 = w3287 & w20793;
assign w6832 = (~pi006 & ~w3273) | (~pi006 & w18666) | (~w3273 & w18666);
assign w6833 = ~w6831 & w6832;
assign w6834 = ~w6830 & w6833;
assign w6835 = ~w6829 & w6834;
assign w6836 = pi088 & ~w6823;
assign w6837 = w6835 & ~w6836;
assign w6838 = ~w6796 & w6815;
assign w6839 = ~w6806 & w6838;
assign w6840 = ~w6837 & ~w6839;
assign w6841 = ~w3318 & ~w6478;
assign w6842 = ~w6311 & w6841;
assign w6843 = ~pi051 & w3296;
assign w6844 = w3286 & w6843;
assign w6845 = ~w3217 & ~w6844;
assign w6846 = (~pi090 & ~w6845) | (~pi090 & w10236) | (~w6845 & w10236);
assign w6847 = w3330 & w6287;
assign w6848 = w6516 & w18667;
assign w6849 = ~w6847 & ~w6848;
assign w6850 = ~w6284 & ~w6525;
assign w6851 = ~pi088 & w6850;
assign w6852 = w6849 & w6851;
assign w6853 = ~w6846 & w6852;
assign w6854 = (pi090 & ~w6842) | (pi090 & w18668) | (~w6842 & w18668);
assign w6855 = w6853 & ~w6854;
assign w6856 = w3220 & ~w3238;
assign w6857 = ~w6403 & ~w6856;
assign w6858 = (~pi090 & ~w6857) | (~pi090 & w18669) | (~w6857 & w18669);
assign w6859 = pi086 & w3238;
assign w6860 = w6287 & w6859;
assign w6861 = w3229 & w3317;
assign w6862 = ~w6860 & ~w6861;
assign w6863 = pi049 & w6461;
assign w6864 = w6862 & ~w6863;
assign w6865 = (pi088 & ~w3221) | (pi088 & w18670) | (~w3221 & w18670);
assign w6866 = w6864 & w18671;
assign w6867 = ~w6858 & w6866;
assign w6868 = ~w6855 & ~w6867;
assign w6869 = ~w6840 & ~w6868;
assign w6870 = ~pi255 & w6869;
assign w6871 = pi255 & ~w6869;
assign w6872 = ~w6870 & ~w6871;
assign w6873 = w6789 & w6872;
assign w6874 = ~w6789 & ~w6872;
assign w6875 = ~w6873 & ~w6874;
assign w6876 = ~w6642 & w6875;
assign w6877 = ~pi529 & ~w6876;
assign w6878 = w6642 & ~w6875;
assign w6879 = w6877 & ~w6878;
assign w6880 = ~pi255 & pi505;
assign w6881 = pi529 & ~w6880;
assign w6882 = pi255 & ~pi505;
assign w6883 = w6881 & ~w6882;
assign w6884 = ~w6879 & ~w6883;
assign w6885 = ~w6316 & ~w6457;
assign w6886 = (pi090 & ~w6885) | (pi090 & w18672) | (~w6885 & w18672);
assign w6887 = w3214 & w3226;
assign w6888 = ~w6281 & ~w6516;
assign w6889 = ~w6887 & w6888;
assign w6890 = w3250 & w6445;
assign w6891 = w6889 & ~w6890;
assign w6892 = (~pi088 & ~w6891) | (~pi088 & w18673) | (~w6891 & w18673);
assign w6893 = ~w3260 & ~w3313;
assign w6894 = ~w6387 & ~w6437;
assign w6895 = w6893 & w6894;
assign w6896 = pi090 & ~w6895;
assign w6897 = ~w3205 & ~w6306;
assign w6898 = (pi088 & ~w6897) | (pi088 & w20794) | (~w6897 & w20794);
assign w6899 = ~w3264 & ~w3296;
assign w6900 = pi019 & ~w6899;
assign w6901 = w3215 & w3251;
assign w6902 = ~w6320 & ~w6901;
assign w6903 = ~w6900 & w6902;
assign w6904 = ~pi090 & ~w6903;
assign w6905 = ~w3219 & ~w6861;
assign w6906 = ~w6904 & w20795;
assign w6907 = (pi006 & ~w18674) | (pi006 & w20796) | (~w18674 & w20796);
assign w6908 = pi051 & w3258;
assign w6909 = ~w6463 & ~w6908;
assign w6910 = w3228 & ~w6909;
assign w6911 = ~w6326 & ~w6330;
assign w6912 = ~w6470 & w6911;
assign w6913 = ~w6910 & w6912;
assign w6914 = ~pi019 & ~w6355;
assign w6915 = ~w3296 & ~w6859;
assign w6916 = w3341 & ~w6915;
assign w6917 = w3248 & w6300;
assign w6918 = ~w3281 & ~w6917;
assign w6919 = ~pi090 & ~w6918;
assign w6920 = w3280 & w6442;
assign w6921 = ~w3253 & ~w6920;
assign w6922 = ~w6916 & ~w6919;
assign w6923 = w6921 & w6922;
assign w6924 = (~pi088 & w6914) | (~pi088 & w18675) | (w6914 & w18675);
assign w6925 = w6923 & ~w6924;
assign w6926 = (~pi006 & ~w6925) | (~pi006 & w18676) | (~w6925 & w18676);
assign w6927 = ~w6793 & ~w6802;
assign w6928 = w3234 & w3250;
assign w6929 = w6927 & ~w6928;
assign w6930 = ~w3344 & ~w6276;
assign w6931 = (pi088 & ~w6929) | (pi088 & w18677) | (~w6929 & w18677);
assign w6932 = ~w3260 & ~w6478;
assign w6933 = pi090 & ~w6379;
assign w6934 = w6932 & w6933;
assign w6935 = ~w6275 & ~w6312;
assign w6936 = ~pi090 & w6935;
assign w6937 = ~w6394 & ~w6525;
assign w6938 = w6936 & w6937;
assign w6939 = ~pi088 & ~w6938;
assign w6940 = w3258 & w18678;
assign w6941 = w3203 & w3248;
assign w6942 = pi112 & w6940;
assign w6943 = w6382 & w6941;
assign w6944 = ~w6942 & ~w6943;
assign w6945 = (w6944 & ~w6939) | (w6944 & w18679) | (~w6939 & w18679);
assign w6946 = ~w6931 & w6945;
assign w6947 = ~w6926 & w6946;
assign w6948 = ~w6907 & w6947;
assign w6949 = ~pi189 & w6948;
assign w6950 = pi189 & ~w6948;
assign w6951 = ~w6949 & ~w6950;
assign w6952 = ~w6265 & w6624;
assign w6953 = w6265 & ~w6624;
assign w6954 = ~w6952 & ~w6953;
assign w6955 = ~w2744 & w2849;
assign w6956 = w2744 & ~w2849;
assign w6957 = ~w6955 & ~w6956;
assign w6958 = w6954 & w6957;
assign w6959 = ~w6954 & ~w6957;
assign w6960 = ~w6958 & ~w6959;
assign w6961 = (~pi529 & ~w6960) | (~pi529 & w18680) | (~w6960 & w18680);
assign w6962 = ~w6951 & ~w6960;
assign w6963 = w6961 & ~w6962;
assign w6964 = pi189 & pi496;
assign w6965 = pi529 & ~w6964;
assign w6966 = ~pi189 & ~pi496;
assign w6967 = w6965 & ~w6966;
assign w6968 = ~w6963 & ~w6967;
assign w6969 = w4144 & w18681;
assign w6970 = ~w4163 & ~w4664;
assign w6971 = (pi113 & ~w6970) | (pi113 & w18682) | (~w6970 & w18682);
assign w6972 = w4126 & w4127;
assign w6973 = ~w4668 & ~w4710;
assign w6974 = ~w6972 & w6973;
assign w6975 = w4150 & w4175;
assign w6976 = w6974 & ~w6975;
assign w6977 = (~pi096 & ~w6976) | (~pi096 & w18683) | (~w6976 & w18683);
assign w6978 = (pi096 & w4145) | (pi096 & w18684) | (w4145 & w18684);
assign w6979 = ~pi124 & w4127;
assign w6980 = ~w4680 & ~w4681;
assign w6981 = ~w4700 & ~w6979;
assign w6982 = w6980 & w6981;
assign w6983 = (~pi113 & ~w6982) | (~pi113 & w18685) | (~w6982 & w18685);
assign w6984 = w4156 & w4183;
assign w6985 = w4127 & w4192;
assign w6986 = ~w6984 & ~w6985;
assign w6987 = w4134 & w18686;
assign w6988 = ~w4571 & ~w6987;
assign w6989 = w6986 & w6988;
assign w6990 = pi113 & ~w6989;
assign w6991 = pi096 & w4627;
assign w6992 = w4138 & w4166;
assign w6993 = ~w4235 & ~w6991;
assign w6994 = ~w6992 & w6993;
assign w6995 = ~w6990 & w6994;
assign w6996 = w6995 & w18687;
assign w6997 = ~pi010 & ~w6996;
assign w6998 = (~w4555 & w4705) | (~w4555 & w18688) | (w4705 & w18688);
assign w6999 = ~pi009 & ~w4735;
assign w7000 = w4158 & w4263;
assign w7001 = ~w4573 & ~w7000;
assign w7002 = ~w4571 & w7001;
assign w7003 = ~pi113 & ~w7002;
assign w7004 = ~w4226 & ~w4546;
assign w7005 = w4632 & ~w7004;
assign w7006 = ~w4159 & ~w4237;
assign w7007 = w4706 & ~w7006;
assign w7008 = ~w7005 & ~w7007;
assign w7009 = ~w7003 & w7008;
assign w7010 = (~pi096 & w6999) | (~pi096 & w18689) | (w6999 & w18689);
assign w7011 = w7009 & ~w7010;
assign w7012 = (pi096 & ~w6998) | (pi096 & w18690) | (~w6998 & w18690);
assign w7013 = (pi010 & ~w7011) | (pi010 & w18691) | (~w7011 & w18691);
assign w7014 = (pi113 & w4265) | (pi113 & w18692) | (w4265 & w18692);
assign w7015 = w4236 & w4701;
assign w7016 = ~w4168 & ~w4578;
assign w7017 = ~w4189 & w4548;
assign w7018 = (pi113 & ~w4701) | (pi113 & w18693) | (~w4701 & w18693);
assign w7019 = ~w7015 & ~w7017;
assign w7020 = w7016 & w7019;
assign w7021 = (~w7014 & w7020) | (~w7014 & w18694) | (w7020 & w18694);
assign w7022 = ~pi096 & ~w7021;
assign w7023 = (~pi113 & ~w4162) | (~pi113 & w4150) | (~w4162 & w4150);
assign w7024 = w4137 & w4188;
assign w7025 = (~w7023 & w4732) | (~w7023 & w18695) | (w4732 & w18695);
assign w7026 = ~pi113 & ~w4552;
assign w7027 = ~w4206 & ~w7026;
assign w7028 = w4138 & w4594;
assign w7029 = ~w4184 & ~w4217;
assign w7030 = ~w7027 & w7029;
assign w7031 = (w7030 & w20797) | (w7030 & w20798) | (w20797 & w20798);
assign w7032 = ~w7022 & w7031;
assign w7033 = ~w7013 & w7032;
assign w7034 = ~w6997 & w7033;
assign w7035 = ~pi139 & w7034;
assign w7036 = pi139 & ~w7034;
assign w7037 = ~w7035 & ~w7036;
assign w7038 = w3663 & ~w4988;
assign w7039 = ~w3663 & w4988;
assign w7040 = ~w7038 & ~w7039;
assign w7041 = (~pi529 & w7040) | (~pi529 & w18697) | (w7040 & w18697);
assign w7042 = ~w7037 & w7040;
assign w7043 = w7041 & ~w7042;
assign w7044 = pi139 & pi418;
assign w7045 = pi529 & ~w7044;
assign w7046 = ~pi139 & ~pi418;
assign w7047 = w7045 & ~w7046;
assign w7048 = ~w7043 & ~w7047;
assign w7049 = ~w3660 & w4440;
assign w7050 = w3660 & ~w4440;
assign w7051 = ~w7049 & ~w7050;
assign w7052 = w3876 & w7051;
assign w7053 = ~w3876 & ~w7051;
assign w7054 = ~w7052 & ~w7053;
assign w7055 = ~pi113 & w4561;
assign w7056 = ~w4133 & ~w7055;
assign w7057 = ~w4167 & ~w4182;
assign w7058 = ~w4164 & w7057;
assign w7059 = w7056 & w7058;
assign w7060 = ~w4194 & ~w4710;
assign w7061 = w4124 & w4213;
assign w7062 = ~pi125 & w4144;
assign w7063 = w4144 & w18698;
assign w7064 = ~w7061 & ~w7063;
assign w7065 = ~w4573 & ~w6984;
assign w7066 = w7064 & w7065;
assign w7067 = pi113 & ~w7066;
assign w7068 = ~w4606 & ~w4618;
assign w7069 = ~w4578 & w7068;
assign w7070 = w4738 & ~w7069;
assign w7071 = pi025 & w7028;
assign w7072 = ~w4168 & ~w4265;
assign w7073 = (~pi010 & ~w7028) | (~pi010 & w18699) | (~w7028 & w18699);
assign w7074 = w7072 & w7073;
assign w7075 = ~w7070 & w7074;
assign w7076 = ~w7067 & w7075;
assign w7077 = (~pi096 & ~w7059) | (~pi096 & w18700) | (~w7059 & w18700);
assign w7078 = w7076 & ~w7077;
assign w7079 = (pi113 & ~w4144) | (pi113 & w4236) | (~w4144 & w4236);
assign w7080 = ~w4214 & w7079;
assign w7081 = ~w4583 & ~w4680;
assign w7082 = w7023 & w7081;
assign w7083 = (~w4692 & w7082) | (~w4692 & w18701) | (w7082 & w18701);
assign w7084 = pi096 & ~w7083;
assign w7085 = w4149 & w18702;
assign w7086 = w4183 & w4241;
assign w7087 = ~w4552 & ~w7086;
assign w7088 = pi010 & ~w4198;
assign w7089 = w4163 & w4236;
assign w7090 = w7088 & ~w7089;
assign w7091 = ~pi096 & ~w7087;
assign w7092 = w7090 & ~w7091;
assign w7093 = ~w7085 & w7092;
assign w7094 = ~w7084 & w7093;
assign w7095 = ~w7078 & ~w7094;
assign w7096 = (~pi113 & ~w4586) | (~pi113 & w18703) | (~w4586 & w18703);
assign w7097 = w4126 & w4207;
assign w7098 = ~w4729 & ~w7097;
assign w7099 = ~w4163 & ~w4662;
assign w7100 = pi113 & w7099;
assign w7101 = ~pi125 & w4559;
assign w7102 = w7100 & ~w7101;
assign w7103 = w7096 & w7098;
assign w7104 = (~w4254 & w7102) | (~w4254 & w18704) | (w7102 & w18704);
assign w7105 = pi096 & ~w7104;
assign w7106 = ~pi125 & w4183;
assign w7107 = ~w4704 & ~w7106;
assign w7108 = ~pi055 & ~w7107;
assign w7109 = ~pi055 & w4204;
assign w7110 = ~w4552 & ~w7109;
assign w7111 = ~w4252 & w7110;
assign w7112 = pi113 & ~w7111;
assign w7113 = ~pi113 & w4167;
assign w7114 = w4137 & w4263;
assign w7115 = ~w6987 & ~w7114;
assign w7116 = ~w7113 & w7115;
assign w7117 = ~w7112 & w7116;
assign w7118 = (~pi096 & ~w7117) | (~pi096 & w18706) | (~w7117 & w18706);
assign w7119 = (pi113 & w4168) | (pi113 & w18707) | (w4168 & w18707);
assign w7120 = ~w7105 & ~w7118;
assign w7121 = ~w4623 & ~w7119;
assign w7122 = w7120 & w7121;
assign w7123 = ~w7095 & w7122;
assign w7124 = ~pi182 & w7123;
assign w7125 = pi182 & ~w7123;
assign w7126 = ~w7124 & ~w7125;
assign w7127 = ~w4540 & w4749;
assign w7128 = w4540 & ~w4749;
assign w7129 = ~w7127 & ~w7128;
assign w7130 = w7126 & w7129;
assign w7131 = ~w7126 & ~w7129;
assign w7132 = ~w7130 & ~w7131;
assign w7133 = w7054 & w7132;
assign w7134 = ~pi529 & ~w7133;
assign w7135 = ~w7054 & ~w7132;
assign w7136 = w7134 & ~w7135;
assign w7137 = ~pi182 & pi436;
assign w7138 = pi529 & ~w7137;
assign w7139 = pi182 & ~pi436;
assign w7140 = w7138 & ~w7139;
assign w7141 = ~w7136 & ~w7140;
assign w7142 = ~pi193 & w7034;
assign w7143 = pi193 & ~w7034;
assign w7144 = ~w7142 & ~w7143;
assign w7145 = ~pi106 & ~w4837;
assign w7146 = w3975 & w4532;
assign w7147 = (~w7145 & ~w7146) | (~w7145 & w18708) | (~w7146 & w18708);
assign w7148 = (pi065 & w7147) | (pi065 & w18709) | (w7147 & w18709);
assign w7149 = ~w3988 & ~w4098;
assign w7150 = (w3973 & ~w7149) | (w3973 & w18711) | (~w7149 & w18711);
assign w7151 = pi106 & w4466;
assign w7152 = w3995 & w4467;
assign w7153 = ~w7151 & ~w7152;
assign w7154 = ~w7150 & w7153;
assign w7155 = (~pi065 & ~w7154) | (~pi065 & w18712) | (~w7154 & w18712);
assign w7156 = pi128 & w3978;
assign w7157 = ~w4841 & ~w7156;
assign w7158 = pi100 & ~w7157;
assign w7159 = ~w4468 & ~w4833;
assign w7160 = (pi106 & w7158) | (pi106 & w18713) | (w7158 & w18713);
assign w7161 = pi031 & w4099;
assign w7162 = ~w4857 & ~w7161;
assign w7163 = ~w7160 & w7162;
assign w7164 = ~w7155 & w7163;
assign w7165 = pi128 & w4060;
assign w7166 = ~w4095 & ~w4852;
assign w7167 = ~w7165 & w7166;
assign w7168 = (~pi065 & ~w7167) | (~pi065 & w18714) | (~w7167 & w18714);
assign w7169 = ~w4839 & ~w4885;
assign w7170 = ~w4001 & w7169;
assign w7171 = (~pi106 & ~w7170) | (~pi106 & w18715) | (~w7170 & w18715);
assign w7172 = ~pi031 & w3977;
assign w7173 = w3977 & w18716;
assign w7174 = ~w4855 & ~w4898;
assign w7175 = (w4015 & ~w7174) | (w4015 & w18717) | (~w7174 & w18717);
assign w7176 = ~w7168 & ~w7171;
assign w7177 = (~pi068 & ~w7176) | (~pi068 & w18718) | (~w7176 & w18718);
assign w7178 = w4044 & w3971;
assign w7179 = (pi128 & w4520) | (pi128 & w18719) | (w4520 & w18719);
assign w7180 = w3973 & w18356;
assign w7181 = w3992 & w4840;
assign w7182 = pi106 & ~w7181;
assign w7183 = ~w7180 & w7182;
assign w7184 = (~pi035 & w7179) | (~pi035 & w20799) | (w7179 & w20799);
assign w7185 = w7183 & ~w7184;
assign w7186 = pi031 & w4467;
assign w7187 = ~w4016 & ~w7186;
assign w7188 = w4873 & w7187;
assign w7189 = (~w7188 & w7900) | (~w7188 & w20800) | (w7900 & w20800);
assign w7190 = ~w3983 & ~w4456;
assign w7191 = ~pi106 & ~w7190;
assign w7192 = pi031 & w3989;
assign w7193 = w4021 & w7192;
assign w7194 = w3969 & w4059;
assign w7195 = pi031 & w3994;
assign w7196 = ~w7193 & ~w7195;
assign w7197 = ~w7191 & w7196;
assign w7198 = pi065 & ~pi068;
assign w7199 = (w7198 & ~w7197) | (w7198 & w18720) | (~w7197 & w18720);
assign w7200 = pi031 & w4031;
assign w7201 = w4031 & w3988;
assign w7202 = w3971 & w4010;
assign w7203 = ~w4020 & w18721;
assign w7204 = w4526 & ~w7203;
assign w7205 = w3981 & w3995;
assign w7206 = (~pi065 & w4452) | (~pi065 & w4529) | (w4452 & w4529);
assign w7207 = ~w4452 & ~w7205;
assign w7208 = w7169 & w7207;
assign w7209 = w7206 & ~w7208;
assign w7210 = ~w4082 & ~w7172;
assign w7211 = ~w4896 & ~w7202;
assign w7212 = w7210 & ~w7211;
assign w7213 = ~pi106 & w7212;
assign w7214 = ~w7209 & ~w7213;
assign w7215 = ~w7204 & w7214;
assign w7216 = ~w7199 & w7215;
assign w7217 = ~w7185 & w7189;
assign w7218 = w7216 & w18722;
assign w7219 = (pi068 & ~w7164) | (pi068 & w20801) | (~w7164 & w20801);
assign w7220 = w7218 & ~w7219;
assign w7221 = ~w4921 & w7220;
assign w7222 = w4921 & ~w7220;
assign w7223 = ~w7221 & ~w7222;
assign w7224 = ~w3517 & w4828;
assign w7225 = w3517 & ~w4828;
assign w7226 = ~w7224 & ~w7225;
assign w7227 = w7223 & w7226;
assign w7228 = ~w7223 & ~w7226;
assign w7229 = ~w7227 & ~w7228;
assign w7230 = (~pi529 & ~w7229) | (~pi529 & w18723) | (~w7229 & w18723);
assign w7231 = ~w7144 & ~w7229;
assign w7232 = w7230 & ~w7231;
assign w7233 = pi193 & pi475;
assign w7234 = pi529 & ~w7233;
assign w7235 = ~pi193 & ~pi475;
assign w7236 = w7234 & ~w7235;
assign w7237 = ~w7232 & ~w7236;
assign w7238 = ~w293 & ~w1047;
assign w7239 = (~w1396 & w7238) | (~w1396 & w18724) | (w7238 & w18724);
assign w7240 = ~pi123 & ~w7239;
assign w7241 = (pi123 & w320) | (pi123 & w18025) | (w320 & w18025);
assign w7242 = w286 & w317;
assign w7243 = ~w278 & ~w1120;
assign w7244 = ~w5028 & ~w7242;
assign w7245 = w7243 & w7244;
assign w7246 = ~w1114 & w7245;
assign w7247 = ~w7241 & w7246;
assign w7248 = ~w7240 & w7247;
assign w7249 = w264 & w304;
assign w7250 = ~w1240 & ~w7249;
assign w7251 = ~pi111 & ~w7250;
assign w7252 = w299 & w343;
assign w7253 = ~w378 & ~w7252;
assign w7254 = ~w7251 & w7253;
assign w7255 = ~pi048 & ~w7254;
assign w7256 = ~w1427 & ~w5045;
assign w7257 = ~w273 & w7256;
assign w7258 = (pi123 & ~w7257) | (pi123 & w18725) | (~w7257 & w18725);
assign w7259 = ~w1097 & ~w1115;
assign w7260 = (~pi123 & ~w7259) | (~pi123 & w7289) | (~w7259 & w7289);
assign w7261 = ~w1089 & ~w7260;
assign w7262 = ~w7255 & w18726;
assign w7263 = pi048 & ~w7248;
assign w7264 = ~pi123 & w324;
assign w7265 = ~w343 & w345;
assign w7266 = ~w7264 & ~w7265;
assign w7267 = (~pi048 & ~w1085) | (~pi048 & w18727) | (~w1085 & w18727);
assign w7268 = ~w361 & w7266;
assign w7269 = w7267 & w7268;
assign w7270 = w1224 & w18728;
assign w7271 = ~w7269 & ~w7270;
assign w7272 = (~pi123 & w1371) | (~pi123 & w18729) | (w1371 & w18729);
assign w7273 = pi023 & w1063;
assign w7274 = (w1420 & ~w1226) | (w1420 & w18730) | (~w1226 & w18730);
assign w7275 = ~w396 & ~w1082;
assign w7276 = w343 & ~w7275;
assign w7277 = ~pi123 & w364;
assign w7278 = ~w5020 & ~w7277;
assign w7279 = ~w7272 & ~w7274;
assign w7280 = ~w7276 & w7278;
assign w7281 = w7279 & w7280;
assign w7282 = (pi020 & w7271) | (pi020 & w18731) | (w7271 & w18731);
assign w7283 = (w386 & ~w5018) | (w386 & w18732) | (~w5018 & w18732);
assign w7284 = w383 & w1047;
assign w7285 = ~w1385 & ~w7284;
assign w7286 = ~w7283 & w7285;
assign w7287 = ~pi048 & ~w7286;
assign w7288 = ~w395 & ~w5382;
assign w7289 = ~pi123 & w312;
assign w7290 = w345 & w386;
assign w7291 = ~w7289 & ~w7290;
assign w7292 = ~w1263 & ~w5372;
assign w7293 = w274 & w1027;
assign w7294 = w7292 & ~w7293;
assign w7295 = (pi048 & ~w7291) | (pi048 & w18733) | (~w7291 & w18733);
assign w7296 = w7294 & ~w7295;
assign w7297 = (w5058 & w7288) | (w5058 & w18734) | (w7288 & w18734);
assign w7298 = w7296 & ~w7297;
assign w7299 = ~w7287 & w7298;
assign w7300 = ~w7282 & w7299;
assign w7301 = (~pi020 & w7263) | (~pi020 & w18735) | (w7263 & w18735);
assign w7302 = w7300 & ~w7301;
assign w7303 = ~w457 & ~w478;
assign w7304 = ~pi114 & ~w7303;
assign w7305 = ~w495 & ~w7304;
assign w7306 = w417 & w413;
assign w7307 = ~w1148 & ~w7306;
assign w7308 = ~w412 & ~w1145;
assign w7309 = w7307 & w7308;
assign w7310 = pi001 & ~w7309;
assign w7311 = pi001 & ~pi114;
assign w7312 = ~pi007 & w405;
assign w7313 = pi007 & w515;
assign w7314 = ~w469 & ~w7312;
assign w7315 = (w7311 & ~w7314) | (w7311 & w18736) | (~w7314 & w18736);
assign w7316 = ~w466 & w524;
assign w7317 = (~pi114 & w7316) | (~pi114 & w18737) | (w7316 & w18737);
assign w7318 = ~pi114 & w467;
assign w7319 = w486 & w941;
assign w7320 = ~w7318 & ~w7319;
assign w7321 = ~w1184 & ~w5133;
assign w7322 = w7320 & w7321;
assign w7323 = ~w7317 & w7322;
assign w7324 = ~w7310 & w7323;
assign w7325 = ~w7315 & w7324;
assign w7326 = w403 & w442;
assign w7327 = ~w972 & ~w5095;
assign w7328 = (~pi114 & ~w7327) | (~pi114 & w18739) | (~w7327 & w18739);
assign w7329 = (pi114 & w438) | (pi114 & w18740) | (w438 & w18740);
assign w7330 = w425 & w1170;
assign w7331 = ~w5101 & ~w7330;
assign w7332 = ~w1013 & ~w5074;
assign w7333 = ~w1008 & w7332;
assign w7334 = w7331 & w7333;
assign w7335 = ~w7328 & ~w7329;
assign w7336 = w7334 & w7335;
assign w7337 = ~pi114 & w426;
assign w7338 = ~w487 & ~w1013;
assign w7339 = ~w452 & ~w7338;
assign w7340 = (pi001 & w7339) | (pi001 & w18741) | (w7339 & w18741);
assign w7341 = (~pi114 & w416) | (~pi114 & w18742) | (w416 & w18742);
assign w7342 = ~w1186 & ~w7341;
assign w7343 = ~w7340 & w7342;
assign w7344 = pi001 & ~pi029;
assign w7345 = ~w7336 & w7344;
assign w7346 = w7343 & ~w7345;
assign w7347 = ~w488 & ~w969;
assign w7348 = (~w467 & w7347) | (~w467 & w18743) | (w7347 & w18743);
assign w7349 = ~pi114 & ~w7348;
assign w7350 = (w486 & ~w5094) | (w486 & w7319) | (~w5094 & w7319);
assign w7351 = w928 & w971;
assign w7352 = ~w498 & ~w7351;
assign w7353 = ~w7350 & w7352;
assign w7354 = ~w7349 & w7353;
assign w7355 = ~pi001 & ~w7354;
assign w7356 = w405 & w976;
assign w7357 = w409 & w5109;
assign w7358 = ~w7356 & ~w7357;
assign w7359 = ~pi013 & ~w991;
assign w7360 = w7358 & ~w7359;
assign w7361 = ~pi001 & ~w7360;
assign w7362 = w405 & w445;
assign w7363 = ~w945 & ~w7362;
assign w7364 = ~w921 & ~w7337;
assign w7365 = w7363 & w7364;
assign w7366 = pi098 & w425;
assign w7367 = ~w5099 & ~w7366;
assign w7368 = ~pi114 & w989;
assign w7369 = w5110 & w7313;
assign w7370 = ~w7368 & ~w7369;
assign w7371 = w536 & ~w7367;
assign w7372 = w7370 & ~w7371;
assign w7373 = w7365 & w7372;
assign w7374 = ~w7361 & w7373;
assign w7375 = ~pi029 & ~w7374;
assign w7376 = ~w7355 & ~w7375;
assign w7377 = w7346 & w7376;
assign w7378 = (pi029 & ~w7325) | (pi029 & w18744) | (~w7325 & w18744);
assign w7379 = w7377 & ~w7378;
assign w7380 = ~w7302 & w7379;
assign w7381 = w7302 & ~w7379;
assign w7382 = ~w7380 & ~w7381;
assign w7383 = ~pi108 & w7;
assign w7384 = ~w34 & ~w7383;
assign w7385 = pi107 & w187;
assign w7386 = w38 & w5230;
assign w7387 = w202 & w7385;
assign w7388 = ~w7386 & ~w7387;
assign w7389 = ~w150 & ~w5308;
assign w7390 = w7388 & w7389;
assign w7391 = (~pi040 & ~w7390) | (~pi040 & w18745) | (~w7390 & w18745);
assign w7392 = ~w58 & ~w191;
assign w7393 = ~w1290 & w7392;
assign w7394 = pi083 & ~w7393;
assign w7395 = w85 & ~w89;
assign w7396 = w5589 & ~w7395;
assign w7397 = ~w7394 & w7396;
assign w7398 = pi040 & ~w7397;
assign w7399 = ~w72 & ~w1352;
assign w7400 = ~pi083 & w7399;
assign w7401 = ~w51 & w5202;
assign w7402 = w213 & w7401;
assign w7403 = ~w7400 & ~w7402;
assign w7404 = ~w7398 & w18746;
assign w7405 = pi078 & ~w7404;
assign w7406 = ~w104 & ~w5582;
assign w7407 = w60 & ~w7406;
assign w7408 = ~w1352 & ~w5636;
assign w7409 = ~pi040 & w7408;
assign w7410 = ~w17 & ~w5179;
assign w7411 = ~w7407 & w7410;
assign w7412 = w7409 & w7411;
assign w7413 = ~w188 & ~w1302;
assign w7414 = w8 & ~w7413;
assign w7415 = (pi040 & ~w29) | (pi040 & w18747) | (~w29 & w18747);
assign w7416 = ~pi107 & w153;
assign w7417 = ~w7414 & w18748;
assign w7418 = w20 & w70;
assign w7419 = ~w190 & ~w7418;
assign w7420 = ~pi107 & w5174;
assign w7421 = w5208 & ~w7420;
assign w7422 = pi083 & ~w5610;
assign w7423 = ~w17 & w7422;
assign w7424 = w7419 & w7421;
assign w7425 = ~w7412 & ~w7417;
assign w7426 = ~w26 & w5615;
assign w7427 = ~w133 & ~w5304;
assign w7428 = ~w215 & w7427;
assign w7429 = ~w5613 & w7428;
assign w7430 = (~pi083 & w7426) | (~pi083 & w18035) | (w7426 & w18035);
assign w7431 = ~pi107 & w13;
assign w7432 = ~w7431 & w18749;
assign w7433 = w88 & ~w7432;
assign w7434 = ~w92 & ~w212;
assign w7435 = w36 & ~w7434;
assign w7436 = w107 & w18750;
assign w7437 = ~w203 & ~w5173;
assign w7438 = ~w7436 & w7437;
assign w7439 = ~w7435 & w7438;
assign w7440 = ~w7433 & w7439;
assign w7441 = (~pi040 & ~w7429) | (~pi040 & w18751) | (~w7429 & w18751);
assign w7442 = w7440 & ~w7441;
assign w7443 = (~pi078 & w7425) | (~pi078 & w18752) | (w7425 & w18752);
assign w7444 = w7442 & ~w7443;
assign w7445 = ~w7405 & w7444;
assign w7446 = ~w613 & ~w779;
assign w7447 = ~w1445 & w7446;
assign w7448 = pi104 & ~w7447;
assign w7449 = pi102 & ~w836;
assign w7450 = ~w1465 & w7449;
assign w7451 = w635 & ~w646;
assign w7452 = w7450 & ~w7451;
assign w7453 = pi127 & w683;
assign w7454 = w593 & w857;
assign w7455 = w689 & w7453;
assign w7456 = ~w7454 & ~w7455;
assign w7457 = ~w599 & ~w738;
assign w7458 = pi104 & ~w7457;
assign w7459 = w622 & w686;
assign w7460 = ~pi102 & ~w722;
assign w7461 = ~w7459 & w7460;
assign w7462 = ~w7458 & w7461;
assign w7463 = ~w7448 & w7452;
assign w7464 = w7456 & w7462;
assign w7465 = ~w7463 & ~w7464;
assign w7466 = ~pi104 & ~w1498;
assign w7467 = ~w653 & w7466;
assign w7468 = ~w608 & w871;
assign w7469 = w768 & w7468;
assign w7470 = ~w7467 & ~w7469;
assign w7471 = (pi012 & w7465) | (pi012 & w18753) | (w7465 & w18753);
assign w7472 = w572 & w585;
assign w7473 = w558 & w593;
assign w7474 = ~w568 & ~w675;
assign w7475 = ~w817 & ~w7473;
assign w7476 = w7474 & w7475;
assign w7477 = ~w1498 & ~w7472;
assign w7478 = ~pi102 & w7477;
assign w7479 = w7476 & w7478;
assign w7480 = ~w746 & ~w1459;
assign w7481 = w755 & ~w7480;
assign w7482 = w703 & w725;
assign w7483 = ~w581 & ~w7482;
assign w7484 = ~w7481 & w7483;
assign w7485 = pi102 & w7484;
assign w7486 = ~w589 & ~w814;
assign w7487 = w829 & ~w7486;
assign w7488 = w585 & w588;
assign w7489 = pi104 & ~w7488;
assign w7490 = ~w568 & w7489;
assign w7491 = ~w747 & w875;
assign w7492 = ~w7487 & w7491;
assign w7493 = ~w7479 & ~w7485;
assign w7494 = ~w585 & w718;
assign w7495 = (~pi104 & w7494) | (~pi104 & w18065) | (w7494 & w18065);
assign w7496 = w639 & w5501;
assign w7497 = ~w713 & ~w7496;
assign w7498 = w1518 & w7497;
assign w7499 = (~pi102 & ~w7498) | (~pi102 & w18754) | (~w7498 & w18754);
assign w7500 = w572 & w620;
assign w7501 = pi033 & w7500;
assign w7502 = ~w7501 & w18755;
assign w7503 = w645 & ~w7502;
assign w7504 = (pi104 & w799) | (pi104 & w18756) | (w799 & w18756);
assign w7505 = ~w759 & ~w813;
assign w7506 = ~w7504 & w7505;
assign w7507 = pi102 & w5518;
assign w7508 = w7506 & ~w7507;
assign w7509 = ~w7499 & w7508;
assign w7510 = ~w7503 & w7509;
assign w7511 = (~pi012 & w7493) | (~pi012 & w18757) | (w7493 & w18757);
assign w7512 = w7510 & ~w7511;
assign w7513 = ~w7471 & w7512;
assign w7514 = ~w7445 & w7513;
assign w7515 = w7445 & ~w7513;
assign w7516 = ~w7514 & ~w7515;
assign w7517 = ~w1049 & ~w5028;
assign w7518 = (pi123 & ~w1375) | (pi123 & w18758) | (~w1375 & w18758);
assign w7519 = ~w1022 & w1027;
assign w7520 = ~w1074 & ~w1223;
assign w7521 = ~w7519 & w7520;
assign w7522 = ~w7518 & w7521;
assign w7523 = pi048 & ~w7522;
assign w7524 = (~pi123 & ~w7259) | (~pi123 & w18759) | (~w7259 & w18759);
assign w7525 = pi093 & w286;
assign w7526 = ~w1259 & ~w7525;
assign w7527 = (~w312 & w7526) | (~w312 & w18760) | (w7526 & w18760);
assign w7528 = ~w7524 & w7527;
assign w7529 = ~pi048 & ~w7528;
assign w7530 = ~pi123 & ~w1422;
assign w7531 = w282 & w270;
assign w7532 = w7530 & ~w7531;
assign w7533 = w325 & ~w1089;
assign w7534 = w5043 & w7533;
assign w7535 = ~w7532 & ~w7534;
assign w7536 = ~w7529 & ~w7535;
assign w7537 = ~w7523 & w7536;
assign w7538 = pi020 & ~w7537;
assign w7539 = w258 & w1063;
assign w7540 = ~w1109 & ~w7539;
assign w7541 = (pi048 & ~w287) | (pi048 & w18761) | (~w287 & w18761);
assign w7542 = pi123 & ~w7540;
assign w7543 = w299 & w318;
assign w7544 = ~w7542 & w18762;
assign w7545 = ~w1276 & ~w1422;
assign w7546 = ~w365 & w7545;
assign w7547 = ~pi048 & w7546;
assign w7548 = (w314 & w1030) | (w314 & w18763) | (w1030 & w18763);
assign w7549 = ~w385 & ~w7548;
assign w7550 = w7547 & w7549;
assign w7551 = ~w7544 & ~w7550;
assign w7552 = w257 & w270;
assign w7553 = ~pi023 & w380;
assign w7554 = ~w7552 & ~w7553;
assign w7555 = pi123 & ~w259;
assign w7556 = ~w365 & w7555;
assign w7557 = w335 & ~w5026;
assign w7558 = w7554 & w7557;
assign w7559 = (~pi020 & w7551) | (~pi020 & w18764) | (w7551 & w18764);
assign w7560 = ~w253 & ~w1068;
assign w7561 = ~pi023 & ~w7560;
assign w7562 = (pi048 & w7561) | (pi048 & w18765) | (w7561 & w18765);
assign w7563 = (pi123 & w7562) | (pi123 & w18766) | (w7562 & w18766);
assign w7564 = ~w258 & w5000;
assign w7565 = ~w1273 & ~w5349;
assign w7566 = pi123 & ~w328;
assign w7567 = w7565 & ~w7566;
assign w7568 = (~pi123 & w7564) | (~pi123 & w18051) | (w7564 & w18051);
assign w7569 = w7567 & ~w7568;
assign w7570 = ~w333 & ~w5035;
assign w7571 = w283 & w18767;
assign w7572 = w7570 & w18768;
assign w7573 = (w7572 & w7569) | (w7572 & w18769) | (w7569 & w18769);
assign w7574 = ~w7563 & w7573;
assign w7575 = ~w7559 & w7574;
assign w7576 = ~w7538 & w7575;
assign w7577 = ~pi153 & w7576;
assign w7578 = pi153 & ~w7576;
assign w7579 = ~w7577 & ~w7578;
assign w7580 = w7516 & w7579;
assign w7581 = ~w7516 & ~w7579;
assign w7582 = ~w7580 & ~w7581;
assign w7583 = (~pi529 & w7582) | (~pi529 & w18770) | (w7582 & w18770);
assign w7584 = ~w7382 & w7582;
assign w7585 = w7583 & ~w7584;
assign w7586 = ~pi153 & pi515;
assign w7587 = pi529 & ~w7586;
assign w7588 = pi153 & ~pi515;
assign w7589 = w7587 & ~w7588;
assign w7590 = ~w7585 & ~w7589;
assign w7591 = ~w5243 & ~w7382;
assign w7592 = w5243 & w7382;
assign w7593 = ~w7591 & ~w7592;
assign w7594 = w560 & w585;
assign w7595 = ~w653 & ~w7594;
assign w7596 = (~pi104 & ~w7595) | (~pi104 & w18771) | (~w7595 & w18771);
assign w7597 = ~w595 & ~w654;
assign w7598 = pi104 & ~w7597;
assign w7599 = ~w708 & ~w750;
assign w7600 = ~w779 & w7599;
assign w7601 = ~w671 & ~w679;
assign w7602 = ~w7598 & w7601;
assign w7603 = w7602 & w18772;
assign w7604 = pi102 & ~w7603;
assign w7605 = w588 & w640;
assign w7606 = ~w752 & ~w7605;
assign w7607 = w566 & w1456;
assign w7608 = w597 & w648;
assign w7609 = ~w7607 & ~w7608;
assign w7610 = w7606 & w7609;
assign w7611 = ~pi102 & ~w7610;
assign w7612 = ~w750 & ~w770;
assign w7613 = ~w835 & w7612;
assign w7614 = (pi104 & ~w7613) | (pi104 & w18773) | (~w7613 & w18773);
assign w7615 = ~w608 & ~w1470;
assign w7616 = w7456 & w7615;
assign w7617 = ~w7611 & w18774;
assign w7618 = ~w7604 & w7617;
assign w7619 = ~pi012 & ~w7618;
assign w7620 = w626 & ~w755;
assign w7621 = w561 & w848;
assign w7622 = ~w7620 & ~w7621;
assign w7623 = (~pi102 & ~w766) | (~pi102 & w18775) | (~w766 & w18775);
assign w7624 = w7622 & w7623;
assign w7625 = pi104 & ~w858;
assign w7626 = w7624 & ~w7625;
assign w7627 = ~w731 & ~w1465;
assign w7628 = w7627 & w18776;
assign w7629 = ~w7626 & ~w7628;
assign w7630 = ~w847 & ~w1455;
assign w7631 = (~pi104 & w1462) | (~pi104 & w18777) | (w1462 & w18777);
assign w7632 = ~w583 & ~w798;
assign w7633 = ~w760 & ~w7632;
assign w7634 = ~w742 & ~w789;
assign w7635 = ~w7633 & w7634;
assign w7636 = pi102 & ~pi104;
assign w7637 = (w7636 & ~w7630) | (w7636 & w18778) | (~w7630 & w18778);
assign w7638 = w7635 & w20802;
assign w7639 = (pi012 & w7629) | (pi012 & w20803) | (w7629 & w20803);
assign w7640 = ~w607 & ~w5542;
assign w7641 = (~pi104 & w7640) | (~pi104 & w18779) | (w7640 & w18779);
assign w7642 = (w571 & ~w739) | (w571 & w18780) | (~w739 & w18780);
assign w7643 = w604 & w652;
assign w7644 = ~w712 & ~w7643;
assign w7645 = ~w7642 & w7644;
assign w7646 = ~w7641 & w7645;
assign w7647 = ~pi102 & ~w7646;
assign w7648 = (~w585 & w1470) | (~w585 & w18781) | (w1470 & w18781);
assign w7649 = (pi102 & w7648) | (pi102 & w18782) | (w7648 & w18782);
assign w7650 = (~pi104 & w884) | (~pi104 & w17985) | (w884 & w17985);
assign w7651 = w604 & w605;
assign w7652 = ~w7650 & ~w7651;
assign w7653 = ~w7649 & w7652;
assign w7654 = ~w7647 & w7653;
assign w7655 = ~w7639 & w7654;
assign w7656 = ~w7619 & w7655;
assign w7657 = w7655 & w18783;
assign w7658 = (pi179 & ~w7655) | (pi179 & w18784) | (~w7655 & w18784);
assign w7659 = ~w7657 & w20804;
assign w7660 = (w901 & w7657) | (w901 & w20805) | (w7657 & w20805);
assign w7661 = ~w7659 & ~w7660;
assign w7662 = (~pi529 & ~w7593) | (~pi529 & w18785) | (~w7593 & w18785);
assign w7663 = ~w7593 & ~w7661;
assign w7664 = w7662 & ~w7663;
assign w7665 = pi179 & pi457;
assign w7666 = pi529 & ~w7665;
assign w7667 = ~pi179 & ~pi457;
assign w7668 = w7666 & ~w7667;
assign w7669 = ~w7664 & ~w7668;
assign w7670 = w7218 & w20806;
assign w7671 = (pi358 & ~w7218) | (pi358 & w20807) | (~w7218 & w20807);
assign w7672 = ~w7670 & ~w7671;
assign w7673 = ~w4120 & w4276;
assign w7674 = w4120 & ~w4276;
assign w7675 = ~w7673 & ~w7674;
assign w7676 = w7672 & w7675;
assign w7677 = ~w7672 & ~w7675;
assign w7678 = ~w7676 & ~w7677;
assign w7679 = ~w3840 & ~w3855;
assign w7680 = ~pi091 & ~w7679;
assign w7681 = ~w3852 & ~w4371;
assign w7682 = pi024 & ~w4384;
assign w7683 = w7681 & w7682;
assign w7684 = ~pi024 & ~w3860;
assign w7685 = ~w3846 & w7684;
assign w7686 = ~pi005 & ~w3773;
assign w7687 = w3631 & ~w7686;
assign w7688 = ~w4788 & ~w7687;
assign w7689 = w7685 & w7688;
assign w7690 = ~w7680 & w7683;
assign w7691 = ~w7689 & ~w7690;
assign w7692 = ~pi091 & ~w3789;
assign w7693 = ~w4814 & w7692;
assign w7694 = ~w4363 & w7693;
assign w7695 = w3524 & w3550;
assign w7696 = ~w3632 & ~w7695;
assign w7697 = ~w3551 & ~w3774;
assign w7698 = (pi091 & ~w3543) | (pi091 & w18786) | (~w3543 & w18786);
assign w7699 = w7697 & w7698;
assign w7700 = w7696 & w7699;
assign w7701 = ~w7694 & ~w7700;
assign w7702 = ~pi091 & w3531;
assign w7703 = (~pi005 & w7702) | (~pi005 & w18283) | (w7702 & w18283);
assign w7704 = ~pi084 & w3520;
assign w7705 = ~w4787 & ~w7704;
assign w7706 = pi091 & ~w7705;
assign w7707 = (pi005 & ~w3518) | (pi005 & w18787) | (~w3518 & w18787);
assign w7708 = ~w7705 & w18788;
assign w7709 = ~w7703 & ~w7708;
assign w7710 = ~pi018 & w7709;
assign w7711 = w3539 & w3801;
assign w7712 = w3568 & w3645;
assign w7713 = ~w3598 & ~w7712;
assign w7714 = ~w7695 & ~w7711;
assign w7715 = ~pi024 & w7714;
assign w7716 = w7713 & w7715;
assign w7717 = w3547 & w3596;
assign w7718 = ~w7717 & w18789;
assign w7719 = ~w7716 & ~w7718;
assign w7720 = pi084 & w3550;
assign w7721 = ~w3530 & w3533;
assign w7722 = ~w7720 & w7721;
assign w7723 = (~w3830 & ~w7722) | (~w3830 & w18790) | (~w7722 & w18790);
assign w7724 = pi024 & ~w7723;
assign w7725 = ~w7719 & ~w7724;
assign w7726 = w7710 & w7725;
assign w7727 = pi018 & ~w7701;
assign w7728 = ~w7691 & w7727;
assign w7729 = ~w7726 & ~w7728;
assign w7730 = ~w3524 & w3545;
assign w7731 = ~w3816 & ~w4814;
assign w7732 = (~pi091 & ~w7731) | (~pi091 & w18791) | (~w7731 & w18791);
assign w7733 = ~w4775 & ~w4807;
assign w7734 = w3801 & w4378;
assign w7735 = (pi024 & ~w3531) | (pi024 & w18792) | (~w3531 & w18792);
assign w7736 = w7733 & w18793;
assign w7737 = ~w7732 & w7736;
assign w7738 = ~w3551 & ~w3624;
assign w7739 = ~w4387 & w7738;
assign w7740 = w3518 & w4780;
assign w7741 = ~w4400 & ~w7740;
assign w7742 = w7739 & w7741;
assign w7743 = pi091 & ~w7742;
assign w7744 = w3565 & ~w3609;
assign w7745 = ~pi005 & w7744;
assign w7746 = ~w4411 & ~w7745;
assign w7747 = ~w3602 & ~w4401;
assign w7748 = ~pi024 & w7747;
assign w7749 = ~pi091 & ~w7746;
assign w7750 = w7748 & ~w7749;
assign w7751 = ~w7743 & w7750;
assign w7752 = ~pi091 & w3630;
assign w7753 = (pi005 & w7752) | (pi005 & w18794) | (w7752 & w18794);
assign w7754 = (~w7753 & w7751) | (~w7753 & w20808) | (w7751 & w20808);
assign w7755 = ~w7729 & w7754;
assign w7756 = ~w3517 & w7755;
assign w7757 = w3517 & ~w7755;
assign w7758 = ~w7756 & ~w7757;
assign w7759 = w4543 & w7758;
assign w7760 = ~w4543 & ~w7758;
assign w7761 = ~w7759 & ~w7760;
assign w7762 = w7678 & w7761;
assign w7763 = ~pi529 & ~w7762;
assign w7764 = ~w7678 & ~w7761;
assign w7765 = w7763 & ~w7764;
assign w7766 = ~pi358 & pi481;
assign w7767 = pi529 & ~w7766;
assign w7768 = pi358 & ~pi481;
assign w7769 = w7767 & ~w7768;
assign w7770 = ~w7765 & ~w7769;
assign w7771 = ~w4828 & w4985;
assign w7772 = w4828 & ~w4985;
assign w7773 = ~w7771 & ~w7772;
assign w7774 = w3663 & ~w7773;
assign w7775 = ~w3663 & w7773;
assign w7776 = ~w7774 & ~w7775;
assign w7777 = ~pi043 & w3481;
assign w7778 = (~pi122 & w7777) | (~pi122 & w18795) | (w7777 & w18795);
assign w7779 = ~w3668 & ~w4944;
assign w7780 = pi122 & ~w7779;
assign w7781 = ~w3762 & ~w3953;
assign w7782 = ~w7780 & w7781;
assign w7783 = ~pi070 & ~w3377;
assign w7784 = ~w4313 & w7783;
assign w7785 = pi076 & w3491;
assign w7786 = ~w3450 & ~w7785;
assign w7787 = pi122 & ~w7786;
assign w7788 = ~w3480 & ~w3925;
assign w7789 = ~w3505 & w7788;
assign w7790 = ~w7787 & w7789;
assign w7791 = (~pi122 & w7784) | (~pi122 & w18796) | (w7784 & w18796);
assign w7792 = ~w3691 & ~w3953;
assign w7793 = ~pi122 & ~w7792;
assign w7794 = (w3721 & w3458) | (w3721 & w18797) | (w3458 & w18797);
assign w7795 = ~w4968 & ~w7794;
assign w7796 = ~w7793 & w18798;
assign w7797 = (pi039 & ~w7790) | (pi039 & w20809) | (~w7790 & w20809);
assign w7798 = w7796 & ~w7797;
assign w7799 = (~pi039 & ~w7782) | (~pi039 & w18799) | (~w7782 & w18799);
assign w7800 = ~w3371 & ~w3395;
assign w7801 = ~pi070 & ~w7800;
assign w7802 = (pi122 & w7801) | (pi122 & w18800) | (w7801 & w18800);
assign w7803 = w4299 & ~w7802;
assign w7804 = w3384 & w3412;
assign w7805 = ~w3475 & ~w7804;
assign w7806 = ~pi043 & w3714;
assign w7807 = w7805 & ~w7806;
assign w7808 = ~w3404 & w3697;
assign w7809 = ~w3445 & ~w3674;
assign w7810 = w3913 & ~w7809;
assign w7811 = ~w3440 & ~w3445;
assign w7812 = ~w3475 & ~w4944;
assign w7813 = w7811 & w7812;
assign w7814 = ~pi122 & ~w7813;
assign w7815 = ~w7810 & ~w7814;
assign w7816 = (~pi039 & ~w7807) | (~pi039 & w18801) | (~w7807 & w18801);
assign w7817 = w7815 & ~w7816;
assign w7818 = (pi017 & ~w7817) | (pi017 & w18802) | (~w7817 & w18802);
assign w7819 = ~w3432 & ~w4931;
assign w7820 = ~w3753 & w7819;
assign w7821 = ~pi122 & ~w7820;
assign w7822 = ~w3948 & ~w4932;
assign w7823 = (~pi039 & w7821) | (~pi039 & w18803) | (w7821 & w18803);
assign w7824 = pi039 & ~pi122;
assign w7825 = w3377 & w3384;
assign w7826 = w3708 & w4340;
assign w7827 = w3382 & w3386;
assign w7828 = ~w7826 & ~w7827;
assign w7829 = ~w3505 & ~w3943;
assign w7830 = w7828 & w7829;
assign w7831 = (w3692 & w3481) | (w3692 & w18804) | (w3481 & w18804);
assign w7832 = ~w3438 & ~w7831;
assign w7833 = w3756 & ~w7832;
assign w7834 = ~w3411 & ~w3684;
assign w7835 = ~w3730 & w7834;
assign w7836 = w3459 & ~w7835;
assign w7837 = ~w3750 & ~w7826;
assign w7838 = w3464 & ~w7837;
assign w7839 = ~w7836 & ~w7838;
assign w7840 = ~w7833 & w7839;
assign w7841 = (w7824 & ~w7830) | (w7824 & w18805) | (~w7830 & w18805);
assign w7842 = w7840 & w18806;
assign w7843 = ~w7818 & w7842;
assign w7844 = (~pi017 & ~w7798) | (~pi017 & w18807) | (~w7798 & w18807);
assign w7845 = w7843 & ~w7844;
assign w7846 = w3989 & w7156;
assign w7847 = (~pi106 & w7846) | (~pi106 & w18808) | (w7846 & w18808);
assign w7848 = ~w4073 & ~w4864;
assign w7849 = pi106 & ~w7848;
assign w7850 = ~w3997 & ~w4531;
assign w7851 = ~w7849 & w7850;
assign w7852 = w3989 & w3982;
assign w7853 = ~pi035 & w4037;
assign w7854 = ~w7172 & ~w7853;
assign w7855 = (~pi106 & ~w7854) | (~pi106 & w18809) | (~w7854 & w18809);
assign w7856 = pi031 & w4059;
assign w7857 = ~w4885 & ~w7856;
assign w7858 = pi106 & ~w7857;
assign w7859 = w3974 & ~w4018;
assign w7860 = ~w7202 & ~w7859;
assign w7861 = ~w7858 & w7860;
assign w7862 = ~w3997 & ~w4469;
assign w7863 = ~pi106 & ~w7862;
assign w7864 = pi106 & w4067;
assign w7865 = ~w4462 & ~w7864;
assign w7866 = ~w4055 & ~w4487;
assign w7867 = ~w7865 & w7866;
assign w7868 = ~w4899 & ~w7867;
assign w7869 = ~w7863 & w7868;
assign w7870 = (pi065 & ~w7861) | (pi065 & w18810) | (~w7861 & w18810);
assign w7871 = w7869 & ~w7870;
assign w7872 = (~pi065 & ~w7851) | (~pi065 & w18811) | (~w7851 & w18811);
assign w7873 = ~w4490 & ~w7181;
assign w7874 = ~w4019 & ~w4850;
assign w7875 = (pi106 & ~w7874) | (pi106 & w18812) | (~w7874 & w18812);
assign w7876 = w7873 & ~w7875;
assign w7877 = w3982 & w4486;
assign w7878 = ~w4872 & ~w7877;
assign w7879 = ~pi035 & w4519;
assign w7880 = w7878 & ~w7879;
assign w7881 = ~w3994 & ~w4898;
assign w7882 = w4061 & ~w7881;
assign w7883 = ~w4864 & ~w4872;
assign w7884 = ~w4898 & ~w7194;
assign w7885 = w7883 & w7884;
assign w7886 = ~pi106 & ~w7885;
assign w7887 = ~w7882 & ~w7886;
assign w7888 = (~pi065 & ~w7880) | (~pi065 & w18813) | (~w7880 & w18813);
assign w7889 = w7887 & ~w7888;
assign w7890 = (pi068 & ~w7889) | (pi068 & w18814) | (~w7889 & w18814);
assign w7891 = ~w4456 & ~w4852;
assign w7892 = ~w4042 & w7891;
assign w7893 = ~pi106 & ~w7892;
assign w7894 = ~w3984 & ~w4848;
assign w7895 = (~pi065 & w7893) | (~pi065 & w18815) | (w7893 & w18815);
assign w7896 = pi065 & ~pi106;
assign w7897 = ~w3978 & ~w4067;
assign w7898 = ~w7173 & w7211;
assign w7899 = (w7896 & ~w7898) | (w7896 & w18816) | (~w7898 & w18816);
assign w7900 = pi065 & pi106;
assign w7901 = ~w7181 & ~w7200;
assign w7902 = pi035 & ~w7901;
assign w7903 = (w7900 & w7902) | (w7900 & w18817) | (w7902 & w18817);
assign w7904 = ~w4462 & ~w4837;
assign w7905 = ~w4504 & w7904;
assign w7906 = w4526 & ~w7905;
assign w7907 = ~w4038 & ~w7173;
assign w7908 = w4015 & ~w7907;
assign w7909 = ~w7899 & ~w7903;
assign w7910 = ~w7906 & ~w7908;
assign w7911 = w7909 & w7910;
assign w7912 = ~w7895 & w7911;
assign w7913 = ~w7890 & w7912;
assign w7914 = (~pi068 & ~w7871) | (~pi068 & w18818) | (~w7871 & w18818);
assign w7915 = w7913 & ~w7914;
assign w7916 = ~w7845 & w7915;
assign w7917 = w7845 & ~w7915;
assign w7918 = ~w7916 & ~w7917;
assign w7919 = ~pi009 & w4126;
assign w7920 = w4137 & w4159;
assign w7921 = ~w7919 & ~w7920;
assign w7922 = pi124 & w4197;
assign w7923 = ~w4226 & ~w7922;
assign w7924 = pi113 & w7923;
assign w7925 = (~pi113 & ~w4263) | (~pi113 & w18819) | (~w4263 & w18819);
assign w7926 = w7921 & w7925;
assign w7927 = ~w7924 & ~w7926;
assign w7928 = ~w4124 & w4213;
assign w7929 = ~pi125 & w4159;
assign w7930 = w4253 & w7929;
assign w7931 = ~w4627 & ~w7930;
assign w7932 = ~w4189 & ~w4631;
assign w7933 = w4231 & ~w7932;
assign w7934 = ~w7061 & ~w7071;
assign w7935 = ~w7933 & w7934;
assign w7936 = (~pi113 & w7930) | (~pi113 & w18821) | (w7930 & w18821);
assign w7937 = (w4188 & w4252) | (w4188 & w18822) | (w4252 & w18822);
assign w7938 = ~pi124 & w4158;
assign w7939 = ~w6969 & ~w7938;
assign w7940 = pi113 & ~w7939;
assign w7941 = ~w4561 & ~w7015;
assign w7942 = ~w7937 & ~w7940;
assign w7943 = w7941 & w7942;
assign w7944 = (~pi096 & ~w7935) | (~pi096 & w18823) | (~w7935 & w18823);
assign w7945 = w7943 & ~w7944;
assign w7946 = (pi010 & ~w7945) | (pi010 & w18824) | (~w7945 & w18824);
assign w7947 = ~w4231 & ~w4621;
assign w7948 = ~w4693 & w7947;
assign w7949 = (~w4729 & w7948) | (~w4729 & w18825) | (w7948 & w18825);
assign w7950 = pi096 & ~w7949;
assign w7951 = w4137 & w4183;
assign w7952 = ~w4242 & ~w7951;
assign w7953 = w4258 & w4662;
assign w7954 = w7952 & ~w7953;
assign w7955 = ~w4242 & ~w4692;
assign w7956 = ~w4701 & ~w6992;
assign w7957 = w7955 & w7956;
assign w7958 = ~w4125 & w4254;
assign w7959 = ~pi009 & w4701;
assign w7960 = ~w7958 & ~w7959;
assign w7961 = ~pi113 & ~w7957;
assign w7962 = w7960 & ~w7961;
assign w7963 = (~pi096 & ~w7954) | (~pi096 & w18826) | (~w7954 & w18826);
assign w7964 = w7962 & ~w7963;
assign w7965 = (~pi010 & ~w7964) | (~pi010 & w18827) | (~w7964 & w18827);
assign w7966 = ~w4559 & ~w6985;
assign w7967 = ~w4179 & w7966;
assign w7968 = ~pi113 & ~w7967;
assign w7969 = ~w4257 & ~w6984;
assign w7970 = (~pi096 & w7968) | (~pi096 & w18828) | (w7968 & w18828);
assign w7971 = ~w4146 & ~w4729;
assign w7972 = pi009 & ~w7971;
assign w7973 = ~pi009 & w4163;
assign w7974 = (w4726 & w7972) | (w4726 & w18829) | (w7972 & w18829);
assign w7975 = w4207 & ~w4237;
assign w7976 = ~w4145 & ~w4545;
assign w7977 = ~w7975 & ~w7976;
assign w7978 = w4138 & w4189;
assign w7979 = (w4738 & w7977) | (w4738 & w18830) | (w7977 & w18830);
assign w7980 = w4253 & w4263;
assign w7981 = ~w4561 & ~w7980;
assign w7982 = ~w4607 & w7981;
assign w7983 = w4632 & ~w7982;
assign w7984 = w4263 & w6979;
assign w7985 = ~w4257 & ~w7984;
assign w7986 = pi113 & ~w7985;
assign w7987 = ~w7974 & ~w7979;
assign w7988 = ~w7983 & ~w7986;
assign w7989 = w7987 & w7988;
assign w7990 = ~w7970 & w7989;
assign w7991 = ~w7965 & w7990;
assign w7992 = ~w7946 & w7991;
assign w7993 = w7991 & w18831;
assign w7994 = (pi302 & ~w7991) | (pi302 & w18832) | (~w7991 & w18832);
assign w7995 = ~w7993 & ~w7994;
assign w7996 = w7918 & w7995;
assign w7997 = ~w7918 & ~w7995;
assign w7998 = ~w7996 & ~w7997;
assign w7999 = ~w7776 & ~w7998;
assign w8000 = ~pi529 & ~w7999;
assign w8001 = w7776 & w7998;
assign w8002 = w8000 & ~w8001;
assign w8003 = pi302 & pi502;
assign w8004 = pi529 & ~w8003;
assign w8005 = ~pi302 & ~pi502;
assign w8006 = w8004 & ~w8005;
assign w8007 = ~w8002 & ~w8006;
assign w8008 = ~w551 & ~w7382;
assign w8009 = w551 & w7382;
assign w8010 = ~w8008 & ~w8009;
assign w8011 = w2 & w26;
assign w8012 = ~w72 & ~w178;
assign w8013 = (~pi083 & ~w8012) | (~pi083 & w18833) | (~w8012 & w18833);
assign w8014 = (pi083 & w5199) | (pi083 & w18834) | (w5199 & w18834);
assign w8015 = ~w16 & ~w125;
assign w8016 = ~w191 & ~w195;
assign w8017 = w8015 & w8016;
assign w8018 = ~w8013 & ~w8014;
assign w8019 = ~w134 & w8017;
assign w8020 = w8018 & w8019;
assign w8021 = pi014 & ~w7413;
assign w8022 = ~w5279 & ~w5631;
assign w8023 = ~w8021 & w8022;
assign w8024 = pi083 & ~w8023;
assign w8025 = w8 & w135;
assign w8026 = w46 & w1299;
assign w8027 = ~w8025 & ~w8026;
assign w8028 = ~w105 & ~w194;
assign w8029 = w8027 & w8028;
assign w8030 = ~pi040 & ~w8029;
assign w8031 = ~pi083 & w150;
assign w8032 = ~pi078 & ~w51;
assign w8033 = ~w8031 & w8032;
assign w8034 = w7388 & w8033;
assign w8035 = ~w8024 & ~w8030;
assign w8036 = w8034 & w8035;
assign w8037 = pi040 & ~w8020;
assign w8038 = w8036 & ~w8037;
assign w8039 = ~w29 & ~w160;
assign w8040 = ~w106 & ~w211;
assign w8041 = ~w5232 & w8040;
assign w8042 = ~w172 & ~w231;
assign w8043 = ~w1341 & ~w5583;
assign w8044 = w8042 & w8043;
assign w8045 = ~w182 & ~w5278;
assign w8046 = pi078 & w8045;
assign w8047 = ~w7413 & w18835;
assign w8048 = w8046 & ~w8047;
assign w8049 = ~w41 & ~w1299;
assign w8050 = (w1348 & ~w8049) | (w1348 & w18836) | (~w8049 & w18836);
assign w8051 = (~pi083 & w1305) | (~pi083 & w18837) | (w1305 & w18837);
assign w8052 = ~w8050 & ~w8051;
assign w8053 = w8048 & w8052;
assign w8054 = pi040 & ~w8044;
assign w8055 = (~pi040 & ~w8041) | (~pi040 & w18838) | (~w8041 & w18838);
assign w8056 = w8053 & w20810;
assign w8057 = (w9 & w180) | (w9 & w18839) | (w180 & w18839);
assign w8058 = ~w166 & ~w1311;
assign w8059 = ~w8057 & w8058;
assign w8060 = ~pi040 & ~w8059;
assign w8061 = w23 & w60;
assign w8062 = ~w30 & w18840;
assign w8063 = w234 & ~w8062;
assign w8064 = ~w1358 & ~w8031;
assign w8065 = pi040 & ~w8064;
assign w8066 = ~pi083 & w16;
assign w8067 = ~w1312 & ~w8066;
assign w8068 = w189 & w18841;
assign w8069 = ~w5271 & ~w8068;
assign w8070 = ~w8065 & w8067;
assign w8071 = w8070 & w18842;
assign w8072 = ~w8060 & w8071;
assign w8073 = ~w8038 & ~w8056;
assign w8074 = (w8072 & w8038) | (w8072 & w20811) | (w8038 & w20811);
assign w8075 = (w18843 & w8038) | (w18843 & w20812) | (w8038 & w20812);
assign w8076 = (~w8038 & w20813) | (~w8038 & w20814) | (w20813 & w20814);
assign w8077 = ~w8075 & ~w8076;
assign w8078 = ~w901 & w8077;
assign w8079 = w901 & ~w8077;
assign w8080 = ~w8078 & ~w8079;
assign w8081 = (~pi529 & ~w8010) | (~pi529 & w18845) | (~w8010 & w18845);
assign w8082 = ~w8010 & ~w8080;
assign w8083 = w8081 & ~w8082;
assign w8084 = pi142 & pi400;
assign w8085 = pi529 & ~w8084;
assign w8086 = ~pi142 & ~pi400;
assign w8087 = w8085 & ~w8086;
assign w8088 = ~w8083 & ~w8087;
assign w8089 = w519 & w969;
assign w8090 = ~w1152 & ~w8089;
assign w8091 = (~w5109 & w8089) | (~w5109 & w18846) | (w8089 & w18846);
assign w8092 = (~pi001 & w8091) | (~pi001 & w18847) | (w8091 & w18847);
assign w8093 = ~w936 & ~w7366;
assign w8094 = w5136 & ~w8093;
assign w8095 = (w5109 & w409) | (w5109 & w18848) | (w409 & w18848);
assign w8096 = ~w8094 & ~w8095;
assign w8097 = (pi001 & w7316) | (pi001 & w18849) | (w7316 & w18849);
assign w8098 = ~w539 & ~w5465;
assign w8099 = (w7311 & ~w8098) | (w7311 & w18850) | (~w8098 & w18850);
assign w8100 = ~w521 & ~w1148;
assign w8101 = ~pi114 & ~w8100;
assign w8102 = ~w449 & ~w1154;
assign w8103 = w1011 & ~w8102;
assign w8104 = ~w8097 & ~w8099;
assign w8105 = ~w8101 & ~w8103;
assign w8106 = w8105 & w18851;
assign w8107 = (~pi029 & ~w8106) | (~pi029 & w18852) | (~w8106 & w18852);
assign w8108 = ~w466 & ~w1170;
assign w8109 = pi021 & ~w8108;
assign w8110 = (w5136 & w8109) | (w5136 & w18853) | (w8109 & w18853);
assign w8111 = ~w942 & ~w5074;
assign w8112 = w437 & ~w8111;
assign w8113 = (pi001 & w5102) | (pi001 & w18854) | (w5102 & w18854);
assign w8114 = ~w8112 & ~w8113;
assign w8115 = w415 & w432;
assign w8116 = ~w516 & ~w8115;
assign w8117 = ~w418 & w5095;
assign w8118 = w8116 & ~w8117;
assign w8119 = ~w516 & ~w922;
assign w8120 = w8119 & w18855;
assign w8121 = ~pi114 & ~w8120;
assign w8122 = (~pi001 & ~w8118) | (~pi001 & w18856) | (~w8118 & w18856);
assign w8123 = ~w8121 & ~w8122;
assign w8124 = ~w8110 & w8114;
assign w8125 = w8123 & w8124;
assign w8126 = pi029 & ~w8125;
assign w8127 = ~w412 & w18857;
assign w8128 = ~pi114 & ~w8127;
assign w8129 = w5081 & w7367;
assign w8130 = w445 & w475;
assign w8131 = ~w7362 & ~w8130;
assign w8132 = (w7311 & w8129) | (w7311 & w18858) | (w8129 & w18858);
assign w8133 = (w446 & w989) | (w446 & w18859) | (w989 & w18859);
assign w8134 = ~w468 & ~w8133;
assign w8135 = w5136 & ~w8134;
assign w8136 = ~w507 & ~w1142;
assign w8137 = pi001 & w5110;
assign w8138 = w409 & w8137;
assign w8139 = ~w946 & ~w8138;
assign w8140 = w507 & w928;
assign w8141 = w8139 & ~w8140;
assign w8142 = ~pi001 & w5109;
assign w8143 = (w8142 & ~w8136) | (w8142 & w18860) | (~w8136 & w18860);
assign w8144 = w8141 & ~w8143;
assign w8145 = ~w8132 & ~w8135;
assign w8146 = w8144 & w8145;
assign w8147 = (~pi001 & w8128) | (~pi001 & w18861) | (w8128 & w18861);
assign w8148 = w8146 & ~w8147;
assign w8149 = ~w8126 & w8148;
assign w8150 = ~w8107 & w8149;
assign w8151 = ~w1128 & w8150;
assign w8152 = w1128 & ~w8150;
assign w8153 = ~w8151 & ~w8152;
assign w8154 = w5651 & w8153;
assign w8155 = ~w5651 & ~w8153;
assign w8156 = ~w8154 & ~w8155;
assign w8157 = w1525 & w18862;
assign w8158 = (pi173 & ~w1525) | (pi173 & w18863) | (~w1525 & w18863);
assign w8159 = ~w8157 & ~w8158;
assign w8160 = ~w145 & w1367;
assign w8161 = w145 & ~w1367;
assign w8162 = ~w8160 & ~w8161;
assign w8163 = w8159 & w8162;
assign w8164 = ~w8159 & ~w8162;
assign w8165 = ~w8163 & ~w8164;
assign w8166 = (~pi529 & ~w8165) | (~pi529 & w18864) | (~w8165 & w18864);
assign w8167 = w8156 & ~w8165;
assign w8168 = w8166 & ~w8167;
assign w8169 = pi173 & pi407;
assign w8170 = pi529 & ~w8169;
assign w8171 = ~pi173 & ~pi407;
assign w8172 = w8170 & ~w8171;
assign w8173 = ~w8168 & ~w8172;
assign w8174 = ~w3972 & ~w4074;
assign w8175 = pi106 & ~w8174;
assign w8176 = ~pi106 & w4834;
assign w8177 = ~w8176 & w18865;
assign w8178 = ~w4048 & ~w4447;
assign w8179 = ~w4839 & w8178;
assign w8180 = w8177 & w8179;
assign w8181 = ~w7865 & ~w8175;
assign w8182 = w8180 & ~w8181;
assign w8183 = ~w4487 & ~w4520;
assign w8184 = ~pi106 & ~w8183;
assign w8185 = w3971 & w4047;
assign w8186 = ~w4897 & ~w8185;
assign w8187 = ~w8184 & w8186;
assign w8188 = pi065 & ~w8187;
assign w8189 = (~pi035 & ~w18866) | (~pi035 & w20799) | (~w18866 & w20799);
assign w8190 = ~w3996 & ~w4530;
assign w8191 = (w4015 & ~w8190) | (w4015 & w4899) | (~w8190 & w4899);
assign w8192 = ~w8188 & w18867;
assign w8193 = ~pi065 & ~w8182;
assign w8194 = w8192 & ~w8193;
assign w8195 = ~w4019 & ~w4485;
assign w8196 = (~w7194 & w8174) | (~w7194 & w20815) | (w8174 & w20815);
assign w8197 = (pi065 & ~w8196) | (pi065 & w18869) | (~w8196 & w18869);
assign w8198 = (~w4056 & ~w4020) | (~w4056 & w18870) | (~w4020 & w18870);
assign w8199 = w4053 & w4486;
assign w8200 = ~w4452 & ~w8199;
assign w8201 = w4097 & w4498;
assign w8202 = ~pi065 & ~w8200;
assign w8203 = ~w8201 & ~w8202;
assign w8204 = w8198 & w8203;
assign w8205 = (~pi068 & ~w8204) | (~pi068 & w20816) | (~w8204 & w20816);
assign w8206 = w3982 & w4037;
assign w8207 = ~w4001 & ~w7178;
assign w8208 = ~w3997 & w4908;
assign w8209 = pi106 & ~w8208;
assign w8210 = w3969 & w4018;
assign w8211 = w4016 & w4098;
assign w8212 = ~w4851 & ~w8210;
assign w8213 = ~w8211 & w8212;
assign w8214 = ~w8209 & w8213;
assign w8215 = (~pi065 & ~w8214) | (~pi065 & w18871) | (~w8214 & w18871);
assign w8216 = w3988 & w4037;
assign w8217 = ~w3994 & ~w8216;
assign w8218 = (pi065 & w3994) | (pi065 & w7896) | (w3994 & w7896);
assign w8219 = (w8218 & ~w7873) | (w8218 & w18872) | (~w7873 & w18872);
assign w8220 = ~w4834 & ~w7156;
assign w8221 = w3973 & w4841;
assign w8222 = w8220 & ~w8221;
assign w8223 = w7900 & ~w8222;
assign w8224 = w4003 & w8185;
assign w8225 = ~w7151 & ~w8224;
assign w8226 = ~w4524 & w8225;
assign w8227 = ~w8223 & w8226;
assign w8228 = ~w8219 & w8227;
assign w8229 = ~w8215 & w8228;
assign w8230 = ~w8205 & w8229;
assign w8231 = pi068 & ~w8194;
assign w8232 = w8230 & ~w8231;
assign w8233 = ~w4357 & w8232;
assign w8234 = w4357 & ~w8232;
assign w8235 = ~w8233 & ~w8234;
assign w8236 = ~w3517 & w3873;
assign w8237 = w3517 & ~w3873;
assign w8238 = ~w8236 & ~w8237;
assign w8239 = w8235 & w8238;
assign w8240 = ~w8235 & ~w8238;
assign w8241 = ~w8239 & ~w8240;
assign w8242 = ~w4540 & w7220;
assign w8243 = w4540 & ~w7220;
assign w8244 = ~w8242 & ~w8243;
assign w8245 = w4639 & w20817;
assign w8246 = (pi132 & ~w4639) | (pi132 & w20818) | (~w4639 & w20818);
assign w8247 = ~w8245 & ~w8246;
assign w8248 = w8244 & w8247;
assign w8249 = ~w8244 & ~w8247;
assign w8250 = ~w8248 & ~w8249;
assign w8251 = w8241 & w8250;
assign w8252 = ~pi529 & ~w8251;
assign w8253 = ~w8241 & ~w8250;
assign w8254 = w8252 & ~w8253;
assign w8255 = ~pi132 & pi447;
assign w8256 = pi529 & ~w8255;
assign w8257 = pi132 & ~pi447;
assign w8258 = w8256 & ~w8257;
assign w8259 = ~w8254 & ~w8258;
assign w8260 = ~w4641 & w4749;
assign w8261 = w4641 & ~w4749;
assign w8262 = ~w8260 & ~w8261;
assign w8263 = ~pi175 & w7123;
assign w8264 = pi175 & ~w7123;
assign w8265 = ~w8263 & ~w8264;
assign w8266 = w8262 & w8265;
assign w8267 = ~w8262 & ~w8265;
assign w8268 = ~w8266 & ~w8267;
assign w8269 = ~w7220 & w8232;
assign w8270 = w7220 & ~w8232;
assign w8271 = ~w8269 & ~w8270;
assign w8272 = w3876 & w8271;
assign w8273 = ~w3876 & ~w8271;
assign w8274 = ~w8272 & ~w8273;
assign w8275 = w8268 & w8274;
assign w8276 = ~pi529 & ~w8275;
assign w8277 = ~w8268 & ~w8274;
assign w8278 = w8276 & ~w8277;
assign w8279 = ~pi175 & pi416;
assign w8280 = pi529 & ~w8279;
assign w8281 = pi175 & ~pi416;
assign w8282 = w8280 & ~w8281;
assign w8283 = ~w8278 & ~w8282;
assign w8284 = ~w567 & ~w654;
assign w8285 = (pi104 & ~w8284) | (pi104 & w18756) | (~w8284 & w18756);
assign w8286 = ~w586 & ~w5540;
assign w8287 = ~w7500 & w8286;
assign w8288 = w1456 & w18873;
assign w8289 = w8287 & ~w8288;
assign w8290 = (~pi102 & ~w8289) | (~pi102 & w18874) | (~w8289 & w18874);
assign w8291 = ~w836 & ~w5536;
assign w8292 = (pi104 & ~w7627) | (pi104 & w18875) | (~w7627 & w18875);
assign w8293 = (~pi104 & w725) | (~pi104 & w18876) | (w725 & w18876);
assign w8294 = (pi102 & w8293) | (pi102 & w18877) | (w8293 & w18877);
assign w8295 = w829 & w863;
assign w8296 = ~w606 & ~w1453;
assign w8297 = ~w8295 & w8296;
assign w8298 = ~pi104 & ~w8297;
assign w8299 = ~w784 & ~w1449;
assign w8300 = ~w8298 & w18878;
assign w8301 = ~w8290 & w8300;
assign w8302 = (pi012 & ~w8301) | (pi012 & w18879) | (~w8301 & w18879);
assign w8303 = ~pi069 & w685;
assign w8304 = w604 & w626;
assign w8305 = w622 & w624;
assign w8306 = ~w8304 & ~w8305;
assign w8307 = ~w559 & ~w600;
assign w8308 = w8306 & ~w8307;
assign w8309 = ~w732 & ~w7488;
assign w8310 = ~pi104 & ~w8309;
assign w8311 = ~w583 & ~w718;
assign w8312 = w668 & ~w8311;
assign w8313 = ~w569 & ~w686;
assign w8314 = w640 & ~w8313;
assign w8315 = ~w1471 & ~w8310;
assign w8316 = ~w8312 & ~w8314;
assign w8317 = w8315 & w8316;
assign w8318 = pi102 & ~w8308;
assign w8319 = w8317 & ~w8318;
assign w8320 = ~w774 & ~w840;
assign w8321 = (~pi104 & ~w8320) | (~pi104 & w18880) | (~w8320 & w18880);
assign w8322 = (pi104 & w5504) | (pi104 & w18881) | (w5504 & w18881);
assign w8323 = w620 & w627;
assign w8324 = ~w7651 & ~w8323;
assign w8325 = ~w8322 & w8324;
assign w8326 = ~w8321 & w8325;
assign w8327 = ~w618 & ~w736;
assign w8328 = w597 & ~w8327;
assign w8329 = ~pi104 & w676;
assign w8330 = ~w884 & ~w8329;
assign w8331 = ~w813 & ~w8328;
assign w8332 = (pi102 & ~w8331) | (pi102 & w18882) | (~w8331 & w18882);
assign w8333 = w585 & w711;
assign w8334 = pi063 & w7473;
assign w8335 = ~w8333 & ~w8334;
assign w8336 = ~w8332 & w8335;
assign w8337 = ~pi102 & ~w8326;
assign w8338 = w8336 & ~w8337;
assign w8339 = (~pi012 & ~w8319) | (~pi012 & w18883) | (~w8319 & w18883);
assign w8340 = w8338 & ~w8339;
assign w8341 = ~w8302 & w8340;
assign w8342 = w8340 & w18884;
assign w8343 = (pi164 & ~w8340) | (pi164 & w18885) | (~w8340 & w18885);
assign w8344 = ~w8342 & ~w8343;
assign w8345 = w1131 & ~w5651;
assign w8346 = ~w1131 & w5651;
assign w8347 = ~w8345 & ~w8346;
assign w8348 = (~pi529 & w8347) | (~pi529 & w18886) | (w8347 & w18886);
assign w8349 = ~w8344 & w8347;
assign w8350 = w8348 & ~w8349;
assign w8351 = pi164 & pi448;
assign w8352 = pi529 & ~w8351;
assign w8353 = ~pi164 & ~pi448;
assign w8354 = w8352 & ~w8353;
assign w8355 = ~w8350 & ~w8354;
assign w8356 = w8340 & w18887;
assign w8357 = (pi154 & ~w8340) | (pi154 & w18888) | (~w8340 & w18888);
assign w8358 = ~w8356 & ~w8357;
assign w8359 = ~w145 & w5648;
assign w8360 = w145 & ~w5648;
assign w8361 = ~w8359 & ~w8360;
assign w8362 = ~w1128 & w1206;
assign w8363 = w1128 & ~w1206;
assign w8364 = ~w8362 & ~w8363;
assign w8365 = w8361 & w8364;
assign w8366 = ~w8361 & ~w8364;
assign w8367 = ~w8365 & ~w8366;
assign w8368 = (~pi529 & ~w8367) | (~pi529 & w18889) | (~w8367 & w18889);
assign w8369 = ~w8358 & ~w8367;
assign w8370 = w8368 & ~w8369;
assign w8371 = pi154 & pi516;
assign w8372 = pi529 & ~w8371;
assign w8373 = ~pi154 & ~pi516;
assign w8374 = w8372 & ~w8373;
assign w8375 = ~w8370 & ~w8374;
assign w8376 = w2071 & w2098;
assign w8377 = ~pi092 & ~w2065;
assign w8378 = pi085 & w2157;
assign w8379 = w8377 & ~w8378;
assign w8380 = pi092 & ~w8376;
assign w8381 = ~w8379 & ~w8380;
assign w8382 = ~w2078 & ~w5792;
assign w8383 = ~pi092 & ~w8382;
assign w8384 = ~pi089 & w2107;
assign w8385 = pi092 & ~w2132;
assign w8386 = w8384 & ~w8385;
assign w8387 = ~w2186 & ~w8386;
assign w8388 = ~w8383 & w8387;
assign w8389 = ~pi053 & w8388;
assign w8390 = w2085 & w18891;
assign w8391 = (~pi089 & w2189) | (~pi089 & w18892) | (w2189 & w18892);
assign w8392 = pi092 & w2095;
assign w8393 = pi085 & w2085;
assign w8394 = (pi087 & w8393) | (pi087 & w18893) | (w8393 & w18893);
assign w8395 = w2085 & w2048;
assign w8396 = w2083 & w2111;
assign w8397 = (~pi092 & w8396) | (~pi092 & w20819) | (w8396 & w20819);
assign w8398 = w8392 & w8394;
assign w8399 = ~w8397 & ~w8398;
assign w8400 = w8389 & w8399;
assign w8401 = w8400 & w18894;
assign w8402 = ~w2115 & ~w5859;
assign w8403 = w2060 & ~w8402;
assign w8404 = ~w5848 & w5868;
assign w8405 = w2056 & w5848;
assign w8406 = ~w2062 & w5854;
assign w8407 = ~w8405 & ~w8406;
assign w8408 = ~w2053 & w8404;
assign w8409 = w8407 & ~w8408;
assign w8410 = (~pi089 & ~w8409) | (~pi089 & w18895) | (~w8409 & w18895);
assign w8411 = pi092 & ~w2124;
assign w8412 = ~w2083 & w8411;
assign w8413 = pi085 & w2073;
assign w8414 = ~pi028 & w2085;
assign w8415 = ~w8413 & ~w8414;
assign w8416 = w8412 & w8415;
assign w8417 = ~pi092 & ~w2180;
assign w8418 = w2053 & w2095;
assign w8419 = (~w8418 & w8416) | (~w8418 & w18896) | (w8416 & w18896);
assign w8420 = pi089 & ~w8419;
assign w8421 = w2092 & w5848;
assign w8422 = w2051 & w2052;
assign w8423 = ~w5786 & ~w8421;
assign w8424 = (pi092 & ~w8423) | (pi092 & w18897) | (~w8423 & w18897);
assign w8425 = (w2092 & w5854) | (w2092 & w2139) | (w5854 & w2139);
assign w8426 = (pi053 & ~w2185) | (pi053 & w18898) | (~w2185 & w18898);
assign w8427 = ~w8425 & w8426;
assign w8428 = ~w8424 & w8427;
assign w8429 = ~w8420 & w8428;
assign w8430 = ~w8410 & w8429;
assign w8431 = ~w8401 & ~w8430;
assign w8432 = w2048 & w2075;
assign w8433 = w2085 & w2163;
assign w8434 = ~w8422 & ~w8432;
assign w8435 = ~pi028 & ~w8433;
assign w8436 = w8434 & w8435;
assign w8437 = w2049 & w2132;
assign w8438 = ~w2109 & ~w8437;
assign w8439 = (w8438 & w8436) | (w8438 & w18899) | (w8436 & w18899);
assign w8440 = ~w2107 & w5848;
assign w8441 = (pi028 & ~w5835) | (pi028 & w18900) | (~w5835 & w18900);
assign w8442 = ~pi092 & ~w8441;
assign w8443 = w2071 & w2077;
assign w8444 = ~w8418 & w18901;
assign w8445 = w2177 & ~w8444;
assign w8446 = ~w2158 & ~w5844;
assign w8447 = w5805 & ~w8446;
assign w8448 = w2115 & w2126;
assign w8449 = ~w2178 & ~w8448;
assign w8450 = ~w8383 & w8449;
assign w8451 = ~pi089 & ~w8450;
assign w8452 = ~w8451 & w18902;
assign w8453 = ~w8439 & ~w8442;
assign w8454 = pi089 & w8453;
assign w8455 = w8452 & ~w8454;
assign w8456 = ~w8431 & w8455;
assign w8457 = ~w2093 & ~w2166;
assign w8458 = w2075 & w2111;
assign w8459 = ~w2063 & ~w8458;
assign w8460 = w2049 & w5823;
assign w8461 = ~w2178 & ~w5806;
assign w8462 = w8459 & w8461;
assign w8463 = ~w8460 & w8462;
assign w8464 = (pi089 & ~w8463) | (pi089 & w18904) | (~w8463 & w18904);
assign w8465 = ~w2059 & ~w5814;
assign w8466 = (pi092 & ~w8465) | (pi092 & w18905) | (~w8465 & w18905);
assign w8467 = w2052 & w2098;
assign w8468 = ~w2065 & ~w8467;
assign w8469 = ~pi092 & ~w8468;
assign w8470 = ~w2090 & ~w5844;
assign w8471 = ~w2159 & w8470;
assign w8472 = ~w8469 & w8471;
assign w8473 = (~pi089 & ~w8472) | (~pi089 & w18906) | (~w8472 & w18906);
assign w8474 = w2098 & w2107;
assign w8475 = ~w2094 & w18907;
assign w8476 = ~pi092 & ~w8475;
assign w8477 = ~w2050 & ~w8432;
assign w8478 = pi050 & w2095;
assign w8479 = w2095 & w2075;
assign w8480 = (pi092 & ~w8477) | (pi092 & w18908) | (~w8477 & w18908);
assign w8481 = w2056 & w2059;
assign w8482 = ~w8480 & ~w8481;
assign w8483 = ~w8476 & w8482;
assign w8484 = ~w8464 & ~w8473;
assign w8485 = (pi053 & ~w8484) | (pi053 & w18909) | (~w8484 & w18909);
assign w8486 = ~pi085 & w2121;
assign w8487 = w2059 & w2092;
assign w8488 = w2107 & w5802;
assign w8489 = ~pi085 & w2078;
assign w8490 = ~pi046 & w8488;
assign w8491 = ~w8489 & ~w8490;
assign w8492 = ~w2112 & ~w5814;
assign w8493 = w8491 & w8492;
assign w8494 = ~w2073 & w2140;
assign w8495 = ~w8474 & ~w8494;
assign w8496 = w2111 & w2127;
assign w8497 = ~w5802 & w8393;
assign w8498 = ~w8496 & ~w8497;
assign w8499 = w8495 & w8498;
assign w8500 = ~pi089 & ~w8499;
assign w8501 = w2049 & w2095;
assign w8502 = ~w2179 & ~w8501;
assign w8503 = w2062 & w2167;
assign w8504 = ~w5834 & ~w8503;
assign w8505 = pi092 & ~w8504;
assign w8506 = pi046 & w2121;
assign w8507 = w2051 & w8506;
assign w8508 = ~w8505 & ~w8507;
assign w8509 = (~pi092 & w2179) | (~pi092 & w18912) | (w2179 & w18912);
assign w8510 = w8508 & ~w8509;
assign w8511 = ~w8500 & w8510;
assign w8512 = (~pi053 & ~w8511) | (~pi053 & w18913) | (~w8511 & w18913);
assign w8513 = w2056 & w20820;
assign w8514 = (pi092 & ~w8459) | (pi092 & w20821) | (~w8459 & w20821);
assign w8515 = w2075 & w2163;
assign w8516 = ~pi085 & w2049;
assign w8517 = ~w8413 & ~w8515;
assign w8518 = (w5823 & ~w8517) | (w5823 & w18914) | (~w8517 & w18914);
assign w8519 = w2126 & w5799;
assign w8520 = (pi089 & ~w18915) | (pi089 & w20822) | (~w18915 & w20822);
assign w8521 = w2060 & w2125;
assign w8522 = ~w2152 & ~w8521;
assign w8523 = w2177 & ~w8522;
assign w8524 = ~w2109 & ~w8432;
assign w8525 = w2187 & ~w8524;
assign w8526 = ~pi089 & ~pi092;
assign w8527 = w2057 & w8526;
assign w8528 = ~w2066 & ~w8527;
assign w8529 = ~w8525 & w8528;
assign w8530 = ~w8523 & w8529;
assign w8531 = ~w8520 & w8530;
assign w8532 = ~w8512 & w8531;
assign w8533 = ~w8485 & w8532;
assign w8534 = ~w8456 & w8533;
assign w8535 = w8456 & ~w8533;
assign w8536 = ~w8534 & ~w8535;
assign w8537 = pi059 & pi115;
assign w8538 = w1767 & w8537;
assign w8539 = ~pi056 & w1744;
assign w8540 = w1744 & w18916;
assign w8541 = w1982 & w1984;
assign w8542 = ~w8540 & ~w8541;
assign w8543 = ~w1729 & ~w8538;
assign w8544 = ~pi026 & w8543;
assign w8545 = w8542 & w8544;
assign w8546 = ~pi115 & w1708;
assign w8547 = w1693 & w1695;
assign w8548 = pi026 & ~w8547;
assign w8549 = ~w1983 & w8548;
assign w8550 = w1702 & w1732;
assign w8551 = w8549 & ~w8550;
assign w8552 = ~w2000 & w8546;
assign w8553 = ~w1705 & w8552;
assign w8554 = w8551 & ~w8553;
assign w8555 = w1693 & w1723;
assign w8556 = ~w1789 & ~w8555;
assign w8557 = pi115 & ~w8556;
assign w8558 = (pi008 & ~w1727) | (pi008 & w18917) | (~w1727 & w18917);
assign w8559 = ~w8556 & w18918;
assign w8560 = w1706 & w1984;
assign w8561 = ~w2010 & ~w8560;
assign w8562 = ~w8559 & w8561;
assign w8563 = (w8562 & w8554) | (w8562 & w18919) | (w8554 & w18919);
assign w8564 = ~pi030 & ~w8563;
assign w8565 = ~w1810 & ~w1820;
assign w8566 = ~pi115 & ~w8565;
assign w8567 = w1708 & w1771;
assign w8568 = ~w2253 & ~w8567;
assign w8569 = (pi026 & ~w2000) | (pi026 & w18920) | (~w2000 & w18920);
assign w8570 = ~w8566 & w8568;
assign w8571 = w8569 & w8570;
assign w8572 = w1736 & ~w2240;
assign w8573 = w1708 & w1715;
assign w8574 = pi115 & w8573;
assign w8575 = w1704 & w1737;
assign w8576 = ~w8572 & ~w8574;
assign w8577 = w8576 & w18921;
assign w8578 = w1695 & w1737;
assign w8579 = ~w2212 & ~w8578;
assign w8580 = ~w2018 & w8579;
assign w8581 = ~pi115 & w8580;
assign w8582 = ~w1806 & ~w8540;
assign w8583 = pi115 & ~w2020;
assign w8584 = ~w1943 & ~w2252;
assign w8585 = w8583 & w8584;
assign w8586 = w8582 & w8585;
assign w8587 = ~w8571 & ~w8577;
assign w8588 = ~w8581 & ~w8586;
assign w8589 = (pi030 & w8587) | (pi030 & w18922) | (w8587 & w18922);
assign w8590 = ~w1775 & ~w1824;
assign w8591 = ~w2262 & w8590;
assign w8592 = ~w2029 & ~w2257;
assign w8593 = w8591 & w8592;
assign w8594 = pi115 & ~w8593;
assign w8595 = w1700 & w1701;
assign w8596 = ~w2241 & ~w8595;
assign w8597 = ~w2215 & w8596;
assign w8598 = ~pi115 & ~w8597;
assign w8599 = ~w1716 & ~w2010;
assign w8600 = ~pi026 & w8599;
assign w8601 = ~w8598 & w8600;
assign w8602 = ~pi059 & w1718;
assign w8603 = w1696 & ~w1723;
assign w8604 = ~w2018 & ~w8603;
assign w8605 = (~pi115 & ~w8604) | (~pi115 & w18923) | (~w8604 & w18923);
assign w8606 = ~w1782 & ~w1965;
assign w8607 = pi026 & w8606;
assign w8608 = ~w8605 & w8607;
assign w8609 = ~w8594 & w8601;
assign w8610 = w1730 & w2009;
assign w8611 = (w2265 & w8610) | (w2265 & w18924) | (w8610 & w18924);
assign w8612 = w1734 & w2007;
assign w8613 = (pi008 & w8612) | (pi008 & w18925) | (w8612 & w18925);
assign w8614 = ~w8611 & ~w8613;
assign w8615 = ~w8564 & ~w8589;
assign w8616 = (w8614 & w8609) | (w8614 & w18926) | (w8609 & w18926);
assign w8617 = w8615 & w8616;
assign w8618 = w1544 & w1634;
assign w8619 = ~pi032 & w1554;
assign w8620 = ~w8618 & ~w8619;
assign w8621 = ~pi117 & ~w8620;
assign w8622 = ~pi105 & w1549;
assign w8623 = w1564 & w8622;
assign w8624 = w1625 & w1634;
assign w8625 = ~w1917 & ~w8623;
assign w8626 = pi002 & ~w8624;
assign w8627 = w8625 & w8626;
assign w8628 = w1543 & w1623;
assign w8629 = ~pi002 & ~w8628;
assign w8630 = ~w1885 & w8629;
assign w8631 = ~pi032 & ~pi117;
assign w8632 = ~pi067 & ~w8631;
assign w8633 = w1559 & ~w8632;
assign w8634 = w1578 & w1634;
assign w8635 = pi117 & w8634;
assign w8636 = ~w8633 & ~w8635;
assign w8637 = w8630 & w8636;
assign w8638 = ~w8621 & w8627;
assign w8639 = ~w8637 & ~w8638;
assign w8640 = ~pi032 & w1558;
assign w8641 = ~w1919 & ~w8622;
assign w8642 = ~w8640 & w8641;
assign w8643 = w1543 & w1555;
assign w8644 = ~pi117 & ~w8643;
assign w8645 = w1554 & w1623;
assign w8646 = ~w1918 & w8644;
assign w8647 = ~w8645 & w8646;
assign w8648 = pi117 & ~w1650;
assign w8649 = w8642 & w8648;
assign w8650 = ~w8647 & ~w8649;
assign w8651 = pi036 & ~w8650;
assign w8652 = ~w8639 & w8651;
assign w8653 = ~w1616 & ~w1679;
assign w8654 = ~pi002 & ~w8653;
assign w8655 = pi117 & ~w1884;
assign w8656 = ~pi064 & w1601;
assign w8657 = w8655 & ~w8656;
assign w8658 = ~w1638 & ~w1878;
assign w8659 = ~w8657 & w8658;
assign w8660 = ~w8654 & ~w8659;
assign w8661 = pi064 & w1623;
assign w8662 = ~w1544 & w1634;
assign w8663 = ~w8661 & w8662;
assign w8664 = pi002 & w8663;
assign w8665 = w1547 & ~w8664;
assign w8666 = ~w8660 & ~w8665;
assign w8667 = w1554 & w1552;
assign w8668 = w1554 & w1878;
assign w8669 = pi105 & w1927;
assign w8670 = w1544 & w8669;
assign w8671 = ~w8670 & w18927;
assign w8672 = pi002 & ~w8671;
assign w8673 = w1554 & w1639;
assign w8674 = w1582 & w1623;
assign w8675 = pi064 & w8673;
assign w8676 = (~pi002 & w8675) | (~pi002 & w18928) | (w8675 & w18928);
assign w8677 = ~pi036 & ~w1663;
assign w8678 = ~w8676 & w8677;
assign w8679 = ~w8672 & w8678;
assign w8680 = ~w8666 & w8679;
assign w8681 = ~w8652 & ~w8680;
assign w8682 = pi032 & pi117;
assign w8683 = w1914 & w8631;
assign w8684 = w1615 & w8682;
assign w8685 = w1567 & w1582;
assign w8686 = ~w1624 & ~w1664;
assign w8687 = ~w8685 & w8686;
assign w8688 = pi067 & w1634;
assign w8689 = w1544 & w8688;
assign w8690 = ~w1903 & ~w8689;
assign w8691 = w8687 & w8690;
assign w8692 = pi117 & ~w8691;
assign w8693 = pi067 & w1543;
assign w8694 = w1677 & w8693;
assign w8695 = w1543 & w1621;
assign w8696 = ~w1550 & ~w8695;
assign w8697 = ~w8694 & w8696;
assign w8698 = ~pi117 & ~w8697;
assign w8699 = ~w1574 & ~w1663;
assign w8700 = ~pi002 & w8699;
assign w8701 = ~w8698 & w8700;
assign w8702 = w1555 & ~w1582;
assign w8703 = ~w1658 & ~w1918;
assign w8704 = (~pi117 & ~w8703) | (~pi117 & w18929) | (~w8703 & w18929);
assign w8705 = w1577 & w1892;
assign w8706 = w1554 & w1915;
assign w8707 = ~w1873 & ~w8706;
assign w8708 = ~w1633 & ~w8705;
assign w8709 = w8707 & w8708;
assign w8710 = pi002 & w8709;
assign w8711 = ~w8692 & w8701;
assign w8712 = ~w8704 & w8710;
assign w8713 = ~w8711 & ~w8712;
assign w8714 = (pi067 & w8683) | (pi067 & w18930) | (w8683 & w18930);
assign w8715 = ~w8713 & ~w8714;
assign w8716 = ~w8681 & w8715;
assign w8717 = ~w8617 & w8716;
assign w8718 = w8617 & ~w8716;
assign w8719 = ~w8717 & ~w8718;
assign w8720 = w8536 & ~w8719;
assign w8721 = ~w8536 & w8719;
assign w8722 = ~w8720 & ~w8721;
assign w8723 = pi110 & w2346;
assign w8724 = ~w2404 & ~w5695;
assign w8725 = ~w5696 & ~w5709;
assign w8726 = ~pi080 & ~w8725;
assign w8727 = w2293 & w2328;
assign w8728 = ~w2348 & ~w8727;
assign w8729 = ~w5748 & w8728;
assign w8730 = ~w8726 & w8729;
assign w8731 = ~pi075 & w2333;
assign w8732 = w2314 & w2328;
assign w8733 = pi080 & ~w8732;
assign w8734 = ~pi080 & ~w2397;
assign w8735 = ~w8731 & w8733;
assign w8736 = ~w8734 & ~w8735;
assign w8737 = w2337 & w2359;
assign w8738 = ~w2350 & ~w8737;
assign w8739 = ~w2400 & w8738;
assign w8740 = ~pi080 & w2295;
assign w8741 = w2359 & w18932;
assign w8742 = ~w8740 & ~w8741;
assign w8743 = w8739 & w8742;
assign w8744 = ~w8736 & w8743;
assign w8745 = pi110 & w2384;
assign w8746 = w2293 & w2376;
assign w8747 = ~w5710 & ~w8746;
assign w8748 = ~w8745 & w8747;
assign w8749 = ~pi080 & ~w8748;
assign w8750 = pi075 & pi080;
assign w8751 = ~w2303 & ~w5733;
assign w8752 = (w8750 & ~w8751) | (w8750 & w18933) | (~w8751 & w18933);
assign w8753 = w2306 & w2326;
assign w8754 = ~w8749 & w18934;
assign w8755 = ~pi073 & ~w8744;
assign w8756 = ~pi071 & ~pi110;
assign w8757 = ~pi075 & w8756;
assign w8758 = w2298 & w5707;
assign w8759 = (pi080 & w8758) | (pi080 & w18936) | (w8758 & w18936);
assign w8760 = w2306 & w5693;
assign w8761 = ~pi042 & w8760;
assign w8762 = ~w5754 & ~w8761;
assign w8763 = ~w2361 & ~w8732;
assign w8764 = w8762 & w8763;
assign w8765 = ~w2316 & w5683;
assign w8766 = pi110 & w8765;
assign w8767 = ~w5710 & ~w8766;
assign w8768 = ~w2325 & ~w8750;
assign w8769 = w2329 & ~w8768;
assign w8770 = w2342 & w2348;
assign w8771 = ~w8769 & ~w8770;
assign w8772 = w8767 & w8771;
assign w8773 = ~pi073 & ~w8772;
assign w8774 = w2299 & w2302;
assign w8775 = ~w2416 & ~w8774;
assign w8776 = (~pi080 & w2416) | (~pi080 & w18937) | (w2416 & w18937);
assign w8777 = w5715 & w8756;
assign w8778 = ~w2343 & ~w8777;
assign w8779 = pi080 & ~w8778;
assign w8780 = w2357 & w5709;
assign w8781 = ~w8779 & ~w8780;
assign w8782 = ~w8776 & w8781;
assign w8783 = ~w8773 & w8782;
assign w8784 = (pi073 & ~w8764) | (pi073 & w18938) | (~w8764 & w18938);
assign w8785 = pi071 & w5715;
assign w8786 = w5715 & w2359;
assign w8787 = (pi080 & ~w8728) | (pi080 & w18939) | (~w8728 & w18939);
assign w8788 = ~pi075 & w2299;
assign w8789 = ~w2369 & ~w5706;
assign w8790 = (w2345 & ~w8789) | (w2345 & w18940) | (~w8789 & w18940);
assign w8791 = ~pi080 & w8732;
assign w8792 = w8732 & w18941;
assign w8793 = ~w8787 & ~w8790;
assign w8794 = (pi073 & ~w8793) | (pi073 & w18942) | (~w8793 & w18942);
assign w8795 = ~w2396 & ~w8780;
assign w8796 = w2415 & ~w8795;
assign w8797 = ~w2358 & ~w2422;
assign w8798 = w2421 & ~w8797;
assign w8799 = w2293 & w5715;
assign w8800 = ~pi073 & ~pi080;
assign w8801 = w8799 & w8800;
assign w8802 = ~w2304 & ~w8801;
assign w8803 = ~w8798 & w8802;
assign w8804 = ~w8796 & w8803;
assign w8805 = ~w8794 & w8804;
assign w8806 = (~pi015 & ~w8783) | (~pi015 & w18943) | (~w8783 & w18943);
assign w8807 = w8805 & ~w8806;
assign w8808 = (w8755 & w20823) | (w8755 & w20824) | (w20823 & w20824);
assign w8809 = w8807 & ~w8808;
assign w8810 = ~w5779 & w8809;
assign w8811 = w5779 & ~w8809;
assign w8812 = ~w8810 & ~w8811;
assign w8813 = ~w2302 & ~w2337;
assign w8814 = (pi071 & ~w5737) | (pi071 & w18945) | (~w5737 & w18945);
assign w8815 = w5733 & ~w8813;
assign w8816 = (pi080 & w8814) | (pi080 & w18946) | (w8814 & w18946);
assign w8817 = ~w5726 & ~w8757;
assign w8818 = ~pi080 & w8817;
assign w8819 = ~w2290 & ~w8799;
assign w8820 = w8818 & ~w8819;
assign w8821 = w2342 & w2370;
assign w8822 = w2410 & w2421;
assign w8823 = ~w8821 & ~w8822;
assign w8824 = ~w5688 & ~w5757;
assign w8825 = w8823 & w8824;
assign w8826 = ~pi073 & w8825;
assign w8827 = ~pi075 & w2329;
assign w8828 = w2294 & w8827;
assign w8829 = w2328 & ~w2329;
assign w8830 = ~w5754 & ~w8828;
assign w8831 = (~pi080 & ~w8830) | (~pi080 & w18947) | (~w8830 & w18947);
assign w8832 = w2421 & w5766;
assign w8833 = ~pi042 & w5746;
assign w8834 = ~w5732 & ~w8832;
assign w8835 = (pi073 & ~w5746) | (pi073 & w18948) | (~w5746 & w18948);
assign w8836 = w8834 & w8835;
assign w8837 = w2299 & w5683;
assign w8838 = pi075 & w8837;
assign w8839 = w8823 & ~w8838;
assign w8840 = w8836 & w8839;
assign w8841 = ~w8831 & w8840;
assign w8842 = w8826 & w18949;
assign w8843 = ~w8841 & ~w8842;
assign w8844 = ~w2325 & w5693;
assign w8845 = ~w8785 & w8844;
assign w8846 = ~pi042 & w8845;
assign w8847 = ~pi079 & w8750;
assign w8848 = w2363 & w8847;
assign w8849 = ~w8774 & ~w8848;
assign w8850 = pi073 & ~w8741;
assign w8851 = ~w8846 & w8849;
assign w8852 = w8850 & w8851;
assign w8853 = ~w2410 & ~w5696;
assign w8854 = pi080 & ~w8853;
assign w8855 = ~pi080 & w2300;
assign w8856 = w2329 & w5715;
assign w8857 = ~pi073 & ~w8856;
assign w8858 = ~w8855 & w8857;
assign w8859 = ~w8854 & w8858;
assign w8860 = pi042 & w2357;
assign w8861 = w2302 & w2329;
assign w8862 = ~w8860 & ~w8861;
assign w8863 = pi080 & ~w8862;
assign w8864 = (pi079 & ~w2329) | (pi079 & w2376) | (~w2329 & w2376);
assign w8865 = ~w8862 & w18950;
assign w8866 = w2306 & w2329;
assign w8867 = w2312 & w5693;
assign w8868 = (~pi079 & w8867) | (~pi079 & w18951) | (w8867 & w18951);
assign w8869 = ~w8865 & ~w8868;
assign w8870 = ~pi015 & w8869;
assign w8871 = ~w8852 & ~w8859;
assign w8872 = w8870 & ~w8871;
assign w8873 = ~w2422 & ~w8788;
assign w8874 = ~pi080 & ~w8873;
assign w8875 = w2333 & w5716;
assign w8876 = w2314 & w2368;
assign w8877 = ~w2396 & ~w8875;
assign w8878 = pi073 & ~w8876;
assign w8879 = w8877 & w8878;
assign w8880 = (~pi073 & ~w8861) | (~pi073 & w2415) | (~w8861 & w2415);
assign w8881 = ~w2393 & ~w8760;
assign w8882 = ~w8799 & w8881;
assign w8883 = pi080 & w2348;
assign w8884 = ~w8874 & w8879;
assign w8885 = w8882 & w18952;
assign w8886 = ~w8884 & ~w8885;
assign w8887 = ~pi110 & w2381;
assign w8888 = ~w2343 & ~w5716;
assign w8889 = w8733 & w8888;
assign w8890 = ~w8887 & w8889;
assign w8891 = ~pi080 & ~w8727;
assign w8892 = w2299 & w5715;
assign w8893 = ~w8828 & w8891;
assign w8894 = ~w8892 & w8893;
assign w8895 = ~w8890 & ~w8894;
assign w8896 = pi015 & ~w8895;
assign w8897 = ~w8886 & w8896;
assign w8898 = ~w8872 & ~w8897;
assign w8899 = ~w8843 & ~w8898;
assign w8900 = ~w8898 & w18953;
assign w8901 = (pi301 & w8898) | (pi301 & w18954) | (w8898 & w18954);
assign w8902 = ~w8900 & ~w8901;
assign w8903 = w8812 & w8902;
assign w8904 = ~w8812 & ~w8902;
assign w8905 = ~w8903 & ~w8904;
assign w8906 = (~pi529 & ~w8905) | (~pi529 & w18955) | (~w8905 & w18955);
assign w8907 = w8722 & ~w8905;
assign w8908 = w8906 & ~w8907;
assign w8909 = ~pi301 & pi512;
assign w8910 = pi529 & ~w8909;
assign w8911 = pi301 & ~pi512;
assign w8912 = w8910 & ~w8911;
assign w8913 = ~w8908 & ~w8912;
assign w8914 = ~w1818 & ~w1982;
assign w8915 = pi115 & w8914;
assign w8916 = ~w1697 & ~w2241;
assign w8917 = ~pi115 & w8916;
assign w8918 = ~w8915 & ~w8917;
assign w8919 = ~w2028 & ~w2222;
assign w8920 = ~w2021 & w8919;
assign w8921 = ~w2257 & w8920;
assign w8922 = ~w8918 & w8921;
assign w8923 = ~pi026 & ~w8922;
assign w8924 = ~w1705 & ~w1760;
assign w8925 = pi099 & ~w8924;
assign w8926 = (pi115 & w8925) | (pi115 & w18956) | (w8925 & w18956);
assign w8927 = ~w2274 & ~w8573;
assign w8928 = w1695 & w1984;
assign w8929 = w8927 & ~w8928;
assign w8930 = ~w1836 & ~w2212;
assign w8931 = w8929 & w8930;
assign w8932 = w1766 & w1783;
assign w8933 = ~w1991 & w18957;
assign w8934 = ~pi115 & ~w8933;
assign w8935 = ~w1940 & ~w2007;
assign w8936 = (w8537 & ~w8935) | (w8537 & w18958) | (~w8935 & w18958);
assign w8937 = pi008 & w2261;
assign w8938 = ~w8936 & ~w8937;
assign w8939 = ~w8934 & w8938;
assign w8940 = (pi026 & ~w8931) | (pi026 & w18959) | (~w8931 & w18959);
assign w8941 = w8939 & ~w8940;
assign w8942 = ~w8923 & w8941;
assign w8943 = pi030 & ~w8942;
assign w8944 = ~pi059 & w1804;
assign w8945 = w1767 & w2252;
assign w8946 = (pi115 & w8945) | (pi115 & w18960) | (w8945 & w18960);
assign w8947 = w1760 & w1766;
assign w8948 = ~pi115 & w8947;
assign w8949 = ~w8602 & ~w8948;
assign w8950 = pi026 & ~w2020;
assign w8951 = ~w2230 & w8950;
assign w8952 = w8949 & w8951;
assign w8953 = w1715 & w8546;
assign w8954 = w8546 & w18961;
assign w8955 = ~w1705 & ~w8537;
assign w8956 = w1723 & ~w8955;
assign w8957 = ~w1727 & w1773;
assign w8958 = pi099 & w8957;
assign w8959 = ~pi026 & ~w8932;
assign w8960 = ~w8956 & ~w8958;
assign w8961 = ~w8946 & w8952;
assign w8962 = w8960 & w18962;
assign w8963 = ~w8961 & ~w8962;
assign w8964 = w1696 & w1744;
assign w8965 = ~w1806 & ~w8964;
assign w8966 = ~w2269 & ~w8547;
assign w8967 = (~pi115 & w2269) | (~pi115 & w18963) | (w2269 & w18963);
assign w8968 = ~w2008 & ~w8967;
assign w8969 = (~pi030 & w8963) | (~pi030 & w18964) | (w8963 & w18964);
assign w8970 = ~w1753 & ~w1810;
assign w8971 = (w1984 & ~w8970) | (w1984 & w18965) | (~w8970 & w18965);
assign w8972 = ~pi056 & w1696;
assign w8973 = w1735 & w8972;
assign w8974 = ~w8574 & ~w8973;
assign w8975 = ~w8971 & w8974;
assign w8976 = pi026 & ~w8975;
assign w8977 = w1773 & w1805;
assign w8978 = ~w2253 & ~w8977;
assign w8979 = w1996 & ~w8978;
assign w8980 = w1737 & w1767;
assign w8981 = ~w2212 & ~w8980;
assign w8982 = ~pi026 & ~pi115;
assign w8983 = w8575 & w8982;
assign w8984 = ~w2216 & ~w8983;
assign w8985 = w1730 & ~w1821;
assign w8986 = w8984 & ~w8985;
assign w8987 = w2265 & ~w8981;
assign w8988 = w8986 & ~w8987;
assign w8989 = ~w8979 & w8988;
assign w8990 = ~w8976 & w8989;
assign w8991 = ~w8969 & w8990;
assign w8992 = ~w8943 & w8991;
assign w8993 = ~pi032 & w1569;
assign w8994 = ~w1919 & ~w8993;
assign w8995 = ~w1556 & ~w8695;
assign w8996 = ~pi117 & ~w8995;
assign w8997 = ~w1662 & ~w1902;
assign w8998 = ~w8668 & w8997;
assign w8999 = ~w8996 & w8998;
assign w9000 = ~w1544 & ~w1608;
assign w9001 = pi105 & ~w9000;
assign w9002 = (pi117 & w9001) | (pi117 & w18966) | (w9001 & w18966);
assign w9003 = ~w1683 & ~w8634;
assign w9004 = ~w8643 & ~w8673;
assign w9005 = w9003 & w9004;
assign w9006 = ~w1867 & w9005;
assign w9007 = (pi002 & ~w9006) | (pi002 & w18967) | (~w9006 & w18967);
assign w9008 = ~w1684 & ~w8693;
assign w9009 = ~w1555 & ~w9008;
assign w9010 = (~pi117 & w9009) | (~pi117 & w18968) | (w9009 & w18968);
assign w9011 = ~w1554 & ~w1634;
assign w9012 = ~pi064 & ~w9011;
assign w9013 = (w8682 & w9012) | (w8682 & w18969) | (w9012 & w18969);
assign w9014 = ~w1906 & ~w9013;
assign w9015 = ~w9010 & w9014;
assign w9016 = ~w9007 & w9015;
assign w9017 = (pi036 & ~w9016) | (pi036 & w18970) | (~w9016 & w18970);
assign w9018 = pi064 & w1543;
assign w9019 = w1552 & w9018;
assign w9020 = w1607 & w1927;
assign w9021 = ~pi032 & w1651;
assign w9022 = w1895 & w8631;
assign w9023 = w1651 & w1625;
assign w9024 = ~w9022 & ~w9023;
assign w9025 = ~w9019 & ~w9020;
assign w9026 = w9024 & w9025;
assign w9027 = w1665 & w8634;
assign w9028 = ~w1544 & ~w8682;
assign w9029 = w1582 & ~w9028;
assign w9030 = ~w1564 & w8669;
assign w9031 = ~w9029 & ~w9030;
assign w9032 = ~w1622 & ~w9027;
assign w9033 = w9031 & w9032;
assign w9034 = ~pi002 & ~w9033;
assign w9035 = w1559 & w1672;
assign w9036 = w1577 & w9021;
assign w9037 = pi117 & w1650;
assign w9038 = ~w9036 & ~w9037;
assign w9039 = w1570 & w1914;
assign w9040 = w9038 & ~w9039;
assign w9041 = (~pi117 & w9035) | (~pi117 & w18972) | (w9035 & w18972);
assign w9042 = w9040 & ~w9041;
assign w9043 = ~w9034 & w9042;
assign w9044 = (~pi036 & ~w9043) | (~pi036 & w18973) | (~w9043 & w18973);
assign w9045 = w1634 & w1677;
assign w9046 = ~w1565 & ~w8619;
assign w9047 = (w1639 & ~w9046) | (w1639 & w18974) | (~w9046 & w18974);
assign w9048 = w1684 & w20825;
assign w9049 = ~w8635 & ~w9048;
assign w9050 = (pi002 & ~w9049) | (pi002 & w18975) | (~w9049 & w18975);
assign w9051 = pi002 & pi117;
assign w9052 = w1623 & w1615;
assign w9053 = ~w8643 & ~w9052;
assign w9054 = w1652 & w1927;
assign w9055 = ~w8623 & ~w9054;
assign w9056 = w1588 & ~w9055;
assign w9057 = ~w1666 & ~w8618;
assign w9058 = w1577 & ~w9057;
assign w9059 = w1544 & w1602;
assign w9060 = ~pi002 & ~pi117;
assign w9061 = w8628 & w9060;
assign w9062 = ~w9059 & ~w9061;
assign w9063 = ~w9058 & w9062;
assign w9064 = ~w9056 & w9063;
assign w9065 = w9051 & ~w9053;
assign w9066 = w9064 & ~w9065;
assign w9067 = ~w9050 & w9066;
assign w9068 = ~w9044 & w9067;
assign w9069 = ~w9017 & w9068;
assign w9070 = ~w8992 & w9069;
assign w9071 = w8992 & ~w9069;
assign w9072 = ~w9070 & ~w9071;
assign w9073 = w1844 & ~w9072;
assign w9074 = ~w1844 & w9072;
assign w9075 = ~w9073 & ~w9074;
assign w9076 = (pi092 & ~w2107) | (pi092 & w18976) | (~w2107 & w18976);
assign w9077 = ~w8432 & ~w8516;
assign w9078 = (~w9076 & ~w9077) | (~w9076 & w18977) | (~w9077 & w18977);
assign w9079 = ~w2152 & ~w5865;
assign w9080 = ~w9078 & w9079;
assign w9081 = pi089 & ~w9080;
assign w9082 = pi092 & ~w5834;
assign w9083 = ~pi085 & w2157;
assign w9084 = ~w5814 & ~w9083;
assign w9085 = ~pi050 & w2092;
assign w9086 = w9084 & ~w9085;
assign w9087 = w2049 & w2056;
assign w9088 = ~w2063 & ~w9087;
assign w9089 = ~w5863 & w9088;
assign w9090 = ~pi092 & w9089;
assign w9091 = w9082 & w9086;
assign w9092 = ~w9090 & ~w9091;
assign w9093 = pi092 & ~w8458;
assign w9094 = ~w5833 & ~w9093;
assign w9095 = pi028 & w2079;
assign w9096 = ~w2057 & ~w8488;
assign w9097 = ~w9095 & w9096;
assign w9098 = ~w9094 & w9097;
assign w9099 = (pi053 & w9098) | (pi053 & w18978) | (w9098 & w18978);
assign w9100 = ~w2048 & w2075;
assign w9101 = ~w5855 & w9100;
assign w9102 = ~pi092 & w9101;
assign w9103 = ~w5820 & ~w8501;
assign w9104 = ~w9102 & w9103;
assign w9105 = w2056 & w2085;
assign w9106 = w2071 & w18979;
assign w9107 = ~pi092 & w2130;
assign w9108 = ~w9106 & ~w9107;
assign w9109 = ~w8390 & ~w9105;
assign w9110 = (~pi089 & ~w9108) | (~pi089 & w18980) | (~w9108 & w18980);
assign w9111 = ~pi087 & w2124;
assign w9112 = ~w5832 & ~w9111;
assign w9113 = (pi028 & ~w2085) | (pi028 & w2132) | (~w2085 & w2132);
assign w9114 = ~w9112 & w18981;
assign w9115 = w2143 & w5823;
assign w9116 = (~pi053 & ~w2100) | (~pi053 & w18982) | (~w2100 & w18982);
assign w9117 = ~w9115 & w9116;
assign w9118 = ~w9114 & w9117;
assign w9119 = ~w9110 & w9118;
assign w9120 = (pi089 & ~w9104) | (pi089 & w18983) | (~w9104 & w18983);
assign w9121 = w9119 & ~w9120;
assign w9122 = ~w9081 & w9099;
assign w9123 = ~w9092 & w9122;
assign w9124 = ~w9121 & ~w9123;
assign w9125 = ~w2166 & ~w8405;
assign w9126 = pi092 & ~w8437;
assign w9127 = w9125 & w9126;
assign w9128 = ~w8376 & ~w8467;
assign w9129 = ~w8396 & w9128;
assign w9130 = w2091 & w9129;
assign w9131 = ~w2159 & ~w5845;
assign w9132 = w9127 & w9131;
assign w9133 = ~w9130 & ~w9132;
assign w9134 = w2062 & ~w2085;
assign w9135 = ~w5863 & ~w8489;
assign w9136 = (~pi092 & ~w9135) | (~pi092 & w18984) | (~w9135 & w18984);
assign w9137 = w2096 & w2187;
assign w9138 = ~w8418 & ~w9137;
assign w9139 = w2060 & w5859;
assign w9140 = (pi089 & ~w5814) | (pi089 & w18985) | (~w5814 & w18985);
assign w9141 = w9138 & w18986;
assign w9142 = ~w9136 & w9141;
assign w9143 = (~pi089 & ~w2100) | (~pi089 & w18987) | (~w2100 & w18987);
assign w9144 = ~w9133 & w9143;
assign w9145 = ~pi092 & w2125;
assign w9146 = (pi028 & w9145) | (pi028 & w18988) | (w9145 & w18988);
assign w9147 = (~w9146 & w9144) | (~w9146 & w20826) | (w9144 & w20826);
assign w9148 = ~w9124 & w9147;
assign w9149 = ~w8617 & w9148;
assign w9150 = w8617 & ~w9148;
assign w9151 = ~w9149 & ~w9150;
assign w9152 = ~w8898 & w18989;
assign w9153 = (pi184 & w8898) | (pi184 & w18990) | (w8898 & w18990);
assign w9154 = ~w9152 & ~w9153;
assign w9155 = w9151 & w9154;
assign w9156 = ~w9151 & ~w9154;
assign w9157 = ~w9155 & ~w9156;
assign w9158 = ~w9075 & w9157;
assign w9159 = ~pi529 & ~w9158;
assign w9160 = w9075 & ~w9157;
assign w9161 = w9159 & ~w9160;
assign w9162 = ~pi184 & pi442;
assign w9163 = pi529 & ~w9162;
assign w9164 = pi184 & ~pi442;
assign w9165 = w9163 & ~w9164;
assign w9166 = ~w9161 & ~w9165;
assign w9167 = w1695 & w1719;
assign w9168 = ~w1761 & ~w2236;
assign w9169 = (~pi115 & ~w9168) | (~pi115 & w18991) | (~w9168 & w18991);
assign w9170 = (pi115 & w8572) | (pi115 & w18992) | (w8572 & w18992);
assign w9171 = w1693 & w1736;
assign w9172 = ~w1809 & ~w2241;
assign w9173 = ~w8947 & ~w9171;
assign w9174 = w9172 & w9173;
assign w9175 = ~w9169 & ~w9170;
assign w9176 = ~w1811 & w9174;
assign w9177 = w9175 & w9176;
assign w9178 = w1773 & w1949;
assign w9179 = w1730 & w1956;
assign w9180 = ~w9178 & ~w9179;
assign w9181 = ~w1941 & ~w8602;
assign w9182 = w9180 & w9181;
assign w9183 = ~pi026 & ~w9182;
assign w9184 = ~w1942 & ~w8595;
assign w9185 = ~pi099 & ~w9184;
assign w9186 = ~w8539 & ~w9171;
assign w9187 = (pi115 & w9185) | (pi115 & w18993) | (w9185 & w18993);
assign w9188 = w1693 & w1804;
assign w9189 = ~w1817 & ~w9188;
assign w9190 = (~pi115 & ~w9189) | (~pi115 & w18994) | (~w9189 & w18994);
assign w9191 = ~w1745 & ~w9190;
assign w9192 = ~w9183 & w18995;
assign w9193 = pi026 & ~w9177;
assign w9194 = w9192 & ~w9193;
assign w9195 = ~w1773 & w1982;
assign w9196 = ~pi115 & w2020;
assign w9197 = ~w9195 & ~w9196;
assign w9198 = (~pi026 & ~w1787) | (~pi026 & w18996) | (~w1787 & w18996);
assign w9199 = ~w8557 & w9197;
assign w9200 = w9198 & w9199;
assign w9201 = (pi026 & ~w1959) | (pi026 & w18997) | (~w1959 & w18997);
assign w9202 = ~w1991 & ~w2253;
assign w9203 = w9202 & w18998;
assign w9204 = (~w2000 & w8925) | (~w2000 & w18999) | (w8925 & w18999);
assign w9205 = (~pi115 & w2205) | (~pi115 & w19000) | (w2205 & w19000);
assign w9206 = ~pi115 & w1706;
assign w9207 = w1702 & w1741;
assign w9208 = ~w9206 & ~w9207;
assign w9209 = ~w8937 & ~w8977;
assign w9210 = w9208 & w9209;
assign w9211 = ~w9205 & w9210;
assign w9212 = w2260 & ~w9204;
assign w9213 = w9211 & ~w9212;
assign w9214 = ~w9200 & ~w9203;
assign w9215 = w9213 & ~w9214;
assign w9216 = w1717 & w1766;
assign w9217 = ~w1706 & ~w9216;
assign w9218 = ~w1716 & w9217;
assign w9219 = ~pi026 & ~w9218;
assign w9220 = (~pi115 & w9219) | (~pi115 & w19001) | (w9219 & w19001);
assign w9221 = (w1702 & ~w8935) | (w1702 & w9207) | (~w8935 & w9207);
assign w9222 = w1731 & w1760;
assign w9223 = ~w2222 & ~w9222;
assign w9224 = ~w9221 & w9223;
assign w9225 = ~pi026 & ~w9224;
assign w9226 = w1759 & w1773;
assign w9227 = ~w8953 & ~w9226;
assign w9228 = pi008 & w1745;
assign w9229 = (pi026 & ~w9227) | (pi026 & w19002) | (~w9227 & w19002);
assign w9230 = ~w2015 & ~w9229;
assign w9231 = ~w9220 & ~w9225;
assign w9232 = w9230 & w9231;
assign w9233 = pi030 & ~w9215;
assign w9234 = w9232 & ~w9233;
assign w9235 = ~pi030 & ~w9194;
assign w9236 = w9234 & ~w9235;
assign w9237 = ~w1573 & ~w1919;
assign w9238 = ~pi117 & w9237;
assign w9239 = ~w8657 & ~w9238;
assign w9240 = pi105 & w8640;
assign w9241 = ~w8623 & ~w9240;
assign w9242 = w1857 & w9241;
assign w9243 = pi002 & ~w9242;
assign w9244 = pi002 & ~pi117;
assign w9245 = ~pi032 & w1564;
assign w9246 = pi032 & w1651;
assign w9247 = ~w8661 & ~w9245;
assign w9248 = (w9244 & ~w9247) | (w9244 & w19004) | (~w9247 & w19004);
assign w9249 = ~w1544 & w1602;
assign w9250 = (~pi117 & w9249) | (~pi117 & w19005) | (w9249 & w19005);
assign w9251 = ~pi117 & w1545;
assign w9252 = w1568 & w8682;
assign w9253 = ~w9251 & ~w9252;
assign w9254 = ~w1906 & ~w9054;
assign w9255 = w9253 & w9254;
assign w9256 = ~w9250 & w9255;
assign w9257 = ~w9243 & w9256;
assign w9258 = w9257 & w19006;
assign w9259 = ~pi067 & w8619;
assign w9260 = ~w1609 & ~w8688;
assign w9261 = ~w9259 & w9260;
assign w9262 = ~pi117 & ~w9261;
assign w9263 = (pi117 & w8633) | (pi117 & w19007) | (w8633 & w19007);
assign w9264 = pi064 & w1586;
assign w9265 = ~w1678 & ~w9264;
assign w9266 = ~w1674 & ~w8695;
assign w9267 = ~w9045 & w9266;
assign w9268 = w9265 & w9267;
assign w9269 = ~w9262 & ~w9263;
assign w9270 = pi067 & w1581;
assign w9271 = ~pi117 & w8634;
assign w9272 = ~w9020 & ~w9270;
assign w9273 = (pi002 & ~w9272) | (pi002 & w19008) | (~w9272 & w19008);
assign w9274 = w1582 & w1677;
assign w9275 = w1665 & w9274;
assign w9276 = ~pi117 & w8695;
assign w9277 = ~w1905 & ~w9276;
assign w9278 = ~w9275 & w9277;
assign w9279 = ~w9273 & w9278;
assign w9280 = pi002 & ~pi036;
assign w9281 = (w9280 & ~w9269) | (w9280 & w19009) | (~w9269 & w19009);
assign w9282 = w9279 & ~w9281;
assign w9283 = w1591 & w1567;
assign w9284 = ~w1574 & w19010;
assign w9285 = ~pi117 & ~w9284;
assign w9286 = (w1915 & w9012) | (w1915 & w19011) | (w9012 & w19011);
assign w9287 = w1553 & w1878;
assign w9288 = ~w1662 & ~w9287;
assign w9289 = ~w9286 & w9288;
assign w9290 = ~w9285 & w9289;
assign w9291 = ~pi002 & ~w9290;
assign w9292 = w1679 & w1927;
assign w9293 = w1577 & w9245;
assign w9294 = ~w9292 & ~w9293;
assign w9295 = w1661 & w9294;
assign w9296 = ~pi002 & ~w9295;
assign w9297 = w1586 & w1878;
assign w9298 = ~pi117 & w1666;
assign w9299 = w1665 & w9246;
assign w9300 = ~w9298 & ~w9299;
assign w9301 = w1582 & w1625;
assign w9302 = ~w1581 & ~w9301;
assign w9303 = ~w1916 & w9302;
assign w9304 = w9300 & w9303;
assign w9305 = ~w9036 & ~w9271;
assign w9306 = ~w9297 & w9305;
assign w9307 = w9304 & w9306;
assign w9308 = ~w9296 & w9307;
assign w9309 = ~pi036 & ~w9308;
assign w9310 = ~w9291 & ~w9309;
assign w9311 = w9282 & w9310;
assign w9312 = pi036 & ~w9258;
assign w9313 = w9311 & ~w9312;
assign w9314 = ~w9236 & w9313;
assign w9315 = w9236 & ~w9313;
assign w9316 = ~w9314 & ~w9315;
assign w9317 = ~w8716 & ~w9316;
assign w9318 = w8716 & w9316;
assign w9319 = ~w9317 & ~w9318;
assign w9320 = (~w2085 & w2100) | (~w2085 & w19012) | (w2100 & w19012);
assign w9321 = (~pi092 & w9320) | (~pi092 & w19013) | (w9320 & w19013);
assign w9322 = ~w5786 & ~w9095;
assign w9323 = pi092 & ~w9322;
assign w9324 = w2079 & w2095;
assign w9325 = ~w2086 & ~w8467;
assign w9326 = ~w8515 & ~w9324;
assign w9327 = w9325 & w9326;
assign w9328 = ~pi028 & w2164;
assign w9329 = w9327 & ~w9328;
assign w9330 = w9329 & w19014;
assign w9331 = pi028 & w2074;
assign w9332 = (pi092 & w9331) | (pi092 & w19015) | (w9331 & w19015);
assign w9333 = ~w5789 & ~w8489;
assign w9334 = ~w9332 & w9333;
assign w9335 = ~pi089 & ~w9334;
assign w9336 = ~w8503 & ~w9324;
assign w9337 = ~w5860 & w9336;
assign w9338 = w2095 & w2121;
assign w9339 = ~w2109 & ~w9338;
assign w9340 = ~pi092 & ~w9339;
assign w9341 = ~pi092 & w8458;
assign w9342 = ~pi053 & ~w2168;
assign w9343 = ~w9341 & w9342;
assign w9344 = ~w9340 & w9343;
assign w9345 = (pi092 & ~w9337) | (pi092 & w9506) | (~w9337 & w9506);
assign w9346 = w9344 & ~w9345;
assign w9347 = ~w9335 & w9346;
assign w9348 = pi089 & ~w9330;
assign w9349 = w9347 & ~w9348;
assign w9350 = w2059 & ~w2060;
assign w9351 = ~w2179 & ~w9350;
assign w9352 = ~pi087 & w2127;
assign w9353 = w9351 & ~w9352;
assign w9354 = (~pi089 & ~w9353) | (~pi089 & w19016) | (~w9353 & w19016);
assign w9355 = ~w2094 & ~w2097;
assign w9356 = ~w2152 & ~w5791;
assign w9357 = w9355 & w9356;
assign w9358 = ~w2080 & ~w8486;
assign w9359 = w2060 & ~w9358;
assign w9360 = ~pi092 & w2143;
assign w9361 = ~w8481 & ~w9360;
assign w9362 = pi053 & w9361;
assign w9363 = ~w9358 & w19017;
assign w9364 = w9362 & ~w9363;
assign w9365 = ~w2074 & ~w5803;
assign w9366 = (w2162 & ~w9365) | (w2162 & w19018) | (~w9365 & w19018);
assign w9367 = (~pi092 & w2084) | (~pi092 & w19019) | (w2084 & w19019);
assign w9368 = ~w9366 & ~w9367;
assign w9369 = w9364 & w9368;
assign w9370 = pi089 & ~w9357;
assign w9371 = w9369 & w19020;
assign w9372 = ~w9349 & ~w9371;
assign w9373 = (w2060 & ~w8477) | (w2060 & w19021) | (~w8477 & w19021);
assign w9374 = w5848 & w8392;
assign w9375 = ~w2090 & ~w9374;
assign w9376 = ~w9373 & w9375;
assign w9377 = ~pi089 & ~w9376;
assign w9378 = ~pi028 & w2107;
assign w9379 = w2107 & w2077;
assign w9380 = ~w8396 & w19022;
assign w9381 = w8526 & ~w9380;
assign w9382 = w2085 & w5790;
assign w9383 = ~w9341 & ~w9382;
assign w9384 = w2059 & w19023;
assign w9385 = (pi089 & ~w9383) | (pi089 & w19024) | (~w9383 & w19024);
assign w9386 = w5864 & w20827;
assign w9387 = w2052 & w5824;
assign w9388 = ~w5853 & ~w9387;
assign w9389 = ~w9381 & ~w9385;
assign w9390 = ~w9386 & w9388;
assign w9391 = w9389 & w9390;
assign w9392 = ~w9377 & w9391;
assign w9393 = ~w9372 & w9392;
assign w9394 = ~w9372 & w19025;
assign w9395 = (pi178 & w9372) | (pi178 & w19026) | (w9372 & w19026);
assign w9396 = ~w9394 & ~w9395;
assign w9397 = ~w8899 & w9396;
assign w9398 = w8899 & ~w9396;
assign w9399 = ~w9397 & ~w9398;
assign w9400 = (~pi529 & ~w9319) | (~pi529 & w19027) | (~w9319 & w19027);
assign w9401 = ~w9319 & w9399;
assign w9402 = w9400 & ~w9401;
assign w9403 = ~pi178 & pi450;
assign w9404 = pi529 & ~w9403;
assign w9405 = pi178 & ~pi450;
assign w9406 = w9404 & ~w9405;
assign w9407 = ~w9402 & ~w9406;
assign w9408 = w1548 & w1657;
assign w9409 = (~w1927 & w9408) | (~w1927 & w19028) | (w9408 & w19028);
assign w9410 = (~pi002 & w9409) | (~pi002 & w19029) | (w9409 & w19029);
assign w9411 = ~w1872 & ~w8643;
assign w9412 = w1588 & ~w9411;
assign w9413 = (w1927 & w1679) | (w1927 & w19030) | (w1679 & w19030);
assign w9414 = pi032 & w1559;
assign w9415 = ~w1568 & ~w9414;
assign w9416 = w9051 & ~w9415;
assign w9417 = ~w9413 & ~w9416;
assign w9418 = ~w1662 & ~w1905;
assign w9419 = ~w9412 & w9418;
assign w9420 = w9417 & w9419;
assign w9421 = w1548 & w1552;
assign w9422 = ~w1659 & ~w9245;
assign w9423 = (w9244 & ~w9422) | (w9244 & w19031) | (~w9422 & w19031);
assign w9424 = ~w1854 & ~w8694;
assign w9425 = ~pi117 & ~w9424;
assign w9426 = (pi002 & w9249) | (pi002 & w19032) | (w9249 & w19032);
assign w9427 = ~w9423 & ~w9425;
assign w9428 = w9420 & w9427;
assign w9429 = (~pi036 & ~w9428) | (~pi036 & w20828) | (~w9428 & w20828);
assign w9430 = ~w1666 & ~w9019;
assign w9431 = (pi117 & ~w9008) | (pi117 & w19034) | (~w9008 & w19034);
assign w9432 = w9430 & ~w9431;
assign w9433 = w1659 & w1677;
assign w9434 = ~w1652 & ~w1855;
assign w9435 = ~w9433 & w9434;
assign w9436 = ~w1625 & w8688;
assign w9437 = ~w1583 & ~w8695;
assign w9438 = w8632 & ~w9437;
assign w9439 = ~w1560 & ~w1583;
assign w9440 = ~w1652 & ~w1872;
assign w9441 = w9439 & w9440;
assign w9442 = ~pi117 & ~w9441;
assign w9443 = ~w9438 & ~w9442;
assign w9444 = (~pi002 & ~w9435) | (~pi002 & w19035) | (~w9435 & w19035);
assign w9445 = w9443 & ~w9444;
assign w9446 = (pi036 & ~w9445) | (pi036 & w19036) | (~w9445 & w19036);
assign w9447 = ~w1556 & ~w1859;
assign w9448 = ~w8623 & w9447;
assign w9449 = ~pi117 & ~w9448;
assign w9450 = ~w1856 & ~w8689;
assign w9451 = (~pi002 & w9449) | (~pi002 & w19037) | (w9449 & w19037);
assign w9452 = w1554 & w1677;
assign w9453 = ~w1581 & ~w1674;
assign w9454 = ~w8685 & ~w9452;
assign w9455 = w9453 & w9454;
assign w9456 = (w9244 & ~w9455) | (w9244 & w19038) | (~w9455 & w19038);
assign w9457 = ~w1616 & ~w1666;
assign w9458 = pi067 & ~w9457;
assign w9459 = (w9051 & w9458) | (w9051 & w19039) | (w9458 & w19039);
assign w9460 = w1621 & w1634;
assign w9461 = ~w1662 & ~w9460;
assign w9462 = ~w9035 & w9461;
assign w9463 = w1588 & ~w9462;
assign w9464 = ~w1581 & ~w8618;
assign w9465 = w1577 & ~w9464;
assign w9466 = ~w9456 & ~w9459;
assign w9467 = ~w9463 & ~w9465;
assign w9468 = w9466 & w9467;
assign w9469 = ~w9451 & w9468;
assign w9470 = ~w9446 & w9469;
assign w9471 = ~w9429 & w9470;
assign w9472 = ~w1841 & w9471;
assign w9473 = w1841 & ~w9471;
assign w9474 = ~w9472 & ~w9473;
assign w9475 = w5881 & w9474;
assign w9476 = ~w5881 & ~w9474;
assign w9477 = ~w9475 & ~w9476;
assign w9478 = ~w8431 & w19040;
assign w9479 = (pi281 & w8431) | (pi281 & w19041) | (w8431 & w19041);
assign w9480 = ~w9478 & ~w9479;
assign w9481 = ~w2198 & w2431;
assign w9482 = w2198 & ~w2431;
assign w9483 = ~w9481 & ~w9482;
assign w9484 = w9480 & w9483;
assign w9485 = ~w9480 & ~w9483;
assign w9486 = ~w9484 & ~w9485;
assign w9487 = ~w9477 & w9486;
assign w9488 = ~pi529 & ~w9487;
assign w9489 = w9477 & ~w9486;
assign w9490 = w9488 & ~w9489;
assign w9491 = pi281 & pi426;
assign w9492 = pi529 & ~w9491;
assign w9493 = ~pi281 & ~pi426;
assign w9494 = w9492 & ~w9493;
assign w9495 = ~w9490 & ~w9494;
assign w9496 = ~pi092 & ~w2090;
assign w9497 = ~w5847 & w9076;
assign w9498 = ~w9496 & ~w9497;
assign w9499 = ~w2057 & ~w2166;
assign w9500 = ~w5792 & w9499;
assign w9501 = ~w5820 & ~w9360;
assign w9502 = w9500 & w9501;
assign w9503 = (~pi089 & ~w9502) | (~pi089 & w19042) | (~w9502 & w19042);
assign w9504 = ~w2092 & ~w8413;
assign w9505 = w8404 & ~w9504;
assign w9506 = w2085 & w19043;
assign w9507 = ~w5856 & ~w9506;
assign w9508 = ~w9505 & w9507;
assign w9509 = (w2187 & w8394) | (w2187 & w19044) | (w8394 & w19044);
assign w9510 = ~w2061 & ~w5845;
assign w9511 = ~w5849 & w9510;
assign w9512 = ~w9509 & w9511;
assign w9513 = ~w9503 & w9512;
assign w9514 = (pi053 & ~w9513) | (pi053 & w19045) | (~w9513 & w19045);
assign w9515 = ~w8414 & ~w9087;
assign w9516 = pi092 & w9515;
assign w9517 = ~w2110 & ~w8486;
assign w9518 = w8377 & w9517;
assign w9519 = ~w9516 & ~w9518;
assign w9520 = (pi089 & w9519) | (pi089 & w19046) | (w9519 & w19046);
assign w9521 = (pi085 & w2064) | (pi085 & w19047) | (w2064 & w19047);
assign w9522 = w2126 & w2138;
assign w9523 = ~w2178 & ~w9522;
assign w9524 = ~pi089 & ~w9523;
assign w9525 = ~w9386 & ~w9524;
assign w9526 = ~w9521 & w9525;
assign w9527 = ~w9520 & w9526;
assign w9528 = ~pi053 & ~w9527;
assign w9529 = ~w8396 & w19048;
assign w9530 = ~pi046 & w2062;
assign w9531 = ~w2178 & ~w9530;
assign w9532 = ~w2058 & w9531;
assign w9533 = pi092 & ~w9532;
assign w9534 = w2096 & w5823;
assign w9535 = ~w2158 & ~w5799;
assign w9536 = ~w9534 & w9535;
assign w9537 = ~w9533 & w9536;
assign w9538 = (~pi089 & ~w9537) | (~pi089 & w19049) | (~w9537 & w19049);
assign w9539 = w2075 & w2092;
assign w9540 = ~w8467 & ~w9539;
assign w9541 = (pi089 & w8467) | (pi089 & w2162) | (w8467 & w2162);
assign w9542 = (w9541 & ~w2113) | (w9541 & w20829) | (~w2113 & w20829);
assign w9543 = w2049 & w5790;
assign w9544 = ~w2143 & ~w9378;
assign w9545 = ~w9543 & w9544;
assign w9546 = w2172 & ~w9545;
assign w9547 = (pi092 & w5849) | (pi092 & w19050) | (w5849 & w19050);
assign w9548 = ~w9546 & ~w9547;
assign w9549 = w9548 & w20830;
assign w9550 = ~w9538 & w9549;
assign w9551 = w9550 & w19051;
assign w9552 = ~w8456 & w9551;
assign w9553 = w8456 & ~w9551;
assign w9554 = ~w9552 & ~w9553;
assign w9555 = w9072 & w9554;
assign w9556 = ~w9072 & ~w9554;
assign w9557 = ~w9555 & ~w9556;
assign w9558 = ~w2307 & ~w2325;
assign w9559 = w5736 & w9558;
assign w9560 = ~w8867 & ~w9559;
assign w9561 = ~w8741 & ~w8837;
assign w9562 = w9560 & w9561;
assign w9563 = ~w5689 & ~w8799;
assign w9564 = (pi080 & ~w2329) | (pi080 & w8750) | (~w2329 & w8750);
assign w9565 = pi073 & ~w9564;
assign w9566 = ~w8753 & w19052;
assign w9567 = w9565 & ~w9566;
assign w9568 = ~w2292 & ~w2375;
assign w9569 = (w2421 & ~w9568) | (w2421 & w19053) | (~w9568 & w19053);
assign w9570 = w2314 & w2337;
assign w9571 = ~pi071 & w9570;
assign w9572 = ~w2301 & ~w5757;
assign w9573 = (pi015 & ~w9570) | (pi015 & w19054) | (~w9570 & w19054);
assign w9574 = w9572 & w9573;
assign w9575 = ~w9569 & w9574;
assign w9576 = ~w9567 & w9575;
assign w9577 = (~pi073 & ~w9562) | (~pi073 & w19055) | (~w9562 & w19055);
assign w9578 = w9576 & ~w9577;
assign w9579 = ~w5736 & ~w8892;
assign w9580 = pi080 & w9579;
assign w9581 = w8817 & w19056;
assign w9582 = ~w9580 & ~w9581;
assign w9583 = (pi073 & w9582) | (pi073 & w18516) | (w9582 & w18516);
assign w9584 = ~pi015 & ~w2348;
assign w9585 = w5726 & w19057;
assign w9586 = w9584 & ~w9585;
assign w9587 = w5716 & w19058;
assign w9588 = w2333 & w2342;
assign w9589 = ~w5748 & ~w9588;
assign w9590 = ~pi073 & ~w9589;
assign w9591 = ~w9587 & ~w9590;
assign w9592 = w9586 & w9591;
assign w9593 = ~w9583 & w9592;
assign w9594 = ~pi110 & w5715;
assign w9595 = (w2290 & w9594) | (w2290 & w19059) | (w9594 & w19059);
assign w9596 = (pi080 & ~w2337) | (pi080 & w18932) | (~w2337 & w18932);
assign w9597 = (~pi080 & ~w2315) | (~pi080 & w18941) | (~w2315 & w18941);
assign w9598 = w2362 & w9597;
assign w9599 = (~w9598 & w20831) | (~w9598 & w20832) | (w20831 & w20832);
assign w9600 = (pi079 & w2343) | (pi079 & w19061) | (w2343 & w19061);
assign w9601 = (pi080 & w9600) | (pi080 & w19062) | (w9600 & w19062);
assign w9602 = w2302 & w2314;
assign w9603 = ~w8866 & ~w9602;
assign w9604 = ~w5688 & w9603;
assign w9605 = ~pi080 & ~w9604;
assign w9606 = w2316 & w2302;
assign w9607 = w2314 & w2357;
assign w9608 = w2345 & w5766;
assign w9609 = ~w9606 & ~w9607;
assign w9610 = ~w9608 & w9609;
assign w9611 = ~w9605 & w19063;
assign w9612 = ~pi073 & ~w9611;
assign w9613 = w5683 & w8866;
assign w9614 = ~w5711 & ~w9613;
assign w9615 = ~w8792 & w9614;
assign w9616 = ~w9612 & w20833;
assign w9617 = ~w9578 & ~w9593;
assign w9618 = w9616 & ~w9617;
assign w9619 = ~pi172 & w9618;
assign w9620 = pi172 & ~w9618;
assign w9621 = ~w9619 & ~w9620;
assign w9622 = w8812 & w9621;
assign w9623 = ~w8812 & ~w9621;
assign w9624 = ~w9622 & ~w9623;
assign w9625 = (~pi529 & ~w9624) | (~pi529 & w19064) | (~w9624 & w19064);
assign w9626 = ~w9557 & ~w9624;
assign w9627 = w9625 & ~w9626;
assign w9628 = ~pi172 & pi484;
assign w9629 = pi529 & ~w9628;
assign w9630 = pi172 & ~pi484;
assign w9631 = w9629 & ~w9630;
assign w9632 = ~w9627 & ~w9631;
assign w9633 = w2293 & w2325;
assign w9634 = ~w2336 & ~w5722;
assign w9635 = (pi080 & ~w9634) | (pi080 & w19065) | (~w9634 & w19065);
assign w9636 = pi071 & ~w2314;
assign w9637 = w5715 & ~w9636;
assign w9638 = w2345 & w2422;
assign w9639 = ~w5689 & ~w9638;
assign w9640 = ~w9637 & w9639;
assign w9641 = (~pi073 & ~w9640) | (~pi073 & w19066) | (~w9640 & w19066);
assign w9642 = ~w2335 & ~w2394;
assign w9643 = ~w8745 & ~w9607;
assign w9644 = w9642 & w9643;
assign w9645 = ~w5701 & ~w5727;
assign w9646 = ~pi080 & w9645;
assign w9647 = (~w9646 & ~w9644) | (~w9646 & w19067) | (~w9644 & w19067);
assign w9648 = (pi073 & w5696) | (pi073 & w19068) | (w5696 & w19068);
assign w9649 = ~w5726 & ~w9594;
assign w9650 = ~w9648 & w9649;
assign w9651 = ~pi080 & ~w9650;
assign w9652 = pi073 & w2292;
assign w9653 = ~w8833 & ~w9652;
assign w9654 = ~w2300 & w9653;
assign w9655 = ~w9651 & w9654;
assign w9656 = ~w9641 & ~w9647;
assign w9657 = (pi015 & ~w9656) | (pi015 & w19069) | (~w9656 & w19069);
assign w9658 = (pi080 & w9571) | (pi080 & w19070) | (w9571 & w19070);
assign w9659 = ~w2306 & w5709;
assign w9660 = ~w5757 & ~w9659;
assign w9661 = w5766 & w19071;
assign w9662 = w5738 & w9588;
assign w9663 = ~w9661 & ~w9662;
assign w9664 = ~pi080 & ~w9660;
assign w9665 = ~w9664 & w19072;
assign w9666 = ~pi073 & ~w9665;
assign w9667 = ~pi079 & ~w5764;
assign w9668 = w8880 & ~w9667;
assign w9669 = ~w2302 & w2329;
assign w9670 = pi073 & ~w9669;
assign w9671 = w2294 & w5693;
assign w9672 = w9670 & ~w9671;
assign w9673 = w2293 & w2302;
assign w9674 = pi080 & w5687;
assign w9675 = ~w9673 & ~w9674;
assign w9676 = w9672 & w9675;
assign w9677 = ~w9668 & ~w9676;
assign w9678 = w2316 & w2337;
assign w9679 = ~w8746 & ~w9678;
assign w9680 = ~pi080 & ~w9679;
assign w9681 = ~w2320 & ~w8723;
assign w9682 = w2415 & ~w9681;
assign w9683 = ~w8860 & ~w8866;
assign w9684 = w2421 & ~w9683;
assign w9685 = ~w9680 & ~w9682;
assign w9686 = ~w2349 & ~w9684;
assign w9687 = w9685 & w9686;
assign w9688 = ~w9677 & w9687;
assign w9689 = ~pi015 & ~w9688;
assign w9690 = ~pi080 & ~w5748;
assign w9691 = ~w8733 & ~w9690;
assign w9692 = ~w5684 & ~w8828;
assign w9693 = ~w9691 & w9692;
assign w9694 = w2342 & w2347;
assign w9695 = w5714 & w19073;
assign w9696 = pi042 & w9694;
assign w9697 = ~w9695 & ~w9696;
assign w9698 = (pi073 & ~w9693) | (pi073 & w19074) | (~w9693 & w19074);
assign w9699 = w9697 & ~w9698;
assign w9700 = ~w9689 & w19075;
assign w9701 = ~w9657 & w9700;
assign w9702 = w9700 & w19076;
assign w9703 = (pi162 & ~w9700) | (pi162 & w19077) | (~w9700 & w19077);
assign w9704 = ~w9702 & ~w9703;
assign w9705 = w1844 & ~w5881;
assign w9706 = ~w1844 & w5881;
assign w9707 = ~w9705 & ~w9706;
assign w9708 = (~pi529 & w9707) | (~pi529 & w19078) | (w9707 & w19078);
assign w9709 = ~w9704 & w9707;
assign w9710 = w9708 & ~w9709;
assign w9711 = pi162 & pi485;
assign w9712 = pi529 & ~w9711;
assign w9713 = ~pi162 & ~pi485;
assign w9714 = w9712 & ~w9713;
assign w9715 = ~w9710 & ~w9714;
assign w9716 = ~w9148 & ~w9316;
assign w9717 = w9148 & w9316;
assign w9718 = ~w9716 & ~w9717;
assign w9719 = ~w5765 & ~w8788;
assign w9720 = (~w2367 & w9719) | (~w2367 & w19079) | (w9719 & w19079);
assign w9721 = ~pi080 & ~w9720;
assign w9722 = ~w2393 & ~w5722;
assign w9723 = pi080 & ~w9722;
assign w9724 = w2347 & w2376;
assign w9725 = ~w2295 & ~w2330;
assign w9726 = ~w2369 & ~w9724;
assign w9727 = w9725 & w9726;
assign w9728 = ~w9723 & w9727;
assign w9729 = ~w5761 & w9728;
assign w9730 = ~w5716 & ~w5736;
assign w9731 = w2307 & ~w9730;
assign w9732 = w5756 & ~w9731;
assign w9733 = ~pi073 & ~w9732;
assign w9734 = ~w8777 & ~w8827;
assign w9735 = ~w9724 & w9734;
assign w9736 = (pi080 & ~w9735) | (pi080 & w19080) | (~w9735 & w19080);
assign w9737 = ~pi080 & w2348;
assign w9738 = ~w2405 & ~w9737;
assign w9739 = w2291 & w2328;
assign w9740 = ~w2358 & ~w9739;
assign w9741 = ~pi080 & ~w9740;
assign w9742 = w9738 & ~w9741;
assign w9743 = ~w9733 & w19081;
assign w9744 = (pi073 & ~w9729) | (pi073 & w20834) | (~w9729 & w20834);
assign w9745 = ~w5683 & w5714;
assign w9746 = ~w8791 & ~w9745;
assign w9747 = (~pi073 & ~w2382) | (~pi073 & w19082) | (~w2382 & w19082);
assign w9748 = ~w8863 & w9746;
assign w9749 = w9747 & w9748;
assign w9750 = w2314 & w5715;
assign w9751 = pi073 & ~w9750;
assign w9752 = ~w2335 & ~w2396;
assign w9753 = ~w8745 & w9751;
assign w9754 = w9752 & w9753;
assign w9755 = ~w9749 & ~w9754;
assign w9756 = pi075 & w8756;
assign w9757 = ~w2317 & ~w8785;
assign w9758 = (w2403 & ~w9757) | (w2403 & w19083) | (~w9757 & w19083);
assign w9759 = (~pi080 & w2327) | (~pi080 & w19084) | (w2327 & w19084);
assign w9760 = ~w2370 & ~w5701;
assign w9761 = w5683 & ~w9760;
assign w9762 = ~w8753 & ~w8867;
assign w9763 = ~w9761 & w9762;
assign w9764 = w9763 & w19085;
assign w9765 = (pi015 & w9755) | (pi015 & w19086) | (w9755 & w19086);
assign w9766 = w2321 & w2337;
assign w9767 = ~w9633 & ~w9766;
assign w9768 = ~w5688 & w9767;
assign w9769 = ~pi080 & ~w9768;
assign w9770 = (w8847 & ~w8751) | (w8847 & w19087) | (~w8751 & w19087);
assign w9771 = w2421 & w5765;
assign w9772 = ~w2350 & ~w9771;
assign w9773 = ~w9769 & w19088;
assign w9774 = ~pi073 & ~w9773;
assign w9775 = (~w2337 & w9737) | (~w2337 & w19089) | (w9737 & w19089);
assign w9776 = ~w9587 & ~w9661;
assign w9777 = ~w8740 & w9776;
assign w9778 = (pi073 & w9775) | (pi073 & w19090) | (w9775 & w19090);
assign w9779 = w9777 & ~w9778;
assign w9780 = ~w9774 & w9779;
assign w9781 = ~w9765 & w9780;
assign w9782 = (~pi015 & w9744) | (~pi015 & w19091) | (w9744 & w19091);
assign w9783 = w9781 & ~w9782;
assign w9784 = ~pi226 & w9783;
assign w9785 = pi226 & ~w9783;
assign w9786 = ~w9784 & ~w9785;
assign w9787 = ~w8899 & w9786;
assign w9788 = w8899 & ~w9786;
assign w9789 = ~w9787 & ~w9788;
assign w9790 = (~pi529 & ~w9718) | (~pi529 & w19092) | (~w9718 & w19092);
assign w9791 = ~w9718 & w9789;
assign w9792 = w9790 & ~w9791;
assign w9793 = ~pi226 & pi445;
assign w9794 = pi529 & ~w9793;
assign w9795 = pi226 & ~pi445;
assign w9796 = w9794 & ~w9795;
assign w9797 = ~w9792 & ~w9796;
assign w9798 = w9700 & w19093;
assign w9799 = (pi192 & ~w9700) | (pi192 & w19094) | (~w9700 & w19094);
assign w9800 = ~w9798 & ~w9799;
assign w9801 = ~w1841 & w8456;
assign w9802 = w1841 & ~w8456;
assign w9803 = ~w9801 & ~w9802;
assign w9804 = ~w1936 & w5878;
assign w9805 = w1936 & ~w5878;
assign w9806 = ~w9804 & ~w9805;
assign w9807 = w9803 & w9806;
assign w9808 = ~w9803 & ~w9806;
assign w9809 = ~w9807 & ~w9808;
assign w9810 = (~pi529 & w9809) | (~pi529 & w19095) | (w9809 & w19095);
assign w9811 = ~w9800 & w9809;
assign w9812 = w9810 & ~w9811;
assign w9813 = ~pi192 & pi453;
assign w9814 = pi529 & ~w9813;
assign w9815 = pi192 & ~pi453;
assign w9816 = w9814 & ~w9815;
assign w9817 = ~w9812 & ~w9816;
assign w9818 = ~pi016 & w5923;
assign w9819 = (~pi120 & w9818) | (~pi120 & w19096) | (w9818 & w19096);
assign w9820 = w2464 & w2526;
assign w9821 = ~w5986 & ~w9820;
assign w9822 = ~w9819 & w9821;
assign w9823 = ~pi003 & ~w9822;
assign w9824 = (w5996 & w5949) | (w5996 & w19097) | (w5949 & w19097);
assign w9825 = ~w2776 & ~w5918;
assign w9826 = w2805 & ~w9825;
assign w9827 = ~w2564 & ~w2819;
assign w9828 = (pi003 & ~w9827) | (pi003 & w19098) | (~w9827 & w19098);
assign w9829 = (w2828 & w2536) | (w2828 & w19099) | (w2536 & w19099);
assign w9830 = ~w2764 & ~w9820;
assign w9831 = ~pi120 & ~w9830;
assign w9832 = pi003 & ~pi120;
assign w9833 = w2448 & w2476;
assign w9834 = ~w2766 & ~w9833;
assign w9835 = ~pi074 & w2522;
assign w9836 = (w9832 & ~w9834) | (w9832 & w19100) | (~w9834 & w19100);
assign w9837 = ~w9831 & ~w9836;
assign w9838 = ~w2823 & ~w9829;
assign w9839 = ~w5925 & w9838;
assign w9840 = w9837 & w9839;
assign w9841 = ~w9824 & ~w9826;
assign w9842 = ~w9828 & w9841;
assign w9843 = w9840 & w19101;
assign w9844 = ~pi044 & ~w9843;
assign w9845 = ~w2518 & ~w2796;
assign w9846 = pi081 & ~w9845;
assign w9847 = ~pi016 & w2459;
assign w9848 = pi045 & w2541;
assign w9849 = ~w2565 & ~w9848;
assign w9850 = ~pi016 & ~pi120;
assign w9851 = ~pi074 & ~w9850;
assign w9852 = ~w2546 & ~w5923;
assign w9853 = w9851 & ~w9852;
assign w9854 = (pi003 & w9848) | (pi003 & w19102) | (w9848 & w19102);
assign w9855 = ~w9853 & ~w9854;
assign w9856 = (w5996 & w9846) | (w5996 & w19103) | (w9846 & w19103);
assign w9857 = w9855 & ~w9856;
assign w9858 = ~pi016 & pi120;
assign w9859 = ~w2569 & ~w2762;
assign w9860 = w2523 & ~w9858;
assign w9861 = w9859 & ~w9860;
assign w9862 = ~w2546 & ~w2569;
assign w9863 = w9862 & w19104;
assign w9864 = ~pi120 & ~w9863;
assign w9865 = (~pi003 & ~w9861) | (~pi003 & w19105) | (~w9861 & w19105);
assign w9866 = ~w9864 & ~w9865;
assign w9867 = w9857 & w9866;
assign w9868 = pi044 & ~w9867;
assign w9869 = ~w2512 & ~w2533;
assign w9870 = ~w5993 & w9869;
assign w9871 = ~pi120 & ~w9870;
assign w9872 = ~w2763 & ~w5926;
assign w9873 = (~pi003 & w9871) | (~pi003 & w19106) | (w9871 & w19106);
assign w9874 = ~w2521 & ~w5983;
assign w9875 = (w5996 & ~w9874) | (w5996 & w19107) | (~w9874 & w19107);
assign w9876 = w2478 & w18205;
assign w9877 = ~w2547 & ~w2577;
assign w9878 = ~w9876 & w9877;
assign w9879 = w2522 & w2748;
assign w9880 = ~w5925 & ~w9879;
assign w9881 = ~w5965 & w9880;
assign w9882 = w2805 & ~w9881;
assign w9883 = ~w9832 & ~w9858;
assign w9884 = w2584 & ~w9883;
assign w9885 = ~w5987 & ~w9884;
assign w9886 = ~w9882 & w9885;
assign w9887 = (w9832 & ~w9878) | (w9832 & w19108) | (~w9878 & w19108);
assign w9888 = w9886 & ~w9887;
assign w9889 = w9888 & w19109;
assign w9890 = ~w9868 & w9889;
assign w9891 = ~w9844 & w9890;
assign w9892 = ~w2744 & w9891;
assign w9893 = w2744 & ~w9891;
assign w9894 = ~w9892 & ~w9893;
assign w9895 = w6627 & w9894;
assign w9896 = ~w6627 & ~w9894;
assign w9897 = ~w9895 & ~w9896;
assign w9898 = ~w6235 & w19110;
assign w9899 = (pi278 & w6235) | (pi278 & w19111) | (w6235 & w19111);
assign w9900 = ~w9898 & ~w9899;
assign w9901 = ~w3102 & w3353;
assign w9902 = w3102 & ~w3353;
assign w9903 = ~w9901 & ~w9902;
assign w9904 = w9900 & w9903;
assign w9905 = ~w9900 & ~w9903;
assign w9906 = ~w9904 & ~w9905;
assign w9907 = ~w9897 & w9906;
assign w9908 = ~pi529 & ~w9907;
assign w9909 = w9897 & ~w9906;
assign w9910 = w9908 & ~w9909;
assign w9911 = pi278 & pi513;
assign w9912 = pi529 & ~w9911;
assign w9913 = ~pi278 & ~pi513;
assign w9914 = w9912 & ~w9913;
assign w9915 = ~w9910 & ~w9914;
assign w9916 = ~w3199 & w9891;
assign w9917 = w3199 & ~w9891;
assign w9918 = ~w9916 & ~w9917;
assign w9919 = w6954 & ~w9918;
assign w9920 = ~w6954 & w9918;
assign w9921 = ~w9919 & ~w9920;
assign w9922 = ~w6367 & w6948;
assign w9923 = w6367 & ~w6948;
assign w9924 = ~w9922 & ~w9923;
assign w9925 = ~pi280 & w3353;
assign w9926 = pi280 & ~w3353;
assign w9927 = ~w9925 & ~w9926;
assign w9928 = w9924 & w9927;
assign w9929 = ~w9924 & ~w9927;
assign w9930 = ~w9928 & ~w9929;
assign w9931 = ~w9921 & ~w9930;
assign w9932 = ~pi529 & ~w9931;
assign w9933 = w9921 & w9930;
assign w9934 = w9932 & ~w9933;
assign w9935 = pi280 & pi470;
assign w9936 = pi529 & ~w9935;
assign w9937 = ~pi280 & ~pi470;
assign w9938 = w9936 & ~w9937;
assign w9939 = ~w9934 & ~w9938;
assign w9940 = ~w2518 & w2522;
assign w9941 = ~w2465 & w9940;
assign w9942 = pi003 & w9941;
assign w9943 = (~pi120 & w9942) | (~pi120 & w19112) | (w9942 & w19112);
assign w9944 = w2464 & w2478;
assign w9945 = w2457 & w5938;
assign w9946 = pi041 & w2468;
assign w9947 = ~w2537 & ~w9946;
assign w9948 = ~w9944 & ~w9945;
assign w9949 = ~pi003 & w9948;
assign w9950 = w9947 & w9949;
assign w9951 = w2459 & w2469;
assign w9952 = ~w2775 & ~w9951;
assign w9953 = pi120 & ~w9952;
assign w9954 = pi003 & ~w2477;
assign w9955 = ~w9953 & w9954;
assign w9956 = ~w9950 & ~w9955;
assign w9957 = w2448 & w2460;
assign w9958 = (pi120 & w2580) | (pi120 & w19113) | (w2580 & w19113);
assign w9959 = ~pi044 & ~w2812;
assign w9960 = ~w9958 & w9959;
assign w9961 = ~w2559 & ~w5974;
assign w9962 = ~pi120 & ~w9961;
assign w9963 = w2522 & w9858;
assign w9964 = ~w2837 & ~w5993;
assign w9965 = pi003 & ~w9963;
assign w9966 = w9964 & w9965;
assign w9967 = w2475 & w2796;
assign w9968 = w2532 & ~w9851;
assign w9969 = ~w5977 & ~w9968;
assign w9970 = ~pi003 & ~w9967;
assign w9971 = ~w2792 & w9970;
assign w9972 = w9969 & w9971;
assign w9973 = ~w9962 & w9966;
assign w9974 = ~w9972 & ~w9973;
assign w9975 = ~pi045 & w2469;
assign w9976 = ~w2777 & ~w9975;
assign w9977 = pi120 & ~w2570;
assign w9978 = ~w5926 & w9976;
assign w9979 = w9977 & w9978;
assign w9980 = ~pi120 & ~w5918;
assign w9981 = ~w2834 & w9980;
assign w9982 = ~w2819 & w9981;
assign w9983 = ~w9979 & ~w9982;
assign w9984 = pi044 & ~w9983;
assign w9985 = ~w9974 & w9984;
assign w9986 = ~w9956 & w19114;
assign w9987 = ~w9985 & ~w9986;
assign w9988 = ~w2817 & ~w5926;
assign w9989 = ~w2466 & ~w2564;
assign w9990 = w9988 & w19115;
assign w9991 = pi120 & ~w9990;
assign w9992 = ~w2510 & ~w5923;
assign w9993 = ~w9820 & w9992;
assign w9994 = ~pi120 & ~w9993;
assign w9995 = w2831 & w9850;
assign w9996 = (pi074 & w9995) | (pi074 & w19116) | (w9995 & w19116);
assign w9997 = ~w2542 & ~w2812;
assign w9998 = ~pi003 & w9997;
assign w9999 = ~w9996 & w9998;
assign w10000 = ~w9994 & w9999;
assign w10001 = ~w9991 & w10000;
assign w10002 = ~w2478 & w5945;
assign w10003 = ~w2834 & ~w5949;
assign w10004 = (~pi120 & ~w10003) | (~pi120 & w19117) | (~w10003 & w19117);
assign w10005 = pi120 & w2447;
assign w10006 = w2499 & w2802;
assign w10007 = ~w2778 & ~w10006;
assign w10008 = w2469 & w10005;
assign w10009 = w10007 & ~w10008;
assign w10010 = (pi003 & ~w2485) | (pi003 & w19118) | (~w2485 & w19118);
assign w10011 = w10009 & w19119;
assign w10012 = ~w10004 & w10011;
assign w10013 = ~w10001 & ~w10012;
assign w10014 = ~w9987 & ~w10013;
assign w10015 = ~w6711 & w10014;
assign w10016 = w6711 & ~w10014;
assign w10017 = ~w10015 & ~w10016;
assign w10018 = w2599 & w2721;
assign w10019 = ~w2633 & ~w3168;
assign w10020 = (~pi118 & ~w10019) | (~pi118 & w19120) | (~w10019 & w19120);
assign w10021 = ~w2635 & ~w6677;
assign w10022 = pi118 & ~w10021;
assign w10023 = w2660 & w2713;
assign w10024 = ~w2711 & ~w3154;
assign w10025 = ~w6126 & ~w10023;
assign w10026 = w10024 & w10025;
assign w10027 = ~w10022 & w10026;
assign w10028 = w10027 & w19121;
assign w10029 = (w2719 & w3105) | (w2719 & w19122) | (w3105 & w19122);
assign w10030 = ~w2739 & ~w10023;
assign w10031 = ~w10029 & w10030;
assign w10032 = pi118 & ~w10031;
assign w10033 = w2648 & w2697;
assign w10034 = ~w6125 & ~w10033;
assign w10035 = ~pi066 & w2689;
assign w10036 = pi119 & w2854;
assign w10037 = ~w10035 & ~w10036;
assign w10038 = w10034 & w10037;
assign w10039 = ~pi034 & ~w10038;
assign w10040 = ~pi118 & w2865;
assign w10041 = ~w3174 & ~w10040;
assign w10042 = ~w2720 & ~w2736;
assign w10043 = ~pi118 & ~w10042;
assign w10044 = w10041 & ~w10043;
assign w10045 = ~w10039 & w19123;
assign w10046 = pi034 & ~w10028;
assign w10047 = w10045 & ~w10046;
assign w10048 = ~w2624 & ~w6662;
assign w10049 = ~w6108 & ~w10048;
assign w10050 = (~pi034 & ~w3105) | (~pi034 & w19124) | (~w3105 & w19124);
assign w10051 = ~w10049 & w10050;
assign w10052 = pi118 & ~w6652;
assign w10053 = w10051 & ~w10052;
assign w10054 = pi034 & ~w2856;
assign w10055 = ~w2863 & w10054;
assign w10056 = ~w2866 & ~w3164;
assign w10057 = w10055 & w10056;
assign w10058 = ~w10053 & ~w10057;
assign w10059 = pi103 & w2719;
assign w10060 = ~w2697 & ~w2918;
assign w10061 = (w3172 & ~w10060) | (w3172 & w19125) | (~w10060 & w19125);
assign w10062 = (~pi118 & w3110) | (~pi118 & w19126) | (w3110 & w19126);
assign w10063 = pi118 & w2632;
assign w10064 = w2664 & w2853;
assign w10065 = w3139 & w10063;
assign w10066 = ~w10064 & ~w10065;
assign w10067 = ~w2919 & ~w6158;
assign w10068 = w10066 & w10067;
assign w10069 = w10068 & w19127;
assign w10070 = (pi038 & w10058) | (pi038 & w19128) | (w10058 & w19128);
assign w10071 = (w10063 & w6117) | (w10063 & w10065) | (w6117 & w10065);
assign w10072 = w2661 & w6131;
assign w10073 = ~w3186 & ~w10072;
assign w10074 = ~w10071 & w10073;
assign w10075 = ~pi034 & ~w10074;
assign w10076 = ~w2627 & ~w2641;
assign w10077 = ~w2614 & ~w10076;
assign w10078 = w2625 & w2922;
assign w10079 = w3147 & w10078;
assign w10080 = w2853 & w6140;
assign w10081 = ~w3128 & ~w10080;
assign w10082 = w2600 & w19129;
assign w10083 = w10081 & w19130;
assign w10084 = pi034 & ~w2721;
assign w10085 = (w10084 & w10040) | (w10084 & w19131) | (w10040 & w19131);
assign w10086 = w10083 & ~w10085;
assign w10087 = (w6164 & w10077) | (w6164 & w19132) | (w10077 & w19132);
assign w10088 = w10086 & ~w10087;
assign w10089 = ~w10075 & w10088;
assign w10090 = ~w10070 & w10089;
assign w10091 = ~pi038 & ~w10047;
assign w10092 = w10090 & ~w10091;
assign w10093 = w2962 & w3006;
assign w10094 = pi011 & w2982;
assign w10095 = ~w3043 & ~w10094;
assign w10096 = (~pi116 & ~w10095) | (~pi116 & w19133) | (~w10095 & w19133);
assign w10097 = ~w6203 & ~w6737;
assign w10098 = pi116 & ~w10097;
assign w10099 = w2957 & w2984;
assign w10100 = w3042 & w6084;
assign w10101 = ~w2993 & ~w3040;
assign w10102 = ~w10099 & ~w10100;
assign w10103 = w10101 & w10102;
assign w10104 = ~w10098 & w10103;
assign w10105 = w10104 & w19134;
assign w10106 = w2980 & w2958;
assign w10107 = (pi116 & w10106) | (pi116 & w18629) | (w10106 & w18629);
assign w10108 = ~w6246 & ~w6713;
assign w10109 = ~w10107 & w10108;
assign w10110 = ~pi058 & ~w10109;
assign w10111 = (w3023 & w3084) | (w3023 & w19135) | (w3084 & w19135);
assign w10112 = ~w6009 & ~w10099;
assign w10113 = ~w10111 & w10112;
assign w10114 = pi116 & ~w10113;
assign w10115 = ~pi022 & w2950;
assign w10116 = w2950 & w2968;
assign w10117 = ~w2954 & ~w10116;
assign w10118 = ~pi116 & ~w10117;
assign w10119 = ~pi116 & w6051;
assign w10120 = ~w10119 & w19136;
assign w10121 = ~w10118 & w10120;
assign w10122 = ~w10114 & w10121;
assign w10123 = ~w10110 & w10122;
assign w10124 = pi058 & ~w10105;
assign w10125 = w10123 & ~w10124;
assign w10126 = ~pi022 & w3028;
assign w10127 = (~w2965 & w10126) | (~w2965 & w19137) | (w10126 & w19137);
assign w10128 = ~w3085 & ~w6776;
assign w10129 = (~pi058 & ~w10128) | (~pi058 & w19138) | (~w10128 & w19138);
assign w10130 = w2982 & w2958;
assign w10131 = ~w3053 & ~w10130;
assign w10132 = ~w2997 & ~w3059;
assign w10133 = w10131 & w10132;
assign w10134 = pi058 & ~w10133;
assign w10135 = w2976 & w6178;
assign w10136 = w3033 & w6744;
assign w10137 = w2965 & w3026;
assign w10138 = ~w10136 & ~w10137;
assign w10139 = ~w6022 & ~w10135;
assign w10140 = w10138 & w10139;
assign w10141 = pi060 & w10140;
assign w10142 = (~pi116 & w2991) | (~pi116 & w19139) | (w2991 & w19139);
assign w10143 = ~w2981 & ~w6765;
assign w10144 = (w3065 & ~w10143) | (w3065 & w19140) | (~w10143 & w19140);
assign w10145 = ~w10134 & w10141;
assign w10146 = ~w10142 & ~w10144;
assign w10147 = w10145 & w19141;
assign w10148 = ~w10125 & ~w10147;
assign w10149 = ~pi022 & w2962;
assign w10150 = ~w6033 & ~w10149;
assign w10151 = ~w3007 & ~w10135;
assign w10152 = w3003 & w3061;
assign w10153 = w10151 & ~w10152;
assign w10154 = w6178 & ~w10150;
assign w10155 = w10153 & ~w10154;
assign w10156 = ~pi058 & ~pi116;
assign w10157 = w6084 & w3031;
assign w10158 = ~w6067 & w19142;
assign w10159 = w10156 & ~w10158;
assign w10160 = (~pi116 & w6057) | (~pi116 & w18654) | (w6057 & w18654);
assign w10161 = w3023 & w6568;
assign w10162 = ~w10119 & ~w10161;
assign w10163 = w3052 & w3076;
assign w10164 = w3052 & w19143;
assign w10165 = ~w3005 & ~w10164;
assign w10166 = pi058 & ~w10162;
assign w10167 = w10165 & ~w10166;
assign w10168 = w10167 & w19144;
assign w10169 = ~pi058 & ~w10155;
assign w10170 = w10168 & ~w10169;
assign w10171 = ~w10148 & w10170;
assign w10172 = ~w10092 & w10171;
assign w10173 = w10092 & ~w10171;
assign w10174 = ~w10172 & ~w10173;
assign w10175 = ~w3289 & ~w3317;
assign w10176 = (~pi090 & ~w10175) | (~pi090 & w19145) | (~w10175 & w19145);
assign w10177 = ~w6316 & ~w6807;
assign w10178 = pi090 & ~w10177;
assign w10179 = w3258 & w3280;
assign w10180 = ~w3239 & ~w3285;
assign w10181 = ~w6401 & ~w10179;
assign w10182 = w10180 & w10181;
assign w10183 = ~w10178 & w10182;
assign w10184 = w10183 & w19146;
assign w10185 = w3214 & w6459;
assign w10186 = ~w6515 & ~w10185;
assign w10187 = ~pi086 & ~w10186;
assign w10188 = w3262 & w3263;
assign w10189 = ~w6403 & ~w10188;
assign w10190 = ~w10187 & w10189;
assign w10191 = ~pi088 & ~w10190;
assign w10192 = ~w6470 & ~w10179;
assign w10193 = ~w6844 & w10192;
assign w10194 = w3220 & w3264;
assign w10195 = (pi090 & ~w10193) | (pi090 & w19147) | (~w10193 & w19147);
assign w10196 = w3251 & w6816;
assign w10197 = ~w3324 & ~w10196;
assign w10198 = ~w3208 & ~w3212;
assign w10199 = ~pi090 & ~w10198;
assign w10200 = w10197 & ~w10199;
assign w10201 = ~w10191 & w19148;
assign w10202 = pi088 & ~w10184;
assign w10203 = w10201 & ~w10202;
assign w10204 = pi112 & w3229;
assign w10205 = ~w6808 & ~w10204;
assign w10206 = ~w3262 & w6283;
assign w10207 = ~pi090 & w3343;
assign w10208 = ~w10206 & ~w10207;
assign w10209 = (~pi088 & ~w3335) | (~pi088 & w19149) | (~w3335 & w19149);
assign w10210 = w10208 & w10209;
assign w10211 = pi090 & ~w10205;
assign w10212 = w10210 & ~w10211;
assign w10213 = pi088 & ~w6887;
assign w10214 = ~w3260 & w10213;
assign w10215 = ~w3311 & ~w6387;
assign w10216 = w10214 & w10215;
assign w10217 = ~w10212 & ~w10216;
assign w10218 = w3231 & ~w3233;
assign w10219 = ~w3275 & ~w6901;
assign w10220 = w3262 & ~w10219;
assign w10221 = ~pi090 & w6457;
assign w10222 = ~w6394 & ~w10221;
assign w10223 = ~w10220 & w10222;
assign w10224 = (~pi090 & w3241) | (~pi090 & w19150) | (w3241 & w19150);
assign w10225 = (w3321 & w10218) | (w3321 & w19151) | (w10218 & w19151);
assign w10226 = w10223 & w20835;
assign w10227 = (pi006 & w10217) | (pi006 & w20836) | (w10217 & w20836);
assign w10228 = ~w3229 & ~w6518;
assign w10229 = (~pi090 & w10228) | (~pi090 & w18594) | (w10228 & w18594);
assign w10230 = (w6817 & w6392) | (w6817 & w19152) | (w6392 & w19152);
assign w10231 = w3272 & w6288;
assign w10232 = ~w3249 & ~w10231;
assign w10233 = ~w10230 & w10232;
assign w10234 = ~w10229 & w10233;
assign w10235 = ~pi088 & ~w10234;
assign w10236 = ~pi090 & w3285;
assign w10237 = ~w6494 & ~w10236;
assign w10238 = w6399 & w19153;
assign w10239 = w10237 & w19154;
assign w10240 = pi088 & ~w3284;
assign w10241 = (w10240 & w10196) | (w10240 & w19155) | (w10196 & w19155);
assign w10242 = w10239 & ~w10241;
assign w10243 = ~w10235 & w10242;
assign w10244 = ~w10227 & w10243;
assign w10245 = ~pi006 & ~w10203;
assign w10246 = w10244 & ~w10245;
assign w10247 = w10244 & w19156;
assign w10248 = (pi141 & ~w10244) | (pi141 & w19157) | (~w10244 & w19157);
assign w10249 = ~w10247 & ~w10248;
assign w10250 = w10174 & w10249;
assign w10251 = ~w10174 & ~w10249;
assign w10252 = ~w10250 & ~w10251;
assign w10253 = (~pi529 & w10252) | (~pi529 & w19158) | (w10252 & w19158);
assign w10254 = ~w10017 & w10252;
assign w10255 = w10253 & ~w10254;
assign w10256 = ~pi141 & pi488;
assign w10257 = pi529 & ~w10256;
assign w10258 = pi141 & ~pi488;
assign w10259 = w10257 & ~w10258;
assign w10260 = ~w10255 & ~w10259;
assign w10261 = ~w2500 & ~w2791;
assign w10262 = pi120 & ~w10261;
assign w10263 = ~w5965 & ~w5978;
assign w10264 = ~w10262 & w10263;
assign w10265 = w2464 & w2522;
assign w10266 = ~w5993 & ~w10265;
assign w10267 = w2765 & w10266;
assign w10268 = pi003 & ~w10267;
assign w10269 = (~pi120 & ~w9827) | (~pi120 & w19159) | (~w9827 & w19159);
assign w10270 = pi016 & w2568;
assign w10271 = ~pi120 & w2520;
assign w10272 = w2526 & w2832;
assign w10273 = ~w10271 & ~w10272;
assign w10274 = ~w5937 & ~w5991;
assign w10275 = w10273 & w10274;
assign w10276 = (w9832 & ~w2767) | (w9832 & w19160) | (~w2767 & w19160);
assign w10277 = w10275 & ~w10276;
assign w10278 = ~w10268 & w10277;
assign w10279 = ~w10269 & w10278;
assign w10280 = w2447 & w2460;
assign w10281 = ~w2496 & ~w2523;
assign w10282 = (~pi120 & ~w10281) | (~pi120 & w19162) | (~w10281 & w19162);
assign w10283 = (w2821 & w2494) | (w2821 & w19163) | (w2494 & w19163);
assign w10284 = w2476 & w2532;
assign w10285 = ~w5950 & ~w10284;
assign w10286 = ~w2584 & ~w5923;
assign w10287 = ~w2578 & w10286;
assign w10288 = w10285 & w10287;
assign w10289 = w10288 & w19164;
assign w10290 = ~pi120 & w5954;
assign w10291 = w2568 & w2777;
assign w10292 = ~w10290 & ~w10291;
assign w10293 = w2775 & w2832;
assign w10294 = w2558 & w5955;
assign w10295 = ~pi120 & w5923;
assign w10296 = ~w10294 & ~w10295;
assign w10297 = ~w2823 & w10296;
assign w10298 = (pi003 & ~w10292) | (pi003 & w19165) | (~w10292 & w19165);
assign w10299 = w10297 & ~w10298;
assign w10300 = pi003 & ~pi044;
assign w10301 = ~w10289 & w10300;
assign w10302 = w10299 & ~w10301;
assign w10303 = ~w2559 & ~w2570;
assign w10304 = ~pi074 & ~w10303;
assign w10305 = w2536 & w2828;
assign w10306 = w2480 & w2801;
assign w10307 = ~w10305 & ~w10306;
assign w10308 = ~w10304 & w10307;
assign w10309 = ~pi003 & ~w10308;
assign w10310 = w2478 & w9858;
assign w10311 = ~w2833 & ~w10290;
assign w10312 = ~w2547 & ~w10310;
assign w10313 = w10311 & w10312;
assign w10314 = ~w2565 & ~w2579;
assign w10315 = ~w5917 & ~w5943;
assign w10316 = ~pi120 & ~w10314;
assign w10317 = w2499 & ~w10315;
assign w10318 = ~w10316 & ~w10317;
assign w10319 = w10313 & w10318;
assign w10320 = ~w10309 & w10319;
assign w10321 = ~pi044 & ~w10320;
assign w10322 = w2460 & w2532;
assign w10323 = ~w2542 & w19166;
assign w10324 = ~pi120 & ~w10323;
assign w10325 = (w2832 & ~w5939) | (w2832 & w10272) | (~w5939 & w10272);
assign w10326 = ~w2822 & ~w5925;
assign w10327 = ~w10325 & w10326;
assign w10328 = ~w10324 & w10327;
assign w10329 = ~pi003 & ~w10328;
assign w10330 = ~w10321 & ~w10329;
assign w10331 = w10302 & w10330;
assign w10332 = (pi044 & ~w10279) | (pi044 & w19167) | (~w10279 & w19167);
assign w10333 = w10331 & ~w10332;
assign w10334 = ~pi118 & ~w3177;
assign w10335 = (pi118 & ~w2599) | (pi118 & w19168) | (~w2599 & w19168);
assign w10336 = pi119 & w2660;
assign w10337 = w10335 & ~w10336;
assign w10338 = w10042 & w10334;
assign w10339 = ~w2600 & ~w6126;
assign w10340 = ~w3116 & w10339;
assign w10341 = pi118 & ~w10340;
assign w10342 = (pi034 & ~w3104) | (pi034 & w19169) | (~w3104 & w19169);
assign w10343 = w2864 & w10342;
assign w10344 = ~w10341 & w10343;
assign w10345 = ~pi034 & ~w2865;
assign w10346 = (w10345 & w10338) | (w10345 & w19170) | (w10338 & w19170);
assign w10347 = ~w10344 & ~w10346;
assign w10348 = w2931 & ~w3174;
assign w10349 = w6139 & w10348;
assign w10350 = ~w2633 & ~w3173;
assign w10351 = (pi038 & w10347) | (pi038 & w19171) | (w10347 & w19171);
assign w10352 = w2719 & w2721;
assign w10353 = ~w2714 & ~w10352;
assign w10354 = (pi034 & ~w2673) | (pi034 & w19172) | (~w2673 & w19172);
assign w10355 = ~pi103 & w2877;
assign w10356 = w10354 & ~w10355;
assign w10357 = pi118 & ~w10353;
assign w10358 = w10356 & ~w10357;
assign w10359 = ~w2716 & ~w2927;
assign w10360 = ~pi034 & ~w3173;
assign w10361 = w10359 & w10360;
assign w10362 = w2669 & w2721;
assign w10363 = ~w2665 & ~w6702;
assign w10364 = w10361 & w10363;
assign w10365 = ~w10362 & w10364;
assign w10366 = ~w2641 & ~w2697;
assign w10367 = w2609 & ~w10366;
assign w10368 = ~w2854 & ~w3118;
assign w10369 = ~w6124 & w10368;
assign w10370 = (~pi118 & ~w10369) | (~pi118 & w19173) | (~w10369 & w19173);
assign w10371 = ~w10358 & ~w10365;
assign w10372 = ~w2666 & ~w2670;
assign w10373 = ~pi118 & ~w2865;
assign w10374 = w10372 & w10373;
assign w10375 = ~w2731 & ~w6648;
assign w10376 = pi118 & w10375;
assign w10377 = ~w10374 & ~w10376;
assign w10378 = w2660 & w2669;
assign w10379 = ~w2722 & ~w10378;
assign w10380 = (~pi034 & w10377) | (~pi034 & w19174) | (w10377 & w19174);
assign w10381 = ~w2626 & ~w2670;
assign w10382 = (~w2680 & w10381) | (~w2680 & w19175) | (w10381 & w19175);
assign w10383 = w3181 & ~w10382;
assign w10384 = w2606 & w3191;
assign w10385 = w2739 & w19176;
assign w10386 = ~w10384 & ~w10385;
assign w10387 = ~w6135 & ~w10035;
assign w10388 = ~w2929 & w10387;
assign w10389 = w10386 & w10388;
assign w10390 = ~w10383 & w10389;
assign w10391 = ~w10380 & w10390;
assign w10392 = (~pi038 & w10371) | (~pi038 & w19177) | (w10371 & w19177);
assign w10393 = w10391 & ~w10392;
assign w10394 = ~w10351 & w10393;
assign w10395 = ~w2494 & ~w5950;
assign w10396 = ~w9818 & w10395;
assign w10397 = pi120 & ~w10396;
assign w10398 = (pi003 & w10397) | (pi003 & w19178) | (w10397 & w19178);
assign w10399 = ~w9876 & w10314;
assign w10400 = (~w10399 & w20837) | (~w10399 & w20838) | (w20837 & w20838);
assign w10401 = ~w5965 & w19180;
assign w10402 = pi120 & ~w10401;
assign w10403 = ~w2485 & ~w2831;
assign w10404 = w2805 & ~w10403;
assign w10405 = ~w2496 & ~w2577;
assign w10406 = ~pi120 & ~w10405;
assign w10407 = ~w2475 & w2748;
assign w10408 = w9832 & w10407;
assign w10409 = ~w2836 & ~w10408;
assign w10410 = ~w10404 & ~w10406;
assign w10411 = w10409 & w10410;
assign w10412 = ~w10402 & w10411;
assign w10413 = ~w10398 & ~w10400;
assign w10414 = w10412 & w10413;
assign w10415 = pi044 & ~w10414;
assign w10416 = ~w2771 & ~w2828;
assign w10417 = ~w10315 & ~w10416;
assign w10418 = w2460 & w2522;
assign w10419 = ~w2589 & ~w10418;
assign w10420 = ~w2521 & ~w2827;
assign w10421 = ~w10006 & w10420;
assign w10422 = ~pi003 & ~w2577;
assign w10423 = w10419 & w10422;
assign w10424 = w10421 & w10423;
assign w10425 = (pi003 & ~w2541) | (pi003 & w19181) | (~w2541 & w19181);
assign w10426 = ~w10417 & w10425;
assign w10427 = ~w10424 & ~w10426;
assign w10428 = ~pi016 & w10002;
assign w10429 = w9980 & ~w10428;
assign w10430 = pi120 & ~w2795;
assign w10431 = ~w2521 & w10430;
assign w10432 = ~w5944 & ~w5992;
assign w10433 = w10429 & w10432;
assign w10434 = (~pi044 & w10427) | (~pi044 & w19182) | (w10427 & w19182);
assign w10435 = ~w2772 & ~w5954;
assign w10436 = (~pi120 & ~w10435) | (~pi120 & w19183) | (~w10435 & w19183);
assign w10437 = w2545 & w2796;
assign w10438 = ~w2816 & ~w10437;
assign w10439 = ~w5966 & w10438;
assign w10440 = w2478 & w2801;
assign w10441 = w10439 & ~w10440;
assign w10442 = (~pi003 & ~w10441) | (~pi003 & w19184) | (~w10441 & w19184);
assign w10443 = pi041 & w10265;
assign w10444 = ~w2540 & ~w5925;
assign w10445 = ~w10443 & w10444;
assign w10446 = w5996 & ~w10445;
assign w10447 = w2499 & w2772;
assign w10448 = ~w10305 & ~w10447;
assign w10449 = ~w2834 & ~w5956;
assign w10450 = w10448 & w10449;
assign w10451 = w2465 & w19185;
assign w10452 = w10450 & ~w10451;
assign w10453 = ~w10446 & w10452;
assign w10454 = ~w10442 & w10453;
assign w10455 = ~w10434 & w10454;
assign w10456 = ~w10415 & w10455;
assign w10457 = ~w10394 & w10456;
assign w10458 = w10394 & ~w10456;
assign w10459 = ~w10457 & ~w10458;
assign w10460 = ~w10333 & ~w10459;
assign w10461 = w10333 & w10459;
assign w10462 = ~w10460 & ~w10461;
assign w10463 = ~w6064 & ~w10149;
assign w10464 = pi116 & ~w10463;
assign w10465 = ~w6051 & ~w6074;
assign w10466 = ~w10464 & w10465;
assign w10467 = ~w6206 & ~w10100;
assign w10468 = ~w2955 & w10467;
assign w10469 = pi116 & ~w10468;
assign w10470 = ~w2953 & w6015;
assign w10471 = ~pi022 & w10470;
assign w10472 = w6559 & ~w10471;
assign w10473 = ~w10469 & w10472;
assign w10474 = pi058 & ~w10473;
assign w10475 = ~w3085 & ~w6769;
assign w10476 = ~w3071 & ~w3095;
assign w10477 = (pi116 & ~w10475) | (pi116 & w19186) | (~w10475 & w19186);
assign w10478 = ~w3043 & ~w3067;
assign w10479 = (pi060 & w10478) | (pi060 & w19187) | (w10478 & w19187);
assign w10480 = ~w10477 & w10479;
assign w10481 = (~pi058 & ~w10466) | (~pi058 & w19188) | (~w10466 & w19188);
assign w10482 = ~w10474 & w20839;
assign w10483 = ~w3081 & ~w6016;
assign w10484 = ~w3067 & ~w6253;
assign w10485 = ~w6615 & w10484;
assign w10486 = ~w6719 & w10485;
assign w10487 = w2980 & w2995;
assign w10488 = ~pi000 & w6712;
assign w10489 = ~w10487 & ~w10488;
assign w10490 = ~w2970 & ~w10163;
assign w10491 = w10489 & w10490;
assign w10492 = ~pi116 & ~w10491;
assign w10493 = w3006 & w3023;
assign w10494 = ~w2996 & ~w10493;
assign w10495 = pi116 & ~w10494;
assign w10496 = w2980 & w6006;
assign w10497 = ~pi000 & w10496;
assign w10498 = ~w6067 & ~w10497;
assign w10499 = ~w10495 & w10498;
assign w10500 = pi058 & ~w10499;
assign w10501 = ~w2981 & ~w3081;
assign w10502 = ~w10492 & ~w10500;
assign w10503 = (~pi060 & w10501) | (~pi060 & w19190) | (w10501 & w19190);
assign w10504 = w10502 & w19191;
assign w10505 = w2958 & w3021;
assign w10506 = ~w3007 & ~w6184;
assign w10507 = ~w10505 & w10506;
assign w10508 = (~w6058 & w10507) | (~w6058 & w19192) | (w10507 & w19192);
assign w10509 = pi058 & ~w10508;
assign w10510 = ~w3006 & w3021;
assign w10511 = pi116 & w6236;
assign w10512 = w2982 & w2984;
assign w10513 = ~w10511 & ~w10512;
assign w10514 = ~w6239 & ~w6581;
assign w10515 = w10513 & w10514;
assign w10516 = (~pi116 & w10510) | (~pi116 & w18227) | (w10510 & w18227);
assign w10517 = w3027 & w6051;
assign w10518 = ~w2965 & ~w3006;
assign w10519 = w3001 & ~w10518;
assign w10520 = ~w10517 & ~w10519;
assign w10521 = w2951 & w3090;
assign w10522 = w10520 & ~w10521;
assign w10523 = (~pi058 & ~w10515) | (~pi058 & w19193) | (~w10515 & w19193);
assign w10524 = w10522 & ~w10523;
assign w10525 = ~w10509 & w10524;
assign w10526 = (w10525 & w10482) | (w10525 & w19194) | (w10482 & w19194);
assign w10527 = (w19194 & w20840) | (w19194 & w20841) | (w20840 & w20841);
assign w10528 = (~w19194 & w20842) | (~w19194 & w20843) | (w20842 & w20843);
assign w10529 = ~w10527 & ~w10528;
assign w10530 = ~w10246 & w10529;
assign w10531 = w10246 & ~w10529;
assign w10532 = ~w10530 & ~w10531;
assign w10533 = (~pi529 & ~w10462) | (~pi529 & w20844) | (~w10462 & w20844);
assign w10534 = ~w10462 & ~w10532;
assign w10535 = w10533 & ~w10534;
assign w10536 = pi272 & pi511;
assign w10537 = pi529 & ~w10536;
assign w10538 = ~pi272 & ~pi511;
assign w10539 = w10537 & ~w10538;
assign w10540 = ~w10535 & ~w10539;
assign w10541 = ~w2626 & ~w6670;
assign w10542 = pi118 & w10541;
assign w10543 = ~w2889 & ~w6123;
assign w10544 = w2607 & w10543;
assign w10545 = ~w10542 & ~w10544;
assign w10546 = (pi034 & w10545) | (pi034 & w18195) | (w10545 & w18195);
assign w10547 = w2653 & w3147;
assign w10548 = ~w2714 & ~w10547;
assign w10549 = ~w2865 & ~w10079;
assign w10550 = w2641 & w2648;
assign w10551 = w10549 & ~w10550;
assign w10552 = ~pi034 & ~w10548;
assign w10553 = w10551 & ~w10552;
assign w10554 = ~w10546 & w10553;
assign w10555 = ~pi038 & ~w10554;
assign w10556 = ~w2641 & ~w3186;
assign w10557 = ~pi118 & w10556;
assign w10558 = ~w2882 & ~w2921;
assign w10559 = pi118 & w10558;
assign w10560 = ~w10557 & ~w10559;
assign w10561 = ~w2678 & ~w2729;
assign w10562 = w10561 & w19195;
assign w10563 = (~pi034 & w10560) | (~pi034 & w19196) | (w10560 & w19196);
assign w10564 = (pi034 & w2739) | (pi034 & w3172) | (w2739 & w3172);
assign w10565 = w2920 & w3106;
assign w10566 = w10564 & ~w10565;
assign w10567 = ~w2666 & ~w2693;
assign w10568 = (w2648 & ~w10567) | (w2648 & w19197) | (~w10567 & w19197);
assign w10569 = ~w2729 & ~w2867;
assign w10570 = ~pi066 & ~w10569;
assign w10571 = ~w2740 & ~w10570;
assign w10572 = ~w10568 & w10571;
assign w10573 = ~w10566 & w10572;
assign w10574 = (pi038 & ~w10573) | (pi038 & w19198) | (~w10573 & w19198);
assign w10575 = ~w10078 & ~w10378;
assign w10576 = ~w2674 & w10575;
assign w10577 = w10334 & w10576;
assign w10578 = pi066 & w2601;
assign w10579 = ~w2714 & ~w10578;
assign w10580 = ~w3122 & w10579;
assign w10581 = pi118 & w10580;
assign w10582 = w2601 & ~w2632;
assign w10583 = ~w2677 & w10582;
assign w10584 = ~w10577 & ~w10581;
assign w10585 = w2669 & w2632;
assign w10586 = ~w3154 & ~w10585;
assign w10587 = (pi034 & w3154) | (pi034 & w3172) | (w3154 & w3172);
assign w10588 = (w10587 & ~w3141) | (w10587 & w19199) | (~w3141 & w19199);
assign w10589 = pi034 & ~w10076;
assign w10590 = ~w2615 & ~w2740;
assign w10591 = ~w10589 & w10590;
assign w10592 = pi118 & ~w10591;
assign w10593 = w2605 & w3181;
assign w10594 = w6150 & w10593;
assign w10595 = ~w6154 & ~w10594;
assign w10596 = ~w10592 & w19200;
assign w10597 = (~pi034 & w10584) | (~pi034 & w20845) | (w10584 & w20845);
assign w10598 = w10596 & ~w10597;
assign w10599 = ~w10555 & ~w10574;
assign w10600 = w10598 & w10599;
assign w10601 = ~w2744 & w10600;
assign w10602 = w2744 & ~w10600;
assign w10603 = ~w10601 & ~w10602;
assign w10604 = w6101 & ~w10603;
assign w10605 = ~w6101 & w10603;
assign w10606 = ~w10604 & ~w10605;
assign w10607 = ~w3095 & ~w6056;
assign w10608 = ~w3040 & ~w3054;
assign w10609 = ~pi116 & ~w10608;
assign w10610 = ~w3007 & ~w6239;
assign w10611 = ~w6020 & w10610;
assign w10612 = ~w10609 & w10611;
assign w10613 = ~w3021 & ~w3068;
assign w10614 = (pi116 & ~w10613) | (pi116 & w19201) | (~w10613 & w19201);
assign w10615 = ~w6051 & ~w6209;
assign w10616 = ~w10496 & w10615;
assign w10617 = ~w2970 & ~w2996;
assign w10618 = w10616 & w10617;
assign w10619 = ~w2997 & w19202;
assign w10620 = ~pi116 & ~w10619;
assign w10621 = (w3094 & ~w10150) | (w3094 & w19203) | (~w10150 & w19203);
assign w10622 = ~w10136 & ~w10621;
assign w10623 = ~w10620 & w10622;
assign w10624 = (pi058 & ~w10618) | (pi058 & w19204) | (~w10618 & w19204);
assign w10625 = w10623 & ~w10624;
assign w10626 = (pi060 & ~w10625) | (pi060 & w19205) | (~w10625 & w19205);
assign w10627 = ~pi116 & w10100;
assign w10628 = ~w6713 & ~w10627;
assign w10629 = ~w3013 & ~w3095;
assign w10630 = w10628 & w10629;
assign w10631 = ~w2961 & ~w3094;
assign w10632 = w2992 & ~w10631;
assign w10633 = w2965 & ~w2980;
assign w10634 = pi097 & w10633;
assign w10635 = ~w10632 & ~w10634;
assign w10636 = ~w6211 & ~w10517;
assign w10637 = w10635 & w10636;
assign w10638 = ~pi058 & ~w10637;
assign w10639 = pi057 & w10493;
assign w10640 = ~w3092 & ~w10511;
assign w10641 = ~w10639 & w10640;
assign w10642 = (~pi116 & w3085) | (~pi116 & w19208) | (w3085 & w19208);
assign w10643 = w10641 & ~w10642;
assign w10644 = ~w10638 & w10643;
assign w10645 = (~pi060 & ~w10644) | (~pi060 & w19209) | (~w10644 & w19209);
assign w10646 = ~w6010 & ~w6744;
assign w10647 = (w6015 & ~w10646) | (w6015 & w19210) | (~w10646 & w19210);
assign w10648 = w2953 & w3033;
assign w10649 = ~w2970 & ~w6051;
assign w10650 = (pi116 & ~w10649) | (pi116 & w19211) | (~w10649 & w19211);
assign w10651 = ~w10647 & ~w10650;
assign w10652 = (pi058 & ~w10651) | (pi058 & w19212) | (~w10651 & w19212);
assign w10653 = ~w2954 & ~w6245;
assign w10654 = w3090 & ~w10653;
assign w10655 = ~w3053 & ~w10639;
assign w10656 = w3083 & ~w10655;
assign w10657 = w6021 & w10156;
assign w10658 = ~w2964 & ~w10657;
assign w10659 = ~w10656 & w19213;
assign w10660 = ~w10652 & w10659;
assign w10661 = ~w10645 & w10660;
assign w10662 = ~w10626 & w10661;
assign w10663 = ~w6265 & w10662;
assign w10664 = w6265 & ~w10662;
assign w10665 = ~w10663 & ~w10664;
assign w10666 = w6452 & w20846;
assign w10667 = (pi130 & ~w6452) | (pi130 & w20847) | (~w6452 & w20847);
assign w10668 = ~w10666 & ~w10667;
assign w10669 = w10665 & w10668;
assign w10670 = ~w10665 & ~w10668;
assign w10671 = ~w10669 & ~w10670;
assign w10672 = w10606 & ~w10671;
assign w10673 = ~pi529 & ~w10672;
assign w10674 = ~w10606 & w10671;
assign w10675 = w10673 & ~w10674;
assign w10676 = ~pi130 & pi506;
assign w10677 = pi529 & ~w10676;
assign w10678 = pi130 & ~pi506;
assign w10679 = w10677 & ~w10678;
assign w10680 = ~w10675 & ~w10679;
assign w10681 = ~pi160 & w6948;
assign w10682 = pi160 & ~w6948;
assign w10683 = ~w10681 & ~w10682;
assign w10684 = w2747 & ~w6627;
assign w10685 = ~w2747 & w6627;
assign w10686 = ~w10684 & ~w10685;
assign w10687 = (~pi529 & w10686) | (~pi529 & w19214) | (w10686 & w19214);
assign w10688 = ~w10683 & w10686;
assign w10689 = w10687 & ~w10688;
assign w10690 = pi160 & pi472;
assign w10691 = pi529 & ~w10690;
assign w10692 = ~pi160 & ~pi472;
assign w10693 = w10691 & ~w10692;
assign w10694 = ~w10689 & ~w10693;
assign w10695 = ~w6265 & w6367;
assign w10696 = w6265 & ~w6367;
assign w10697 = ~w10695 & ~w10696;
assign w10698 = ~w2708 & w19215;
assign w10699 = (pi161 & w2708) | (pi161 & w19216) | (w2708 & w19216);
assign w10700 = ~w10698 & ~w10699;
assign w10701 = w10697 & w10700;
assign w10702 = ~w10697 & ~w10700;
assign w10703 = ~w10701 & ~w10702;
assign w10704 = (~pi529 & w10703) | (~pi529 & w19217) | (w10703 & w19217);
assign w10705 = ~w10459 & w10703;
assign w10706 = w10704 & ~w10705;
assign w10707 = ~pi161 & pi409;
assign w10708 = pi529 & ~w10707;
assign w10709 = pi161 & ~pi409;
assign w10710 = w10708 & ~w10709;
assign w10711 = ~w10706 & ~w10710;
assign w10712 = ~w4468 & ~w4474;
assign w10713 = (~pi106 & ~w10712) | (~pi106 & w19218) | (~w10712 & w19218);
assign w10714 = (pi106 & w4062) | (pi106 & w19219) | (w4062 & w19219);
assign w10715 = ~w3994 & ~w4489;
assign w10716 = ~w4519 & ~w7202;
assign w10717 = w10715 & w10716;
assign w10718 = ~w10713 & ~w10714;
assign w10719 = ~w4904 & w10717;
assign w10720 = w10718 & w10719;
assign w10721 = ~w4038 & ~w4095;
assign w10722 = ~pi035 & ~w10721;
assign w10723 = w4015 & w7172;
assign w10724 = ~w4008 & ~w10723;
assign w10725 = ~w10722 & w10724;
assign w10726 = ~pi065 & ~w10725;
assign w10727 = ~w4485 & ~w7856;
assign w10728 = pi035 & ~w10727;
assign w10729 = ~w3991 & ~w4002;
assign w10730 = ~w10728 & w10729;
assign w10731 = pi106 & ~w10730;
assign w10732 = w4448 & w4838;
assign w10733 = ~w7173 & ~w10732;
assign w10734 = pi031 & w4484;
assign w10735 = w3989 & w7165;
assign w10736 = w4053 & w10734;
assign w10737 = ~w10735 & ~w10736;
assign w10738 = ~w10726 & ~w10731;
assign w10739 = w10733 & w10737;
assign w10740 = w10738 & w10739;
assign w10741 = w4000 & ~w4021;
assign w10742 = ~w4523 & ~w10741;
assign w10743 = (~pi065 & ~w4487) | (~pi065 & w19220) | (~w4487 & w19220);
assign w10744 = w10742 & w10743;
assign w10745 = pi106 & ~w4109;
assign w10746 = w10744 & ~w10745;
assign w10747 = w4849 & w19221;
assign w10748 = ~w10746 & ~w10747;
assign w10749 = (w7896 & ~w7210) | (w7896 & w19222) | (~w7210 & w19222);
assign w10750 = (~pi106 & w7859) | (~pi106 & w19223) | (w7859 & w19223);
assign w10751 = ~w4855 & ~w4872;
assign w10752 = w4021 & ~w10751;
assign w10753 = ~w4478 & ~w8176;
assign w10754 = ~w10752 & w10753;
assign w10755 = w10754 & w19224;
assign w10756 = (pi068 & w10748) | (pi068 & w19225) | (w10748 & w19225);
assign w10757 = w4015 & w7186;
assign w10758 = ~w4462 & ~w10757;
assign w10759 = pi031 & w4021;
assign w10760 = (w10759 & w4476) | (w10759 & w19226) | (w4476 & w19226);
assign w10761 = w10758 & ~w10760;
assign w10762 = ~w4840 & ~w8220;
assign w10763 = ~w4112 & ~w4899;
assign w10764 = w4487 & w19227;
assign w10765 = w10763 & w19228;
assign w10766 = pi065 & ~w3993;
assign w10767 = (w10766 & w10732) | (w10766 & w19229) | (w10732 & w19229);
assign w10768 = w10765 & ~w10767;
assign w10769 = (w4529 & w10762) | (w4529 & w19230) | (w10762 & w19230);
assign w10770 = w10768 & ~w10769;
assign w10771 = ~pi065 & ~w10761;
assign w10772 = w10770 & ~w10771;
assign w10773 = ~w10756 & w10772;
assign w10774 = (~pi068 & ~w10740) | (~pi068 & w19231) | (~w10740 & w19231);
assign w10775 = w10773 & ~w10774;
assign w10776 = ~w3417 & ~w3714;
assign w10777 = ~w7777 & w10776;
assign w10778 = pi122 & ~w10777;
assign w10779 = (pi039 & ~w7783) | (pi039 & w19232) | (~w7783 & w19232);
assign w10780 = w4933 & w10779;
assign w10781 = ~w10778 & w10780;
assign w10782 = ~w3732 & ~w3947;
assign w10783 = pi122 & ~w10782;
assign w10784 = ~w3481 & ~w3499;
assign w10785 = ~pi122 & ~w10784;
assign w10786 = w3418 & w3486;
assign w10787 = ~pi039 & ~w3669;
assign w10788 = ~w10786 & w10787;
assign w10789 = ~w10785 & w10788;
assign w10790 = ~w10783 & w10789;
assign w10791 = ~w10781 & ~w10790;
assign w10792 = ~w3388 & ~w7825;
assign w10793 = w3919 & ~w7826;
assign w10794 = w3731 & w10793;
assign w10795 = (pi017 & w10791) | (pi017 & w19233) | (w10791 & w19233);
assign w10796 = ~w3376 & ~w3385;
assign w10797 = ~pi043 & ~w10796;
assign w10798 = pi076 & ~w3381;
assign w10799 = w3935 & ~w10798;
assign w10800 = pi122 & ~w4957;
assign w10801 = ~w3438 & w10800;
assign w10802 = ~pi122 & ~w10799;
assign w10803 = ~w10797 & w10802;
assign w10804 = ~w3493 & ~w3881;
assign w10805 = ~pi039 & ~w7825;
assign w10806 = w10804 & w10805;
assign w10807 = w3412 & w19234;
assign w10808 = ~w3438 & ~w3960;
assign w10809 = w10806 & w10808;
assign w10810 = ~w10807 & w10809;
assign w10811 = ~w3709 & ~w7785;
assign w10812 = w3721 & ~w10811;
assign w10813 = ~pi122 & w7826;
assign w10814 = ~w3448 & ~w10813;
assign w10815 = ~w10812 & w10814;
assign w10816 = pi039 & w10815;
assign w10817 = ~w10810 & ~w10816;
assign w10818 = ~w3440 & ~w3669;
assign w10819 = (~pi122 & ~w10818) | (~pi122 & w18795) | (~w10818 & w18795);
assign w10820 = w3369 & w3420;
assign w10821 = w3412 & w3409;
assign w10822 = ~w10820 & ~w10821;
assign w10823 = ~w3685 & ~w3734;
assign w10824 = w10822 & w10823;
assign w10825 = ~pi077 & w4931;
assign w10826 = ~w3454 & ~w3684;
assign w10827 = ~w10825 & w10826;
assign w10828 = w3756 & ~w10827;
assign w10829 = ~w3394 & ~w4957;
assign w10830 = ~w3374 & ~w10829;
assign w10831 = w3398 & w19235;
assign w10832 = ~w3720 & ~w10831;
assign w10833 = ~w10828 & w19236;
assign w10834 = (~pi039 & ~w10824) | (~pi039 & w20848) | (~w10824 & w20848);
assign w10835 = w10833 & ~w10834;
assign w10836 = (~pi017 & w10817) | (~pi017 & w19237) | (w10817 & w19237);
assign w10837 = w10835 & ~w10836;
assign w10838 = ~w10795 & w10837;
assign w10839 = ~pi084 & w3561;
assign w10840 = ~w3541 & ~w3841;
assign w10841 = ~w10839 & w10840;
assign w10842 = pi091 & ~w10841;
assign w10843 = (pi024 & w10842) | (pi024 & w19238) | (w10842 & w19238);
assign w10844 = pi004 & w3648;
assign w10845 = ~pi091 & w3625;
assign w10846 = w3822 & w10844;
assign w10847 = ~w10845 & ~w10846;
assign w10848 = ~w3788 & ~w4417;
assign w10849 = w10847 & w10848;
assign w10850 = ~pi024 & ~w10849;
assign w10851 = ~w3829 & w19239;
assign w10852 = pi091 & ~w10851;
assign w10853 = ~w3803 & ~w4780;
assign w10854 = w3652 & ~w10853;
assign w10855 = w3522 & w3620;
assign w10856 = ~w3559 & ~w10855;
assign w10857 = ~pi091 & ~w10856;
assign w10858 = pi024 & ~pi091;
assign w10859 = ~w3520 & w3534;
assign w10860 = w10858 & w10859;
assign w10861 = ~w4813 & ~w10860;
assign w10862 = ~w10854 & ~w10857;
assign w10863 = w10861 & w10862;
assign w10864 = ~w10852 & w10863;
assign w10865 = w10864 & w19240;
assign w10866 = pi018 & ~w10865;
assign w10867 = pi004 & w3631;
assign w10868 = ~w3811 & ~w10867;
assign w10869 = w3547 & ~w10868;
assign w10870 = (pi024 & ~w3541) | (pi024 & w19241) | (~w3541 & w19241);
assign w10871 = w3597 & w3773;
assign w10872 = ~w10869 & w19242;
assign w10873 = ~w3639 & ~w4422;
assign w10874 = ~w4820 & ~w10855;
assign w10875 = ~pi024 & w10874;
assign w10876 = ~w3585 & ~w4807;
assign w10877 = w10875 & w10876;
assign w10878 = w3593 & ~w10873;
assign w10879 = w10877 & ~w10878;
assign w10880 = w3518 & w3543;
assign w10881 = ~w3813 & ~w10880;
assign w10882 = ~pi004 & w7730;
assign w10883 = w7692 & ~w10882;
assign w10884 = pi091 & ~w4790;
assign w10885 = ~w3585 & w10884;
assign w10886 = w10881 & w10883;
assign w10887 = ~w10872 & ~w10879;
assign w10888 = ~w3560 & w3784;
assign w10889 = ~w3779 & ~w4408;
assign w10890 = pi091 & ~w7696;
assign w10891 = w10889 & ~w10890;
assign w10892 = (~pi091 & w10888) | (~pi091 & w19243) | (w10888 & w19243);
assign w10893 = ~w7720 & ~w10844;
assign w10894 = ~w3842 & ~w10893;
assign w10895 = w3547 & w3597;
assign w10896 = w3523 & w19244;
assign w10897 = w4370 & w19245;
assign w10898 = ~w10896 & ~w10897;
assign w10899 = ~w3823 & ~w4814;
assign w10900 = ~w10895 & w10899;
assign w10901 = w10898 & w10900;
assign w10902 = (w3858 & w10894) | (w3858 & w19246) | (w10894 & w19246);
assign w10903 = w10901 & ~w10902;
assign w10904 = (~pi024 & ~w10891) | (~pi024 & w19247) | (~w10891 & w19247);
assign w10905 = w10903 & ~w10904;
assign w10906 = (~pi018 & w10887) | (~pi018 & w19248) | (w10887 & w19248);
assign w10907 = w10905 & ~w10906;
assign w10908 = ~w10866 & w10907;
assign w10909 = ~w10838 & w10908;
assign w10910 = w10838 & ~w10908;
assign w10911 = ~w10909 & ~w10910;
assign w10912 = ~w10775 & ~w10911;
assign w10913 = w10775 & w10911;
assign w10914 = ~w10912 & ~w10913;
assign w10915 = w4158 & w4138;
assign w10916 = ~w4234 & ~w4663;
assign w10917 = (~pi113 & ~w10916) | (~pi113 & w19249) | (~w10916 & w19249);
assign w10918 = ~w4193 & ~w4664;
assign w10919 = pi113 & ~w10918;
assign w10920 = w4137 & w4192;
assign w10921 = ~w4254 & ~w4588;
assign w10922 = ~w4719 & ~w10920;
assign w10923 = w10921 & w10922;
assign w10924 = ~w10919 & w10923;
assign w10925 = w10924 & w19250;
assign w10926 = pi096 & ~w10925;
assign w10927 = ~w4149 & ~w4658;
assign w10928 = w4631 & ~w10927;
assign w10929 = ~w4728 & ~w10928;
assign w10930 = ~pi096 & ~w10929;
assign w10931 = w4127 & w4155;
assign w10932 = ~w7062 & ~w10920;
assign w10933 = ~w4251 & w10932;
assign w10934 = pi125 & w4155;
assign w10935 = w4233 & w4625;
assign w10936 = w4241 & w10934;
assign w10937 = ~w10935 & ~w10936;
assign w10938 = ~pi113 & w4198;
assign w10939 = w4144 & w4233;
assign w10940 = ~w10938 & ~w10939;
assign w10941 = w10937 & w10940;
assign w10942 = (pi113 & ~w10933) | (pi113 & w19251) | (~w10933 & w19251);
assign w10943 = w10941 & ~w10942;
assign w10944 = ~w10930 & w10943;
assign w10945 = ~w10926 & w10944;
assign w10946 = pi010 & ~w10945;
assign w10947 = ~pi113 & ~w4205;
assign w10948 = ~w4195 & ~w7929;
assign w10949 = pi113 & w10948;
assign w10950 = ~w10947 & ~w10949;
assign w10951 = w4132 & ~w4594;
assign w10952 = ~w4607 & ~w10951;
assign w10953 = ~pi096 & w10952;
assign w10954 = ~w10950 & w10953;
assign w10955 = ~w4571 & ~w6984;
assign w10956 = w10955 & w19252;
assign w10957 = ~w10954 & ~w10956;
assign w10958 = ~w4128 & ~w4264;
assign w10959 = (w4738 & ~w10958) | (w4738 & w19253) | (~w10958 & w19253);
assign w10960 = (~pi113 & w7928) | (~pi113 & w19254) | (w7928 & w19254);
assign w10961 = ~w4242 & ~w4700;
assign w10962 = w4594 & ~w10961;
assign w10963 = ~w4164 & ~w4578;
assign w10964 = ~w10962 & w10963;
assign w10965 = w10964 & w19255;
assign w10966 = (~pi010 & w10957) | (~pi010 & w19256) | (w10957 & w19256);
assign w10967 = ~w4233 & ~w7099;
assign w10968 = (~pi113 & w10967) | (~pi113 & w18705) | (w10967 & w18705);
assign w10969 = (w4136 & w4580) | (w4136 & w19257) | (w4580 & w19257);
assign w10970 = w4236 & w4570;
assign w10971 = ~w4561 & ~w10970;
assign w10972 = ~w10969 & w10971;
assign w10973 = ~w10968 & w10972;
assign w10974 = ~pi096 & ~w10973;
assign w10975 = ~w7984 & ~w10938;
assign w10976 = pi096 & ~w10975;
assign w10977 = ~w4556 & ~w7015;
assign w10978 = w4548 & w19258;
assign w10979 = w10977 & w19259;
assign w10980 = ~w10976 & w10979;
assign w10981 = ~w10974 & w10980;
assign w10982 = ~w10966 & w10981;
assign w10983 = ~w10946 & w10982;
assign w10984 = ~w4588 & ~w4664;
assign w10985 = (pi113 & ~w7931) | (pi113 & w19260) | (~w7931 & w19260);
assign w10986 = ~w4657 & w4677;
assign w10987 = w6986 & ~w10986;
assign w10988 = ~w10985 & w10987;
assign w10989 = pi096 & ~w10988;
assign w10990 = ~w4250 & ~w4704;
assign w10991 = pi113 & ~w10990;
assign w10992 = w10937 & ~w10991;
assign w10993 = ~w4663 & ~w7978;
assign w10994 = ~pi113 & w10993;
assign w10995 = w4206 & ~w10939;
assign w10996 = w4608 & w10995;
assign w10997 = ~w10994 & ~w10996;
assign w10998 = (~pi096 & ~w10992) | (~pi096 & w19261) | (~w10992 & w19261);
assign w10999 = ~w10997 & ~w10998;
assign w11000 = ~w10989 & w10999;
assign w11001 = ~pi010 & ~w11000;
assign w11002 = ~w4583 & ~w7922;
assign w11003 = w4594 & ~w11002;
assign w11004 = ~pi113 & w10939;
assign w11005 = ~w4269 & ~w11004;
assign w11006 = ~w11003 & w11005;
assign w11007 = pi096 & w11006;
assign w11008 = pi124 & w4204;
assign w11009 = ~w7919 & ~w11008;
assign w11010 = ~w7024 & ~w7978;
assign w11011 = ~pi096 & w11010;
assign w11012 = ~w4238 & ~w7973;
assign w11013 = w11011 & w11012;
assign w11014 = ~pi125 & ~w11009;
assign w11015 = w11013 & ~w11014;
assign w11016 = ~pi125 & w4228;
assign w11017 = w4263 & w4207;
assign w11018 = ~w11016 & ~w11017;
assign w11019 = pi113 & ~w7000;
assign w11020 = ~w7973 & w11019;
assign w11021 = w4216 & ~w4584;
assign w11022 = w11018 & w11021;
assign w11023 = ~w11007 & ~w11015;
assign w11024 = ~w4158 & w4546;
assign w11025 = w4137 & w4126;
assign w11026 = ~w4707 & ~w11025;
assign w11027 = ~w4560 & ~w4609;
assign w11028 = w11026 & w11027;
assign w11029 = (~pi113 & w11024) | (~pi113 & w18821) | (w11024 & w18821);
assign w11030 = (pi113 & w7061) | (pi113 & w18682) | (w7061 & w18682);
assign w11031 = w4127 & w4546;
assign w11032 = ~w4178 & ~w4561;
assign w11033 = ~w11031 & w11032;
assign w11034 = w4726 & ~w11033;
assign w11035 = w4149 & w19262;
assign w11036 = ~w4217 & ~w4601;
assign w11037 = ~w11035 & w11036;
assign w11038 = ~w11034 & w11037;
assign w11039 = ~w11030 & w11038;
assign w11040 = (~pi096 & ~w11028) | (~pi096 & w19263) | (~w11028 & w19263);
assign w11041 = w11039 & ~w11040;
assign w11042 = (pi010 & w11023) | (pi010 & w19264) | (w11023 & w19264);
assign w11043 = w11041 & ~w11042;
assign w11044 = ~w11001 & w11043;
assign w11045 = ~pi215 & w11044;
assign w11046 = pi215 & ~w11044;
assign w11047 = ~w11045 & ~w11046;
assign w11048 = ~w10983 & w11047;
assign w11049 = w10983 & ~w11047;
assign w11050 = ~w11048 & ~w11049;
assign w11051 = w10914 & ~w11050;
assign w11052 = ~pi529 & ~w11051;
assign w11053 = ~w10914 & w11050;
assign w11054 = w11052 & ~w11053;
assign w11055 = ~pi215 & pi401;
assign w11056 = pi529 & ~w11055;
assign w11057 = pi215 & ~pi401;
assign w11058 = w11056 & ~w11057;
assign w11059 = ~w11054 & ~w11058;
assign w11060 = w3401 & w3382;
assign w11061 = ~w3388 & ~w3697;
assign w11062 = (~pi122 & ~w11061) | (~pi122 & w19265) | (~w11061 & w19265);
assign w11063 = (pi122 & w3914) | (pi122 & w19266) | (w3914 & w19266);
assign w11064 = ~w3505 & ~w3674;
assign w11065 = ~w3712 & ~w3714;
assign w11066 = w11064 & w11065;
assign w11067 = ~w11062 & ~w11063;
assign w11068 = ~w3502 & w11066;
assign w11069 = w11067 & w11068;
assign w11070 = pi039 & ~w11069;
assign w11071 = ~w3370 & ~w3920;
assign w11072 = w3394 & ~w11071;
assign w11073 = ~w3485 & ~w3711;
assign w11074 = ~w11072 & w11073;
assign w11075 = ~pi039 & ~w11074;
assign w11076 = w3401 & w3410;
assign w11077 = ~w3709 & ~w11076;
assign w11078 = ~w3382 & ~w11077;
assign w11079 = ~w3712 & ~w3923;
assign w11080 = (pi122 & w11078) | (pi122 & w19267) | (w11078 & w19267);
assign w11081 = ~pi122 & w3669;
assign w11082 = ~w7826 & ~w11081;
assign w11083 = ~w10785 & w11082;
assign w11084 = ~w11080 & w11083;
assign w11085 = ~w11075 & w11084;
assign w11086 = ~w11070 & w11085;
assign w11087 = ~pi017 & ~w11086;
assign w11088 = ~pi076 & w3419;
assign w11089 = ~pi122 & ~w3679;
assign w11090 = ~w3911 & ~w11088;
assign w11091 = pi122 & w11090;
assign w11092 = ~w11089 & ~w11091;
assign w11093 = w3402 & ~w3721;
assign w11094 = ~w3730 & ~w11093;
assign w11095 = ~pi039 & w11094;
assign w11096 = ~w11092 & w11095;
assign w11097 = ~w3753 & ~w4932;
assign w11098 = w3409 & w3397;
assign w11099 = (pi039 & ~w3669) | (pi039 & w19268) | (~w3669 & w19268);
assign w11100 = w11097 & w19269;
assign w11101 = ~w11096 & ~w11100;
assign w11102 = (~pi122 & ~w7788) | (~pi122 & w19270) | (~w7788 & w19270);
assign w11103 = ~pi076 & ~w3449;
assign w11104 = ~w3708 & ~w11103;
assign w11105 = ~w3475 & ~w4940;
assign w11106 = w3721 & ~w11105;
assign w11107 = ~w3703 & ~w4307;
assign w11108 = ~w11106 & w11107;
assign w11109 = w7824 & ~w11088;
assign w11110 = ~w11104 & w11109;
assign w11111 = w11108 & w19271;
assign w11112 = (pi017 & w11101) | (pi017 & w19272) | (w11101 & w19272);
assign w11113 = (w3435 & w3699) | (w3435 & w19273) | (w3699 & w19273);
assign w11114 = w3431 & w4306;
assign w11115 = ~w3684 & ~w11114;
assign w11116 = ~w11113 & w11115;
assign w11117 = ~pi039 & ~w11116;
assign w11118 = w3417 & w19274;
assign w11119 = ~pi122 & w3674;
assign w11120 = ~w4341 & ~w11119;
assign w11121 = w3708 & w3920;
assign w11122 = ~w11081 & ~w11121;
assign w11123 = w3759 & ~w11103;
assign w11124 = ~w3480 & w4344;
assign w11125 = w11123 & ~w11124;
assign w11126 = pi039 & ~w11122;
assign w11127 = ~w11125 & ~w11126;
assign w11128 = ~w4968 & ~w11118;
assign w11129 = w11120 & w11128;
assign w11130 = w11127 & w11129;
assign w11131 = ~w11117 & w11130;
assign w11132 = ~w11112 & w11131;
assign w11133 = ~w11087 & w11132;
assign w11134 = ~w10775 & w11133;
assign w11135 = w10775 & ~w11133;
assign w11136 = ~w11134 & ~w11135;
assign w11137 = ~w10908 & ~w11136;
assign w11138 = w10908 & w11136;
assign w11139 = ~w11137 & ~w11138;
assign w11140 = pi128 & w3982;
assign w11141 = ~w3990 & ~w11140;
assign w11142 = pi106 & ~w11141;
assign w11143 = w10737 & ~w11142;
assign w11144 = ~w4022 & ~w4519;
assign w11145 = ~w7846 & w11144;
assign w11146 = pi106 & ~w11145;
assign w11147 = w4035 & ~w4106;
assign w11148 = ~pi035 & w11147;
assign w11149 = ~w4848 & ~w11148;
assign w11150 = ~w4852 & w11149;
assign w11151 = ~w11146 & w11150;
assign w11152 = ~w4065 & ~w7173;
assign w11153 = (pi106 & ~w4505) | (pi106 & w19275) | (~w4505 & w19275);
assign w11154 = ~w4468 & ~w4896;
assign w11155 = (pi068 & w11154) | (pi068 & w19276) | (w11154 & w19276);
assign w11156 = ~w11153 & w11155;
assign w11157 = pi065 & ~w11151;
assign w11158 = (~pi065 & ~w11143) | (~pi065 & w19277) | (~w11143 & w19277);
assign w11159 = ~w11157 & w20849;
assign w11160 = w3982 & w19278;
assign w11161 = w4037 & w3978;
assign w11162 = ~w7195 & w19279;
assign w11163 = ~w4896 & ~w7205;
assign w11164 = ~w4017 & w11163;
assign w11165 = w11162 & w11164;
assign w11166 = ~w4021 & ~w4451;
assign w11167 = ~w10727 & ~w11166;
assign w11168 = (pi065 & w11167) | (pi065 & w19280) | (w11167 & w19280);
assign w11169 = w3977 & w3988;
assign w11170 = ~pi031 & w4011;
assign w11171 = ~w11169 & ~w11170;
assign w11172 = ~w4073 & ~w4488;
assign w11173 = w11171 & w11172;
assign w11174 = ~pi106 & ~w11173;
assign w11175 = ~w4834 & ~w7172;
assign w11176 = ~w11168 & ~w11174;
assign w11177 = (~pi068 & w11175) | (~pi068 & w19281) | (w11175 & w19281);
assign w11178 = w11176 & w19282;
assign w11179 = w4037 & w4082;
assign w11180 = ~w4041 & ~w4462;
assign w11181 = ~w11179 & w11180;
assign w11182 = (~w11181 & w20944) | (~w11181 & w20945) | (w20944 & w20945);
assign w11183 = ~w4056 & ~w4530;
assign w11184 = (~pi106 & ~w11183) | (~pi106 & w19284) | (~w11183 & w19284);
assign w11185 = ~w4463 & ~w8206;
assign w11186 = ~w4507 & w11185;
assign w11187 = w4002 & w4015;
assign w11188 = w11186 & ~w11187;
assign w11189 = (~pi065 & ~w11188) | (~pi065 & w19285) | (~w11188 & w19285);
assign w11190 = w4832 & ~w4838;
assign w11191 = ~w4499 & ~w11190;
assign w11192 = w4530 & w4015;
assign w11193 = w11191 & ~w11192;
assign w11194 = ~w11189 & w20946;
assign w11195 = (w11194 & w11159) | (w11194 & w19286) | (w11159 & w19286);
assign w11196 = (w19286 & w20850) | (w19286 & w20851) | (w20850 & w20851);
assign w11197 = (~w19286 & w20852) | (~w19286 & w20853) | (w20852 & w20853);
assign w11198 = ~w11196 & ~w11197;
assign w11199 = ~w11044 & w11198;
assign w11200 = w11044 & ~w11198;
assign w11201 = ~w11199 & ~w11200;
assign w11202 = (~pi529 & ~w11139) | (~pi529 & w20854) | (~w11139 & w20854);
assign w11203 = ~w11139 & w11201;
assign w11204 = w11202 & ~w11203;
assign w11205 = ~pi275 & pi523;
assign w11206 = pi529 & ~w11205;
assign w11207 = pi275 & ~pi523;
assign w11208 = w11206 & ~w11207;
assign w11209 = ~w11204 & ~w11208;
assign w11210 = (~pi091 & w10839) | (~pi091 & w19243) | (w10839 & w19243);
assign w11211 = ~w3861 & ~w4411;
assign w11212 = ~w11210 & w11211;
assign w11213 = ~pi024 & ~w11212;
assign w11214 = (w3858 & w3816) | (w3858 & w19287) | (w3816 & w19287);
assign w11215 = w3530 & w3623;
assign w11216 = ~pi004 & w3518;
assign w11217 = ~w4422 & ~w11215;
assign w11218 = (w10858 & ~w11217) | (w10858 & w19288) | (~w11217 & w19288);
assign w11219 = (w3652 & w4402) | (w3652 & w19289) | (w4402 & w19289);
assign w11220 = (w3547 & w3597) | (w3547 & w19290) | (w3597 & w19290);
assign w11221 = ~w4808 & ~w11220;
assign w11222 = ~w3778 & w11221;
assign w11223 = w3523 & ~w3530;
assign w11224 = (pi024 & w11223) | (pi024 & w19291) | (w11223 & w19291);
assign w11225 = ~w3795 & ~w4411;
assign w11226 = ~pi091 & ~w11225;
assign w11227 = ~w11224 & ~w11226;
assign w11228 = w11222 & w11227;
assign w11229 = ~w11214 & ~w11218;
assign w11230 = ~w11219 & w11229;
assign w11231 = w11228 & w19292;
assign w11232 = ~pi018 & ~w11231;
assign w11233 = ~w4360 & ~w4399;
assign w11234 = (w3858 & ~w11233) | (w3858 & w19293) | (~w11233 & w19293);
assign w11235 = ~w3771 & ~w4396;
assign w11236 = w7686 & ~w11235;
assign w11237 = (pi024 & w3817) | (pi024 & w19294) | (w3817 & w19294);
assign w11238 = ~w11236 & ~w11237;
assign w11239 = w3593 & w3783;
assign w11240 = w3570 & w3580;
assign w11241 = ~w3630 & ~w11240;
assign w11242 = w3805 & ~w4383;
assign w11243 = w11241 & ~w11242;
assign w11244 = (~pi024 & ~w11243) | (~pi024 & w19295) | (~w11243 & w19295);
assign w11245 = ~w3587 & ~w3630;
assign w11246 = w11245 & w19296;
assign w11247 = ~pi091 & ~w11246;
assign w11248 = ~w11244 & ~w11247;
assign w11249 = ~w11234 & w11238;
assign w11250 = w11248 & w11249;
assign w11251 = pi018 & ~w11250;
assign w11252 = ~w3582 & ~w4767;
assign w11253 = ~w3852 & w11252;
assign w11254 = ~pi091 & ~w11253;
assign w11255 = ~w4768 & ~w7740;
assign w11256 = (~pi024 & w11254) | (~pi024 & w19297) | (w11254 & w19297);
assign w11257 = ~w3610 & ~w3649;
assign w11258 = ~w10855 & w11257;
assign w11259 = ~w4387 & ~w11239;
assign w11260 = w11258 & w11259;
assign w11261 = w10858 & ~w11260;
assign w11262 = ~w3540 & ~w3625;
assign w11263 = pi005 & ~w11262;
assign w11264 = (w3858 & w11263) | (w3858 & w19298) | (w11263 & w19298);
assign w11265 = ~w3610 & ~w3855;
assign w11266 = w3566 & ~w11265;
assign w11267 = ~w3535 & ~w3778;
assign w11268 = ~w3829 & w11267;
assign w11269 = w3652 & ~w11268;
assign w11270 = ~w11261 & ~w11264;
assign w11271 = ~w11266 & ~w11269;
assign w11272 = w11270 & w19299;
assign w11273 = ~w11251 & w11272;
assign w11274 = ~w11232 & w11273;
assign w11275 = ~w3517 & w11274;
assign w11276 = w3517 & ~w11274;
assign w11277 = ~w11275 & ~w11276;
assign w11278 = w4988 & w11277;
assign w11279 = ~w4988 & ~w11277;
assign w11280 = ~w11278 & ~w11279;
assign w11281 = ~w7220 & w7915;
assign w11282 = w7220 & ~w7915;
assign w11283 = ~w11281 & ~w11282;
assign w11284 = w7991 & w19300;
assign w11285 = (pi284 & ~w7991) | (pi284 & w19301) | (~w7991 & w19301);
assign w11286 = ~w11284 & ~w11285;
assign w11287 = w11283 & w11286;
assign w11288 = ~w11283 & ~w11286;
assign w11289 = ~w11287 & ~w11288;
assign w11290 = ~w11280 & w11289;
assign w11291 = ~pi529 & ~w11290;
assign w11292 = w11280 & ~w11289;
assign w11293 = w11291 & ~w11292;
assign w11294 = pi284 & pi414;
assign w11295 = pi529 & ~w11294;
assign w11296 = ~pi284 & ~pi414;
assign w11297 = w11295 & ~w11296;
assign w11298 = ~w11293 & ~w11297;
assign w11299 = ~w3968 & w7755;
assign w11300 = w3968 & ~w7755;
assign w11301 = ~w11299 & ~w11300;
assign w11302 = ~w3660 & w3873;
assign w11303 = w3660 & ~w3873;
assign w11304 = ~w11302 & ~w11303;
assign w11305 = w11301 & w11304;
assign w11306 = ~w11301 & ~w11304;
assign w11307 = ~w11305 & ~w11306;
assign w11308 = ~pi321 & w4120;
assign w11309 = pi321 & ~w4120;
assign w11310 = ~w11308 & ~w11309;
assign w11311 = w8262 & w11310;
assign w11312 = ~w8262 & ~w11310;
assign w11313 = ~w11311 & ~w11312;
assign w11314 = w11307 & w11313;
assign w11315 = ~pi529 & ~w11314;
assign w11316 = ~w11307 & ~w11313;
assign w11317 = w11315 & ~w11316;
assign w11318 = ~pi321 & pi494;
assign w11319 = pi529 & ~w11318;
assign w11320 = pi321 & ~pi494;
assign w11321 = w11319 & ~w11320;
assign w11322 = ~w11317 & ~w11321;
assign w11323 = w3663 & w11195;
assign w11324 = ~w3663 & ~w11195;
assign w11325 = ~w11323 & ~w11324;
assign w11326 = w4747 & w19302;
assign w11327 = (pi233 & ~w4747) | (pi233 & w19303) | (~w4747 & w19303);
assign w11328 = ~w11326 & ~w11327;
assign w11329 = ~w11044 & w11328;
assign w11330 = w11044 & ~w11328;
assign w11331 = ~w11329 & ~w11330;
assign w11332 = (~pi529 & ~w11325) | (~pi529 & w19304) | (~w11325 & w19304);
assign w11333 = ~w11325 & w11331;
assign w11334 = w11332 & ~w11333;
assign w11335 = ~pi233 & pi477;
assign w11336 = pi529 & ~w11335;
assign w11337 = pi233 & ~pi477;
assign w11338 = w11336 & ~w11337;
assign w11339 = ~w11334 & ~w11338;
assign w11340 = w3663 & w10908;
assign w11341 = ~w3663 & ~w10908;
assign w11342 = ~w11340 & ~w11341;
assign w11343 = ~pi342 & w11044;
assign w11344 = pi342 & ~w11044;
assign w11345 = ~w11343 & ~w11344;
assign w11346 = ~w7220 & w11345;
assign w11347 = w7220 & ~w11345;
assign w11348 = ~w11346 & ~w11347;
assign w11349 = w11342 & ~w11348;
assign w11350 = ~pi529 & ~w11349;
assign w11351 = ~w11342 & w11348;
assign w11352 = w11350 & ~w11351;
assign w11353 = ~pi342 & pi467;
assign w11354 = pi529 & ~w11353;
assign w11355 = pi342 & ~pi467;
assign w11356 = w11354 & ~w11355;
assign w11357 = ~w11352 & ~w11356;
assign w11358 = ~w10838 & w11195;
assign w11359 = w10838 & ~w11195;
assign w11360 = ~w11358 & ~w11359;
assign w11361 = ~w3829 & ~w3844;
assign w11362 = ~w7706 & w11361;
assign w11363 = ~w3795 & ~w3852;
assign w11364 = ~w4755 & ~w4768;
assign w11365 = w11363 & w11364;
assign w11366 = (~pi091 & w11223) | (~pi091 & w19305) | (w11223 & w19305);
assign w11367 = (w10858 & ~w10893) | (w10858 & w19288) | (~w10893 & w19288);
assign w11368 = w3588 & w3604;
assign w11369 = ~w7702 & ~w11368;
assign w11370 = ~w3807 & ~w3850;
assign w11371 = w11369 & w11370;
assign w11372 = w11371 & w19306;
assign w11373 = pi024 & ~w11365;
assign w11374 = w11372 & ~w11373;
assign w11375 = ~w3559 & ~w3805;
assign w11376 = (~pi091 & ~w11375) | (~pi091 & w19308) | (~w11375 & w19308);
assign w11377 = ~w3558 & ~w7687;
assign w11378 = pi091 & ~w11377;
assign w11379 = w3580 & w3631;
assign w11380 = ~w3649 & ~w3771;
assign w11381 = ~w3841 & ~w11379;
assign w11382 = w11380 & w11381;
assign w11383 = ~w11376 & ~w11378;
assign w11384 = ~pi091 & w3788;
assign w11385 = ~pi004 & w3649;
assign w11386 = ~w11384 & ~w11385;
assign w11387 = w3540 & w19309;
assign w11388 = (~pi091 & w4371) | (~pi091 & w19310) | (w4371 & w19310);
assign w11389 = ~w4808 & ~w11388;
assign w11390 = (pi024 & ~w11386) | (pi024 & w19311) | (~w11386 & w19311);
assign w11391 = w11389 & ~w11390;
assign w11392 = ~pi018 & pi024;
assign w11393 = (w11392 & ~w11383) | (w11392 & w19312) | (~w11383 & w19312);
assign w11394 = w11391 & ~w11393;
assign w11395 = ~w3546 & ~w4433;
assign w11396 = (~pi091 & w11395) | (~pi091 & w19313) | (w11395 & w19313);
assign w11397 = (w3588 & ~w3804) | (w3588 & w11368) | (~w3804 & w11368);
assign w11398 = w3608 & w4806;
assign w11399 = ~w3778 & ~w11398;
assign w11400 = ~w11397 & w11399;
assign w11401 = ~w11396 & w11400;
assign w11402 = ~pi024 & ~w11401;
assign w11403 = ~w3530 & ~w4806;
assign w11404 = ~w10873 & ~w11403;
assign w11405 = ~w3816 & ~w10895;
assign w11406 = ~w11404 & w11405;
assign w11407 = ~pi024 & ~w11406;
assign w11408 = ~w3832 & ~w4812;
assign w11409 = ~w3610 & ~w11384;
assign w11410 = w11408 & w11409;
assign w11411 = ~w4391 & ~w11379;
assign w11412 = pi091 & ~w11411;
assign w11413 = w10847 & ~w11412;
assign w11414 = w11410 & w11413;
assign w11415 = ~w11407 & w11414;
assign w11416 = ~pi018 & ~w11415;
assign w11417 = ~w11402 & ~w11416;
assign w11418 = w11394 & w11417;
assign w11419 = (pi018 & ~w11374) | (pi018 & w19314) | (~w11374 & w19314);
assign w11420 = w11417 & w20855;
assign w11421 = ~w11133 & w11420;
assign w11422 = w11133 & ~w11420;
assign w11423 = ~w11421 & ~w11422;
assign w11424 = ~pi147 & w11044;
assign w11425 = pi147 & ~w11044;
assign w11426 = ~w11424 & ~w11425;
assign w11427 = w11423 & w11426;
assign w11428 = ~w11423 & ~w11426;
assign w11429 = ~w11427 & ~w11428;
assign w11430 = (~pi529 & w11429) | (~pi529 & w19315) | (w11429 & w19315);
assign w11431 = ~w11360 & w11429;
assign w11432 = w11430 & ~w11431;
assign w11433 = ~pi147 & pi463;
assign w11434 = pi529 & ~w11433;
assign w11435 = pi147 & ~pi463;
assign w11436 = w11434 & ~w11435;
assign w11437 = ~w11432 & ~w11436;
assign w11438 = ~pi234 & w7034;
assign w11439 = pi234 & ~w7034;
assign w11440 = ~w11438 & ~w11439;
assign w11441 = ~w4749 & w7220;
assign w11442 = w4749 & ~w7220;
assign w11443 = ~w11441 & ~w11442;
assign w11444 = w7773 & ~w11443;
assign w11445 = ~w7773 & w11443;
assign w11446 = ~w11444 & ~w11445;
assign w11447 = (~pi529 & ~w11446) | (~pi529 & w19316) | (~w11446 & w19316);
assign w11448 = ~w11440 & ~w11446;
assign w11449 = w11447 & ~w11448;
assign w11450 = ~pi234 & pi428;
assign w11451 = pi529 & ~w11450;
assign w11452 = pi234 & ~pi428;
assign w11453 = w11451 & ~w11452;
assign w11454 = ~w11449 & ~w11453;
assign w11455 = ~w7302 & w8074;
assign w11456 = w7302 & ~w8074;
assign w11457 = ~w11455 & ~w11456;
assign w11458 = w7655 & w19317;
assign w11459 = (pi140 & ~w7655) | (pi140 & w19318) | (~w7655 & w19318);
assign w11460 = ~w11458 & ~w11459;
assign w11461 = w11457 & w11460;
assign w11462 = ~w11457 & ~w11460;
assign w11463 = ~w11461 & ~w11462;
assign w11464 = (~pi529 & w11463) | (~pi529 & w19319) | (w11463 & w19319);
assign w11465 = ~w554 & w11463;
assign w11466 = w11464 & ~w11465;
assign w11467 = ~pi140 & pi423;
assign w11468 = pi529 & ~w11467;
assign w11469 = pi140 & ~pi423;
assign w11470 = w11468 & ~w11469;
assign w11471 = ~w11466 & ~w11470;
assign w11472 = ~w973 & ~w5101;
assign w11473 = (pi001 & ~w8090) | (pi001 & w19320) | (~w8090 & w19320);
assign w11474 = ~w5118 & w20856;
assign w11475 = (pi114 & w11473) | (pi114 & w20857) | (w11473 & w20857);
assign w11476 = ~w426 & ~w5441;
assign w11477 = w7370 & w11476;
assign w11478 = ~pi001 & ~w11477;
assign w11479 = ~w972 & ~w8130;
assign w11480 = ~pi114 & ~w11479;
assign w11481 = ~w920 & ~w1160;
assign w11482 = w1011 & ~w11481;
assign w11483 = ~w453 & w5073;
assign w11484 = w7311 & w11483;
assign w11485 = ~w1191 & ~w11484;
assign w11486 = ~w11480 & ~w11482;
assign w11487 = (pi001 & w1145) | (pi001 & w19321) | (w1145 & w19321);
assign w11488 = w11486 & w19322;
assign w11489 = ~w11478 & w11488;
assign w11490 = (pi029 & ~w11489) | (pi029 & w20858) | (~w11489 & w20858);
assign w11491 = w417 & w442;
assign w11492 = ~w468 & ~w537;
assign w11493 = ~pi001 & ~w1005;
assign w11494 = w11492 & w11493;
assign w11495 = ~w1196 & ~w8130;
assign w11496 = ~w11491 & w11495;
assign w11497 = w11494 & w11496;
assign w11498 = ~w7367 & w19323;
assign w11499 = pi001 & ~w525;
assign w11500 = ~w11498 & w11499;
assign w11501 = ~w11497 & ~w11500;
assign w11502 = ~w406 & ~w533;
assign w11503 = ~w508 & ~w11502;
assign w11504 = pi114 & ~w443;
assign w11505 = ~w468 & w11504;
assign w11506 = w450 & ~w5100;
assign w11507 = ~w11503 & w11506;
assign w11508 = (~pi029 & w11501) | (~pi029 & w19324) | (w11501 & w19324);
assign w11509 = ~w426 & ~w922;
assign w11510 = (~pi114 & ~w11509) | (~pi114 & w19325) | (~w11509 & w19325);
assign w11511 = ~w531 & ~w5433;
assign w11512 = ~w5119 & w11511;
assign w11513 = w408 & w976;
assign w11514 = w11512 & ~w11513;
assign w11515 = (~pi001 & ~w11514) | (~pi001 & w19326) | (~w11514 & w19326);
assign w11516 = ~w922 & ~w950;
assign w11517 = (~w938 & w11516) | (~w938 & w19327) | (w11516 & w19327);
assign w11518 = w5136 & ~w11517;
assign w11519 = (pi114 & w5142) | (pi114 & w19328) | (w5142 & w19328);
assign w11520 = w993 & w8137;
assign w11521 = ~w444 & ~w5111;
assign w11522 = ~w11520 & w11521;
assign w11523 = ~w11519 & w11522;
assign w11524 = ~w11518 & w11523;
assign w11525 = ~w11515 & w11524;
assign w11526 = ~w11508 & w11525;
assign w11527 = ~w11490 & w11526;
assign w11528 = ~w7576 & w11527;
assign w11529 = w7576 & ~w11527;
assign w11530 = ~w11528 & ~w11529;
assign w11531 = ~w7379 & ~w11530;
assign w11532 = w7379 & w11530;
assign w11533 = ~w11531 & ~w11532;
assign w11534 = w7655 & w19329;
assign w11535 = (pi169 & ~w7655) | (pi169 & w19330) | (~w7655 & w19330);
assign w11536 = ~w11534 & ~w11535;
assign w11537 = ~w7445 & w11536;
assign w11538 = w7445 & ~w11536;
assign w11539 = ~w11537 & ~w11538;
assign w11540 = (~pi529 & ~w11533) | (~pi529 & w20859) | (~w11533 & w20859);
assign w11541 = ~w11533 & ~w11539;
assign w11542 = w11540 & ~w11541;
assign w11543 = pi169 & pi525;
assign w11544 = pi529 & ~w11543;
assign w11545 = ~pi169 & ~pi525;
assign w11546 = w11544 & ~w11545;
assign w11547 = ~w11542 & ~w11546;
assign w11548 = w11457 & w11527;
assign w11549 = ~w11457 & ~w11527;
assign w11550 = ~w11548 & ~w11549;
assign w11551 = ~pi168 & ~w7516;
assign w11552 = pi168 & w7516;
assign w11553 = ~w11551 & ~w11552;
assign w11554 = (~pi529 & ~w11550) | (~pi529 & w19331) | (~w11550 & w19331);
assign w11555 = ~w11550 & ~w11553;
assign w11556 = w11554 & ~w11555;
assign w11557 = ~pi168 & pi411;
assign w11558 = pi529 & ~w11557;
assign w11559 = pi168 & ~pi411;
assign w11560 = w11558 & ~w11559;
assign w11561 = ~w11556 & ~w11560;
assign w11562 = ~w8074 & ~w11530;
assign w11563 = w8074 & w11530;
assign w11564 = ~w11562 & ~w11563;
assign w11565 = w7512 & w19332;
assign w11566 = (pi152 & ~w7512) | (pi152 & w19333) | (~w7512 & w19333);
assign w11567 = ~w11565 & ~w11566;
assign w11568 = ~w7656 & w11567;
assign w11569 = w7656 & ~w11567;
assign w11570 = ~w11568 & ~w11569;
assign w11571 = (~pi529 & ~w11564) | (~pi529 & w19334) | (~w11564 & w19334);
assign w11572 = ~w11564 & ~w11570;
assign w11573 = w11571 & ~w11572;
assign w11574 = pi152 & pi421;
assign w11575 = pi529 & ~w11574;
assign w11576 = ~pi152 & ~pi421;
assign w11577 = w11575 & ~w11576;
assign w11578 = ~w11573 & ~w11577;
assign w11579 = ~w1440 & w8150;
assign w11580 = w1440 & ~w8150;
assign w11581 = ~w11579 & ~w11580;
assign w11582 = w8361 & ~w11581;
assign w11583 = ~w8361 & w11581;
assign w11584 = ~w11582 & ~w11583;
assign w11585 = ~w702 & w8341;
assign w11586 = w702 & ~w8341;
assign w11587 = ~w11585 & ~w11586;
assign w11588 = w1525 & w19335;
assign w11589 = (pi174 & ~w1525) | (pi174 & w19336) | (~w1525 & w19336);
assign w11590 = ~w11588 & ~w11589;
assign w11591 = w11587 & w11590;
assign w11592 = ~w11587 & ~w11590;
assign w11593 = ~w11591 & ~w11592;
assign w11594 = (~pi529 & w11584) | (~pi529 & w19337) | (w11584 & w19337);
assign w11595 = w11584 & w11593;
assign w11596 = w11594 & ~w11595;
assign w11597 = pi174 & pi479;
assign w11598 = pi529 & ~w11597;
assign w11599 = ~pi174 & ~pi479;
assign w11600 = w11598 & ~w11599;
assign w11601 = ~w11596 & ~w11600;
assign w11602 = ~pi220 & w5243;
assign w11603 = pi220 & ~w5243;
assign w11604 = ~w11602 & ~w11603;
assign w11605 = ~w145 & w901;
assign w11606 = w145 & ~w901;
assign w11607 = ~w11605 & ~w11606;
assign w11608 = w11604 & w11607;
assign w11609 = ~w11604 & ~w11607;
assign w11610 = ~w11608 & ~w11609;
assign w11611 = ~w551 & w1128;
assign w11612 = w551 & ~w1128;
assign w11613 = ~w11611 & ~w11612;
assign w11614 = w5899 & w11613;
assign w11615 = ~w5899 & ~w11613;
assign w11616 = ~w11614 & ~w11615;
assign w11617 = (~pi529 & ~w11610) | (~pi529 & w19338) | (~w11610 & w19338);
assign w11618 = ~w11610 & ~w11616;
assign w11619 = w11617 & ~w11618;
assign w11620 = ~pi220 & pi458;
assign w11621 = pi529 & ~w11620;
assign w11622 = pi220 & ~pi458;
assign w11623 = w11621 & ~w11622;
assign w11624 = ~w11619 & ~w11623;
assign w11625 = w8340 & w19339;
assign w11626 = (pi155 & ~w8340) | (pi155 & w19340) | (~w8340 & w19340);
assign w11627 = ~w11625 & ~w11626;
assign w11628 = ~w145 & w702;
assign w11629 = w145 & ~w702;
assign w11630 = ~w11628 & ~w11629;
assign w11631 = w1285 & ~w11630;
assign w11632 = ~w1285 & w11630;
assign w11633 = ~w11631 & ~w11632;
assign w11634 = (~pi529 & ~w11633) | (~pi529 & w19341) | (~w11633 & w19341);
assign w11635 = ~w11627 & ~w11633;
assign w11636 = w11634 & ~w11635;
assign w11637 = ~pi155 & pi476;
assign w11638 = pi529 & ~w11637;
assign w11639 = pi155 & ~pi476;
assign w11640 = w11638 & ~w11639;
assign w11641 = ~w11636 & ~w11640;
assign w11642 = (w1766 & w2199) | (w1766 & w19342) | (w2199 & w19342);
assign w11643 = ~w1707 & ~w2032;
assign w11644 = ~w2261 & ~w8610;
assign w11645 = w11643 & w11644;
assign w11646 = (~pi026 & ~w11645) | (~pi026 & w19343) | (~w11645 & w19343);
assign w11647 = ~w1723 & w1942;
assign w11648 = w1701 & w1727;
assign w11649 = ~w2212 & ~w11648;
assign w11650 = ~w8945 & ~w11647;
assign w11651 = (~pi115 & ~w11650) | (~pi115 & w19344) | (~w11650 & w19344);
assign w11652 = w1734 & w1949;
assign w11653 = ~w1716 & ~w11652;
assign w11654 = ~w2019 & ~w8944;
assign w11655 = pi026 & ~w11654;
assign w11656 = ~w1706 & ~w1956;
assign w11657 = (w1773 & w11655) | (w1773 & w19345) | (w11655 & w19345);
assign w11658 = pi026 & ~w11653;
assign w11659 = ~w11657 & ~w11658;
assign w11660 = ~w11646 & w11659;
assign w11661 = (~pi030 & ~w11660) | (~pi030 & w19346) | (~w11660 & w19346);
assign w11662 = (~pi115 & ~w9189) | (~pi115 & w19347) | (~w9189 & w19347);
assign w11663 = ~w1979 & ~w2007;
assign w11664 = pi115 & ~w11663;
assign w11665 = ~pi026 & ~w8573;
assign w11666 = ~w11664 & w11665;
assign w11667 = ~w11662 & w11666;
assign w11668 = ~w1769 & ~w8947;
assign w11669 = ~w2210 & w11668;
assign w11670 = pi115 & ~w11669;
assign w11671 = w1984 & w2200;
assign w11672 = ~w1738 & ~w11671;
assign w11673 = w9201 & w11672;
assign w11674 = ~w11670 & w11673;
assign w11675 = ~w11667 & ~w11674;
assign w11676 = ~w1761 & ~w2261;
assign w11677 = ~w1745 & w8583;
assign w11678 = w8966 & w11677;
assign w11679 = (pi030 & w11675) | (pi030 & w19348) | (w11675 & w19348);
assign w11680 = ~w1719 & w1997;
assign w11681 = w1693 & w1708;
assign w11682 = ~w2028 & ~w11681;
assign w11683 = pi115 & ~w8582;
assign w11684 = w11682 & ~w11683;
assign w11685 = (~pi115 & w11680) | (~pi115 & w18149) | (w11680 & w18149);
assign w11686 = (~pi026 & ~w11684) | (~pi026 & w19349) | (~w11684 & w19349);
assign w11687 = (~pi115 & ~w2000) | (~pi115 & w20860) | (~w2000 & w20860);
assign w11688 = (~w2260 & ~w1697) | (~w2260 & w19350) | (~w1697 & w19350);
assign w11689 = ~w11687 & ~w11688;
assign w11690 = w1709 & w1964;
assign w11691 = ~w1724 & ~w2222;
assign w11692 = ~w11690 & w11691;
assign w11693 = w2265 & ~w11692;
assign w11694 = ~w2018 & ~w9178;
assign w11695 = ~w8954 & w11694;
assign w11696 = ~w11693 & w11695;
assign w11697 = ~w11689 & w11696;
assign w11698 = ~w11686 & w11697;
assign w11699 = ~w11679 & w11698;
assign w11700 = ~w11661 & w11699;
assign w11701 = w2115 & ~w8422;
assign w11702 = w2095 & w18529;
assign w11703 = ~w2144 & ~w9137;
assign w11704 = w2165 & w11703;
assign w11705 = ~pi085 & w5806;
assign w11706 = ~w8396 & ~w11705;
assign w11707 = ~w9359 & w11706;
assign w11708 = pi089 & ~w11707;
assign w11709 = ~w2063 & ~w2151;
assign w11710 = ~w8487 & w11709;
assign w11711 = (~pi092 & ~w11710) | (~pi092 & w19351) | (~w11710 & w19351);
assign w11712 = ~w2074 & ~w2143;
assign w11713 = (~pi053 & w11712) | (~pi053 & w19352) | (w11712 & w19352);
assign w11714 = ~w11708 & w20861;
assign w11715 = (~pi089 & ~w11704) | (~pi089 & w19353) | (~w11704 & w19353);
assign w11716 = w11714 & ~w11715;
assign w11717 = ~w5859 & ~w8515;
assign w11718 = ~w2054 & w11717;
assign w11719 = pi092 & ~w11718;
assign w11720 = ~w2124 & w5824;
assign w11721 = w5798 & ~w11720;
assign w11722 = ~w11719 & w11721;
assign w11723 = pi089 & ~w11722;
assign w11724 = ~w8478 & ~w8506;
assign w11725 = pi092 & ~w11724;
assign w11726 = ~w9340 & ~w11725;
assign w11727 = ~w2168 & ~w5814;
assign w11728 = (pi092 & ~w8502) | (pi092 & w19354) | (~w8502 & w19354);
assign w11729 = ~w2164 & ~w8421;
assign w11730 = (pi053 & w11729) | (pi053 & w19355) | (w11729 & w19355);
assign w11731 = ~w11728 & w11730;
assign w11732 = (~pi089 & ~w11726) | (~pi089 & w19356) | (~w11726 & w19356);
assign w11733 = w11731 & ~w11732;
assign w11734 = ~w11723 & w11733;
assign w11735 = ~pi092 & ~w2050;
assign w11736 = ~w2051 & w2093;
assign w11737 = w11735 & ~w11736;
assign w11738 = w9082 & ~w9105;
assign w11739 = ~w11737 & ~w11738;
assign w11740 = ~w5844 & ~w8479;
assign w11741 = (~pi089 & w11739) | (~pi089 & w19357) | (w11739 & w19357);
assign w11742 = w2075 & w5855;
assign w11743 = ~w8395 & ~w11742;
assign w11744 = (w2172 & ~w11743) | (w2172 & w19358) | (~w11743 & w19358);
assign w11745 = (~w5868 & w2066) | (~w5868 & w19359) | (w2066 & w19359);
assign w11746 = (~w8496 & ~w9386) | (~w8496 & w19360) | (~w9386 & w19360);
assign w11747 = ~w11744 & w11746;
assign w11748 = ~w11741 & w11747;
assign w11749 = ~w11745 & w11748;
assign w11750 = (w11749 & w11716) | (w11749 & w19361) | (w11716 & w19361);
assign w11751 = ~w11700 & w11750;
assign w11752 = w11700 & ~w11750;
assign w11753 = ~w11751 & ~w11752;
assign w11754 = ~w2369 & ~w5707;
assign w11755 = ~w2296 & w11754;
assign w11756 = pi080 & ~w11755;
assign w11757 = w2345 & ~w5738;
assign w11758 = (pi073 & ~w11757) | (pi073 & w19362) | (~w11757 & w19362);
assign w11759 = w9642 & w11758;
assign w11760 = ~w11756 & w11759;
assign w11761 = ~w2303 & ~w2360;
assign w11762 = pi080 & ~w11761;
assign w11763 = ~pi073 & ~w2348;
assign w11764 = ~w9608 & w11763;
assign w11765 = ~w9741 & w11764;
assign w11766 = ~w11762 & w11765;
assign w11767 = ~w11760 & ~w11766;
assign w11768 = ~w2384 & ~w2406;
assign w11769 = ~w2405 & w8733;
assign w11770 = w8775 & w11769;
assign w11771 = (pi015 & w11767) | (pi015 & w19363) | (w11767 & w19363);
assign w11772 = ~w5706 & ~w8829;
assign w11773 = w8813 & ~w11772;
assign w11774 = ~w8758 & w8891;
assign w11775 = ~w11773 & w11774;
assign w11776 = pi080 & ~w9678;
assign w11777 = ~w2413 & w11776;
assign w11778 = ~pi073 & ~w2406;
assign w11779 = ~w2413 & ~w8832;
assign w11780 = w11778 & w11779;
assign w11781 = ~w5746 & ~w9570;
assign w11782 = ~w9694 & w11781;
assign w11783 = w11780 & w11782;
assign w11784 = ~w2322 & ~w8757;
assign w11785 = w5683 & ~w11784;
assign w11786 = (pi073 & ~w5687) | (pi073 & w19364) | (~w5687 & w19364);
assign w11787 = ~pi080 & w2405;
assign w11788 = ~w11785 & w19365;
assign w11789 = ~w11783 & ~w11788;
assign w11790 = ~w2292 & ~w2348;
assign w11791 = (~pi080 & ~w11790) | (~pi080 & w19366) | (~w11790 & w19366);
assign w11792 = ~w2343 & ~w8856;
assign w11793 = pi080 & ~w11792;
assign w11794 = ~w8737 & ~w9602;
assign w11795 = ~w11793 & w11794;
assign w11796 = pi079 & w2369;
assign w11797 = ~w2350 & ~w2395;
assign w11798 = ~w11796 & w11797;
assign w11799 = w2409 & ~w11798;
assign w11800 = (pi080 & w2304) | (pi080 & w19367) | (w2304 & w19367);
assign w11801 = pi073 & w9587;
assign w11802 = ~w11800 & ~w11801;
assign w11803 = ~w8770 & ~w8828;
assign w11804 = ~w11799 & w11803;
assign w11805 = w11802 & w11804;
assign w11806 = (~pi073 & ~w11795) | (~pi073 & w19368) | (~w11795 & w19368);
assign w11807 = w11805 & ~w11806;
assign w11808 = (~pi015 & w11789) | (~pi015 & w19369) | (w11789 & w19369);
assign w11809 = w11807 & ~w11808;
assign w11810 = ~w11771 & w11809;
assign w11811 = w11809 & w19370;
assign w11812 = (pi146 & ~w11809) | (pi146 & w19371) | (~w11809 & w19371);
assign w11813 = ~w11811 & ~w11812;
assign w11814 = w11753 & w11813;
assign w11815 = ~w11753 & ~w11813;
assign w11816 = ~w11814 & ~w11815;
assign w11817 = (~pi529 & w11816) | (~pi529 & w19372) | (w11816 & w19372);
assign w11818 = ~w9316 & w11816;
assign w11819 = w11817 & ~w11818;
assign w11820 = ~pi146 & pi514;
assign w11821 = pi529 & ~w11820;
assign w11822 = pi146 & ~pi514;
assign w11823 = w11821 & ~w11822;
assign w11824 = ~w11819 & ~w11823;
assign w11825 = ~w1617 & ~w9045;
assign w11826 = ~w9408 & w11825;
assign w11827 = pi002 & ~w11826;
assign w11828 = ~w9035 & w19373;
assign w11829 = (pi117 & w11827) | (pi117 & w19374) | (w11827 & w19374);
assign w11830 = w1639 & w1892;
assign w11831 = ~w8634 & ~w11830;
assign w11832 = w9300 & w11831;
assign w11833 = ~pi002 & ~w11832;
assign w11834 = ~w1601 & w1635;
assign w11835 = w1855 & w19375;
assign w11836 = ~w1920 & ~w11835;
assign w11837 = ~w1609 & ~w9452;
assign w11838 = ~pi117 & ~w11837;
assign w11839 = ~w1586 & ~w1914;
assign w11840 = w1588 & ~w11839;
assign w11841 = ~w11838 & ~w11840;
assign w11842 = (pi002 & w11834) | (pi002 & w19376) | (w11834 & w19376);
assign w11843 = w11841 & w20862;
assign w11844 = (pi036 & ~w19377) | (pi036 & w20863) | (~w19377 & w20863);
assign w11845 = ~w1683 & ~w9021;
assign w11846 = w1927 & ~w11845;
assign w11847 = w1679 & w8631;
assign w11848 = ~w1574 & ~w11847;
assign w11849 = ~w11846 & w11848;
assign w11850 = pi002 & w11849;
assign w11851 = (w1591 & w1659) | (w1591 & w19378) | (w1659 & w19378);
assign w11852 = ~pi002 & ~w9452;
assign w11853 = ~w1546 & w11852;
assign w11854 = ~w1926 & ~w8705;
assign w11855 = ~w11851 & w11854;
assign w11856 = w11853 & w11855;
assign w11857 = ~pi032 & w8702;
assign w11858 = w8644 & ~w11857;
assign w11859 = w1549 & ~w1614;
assign w11860 = w11858 & ~w11859;
assign w11861 = pi117 & ~w1887;
assign w11862 = ~w1546 & w11861;
assign w11863 = ~w11850 & ~w11856;
assign w11864 = ~w1570 & w1895;
assign w11865 = w1552 & w1634;
assign w11866 = ~w1902 & ~w11865;
assign w11867 = ~w9037 & w11866;
assign w11868 = w1582 & w1638;
assign w11869 = w11867 & ~w11868;
assign w11870 = (~pi117 & w11864) | (~pi117 & w19379) | (w11864 & w19379);
assign w11871 = ~pi032 & w1560;
assign w11872 = ~w11871 & w19380;
assign w11873 = w9051 & ~w11872;
assign w11874 = (pi117 & w9059) | (pi117 & w18103) | (w9059 & w18103);
assign w11875 = w9274 & w20864;
assign w11876 = ~w1918 & ~w9027;
assign w11877 = ~w11875 & w11876;
assign w11878 = ~w11874 & w11877;
assign w11879 = ~w11873 & w11878;
assign w11880 = (~pi002 & ~w11869) | (~pi002 & w19381) | (~w11869 & w19381);
assign w11881 = w11879 & ~w11880;
assign w11882 = (~pi036 & w11863) | (~pi036 & w19382) | (w11863 & w19382);
assign w11883 = w11881 & ~w11882;
assign w11884 = ~w11844 & w11883;
assign w11885 = ~w9236 & w9393;
assign w11886 = w9236 & ~w9393;
assign w11887 = ~w11885 & ~w11886;
assign w11888 = ~w11884 & ~w11887;
assign w11889 = w11884 & w11887;
assign w11890 = ~w11888 & ~w11889;
assign w11891 = w11809 & w19383;
assign w11892 = (pi273 & ~w11809) | (pi273 & w19384) | (~w11809 & w19384);
assign w11893 = ~w11891 & ~w11892;
assign w11894 = ~w11750 & w11893;
assign w11895 = w11750 & ~w11893;
assign w11896 = ~w11894 & ~w11895;
assign w11897 = (~pi529 & ~w11890) | (~pi529 & w19385) | (~w11890 & w19385);
assign w11898 = ~w11890 & w11896;
assign w11899 = w11897 & ~w11898;
assign w11900 = ~pi273 & pi427;
assign w11901 = pi529 & ~w11900;
assign w11902 = pi273 & ~pi427;
assign w11903 = w11901 & ~w11902;
assign w11904 = ~w11899 & ~w11903;
assign w11905 = ~w11700 & w11884;
assign w11906 = w11700 & ~w11884;
assign w11907 = ~w11905 & ~w11906;
assign w11908 = ~w9313 & ~w11907;
assign w11909 = w9313 & w11907;
assign w11910 = ~w11908 & ~w11909;
assign w11911 = (w19361 & w20865) | (w19361 & w20866) | (w20865 & w20866);
assign w11912 = (~w19361 & w20867) | (~w19361 & w20868) | (w20867 & w20868);
assign w11913 = ~w11911 & ~w11912;
assign w11914 = ~w9783 & w11913;
assign w11915 = w9783 & ~w11913;
assign w11916 = ~w11914 & ~w11915;
assign w11917 = (~pi529 & ~w11910) | (~pi529 & w20869) | (~w11910 & w20869);
assign w11918 = ~w11910 & ~w11916;
assign w11919 = w11917 & ~w11918;
assign w11920 = pi274 & pi440;
assign w11921 = pi529 & ~w11920;
assign w11922 = ~pi274 & ~pi440;
assign w11923 = w11921 & ~w11922;
assign w11924 = ~w11919 & ~w11923;
assign w11925 = ~pi144 & w9783;
assign w11926 = pi144 & ~w9783;
assign w11927 = ~w11925 & ~w11926;
assign w11928 = w11887 & w11927;
assign w11929 = ~w11887 & ~w11927;
assign w11930 = ~w11928 & ~w11929;
assign w11931 = (~pi529 & w11930) | (~pi529 & w19386) | (w11930 & w19386);
assign w11932 = ~w8719 & w11930;
assign w11933 = w11931 & ~w11932;
assign w11934 = ~pi144 & pi497;
assign w11935 = pi529 & ~w11934;
assign w11936 = pi144 & ~pi497;
assign w11937 = w11935 & ~w11936;
assign w11938 = ~w11933 & ~w11937;
assign w11939 = ~w2286 & w9471;
assign w11940 = w2286 & ~w9471;
assign w11941 = ~w11939 & ~w11940;
assign w11942 = ~w5878 & w8456;
assign w11943 = w5878 & ~w8456;
assign w11944 = ~w11942 & ~w11943;
assign w11945 = w11941 & w11944;
assign w11946 = ~w11941 & ~w11944;
assign w11947 = ~w11945 & ~w11946;
assign w11948 = ~w5779 & w9701;
assign w11949 = w5779 & ~w9701;
assign w11950 = ~w11948 & ~w11949;
assign w11951 = w2429 & w19387;
assign w11952 = (pi283 & ~w2429) | (pi283 & w19388) | (~w2429 & w19388);
assign w11953 = ~w11951 & ~w11952;
assign w11954 = w11950 & w11953;
assign w11955 = ~w11950 & ~w11953;
assign w11956 = ~w11954 & ~w11955;
assign w11957 = (~pi529 & ~w11956) | (~pi529 & w19389) | (~w11956 & w19389);
assign w11958 = w11947 & ~w11956;
assign w11959 = w11957 & ~w11958;
assign w11960 = pi283 & pi498;
assign w11961 = pi529 & ~w11960;
assign w11962 = ~pi283 & ~pi498;
assign w11963 = w11961 & ~w11962;
assign w11964 = ~w11959 & ~w11963;
assign w11965 = ~w1706 & ~w2222;
assign w11966 = ~pi115 & w11965;
assign w11967 = ~w1772 & ~w1964;
assign w11968 = pi115 & w11967;
assign w11969 = ~w11966 & ~w11968;
assign w11970 = ~w1721 & ~w2262;
assign w11971 = w11970 & w19390;
assign w11972 = (~pi026 & w11969) | (~pi026 & w19391) | (w11969 & w19391);
assign w11973 = ~pi115 & w2201;
assign w11974 = (pi115 & ~w1744) | (pi115 & w19392) | (~w1744 & w19392);
assign w11975 = (~w11974 & ~w2201) | (~w11974 & w19393) | (~w2201 & w19393);
assign w11976 = (pi026 & w11975) | (pi026 & w19394) | (w11975 & w19394);
assign w11977 = (w1730 & ~w1743) | (w1730 & w19395) | (~w1743 & w19395);
assign w11978 = ~pi008 & w1983;
assign w11979 = ~w2010 & ~w2029;
assign w11980 = ~w11978 & w11979;
assign w11981 = ~w11972 & ~w11976;
assign w11982 = (pi030 & ~w11981) | (pi030 & w19396) | (~w11981 & w19396);
assign w11983 = ~w1781 & ~w1804;
assign w11984 = w11973 & ~w11983;
assign w11985 = ~w1754 & ~w8578;
assign w11986 = (~w1710 & w11985) | (~w1710 & w19397) | (w11985 & w19397);
assign w11987 = (pi026 & w11984) | (pi026 & w19398) | (w11984 & w19398);
assign w11988 = ~w1829 & ~w11687;
assign w11989 = ~w1836 & ~w2013;
assign w11990 = (~w8573 & w11989) | (~w8573 & w19399) | (w11989 & w19399);
assign w11991 = ~w11988 & w11990;
assign w11992 = ~w2262 & ~w11681;
assign w11993 = ~pi115 & w11992;
assign w11994 = ~w1836 & ~w8972;
assign w11995 = ~w2215 & w11994;
assign w11996 = pi115 & w11995;
assign w11997 = ~w1716 & ~w1819;
assign w11998 = w11993 & w11997;
assign w11999 = ~w11996 & ~w11998;
assign w12000 = ~w1701 & w1727;
assign w12001 = w1708 & w1701;
assign w12002 = ~w2241 & ~w12001;
assign w12003 = (pi026 & w2241) | (pi026 & w2260) | (w2241 & w2260);
assign w12004 = (w12003 & ~w2231) | (w12003 & w19400) | (~w2231 & w19400);
assign w12005 = ~w1732 & ~w2009;
assign w12006 = w2031 & ~w12005;
assign w12007 = ~w1706 & ~w1758;
assign w12008 = w2265 & ~w12007;
assign w12009 = pi115 & w2273;
assign w12010 = w1805 & w12009;
assign w12011 = ~w8973 & ~w12010;
assign w12012 = ~w12006 & ~w12008;
assign w12013 = w12011 & w12012;
assign w12014 = ~w12004 & w12013;
assign w12015 = (~pi026 & w11999) | (~pi026 & w19401) | (w11999 & w19401);
assign w12016 = w12014 & ~w12015;
assign w12017 = (~pi030 & w11987) | (~pi030 & w20870) | (w11987 & w20870);
assign w12018 = w12016 & ~w12017;
assign w12019 = ~w11982 & w12018;
assign w12020 = ~w9551 & w12019;
assign w12021 = w9551 & ~w12019;
assign w12022 = ~w12020 & ~w12021;
assign w12023 = ~w1841 & w9069;
assign w12024 = w1841 & ~w9069;
assign w12025 = ~w12023 & ~w12024;
assign w12026 = w12022 & w12025;
assign w12027 = ~w12022 & ~w12025;
assign w12028 = ~w12026 & ~w12027;
assign w12029 = w8807 & w20871;
assign w12030 = (pi131 & ~w8807) | (pi131 & w20872) | (~w8807 & w20872);
assign w12031 = ~w12029 & ~w12030;
assign w12032 = w8536 & w12031;
assign w12033 = ~w8536 & ~w12031;
assign w12034 = ~w12032 & ~w12033;
assign w12035 = w12028 & w12034;
assign w12036 = ~pi529 & ~w12035;
assign w12037 = ~w12028 & ~w12034;
assign w12038 = w12036 & ~w12037;
assign w12039 = ~pi131 & pi524;
assign w12040 = pi529 & ~w12039;
assign w12041 = pi131 & ~pi524;
assign w12042 = w12040 & ~w12041;
assign w12043 = ~w12038 & ~w12042;
assign w12044 = ~w1545 & ~w1662;
assign w12045 = ~w1571 & ~w8624;
assign w12046 = ~w8628 & ~w8685;
assign w12047 = w12045 & w12046;
assign w12048 = w1554 & ~w1555;
assign w12049 = pi117 & w12048;
assign w12050 = w12047 & ~w12049;
assign w12051 = (~pi002 & ~w12050) | (~pi002 & w19402) | (~w12050 & w19402);
assign w12052 = ~w1565 & ~w1672;
assign w12053 = ~w1906 & w12052;
assign w12054 = (~w12053 & w20873) | (~w12053 & w20874) | (w20873 & w20874);
assign w12055 = ~w1583 & ~w1868;
assign w12056 = (w1577 & ~w12055) | (w1577 & w19404) | (~w12055 & w19404);
assign w12057 = ~w1663 & ~w1903;
assign w12058 = ~w1928 & w12057;
assign w12059 = ~w12051 & ~w12054;
assign w12060 = (pi036 & ~w12059) | (pi036 & w19405) | (~w12059 & w19405);
assign w12061 = ~pi117 & w12052;
assign w12062 = ~w1651 & ~w8693;
assign w12063 = w12061 & ~w12062;
assign w12064 = ~w1603 & ~w8645;
assign w12065 = (~w1560 & w12064) | (~w1560 & w19406) | (w12064 & w19406);
assign w12066 = (pi002 & w12063) | (pi002 & w19407) | (w12063 & w19407);
assign w12067 = w1569 & w1665;
assign w12068 = ~w1683 & ~w12067;
assign w12069 = ~w8634 & ~w9275;
assign w12070 = w1545 & w1577;
assign w12071 = w12069 & ~w12070;
assign w12072 = ~pi002 & ~w12068;
assign w12073 = w12071 & ~w12072;
assign w12074 = ~w12066 & w12073;
assign w12075 = ~pi036 & ~w12074;
assign w12076 = ~pi064 & w1558;
assign w12077 = ~w1683 & ~w12076;
assign w12078 = ~w8694 & w12077;
assign w12079 = ~w9274 & ~w11865;
assign w12080 = ~w1574 & w12079;
assign w12081 = ~pi117 & ~w12080;
assign w12082 = w1558 & w1544;
assign w12083 = ~w11830 & w19408;
assign w12084 = ~w12081 & w12083;
assign w12085 = (~pi002 & ~w12084) | (~pi002 & w19409) | (~w12084 & w19409);
assign w12086 = w1634 & w1549;
assign w12087 = ~w8695 & ~w12086;
assign w12088 = (pi002 & w8695) | (pi002 & w9244) | (w8695 & w9244);
assign w12089 = (w12088 & ~w9430) | (w12088 & w20875) | (~w9430 & w20875);
assign w12090 = (pi117 & w1663) | (pi117 & w1629) | (w1663 & w1629);
assign w12091 = ~w1545 & ~w1657;
assign w12092 = w9051 & ~w12091;
assign w12093 = pi002 & w1577;
assign w12094 = w1652 & w12093;
assign w12095 = ~w9048 & ~w12094;
assign w12096 = ~w12090 & w12095;
assign w12097 = ~w12089 & w12096;
assign w12098 = ~w12092 & w12097;
assign w12099 = ~w12085 & w12098;
assign w12100 = w12099 & w19410;
assign w12101 = ~w12019 & w12100;
assign w12102 = w12019 & ~w12100;
assign w12103 = ~w12101 & ~w12102;
assign w12104 = w1844 & ~w12103;
assign w12105 = ~w1844 & w12103;
assign w12106 = ~w12104 & ~w12105;
assign w12107 = ~w8533 & w8992;
assign w12108 = w8533 & ~w8992;
assign w12109 = ~w12107 & ~w12108;
assign w12110 = w8807 & w20876;
assign w12111 = (pi135 & ~w8807) | (pi135 & w20877) | (~w8807 & w20877);
assign w12112 = ~w12110 & ~w12111;
assign w12113 = w12109 & w12112;
assign w12114 = ~w12109 & ~w12112;
assign w12115 = ~w12113 & ~w12114;
assign w12116 = ~w12106 & w12115;
assign w12117 = ~pi529 & ~w12116;
assign w12118 = w12106 & ~w12115;
assign w12119 = w12117 & ~w12118;
assign w12120 = ~pi135 & pi430;
assign w12121 = pi529 & ~w12120;
assign w12122 = pi135 & ~pi430;
assign w12123 = w12121 & ~w12122;
assign w12124 = ~w12119 & ~w12123;
assign w12125 = w9700 & w19411;
assign w12126 = (pi230 & ~w9700) | (pi230 & w19412) | (~w9700 & w19412);
assign w12127 = ~w12125 & ~w12126;
assign w12128 = ~w5779 & w8456;
assign w12129 = w5779 & ~w8456;
assign w12130 = ~w12128 & ~w12129;
assign w12131 = w2044 & ~w12130;
assign w12132 = ~w2044 & w12130;
assign w12133 = ~w12131 & ~w12132;
assign w12134 = (~pi529 & ~w12133) | (~pi529 & w19413) | (~w12133 & w19413);
assign w12135 = ~w12127 & ~w12133;
assign w12136 = w12134 & ~w12135;
assign w12137 = ~pi230 & pi491;
assign w12138 = pi529 & ~w12137;
assign w12139 = pi230 & ~pi491;
assign w12140 = w12138 & ~w12139;
assign w12141 = ~w12136 & ~w12140;
assign w12142 = ~w1692 & w12100;
assign w12143 = w1692 & ~w12100;
assign w12144 = ~w12142 & ~w12143;
assign w12145 = w9072 & w12144;
assign w12146 = ~w9072 & ~w12144;
assign w12147 = ~w12145 & ~w12146;
assign w12148 = ~pi180 & w9618;
assign w12149 = pi180 & ~w9618;
assign w12150 = ~w12148 & ~w12149;
assign w12151 = ~w5779 & w8533;
assign w12152 = w5779 & ~w8533;
assign w12153 = ~w12151 & ~w12152;
assign w12154 = w12150 & w12153;
assign w12155 = ~w12150 & ~w12153;
assign w12156 = ~w12154 & ~w12155;
assign w12157 = (~pi529 & ~w12156) | (~pi529 & w19414) | (~w12156 & w19414);
assign w12158 = ~w12147 & ~w12156;
assign w12159 = w12157 & ~w12158;
assign w12160 = ~pi180 & pi402;
assign w12161 = pi529 & ~w12160;
assign w12162 = pi180 & ~pi402;
assign w12163 = w12161 & ~w12162;
assign w12164 = ~w12159 & ~w12163;
assign w12165 = w6789 & w10333;
assign w12166 = ~w6789 & ~w10333;
assign w12167 = ~w12165 & ~w12166;
assign w12168 = w10244 & w19415;
assign w12169 = (pi148 & ~w10244) | (pi148 & w19416) | (~w10244 & w19416);
assign w12170 = ~w12168 & ~w12169;
assign w12171 = ~w10171 & w12170;
assign w12172 = w10171 & ~w12170;
assign w12173 = ~w12171 & ~w12172;
assign w12174 = (~pi529 & ~w12167) | (~pi529 & w20878) | (~w12167 & w20878);
assign w12175 = ~w12167 & w12173;
assign w12176 = w12174 & ~w12175;
assign w12177 = ~pi148 & pi519;
assign w12178 = pi529 & ~w12177;
assign w12179 = pi148 & ~pi519;
assign w12180 = w12178 & ~w12179;
assign w12181 = ~w12176 & ~w12180;
assign w12182 = ~w10092 & w10333;
assign w12183 = w10092 & ~w10333;
assign w12184 = ~w12182 & ~w12183;
assign w12185 = ~w10014 & ~w12184;
assign w12186 = w10014 & w12184;
assign w12187 = ~w12185 & ~w12186;
assign w12188 = ~w10148 & w19417;
assign w12189 = (pi167 & w10148) | (pi167 & w19418) | (w10148 & w19418);
assign w12190 = ~w12188 & ~w12189;
assign w12191 = ~w6869 & w12190;
assign w12192 = w6869 & ~w12190;
assign w12193 = ~w12191 & ~w12192;
assign w12194 = (~pi529 & ~w12187) | (~pi529 & w19419) | (~w12187 & w19419);
assign w12195 = ~w12187 & ~w12193;
assign w12196 = w12194 & ~w12195;
assign w12197 = pi167 & pi492;
assign w12198 = pi529 & ~w12197;
assign w12199 = ~pi167 & ~pi492;
assign w12200 = w12198 & ~w12199;
assign w12201 = ~w12196 & ~w12200;
assign w12202 = ~w6786 & ~w12184;
assign w12203 = w6786 & w12184;
assign w12204 = ~w12202 & ~w12203;
assign w12205 = w10244 & w19420;
assign w12206 = (pi223 & ~w10244) | (pi223 & w19421) | (~w10244 & w19421);
assign w12207 = ~w12205 & ~w12206;
assign w12208 = ~w6869 & w12207;
assign w12209 = w6869 & ~w12207;
assign w12210 = ~w12208 & ~w12209;
assign w12211 = (~pi529 & ~w12204) | (~pi529 & w19422) | (~w12204 & w19422);
assign w12212 = ~w12204 & ~w12210;
assign w12213 = w12211 & ~w12212;
assign w12214 = pi223 & pi518;
assign w12215 = pi529 & ~w12214;
assign w12216 = ~pi223 & ~pi518;
assign w12217 = w12215 & ~w12216;
assign w12218 = ~w12213 & ~w12217;
assign w12219 = w6551 & ~w9918;
assign w12220 = ~w6551 & w9918;
assign w12221 = ~w12219 & ~w12220;
assign w12222 = w3101 & w19423;
assign w12223 = (pi376 & ~w3101) | (pi376 & w19424) | (~w3101 & w19424);
assign w12224 = ~w12222 & ~w12223;
assign w12225 = w9924 & w12224;
assign w12226 = ~w9924 & ~w12224;
assign w12227 = ~w12225 & ~w12226;
assign w12228 = ~w12221 & ~w12227;
assign w12229 = ~pi529 & ~w12228;
assign w12230 = w12221 & w12227;
assign w12231 = w12229 & ~w12230;
assign w12232 = pi376 & pi459;
assign w12233 = pi529 & ~w12232;
assign w12234 = ~pi376 & ~pi459;
assign w12235 = w12233 & ~w12234;
assign w12236 = ~w12231 & ~w12235;
assign w12237 = ~w2520 & ~w5925;
assign w12238 = ~pi120 & ~w12237;
assign w12239 = ~w2753 & ~w9963;
assign w12240 = ~w9967 & w12239;
assign w12241 = ~w12238 & w12240;
assign w12242 = w2453 & ~w2563;
assign w12243 = ~w2820 & ~w12242;
assign w12244 = (pi003 & ~w12243) | (pi003 & w19427) | (~w12243 & w19427);
assign w12245 = w2752 & ~w5927;
assign w12246 = ~w2812 & ~w2817;
assign w12247 = pi120 & w2776;
assign w12248 = w12246 & ~w12247;
assign w12249 = (w2499 & w12245) | (w2499 & w10447) | (w12245 & w10447);
assign w12250 = w12248 & ~w12249;
assign w12251 = ~w12244 & w12250;
assign w12252 = (pi044 & ~w12251) | (pi044 & w19428) | (~w12251 & w19428);
assign w12253 = ~w2558 & ~w10437;
assign w12254 = ~pi120 & w12253;
assign w12255 = ~w2588 & ~w5946;
assign w12256 = ~w9820 & w12255;
assign w12257 = pi120 & w12256;
assign w12258 = ~w2542 & ~w9876;
assign w12259 = w12254 & w12258;
assign w12260 = ~w12257 & ~w12259;
assign w12261 = ~w2449 & ~w2469;
assign w12262 = (~pi003 & w12260) | (~pi003 & w19429) | (w12260 & w19429);
assign w12263 = ~w2479 & ~w2819;
assign w12264 = pi120 & ~w12263;
assign w12265 = ~w2449 & ~w2563;
assign w12266 = w2456 & ~w12265;
assign w12267 = ~w2524 & ~w12266;
assign w12268 = ~w12264 & w12267;
assign w12269 = pi003 & ~w12268;
assign w12270 = w2455 & w5955;
assign w12271 = ~w2588 & ~w12270;
assign w12272 = ~w5954 & ~w10294;
assign w12273 = ~pi003 & ~w12271;
assign w12274 = w12272 & ~w12273;
assign w12275 = w2485 & w19430;
assign w12276 = w12274 & ~w12275;
assign w12277 = ~w12269 & w12276;
assign w12278 = ~pi044 & ~w12277;
assign w12279 = (pi003 & w5923) | (pi003 & w9832) | (w5923 & w9832);
assign w12280 = ~w2764 & ~w9951;
assign w12281 = w9849 & w12280;
assign w12282 = w12279 & ~w12281;
assign w12283 = (pi120 & w2812) | (pi120 & w19431) | (w2812 & w19431);
assign w12284 = ~w2492 & ~w2520;
assign w12285 = w5996 & ~w12284;
assign w12286 = pi003 & w2499;
assign w12287 = w2569 & w12286;
assign w12288 = ~w5979 & ~w12287;
assign w12289 = ~w12283 & w12288;
assign w12290 = ~w12282 & w19432;
assign w12291 = ~w12262 & ~w12278;
assign w12292 = w12291 & w19433;
assign w12293 = ~w2596 & w12292;
assign w12294 = w2596 & ~w12292;
assign w12295 = ~w12293 & ~w12294;
assign w12296 = w10603 & ~w12295;
assign w12297 = ~w10603 & w12295;
assign w12298 = ~w12296 & ~w12297;
assign w12299 = ~w6175 & w10662;
assign w12300 = w6175 & ~w10662;
assign w12301 = ~w12299 & ~w12300;
assign w12302 = w6452 & w20879;
assign w12303 = (pi134 & ~w6452) | (pi134 & w20880) | (~w6452 & w20880);
assign w12304 = ~w12302 & ~w12303;
assign w12305 = w12301 & w12304;
assign w12306 = ~w12301 & ~w12304;
assign w12307 = ~w12305 & ~w12306;
assign w12308 = ~w12298 & w12307;
assign w12309 = ~pi529 & ~w12308;
assign w12310 = w12298 & ~w12307;
assign w12311 = w12309 & ~w12310;
assign w12312 = ~pi134 & pi417;
assign w12313 = pi529 & ~w12312;
assign w12314 = pi134 & ~pi417;
assign w12315 = w12313 & ~w12314;
assign w12316 = ~w12311 & ~w12315;
assign w12317 = ~pi319 & w6786;
assign w12318 = pi319 & ~w6786;
assign w12319 = ~w12317 & ~w12318;
assign w12320 = w6456 & w12319;
assign w12321 = ~w6456 & ~w12319;
assign w12322 = ~w12320 & ~w12321;
assign w12323 = ~w2596 & w6005;
assign w12324 = w2596 & ~w6005;
assign w12325 = ~w12323 & ~w12324;
assign w12326 = w10017 & w12325;
assign w12327 = ~w10017 & ~w12325;
assign w12328 = ~w12326 & ~w12327;
assign w12329 = w12322 & w12328;
assign w12330 = ~pi529 & ~w12329;
assign w12331 = ~w12322 & ~w12328;
assign w12332 = w12330 & ~w12331;
assign w12333 = ~pi319 & pi500;
assign w12334 = pi529 & ~w12333;
assign w12335 = pi319 & ~pi500;
assign w12336 = w12334 & ~w12335;
assign w12337 = ~w12332 & ~w12336;
assign w12338 = ~w6265 & w6786;
assign w12339 = w6265 & ~w6786;
assign w12340 = ~w12338 & ~w12339;
assign w12341 = ~pi356 & w6869;
assign w12342 = pi356 & ~w6869;
assign w12343 = ~w12341 & ~w12342;
assign w12344 = w12340 & w12343;
assign w12345 = ~w12340 & ~w12343;
assign w12346 = ~w12344 & ~w12345;
assign w12347 = ~w2744 & w10014;
assign w12348 = w2744 & ~w10014;
assign w12349 = ~w12347 & ~w12348;
assign w12350 = w12301 & w12349;
assign w12351 = ~w12301 & ~w12349;
assign w12352 = ~w12350 & ~w12351;
assign w12353 = w12346 & w12352;
assign w12354 = ~pi529 & ~w12353;
assign w12355 = ~w12346 & ~w12352;
assign w12356 = w12354 & ~w12355;
assign w12357 = ~pi356 & pi398;
assign w12358 = pi529 & ~w12357;
assign w12359 = pi356 & ~pi398;
assign w12360 = w12358 & ~w12359;
assign w12361 = ~w12356 & ~w12360;
assign w12362 = w10174 & w10456;
assign w12363 = ~w10174 & ~w10456;
assign w12364 = ~w12362 & ~w12363;
assign w12365 = ~w6843 & ~w6908;
assign w12366 = pi090 & ~w12365;
assign w12367 = w3250 & w6859;
assign w12368 = ~w3252 & ~w12367;
assign w12369 = ~w12366 & w12368;
assign w12370 = (~pi088 & ~w12369) | (~pi088 & w19434) | (~w12369 & w19434);
assign w12371 = pi049 & w3203;
assign w12372 = ~w6401 & ~w12371;
assign w12373 = ~w3209 & w12372;
assign w12374 = pi090 & ~w12373;
assign w12375 = w3231 & w3250;
assign w12376 = w6893 & ~w12375;
assign w12377 = ~w12374 & w12376;
assign w12378 = pi088 & ~w12377;
assign w12379 = ~w3324 & ~w3343;
assign w12380 = pi090 & w12379;
assign w12381 = w6418 & w12380;
assign w12382 = ~w3289 & ~w3322;
assign w12383 = ~pi090 & w12382;
assign w12384 = ~w12381 & ~w12383;
assign w12385 = ~w12378 & w19435;
assign w12386 = pi006 & ~w12385;
assign w12387 = ~w3234 & ~w6398;
assign w12388 = w3262 & ~w12387;
assign w12389 = ~pi090 & w3324;
assign w12390 = ~w6284 & ~w12389;
assign w12391 = ~w12388 & w12390;
assign w12392 = pi088 & w12391;
assign w12393 = w3226 & w3248;
assign w12394 = ~w6940 & ~w12393;
assign w12395 = ~w3329 & ~w6860;
assign w12396 = w12394 & w12395;
assign w12397 = ~w3322 & ~w6347;
assign w12398 = ~pi088 & w12397;
assign w12399 = w12396 & w12398;
assign w12400 = (w3286 & w6283) | (w3286 & w19436) | (w6283 & w19436);
assign w12401 = ~w3238 & w6516;
assign w12402 = w6803 & ~w12401;
assign w12403 = pi090 & ~w6917;
assign w12404 = ~w3329 & w12403;
assign w12405 = ~w12400 & w12402;
assign w12406 = ~w12392 & ~w12399;
assign w12407 = ~w3205 & ~w3252;
assign w12408 = (~pi090 & ~w12407) | (~pi090 & w19437) | (~w12407 & w19437);
assign w12409 = ~w6379 & ~w6504;
assign w12410 = ~w6419 & w12409;
assign w12411 = w6287 & w6470;
assign w12412 = w12410 & ~w12411;
assign w12413 = (~pi088 & ~w12412) | (~pi088 & w19438) | (~w12412 & w19438);
assign w12414 = ~w3213 & ~w6357;
assign w12415 = ~w6503 & ~w12414;
assign w12416 = ~w3211 & ~w3313;
assign w12417 = (~w3249 & w12416) | (~w3249 & w19439) | (w12416 & w19439);
assign w12418 = w3295 & ~w12417;
assign w12419 = ~w6410 & ~w6802;
assign w12420 = ~w10188 & w12419;
assign w12421 = ~w12418 & w12420;
assign w12422 = ~w12413 & w12421;
assign w12423 = ~w12415 & w12422;
assign w12424 = (~pi006 & w12406) | (~pi006 & w19440) | (w12406 & w19440);
assign w12425 = w12423 & ~w12424;
assign w12426 = ~w12386 & w12425;
assign w12427 = ~pi271 & w12426;
assign w12428 = pi271 & ~w12426;
assign w12429 = ~w12427 & ~w12428;
assign w12430 = ~w10526 & w12429;
assign w12431 = w10526 & ~w12429;
assign w12432 = ~w12430 & ~w12431;
assign w12433 = w12364 & ~w12432;
assign w12434 = ~pi529 & ~w12433;
assign w12435 = ~w12364 & w12432;
assign w12436 = w12434 & ~w12435;
assign w12437 = ~pi271 & pi437;
assign w12438 = pi529 & ~w12437;
assign w12439 = pi271 & ~pi437;
assign w12440 = w12438 & ~w12439;
assign w12441 = ~w12436 & ~w12440;
assign w12442 = ~pi225 & w6948;
assign w12443 = pi225 & ~w6948;
assign w12444 = ~w12442 & ~w12443;
assign w12445 = w2945 & ~w10697;
assign w12446 = ~w2945 & w10697;
assign w12447 = ~w12445 & ~w12446;
assign w12448 = (~pi529 & ~w12447) | (~pi529 & w19441) | (~w12447 & w19441);
assign w12449 = ~w12444 & ~w12447;
assign w12450 = w12448 & ~w12449;
assign w12451 = ~pi225 & pi464;
assign w12452 = pi529 & ~w12451;
assign w12453 = pi225 & ~pi464;
assign w12454 = w12452 & ~w12453;
assign w12455 = ~w12450 & ~w12454;
assign w12456 = w6639 & ~w12295;
assign w12457 = ~w6639 & w12295;
assign w12458 = ~w12456 & ~w12457;
assign w12459 = w10661 & w19442;
assign w12460 = (pi181 & ~w10661) | (pi181 & w19443) | (~w10661 & w19443);
assign w12461 = ~w12459 & ~w12460;
assign w12462 = ~w6367 & w6530;
assign w12463 = w6367 & ~w6530;
assign w12464 = ~w12462 & ~w12463;
assign w12465 = w12461 & w12464;
assign w12466 = ~w12461 & ~w12464;
assign w12467 = ~w12465 & ~w12466;
assign w12468 = ~w12458 & w12467;
assign w12469 = ~pi529 & ~w12468;
assign w12470 = w12458 & ~w12467;
assign w12471 = w12469 & ~w12470;
assign w12472 = ~pi181 & pi429;
assign w12473 = pi529 & ~w12472;
assign w12474 = pi181 & ~pi429;
assign w12475 = w12473 & ~w12474;
assign w12476 = ~w12471 & ~w12475;
assign w12477 = ~w10600 & w12292;
assign w12478 = w10600 & ~w12292;
assign w12479 = ~w12477 & ~w12478;
assign w12480 = ~w9891 & ~w12479;
assign w12481 = w9891 & w12479;
assign w12482 = ~w12480 & ~w12481;
assign w12483 = ~pi349 & w6098;
assign w12484 = pi349 & ~w6098;
assign w12485 = ~w12483 & ~w12484;
assign w12486 = ~w3353 & w12485;
assign w12487 = w3353 & ~w12485;
assign w12488 = ~w12486 & ~w12487;
assign w12489 = w12482 & ~w12488;
assign w12490 = ~pi529 & ~w12489;
assign w12491 = ~w12482 & w12488;
assign w12492 = w12490 & ~w12491;
assign w12493 = ~pi349 & pi507;
assign w12494 = pi529 & ~w12493;
assign w12495 = pi349 & ~pi507;
assign w12496 = w12494 & ~w12495;
assign w12497 = ~w12492 & ~w12496;
assign w12498 = ~w10394 & w10526;
assign w12499 = w10394 & ~w10526;
assign w12500 = ~w12498 & ~w12499;
assign w12501 = ~pi145 & w12426;
assign w12502 = pi145 & ~w12426;
assign w12503 = ~w12501 & ~w12502;
assign w12504 = w12184 & w12503;
assign w12505 = ~w12184 & ~w12503;
assign w12506 = ~w12504 & ~w12505;
assign w12507 = (~pi529 & w12506) | (~pi529 & w19444) | (w12506 & w19444);
assign w12508 = ~w12500 & w12506;
assign w12509 = w12507 & ~w12508;
assign w12510 = ~pi145 & pi469;
assign w12511 = pi529 & ~w12510;
assign w12512 = pi145 & ~pi469;
assign w12513 = w12511 & ~w12512;
assign w12514 = ~w12509 & ~w12513;
assign w12515 = ~w10171 & ~w10459;
assign w12516 = w10171 & w10459;
assign w12517 = ~w12515 & ~w12516;
assign w12518 = ~pi256 & w12426;
assign w12519 = pi256 & ~w12426;
assign w12520 = ~w12518 & ~w12519;
assign w12521 = ~w10246 & w12520;
assign w12522 = w10246 & ~w12520;
assign w12523 = ~w12521 & ~w12522;
assign w12524 = w12517 & ~w12523;
assign w12525 = ~pi529 & ~w12524;
assign w12526 = ~w12517 & w12523;
assign w12527 = w12525 & ~w12526;
assign w12528 = ~pi256 & pi462;
assign w12529 = pi529 & ~w12528;
assign w12530 = pi256 & ~pi462;
assign w12531 = w12529 & ~w12530;
assign w12532 = ~w12527 & ~w12531;
assign w12533 = ~w3102 & ~w12479;
assign w12534 = w3102 & w12479;
assign w12535 = ~w12533 & ~w12534;
assign w12536 = ~pi222 & w6530;
assign w12537 = pi222 & ~w6530;
assign w12538 = ~w12536 & ~w12537;
assign w12539 = ~w3353 & w12538;
assign w12540 = w3353 & ~w12538;
assign w12541 = ~w12539 & ~w12540;
assign w12542 = w12535 & ~w12541;
assign w12543 = ~pi529 & ~w12542;
assign w12544 = ~w12535 & w12541;
assign w12545 = w12543 & ~w12544;
assign w12546 = ~pi222 & pi493;
assign w12547 = pi529 & ~w12546;
assign w12548 = pi222 & ~pi493;
assign w12549 = w12547 & ~w12548;
assign w12550 = ~w12545 & ~w12549;
assign w12551 = ~pi129 & w10983;
assign w12552 = pi129 & ~w10983;
assign w12553 = ~w12551 & ~w12552;
assign w12554 = w11136 & w12553;
assign w12555 = ~w11136 & ~w12553;
assign w12556 = ~w12554 & ~w12555;
assign w12557 = (~pi529 & ~w12556) | (~pi529 & w19445) | (~w12556 & w19445);
assign w12558 = ~w11301 & ~w12556;
assign w12559 = w12557 & ~w12558;
assign w12560 = pi129 & pi420;
assign w12561 = pi529 & ~w12560;
assign w12562 = ~pi129 & ~pi420;
assign w12563 = w12561 & ~w12562;
assign w12564 = ~w12559 & ~w12563;
assign w12565 = w8244 & ~w11301;
assign w12566 = ~w8244 & w11301;
assign w12567 = ~w12565 & ~w12566;
assign w12568 = ~pi270 & w4276;
assign w12569 = pi270 & ~w4276;
assign w12570 = ~w12568 & ~w12569;
assign w12571 = w8262 & w12570;
assign w12572 = ~w8262 & ~w12570;
assign w12573 = ~w12571 & ~w12572;
assign w12574 = ~w12567 & w12573;
assign w12575 = ~pi529 & ~w12574;
assign w12576 = w12567 & ~w12573;
assign w12577 = w12575 & ~w12576;
assign w12578 = ~pi270 & pi451;
assign w12579 = pi529 & ~w12578;
assign w12580 = pi270 & ~pi451;
assign w12581 = w12579 & ~w12580;
assign w12582 = ~w12577 & ~w12581;
assign w12583 = ~w7755 & ~w11423;
assign w12584 = w7755 & w11423;
assign w12585 = ~w12583 & ~w12584;
assign w12586 = ~pi170 & w10775;
assign w12587 = pi170 & ~w10775;
assign w12588 = ~w12586 & ~w12587;
assign w12589 = ~w4276 & w12588;
assign w12590 = w4276 & ~w12588;
assign w12591 = ~w12589 & ~w12590;
assign w12592 = (~pi529 & ~w12585) | (~pi529 & w19446) | (~w12585 & w19446);
assign w12593 = ~w12585 & ~w12591;
assign w12594 = w12592 & ~w12593;
assign w12595 = pi170 & pi522;
assign w12596 = pi529 & ~w12595;
assign w12597 = ~pi170 & ~pi522;
assign w12598 = w12596 & ~w12597;
assign w12599 = ~w12594 & ~w12598;
assign w12600 = ~w4120 & ~w11423;
assign w12601 = w4120 & w11423;
assign w12602 = ~w12600 & ~w12601;
assign w12603 = ~pi232 & w10983;
assign w12604 = pi232 & ~w10983;
assign w12605 = ~w12603 & ~w12604;
assign w12606 = ~w4276 & w12605;
assign w12607 = w4276 & ~w12605;
assign w12608 = ~w12606 & ~w12607;
assign w12609 = (~pi529 & ~w12602) | (~pi529 & w19447) | (~w12602 & w19447);
assign w12610 = ~w12602 & ~w12608;
assign w12611 = w12609 & ~w12610;
assign w12612 = pi232 & pi471;
assign w12613 = pi529 & ~w12612;
assign w12614 = ~pi232 & ~pi471;
assign w12615 = w12613 & ~w12614;
assign w12616 = ~w12611 & ~w12615;
assign w12617 = ~w7845 & w11274;
assign w12618 = w7845 & ~w11274;
assign w12619 = ~w12617 & ~w12618;
assign w12620 = w4831 & ~w12619;
assign w12621 = ~w4831 & w12619;
assign w12622 = ~w12620 & ~w12621;
assign w12623 = ~w4749 & w7034;
assign w12624 = w4749 & ~w7034;
assign w12625 = ~w12623 & ~w12624;
assign w12626 = w7913 & w19448;
assign w12627 = (pi372 & ~w7913) | (pi372 & w19449) | (~w7913 & w19449);
assign w12628 = ~w12626 & ~w12627;
assign w12629 = w12625 & w12628;
assign w12630 = ~w12625 & ~w12628;
assign w12631 = ~w12629 & ~w12630;
assign w12632 = ~w12622 & ~w12631;
assign w12633 = ~pi529 & ~w12632;
assign w12634 = w12622 & w12631;
assign w12635 = w12633 & ~w12634;
assign w12636 = pi372 & pi446;
assign w12637 = pi529 & ~w12636;
assign w12638 = ~pi372 & ~pi446;
assign w12639 = w12637 & ~w12638;
assign w12640 = ~w12635 & ~w12639;
assign w12641 = w7223 & ~w12619;
assign w12642 = ~w7223 & w12619;
assign w12643 = ~w12641 & ~w12642;
assign w12644 = w7991 & w19450;
assign w12645 = (pi285 & ~w7991) | (pi285 & w19451) | (~w7991 & w19451);
assign w12646 = ~w12644 & ~w12645;
assign w12647 = w12625 & w12646;
assign w12648 = ~w12625 & ~w12646;
assign w12649 = ~w12647 & ~w12648;
assign w12650 = ~w12643 & ~w12649;
assign w12651 = ~pi529 & ~w12650;
assign w12652 = w12643 & w12649;
assign w12653 = w12651 & ~w12652;
assign w12654 = pi285 & pi455;
assign w12655 = pi529 & ~w12654;
assign w12656 = ~pi285 & ~pi455;
assign w12657 = w12655 & ~w12656;
assign w12658 = ~w12653 & ~w12657;
assign w12659 = w4443 & w11274;
assign w12660 = ~w4443 & ~w11274;
assign w12661 = ~w12659 & ~w12660;
assign w12662 = ~pi352 & w8232;
assign w12663 = pi352 & ~w8232;
assign w12664 = ~w12662 & ~w12663;
assign w12665 = ~w7992 & w12664;
assign w12666 = w7992 & ~w12664;
assign w12667 = ~w12665 & ~w12666;
assign w12668 = w12661 & w12667;
assign w12669 = ~pi529 & ~w12668;
assign w12670 = ~w12661 & ~w12667;
assign w12671 = w12669 & ~w12670;
assign w12672 = pi352 & pi489;
assign w12673 = pi529 & ~w12672;
assign w12674 = ~pi352 & ~pi489;
assign w12675 = w12673 & ~w12674;
assign w12676 = ~w12671 & ~w12675;
assign w12677 = ~pi207 & w7123;
assign w12678 = pi207 & ~w7123;
assign w12679 = ~w12677 & ~w12678;
assign w12680 = w8235 & w12679;
assign w12681 = ~w8235 & ~w12679;
assign w12682 = ~w12680 & ~w12681;
assign w12683 = (~pi529 & w12682) | (~pi529 & w19452) | (w12682 & w19452);
assign w12684 = ~w12619 & w12682;
assign w12685 = w12683 & ~w12684;
assign w12686 = ~pi207 & pi419;
assign w12687 = pi529 & ~w12686;
assign w12688 = pi207 & ~pi419;
assign w12689 = w12687 & ~w12688;
assign w12690 = ~w12685 & ~w12689;
assign w12691 = w4443 & w7915;
assign w12692 = ~w4443 & ~w7915;
assign w12693 = ~w12691 & ~w12692;
assign w12694 = ~pi231 & w7123;
assign w12695 = pi231 & ~w7123;
assign w12696 = ~w12694 & ~w12695;
assign w12697 = ~w7992 & w12696;
assign w12698 = w7992 & ~w12696;
assign w12699 = ~w12697 & ~w12698;
assign w12700 = w12693 & ~w12699;
assign w12701 = ~pi529 & ~w12700;
assign w12702 = ~w12693 & w12699;
assign w12703 = w12701 & ~w12702;
assign w12704 = ~pi231 & pi460;
assign w12705 = pi529 & ~w12704;
assign w12706 = pi231 & ~pi460;
assign w12707 = w12705 & ~w12706;
assign w12708 = ~w12703 & ~w12707;
assign w12709 = ~w3660 & ~w11360;
assign w12710 = w3660 & w11360;
assign w12711 = ~w12709 & ~w12710;
assign w12712 = ~pi354 & ~w11443;
assign w12713 = pi354 & w11443;
assign w12714 = ~w12712 & ~w12713;
assign w12715 = w12711 & w12714;
assign w12716 = ~pi529 & ~w12715;
assign w12717 = ~w12711 & ~w12714;
assign w12718 = w12716 & ~w12717;
assign w12719 = ~pi354 & pi434;
assign w12720 = pi529 & ~w12719;
assign w12721 = pi354 & ~pi434;
assign w12722 = w12720 & ~w12721;
assign w12723 = ~w12718 & ~w12722;
assign w12724 = w3515 & w19453;
assign w12725 = (pi166 & ~w3515) | (pi166 & w19454) | (~w3515 & w19454);
assign w12726 = ~w12724 & ~w12725;
assign w12727 = w10911 & w12726;
assign w12728 = ~w10911 & ~w12726;
assign w12729 = ~w12727 & ~w12728;
assign w12730 = (~pi529 & w12729) | (~pi529 & w19455) | (w12729 & w19455);
assign w12731 = ~w11443 & w12729;
assign w12732 = w12730 & ~w12731;
assign w12733 = ~pi166 & pi508;
assign w12734 = pi529 & ~w12733;
assign w12735 = pi166 & ~pi508;
assign w12736 = w12734 & ~w12735;
assign w12737 = ~w12732 & ~w12736;
assign w12738 = w5246 & w7379;
assign w12739 = ~w5246 & ~w7379;
assign w12740 = ~w12738 & ~w12739;
assign w12741 = w7655 & w19456;
assign w12742 = (pi133 & ~w7655) | (pi133 & w19457) | (~w7655 & w19457);
assign w12743 = ~w12741 & ~w12742;
assign w12744 = ~w8074 & w12743;
assign w12745 = w8074 & ~w12743;
assign w12746 = ~w12744 & ~w12745;
assign w12747 = (~pi529 & ~w12740) | (~pi529 & w20881) | (~w12740 & w20881);
assign w12748 = ~w12740 & w12746;
assign w12749 = w12747 & ~w12748;
assign w12750 = ~pi133 & pi456;
assign w12751 = pi529 & ~w12750;
assign w12752 = pi133 & ~pi456;
assign w12753 = w12751 & ~w12752;
assign w12754 = ~w12749 & ~w12753;
assign w12755 = w5578 & ~w11581;
assign w12756 = ~w5578 & w11581;
assign w12757 = ~w12755 & ~w12756;
assign w12758 = w1365 & w20882;
assign w12759 = (pi257 & ~w1365) | (pi257 & w20883) | (~w1365 & w20883);
assign w12760 = ~w12758 & ~w12759;
assign w12761 = w11587 & w12760;
assign w12762 = ~w11587 & ~w12760;
assign w12763 = ~w12761 & ~w12762;
assign w12764 = ~w12757 & ~w12763;
assign w12765 = ~pi529 & ~w12764;
assign w12766 = w12757 & w12763;
assign w12767 = w12765 & ~w12766;
assign w12768 = pi257 & pi486;
assign w12769 = pi529 & ~w12768;
assign w12770 = ~pi257 & ~pi486;
assign w12771 = w12769 & ~w12770;
assign w12772 = ~w12767 & ~w12771;
assign w12773 = w1131 & w7445;
assign w12774 = ~w1131 & ~w7445;
assign w12775 = ~w12773 & ~w12774;
assign w12776 = w700 & w19458;
assign w12777 = (pi156 & ~w700) | (pi156 & w19459) | (~w700 & w19459);
assign w12778 = ~w12776 & ~w12777;
assign w12779 = ~w7513 & w12778;
assign w12780 = w7513 & ~w12778;
assign w12781 = ~w12779 & ~w12780;
assign w12782 = (~pi529 & ~w12775) | (~pi529 & w19460) | (~w12775 & w19460);
assign w12783 = ~w12775 & w12781;
assign w12784 = w12782 & ~w12783;
assign w12785 = ~pi156 & pi403;
assign w12786 = pi529 & ~w12785;
assign w12787 = pi156 & ~pi403;
assign w12788 = w12786 & ~w12787;
assign w12789 = ~w12784 & ~w12788;
assign w12790 = ~w1127 & w19461;
assign w12791 = (pi165 & w1127) | (pi165 & w19462) | (w1127 & w19462);
assign w12792 = ~w12790 & ~w12791;
assign w12793 = w11630 & w12792;
assign w12794 = ~w11630 & ~w12792;
assign w12795 = ~w12793 & ~w12794;
assign w12796 = (~pi529 & w12795) | (~pi529 & w19463) | (w12795 & w19463);
assign w12797 = ~w11530 & w12795;
assign w12798 = w12796 & ~w12797;
assign w12799 = ~pi165 & pi424;
assign w12800 = pi529 & ~w12799;
assign w12801 = pi165 & ~pi424;
assign w12802 = w12800 & ~w12801;
assign w12803 = ~w12798 & ~w12802;
assign w12804 = ~pi219 & ~w11630;
assign w12805 = pi219 & w11630;
assign w12806 = ~w12804 & ~w12805;
assign w12807 = ~w1021 & w7445;
assign w12808 = w1021 & ~w7445;
assign w12809 = ~w12807 & ~w12808;
assign w12810 = ~w7576 & w12809;
assign w12811 = w7576 & ~w12809;
assign w12812 = ~w12810 & ~w12811;
assign w12813 = (~pi529 & ~w12806) | (~pi529 & w19464) | (~w12806 & w19464);
assign w12814 = ~w12806 & w12812;
assign w12815 = w12813 & ~w12814;
assign w12816 = ~pi219 & pi422;
assign w12817 = pi529 & ~w12816;
assign w12818 = pi219 & ~pi422;
assign w12819 = w12817 & ~w12818;
assign w12820 = ~w12815 & ~w12819;
assign w12821 = ~w9393 & ~w11907;
assign w12822 = w9393 & w11907;
assign w12823 = ~w12821 & ~w12822;
assign w12824 = w11809 & w19465;
assign w12825 = (pi227 & ~w11809) | (pi227 & w19466) | (~w11809 & w19466);
assign w12826 = ~w12824 & ~w12825;
assign w12827 = ~w9783 & w12826;
assign w12828 = w9783 & ~w12826;
assign w12829 = ~w12827 & ~w12828;
assign w12830 = (~pi529 & ~w12823) | (~pi529 & w19467) | (~w12823 & w19467);
assign w12831 = ~w12823 & w12829;
assign w12832 = w12830 & ~w12831;
assign w12833 = ~pi227 & pi425;
assign w12834 = pi529 & ~w12833;
assign w12835 = pi227 & ~pi425;
assign w12836 = w12834 & ~w12835;
assign w12837 = ~w12832 & ~w12836;
assign w12838 = w9151 & w9313;
assign w12839 = ~w9151 & ~w9313;
assign w12840 = ~w12838 & ~w12839;
assign w12841 = ~pi149 & w9783;
assign w12842 = pi149 & ~w9783;
assign w12843 = ~w12841 & ~w12842;
assign w12844 = ~w9393 & w12843;
assign w12845 = w9393 & ~w12843;
assign w12846 = ~w12844 & ~w12845;
assign w12847 = w12840 & ~w12846;
assign w12848 = ~pi529 & ~w12847;
assign w12849 = ~w12840 & w12846;
assign w12850 = w12848 & ~w12849;
assign w12851 = ~pi149 & pi452;
assign w12852 = pi529 & ~w12851;
assign w12853 = pi149 & ~pi452;
assign w12854 = w12852 & ~w12853;
assign w12855 = ~w12850 & ~w12854;
assign w12856 = w5785 & ~w11941;
assign w12857 = ~w5785 & w11941;
assign w12858 = ~w12856 & ~w12857;
assign w12859 = w2196 & w19468;
assign w12860 = (pi373 & ~w2196) | (pi373 & w19469) | (~w2196 & w19469);
assign w12861 = ~w12859 & ~w12860;
assign w12862 = w11950 & w12861;
assign w12863 = ~w11950 & ~w12861;
assign w12864 = ~w12862 & ~w12863;
assign w12865 = (~pi529 & w12864) | (~pi529 & w19470) | (w12864 & w19470);
assign w12866 = w12858 & w12864;
assign w12867 = w12865 & ~w12866;
assign w12868 = pi373 & pi465;
assign w12869 = pi529 & ~w12868;
assign w12870 = ~pi373 & ~pi465;
assign w12871 = w12869 & ~w12870;
assign w12872 = ~w12867 & ~w12871;
assign w12873 = ~w9124 & w20884;
assign w12874 = (pi357 & w9124) | (pi357 & w20885) | (w9124 & w20885);
assign w12875 = ~w12873 & ~w12874;
assign w12876 = ~w8456 & w8899;
assign w12877 = w8456 & ~w8899;
assign w12878 = ~w12876 & ~w12877;
assign w12879 = w12875 & w12878;
assign w12880 = ~w12875 & ~w12878;
assign w12881 = ~w12879 & ~w12880;
assign w12882 = ~w1841 & w8716;
assign w12883 = w1841 & ~w8716;
assign w12884 = ~w12882 & ~w12883;
assign w12885 = w12109 & w12884;
assign w12886 = ~w12109 & ~w12884;
assign w12887 = ~w12885 & ~w12886;
assign w12888 = w12881 & w12887;
assign w12889 = ~pi529 & ~w12888;
assign w12890 = ~w12881 & ~w12887;
assign w12891 = w12889 & ~w12890;
assign w12892 = ~pi357 & pi473;
assign w12893 = pi529 & ~w12892;
assign w12894 = pi357 & ~pi473;
assign w12895 = w12893 & ~w12894;
assign w12896 = ~w12891 & ~w12895;
assign w12897 = ~w9471 & ~w12103;
assign w12898 = w9471 & w12103;
assign w12899 = ~w12897 & ~w12898;
assign w12900 = w19051 & w20886;
assign w12901 = (pi350 & ~w19051) | (pi350 & w20887) | (~w19051 & w20887);
assign w12902 = ~w12900 & ~w12901;
assign w12903 = ~w2431 & w12902;
assign w12904 = w2431 & ~w12902;
assign w12905 = ~w12903 & ~w12904;
assign w12906 = (~pi529 & ~w12899) | (~pi529 & w20888) | (~w12899 & w20888);
assign w12907 = ~w12899 & ~w12905;
assign w12908 = w12906 & ~w12907;
assign w12909 = pi350 & pi454;
assign w12910 = pi529 & ~w12909;
assign w12911 = ~pi350 & ~pi454;
assign w12912 = w12910 & ~w12911;
assign w12913 = ~w12908 & ~w12912;
assign w12914 = w5777 & w19471;
assign w12915 = (pi163 & ~w5777) | (pi163 & w19472) | (~w5777 & w19472);
assign w12916 = ~w12914 & ~w12915;
assign w12917 = w9803 & ~w11907;
assign w12918 = ~w9803 & w11907;
assign w12919 = ~w12917 & ~w12918;
assign w12920 = (~pi529 & ~w12919) | (~pi529 & w19473) | (~w12919 & w19473);
assign w12921 = ~w12916 & ~w12919;
assign w12922 = w12920 & ~w12921;
assign w12923 = ~pi163 & pi504;
assign w12924 = pi529 & ~w12923;
assign w12925 = pi163 & ~pi504;
assign w12926 = w12924 & ~w12925;
assign w12927 = ~w12922 & ~w12926;
assign w12928 = ~w2198 & ~w12103;
assign w12929 = w2198 & w12103;
assign w12930 = ~w12928 & ~w12929;
assign w12931 = ~w9617 & w20889;
assign w12932 = (pi229 & w9617) | (pi229 & w20890) | (w9617 & w20890);
assign w12933 = ~w12931 & ~w12932;
assign w12934 = ~w2431 & w12933;
assign w12935 = w2431 & ~w12933;
assign w12936 = ~w12934 & ~w12935;
assign w12937 = (~pi529 & ~w12930) | (~pi529 & w20891) | (~w12930 & w20891);
assign w12938 = ~w12930 & w12936;
assign w12939 = w12937 & ~w12938;
assign w12940 = ~pi229 & pi474;
assign w12941 = pi529 & ~w12940;
assign w12942 = pi229 & ~pi474;
assign w12943 = w12941 & ~w12942;
assign w12944 = ~w12939 & ~w12943;
assign w12945 = w10017 & ~w10665;
assign w12946 = ~w10017 & w10665;
assign w12947 = ~w12945 & ~w12946;
assign w12948 = ~pi269 & w6869;
assign w12949 = pi269 & ~w6869;
assign w12950 = ~w12948 & ~w12949;
assign w12951 = w6456 & w12950;
assign w12952 = ~w6456 & ~w12950;
assign w12953 = ~w12951 & ~w12952;
assign w12954 = ~w12947 & w12953;
assign w12955 = ~pi529 & ~w12954;
assign w12956 = w12947 & ~w12953;
assign w12957 = w12955 & ~w12956;
assign w12958 = ~pi269 & pi415;
assign w12959 = pi529 & ~w12958;
assign w12960 = pi269 & ~pi415;
assign w12961 = w12959 & ~w12960;
assign w12962 = ~w12957 & ~w12961;
assign w12963 = w2747 & w10526;
assign w12964 = ~w2747 & ~w10526;
assign w12965 = ~w12963 & ~w12964;
assign w12966 = w6366 & w19474;
assign w12967 = (pi224 & ~w6366) | (pi224 & w19475) | (~w6366 & w19475);
assign w12968 = ~w12966 & ~w12967;
assign w12969 = ~w12426 & w12968;
assign w12970 = w12426 & ~w12968;
assign w12971 = ~w12969 & ~w12970;
assign w12972 = (~pi529 & ~w12965) | (~pi529 & w19476) | (~w12965 & w19476);
assign w12973 = ~w12965 & w12971;
assign w12974 = w12972 & ~w12973;
assign w12975 = ~pi224 & pi399;
assign w12976 = pi529 & ~w12975;
assign w12977 = pi224 & ~pi399;
assign w12978 = w12976 & ~w12977;
assign w12979 = ~w12974 & ~w12978;
assign w12980 = ~w2596 & ~w12500;
assign w12981 = w2596 & w12500;
assign w12982 = ~w12980 & ~w12981;
assign w12983 = ~pi353 & ~w10697;
assign w12984 = pi353 & w10697;
assign w12985 = ~w12983 & ~w12984;
assign w12986 = w12982 & w12985;
assign w12987 = ~pi529 & ~w12986;
assign w12988 = ~w12982 & ~w12985;
assign w12989 = w12987 & ~w12988;
assign w12990 = ~pi353 & pi510;
assign w12991 = pi529 & ~w12990;
assign w12992 = pi353 & ~pi510;
assign w12993 = w12991 & ~w12992;
assign w12994 = ~w12989 & ~w12993;
assign w12995 = w2747 & w10456;
assign w12996 = ~w2747 & ~w10456;
assign w12997 = ~w12995 & ~w12996;
assign w12998 = ~pi370 & w12426;
assign w12999 = pi370 & ~w12426;
assign w13000 = ~w12998 & ~w12999;
assign w13001 = ~w6265 & w13000;
assign w13002 = w6265 & ~w13000;
assign w13003 = ~w13001 & ~w13002;
assign w13004 = w12997 & ~w13003;
assign w13005 = ~pi529 & ~w13004;
assign w13006 = ~w12997 & w13003;
assign w13007 = w13005 & ~w13006;
assign w13008 = ~pi370 & pi433;
assign w13009 = pi529 & ~w13008;
assign w13010 = pi370 & ~pi433;
assign w13011 = w13009 & ~w13010;
assign w13012 = ~w13007 & ~w13011;
assign w13013 = w4123 & w11420;
assign w13014 = ~w4123 & ~w11420;
assign w13015 = ~w13013 & ~w13014;
assign w13016 = ~pi157 & w10983;
assign w13017 = pi157 & ~w10983;
assign w13018 = ~w13016 & ~w13017;
assign w13019 = ~w10775 & w13018;
assign w13020 = w10775 & ~w13018;
assign w13021 = ~w13019 & ~w13020;
assign w13022 = w13015 & ~w13021;
assign w13023 = ~pi529 & ~w13022;
assign w13024 = ~w13015 & w13021;
assign w13025 = w13023 & ~w13024;
assign w13026 = ~pi157 & pi521;
assign w13027 = pi529 & ~w13026;
assign w13028 = pi157 & ~pi521;
assign w13029 = w13027 & ~w13028;
assign w13030 = ~w13025 & ~w13029;
assign w13031 = w10911 & w11420;
assign w13032 = ~w10911 & ~w11420;
assign w13033 = ~w13031 & ~w13032;
assign w13034 = (w19286 & w20892) | (w19286 & w20893) | (w20892 & w20893);
assign w13035 = (~w19286 & w20894) | (~w19286 & w20895) | (w20894 & w20895);
assign w13036 = ~w13034 & ~w13035;
assign w13037 = ~w10983 & w13036;
assign w13038 = w10983 & ~w13036;
assign w13039 = ~w13037 & ~w13038;
assign w13040 = (~pi529 & ~w13033) | (~pi529 & w20896) | (~w13033 & w20896);
assign w13041 = ~w13033 & w13039;
assign w13042 = w13040 & ~w13041;
assign w13043 = ~pi276 & pi413;
assign w13044 = pi529 & ~w13043;
assign w13045 = pi276 & ~pi413;
assign w13046 = w13044 & ~w13045;
assign w13047 = ~w13042 & ~w13046;
assign w13048 = w5893 & w8150;
assign w13049 = ~w5893 & ~w8150;
assign w13050 = ~w13048 & ~w13049;
assign w13051 = w5328 & w19477;
assign w13052 = (pi218 & ~w5328) | (pi218 & w19478) | (~w5328 & w19478);
assign w13053 = ~w13051 & ~w13052;
assign w13054 = ~w1527 & w13053;
assign w13055 = w1527 & ~w13053;
assign w13056 = ~w13054 & ~w13055;
assign w13057 = (~pi529 & ~w13050) | (~pi529 & w19479) | (~w13050 & w19479);
assign w13058 = ~w13050 & ~w13056;
assign w13059 = w13057 & ~w13058;
assign w13060 = pi218 & pi461;
assign w13061 = pi529 & ~w13060;
assign w13062 = ~pi218 & ~pi461;
assign w13063 = w13061 & ~w13062;
assign w13064 = ~w13059 & ~w13063;
assign w13065 = ~pi209 & w5554;
assign w13066 = pi209 & ~w5554;
assign w13067 = ~w13065 & ~w13066;
assign w13068 = w5396 & w13067;
assign w13069 = ~w5396 & ~w13067;
assign w13070 = ~w13068 & ~w13069;
assign w13071 = (~pi529 & w13070) | (~pi529 & w19480) | (w13070 & w19480);
assign w13072 = ~w11581 & w13070;
assign w13073 = w13071 & ~w13072;
assign w13074 = ~pi209 & pi435;
assign w13075 = pi529 & ~w13074;
assign w13076 = pi209 & ~pi435;
assign w13077 = w13075 & ~w13076;
assign w13078 = ~w13073 & ~w13077;
assign w13079 = w1443 & w5482;
assign w13080 = ~w1443 & ~w5482;
assign w13081 = ~w13079 & ~w13080;
assign w13082 = ~pi217 & w5554;
assign w13083 = pi217 & ~w5554;
assign w13084 = ~w13082 & ~w13083;
assign w13085 = ~w5329 & w13084;
assign w13086 = w5329 & ~w13084;
assign w13087 = ~w13085 & ~w13086;
assign w13088 = w13081 & ~w13087;
assign w13089 = ~pi529 & ~w13088;
assign w13090 = ~w13081 & w13087;
assign w13091 = w13089 & ~w13090;
assign w13092 = ~pi217 & pi499;
assign w13093 = pi529 & ~w13092;
assign w13094 = pi217 & ~pi499;
assign w13095 = w13093 & ~w13094;
assign w13096 = ~w13091 & ~w13095;
assign w13097 = ~w1367 & ~w5893;
assign w13098 = w1367 & w5893;
assign w13099 = ~w13097 & ~w13098;
assign w13100 = ~pi151 & w5554;
assign w13101 = pi151 & ~w5554;
assign w13102 = ~w13100 & ~w13101;
assign w13103 = ~w1527 & w13102;
assign w13104 = w1527 & ~w13102;
assign w13105 = ~w13103 & ~w13104;
assign w13106 = w13099 & ~w13105;
assign w13107 = ~pi529 & ~w13106;
assign w13108 = ~w13099 & w13105;
assign w13109 = w13107 & ~w13108;
assign w13110 = ~pi151 & pi408;
assign w13111 = pi529 & ~w13110;
assign w13112 = pi151 & ~pi408;
assign w13113 = w13111 & ~w13112;
assign w13114 = ~w13109 & ~w13113;
assign w13115 = ~pi208 & w9618;
assign w13116 = pi208 & ~w9618;
assign w13117 = ~w13115 & ~w13116;
assign w13118 = w12022 & w13117;
assign w13119 = ~w12022 & ~w13117;
assign w13120 = ~w13118 & ~w13119;
assign w13121 = (~pi529 & w13120) | (~pi529 & w19481) | (w13120 & w19481);
assign w13122 = ~w11941 & w13120;
assign w13123 = w13121 & ~w13122;
assign w13124 = ~pi208 & pi449;
assign w13125 = pi529 & ~w13124;
assign w13126 = pi208 & ~pi449;
assign w13127 = w13125 & ~w13126;
assign w13128 = ~w13123 & ~w13127;
assign w13129 = w2289 & w12100;
assign w13130 = ~w2289 & ~w12100;
assign w13131 = ~w13129 & ~w13130;
assign w13132 = ~w9617 & w20897;
assign w13133 = (pi346 & w9617) | (pi346 & w20898) | (w9617 & w20898);
assign w13134 = ~w13132 & ~w13133;
assign w13135 = ~w9551 & w13134;
assign w13136 = w9551 & ~w13134;
assign w13137 = ~w13135 & ~w13136;
assign w13138 = (~pi529 & ~w13131) | (~pi529 & w20899) | (~w13131 & w20899);
assign w13139 = ~w13131 & w13137;
assign w13140 = w13138 & ~w13139;
assign w13141 = ~pi346 & pi468;
assign w13142 = pi529 & ~w13141;
assign w13143 = pi346 & ~pi468;
assign w13144 = w13142 & ~w13143;
assign w13145 = ~w13140 & ~w13144;
assign w13146 = ~w1692 & ~w11753;
assign w13147 = w1692 & w11753;
assign w13148 = ~w13146 & ~w13147;
assign w13149 = ~pi375 & ~w12130;
assign w13150 = pi375 & w12130;
assign w13151 = ~w13149 & ~w13150;
assign w13152 = (~pi529 & ~w13151) | (~pi529 & w19482) | (~w13151 & w19482);
assign w13153 = ~w13148 & ~w13151;
assign w13154 = w13152 & ~w13153;
assign w13155 = ~pi375 & pi528;
assign w13156 = pi529 & ~w13155;
assign w13157 = pi375 & ~pi528;
assign w13158 = w13156 & ~w13157;
assign w13159 = ~w13154 & ~w13158;
assign w13160 = ~w6098 & w6530;
assign w13161 = w6098 & ~w6530;
assign w13162 = ~w13160 & ~w13161;
assign w13163 = ~pi210 & w10600;
assign w13164 = pi210 & ~w10600;
assign w13165 = ~w13163 & ~w13164;
assign w13166 = w13162 & w13165;
assign w13167 = ~w13162 & ~w13165;
assign w13168 = ~w13166 & ~w13167;
assign w13169 = (~pi529 & w13168) | (~pi529 & w19483) | (w13168 & w19483);
assign w13170 = ~w9918 & w13168;
assign w13171 = w13169 & ~w13170;
assign w13172 = ~pi210 & pi509;
assign w13173 = pi529 & ~w13172;
assign w13174 = pi210 & ~pi509;
assign w13175 = w13173 & ~w13174;
assign w13176 = ~w13171 & ~w13175;
assign w13177 = ~pi121 & pi130;
assign w13178 = pi121 & ~pi130;
assign w13179 = ~w13177 & ~w13178;
assign w13180 = pi232 & ~pi233;
assign w13181 = ~pi270 & w13180;
assign w13182 = ~pi215 & ~pi232;
assign w13183 = pi175 & pi233;
assign w13184 = w13182 & w13183;
assign w13185 = pi215 & ~pi233;
assign w13186 = pi232 & w13185;
assign w13187 = ~w13181 & ~w13184;
assign w13188 = (pi231 & ~w13187) | (pi231 & w14925) | (~w13187 & w14925);
assign w13189 = ~pi232 & pi233;
assign w13190 = ~pi175 & ~pi231;
assign w13191 = w13189 & w13190;
assign w13192 = pi215 & w13191;
assign w13193 = (~pi285 & ~w13191) | (~pi285 & w19484) | (~w13191 & w19484);
assign w13194 = pi175 & pi270;
assign w13195 = ~pi215 & w13194;
assign w13196 = w13189 & w13195;
assign w13197 = pi215 & ~pi232;
assign w13198 = pi175 & ~pi233;
assign w13199 = w13197 & w13198;
assign w13200 = ~pi175 & ~pi270;
assign w13201 = pi215 & pi232;
assign w13202 = w13200 & w13201;
assign w13203 = ~pi215 & ~pi233;
assign w13204 = w13200 & w13203;
assign w13205 = ~w13202 & ~w13204;
assign w13206 = ~pi231 & w13199;
assign w13207 = w13205 & ~w13206;
assign w13208 = w13193 & w13207;
assign w13209 = w13208 & w19485;
assign w13210 = ~pi175 & w13185;
assign w13211 = ~pi232 & w13203;
assign w13212 = (~pi231 & ~w13203) | (~pi231 & w19486) | (~w13203 & w19486);
assign w13213 = ~pi215 & pi232;
assign w13214 = pi270 & w13189;
assign w13215 = (pi231 & ~w13189) | (pi231 & w15594) | (~w13189 & w15594);
assign w13216 = ~w13198 & w13213;
assign w13217 = w13215 & ~w13216;
assign w13218 = ~w13210 & w13212;
assign w13219 = ~w13217 & ~w13218;
assign w13220 = pi270 & w13213;
assign w13221 = w13213 & w19487;
assign w13222 = w13183 & w13197;
assign w13223 = ~w13221 & ~w13222;
assign w13224 = pi232 & pi233;
assign w13225 = pi270 & w13224;
assign w13226 = w13224 & w13249;
assign w13227 = pi285 & ~w13226;
assign w13228 = w13223 & w13227;
assign w13229 = ~w13219 & w13228;
assign w13230 = w13189 & w13200;
assign w13231 = w13183 & w13201;
assign w13232 = ~w13230 & ~w13231;
assign w13233 = ~pi215 & w13226;
assign w13234 = w13232 & ~w13233;
assign w13235 = ~pi231 & ~w13234;
assign w13236 = pi231 & pi270;
assign w13237 = ~pi215 & pi233;
assign w13238 = ~w13185 & ~w13237;
assign w13239 = ~pi232 & ~w13238;
assign w13240 = pi233 & w13194;
assign w13241 = w13194 & w13237;
assign w13242 = (w13236 & w13239) | (w13236 & w19488) | (w13239 & w19488);
assign w13243 = pi175 & pi215;
assign w13244 = w13181 & w13243;
assign w13245 = ~w13242 & ~w13244;
assign w13246 = ~w13235 & w13245;
assign w13247 = ~w13209 & ~w13229;
assign w13248 = ~pi233 & ~pi270;
assign w13249 = ~pi175 & pi270;
assign w13250 = w13201 & w13249;
assign w13251 = ~pi233 & w13250;
assign w13252 = (pi231 & w13251) | (pi231 & w19489) | (w13251 & w19489);
assign w13253 = pi233 & w13201;
assign w13254 = w13194 & w13253;
assign w13255 = pi233 & ~pi270;
assign w13256 = ~pi231 & w13255;
assign w13257 = w13200 & w13253;
assign w13258 = w13213 & w13256;
assign w13259 = ~w13257 & ~w13258;
assign w13260 = pi285 & ~w13184;
assign w13261 = ~w13254 & w13260;
assign w13262 = w13259 & w13261;
assign w13263 = ~pi231 & w13221;
assign w13264 = w13221 & w13296;
assign w13265 = ~pi175 & pi231;
assign w13266 = ~pi232 & pi270;
assign w13267 = ~w13236 & ~w13266;
assign w13268 = w13203 & ~w13267;
assign w13269 = ~pi285 & ~w13230;
assign w13270 = ~w13268 & w13269;
assign w13271 = ~w13182 & w13265;
assign w13272 = pi233 & w13271;
assign w13273 = ~w13252 & w13262;
assign w13274 = w13270 & w19490;
assign w13275 = ~w13273 & ~w13274;
assign w13276 = w13248 & w19491;
assign w13277 = w13201 & w13255;
assign w13278 = ~w13276 & ~w13277;
assign w13279 = ~pi232 & w13185;
assign w13280 = pi233 & w13250;
assign w13281 = ~pi233 & pi270;
assign w13282 = w13243 & w13281;
assign w13283 = ~w13280 & ~w13282;
assign w13284 = w13200 & w13279;
assign w13285 = (~pi231 & w13280) | (~pi231 & w19492) | (w13280 & w19492);
assign w13286 = ~w13284 & ~w13285;
assign w13287 = (~pi234 & w13275) | (~pi234 & w19493) | (w13275 & w19493);
assign w13288 = pi231 & ~w13223;
assign w13289 = w13213 & w13255;
assign w13290 = pi270 & w13182;
assign w13291 = pi215 & w13248;
assign w13292 = ~w13290 & ~w13291;
assign w13293 = (w13190 & ~w13292) | (w13190 & w19494) | (~w13292 & w19494);
assign w13294 = pi175 & pi231;
assign w13295 = ~pi270 & w13294;
assign w13296 = pi175 & ~pi231;
assign w13297 = w13237 & w19495;
assign w13298 = w13296 & w13297;
assign w13299 = w13201 & w13295;
assign w13300 = ~w13298 & ~w13299;
assign w13301 = ~w13288 & ~w13293;
assign w13302 = (pi285 & ~w13301) | (pi285 & w19496) | (~w13301 & w19496);
assign w13303 = pi231 & ~pi285;
assign w13304 = w13248 & w13265;
assign w13305 = w13197 & w13304;
assign w13306 = w13211 & w13249;
assign w13307 = ~w13305 & ~w13306;
assign w13308 = w13303 & ~w13307;
assign w13309 = pi231 & w13222;
assign w13310 = pi215 & pi233;
assign w13311 = w13296 & w13310;
assign w13312 = ~pi285 & w13311;
assign w13313 = ~w13309 & ~w13312;
assign w13314 = ~pi270 & ~w13313;
assign w13315 = w13185 & w13266;
assign w13316 = pi175 & w13315;
assign w13317 = w13214 & w13294;
assign w13318 = w13214 & w19497;
assign w13319 = ~w13308 & ~w13314;
assign w13320 = ~w13316 & ~w13318;
assign w13321 = w13319 & w13320;
assign w13322 = ~w13302 & w13321;
assign w13323 = ~w13287 & w13322;
assign w13324 = (pi234 & w13247) | (pi234 & w19498) | (w13247 & w19498);
assign w13325 = w13323 & w19499;
assign w13326 = (pi131 & ~w13323) | (pi131 & w19500) | (~w13323 & w19500);
assign w13327 = ~w13325 & ~w13326;
assign w13328 = ~w13179 & ~w13327;
assign w13329 = w13179 & w13327;
assign w13330 = pi532 & pi584;
assign w13331 = ~w13328 & ~w13329;
assign w13332 = ~pi532 & w13331;
assign w13333 = ~w13330 & ~w13332;
assign w13334 = w3202 & w12292;
assign w13335 = ~w3202 & ~w12292;
assign w13336 = ~w13334 & ~w13335;
assign w13337 = ~pi371 & ~w13162;
assign w13338 = pi371 & w13162;
assign w13339 = ~w13337 & ~w13338;
assign w13340 = w13336 & w13339;
assign w13341 = ~pi529 & ~w13340;
assign w13342 = ~w13336 & ~w13339;
assign w13343 = w13341 & ~w13342;
assign w13344 = ~pi371 & pi501;
assign w13345 = pi529 & ~w13344;
assign w13346 = pi371 & ~pi501;
assign w13347 = w13345 & ~w13346;
assign w13348 = ~w13343 & ~w13347;
assign w13349 = ~w4440 & ~w7918;
assign w13350 = w4440 & w7918;
assign w13351 = ~w13349 & ~w13350;
assign w13352 = ~pi351 & w7123;
assign w13353 = pi351 & ~w7123;
assign w13354 = ~w13352 & ~w13353;
assign w13355 = ~w8232 & w13354;
assign w13356 = w8232 & ~w13354;
assign w13357 = ~w13355 & ~w13356;
assign w13358 = w13351 & ~w13357;
assign w13359 = ~pi529 & ~w13358;
assign w13360 = ~w13351 & w13357;
assign w13361 = w13359 & ~w13360;
assign w13362 = ~pi351 & pi404;
assign w13363 = pi529 & ~w13362;
assign w13364 = pi351 & ~pi404;
assign w13365 = w13363 & ~w13364;
assign w13366 = ~w13361 & ~w13365;
assign w13367 = w1131 & w11527;
assign w13368 = ~w1131 & ~w11527;
assign w13369 = ~w13367 & ~w13368;
assign w13370 = w7512 & w19501;
assign w13371 = (pi258 & ~w7512) | (pi258 & w19502) | (~w7512 & w19502);
assign w13372 = ~w13370 & ~w13371;
assign w13373 = ~w145 & w13372;
assign w13374 = w145 & ~w13372;
assign w13375 = ~w13373 & ~w13374;
assign w13376 = (~pi529 & ~w13369) | (~pi529 & w19503) | (~w13369 & w19503);
assign w13377 = ~w13369 & w13375;
assign w13378 = w13376 & ~w13377;
assign w13379 = ~pi258 & pi431;
assign w13380 = pi529 & ~w13379;
assign w13381 = pi258 & ~pi431;
assign w13382 = w13380 & ~w13381;
assign w13383 = ~w13378 & ~w13382;
assign w13384 = ~w1021 & w5152;
assign w13385 = w1021 & ~w5152;
assign w13386 = ~w13384 & ~w13385;
assign w13387 = w554 & w13386;
assign w13388 = ~w554 & ~w13386;
assign w13389 = ~w13387 & ~w13388;
assign w13390 = ~pi183 & w5243;
assign w13391 = pi183 & ~w5243;
assign w13392 = ~w13390 & ~w13391;
assign w13393 = w811 & w13392;
assign w13394 = ~w811 & ~w13392;
assign w13395 = ~w13393 & ~w13394;
assign w13396 = w13389 & w13395;
assign w13397 = ~pi529 & ~w13396;
assign w13398 = ~w13389 & ~w13395;
assign w13399 = w13397 & ~w13398;
assign w13400 = ~pi183 & pi480;
assign w13401 = pi529 & ~w13400;
assign w13402 = pi183 & ~pi480;
assign w13403 = w13401 & ~w13402;
assign w13404 = ~w13399 & ~w13403;
assign w13405 = w1844 & w11884;
assign w13406 = ~w1844 & ~w11884;
assign w13407 = ~w13405 & ~w13406;
assign w13408 = w11809 & w19504;
assign w13409 = (pi348 & ~w11809) | (pi348 & w19505) | (~w11809 & w19505);
assign w13410 = ~w13408 & ~w13409;
assign w13411 = ~w8456 & w13410;
assign w13412 = w8456 & ~w13410;
assign w13413 = ~w13411 & ~w13412;
assign w13414 = (~pi529 & ~w13407) | (~pi529 & w19506) | (~w13407 & w19506);
assign w13415 = ~w13407 & w13413;
assign w13416 = w13414 & ~w13415;
assign w13417 = ~pi348 & pi526;
assign w13418 = pi529 & ~w13417;
assign w13419 = pi348 & ~pi526;
assign w13420 = w13418 & ~w13419;
assign w13421 = ~w13416 & ~w13420;
assign w13422 = ~w1692 & w9069;
assign w13423 = w1692 & ~w9069;
assign w13424 = ~w13422 & ~w13423;
assign w13425 = w8719 & w13424;
assign w13426 = ~w8719 & ~w13424;
assign w13427 = ~w13425 & ~w13426;
assign w13428 = ~pi320 & w9148;
assign w13429 = pi320 & ~w9148;
assign w13430 = ~w13428 & ~w13429;
assign w13431 = w8812 & w13430;
assign w13432 = ~w8812 & ~w13430;
assign w13433 = ~w13431 & ~w13432;
assign w13434 = (~pi529 & ~w13433) | (~pi529 & w19507) | (~w13433 & w19507);
assign w13435 = ~w13427 & ~w13433;
assign w13436 = w13434 & ~w13435;
assign w13437 = ~pi320 & pi406;
assign w13438 = pi529 & ~w13437;
assign w13439 = pi320 & ~pi406;
assign w13440 = w13438 & ~w13439;
assign w13441 = ~w13436 & ~w13440;
assign w13442 = w1844 & w11750;
assign w13443 = ~w1844 & ~w11750;
assign w13444 = ~w13442 & ~w13443;
assign w13445 = w5777 & w19508;
assign w13446 = (pi228 & ~w5777) | (pi228 & w19509) | (~w5777 & w19509);
assign w13447 = ~w13445 & ~w13446;
assign w13448 = ~w11810 & w13447;
assign w13449 = w11810 & ~w13447;
assign w13450 = ~w13448 & ~w13449;
assign w13451 = (~pi529 & ~w13444) | (~pi529 & w20900) | (~w13444 & w20900);
assign w13452 = ~w13444 & w13450;
assign w13453 = w13451 & ~w13452;
assign w13454 = ~pi228 & pi466;
assign w13455 = pi529 & ~w13454;
assign w13456 = pi228 & ~pi466;
assign w13457 = w13455 & ~w13456;
assign w13458 = ~w13453 & ~w13457;
assign w13459 = pi275 & ~pi354;
assign w13460 = pi157 & w13459;
assign w13461 = w13459 & w19510;
assign w13462 = ~pi284 & ~w13461;
assign w13463 = w13459 & w19511;
assign w13464 = ~pi157 & ~pi275;
assign w13465 = pi132 & pi354;
assign w13466 = w13464 & w13465;
assign w13467 = ~pi351 & w13466;
assign w13468 = ~w13463 & ~w13467;
assign w13469 = w13462 & w13468;
assign w13470 = pi157 & pi354;
assign w13471 = pi358 & w13470;
assign w13472 = w13470 & w13550;
assign w13473 = pi275 & w13472;
assign w13474 = pi275 & ~pi358;
assign w13475 = ~pi157 & w13474;
assign w13476 = ~pi275 & ~pi354;
assign w13477 = pi132 & pi358;
assign w13478 = w13476 & w13477;
assign w13479 = ~w13475 & ~w13478;
assign w13480 = pi351 & ~w13479;
assign w13481 = ~pi275 & pi354;
assign w13482 = pi132 & w13481;
assign w13483 = w13481 & w13502;
assign w13484 = pi157 & ~pi354;
assign w13485 = w13477 & w13484;
assign w13486 = ~pi275 & w13485;
assign w13487 = ~w13486 & w19512;
assign w13488 = ~pi132 & w13476;
assign w13489 = w13476 & w19513;
assign w13490 = pi358 & w13489;
assign w13491 = ~pi275 & w13472;
assign w13492 = ~w13490 & ~w13491;
assign w13493 = w13487 & w13492;
assign w13494 = ~w13473 & ~w13480;
assign w13495 = w13469 & w13494;
assign w13496 = ~w13493 & ~w13495;
assign w13497 = pi132 & ~pi354;
assign w13498 = w13474 & w13497;
assign w13499 = ~w13463 & ~w13498;
assign w13500 = ~pi358 & w13484;
assign w13501 = (~pi351 & ~w13499) | (~pi351 & w19514) | (~w13499 & w19514);
assign w13502 = pi132 & ~pi358;
assign w13503 = ~pi157 & pi354;
assign w13504 = pi358 & w13503;
assign w13505 = ~pi157 & ~w13474;
assign w13506 = pi157 & w13502;
assign w13507 = ~w13504 & w13505;
assign w13508 = pi284 & ~pi351;
assign w13509 = ~pi132 & pi351;
assign w13510 = ~pi354 & ~pi358;
assign w13511 = ~pi157 & w13510;
assign w13512 = ~w13471 & ~w13511;
assign w13513 = w13509 & ~w13512;
assign w13514 = pi275 & pi354;
assign w13515 = ~pi157 & w13514;
assign w13516 = w13514 & w19515;
assign w13517 = ~pi351 & w13516;
assign w13518 = w13460 & w13502;
assign w13519 = ~w13517 & ~w13518;
assign w13520 = ~w13512 & w19516;
assign w13521 = w13519 & ~w13520;
assign w13522 = (w13508 & w13507) | (w13508 & w19517) | (w13507 & w19517);
assign w13523 = ~w13496 & w19518;
assign w13524 = pi193 & ~w13523;
assign w13525 = pi157 & w13481;
assign w13526 = w13481 & w19519;
assign w13527 = ~pi351 & w13526;
assign w13528 = pi157 & pi275;
assign w13529 = pi358 & w13528;
assign w13530 = ~pi358 & w13476;
assign w13531 = w13476 & w13502;
assign w13532 = w13528 & w19520;
assign w13533 = ~w13531 & ~w13532;
assign w13534 = ~pi157 & w13502;
assign w13535 = ~pi132 & w13459;
assign w13536 = ~w13534 & ~w13535;
assign w13537 = ~w13533 & ~w13536;
assign w13538 = (pi284 & w13537) | (pi284 & w19521) | (w13537 & w19521);
assign w13539 = pi157 & w13476;
assign w13540 = w13539 & w19522;
assign w13541 = pi132 & pi351;
assign w13542 = w13539 & w13541;
assign w13543 = w13539 & w19523;
assign w13544 = ~pi132 & ~pi351;
assign w13545 = w13503 & w13544;
assign w13546 = pi275 & w13545;
assign w13547 = ~w13540 & ~w13543;
assign w13548 = ~w13546 & w13547;
assign w13549 = ~w13538 & w13548;
assign w13550 = ~pi132 & pi358;
assign w13551 = ~pi157 & ~w13550;
assign w13552 = ~pi275 & w13477;
assign w13553 = w13503 & w19524;
assign w13554 = ~pi157 & pi275;
assign w13555 = ~pi354 & pi358;
assign w13556 = w13554 & w13555;
assign w13557 = ~w13553 & ~w13556;
assign w13558 = (~w13551 & ~w13557) | (~w13551 & w19525) | (~w13557 & w19525);
assign w13559 = (pi351 & w13558) | (pi351 & w19526) | (w13558 & w19526);
assign w13560 = ~pi358 & w13470;
assign w13561 = w13544 & w13560;
assign w13562 = pi132 & ~pi351;
assign w13563 = w13528 & w13555;
assign w13564 = w13562 & w13563;
assign w13565 = ~pi132 & ~pi358;
assign w13566 = w13476 & w13565;
assign w13567 = ~w13561 & ~w13564;
assign w13568 = w13567 & w19527;
assign w13569 = ~w13559 & w13568;
assign w13570 = ~pi284 & ~w13569;
assign w13571 = pi157 & ~pi275;
assign w13572 = w13550 & w13571;
assign w13573 = ~pi351 & ~w13572;
assign w13574 = w13459 & w13565;
assign w13575 = ~w13482 & ~w13574;
assign w13576 = pi351 & ~w13563;
assign w13577 = w13573 & w13575;
assign w13578 = ~w13576 & ~w13577;
assign w13579 = w13528 & w13565;
assign w13580 = ~pi354 & w13579;
assign w13581 = w13464 & w13497;
assign w13582 = ~w13477 & ~w13541;
assign w13583 = w13470 & ~w13582;
assign w13584 = w13514 & w19513;
assign w13585 = w13470 & w19528;
assign w13586 = ~w13583 & w19529;
assign w13587 = pi284 & ~w13581;
assign w13588 = ~w13580 & w13587;
assign w13589 = w13586 & w13588;
assign w13590 = ~pi157 & w13476;
assign w13591 = w13476 & w19530;
assign w13592 = pi354 & ~pi358;
assign w13593 = w13528 & w13592;
assign w13594 = ~w13553 & ~w13591;
assign w13595 = (~pi132 & ~w13594) | (~pi132 & w19531) | (~w13594 & w19531);
assign w13596 = ~pi358 & w13541;
assign w13597 = w13541 & w19528;
assign w13598 = (~pi284 & ~w13597) | (~pi284 & w19532) | (~w13597 & w19532);
assign w13599 = ~w13578 & w13589;
assign w13600 = ~w13595 & w13598;
assign w13601 = ~w13599 & ~w13600;
assign w13602 = w13464 & w13510;
assign w13603 = ~pi351 & ~w13526;
assign w13604 = w13497 & w19515;
assign w13605 = w13474 & w13503;
assign w13606 = ~w13604 & ~w13605;
assign w13607 = ~pi157 & w13459;
assign w13608 = pi354 & w13477;
assign w13609 = ~w13607 & ~w13608;
assign w13610 = w13497 & w19533;
assign w13611 = pi351 & ~w13530;
assign w13612 = ~w13610 & w13611;
assign w13613 = ~w13551 & ~w13609;
assign w13614 = w13612 & ~w13613;
assign w13615 = w13603 & w13606;
assign w13616 = (~w13602 & w13614) | (~w13602 & w19534) | (w13614 & w19534);
assign w13617 = (~pi193 & w13601) | (~pi193 & w19535) | (w13601 & w19535);
assign w13618 = ~w13524 & ~w13570;
assign w13619 = w13618 & w19536;
assign w13620 = (pi388 & ~w13618) | (pi388 & w19537) | (~w13618 & w19537);
assign w13621 = ~w13619 & ~w13620;
assign w13622 = ~pi140 & pi141;
assign w13623 = pi140 & ~pi141;
assign w13624 = ~w13622 & ~w13623;
assign w13625 = ~pi129 & pi144;
assign w13626 = pi129 & ~pi144;
assign w13627 = ~w13625 & ~w13626;
assign w13628 = w13624 & w13627;
assign w13629 = ~w13624 & ~w13627;
assign w13630 = ~w13628 & ~w13629;
assign w13631 = w13621 & ~w13630;
assign w13632 = ~w13621 & w13630;
assign w13633 = pi532 & pi562;
assign w13634 = ~w13631 & ~w13632;
assign w13635 = ~pi532 & w13634;
assign w13636 = ~w13633 & ~w13635;
assign w13637 = w13323 & w19538;
assign w13638 = (pi130 & ~w13323) | (pi130 & w19539) | (~w13323 & w19539);
assign w13639 = ~w13637 & ~w13638;
assign w13640 = pi532 & ~pi648;
assign w13641 = ~pi532 & ~w13639;
assign w13642 = ~w13640 & ~w13641;
assign w13643 = pi131 & ~w13639;
assign w13644 = ~pi131 & w13639;
assign w13645 = pi532 & pi616;
assign w13646 = ~w13643 & ~w13644;
assign w13647 = ~pi532 & w13646;
assign w13648 = ~w13645 & ~w13647;
assign w13649 = ~pi131 & pi132;
assign w13650 = pi131 & ~pi132;
assign w13651 = ~w13649 & ~w13650;
assign w13652 = w13179 & w13651;
assign w13653 = ~w13179 & ~w13651;
assign w13654 = ~w13652 & ~w13653;
assign w13655 = (~w13654 & ~w13323) | (~w13654 & w19540) | (~w13323 & w19540);
assign w13656 = w13323 & w19541;
assign w13657 = pi532 & pi552;
assign w13658 = ~w13655 & ~w13656;
assign w13659 = ~pi532 & w13658;
assign w13660 = ~w13657 & ~w13659;
assign w13661 = ~pi133 & pi148;
assign w13662 = pi133 & ~pi148;
assign w13663 = ~w13661 & ~w13662;
assign w13664 = w13203 & w19542;
assign w13665 = w13189 & w19543;
assign w13666 = ~w13664 & ~w13665;
assign w13667 = (~pi175 & ~w13666) | (~pi175 & w19544) | (~w13666 & w19544);
assign w13668 = w13185 & w13200;
assign w13669 = w13213 & w13249;
assign w13670 = pi175 & w13237;
assign w13671 = ~w13668 & ~w13669;
assign w13672 = (~pi231 & ~w13671) | (~pi231 & w19545) | (~w13671 & w19545);
assign w13673 = w13186 & w13236;
assign w13674 = ~w13194 & ~w13294;
assign w13675 = w13224 & ~w13674;
assign w13676 = w13203 & w19491;
assign w13677 = w13185 & w19546;
assign w13678 = ~pi270 & w13677;
assign w13679 = ~pi232 & w13310;
assign w13680 = w13310 & w19547;
assign w13681 = ~w13289 & ~w13680;
assign w13682 = ~w13678 & w13681;
assign w13683 = ~w13673 & ~w13675;
assign w13684 = ~w13676 & w13683;
assign w13685 = w13684 & w19548;
assign w13686 = pi285 & ~w13685;
assign w13687 = ~pi232 & ~w13249;
assign w13688 = ~w13240 & ~w13279;
assign w13689 = ~w13687 & ~w13688;
assign w13690 = ~pi270 & w13203;
assign w13691 = ~w13276 & ~w13690;
assign w13692 = (pi231 & w13689) | (pi231 & w19549) | (w13689 & w19549);
assign w13693 = w13182 & w13248;
assign w13694 = ~w13263 & ~w13693;
assign w13695 = w13197 & w13255;
assign w13696 = w13198 & w13266;
assign w13697 = ~w13695 & ~w13696;
assign w13698 = ~pi231 & ~w13697;
assign w13699 = w13694 & ~w13698;
assign w13700 = ~w13692 & w13699;
assign w13701 = ~w13686 & w13700;
assign w13702 = pi270 & w13201;
assign w13703 = w13198 & w13702;
assign w13704 = w13266 & w13310;
assign w13705 = ~pi231 & ~w13704;
assign w13706 = w13200 & w13224;
assign w13707 = w13705 & ~w13706;
assign w13708 = (~w13687 & w13239) | (~w13687 & w19551) | (w13239 & w19551);
assign w13709 = pi231 & ~w13280;
assign w13710 = ~w13708 & w13709;
assign w13711 = ~w13703 & w13707;
assign w13712 = ~w13710 & ~w13711;
assign w13713 = (~pi285 & w13712) | (~pi285 & w19552) | (w13712 & w19552);
assign w13714 = (~pi231 & ~w13185) | (~pi231 & w20901) | (~w13185 & w20901);
assign w13715 = ~pi270 & w13197;
assign w13716 = w13194 & w13203;
assign w13717 = ~w13715 & ~w13716;
assign w13718 = ~w13184 & w13714;
assign w13719 = pi231 & w13717;
assign w13720 = ~w13718 & ~w13719;
assign w13721 = w13180 & w13243;
assign w13722 = ~pi285 & ~w13721;
assign w13723 = ~w13280 & w13722;
assign w13724 = ~w13720 & w13723;
assign w13725 = w13180 & w13195;
assign w13726 = ~w13233 & ~w13725;
assign w13727 = w13237 & w13745;
assign w13728 = ~w13306 & w19553;
assign w13729 = w13726 & w13728;
assign w13730 = pi215 & ~pi270;
assign w13731 = w13198 & w13730;
assign w13732 = ~w13721 & ~w13731;
assign w13733 = ~w13181 & ~w13704;
assign w13734 = w13732 & w13733;
assign w13735 = ~pi231 & ~w13734;
assign w13736 = w13197 & w13248;
assign w13737 = w13201 & w19487;
assign w13738 = ~w13736 & ~w13737;
assign w13739 = w13265 & ~w13738;
assign w13740 = ~pi232 & ~w13730;
assign w13741 = ~pi231 & pi285;
assign w13742 = ~w13214 & w13740;
assign w13743 = w13741 & w13742;
assign w13744 = ~w13185 & ~w13741;
assign w13745 = pi175 & ~pi270;
assign w13746 = pi232 & w13745;
assign w13747 = ~w13744 & w13746;
assign w13748 = ~w13743 & ~w13747;
assign w13749 = ~w13735 & ~w13739;
assign w13750 = w13748 & w13749;
assign w13751 = ~w13724 & ~w13729;
assign w13752 = w13750 & ~w13751;
assign w13753 = w13250 & w19554;
assign w13754 = ~w13725 & ~w13753;
assign w13755 = w13213 & w13745;
assign w13756 = ~pi233 & w13755;
assign w13757 = w13755 & w19555;
assign w13758 = ~w13192 & ~w13757;
assign w13759 = pi231 & ~w13754;
assign w13760 = pi285 & ~w13200;
assign w13761 = (w13760 & w13263) | (w13760 & w19556) | (w13263 & w19556);
assign w13762 = ~w13759 & w19557;
assign w13763 = (w13762 & w13752) | (w13762 & w19558) | (w13752 & w19558);
assign w13764 = ~w13713 & w13763;
assign w13765 = (~pi234 & ~w13701) | (~pi234 & w19559) | (~w13701 & w19559);
assign w13766 = w13764 & w19560;
assign w13767 = (pi149 & ~w13764) | (pi149 & w19561) | (~w13764 & w19561);
assign w13768 = ~w13766 & ~w13767;
assign w13769 = ~w13663 & ~w13768;
assign w13770 = w13663 & w13768;
assign w13771 = pi532 & pi586;
assign w13772 = ~w13769 & ~w13770;
assign w13773 = ~pi532 & w13772;
assign w13774 = ~w13771 & ~w13773;
assign w13775 = pi275 & w13550;
assign w13776 = w13484 & w13775;
assign w13777 = pi132 & w13514;
assign w13778 = w13514 & w19511;
assign w13779 = pi358 & w13778;
assign w13780 = ~pi132 & w13592;
assign w13781 = w13528 & w13780;
assign w13782 = ~w13466 & ~w13781;
assign w13783 = ~pi351 & w13585;
assign w13784 = w13782 & w19563;
assign w13785 = pi132 & w13527;
assign w13786 = ~pi132 & pi354;
assign w13787 = w13476 & w19519;
assign w13788 = ~w13464 & w13786;
assign w13789 = ~w13787 & ~w13788;
assign w13790 = pi351 & ~w13789;
assign w13791 = pi358 & w13464;
assign w13792 = w13464 & w13555;
assign w13793 = w13592 & w19513;
assign w13794 = ~w13785 & ~w13790;
assign w13795 = ~w13792 & ~w13793;
assign w13796 = pi358 & w13459;
assign w13797 = w13459 & w13477;
assign w13798 = ~w13473 & ~w13797;
assign w13799 = w13565 & w13607;
assign w13800 = ~w13593 & ~w13610;
assign w13801 = pi351 & ~w13800;
assign w13802 = ~w13799 & ~w13801;
assign w13803 = (~pi351 & w13473) | (~pi351 & w19565) | (w13473 & w19565);
assign w13804 = w13802 & ~w13803;
assign w13805 = (~pi284 & ~w13794) | (~pi284 & w19566) | (~w13794 & w19566);
assign w13806 = w13804 & ~w13805;
assign w13807 = pi351 & ~w13504;
assign w13808 = ~w13497 & w13571;
assign w13809 = w13807 & ~w13808;
assign w13810 = ~w13535 & ~w13590;
assign w13811 = ~pi351 & w13810;
assign w13812 = ~w13809 & ~w13811;
assign w13813 = w13465 & w13554;
assign w13814 = ~w13526 & ~w13813;
assign w13815 = pi284 & ~w13472;
assign w13816 = w13814 & w13815;
assign w13817 = ~w13812 & w13816;
assign w13818 = w13465 & w13791;
assign w13819 = ~w13460 & ~w13466;
assign w13820 = ~w13500 & w13819;
assign w13821 = (~pi351 & ~w13791) | (~pi351 & w19568) | (~w13791 & w19568);
assign w13822 = ~w13820 & ~w13821;
assign w13823 = ~pi157 & w13562;
assign w13824 = w13459 & w13823;
assign w13825 = ~w13546 & ~w13824;
assign w13826 = ~w13566 & ~w13579;
assign w13827 = ~pi284 & w13826;
assign w13828 = w13825 & w13827;
assign w13829 = ~w13822 & w13828;
assign w13830 = ~w13817 & ~w13829;
assign w13831 = w13477 & w13481;
assign w13832 = ~w13778 & ~w13793;
assign w13833 = ~pi351 & w13832;
assign w13834 = pi351 & ~w13831;
assign w13835 = w13557 & w13834;
assign w13836 = ~w13833 & ~w13835;
assign w13837 = w13526 & w13544;
assign w13838 = ~w13518 & ~w13837;
assign w13839 = (pi193 & w13830) | (pi193 & w19569) | (w13830 & w19569);
assign w13840 = pi351 & ~w13814;
assign w13841 = ~pi358 & w13459;
assign w13842 = ~w13791 & ~w13841;
assign w13843 = (w13544 & ~w13842) | (w13544 & w19570) | (~w13842 & w19570);
assign w13844 = w13466 & w20461;
assign w13845 = w13528 & w13596;
assign w13846 = ~w13844 & ~w13845;
assign w13847 = ~w13840 & ~w13843;
assign w13848 = w13846 & w13847;
assign w13849 = pi284 & ~w13848;
assign w13850 = ~pi284 & pi351;
assign w13851 = ~w13490 & ~w13799;
assign w13852 = w13850 & ~w13851;
assign w13853 = ~pi284 & w13562;
assign w13854 = w13515 & w13541;
assign w13855 = w13465 & w13474;
assign w13856 = (w13855 & w13854) | (w13855 & w19571) | (w13854 & w19571);
assign w13857 = w13504 & w13541;
assign w13858 = w13504 & w19572;
assign w13859 = ~pi157 & w13797;
assign w13860 = ~w13858 & ~w13859;
assign w13861 = ~w13856 & w13860;
assign w13862 = ~w13852 & w13861;
assign w13863 = ~w13849 & w13862;
assign w13864 = ~w13839 & w13863;
assign w13865 = w13864 & w19573;
assign w13866 = (pi386 & ~w13864) | (pi386 & w19574) | (~w13864 & w19574);
assign w13867 = ~w13865 & ~w13866;
assign w13868 = ~pi134 & ~w13867;
assign w13869 = pi134 & w13867;
assign w13870 = pi532 & pi656;
assign w13871 = ~w13868 & ~w13869;
assign w13872 = ~pi532 & w13871;
assign w13873 = ~w13870 & ~w13872;
assign w13874 = ~pi134 & pi135;
assign w13875 = pi134 & ~pi135;
assign w13876 = ~w13874 & ~w13875;
assign w13877 = ~w13867 & ~w13876;
assign w13878 = w13867 & w13876;
assign w13879 = pi532 & pi624;
assign w13880 = ~w13877 & ~w13878;
assign w13881 = ~pi532 & w13880;
assign w13882 = ~w13879 & ~w13881;
assign w13883 = ~pi134 & pi136;
assign w13884 = pi134 & ~pi136;
assign w13885 = ~w13883 & ~w13884;
assign w13886 = ~pi386 & ~w13885;
assign w13887 = pi386 & w13885;
assign w13888 = ~w13886 & ~w13887;
assign w13889 = w13864 & w19575;
assign w13890 = (pi135 & ~w13864) | (pi135 & w19576) | (~w13864 & w19576);
assign w13891 = ~w13889 & ~w13890;
assign w13892 = ~w13888 & ~w13891;
assign w13893 = w13888 & w13891;
assign w13894 = pi532 & pi592;
assign w13895 = ~w13892 & ~w13893;
assign w13896 = ~pi532 & w13895;
assign w13897 = ~w13894 & ~w13896;
assign w13898 = ~pi137 & pi171;
assign w13899 = pi137 & ~pi171;
assign w13900 = ~w13898 & ~w13899;
assign w13901 = ~pi172 & ~w13900;
assign w13902 = pi172 & w13900;
assign w13903 = ~w13901 & ~w13902;
assign w13904 = pi182 & pi342;
assign w13905 = pi170 & pi276;
assign w13906 = pi170 & ~pi276;
assign w13907 = pi321 & w13906;
assign w13908 = w13906 & w14008;
assign w13909 = pi342 & w13908;
assign w13910 = w13904 & w13905;
assign w13911 = ~pi170 & pi342;
assign w13912 = ~pi182 & ~pi321;
assign w13913 = w13911 & w13912;
assign w13914 = ~w13909 & w19577;
assign w13915 = ~pi352 & ~w13914;
assign w13916 = ~pi276 & ~pi342;
assign w13917 = ~pi170 & w13916;
assign w13918 = ~pi182 & ~pi342;
assign w13919 = pi276 & w13918;
assign w13920 = ~w13917 & ~w13919;
assign w13921 = ~pi352 & w13920;
assign w13922 = pi321 & w13911;
assign w13923 = pi182 & ~pi342;
assign w13924 = w13906 & ~w13923;
assign w13925 = pi352 & ~w13924;
assign w13926 = ~w13922 & w13925;
assign w13927 = ~w13921 & ~w13926;
assign w13928 = pi321 & pi342;
assign w13929 = w13906 & w13928;
assign w13930 = ~pi170 & pi276;
assign w13931 = w13904 & w13930;
assign w13932 = ~w13929 & ~w13931;
assign w13933 = pi170 & pi342;
assign w13934 = pi321 & w13933;
assign w13935 = w13933 & w14008;
assign w13936 = w13932 & w19578;
assign w13937 = ~w13927 & w13936;
assign w13938 = ~pi182 & ~pi352;
assign w13939 = w13911 & w13938;
assign w13940 = pi276 & w13939;
assign w13941 = w13923 & w13930;
assign w13942 = w13912 & w13916;
assign w13943 = ~pi372 & ~w13942;
assign w13944 = ~pi352 & w13941;
assign w13945 = w13943 & ~w13944;
assign w13946 = ~pi276 & pi342;
assign w13947 = pi182 & pi321;
assign w13948 = w13946 & w13947;
assign w13949 = ~pi352 & ~w13948;
assign w13950 = pi170 & ~pi342;
assign w13951 = ~pi321 & w13950;
assign w13952 = pi182 & ~pi276;
assign w13953 = w13911 & w13952;
assign w13954 = ~w13951 & ~w13953;
assign w13955 = ~w13949 & ~w13954;
assign w13956 = pi276 & ~pi342;
assign w13957 = pi170 & w13956;
assign w13958 = w13956 & w19579;
assign w13959 = w13905 & w13912;
assign w13960 = ~w13958 & ~w13959;
assign w13961 = ~w13955 & w13960;
assign w13962 = ~w13940 & w13945;
assign w13963 = w13961 & w13962;
assign w13964 = ~w13937 & ~w13963;
assign w13965 = pi321 & pi352;
assign w13966 = ~pi342 & w13930;
assign w13967 = ~pi170 & w13946;
assign w13968 = ~w13966 & ~w13967;
assign w13969 = (w13965 & ~w13968) | (w13965 & w19580) | (~w13968 & w19580);
assign w13970 = w13905 & w13923;
assign w13971 = ~pi321 & w13970;
assign w13972 = (pi191 & ~w13970) | (pi191 & w19581) | (~w13970 & w19581);
assign w13973 = ~w13969 & w13972;
assign w13974 = w13916 & w13965;
assign w13975 = w13916 & w19582;
assign w13976 = pi321 & ~pi352;
assign w13977 = w13933 & w13952;
assign w13978 = w13976 & w13977;
assign w13979 = ~pi182 & pi352;
assign w13980 = ~pi170 & ~pi276;
assign w13981 = w13979 & ~w13980;
assign w13982 = pi342 & w13981;
assign w13983 = ~w13975 & ~w13978;
assign w13984 = ~w13982 & w13983;
assign w13985 = ~w13913 & ~w13974;
assign w13986 = ~pi372 & w13985;
assign w13987 = w13984 & w13986;
assign w13988 = ~pi170 & ~pi342;
assign w13989 = ~pi321 & w13988;
assign w13990 = pi321 & w13918;
assign w13991 = w13905 & w13990;
assign w13992 = (pi352 & w13991) | (pi352 & w19583) | (w13991 & w19583);
assign w13993 = ~pi321 & w13933;
assign w13994 = w13933 & w19584;
assign w13995 = pi342 & w13947;
assign w13996 = w13905 & w13995;
assign w13997 = (pi372 & ~w13995) | (pi372 & w19585) | (~w13995 & w19585);
assign w13998 = pi342 & w13959;
assign w13999 = ~w13953 & ~w13998;
assign w14000 = ~pi352 & w13994;
assign w14001 = w13999 & w19586;
assign w14002 = ~w13992 & w14001;
assign w14003 = ~w13987 & ~w14002;
assign w14004 = ~pi321 & pi342;
assign w14005 = w13905 & w14004;
assign w14006 = pi352 & ~w14005;
assign w14007 = w13947 & w13956;
assign w14008 = ~pi182 & pi321;
assign w14009 = pi342 & w13905;
assign w14010 = w14008 & w14009;
assign w14011 = ~w14007 & ~w14010;
assign w14012 = ~w14010 & w19587;
assign w14013 = ~w14006 & ~w14012;
assign w14014 = pi182 & pi352;
assign w14015 = w13989 & w14014;
assign w14016 = w13912 & w13966;
assign w14017 = ~w14015 & ~w14016;
assign w14018 = ~pi191 & w14017;
assign w14019 = ~w14013 & w14018;
assign w14020 = ~w13964 & w19588;
assign w14021 = ~w14003 & w14019;
assign w14022 = ~w14020 & ~w14021;
assign w14023 = pi182 & ~pi321;
assign w14024 = w14023 & w13905;
assign w14025 = (pi352 & ~w13932) | (pi352 & w19589) | (~w13932 & w19589);
assign w14026 = ~pi321 & w13956;
assign w14027 = pi321 & w13980;
assign w14028 = ~w14026 & ~w14027;
assign w14029 = (w13938 & ~w14028) | (w13938 & w19590) | (~w14028 & w19590);
assign w14030 = pi182 & ~pi352;
assign w14031 = w13980 & w14004;
assign w14032 = w14030 & w14031;
assign w14033 = ~w14025 & ~w14029;
assign w14034 = (pi372 & ~w14033) | (pi372 & w19591) | (~w14033 & w19591);
assign w14035 = pi352 & ~pi372;
assign w14036 = w13980 & w13990;
assign w14037 = ~w14016 & ~w14036;
assign w14038 = w14035 & ~w14037;
assign w14039 = pi182 & w13930;
assign w14040 = ~pi321 & pi352;
assign w14041 = w14039 & w14040;
assign w14042 = ~pi352 & ~pi372;
assign w14043 = w14004 & w14042;
assign w14044 = pi276 & ~pi321;
assign w14045 = w13904 & w14044;
assign w14046 = (w14045 & w14041) | (w14045 & w19592) | (w14041 & w19592);
assign w14047 = w13922 & w14014;
assign w14048 = w13947 & w13966;
assign w14049 = w13922 & w19593;
assign w14050 = ~w14048 & ~w14049;
assign w14051 = ~w14038 & w19594;
assign w14052 = ~w14034 & w14051;
assign w14053 = ~w14022 & w19595;
assign w14054 = (~w13903 & w14022) | (~w13903 & w19596) | (w14022 & w19596);
assign w14055 = pi532 & pi576;
assign w14056 = ~w14053 & ~w14054;
assign w14057 = ~pi532 & w14056;
assign w14058 = ~w14055 & ~w14057;
assign w14059 = ~pi135 & pi138;
assign w14060 = pi135 & ~pi138;
assign w14061 = ~w14059 & ~w14060;
assign w14062 = w13885 & w14061;
assign w14063 = ~w13885 & ~w14061;
assign w14064 = ~w14062 & ~w14063;
assign w14065 = w13867 & ~w14064;
assign w14066 = ~w13867 & w14064;
assign w14067 = pi532 & pi560;
assign w14068 = ~w14065 & ~w14066;
assign w14069 = ~pi532 & w14068;
assign w14070 = ~w14067 & ~w14069;
assign w14071 = pi351 & w13463;
assign w14072 = ~w13476 & ~w13608;
assign w14073 = ~w13552 & ~w14072;
assign w14074 = ~w14073 & w19597;
assign w14075 = pi284 & ~w14074;
assign w14076 = w13464 & w13565;
assign w14077 = ~w13778 & ~w14076;
assign w14078 = ~w13491 & w14077;
assign w14079 = ~pi351 & ~w14078;
assign w14080 = w13510 & w13554;
assign w14081 = ~w13593 & ~w14080;
assign w14082 = ~pi351 & w13478;
assign w14083 = ~pi132 & ~w14081;
assign w14084 = ~w14082 & ~w14083;
assign w14085 = ~w13539 & ~w13554;
assign w14086 = w13596 & ~w14085;
assign w14087 = w13525 & w13850;
assign w14088 = ~pi284 & w13509;
assign w14089 = (~pi193 & ~w14088) | (~pi193 & w19598) | (~w14088 & w19598);
assign w14090 = ~w14086 & w19599;
assign w14091 = ~pi284 & ~w14084;
assign w14092 = w14090 & ~w14091;
assign w14093 = ~w13489 & ~w13516;
assign w14094 = (pi351 & ~w14093) | (pi351 & w19600) | (~w14093 & w19600);
assign w14095 = w13484 & w13565;
assign w14096 = ~w13534 & ~w14095;
assign w14097 = w14096 & w19601;
assign w14098 = w13544 & w13553;
assign w14099 = w14097 & ~w14098;
assign w14100 = ~w13528 & ~w13590;
assign w14101 = pi284 & ~w13556;
assign w14102 = (~pi351 & w13590) | (~pi351 & w19602) | (w13590 & w19602);
assign w14103 = w14101 & ~w14102;
assign w14104 = (~w14103 & ~w14099) | (~w14103 & w19603) | (~w14099 & w19603);
assign w14105 = pi132 & w13560;
assign w14106 = ~w13486 & ~w14105;
assign w14107 = w13464 & w13592;
assign w14108 = pi351 & ~w14107;
assign w14109 = w14106 & w19604;
assign w14110 = (~w13555 & w13529) | (~w13555 & w19605) | (w13529 & w19605);
assign w14111 = (~pi351 & ~w13554) | (~pi351 & w13544) | (~w13554 & w13544);
assign w14112 = ~pi358 & w13466;
assign w14113 = w13484 & w13550;
assign w14114 = w14111 & ~w14112;
assign w14115 = w14114 & w19606;
assign w14116 = ~w14109 & ~w14115;
assign w14117 = w13459 & w19607;
assign w14118 = pi193 & ~w14117;
assign w14119 = ~w14116 & w14118;
assign w14120 = ~w14104 & w14119;
assign w14121 = w14092 & w19608;
assign w14122 = ~w14120 & ~w14121;
assign w14123 = w13477 & w19609;
assign w14124 = w13500 & w13509;
assign w14125 = pi351 & w13466;
assign w14126 = w13509 & w13555;
assign w14127 = w13554 & w14126;
assign w14128 = ~w14125 & ~w14127;
assign w14129 = w13471 & w13544;
assign w14130 = w14128 & ~w14129;
assign w14131 = ~pi358 & w13489;
assign w14132 = (pi284 & ~w13539) | (pi284 & w19610) | (~w13539 & w19610);
assign w14133 = w13464 & w13786;
assign w14134 = ~pi358 & w14133;
assign w14135 = ~w13486 & ~w14134;
assign w14136 = (pi351 & ~w14135) | (pi351 & w19611) | (~w14135 & w19611);
assign w14137 = w13484 & w19528;
assign w14138 = ~w13607 & ~w13796;
assign w14139 = ~w14137 & w14138;
assign w14140 = w13544 & ~w14139;
assign w14141 = w13460 & w19522;
assign w14142 = ~pi284 & ~w14141;
assign w14143 = ~w14140 & w14142;
assign w14144 = ~w14136 & w14143;
assign w14145 = ~w14131 & w14132;
assign w14146 = w14130 & w14145;
assign w14147 = ~w14144 & ~w14146;
assign w14148 = (pi275 & w14124) | (pi275 & w19612) | (w14124 & w19612);
assign w14149 = ~w14147 & ~w14148;
assign w14150 = ~w14122 & w14149;
assign w14151 = ~pi394 & w14150;
assign w14152 = pi394 & ~w14150;
assign w14153 = ~w14151 & ~w14152;
assign w14154 = ~pi160 & pi164;
assign w14155 = pi160 & ~pi164;
assign w14156 = ~w14154 & ~w14155;
assign w14157 = ~pi139 & pi162;
assign w14158 = pi139 & ~pi162;
assign w14159 = ~w14157 & ~w14158;
assign w14160 = w14156 & w14159;
assign w14161 = ~w14156 & ~w14159;
assign w14162 = ~w14160 & ~w14161;
assign w14163 = ~w14153 & ~w14162;
assign w14164 = w14153 & w14162;
assign w14165 = pi532 & pi557;
assign w14166 = ~w14163 & ~w14164;
assign w14167 = ~pi532 & w14166;
assign w14168 = ~w14165 & ~w14167;
assign w14169 = ~pi388 & ~w13624;
assign w14170 = pi388 & w13624;
assign w14171 = ~w14169 & ~w14170;
assign w14172 = w13618 & w19613;
assign w14173 = (pi144 & ~w13618) | (pi144 & w19614) | (~w13618 & w19614);
assign w14174 = ~w14172 & ~w14173;
assign w14175 = ~w14171 & ~w14174;
assign w14176 = w14171 & w14174;
assign w14177 = pi532 & pi594;
assign w14178 = ~w14175 & ~w14176;
assign w14179 = ~pi532 & w14178;
assign w14180 = ~w14177 & ~w14179;
assign w14181 = ~pi141 & ~w13621;
assign w14182 = pi141 & w13621;
assign w14183 = ~w14181 & ~w14182;
assign w14184 = pi532 & ~pi658;
assign w14185 = ~pi532 & ~w14183;
assign w14186 = ~w14184 & ~w14185;
assign w14187 = ~pi142 & pi167;
assign w14188 = pi142 & ~pi167;
assign w14189 = ~w14187 & ~w14188;
assign w14190 = ~pi138 & ~pi185;
assign w14191 = pi147 & ~pi166;
assign w14192 = w14190 & w14191;
assign w14193 = ~pi138 & pi185;
assign w14194 = pi129 & ~pi147;
assign w14195 = w14193 & w14194;
assign w14196 = ~pi147 & pi166;
assign w14197 = pi138 & w14196;
assign w14198 = ~w14192 & ~w14195;
assign w14199 = (~pi207 & ~w14198) | (~pi207 & w19615) | (~w14198 & w19615);
assign w14200 = pi166 & ~pi185;
assign w14201 = w14194 & w14200;
assign w14202 = ~pi129 & pi147;
assign w14203 = ~pi138 & pi166;
assign w14204 = w14202 & w14203;
assign w14205 = ~pi129 & ~pi147;
assign w14206 = pi138 & ~pi166;
assign w14207 = w14205 & w14206;
assign w14208 = pi129 & pi166;
assign w14209 = pi138 & pi185;
assign w14210 = pi138 & pi207;
assign w14211 = ~w14209 & ~w14210;
assign w14212 = w14208 & ~w14211;
assign w14213 = pi129 & pi147;
assign w14214 = ~pi166 & pi185;
assign w14215 = w14213 & w14214;
assign w14216 = pi207 & w14215;
assign w14217 = pi129 & w14191;
assign w14218 = w14190 & w14217;
assign w14219 = ~w14212 & ~w14216;
assign w14220 = ~w14218 & w14219;
assign w14221 = ~w14201 & ~w14204;
assign w14222 = ~w14207 & w14221;
assign w14223 = w14220 & w19616;
assign w14224 = ~pi185 & w14210;
assign w14225 = w14210 & w19617;
assign w14226 = ~pi147 & w14203;
assign w14227 = w14203 & w19618;
assign w14228 = ~w14225 & ~w14227;
assign w14229 = ~pi129 & ~w14228;
assign w14230 = w14190 & w14213;
assign w14231 = pi166 & w14230;
assign w14232 = ~pi138 & pi207;
assign w14233 = ~pi147 & ~pi166;
assign w14234 = ~pi129 & w14233;
assign w14235 = w14232 & w14234;
assign w14236 = ~w14231 & ~w14235;
assign w14237 = ~w14229 & w14236;
assign w14238 = ~pi302 & ~w14237;
assign w14239 = pi185 & w14208;
assign w14240 = ~pi166 & ~pi185;
assign w14241 = ~pi129 & w14240;
assign w14242 = ~w14239 & ~w14241;
assign w14243 = ~pi185 & w14233;
assign w14244 = ~pi166 & w14193;
assign w14245 = w14202 & w14244;
assign w14246 = ~w14243 & ~w14245;
assign w14247 = pi138 & ~w14242;
assign w14248 = w14246 & ~w14247;
assign w14249 = ~pi129 & pi138;
assign w14250 = w14214 & w14249;
assign w14251 = pi147 & ~pi185;
assign w14252 = ~pi129 & pi166;
assign w14253 = w14251 & w14252;
assign w14254 = ~w14250 & ~w14253;
assign w14255 = ~pi207 & ~w14254;
assign w14256 = pi129 & w14196;
assign w14257 = w14196 & w19619;
assign w14258 = ~pi207 & w14257;
assign w14259 = w14233 & w19620;
assign w14260 = ~w14255 & w19621;
assign w14261 = pi207 & ~w14248;
assign w14262 = w14260 & ~w14261;
assign w14263 = ~w14238 & w14262;
assign w14264 = w14209 & w14233;
assign w14265 = ~pi129 & w14251;
assign w14266 = ~w14264 & ~w14265;
assign w14267 = pi207 & ~w14266;
assign w14268 = pi147 & w14208;
assign w14269 = w14193 & w14268;
assign w14270 = pi138 & pi166;
assign w14271 = w14205 & w14270;
assign w14272 = w14217 & ~w14232;
assign w14273 = ~pi207 & w14271;
assign w14274 = ~w14272 & ~w14273;
assign w14275 = (~pi302 & ~w14268) | (~pi302 & w19623) | (~w14268 & w19623);
assign w14276 = ~w14267 & w14274;
assign w14277 = w14275 & w14276;
assign w14278 = w14205 & w14214;
assign w14279 = ~pi138 & w14278;
assign w14280 = (pi302 & ~w14278) | (pi302 & w19624) | (~w14278 & w19624);
assign w14281 = w14196 & w14306;
assign w14282 = pi166 & w14195;
assign w14283 = ~pi147 & w14209;
assign w14284 = pi129 & ~pi166;
assign w14285 = w14283 & w14284;
assign w14286 = ~w14281 & ~w14282;
assign w14287 = w14286 & w19625;
assign w14288 = ~w14277 & ~w14287;
assign w14289 = w14206 & w14213;
assign w14290 = w14206 & w14251;
assign w14291 = ~w14289 & ~w14290;
assign w14292 = pi147 & pi166;
assign w14293 = pi185 & w14292;
assign w14294 = w14292 & w19626;
assign w14295 = ~pi185 & w14284;
assign w14296 = (~pi207 & ~w14284) | (~pi207 & w19627) | (~w14284 & w19627);
assign w14297 = w14291 & w19628;
assign w14298 = ~pi166 & w14202;
assign w14299 = w14190 & w14298;
assign w14300 = ~w14269 & ~w14299;
assign w14301 = pi207 & w14300;
assign w14302 = ~w14297 & ~w14301;
assign w14303 = ~pi129 & ~w14251;
assign w14304 = ~pi207 & pi302;
assign w14305 = pi185 & w14252;
assign w14306 = pi138 & ~pi185;
assign w14307 = pi129 & w14306;
assign w14308 = ~w14191 & ~w14304;
assign w14309 = w14307 & ~w14308;
assign w14310 = w14303 & ~w14305;
assign w14311 = w14304 & w14310;
assign w14312 = ~w14309 & ~w14311;
assign w14313 = ~w14302 & w14312;
assign w14314 = ~w14288 & w14313;
assign w14315 = pi139 & ~w14314;
assign w14316 = w14202 & w14214;
assign w14317 = ~pi129 & w14196;
assign w14318 = w14196 & w19626;
assign w14319 = ~w14316 & ~w14318;
assign w14320 = w14209 & w14194;
assign w14321 = ~w14269 & ~w14320;
assign w14322 = w14193 & ~w14319;
assign w14323 = w14321 & ~w14322;
assign w14324 = pi166 & w14190;
assign w14325 = ~pi207 & w14200;
assign w14326 = w14200 & w19629;
assign w14327 = ~pi207 & w14294;
assign w14328 = w14190 & w14233;
assign w14329 = pi138 & ~pi207;
assign w14330 = w14215 & w14329;
assign w14331 = ~w14328 & ~w14330;
assign w14332 = w14324 & w14326;
assign w14333 = w14331 & w19630;
assign w14334 = pi207 & ~w14323;
assign w14335 = (~pi302 & w14334) | (~pi302 & w19631) | (w14334 & w19631);
assign w14336 = pi207 & ~w14285;
assign w14337 = w14194 & w14240;
assign w14338 = pi138 & w14337;
assign w14339 = (~pi207 & ~w14337) | (~pi207 & w14436) | (~w14337 & w14436);
assign w14340 = ~w14204 & w14339;
assign w14341 = ~w14336 & ~w14340;
assign w14342 = w14233 & w14306;
assign w14343 = ~pi129 & w14342;
assign w14344 = w14215 & w14232;
assign w14345 = ~w14258 & ~w14343;
assign w14346 = (pi302 & ~w14345) | (pi302 & w19632) | (~w14345 & w19632);
assign w14347 = ~w14341 & ~w14346;
assign w14348 = ~w14315 & w19633;
assign w14349 = w14348 & w19634;
assign w14350 = (pi178 & ~w14348) | (pi178 & w19635) | (~w14348 & w19635);
assign w14351 = ~w14349 & ~w14350;
assign w14352 = ~w14189 & ~w14351;
assign w14353 = w14189 & w14351;
assign w14354 = pi532 & pi570;
assign w14355 = ~w14352 & ~w14353;
assign w14356 = ~pi532 & w14355;
assign w14357 = ~w14354 & ~w14356;
assign w14358 = ~pi143 & pi181;
assign w14359 = pi143 & ~pi181;
assign w14360 = ~w14358 & ~w14359;
assign w14361 = ~pi180 & ~w14360;
assign w14362 = pi180 & w14360;
assign w14363 = ~w14361 & ~w14362;
assign w14364 = w14202 & w14206;
assign w14365 = pi207 & ~w14271;
assign w14366 = ~w14217 & ~w14295;
assign w14367 = w14365 & w14366;
assign w14368 = ~w14204 & ~w14364;
assign w14369 = ~pi207 & w14368;
assign w14370 = ~w14367 & ~w14369;
assign w14371 = pi166 & w14209;
assign w14372 = w14205 & w14371;
assign w14373 = (~pi302 & ~w14371) | (~pi302 & w19636) | (~w14371 & w19636);
assign w14374 = ~w14230 & ~w14328;
assign w14375 = w14373 & w14374;
assign w14376 = ~w14370 & w14375;
assign w14377 = ~pi138 & w14191;
assign w14378 = (pi207 & ~w14252) | (pi207 & w16325) | (~w14252 & w16325);
assign w14379 = w14194 & ~w14206;
assign w14380 = w14378 & ~w14379;
assign w14381 = ~w14234 & ~w14377;
assign w14382 = ~pi207 & w14381;
assign w14383 = ~w14380 & ~w14382;
assign w14384 = w14202 & w14270;
assign w14385 = ~w14257 & ~w14384;
assign w14386 = w14193 & w14208;
assign w14387 = pi302 & ~w14386;
assign w14388 = w14385 & w14387;
assign w14389 = ~w14383 & w14388;
assign w14390 = w14190 & w14252;
assign w14391 = w14213 & w14270;
assign w14392 = w14209 & w14196;
assign w14393 = pi207 & ~w14392;
assign w14394 = w14319 & w14393;
assign w14395 = ~w14390 & ~w14391;
assign w14396 = ~pi207 & w14395;
assign w14397 = ~w14394 & ~w14396;
assign w14398 = w14195 & w19637;
assign w14399 = (pi139 & ~w14290) | (pi139 & w19638) | (~w14290 & w19638);
assign w14400 = ~w14398 & w14399;
assign w14401 = ~w14397 & w14400;
assign w14402 = ~w14376 & ~w14389;
assign w14403 = w14401 & ~w14402;
assign w14404 = w14257 & w14329;
assign w14405 = w14194 & w14214;
assign w14406 = w14203 & ~w14205;
assign w14407 = ~w14405 & ~w14406;
assign w14408 = ~w14278 & ~w14390;
assign w14409 = ~pi302 & w14408;
assign w14410 = pi207 & ~w14407;
assign w14411 = w14409 & ~w14410;
assign w14412 = pi185 & w14213;
assign w14413 = w14270 & w14412;
assign w14414 = ~pi207 & w14201;
assign w14415 = ~w14413 & ~w14414;
assign w14416 = w14240 & w19639;
assign w14417 = w14415 & ~w14416;
assign w14418 = pi302 & ~w14271;
assign w14419 = ~w14231 & w14418;
assign w14420 = ~w14344 & w14419;
assign w14421 = ~w14404 & w14411;
assign w14422 = w14417 & w14420;
assign w14423 = ~w14421 & ~w14422;
assign w14424 = pi138 & w14191;
assign w14425 = w14191 & w14209;
assign w14426 = ~w14269 & ~w14425;
assign w14427 = w14208 & w14251;
assign w14428 = pi207 & ~w14427;
assign w14429 = w14240 & w14249;
assign w14430 = w14428 & ~w14429;
assign w14431 = ~w14269 & w19640;
assign w14432 = ~w14430 & ~w14431;
assign w14433 = (~pi139 & ~w14298) | (~pi139 & w19641) | (~w14298 & w19641);
assign w14434 = ~w14432 & w14433;
assign w14435 = ~w14423 & w14434;
assign w14436 = ~pi138 & ~pi207;
assign w14437 = ~pi185 & w14191;
assign w14438 = pi185 & w14205;
assign w14439 = ~w14201 & ~w14437;
assign w14440 = (w14436 & ~w14439) | (w14436 & w19642) | (~w14439 & w19642);
assign w14441 = w14200 & w14205;
assign w14442 = w14329 & w14441;
assign w14443 = w14213 & w14224;
assign w14444 = ~w14442 & ~w14443;
assign w14445 = pi207 & ~w14385;
assign w14446 = w14444 & ~w14445;
assign w14447 = (pi302 & ~w14446) | (pi302 & w19643) | (~w14446 & w19643);
assign w14448 = pi207 & ~pi302;
assign w14449 = ~w14279 & ~w14299;
assign w14450 = w14448 & ~w14449;
assign w14451 = w14210 & w14265;
assign w14452 = w14200 & w19644;
assign w14453 = w14251 & w14270;
assign w14454 = (w14453 & w14451) | (w14453 & w19645) | (w14451 & w19645);
assign w14455 = w14371 & w20902;
assign w14456 = pi147 & w14250;
assign w14457 = ~w14450 & ~w14454;
assign w14458 = ~w14455 & ~w14456;
assign w14459 = w14457 & w14458;
assign w14460 = ~w14403 & ~w14435;
assign w14461 = ~w14460 & w19646;
assign w14462 = (~w14363 & w14460) | (~w14363 & w19647) | (w14460 & w19647);
assign w14463 = pi532 & pi568;
assign w14464 = ~w14461 & ~w14462;
assign w14465 = ~pi532 & w14464;
assign w14466 = ~w14463 & ~w14465;
assign w14467 = ~pi144 & ~w14183;
assign w14468 = pi144 & w14183;
assign w14469 = ~w14467 & ~w14468;
assign w14470 = w13476 & w19607;
assign w14471 = ~pi351 & w14470;
assign w14472 = ~w13526 & ~w14471;
assign w14473 = pi351 & ~w13609;
assign w14474 = w14472 & ~w14473;
assign w14475 = (~pi284 & ~w14474) | (~pi284 & w19648) | (~w14474 & w19648);
assign w14476 = w13475 & w13786;
assign w14477 = ~w14476 & w19649;
assign w14478 = pi351 & ~w14477;
assign w14479 = w13505 & w13544;
assign w14480 = w14106 & ~w14479;
assign w14481 = ~w14478 & w14480;
assign w14482 = pi284 & ~w14481;
assign w14483 = w13510 & w13528;
assign w14484 = ~w13466 & ~w13602;
assign w14485 = pi351 & w14484;
assign w14486 = w13798 & w14485;
assign w14487 = w13573 & ~w14483;
assign w14488 = ~w14486 & ~w14487;
assign w14489 = ~w14482 & w19650;
assign w14490 = pi193 & ~w14489;
assign w14491 = w13515 & w13550;
assign w14492 = ~w14123 & ~w14491;
assign w14493 = w13514 & w13534;
assign w14494 = w14492 & ~w14493;
assign w14495 = ~w13542 & ~w14112;
assign w14496 = w13481 & w13565;
assign w14497 = ~w14483 & ~w14496;
assign w14498 = ~pi284 & w14497;
assign w14499 = w14495 & w14498;
assign w14500 = ~pi351 & w13602;
assign w14501 = w13477 & w13528;
assign w14502 = ~pi354 & w14501;
assign w14503 = ~w14500 & ~w14502;
assign w14504 = ~w13513 & w14503;
assign w14505 = pi284 & w14504;
assign w14506 = w14494 & w14499;
assign w14507 = ~w14505 & ~w14506;
assign w14508 = ~w13476 & w13534;
assign w14509 = w13464 & w13550;
assign w14510 = ~w14508 & ~w14509;
assign w14511 = ~w13776 & ~w13813;
assign w14512 = w14510 & w14511;
assign w14513 = pi351 & ~w14076;
assign w14514 = ~w14491 & w14513;
assign w14515 = (~w14514 & ~w14512) | (~w14514 & w19651) | (~w14512 & w19651);
assign w14516 = (~pi193 & w14507) | (~pi193 & w19652) | (w14507 & w19652);
assign w14517 = w13465 & w13571;
assign w14518 = pi351 & ~w13593;
assign w14519 = ~w13531 & w14518;
assign w14520 = ~w13556 & ~w14517;
assign w14521 = w13603 & w14520;
assign w14522 = ~w14519 & ~w14521;
assign w14523 = ~w13579 & ~w13831;
assign w14524 = (~pi284 & w14522) | (~pi284 & w19653) | (w14522 & w19653);
assign w14525 = ~pi351 & ~w13566;
assign w14526 = ~w13489 & ~w13859;
assign w14527 = ~w14525 & ~w14526;
assign w14528 = pi284 & pi351;
assign w14529 = ~w13488 & ~w14517;
assign w14530 = (~w13792 & w14529) | (~w13792 & w19654) | (w14529 & w19654);
assign w14531 = w14528 & ~w14530;
assign w14532 = w13539 & w19655;
assign w14533 = ~w13785 & ~w14532;
assign w14534 = ~w14527 & ~w14531;
assign w14535 = w14533 & w14534;
assign w14536 = ~w14524 & w14535;
assign w14537 = ~w14516 & w14536;
assign w14538 = ~w14490 & w14537;
assign w14539 = ~pi391 & w14538;
assign w14540 = pi391 & ~w14538;
assign w14541 = ~w14539 & ~w14540;
assign w14542 = ~pi145 & ~w14541;
assign w14543 = pi145 & w14541;
assign w14544 = pi532 & pi659;
assign w14545 = ~w14542 & ~w14543;
assign w14546 = ~pi532 & w14545;
assign w14547 = ~w14544 & ~w14546;
assign w14548 = ~pi145 & pi146;
assign w14549 = pi145 & ~pi146;
assign w14550 = ~w14548 & ~w14549;
assign w14551 = ~w14541 & ~w14550;
assign w14552 = w14541 & w14550;
assign w14553 = pi532 & pi627;
assign w14554 = ~w14551 & ~w14552;
assign w14555 = ~pi532 & w14554;
assign w14556 = ~w14553 & ~w14555;
assign w14557 = ~pi145 & pi153;
assign w14558 = pi145 & ~pi153;
assign w14559 = ~w14557 & ~w14558;
assign w14560 = ~pi146 & pi147;
assign w14561 = pi146 & ~pi147;
assign w14562 = ~w14560 & ~w14561;
assign w14563 = w14559 & w14562;
assign w14564 = ~w14559 & ~w14562;
assign w14565 = ~w14563 & ~w14564;
assign w14566 = w14541 & ~w14565;
assign w14567 = ~w14541 & w14565;
assign w14568 = pi532 & pi563;
assign w14569 = ~w14566 & ~w14567;
assign w14570 = ~pi532 & w14569;
assign w14571 = ~w14568 & ~w14570;
assign w14572 = w13764 & w19656;
assign w14573 = (pi148 & ~w13764) | (pi148 & w19657) | (~w13764 & w19657);
assign w14574 = ~w14572 & ~w14573;
assign w14575 = pi532 & ~pi650;
assign w14576 = ~pi532 & ~w14574;
assign w14577 = ~w14575 & ~w14576;
assign w14578 = pi149 & ~w14574;
assign w14579 = ~pi149 & w14574;
assign w14580 = pi532 & pi618;
assign w14581 = ~w14578 & ~w14579;
assign w14582 = ~pi532 & w14581;
assign w14583 = ~w14580 & ~w14582;
assign w14584 = ~pi150 & pi187;
assign w14585 = pi150 & ~pi187;
assign w14586 = ~w14584 & ~w14585;
assign w14587 = w14233 & w19658;
assign w14588 = ~w14294 & ~w14587;
assign w14589 = (pi207 & ~w14588) | (pi207 & w14216) | (~w14588 & w14216);
assign w14590 = w14252 & w14436;
assign w14591 = ~pi147 & w14590;
assign w14592 = pi129 & ~w14196;
assign w14593 = w14284 & w14190;
assign w14594 = ~pi302 & ~w14593;
assign w14595 = w14306 & ~w14592;
assign w14596 = w14594 & ~w14595;
assign w14597 = w14590 & w19618;
assign w14598 = w14596 & ~w14597;
assign w14599 = ~pi129 & ~w14233;
assign w14600 = ~pi207 & ~w14194;
assign w14601 = ~w14599 & w14600;
assign w14602 = pi302 & ~w14316;
assign w14603 = ~w14601 & w14602;
assign w14604 = (~w14603 & ~w14598) | (~w14603 & w19659) | (~w14598 & w19659);
assign w14605 = pi129 & ~pi185;
assign w14606 = w14270 & w14605;
assign w14607 = ~w14285 & ~w14606;
assign w14608 = pi207 & ~w14441;
assign w14609 = ~w14282 & w14608;
assign w14610 = w14607 & w14609;
assign w14611 = w14208 & w19660;
assign w14612 = w14193 & w14284;
assign w14613 = ~pi166 & w14306;
assign w14614 = ~w14612 & ~w14613;
assign w14615 = (~pi207 & ~w14202) | (~pi207 & w14436) | (~w14202 & w14436);
assign w14616 = w14306 & w14317;
assign w14617 = ~w14611 & w14614;
assign w14618 = w14615 & ~w14616;
assign w14619 = w14617 & w14618;
assign w14620 = w14191 & w19661;
assign w14621 = ~w14610 & ~w14619;
assign w14622 = ~w14620 & ~w14621;
assign w14623 = (pi139 & ~w14622) | (pi139 & w19662) | (~w14622 & w19662);
assign w14624 = w14191 & w20531;
assign w14625 = ~w14293 & ~w14624;
assign w14626 = ~w14209 & w14233;
assign w14627 = ~w14590 & ~w14626;
assign w14628 = (pi138 & w14624) | (pi138 & w19663) | (w14624 & w19663);
assign w14629 = ~pi207 & w14264;
assign w14630 = w14202 & w14240;
assign w14631 = ~w14427 & ~w14630;
assign w14632 = ~pi138 & ~w14631;
assign w14633 = w14190 & w14205;
assign w14634 = ~w14391 & ~w14633;
assign w14635 = ~w14282 & w14634;
assign w14636 = ~pi207 & ~w14635;
assign w14637 = ~pi166 & w14194;
assign w14638 = ~w14202 & ~w14637;
assign w14639 = w14224 & ~w14638;
assign w14640 = ~w14196 & ~w14203;
assign w14641 = pi129 & w14448;
assign w14642 = ~w14640 & w14641;
assign w14643 = ~w14639 & ~w14642;
assign w14644 = ~w14636 & w14643;
assign w14645 = (~pi302 & w14632) | (~pi302 & w19664) | (w14632 & w19664);
assign w14646 = w14644 & ~w14645;
assign w14647 = (pi302 & w14628) | (pi302 & w19665) | (w14628 & w19665);
assign w14648 = w14205 & w14324;
assign w14649 = ~w14285 & ~w14648;
assign w14650 = (pi207 & ~w14649) | (pi207 & w19666) | (~w14649 & w19666);
assign w14651 = w14191 & ~w14605;
assign w14652 = ~w14337 & ~w14651;
assign w14653 = w14290 & w19629;
assign w14654 = w14436 & ~w14652;
assign w14655 = ~w14653 & ~w14654;
assign w14656 = ~w14650 & w14655;
assign w14657 = ~pi302 & ~w14656;
assign w14658 = w14209 & w19637;
assign w14659 = ~w14192 & ~w14658;
assign w14660 = ~w14625 & ~w14659;
assign w14661 = w14232 & w14316;
assign w14662 = pi207 & w14271;
assign w14663 = ~pi166 & w14633;
assign w14664 = ~w14662 & ~w14663;
assign w14665 = w14239 & w14436;
assign w14666 = w14664 & ~w14665;
assign w14667 = ~w14338 & ~w14661;
assign w14668 = (pi302 & ~w14666) | (pi302 & w19667) | (~w14666 & w19667);
assign w14669 = ~w14660 & ~w14668;
assign w14670 = ~w14657 & w14669;
assign w14671 = (~pi139 & ~w14646) | (~pi139 & w19668) | (~w14646 & w19668);
assign w14672 = w14670 & ~w14671;
assign w14673 = w14672 & w19669;
assign w14674 = (pi190 & ~w14672) | (pi190 & w19670) | (~w14672 & w19670);
assign w14675 = ~w14673 & ~w14674;
assign w14676 = ~w14586 & ~w14675;
assign w14677 = w14586 & w14675;
assign w14678 = pi532 & pi565;
assign w14679 = ~w14676 & ~w14677;
assign w14680 = ~pi532 & w14679;
assign w14681 = ~w14678 & ~w14680;
assign w14682 = ~pi151 & pi222;
assign w14683 = pi151 & ~pi222;
assign w14684 = ~w14682 & ~w14683;
assign w14685 = ~pi229 & ~w14684;
assign w14686 = pi229 & w14684;
assign w14687 = ~w14685 & ~w14686;
assign w14688 = w13911 & w14044;
assign w14689 = w13946 & w14008;
assign w14690 = ~w14688 & ~w14689;
assign w14691 = ~w13996 & w14690;
assign w14692 = ~pi352 & ~w14691;
assign w14693 = w13989 & w19671;
assign w14694 = pi276 & pi342;
assign w14695 = ~pi170 & w14694;
assign w14696 = w14694 & w19672;
assign w14697 = pi372 & ~w14696;
assign w14698 = ~w14693 & w14697;
assign w14699 = ~w14692 & w14698;
assign w14700 = ~w14005 & w19673;
assign w14701 = ~pi182 & w13906;
assign w14702 = w13906 & w13918;
assign w14703 = w13950 & w19584;
assign w14704 = w13947 & w13950;
assign w14705 = pi276 & w14704;
assign w14706 = w13949 & ~w14702;
assign w14707 = ~w14703 & ~w14705;
assign w14708 = w14706 & w14707;
assign w14709 = (~w13935 & w14700) | (~w13935 & w19674) | (w14700 & w19674);
assign w14710 = ~w14708 & ~w14709;
assign w14711 = ~w13947 & ~w14004;
assign w14712 = (~pi372 & w14711) | (~pi372 & w19675) | (w14711 & w19675);
assign w14713 = ~w14710 & w14712;
assign w14714 = w13950 & w14044;
assign w14715 = w14030 & w14714;
assign w14716 = ~pi321 & w13916;
assign w14717 = w13916 & w14040;
assign w14718 = pi372 & ~w14717;
assign w14719 = (pi352 & ~w13946) | (pi352 & w13965) | (~w13946 & w13965);
assign w14720 = w13928 & w13930;
assign w14721 = ~w13942 & ~w14720;
assign w14722 = ~pi352 & w14721;
assign w14723 = ~w13919 & ~w13957;
assign w14724 = w14719 & w14723;
assign w14725 = ~w14722 & ~w14724;
assign w14726 = w13950 & w13912;
assign w14727 = ~pi372 & ~w14045;
assign w14728 = ~w14702 & ~w14726;
assign w14729 = w14727 & w14728;
assign w14730 = ~w14715 & w14718;
assign w14731 = (~w14730 & w14725) | (~w14730 & w19676) | (w14725 & w19676);
assign w14732 = pi170 & w13916;
assign w14733 = w13916 & w19677;
assign w14734 = w13930 & w19678;
assign w14735 = ~w14733 & ~w14734;
assign w14736 = (w14014 & ~w14735) | (w14014 & w19679) | (~w14735 & w19679);
assign w14737 = w13905 & w13918;
assign w14738 = pi352 & w14737;
assign w14739 = ~pi182 & w14004;
assign w14740 = w13980 & w14739;
assign w14741 = pi276 & w14008;
assign w14742 = ~w14027 & ~w14741;
assign w14743 = ~pi352 & pi372;
assign w14744 = ~pi276 & w14726;
assign w14745 = ~w14742 & w14743;
assign w14746 = ~w14744 & ~w14745;
assign w14747 = ~w14738 & ~w14740;
assign w14748 = pi191 & w14747;
assign w14749 = w14746 & w14748;
assign w14750 = ~w14736 & w14749;
assign w14751 = ~w14731 & w14750;
assign w14752 = (~pi352 & ~w13930) | (~pi352 & w13938) | (~w13930 & w13938);
assign w14753 = pi182 & w14694;
assign w14754 = w13956 & w14023;
assign w14755 = ~pi182 & w13916;
assign w14756 = ~w14754 & ~w14755;
assign w14757 = pi352 & w14756;
assign w14758 = ~w13989 & ~w14753;
assign w14759 = w14752 & w14758;
assign w14760 = ~w14757 & ~w14759;
assign w14761 = (pi372 & w14760) | (pi372 & w19680) | (w14760 & w19680);
assign w14762 = w13950 & w14030;
assign w14763 = ~w13935 & ~w14762;
assign w14764 = w14030 & w14703;
assign w14765 = w13931 & w13965;
assign w14766 = ~pi191 & ~w13929;
assign w14767 = ~w14765 & w14766;
assign w14768 = ~w14764 & w14767;
assign w14769 = ~pi372 & ~w14763;
assign w14770 = w14768 & ~w14769;
assign w14771 = ~w14761 & w14770;
assign w14772 = ~w13913 & ~w14702;
assign w14773 = w14040 & ~w14772;
assign w14774 = pi352 & pi372;
assign w14775 = ~w14720 & ~w14739;
assign w14776 = w14774 & ~w14775;
assign w14777 = ~w14032 & ~w14776;
assign w14778 = ~w14773 & w14777;
assign w14779 = (w14778 & w14751) | (w14778 & w19681) | (w14751 & w19681);
assign w14780 = w14779 & w19682;
assign w14781 = (~w14687 & ~w14779) | (~w14687 & w19683) | (~w14779 & w19683);
assign w14782 = pi532 & pi575;
assign w14783 = ~w14780 & ~w14781;
assign w14784 = ~pi532 & w14783;
assign w14785 = ~w14782 & ~w14784;
assign w14786 = ~pi170 & w14023;
assign w14787 = ~pi182 & w13946;
assign w14788 = ~w14786 & ~w14787;
assign w14789 = w14004 & ~w14788;
assign w14790 = w13904 & w13976;
assign w14791 = ~w14714 & ~w14790;
assign w14792 = ~pi372 & w14791;
assign w14793 = w14008 & w14695;
assign w14794 = w14014 & w14732;
assign w14795 = ~w14789 & w14792;
assign w14796 = ~w14793 & ~w14794;
assign w14797 = w14795 & w14796;
assign w14798 = ~w13934 & ~w13989;
assign w14799 = w13979 & ~w14798;
assign w14800 = w13988 & w19584;
assign w14801 = ~pi352 & w14800;
assign w14802 = (pi372 & ~w14704) | (pi372 & w19684) | (~w14704 & w19684);
assign w14803 = ~w14799 & w19685;
assign w14804 = ~w13916 & w14786;
assign w14805 = w13980 & w14008;
assign w14806 = ~w13931 & ~w14805;
assign w14807 = ~w13991 & ~w14804;
assign w14808 = (~pi352 & ~w14807) | (~pi352 & w19686) | (~w14807 & w19686);
assign w14809 = w13912 & w13980;
assign w14810 = (pi352 & w14793) | (pi352 & w19687) | (w14793 & w19687);
assign w14811 = ~pi191 & ~w14810;
assign w14812 = ~w14808 & w14811;
assign w14813 = ~w14797 & ~w14803;
assign w14814 = w14812 & ~w14813;
assign w14815 = w13930 & w14739;
assign w14816 = pi321 & w13956;
assign w14817 = ~w14815 & w19688;
assign w14818 = pi352 & ~w14817;
assign w14819 = pi321 & w13952;
assign w14820 = w13950 & w14819;
assign w14821 = w13933 & w14023;
assign w14822 = ~pi170 & ~w14044;
assign w14823 = w13938 & w14822;
assign w14824 = ~w14821 & ~w14823;
assign w14825 = ~w14820 & w14824;
assign w14826 = ~w14818 & w14825;
assign w14827 = pi372 & ~w14826;
assign w14828 = w13947 & w13988;
assign w14829 = ~w14688 & ~w14828;
assign w14830 = (~pi352 & ~w14829) | (~pi352 & w19689) | (~w14829 & w19689);
assign w14831 = ~w13966 & ~w13995;
assign w14832 = (~w13929 & w14831) | (~w13929 & w14844) | (w14831 & w14844);
assign w14833 = ~w14830 & w14832;
assign w14834 = ~pi372 & ~w14833;
assign w14835 = pi352 & ~w13953;
assign w14836 = ~pi352 & ~w14714;
assign w14837 = ~w14800 & w14835;
assign w14838 = w14011 & w14837;
assign w14839 = (pi191 & w14838) | (pi191 & w19690) | (w14838 & w19690);
assign w14840 = ~w14834 & w14839;
assign w14841 = ~w14827 & w14840;
assign w14842 = ~pi321 & w13923;
assign w14843 = w13923 & w19584;
assign w14844 = ~pi352 & ~w13929;
assign w14845 = w14844 & w19691;
assign w14846 = w14006 & ~w14843;
assign w14847 = ~w14845 & ~w14846;
assign w14848 = ~w13948 & ~w13959;
assign w14849 = ~pi372 & w14848;
assign w14850 = ~w14847 & w14849;
assign w14851 = pi170 & w13946;
assign w14852 = w14023 & w14851;
assign w14853 = ~w14852 & w19692;
assign w14854 = (pi372 & ~w14703) | (pi372 & w19693) | (~w14703 & w19693);
assign w14855 = (w14854 & w14853) | (w14854 & w19694) | (w14853 & w19694);
assign w14856 = w13918 & w13980;
assign w14857 = (~w13976 & w14048) | (~w13976 & w19695) | (w14048 & w19695);
assign w14858 = ~w13978 & ~w14857;
assign w14859 = (w14858 & w14850) | (w14858 & w19696) | (w14850 & w19696);
assign w14860 = ~w14814 & ~w14841;
assign w14861 = ~w14860 & w19697;
assign w14862 = (pi256 & w14860) | (pi256 & w19698) | (w14860 & w19698);
assign w14863 = ~w14861 & ~w14862;
assign w14864 = ~pi152 & pi227;
assign w14865 = pi152 & ~pi227;
assign w14866 = ~w14864 & ~w14865;
assign w14867 = ~w14863 & w14866;
assign w14868 = w14863 & ~w14866;
assign w14869 = ~w14867 & ~w14868;
assign w14870 = pi532 & ~pi579;
assign w14871 = ~pi532 & ~w14869;
assign w14872 = ~w14870 & ~w14871;
assign w14873 = ~pi391 & ~w14559;
assign w14874 = pi391 & w14559;
assign w14875 = ~w14873 & ~w14874;
assign w14876 = ~pi146 & w14538;
assign w14877 = pi146 & ~w14538;
assign w14878 = ~w14876 & ~w14877;
assign w14879 = ~w14875 & ~w14878;
assign w14880 = w14875 & w14878;
assign w14881 = pi532 & pi595;
assign w14882 = ~w14879 & ~w14880;
assign w14883 = ~pi532 & w14882;
assign w14884 = ~w14881 & ~w14883;
assign w14885 = ~pi154 & pi189;
assign w14886 = pi154 & ~pi189;
assign w14887 = ~w14885 & ~w14886;
assign w14888 = ~w13186 & ~w13679;
assign w14889 = ~pi175 & w13203;
assign w14890 = w13203 & w19547;
assign w14891 = (~w14890 & w14888) | (~w14890 & w19699) | (w14888 & w19699);
assign w14892 = pi231 & ~w14891;
assign w14893 = ~pi215 & w13191;
assign w14894 = pi232 & ~w13237;
assign w14895 = w13180 & w13200;
assign w14896 = w13745 & ~w14894;
assign w14897 = ~w14895 & ~w14896;
assign w14898 = w13191 & w19543;
assign w14899 = w14897 & ~w14898;
assign w14900 = ~w14892 & w14899;
assign w14901 = ~pi285 & ~w14900;
assign w14902 = ~pi270 & w13224;
assign w14903 = w13224 & w13745;
assign w14904 = ~w13297 & ~w14903;
assign w14905 = pi231 & w14904;
assign w14906 = w13726 & w14905;
assign w14907 = ~pi233 & w13249;
assign w14908 = w13249 & w13180;
assign w14909 = ~w13197 & ~w13248;
assign w14910 = ~w13737 & ~w14908;
assign w14911 = (~pi231 & w14909) | (~pi231 & w13190) | (w14909 & w13190);
assign w14912 = w14910 & w14911;
assign w14913 = ~pi232 & ~w13203;
assign w14914 = ~pi231 & ~w13213;
assign w14915 = ~w14913 & w14914;
assign w14916 = pi175 & w13297;
assign w14917 = pi234 & ~w13677;
assign w14918 = ~w14916 & w14917;
assign w14919 = (pi285 & w14915) | (pi285 & w19700) | (w14915 & w19700);
assign w14920 = w14918 & ~w14919;
assign w14921 = ~w14906 & ~w14912;
assign w14922 = w14920 & ~w14921;
assign w14923 = ~pi270 & w13310;
assign w14924 = (pi175 & ~w13310) | (pi175 & w13194) | (~w13310 & w13194);
assign w14925 = w13185 & w19701;
assign w14926 = ~w13310 & ~w14925;
assign w14927 = w14924 & ~w14926;
assign w14928 = ~w13194 & w13203;
assign w14929 = ~w13191 & ~w14928;
assign w14930 = pi285 & w14929;
assign w14931 = ~w14927 & w14930;
assign w14932 = ~w13277 & ~w13736;
assign w14933 = w13224 & ~w13243;
assign w14934 = (~pi285 & ~w14933) | (~pi285 & w19702) | (~w14933 & w19702);
assign w14935 = ~pi175 & ~w14932;
assign w14936 = w14934 & ~w14935;
assign w14937 = ~pi285 & w13716;
assign w14938 = w13182 & w13200;
assign w14939 = ~w13231 & ~w14938;
assign w14940 = ~w14937 & w14939;
assign w14941 = ~w13233 & w14940;
assign w14942 = pi232 & w13203;
assign w14943 = ~w13197 & ~w14942;
assign w14944 = (~pi234 & w14943) | (~pi234 & w19703) | (w14943 & w19703);
assign w14945 = (w14944 & w14941) | (w14944 & w19704) | (w14941 & w19704);
assign w14946 = ~w14931 & ~w14936;
assign w14947 = w14945 & ~w14946;
assign w14948 = ~w14901 & w14922;
assign w14949 = ~w14947 & ~w14948;
assign w14950 = w13201 & w13248;
assign w14951 = w13194 & w19705;
assign w14952 = ~w14950 & ~w14951;
assign w14953 = ~w13265 & ~w13310;
assign w14954 = ~w14952 & ~w14953;
assign w14955 = (~pi231 & ~w13181) | (~pi231 & w19706) | (~w13181 & w19706);
assign w14956 = ~pi175 & w13237;
assign w14957 = w13237 & w19547;
assign w14958 = ~pi270 & w14957;
assign w14959 = pi231 & ~w13202;
assign w14960 = ~w13725 & w14959;
assign w14961 = w13213 & w13248;
assign w14962 = pi270 & w13185;
assign w14963 = ~w13279 & ~w14961;
assign w14964 = (w13190 & ~w14963) | (w13190 & w16424) | (~w14963 & w16424);
assign w14965 = ~pi285 & ~w14964;
assign w14966 = (~w14955 & ~w14960) | (~w14955 & w19707) | (~w14960 & w19707);
assign w14967 = w14965 & ~w14966;
assign w14968 = pi231 & ~w13184;
assign w14969 = ~pi231 & ~w13226;
assign w14970 = ~w14968 & ~w14969;
assign w14971 = w13210 & w13236;
assign w14972 = w13210 & w19708;
assign w14973 = ~pi233 & w14938;
assign w14974 = ~w13756 & ~w14973;
assign w14975 = w14974 & w19709;
assign w14976 = ~w14970 & w14975;
assign w14977 = ~w14967 & ~w14976;
assign w14978 = ~w14949 & w19710;
assign w14979 = (pi192 & w14949) | (pi192 & w19711) | (w14949 & w19711);
assign w14980 = ~w14978 & ~w14979;
assign w14981 = ~w14887 & ~w14980;
assign w14982 = w14887 & w14980;
assign w14983 = pi532 & pi581;
assign w14984 = ~w14981 & ~w14982;
assign w14985 = ~pi532 & w14984;
assign w14986 = ~w14983 & ~w14985;
assign w14987 = ~pi155 & pi225;
assign w14988 = pi155 & ~pi225;
assign w14989 = ~w14987 & ~w14988;
assign w14990 = ~pi230 & ~w14989;
assign w14991 = pi230 & w14989;
assign w14992 = ~w14990 & ~w14991;
assign w14993 = ~w13909 & w19712;
assign w14994 = ~pi352 & ~w14993;
assign w14995 = w13906 & w14842;
assign w14996 = w14842 & w19713;
assign w14997 = (~pi191 & ~w14039) | (~pi191 & w19714) | (~w14039 & w19714);
assign w14998 = ~w14996 & w14997;
assign w14999 = ~w14994 & w14998;
assign w15000 = pi352 & ~w14696;
assign w15001 = ~w13982 & ~w14851;
assign w15002 = w15000 & ~w15001;
assign w15003 = w13916 & w13947;
assign w15004 = ~pi352 & w15003;
assign w15005 = w13988 & w14044;
assign w15006 = ~w14005 & ~w15005;
assign w15007 = ~pi182 & ~w15006;
assign w15008 = ~w15004 & ~w15007;
assign w15009 = ~w13909 & ~w14820;
assign w15010 = ~w14031 & ~w14821;
assign w15011 = pi352 & w15010;
assign w15012 = w15009 & w15011;
assign w15013 = w13950 & w14008;
assign w15014 = w13905 & w13928;
assign w15015 = ~w14842 & ~w15013;
assign w15016 = w15015 & w19715;
assign w15017 = pi191 & ~w14737;
assign w15018 = pi182 & w14031;
assign w15019 = w15017 & ~w15018;
assign w15020 = (w15019 & w15012) | (w15019 & w19716) | (w15012 & w19716);
assign w15021 = pi321 & w13957;
assign w15022 = ~w14720 & ~w14856;
assign w15023 = ~w15021 & w15022;
assign w15024 = pi352 & ~w15023;
assign w15025 = w13928 & w13980;
assign w15026 = w13952 & w14004;
assign w15027 = ~w14786 & ~w15026;
assign w15028 = ~w14726 & w15027;
assign w15029 = w13938 & w15025;
assign w15030 = w15028 & ~w15029;
assign w15031 = ~w15024 & w15030;
assign w15032 = w15020 & w15031;
assign w15033 = ~w15002 & w15008;
assign w15034 = w14999 & w15033;
assign w15035 = ~w15032 & ~w15034;
assign w15036 = ~w14740 & ~w14820;
assign w15037 = (pi352 & ~w15036) | (pi352 & w19717) | (~w15036 & w19717);
assign w15038 = ~w13966 & ~w14816;
assign w15039 = (w13938 & ~w15038) | (w13938 & w19718) | (~w15038 & w19718);
assign w15040 = ~pi372 & ~w14715;
assign w15041 = ~w15039 & w15040;
assign w15042 = ~w15037 & w15041;
assign w15043 = (~pi352 & w13917) | (~pi352 & w19719) | (w13917 & w19719);
assign w15044 = ~w13916 & ~w13995;
assign w15045 = ~w14819 & ~w15044;
assign w15046 = pi352 & w13970;
assign w15047 = ~w13939 & ~w15046;
assign w15048 = ~w15045 & w15047;
assign w15049 = w14999 & w15048;
assign w15050 = ~w14734 & ~w15043;
assign w15051 = w15020 & w15050;
assign w15052 = ~w15049 & ~w15051;
assign w15053 = ~pi352 & ~w13935;
assign w15054 = ~w14835 & ~w15053;
assign w15055 = pi321 & w13930;
assign w15056 = w13979 & w15055;
assign w15057 = w13906 & w14023;
assign w15058 = (~pi342 & w15056) | (~pi342 & w19720) | (w15056 & w19720);
assign w15059 = ~pi170 & w13942;
assign w15060 = ~w15054 & ~w15058;
assign w15061 = (pi372 & ~w13942) | (pi372 & w19721) | (~w13942 & w19721);
assign w15062 = w15060 & w15061;
assign w15063 = ~w15035 & w15042;
assign w15064 = ~w15052 & w15062;
assign w15065 = ~w15063 & ~w15064;
assign w15066 = w13951 & w13979;
assign w15067 = (pi276 & w15066) | (pi276 & w19722) | (w15066 & w19722);
assign w15068 = ~w15065 & w19723;
assign w15069 = (~w14992 & w15065) | (~w14992 & w19724) | (w15065 & w19724);
assign w15070 = pi532 & pi573;
assign w15071 = ~w15068 & ~w15069;
assign w15072 = ~pi532 & w15071;
assign w15073 = ~w15070 & ~w15072;
assign w15074 = ~pi156 & pi224;
assign w15075 = pi156 & ~pi224;
assign w15076 = ~w15074 & ~w15075;
assign w15077 = ~pi228 & ~w15076;
assign w15078 = pi228 & w15076;
assign w15079 = ~w15077 & ~w15078;
assign w15080 = ~w14007 & ~w14027;
assign w15081 = ~w14044 & ~w14755;
assign w15082 = w15080 & w15081;
assign w15083 = pi372 & ~w15082;
assign w15084 = ~pi321 & w14694;
assign w15085 = ~w13907 & ~w15084;
assign w15086 = ~pi182 & ~w15085;
assign w15087 = ~w15021 & ~w15086;
assign w15088 = ~w15083 & w15087;
assign w15089 = pi352 & ~w15088;
assign w15090 = pi182 & w14720;
assign w15091 = (pi372 & ~w14720) | (pi372 & w19725) | (~w14720 & w19725);
assign w15092 = ~pi276 & w13939;
assign w15093 = w15091 & ~w15092;
assign w15094 = w13905 & ~w14004;
assign w15095 = ~w14816 & ~w15094;
assign w15096 = pi352 & ~w13913;
assign w15097 = (~pi352 & ~w13980) | (~pi352 & w19726) | (~w13980 & w19726);
assign w15098 = w15095 & w15097;
assign w15099 = ~w15096 & ~w15098;
assign w15100 = w13918 & w14040;
assign w15101 = ~w13942 & ~w15100;
assign w15102 = w13919 & w15101;
assign w15103 = ~pi372 & ~w15057;
assign w15104 = ~w15102 & w15103;
assign w15105 = ~w15099 & w15104;
assign w15106 = pi191 & ~w15013;
assign w15107 = ~w14041 & w15106;
assign w15108 = w13919 & w13976;
assign w15109 = w15107 & ~w15108;
assign w15110 = (w15109 & w15105) | (w15109 & w19727) | (w15105 & w19727);
assign w15111 = ~w13941 & ~w14819;
assign w15112 = ~pi352 & ~w15111;
assign w15113 = pi372 & ~w13977;
assign w15114 = ~w14793 & ~w15056;
assign w15115 = w15113 & w15114;
assign w15116 = w13916 & w19728;
assign w15117 = ~w14047 & w19729;
assign w15118 = (~w15117 & ~w15115) | (~w15117 & w19730) | (~w15115 & w19730);
assign w15119 = ~w14733 & ~w14800;
assign w15120 = (w14014 & ~w15119) | (w14014 & w19731) | (~w15119 & w19731);
assign w15121 = ~w13917 & ~w13970;
assign w15122 = w13976 & ~w15121;
assign w15123 = ~w13951 & ~w14009;
assign w15124 = w13938 & ~w15123;
assign w15125 = ~pi372 & w14821;
assign w15126 = ~pi191 & ~w14043;
assign w15127 = ~w15125 & w15126;
assign w15128 = ~w15124 & w15127;
assign w15129 = w15128 & w19732;
assign w15130 = ~w15118 & w15129;
assign w15131 = ~w15089 & w15110;
assign w15132 = ~w15130 & ~w15131;
assign w15133 = w13906 & ~w14004;
assign w15134 = (pi182 & ~w15006) | (pi182 & w19733) | (~w15006 & w19733);
assign w15135 = ~pi352 & ~w15134;
assign w15136 = ~pi182 & ~w15025;
assign w15137 = w15136 & w19734;
assign w15138 = ~w13970 & ~w14688;
assign w15139 = (w15138 & w15137) | (w15138 & w19735) | (w15137 & w19735);
assign w15140 = ~w15135 & ~w15139;
assign w15141 = ~pi321 & w13911;
assign w15142 = w14030 & w15141;
assign w15143 = ~w13935 & ~w15142;
assign w15144 = ~w15124 & w15143;
assign w15145 = ~pi372 & w15144;
assign w15146 = pi372 & ~w15140;
assign w15147 = w13952 & w13988;
assign w15148 = (w14035 & w15090) | (w14035 & w19736) | (w15090 & w19736);
assign w15149 = ~pi372 & w13979;
assign w15150 = w13905 & w13965;
assign w15151 = w13938 & w14714;
assign w15152 = w15149 & w15150;
assign w15153 = ~w15151 & ~w15152;
assign w15154 = w15003 & w19737;
assign w15155 = w15153 & ~w15154;
assign w15156 = ~w15148 & w15155;
assign w15157 = ~w15132 & w19738;
assign w15158 = w15079 & w15157;
assign w15159 = ~w15079 & ~w15157;
assign w15160 = pi532 & pi580;
assign w15161 = ~w15158 & ~w15159;
assign w15162 = ~pi532 & w15161;
assign w15163 = ~w15160 & ~w15162;
assign w15164 = ~pi149 & pi157;
assign w15165 = pi149 & ~pi157;
assign w15166 = ~w15164 & ~w15165;
assign w15167 = w13663 & w15166;
assign w15168 = ~w13663 & ~w15166;
assign w15169 = ~w15167 & ~w15168;
assign w15170 = (~w15169 & ~w13764) | (~w15169 & w19739) | (~w13764 & w19739);
assign w15171 = w13764 & w19740;
assign w15172 = pi532 & pi554;
assign w15173 = ~w15170 & ~w15171;
assign w15174 = ~pi532 & w15173;
assign w15175 = ~w15172 & ~w15174;
assign w15176 = ~pi270 & w4120;
assign w15177 = pi270 & ~w4120;
assign w15178 = ~w15176 & ~w15177;
assign w15179 = ~pi159 & pi269;
assign w15180 = pi159 & ~pi269;
assign w15181 = ~w15179 & ~w15180;
assign w15182 = ~pi352 & ~w15005;
assign w15183 = w13905 & w13947;
assign w15184 = ~w14030 & ~w15183;
assign w15185 = ~w15182 & ~w15184;
assign w15186 = ~pi372 & w13929;
assign w15187 = ~w13953 & ~w13990;
assign w15188 = ~w15186 & w15187;
assign w15189 = pi352 & ~w15188;
assign w15190 = ~w13931 & ~w14754;
assign w15191 = ~w15059 & w15190;
assign w15192 = ~pi352 & ~w15191;
assign w15193 = (w14040 & w14005) | (w14040 & w19741) | (w14005 & w19741);
assign w15194 = ~w15189 & ~w15192;
assign w15195 = pi191 & ~w15193;
assign w15196 = ~w13993 & ~w15003;
assign w15197 = ~pi352 & ~w15196;
assign w15198 = w13904 & ~w14822;
assign w15199 = ~w15197 & ~w15198;
assign w15200 = ~pi321 & w13930;
assign w15201 = pi352 & ~w14023;
assign w15202 = ~w15147 & ~w15200;
assign w15203 = w15201 & ~w15202;
assign w15204 = w13939 & w19742;
assign w15205 = (~pi191 & ~w14726) | (~pi191 & w19743) | (~w14726 & w19743);
assign w15206 = ~w15203 & w19744;
assign w15207 = ~pi352 & w14737;
assign w15208 = ~w15116 & ~w15207;
assign w15209 = ~w14843 & ~w15150;
assign w15210 = w15208 & w15209;
assign w15211 = w15206 & w15210;
assign w15212 = w15194 & w19745;
assign w15213 = ~w15211 & ~w15212;
assign w15214 = pi352 & ~w13970;
assign w15215 = w13980 & w13995;
assign w15216 = ~w15057 & ~w15215;
assign w15217 = ~w14740 & w15214;
assign w15218 = w15216 & w15217;
assign w15219 = w13918 & w15055;
assign w15220 = w14009 & w14023;
assign w15221 = ~w14696 & ~w15219;
assign w15222 = (~pi352 & ~w14009) | (~pi352 & w19746) | (~w14009 & w19746);
assign w15223 = w15221 & w15222;
assign w15224 = (~pi372 & ~w14704) | (~pi372 & w19747) | (~w14704 & w19747);
assign w15225 = ~w13976 & w14702;
assign w15226 = w15224 & ~w15225;
assign w15227 = ~w15218 & ~w15223;
assign w15228 = w15226 & ~w15227;
assign w15229 = ~w14026 & ~w15025;
assign w15230 = (~w14719 & ~w15229) | (~w14719 & w19748) | (~w15229 & w19748);
assign w15231 = ~w14036 & ~w14995;
assign w15232 = ~w15230 & w15231;
assign w15233 = w15194 & w19749;
assign w15234 = ~w14023 & w14851;
assign w15235 = ~w13958 & ~w14007;
assign w15236 = w13922 & w13979;
assign w15237 = w15235 & ~w15236;
assign w15238 = (~pi352 & w15234) | (~pi352 & w19750) | (w15234 & w19750);
assign w15239 = w15237 & ~w15238;
assign w15240 = w15206 & w15239;
assign w15241 = ~w15233 & ~w15240;
assign w15242 = ~w13998 & ~w15059;
assign w15243 = ~pi352 & ~w15242;
assign w15244 = ~w13916 & w14030;
assign w15245 = ~w15026 & ~w15244;
assign w15246 = ~pi170 & ~w15245;
assign w15247 = w13979 & w14816;
assign w15248 = ~w14794 & ~w15247;
assign w15249 = w15091 & ~w15246;
assign w15250 = ~w15243 & w15249;
assign w15251 = w15248 & w15250;
assign w15252 = ~w15213 & w15228;
assign w15253 = ~w15241 & w15251;
assign w15254 = ~w15252 & ~w15253;
assign w15255 = ~w15254 & w19751;
assign w15256 = (pi301 & w15254) | (pi301 & w19752) | (w15254 & w19752);
assign w15257 = ~w15255 & ~w15256;
assign w15258 = w15181 & ~w15257;
assign w15259 = ~w15181 & w15257;
assign w15260 = pi532 & pi577;
assign w15261 = ~w15258 & ~w15259;
assign w15262 = ~pi532 & w15261;
assign w15263 = ~w15260 & ~w15262;
assign w15264 = ~pi160 & ~w14153;
assign w15265 = pi160 & w14153;
assign w15266 = ~w15264 & ~w15265;
assign w15267 = pi532 & ~pi653;
assign w15268 = ~pi532 & ~w15266;
assign w15269 = ~w15267 & ~w15268;
assign w15270 = w13554 & w13608;
assign w15271 = (pi284 & ~w13608) | (pi284 & w19753) | (~w13608 & w19753);
assign w15272 = (pi351 & ~w13476) | (pi351 & w13541) | (~w13476 & w13541);
assign w15273 = ~w13474 & ~w13791;
assign w15274 = ~w13797 & w15272;
assign w15275 = w15273 & w15274;
assign w15276 = ~pi351 & ~w14133;
assign w15277 = ~w15275 & ~w15276;
assign w15278 = ~w13529 & ~w13791;
assign w15279 = (~pi351 & ~w15278) | (~pi351 & w19754) | (~w15278 & w19754);
assign w15280 = w13502 & w13571;
assign w15281 = w13509 & w13510;
assign w15282 = ~w13566 & ~w15281;
assign w15283 = pi351 & w13793;
assign w15284 = w13535 & w15282;
assign w15285 = ~w15283 & ~w15284;
assign w15286 = w13462 & ~w15280;
assign w15287 = w15285 & w19755;
assign w15288 = w15271 & ~w15277;
assign w15289 = ~w15287 & ~w15288;
assign w15290 = ~pi275 & w13592;
assign w15291 = ~w13572 & ~w13780;
assign w15292 = (~w13563 & w15291) | (~w13563 & w19756) | (w15291 & w19756);
assign w15293 = pi351 & ~w15292;
assign w15294 = w13554 & w13596;
assign w15295 = ~w14113 & ~w15294;
assign w15296 = w13544 & w13796;
assign w15297 = w15295 & ~w15296;
assign w15298 = ~w15293 & w15297;
assign w15299 = (pi193 & w15289) | (pi193 & w19757) | (w15289 & w19757);
assign w15300 = w13571 & ~w13592;
assign w15301 = (pi354 & w13791) | (pi354 & w19758) | (w13791 & w19758);
assign w15302 = ~w14137 & ~w15301;
assign w15303 = ~w13463 & ~w13605;
assign w15304 = (w15303 & w15302) | (w15303 & w19759) | (w15302 & w19759);
assign w15305 = pi351 & ~w15304;
assign w15306 = (w13562 & ~w14081) | (w13562 & w19760) | (~w14081 & w19760);
assign w15307 = w13554 & w13497;
assign w15308 = ~w13552 & ~w15307;
assign w15309 = ~pi351 & ~w15308;
assign w15310 = ~w14127 & ~w14491;
assign w15311 = pi284 & ~w14517;
assign w15312 = w15310 & w15311;
assign w15313 = ~w13591 & ~w13857;
assign w15314 = (~pi284 & ~w13560) | (~pi284 & w19761) | (~w13560 & w19761);
assign w15315 = w15313 & w15314;
assign w15316 = ~w15309 & w15312;
assign w15317 = ~w15315 & ~w15316;
assign w15318 = (pi351 & ~w13485) | (pi351 & w19762) | (~w13485 & w19762);
assign w15319 = ~w13779 & w15318;
assign w15320 = (~pi351 & ~w13592) | (~pi351 & w13508) | (~w13592 & w13508);
assign w15321 = ~w13792 & w15320;
assign w15322 = ~w15319 & ~w15321;
assign w15323 = pi157 & w13514;
assign w15324 = ~w13500 & ~w15323;
assign w15325 = w13544 & ~w15324;
assign w15326 = w13541 & w13602;
assign w15327 = ~w13564 & ~w15326;
assign w15328 = ~w15325 & w15327;
assign w15329 = ~w15322 & w15328;
assign w15330 = (~pi193 & w15317) | (~pi193 & w19763) | (w15317 & w19763);
assign w15331 = w13592 & w13823;
assign w15332 = ~w13472 & ~w15331;
assign w15333 = ~w15325 & w15332;
assign w15334 = ~pi284 & ~w15333;
assign w15335 = ~pi275 & w13604;
assign w15336 = ~w13580 & ~w15335;
assign w15337 = (w13850 & w15270) | (w13850 & w19764) | (w15270 & w19764);
assign w15338 = w13529 & w14088;
assign w15339 = ~w15337 & ~w15338;
assign w15340 = ~pi351 & ~w15336;
assign w15341 = w15339 & ~w15340;
assign w15342 = ~w15334 & w15341;
assign w15343 = ~w15330 & w15342;
assign w15344 = (pi284 & w15305) | (pi284 & w19765) | (w15305 & w19765);
assign w15345 = w15343 & w19766;
assign w15346 = ~pi392 & w15345;
assign w15347 = pi392 & ~w15345;
assign w15348 = ~w15346 & ~w15347;
assign w15349 = ~pi161 & ~w15348;
assign w15350 = pi161 & w15348;
assign w15351 = pi532 & pi660;
assign w15352 = ~w15349 & ~w15350;
assign w15353 = ~pi532 & w15352;
assign w15354 = ~w15351 & ~w15353;
assign w15355 = ~pi162 & ~w15266;
assign w15356 = pi162 & w15266;
assign w15357 = ~w15355 & ~w15356;
assign w15358 = ~pi161 & pi163;
assign w15359 = pi161 & ~pi163;
assign w15360 = ~w15358 & ~w15359;
assign w15361 = ~w15348 & ~w15360;
assign w15362 = w15348 & w15360;
assign w15363 = pi532 & pi628;
assign w15364 = ~w15361 & ~w15362;
assign w15365 = ~pi532 & w15364;
assign w15366 = ~w15363 & ~w15365;
assign w15367 = ~pi394 & ~w14156;
assign w15368 = pi394 & w14156;
assign w15369 = ~w15367 & ~w15368;
assign w15370 = ~pi162 & w14150;
assign w15371 = pi162 & ~w14150;
assign w15372 = ~w15370 & ~w15371;
assign w15373 = w15369 & ~w15372;
assign w15374 = ~w15369 & w15372;
assign w15375 = pi532 & pi589;
assign w15376 = ~w15373 & ~w15374;
assign w15377 = ~pi532 & w15376;
assign w15378 = ~w15375 & ~w15377;
assign w15379 = ~pi161 & pi165;
assign w15380 = pi161 & ~pi165;
assign w15381 = ~w15379 & ~w15380;
assign w15382 = ~pi392 & ~w15381;
assign w15383 = pi392 & w15381;
assign w15384 = ~w15382 & ~w15383;
assign w15385 = ~pi163 & w15345;
assign w15386 = pi163 & ~w15345;
assign w15387 = ~w15385 & ~w15386;
assign w15388 = ~w15384 & ~w15387;
assign w15389 = w15384 & w15387;
assign w15390 = pi532 & pi596;
assign w15391 = ~w15388 & ~w15389;
assign w15392 = ~pi532 & w15391;
assign w15393 = ~w15390 & ~w15392;
assign w15394 = ~pi163 & pi166;
assign w15395 = pi163 & ~pi166;
assign w15396 = ~w15394 & ~w15395;
assign w15397 = w15381 & w15396;
assign w15398 = ~w15381 & ~w15396;
assign w15399 = ~w15397 & ~w15398;
assign w15400 = w15348 & ~w15399;
assign w15401 = ~w15348 & w15399;
assign w15402 = pi532 & pi564;
assign w15403 = ~w15400 & ~w15401;
assign w15404 = ~pi532 & w15403;
assign w15405 = ~w15402 & ~w15404;
assign w15406 = w14348 & w19767;
assign w15407 = (pi167 & ~w14348) | (pi167 & w19768) | (~w14348 & w19768);
assign w15408 = ~w15406 & ~w15407;
assign w15409 = pi532 & ~pi634;
assign w15410 = ~pi532 & ~w15408;
assign w15411 = ~w15409 & ~w15410;
assign w15412 = ~pi168 & pi271;
assign w15413 = pi168 & ~pi271;
assign w15414 = ~w15412 & ~w15413;
assign w15415 = ~pi273 & ~w15414;
assign w15416 = pi273 & w15414;
assign w15417 = ~w15415 & ~w15416;
assign w15418 = (~w13294 & w13305) | (~w13294 & w19769) | (w13305 & w19769);
assign w15419 = pi231 & w13226;
assign w15420 = ~w13703 & ~w15419;
assign w15421 = ~w15418 & w15420;
assign w15422 = pi285 & ~w15421;
assign w15423 = w13249 & w13679;
assign w15424 = (pi231 & ~w13679) | (pi231 & w19770) | (~w13679 & w19770);
assign w15425 = w13182 & w13249;
assign w15426 = ~w13251 & ~w15425;
assign w15427 = ~pi231 & ~w13222;
assign w15428 = w13745 & w14913;
assign w15429 = w15427 & ~w15428;
assign w15430 = ~w14938 & w15424;
assign w15431 = w15426 & w15429;
assign w15432 = ~w15430 & ~w15431;
assign w15433 = w13189 & w13745;
assign w15434 = w13294 & w14942;
assign w15435 = w13237 & w13200;
assign w15436 = ~w15434 & ~w15435;
assign w15437 = w14952 & w15436;
assign w15438 = (~pi285 & ~w15437) | (~pi285 & w19771) | (~w15437 & w19771);
assign w15439 = ~w15432 & ~w15438;
assign w15440 = (~pi234 & ~w15439) | (~pi234 & w19772) | (~w15439 & w19772);
assign w15441 = ~pi231 & ~w14950;
assign w15442 = ~w13693 & w14968;
assign w15443 = w13283 & w15442;
assign w15444 = w13200 & w13679;
assign w15445 = ~w13289 & ~w14962;
assign w15446 = ~w15444 & w15445;
assign w15447 = pi231 & ~w15446;
assign w15448 = w13190 & w13740;
assign w15449 = ~w14903 & ~w15448;
assign w15450 = (pi285 & ~w13195) | (pi285 & w19773) | (~w13195 & w19773);
assign w15451 = w15449 & w15450;
assign w15452 = ~w15447 & w15451;
assign w15453 = w13190 & w14942;
assign w15454 = pi231 & ~w13688;
assign w15455 = ~w13698 & ~w15454;
assign w15456 = ~w15453 & w19774;
assign w15457 = w15455 & w15456;
assign w15458 = ~w15452 & ~w15457;
assign w15459 = w13183 & w13213;
assign w15460 = ~pi231 & ~w15459;
assign w15461 = w13203 & w13745;
assign w15462 = ~w13277 & ~w15461;
assign w15463 = pi231 & w15462;
assign w15464 = w15460 & w19775;
assign w15465 = ~w15463 & ~w15464;
assign w15466 = ~pi285 & ~w13202;
assign w15467 = ~w13241 & w15466;
assign w15468 = ~w15465 & w15467;
assign w15469 = ~pi270 & w15459;
assign w15470 = w13182 & w13281;
assign w15471 = ~w13204 & ~w15470;
assign w15472 = ~w15469 & w15471;
assign w15473 = (pi285 & ~w13755) | (pi285 & w19776) | (~w13755 & w19776);
assign w15474 = (w15473 & w15472) | (w15473 & w19777) | (w15472 & w19777);
assign w15475 = ~w15468 & ~w15474;
assign w15476 = (w13236 & w13306) | (w13236 & w19778) | (w13306 & w19778);
assign w15477 = ~w15476 & w19779;
assign w15478 = ~w15475 & w15477;
assign w15479 = (pi234 & w15458) | (pi234 & w19780) | (w15458 & w19780);
assign w15480 = w15478 & ~w15479;
assign w15481 = w15480 & w19781;
assign w15482 = (~w15417 & ~w15480) | (~w15417 & w19782) | (~w15480 & w19782);
assign w15483 = pi532 & pi587;
assign w15484 = ~w15481 & ~w15482;
assign w15485 = ~pi532 & w15484;
assign w15486 = ~w15483 & ~w15485;
assign w15487 = ~pi169 & pi272;
assign w15488 = pi169 & ~pi272;
assign w15489 = ~w15487 & ~w15488;
assign w15490 = ~pi274 & ~w15489;
assign w15491 = pi274 & w15489;
assign w15492 = ~w15490 & ~w15491;
assign w15493 = w14251 & w14284;
assign w15494 = ~w14259 & w14365;
assign w15495 = w14426 & w15494;
assign w15496 = ~w14195 & ~w15493;
assign w15497 = ~pi207 & w15496;
assign w15498 = (pi147 & w14390) | (pi147 & w19783) | (w14390 & w19783);
assign w15499 = (pi207 & w15498) | (pi207 & w19784) | (w15498 & w19784);
assign w15500 = (pi302 & ~w14303) | (pi302 & w19785) | (~w14303 & w19785);
assign w15501 = w14436 & w14637;
assign w15502 = ~w15501 & w19786;
assign w15503 = ~w14298 & ~w14371;
assign w15504 = pi207 & ~w15503;
assign w15505 = ~w14255 & ~w15504;
assign w15506 = w15502 & w15505;
assign w15507 = w14607 & w15500;
assign w15508 = ~w15499 & w15507;
assign w15509 = ~w15506 & ~w15508;
assign w15510 = (pi139 & w15509) | (pi139 & w19787) | (w15509 & w19787);
assign w15511 = ~pi138 & w14233;
assign w15512 = w14194 & w14270;
assign w15513 = ~w15511 & ~w15512;
assign w15514 = ~pi185 & ~w15513;
assign w15515 = pi207 & ~w14278;
assign w15516 = (~w14339 & w15514) | (~w14339 & w19788) | (w15514 & w19788);
assign w15517 = w14206 & w14412;
assign w15518 = ~pi207 & w14259;
assign w15519 = ~w15517 & ~w15518;
assign w15520 = w14232 & ~w14242;
assign w15521 = w15519 & ~w15520;
assign w15522 = ~pi139 & ~w15521;
assign w15523 = (w14200 & w14226) | (w14200 & w19789) | (w14226 & w19789);
assign w15524 = w14210 & w14637;
assign w15525 = ~pi129 & w14292;
assign w15526 = w14193 & w15525;
assign w15527 = ~w15493 & ~w15526;
assign w15528 = ~w14658 & ~w15524;
assign w15529 = w15527 & w15528;
assign w15530 = (~pi139 & ~w15529) | (~pi139 & w19790) | (~w15529 & w19790);
assign w15531 = ~pi207 & ~w14316;
assign w15532 = ~w14190 & w14256;
assign w15533 = w15531 & ~w15532;
assign w15534 = ~w14342 & w14428;
assign w15535 = ~w15533 & ~w15534;
assign w15536 = ~w14230 & ~w14392;
assign w15537 = ~w15535 & w15536;
assign w15538 = ~w15530 & w15537;
assign w15539 = ~w14215 & ~w14438;
assign w15540 = ~pi138 & ~w15539;
assign w15541 = ~pi207 & ~w14384;
assign w15542 = w14306 & w14599;
assign w15543 = w15541 & ~w15542;
assign w15544 = pi207 & ~w14633;
assign w15545 = ~w15526 & w15544;
assign w15546 = ~pi139 & ~w15545;
assign w15547 = ~w15540 & w15543;
assign w15548 = w15546 & ~w15547;
assign w15549 = ~pi207 & ~w14328;
assign w15550 = ~w14456 & ~w14587;
assign w15551 = (~w14404 & w15550) | (~w14404 & w19791) | (w15550 & w19791);
assign w15552 = ~w15548 & w15551;
assign w15553 = ~pi302 & ~w15538;
assign w15554 = w15552 & ~w15553;
assign w15555 = (pi302 & w15522) | (pi302 & w19792) | (w15522 & w19792);
assign w15556 = w15554 & w19793;
assign w15557 = w15492 & w15556;
assign w15558 = ~w15492 & ~w15556;
assign w15559 = pi532 & pi571;
assign w15560 = ~w15557 & ~w15558;
assign w15561 = ~pi532 & w15560;
assign w15562 = ~w15559 & ~w15561;
assign w15563 = ~pi170 & pi178;
assign w15564 = pi170 & ~pi178;
assign w15565 = ~w15563 & ~w15564;
assign w15566 = w14189 & w15565;
assign w15567 = ~w14189 & ~w15565;
assign w15568 = ~w15566 & ~w15567;
assign w15569 = (~w15568 & ~w14348) | (~w15568 & w19794) | (~w14348 & w19794);
assign w15570 = w14348 & w19795;
assign w15571 = pi532 & pi538;
assign w15572 = ~w15569 & ~w15570;
assign w15573 = ~pi532 & w15572;
assign w15574 = ~w15571 & ~w15573;
assign w15575 = ~w14022 & w19796;
assign w15576 = (pi171 & w14022) | (pi171 & w19797) | (w14022 & w19797);
assign w15577 = ~w15575 & ~w15576;
assign w15578 = pi532 & ~pi640;
assign w15579 = ~pi532 & ~w15577;
assign w15580 = ~w15578 & ~w15579;
assign w15581 = ~pi172 & ~w15577;
assign w15582 = pi172 & w15577;
assign w15583 = pi532 & pi608;
assign w15584 = ~w15581 & ~w15582;
assign w15585 = ~pi532 & w15584;
assign w15586 = ~w15583 & ~w15585;
assign w15587 = ~pi173 & pi278;
assign w15588 = pi173 & ~pi278;
assign w15589 = ~w15587 & ~w15588;
assign w15590 = ~pi281 & ~w15589;
assign w15591 = pi281 & w15589;
assign w15592 = ~w15590 & ~w15591;
assign w15593 = w13180 & w13194;
assign w15594 = pi231 & ~pi270;
assign w15595 = ~pi175 & w13289;
assign w15596 = w13670 & ~w15594;
assign w15597 = ~w15595 & ~w15596;
assign w15598 = ~w13736 & ~w15593;
assign w15599 = ~pi285 & w15598;
assign w15600 = w15597 & w15599;
assign w15601 = pi270 & w13197;
assign w15602 = ~w15433 & ~w15601;
assign w15603 = w13232 & w15602;
assign w15604 = pi231 & ~w15603;
assign w15605 = ~w13254 & ~w13695;
assign w15606 = ~w13254 & w19798;
assign w15607 = ~w15604 & w15606;
assign w15608 = ~w15600 & ~w15607;
assign w15609 = pi231 & ~w13680;
assign w15610 = w13213 & w13281;
assign w15611 = ~w13736 & ~w15610;
assign w15612 = ~w13677 & w15460;
assign w15613 = (~w15609 & ~w15612) | (~w15609 & w19799) | (~w15612 & w19799);
assign w15614 = ~w13679 & ~w14942;
assign w15615 = (pi234 & w15614) | (pi234 & w19800) | (w15614 & w19800);
assign w15616 = ~w15613 & w15615;
assign w15617 = ~w15608 & w15616;
assign w15618 = (~pi231 & w15444) | (~pi231 & w19801) | (w15444 & w19801);
assign w15619 = w13186 & w13265;
assign w15620 = w13243 & w14902;
assign w15621 = ~w13316 & ~w15620;
assign w15622 = ~w13309 & ~w15619;
assign w15623 = w15621 & w15622;
assign w15624 = pi270 & ~w13213;
assign w15625 = ~w13243 & w15624;
assign w15626 = (~w14956 & w15625) | (~w14956 & w19802) | (w15625 & w19802);
assign w15627 = (pi231 & w13257) | (pi231 & w19803) | (w13257 & w19803);
assign w15628 = w13732 & w19804;
assign w15629 = ~w15627 & w15628;
assign w15630 = ~pi231 & ~w15626;
assign w15631 = w15629 & ~w15630;
assign w15632 = w15623 & w19805;
assign w15633 = ~w15631 & ~w15632;
assign w15634 = (pi231 & w13725) | (pi231 & w19806) | (w13725 & w19806);
assign w15635 = w13277 & w13296;
assign w15636 = ~w13204 & ~w13304;
assign w15637 = ~w15635 & w15636;
assign w15638 = w15637 & w19807;
assign w15639 = ~w15634 & w15638;
assign w15640 = ~w15633 & w15639;
assign w15641 = ~w15617 & ~w15640;
assign w15642 = ~w13695 & ~w13702;
assign w15643 = pi175 & ~w15642;
assign w15644 = ~w13289 & ~w14942;
assign w15645 = ~pi175 & ~w15644;
assign w15646 = ~w13676 & w15441;
assign w15647 = ~w15645 & w15646;
assign w15648 = ~w13693 & w15647;
assign w15649 = ~w13306 & w19808;
assign w15650 = ~pi231 & ~w15649;
assign w15651 = ~w13196 & ~w13725;
assign w15652 = ~pi285 & w15651;
assign w15653 = ~w15650 & w15652;
assign w15654 = (pi285 & w15648) | (pi285 & w19809) | (w15648 & w19809);
assign w15655 = ~w13280 & w19810;
assign w15656 = w13303 & ~w15655;
assign w15657 = w13211 & w13295;
assign w15658 = ~w13318 & ~w15657;
assign w15659 = ~w15656 & w15658;
assign w15660 = (w15659 & w15654) | (w15659 & w19811) | (w15654 & w19811);
assign w15661 = ~w15641 & w19812;
assign w15662 = (~w15592 & w15641) | (~w15592 & w19813) | (w15641 & w19813);
assign w15663 = pi532 & pi582;
assign w15664 = ~w15661 & ~w15662;
assign w15665 = ~pi532 & w15664;
assign w15666 = ~w15663 & ~w15665;
assign w15667 = (~w14787 & ~w14742) | (~w14787 & w19814) | (~w14742 & w19814);
assign w15668 = (pi352 & w13998) | (pi352 & w19815) | (w13998 & w19815);
assign w15669 = ~w13970 & ~w14754;
assign w15670 = ~w15147 & w15669;
assign w15671 = ~w15668 & w15670;
assign w15672 = ~pi352 & ~w15667;
assign w15673 = w15671 & ~w15672;
assign w15674 = ~w13931 & ~w14737;
assign w15675 = pi352 & w15674;
assign w15676 = ~w14815 & w19816;
assign w15677 = ~w15675 & ~w15676;
assign w15678 = ~w14048 & ~w15220;
assign w15679 = (~pi372 & w15677) | (~pi372 & w19817) | (w15677 & w19817);
assign w15680 = ~w13909 & ~w15220;
assign w15681 = ~pi352 & ~w15680;
assign w15682 = w14732 & w19818;
assign w15683 = w13917 & w13979;
assign w15684 = w15101 & ~w15683;
assign w15685 = ~w15682 & w15684;
assign w15686 = ~w15681 & w15685;
assign w15687 = ~w15679 & w15686;
assign w15688 = pi372 & ~w15673;
assign w15689 = w15687 & ~w15688;
assign w15690 = pi182 & w13946;
assign w15691 = w13906 & w14739;
assign w15692 = ~w14040 & w15690;
assign w15693 = ~w15691 & ~w15692;
assign w15694 = ~w14704 & ~w15005;
assign w15695 = ~pi372 & w15694;
assign w15696 = w15693 & w15695;
assign w15697 = ~w14753 & ~w15055;
assign w15698 = (pi352 & ~w15697) | (pi352 & w19819) | (~w15697 & w19819);
assign w15699 = w13997 & ~w14688;
assign w15700 = ~w15698 & w15699;
assign w15701 = ~w15696 & ~w15700;
assign w15702 = ~w14695 & ~w14732;
assign w15703 = w14008 & ~w15702;
assign w15704 = ~w13977 & ~w14737;
assign w15705 = ~w14733 & w15704;
assign w15706 = (~w15000 & ~w15705) | (~w15000 & w19820) | (~w15705 & w19820);
assign w15707 = ~w15703 & ~w15706;
assign w15708 = ~w15701 & w15707;
assign w15709 = pi191 & ~w15708;
assign w15710 = ~w13941 & ~w14821;
assign w15711 = ~w14036 & w15710;
assign w15712 = ~pi352 & ~w15711;
assign w15713 = ~w14820 & ~w15215;
assign w15714 = (~pi372 & w15712) | (~pi372 & w19821) | (w15712 & w19821);
assign w15715 = w14694 & w14786;
assign w15716 = ~w14793 & ~w15715;
assign w15717 = (w14774 & ~w15716) | (w14774 & w19822) | (~w15716 & w19822);
assign w15718 = ~w13928 & w14701;
assign w15719 = ~w14714 & ~w15718;
assign w15720 = (w14743 & ~w15719) | (w14743 & w19823) | (~w15719 & w19823);
assign w15721 = ~w14800 & ~w15025;
assign w15722 = w14014 & ~w15721;
assign w15723 = ~w13967 & ~w14716;
assign w15724 = (w15149 & ~w15723) | (w15149 & w19824) | (~w15723 & w19824);
assign w15725 = ~w15717 & ~w15720;
assign w15726 = ~w15722 & ~w15724;
assign w15727 = w15725 & w15726;
assign w15728 = ~w15714 & w15727;
assign w15729 = ~w15709 & w15728;
assign w15730 = ~pi191 & ~w15689;
assign w15731 = w15729 & ~w15730;
assign w15732 = ~pi174 & pi280;
assign w15733 = pi174 & ~pi280;
assign w15734 = ~w15732 & ~w15733;
assign w15735 = ~pi283 & ~w15734;
assign w15736 = pi283 & w15734;
assign w15737 = ~w15735 & ~w15736;
assign w15738 = w15731 & w15737;
assign w15739 = ~w15731 & ~w15737;
assign w15740 = pi532 & pi574;
assign w15741 = ~w15738 & ~w15739;
assign w15742 = ~pi532 & w15741;
assign w15743 = ~w15740 & ~w15742;
assign w15744 = ~pi175 & w13903;
assign w15745 = pi175 & ~w13903;
assign w15746 = ~w15744 & ~w15745;
assign w15747 = ~w14022 & w19825;
assign w15748 = (w15746 & w14022) | (w15746 & w19826) | (w14022 & w19826);
assign w15749 = pi532 & pi544;
assign w15750 = ~w15747 & ~w15748;
assign w15751 = ~pi532 & w15750;
assign w15752 = ~w15749 & ~w15751;
assign w15753 = w10331 & w19827;
assign w15754 = (pi141 & ~w10331) | (pi141 & w19828) | (~w10331 & w19828);
assign w15755 = ~w15753 & ~w15754;
assign w15756 = ~pi159 & w5243;
assign w15757 = pi159 & ~w5243;
assign w15758 = ~w15756 & ~w15757;
assign w15759 = pi178 & ~w15408;
assign w15760 = ~pi178 & w15408;
assign w15761 = pi532 & pi602;
assign w15762 = ~w15759 & ~w15760;
assign w15763 = ~pi532 & w15762;
assign w15764 = ~w15761 & ~w15763;
assign w15765 = ~pi179 & pi223;
assign w15766 = pi179 & ~pi223;
assign w15767 = ~w15765 & ~w15766;
assign w15768 = w13956 & w13912;
assign w15769 = ~w13908 & ~w15768;
assign w15770 = (~pi352 & ~w15769) | (~pi352 & w19829) | (~w15769 & w19829);
assign w15771 = ~w13959 & ~w15150;
assign w15772 = ~pi342 & ~w15771;
assign w15773 = pi372 & ~w15147;
assign w15774 = ~w13994 & w15773;
assign w15775 = ~w13947 & ~w14014;
assign w15776 = w13933 & ~w15775;
assign w15777 = ~w15772 & w15774;
assign w15778 = ~w14696 & ~w15776;
assign w15779 = w15777 & w15778;
assign w15780 = w13980 & w14040;
assign w15781 = pi182 & ~w15780;
assign w15782 = ~w15116 & w15136;
assign w15783 = (~pi372 & ~w13959) | (~pi372 & w19830) | (~w13959 & w19830);
assign w15784 = (w15783 & w15782) | (w15783 & w19831) | (w15782 & w19831);
assign w15785 = (~w15784 & ~w15779) | (~w15784 & w19832) | (~w15779 & w19832);
assign w15786 = pi352 & ~w14716;
assign w15787 = ~w15219 & w15786;
assign w15788 = pi182 & ~w14798;
assign w15789 = w15787 & ~w15788;
assign w15790 = w14829 & w14844;
assign w15791 = (~w14800 & w15789) | (~w14800 & w19833) | (w15789 & w19833);
assign w15792 = (~pi191 & w15785) | (~pi191 & w19834) | (w15785 & w19834);
assign w15793 = ~w13953 & ~w13957;
assign w15794 = ~w15214 & ~w15793;
assign w15795 = ~w15003 & ~w15200;
assign w15796 = pi352 & ~w15795;
assign w15797 = (~pi372 & ~w14009) | (~pi372 & w19835) | (~w14009 & w19835);
assign w15798 = ~w15794 & ~w15796;
assign w15799 = w15797 & w15798;
assign w15800 = pi372 & ~w15026;
assign w15801 = ~w14036 & w15800;
assign w15802 = w15009 & w15801;
assign w15803 = ~w13928 & w14822;
assign w15804 = ~w13951 & ~w14720;
assign w15805 = w15669 & w15804;
assign w15806 = (pi372 & w15803) | (pi372 & w19836) | (w15803 & w19836);
assign w15807 = w15805 & ~w15806;
assign w15808 = ~w14798 & w19837;
assign w15809 = ~w13971 & ~w15808;
assign w15810 = ~pi352 & ~w15807;
assign w15811 = w15809 & ~w15810;
assign w15812 = ~w15799 & ~w15802;
assign w15813 = w15811 & ~w15812;
assign w15814 = w13906 & w13947;
assign w15815 = ~w14010 & ~w15814;
assign w15816 = ~w13968 & w14008;
assign w15817 = w15815 & ~w15816;
assign w15818 = pi352 & ~w15817;
assign w15819 = ~w13970 & ~w14695;
assign w15820 = w13976 & ~w15819;
assign w15821 = w13938 & w13993;
assign w15822 = w13943 & ~w15821;
assign w15823 = (pi372 & ~w13917) | (pi372 & w19838) | (~w13917 & w19838);
assign w15824 = ~pi352 & w13929;
assign w15825 = w15823 & ~w15824;
assign w15826 = ~w15820 & w15822;
assign w15827 = (~w15825 & w15818) | (~w15825 & w19839) | (w15818 & w19839);
assign w15828 = w13991 & w14774;
assign w15829 = ~w15682 & ~w15828;
assign w15830 = ~w13940 & ~w14764;
assign w15831 = w15829 & w15830;
assign w15832 = ~w15827 & w15831;
assign w15833 = pi191 & ~w15813;
assign w15834 = ~w15833 & w19840;
assign w15835 = ~pi226 & w15834;
assign w15836 = pi226 & ~w15834;
assign w15837 = ~w15835 & ~w15836;
assign w15838 = ~w15767 & ~w15837;
assign w15839 = w15767 & w15837;
assign w15840 = pi532 & pi578;
assign w15841 = ~w15838 & ~w15839;
assign w15842 = ~pi532 & w15841;
assign w15843 = ~w15840 & ~w15842;
assign w15844 = ~w14460 & w19841;
assign w15845 = (pi181 & w14460) | (pi181 & w19842) | (w14460 & w19842);
assign w15846 = ~w15844 & ~w15845;
assign w15847 = ~pi180 & ~w15846;
assign w15848 = pi180 & w15846;
assign w15849 = pi532 & pi600;
assign w15850 = ~w15847 & ~w15848;
assign w15851 = ~pi532 & w15850;
assign w15852 = ~w15849 & ~w15851;
assign w15853 = pi532 & ~pi632;
assign w15854 = ~pi532 & ~w15846;
assign w15855 = ~w15853 & ~w15854;
assign w15856 = ~pi182 & w14363;
assign w15857 = pi182 & ~w14363;
assign w15858 = ~w15856 & ~w15857;
assign w15859 = ~w14460 & w19843;
assign w15860 = (w15858 & w14460) | (w15858 & w19844) | (w14460 & w19844);
assign w15861 = pi532 & pi536;
assign w15862 = ~w15859 & ~w15860;
assign w15863 = ~pi532 & w15862;
assign w15864 = ~w15861 & ~w15863;
assign w15865 = ~pi183 & pi319;
assign w15866 = pi183 & ~pi319;
assign w15867 = ~w15865 & ~w15866;
assign w15868 = ~pi320 & ~w15867;
assign w15869 = pi320 & w15867;
assign w15870 = ~w15868 & ~w15869;
assign w15871 = ~w14233 & w14249;
assign w15872 = ~w14231 & ~w14663;
assign w15873 = (~pi207 & ~w15872) | (~pi207 & w19845) | (~w15872 & w19845);
assign w15874 = w14249 & w14293;
assign w15875 = pi185 & w14191;
assign w15876 = w14232 & w15875;
assign w15877 = ~w15524 & ~w15876;
assign w15878 = ~w14616 & ~w15874;
assign w15879 = w15877 & w15878;
assign w15880 = pi302 & w15879;
assign w15881 = ~w14424 & ~w15511;
assign w15882 = w14194 & w14306;
assign w15883 = ~w14372 & ~w14648;
assign w15884 = ~w15882 & w15883;
assign w15885 = w14329 & w14427;
assign w15886 = pi129 & w14328;
assign w15887 = w14202 & ~w14240;
assign w15888 = w14436 & w15887;
assign w15889 = ~w15886 & ~w15888;
assign w15890 = ~w15517 & ~w15885;
assign w15891 = w15889 & w15890;
assign w15892 = ~pi302 & w15891;
assign w15893 = (pi207 & ~w15884) | (pi207 & w19846) | (~w15884 & w19846);
assign w15894 = w15892 & ~w15893;
assign w15895 = ~w15873 & w15880;
assign w15896 = ~w15894 & ~w15895;
assign w15897 = ~pi207 & ~w14630;
assign w15898 = w14209 & w14213;
assign w15899 = ~w14329 & ~w15898;
assign w15900 = ~w15897 & ~w15899;
assign w15901 = w14270 & ~w14303;
assign w15902 = ~w14629 & ~w15901;
assign w15903 = (pi207 & ~w14196) | (pi207 & w19847) | (~w14196 & w19847);
assign w15904 = ~pi207 & ~w14437;
assign w15905 = (~w15903 & ~w15904) | (~w15903 & w19848) | (~w15904 & w19848);
assign w15906 = w14280 & ~w14338;
assign w15907 = ~w15905 & w15906;
assign w15908 = ~pi302 & ~w14326;
assign w15909 = w15902 & w15908;
assign w15910 = ~w15907 & ~w15909;
assign w15911 = ~w14663 & w15541;
assign w15912 = ~w14290 & w15911;
assign w15913 = ~w14244 & w14428;
assign w15914 = ~w15912 & ~w15913;
assign w15915 = ~w14662 & w19849;
assign w15916 = w14257 & w14448;
assign w15917 = w15915 & ~w15916;
assign w15918 = w14256 & ~w14306;
assign w15919 = w14232 & w14305;
assign w15920 = ~w14624 & ~w15919;
assign w15921 = pi302 & ~w14425;
assign w15922 = w15920 & w15921;
assign w15923 = (~pi207 & w15918) | (~pi207 & w19850) | (w15918 & w19850);
assign w15924 = w15922 & ~w15923;
assign w15925 = w14233 & w19639;
assign w15926 = w14213 & w19847;
assign w15927 = w14217 & w14436;
assign w15928 = ~w15926 & ~w15927;
assign w15929 = ~w14342 & ~w15925;
assign w15930 = w15928 & w19851;
assign w15931 = pi138 & ~w14234;
assign w15932 = w14267 & ~w15931;
assign w15933 = w15525 & w19852;
assign w15934 = (~pi139 & ~w14328) | (~pi139 & w19853) | (~w14328 & w19853);
assign w15935 = ~w15933 & w15934;
assign w15936 = ~w15932 & w15935;
assign w15937 = ~w15924 & ~w15930;
assign w15938 = w15936 & ~w15937;
assign w15939 = ~w15914 & w15917;
assign w15940 = ~w15910 & w15939;
assign w15941 = ~w15938 & ~w15940;
assign w15942 = ~w15941 & w19854;
assign w15943 = w15870 & w15942;
assign w15944 = ~w15870 & ~w15942;
assign w15945 = pi532 & pi569;
assign w15946 = ~w15943 & ~w15944;
assign w15947 = ~pi532 & w15946;
assign w15948 = ~w15945 & ~w15947;
assign w15949 = ~w13818 & ~w14134;
assign w15950 = ~w13463 & ~w15280;
assign w15951 = w15949 & w19855;
assign w15952 = pi351 & ~w15951;
assign w15953 = pi132 & w13593;
assign w15954 = w13593 & w13562;
assign w15955 = ~pi275 & w14095;
assign w15956 = ~w13510 & w13554;
assign w15957 = w13544 & w15956;
assign w15958 = ~w15955 & ~w15957;
assign w15959 = (~pi284 & ~w14501) | (~pi284 & w19856) | (~w14501 & w19856);
assign w15960 = w15958 & w19857;
assign w15961 = ~w13781 & ~w14131;
assign w15962 = ~pi351 & ~w15961;
assign w15963 = ~w13823 & ~w14126;
assign w15964 = ~w13476 & ~w15963;
assign w15965 = w14495 & w15271;
assign w15966 = ~w15964 & w15965;
assign w15967 = ~w15962 & w15966;
assign w15968 = ~w15952 & w15960;
assign w15969 = ~w15967 & ~w15968;
assign w15970 = ~w13478 & ~w13560;
assign w15971 = ~pi351 & ~w15970;
assign w15972 = (~pi284 & w13505) | (~pi284 & w19858) | (w13505 & w19858);
assign w15973 = (pi351 & ~w13592) | (pi351 & w19762) | (~w13592 & w19762);
assign w15974 = (~pi351 & ~w13459) | (~pi351 & w19859) | (~w13459 & w19859);
assign w15975 = ~w13553 & w15974;
assign w15976 = ~w15973 & ~w15975;
assign w15977 = ~w13490 & w14132;
assign w15978 = ~w15976 & w15977;
assign w15979 = ~w15971 & w15972;
assign w15980 = ~w15978 & ~w15979;
assign w15981 = ~w13498 & ~w13813;
assign w15982 = ~w14131 & w15981;
assign w15983 = ~pi351 & ~w15982;
assign w15984 = (w15973 & w14087) | (w15973 & w20903) | (w14087 & w20903);
assign w15985 = ~w13597 & ~w14125;
assign w15986 = pi193 & ~w14126;
assign w15987 = w15985 & w15986;
assign w15988 = ~w15984 & w15987;
assign w15989 = ~w15983 & w15988;
assign w15990 = ~w15980 & w15989;
assign w15991 = ~w13502 & w13525;
assign w15992 = w13459 & w19860;
assign w15993 = w13504 & w13509;
assign w15994 = ~w15992 & ~w15993;
assign w15995 = pi284 & ~w13797;
assign w15996 = w15994 & w15995;
assign w15997 = (~pi351 & w15991) | (~pi351 & w19861) | (w15991 & w19861);
assign w15998 = w15996 & ~w15997;
assign w15999 = ~w13462 & ~w13853;
assign w16000 = w13533 & ~w13591;
assign w16001 = ~w15999 & w16000;
assign w16002 = (pi132 & ~w13476) | (pi132 & w19511) | (~w13476 & w19511);
assign w16003 = ~w13479 & w19862;
assign w16004 = w13516 & w13544;
assign w16005 = (~pi193 & ~w14095) | (~pi193 & w19863) | (~w14095 & w19863);
assign w16006 = ~w16003 & w19864;
assign w16007 = (w16006 & w15998) | (w16006 & w20904) | (w15998 & w20904);
assign w16008 = ~w15990 & ~w16007;
assign w16009 = ~pi351 & ~w14080;
assign w16010 = ~w13562 & ~w14501;
assign w16011 = ~w16009 & ~w16010;
assign w16012 = ~w16008 & w19865;
assign w16013 = ~pi184 & w16012;
assign w16014 = pi184 & ~w16012;
assign w16015 = ~w16013 & ~w16014;
assign w16016 = ~pi255 & pi384;
assign w16017 = pi255 & ~pi384;
assign w16018 = ~w16016 & ~w16017;
assign w16019 = w16015 & w16018;
assign w16020 = ~w16015 & ~w16018;
assign w16021 = ~w16019 & ~w16020;
assign w16022 = pi532 & pi625;
assign w16023 = ~pi532 & ~w16021;
assign w16024 = ~w16022 & ~w16023;
assign w16025 = ~pi185 & pi221;
assign w16026 = pi185 & ~pi221;
assign w16027 = ~w16025 & ~w16026;
assign w16028 = w16021 & w16027;
assign w16029 = ~w16021 & ~w16027;
assign w16030 = pi532 & pi561;
assign w16031 = ~w16028 & ~w16029;
assign w16032 = ~pi532 & w16031;
assign w16033 = ~w16030 & ~w16032;
assign w16034 = w9311 & w19866;
assign w16035 = (pi144 & ~w9311) | (pi144 & w19867) | (~w9311 & w19867);
assign w16036 = ~w16034 & ~w16035;
assign w16037 = w14672 & w19868;
assign w16038 = (pi187 & ~w14672) | (pi187 & w19869) | (~w14672 & w19869);
assign w16039 = ~w16037 & ~w16038;
assign w16040 = pi532 & ~pi629;
assign w16041 = ~pi532 & ~w16039;
assign w16042 = ~w16040 & ~w16041;
assign w16043 = w7377 & w19870;
assign w16044 = (pi140 & ~w7377) | (pi140 & w19871) | (~w7377 & w19871);
assign w16045 = ~w16043 & ~w16044;
assign w16046 = ~w14949 & w19872;
assign w16047 = (pi189 & w14949) | (pi189 & w19873) | (w14949 & w19873);
assign w16048 = ~w16046 & ~w16047;
assign w16049 = pi532 & ~pi645;
assign w16050 = ~pi532 & ~w16048;
assign w16051 = ~w16049 & ~w16050;
assign w16052 = pi190 & ~w16039;
assign w16053 = ~pi190 & w16039;
assign w16054 = pi532 & pi597;
assign w16055 = ~w16052 & ~w16053;
assign w16056 = ~pi532 & w16055;
assign w16057 = ~w16054 & ~w16056;
assign w16058 = ~pi190 & pi191;
assign w16059 = pi190 & ~pi191;
assign w16060 = ~w16058 & ~w16059;
assign w16061 = w14586 & w16060;
assign w16062 = ~w14586 & ~w16060;
assign w16063 = ~w16061 & ~w16062;
assign w16064 = (~w16063 & ~w14672) | (~w16063 & w19874) | (~w14672 & w19874);
assign w16065 = w14672 & w19875;
assign w16066 = pi532 & pi533;
assign w16067 = ~w16064 & ~w16065;
assign w16068 = ~pi532 & w16067;
assign w16069 = ~w16066 & ~w16068;
assign w16070 = pi192 & ~w16048;
assign w16071 = ~pi192 & w16048;
assign w16072 = pi532 & pi613;
assign w16073 = ~w16070 & ~w16071;
assign w16074 = ~pi532 & w16073;
assign w16075 = ~w16072 & ~w16074;
assign w16076 = ~pi192 & pi193;
assign w16077 = pi192 & ~pi193;
assign w16078 = ~w16076 & ~w16077;
assign w16079 = w14887 & w16078;
assign w16080 = ~w14887 & ~w16078;
assign w16081 = ~w16079 & ~w16080;
assign w16082 = (~w16081 & w14949) | (~w16081 & w19876) | (w14949 & w19876);
assign w16083 = ~w14949 & w19877;
assign w16084 = pi532 & pi549;
assign w16085 = ~w16082 & ~w16083;
assign w16086 = ~pi532 & w16085;
assign w16087 = ~w16084 & ~w16086;
assign w16088 = w10244 & w19878;
assign w16089 = (pi167 & ~w10244) | (pi167 & w19879) | (~w10244 & w19879);
assign w16090 = ~w16088 & ~w16089;
assign w16091 = ~pi269 & w6786;
assign w16092 = pi269 & ~w6786;
assign w16093 = ~w16091 & ~w16092;
assign w16094 = w246 & w19880;
assign w16095 = (pi137 & ~w246) | (pi137 & w19881) | (~w246 & w19881);
assign w16096 = ~w16094 & ~w16095;
assign w16097 = ~w10148 & w19882;
assign w16098 = (pi223 & w10148) | (pi223 & w19883) | (w10148 & w19883);
assign w16099 = ~w16097 & ~w16098;
assign w16100 = ~pi148 & w10092;
assign w16101 = pi148 & ~w10092;
assign w16102 = ~w16100 & ~w16101;
assign w16103 = ~pi301 & w9148;
assign w16104 = pi301 & ~w9148;
assign w16105 = ~w16103 & ~w16104;
assign w16106 = ~w6235 & w19884;
assign w16107 = (pi224 & w6235) | (pi224 & w19885) | (w6235 & w19885);
assign w16108 = ~w16106 & ~w16107;
assign w16109 = ~pi154 & w1282;
assign w16110 = pi154 & ~w1282;
assign w16111 = ~w16109 & ~w16110;
assign w16112 = ~pi192 & w2041;
assign w16113 = pi192 & ~w2041;
assign w16114 = ~w16112 & ~w16113;
assign w16115 = ~pi189 & w2942;
assign w16116 = pi189 & ~w2942;
assign w16117 = ~w16115 & ~w16116;
assign w16118 = ~pi152 & w7445;
assign w16119 = pi152 & ~w7445;
assign w16120 = ~w16118 & ~w16119;
assign w16121 = ~pi145 & w10456;
assign w16122 = pi145 & ~w10456;
assign w16123 = ~w16121 & ~w16122;
assign w16124 = ~pi231 & w8232;
assign w16125 = pi231 & ~w8232;
assign w16126 = ~w16124 & ~w16125;
assign w16127 = ~pi207 & pi209;
assign w16128 = pi207 & ~pi209;
assign w16129 = ~w16127 & ~w16128;
assign w16130 = ~w13535 & w15973;
assign w16131 = ~w14525 & ~w16130;
assign w16132 = ~w13855 & ~w14095;
assign w16133 = w16132 & w19886;
assign w16134 = (~pi284 & ~w19887) | (~pi284 & w20905) | (~w19887 & w20905);
assign w16135 = w13476 & w19888;
assign w16136 = (pi284 & w14141) | (pi284 & w19889) | (w14141 & w19889);
assign w16137 = ~w13556 & ~w15323;
assign w16138 = (w13541 & ~w16137) | (w13541 & w19890) | (~w16137 & w19890);
assign w16139 = ~w13775 & ~w13791;
assign w16140 = w13460 & w13509;
assign w16141 = ~w14134 & ~w15955;
assign w16142 = ~w16140 & w16141;
assign w16143 = w13508 & ~w16139;
assign w16144 = w16142 & w19891;
assign w16145 = ~w16138 & w16144;
assign w16146 = ~w13511 & ~w13777;
assign w16147 = w14111 & w16146;
assign w16148 = ~w13498 & w15272;
assign w16149 = (~w14517 & w16147) | (~w14517 & w19892) | (w16147 & w19892);
assign w16150 = pi284 & ~w16149;
assign w16151 = (pi358 & w13854) | (pi358 & w19893) | (w13854 & w19893);
assign w16152 = w13484 & w13562;
assign w16153 = ~w13472 & ~w16152;
assign w16154 = ~pi284 & ~w16153;
assign w16155 = ~w13540 & ~w16154;
assign w16156 = ~w16151 & w16155;
assign w16157 = ~w16150 & w16156;
assign w16158 = ~pi193 & ~w16157;
assign w16159 = ~w13831 & ~w14137;
assign w16160 = (~pi351 & ~w16159) | (~pi351 & w19894) | (~w16159 & w19894);
assign w16161 = (w13541 & w13593) | (w13541 & w19895) | (w13593 & w19895);
assign w16162 = w13464 & ~w13510;
assign w16163 = ~w13550 & w16162;
assign w16164 = w13471 & w13509;
assign w16165 = ~w16163 & ~w16164;
assign w16166 = ~w14471 & ~w16161;
assign w16167 = w16165 & w16166;
assign w16168 = ~w13605 & ~w13779;
assign w16169 = ~pi275 & w13786;
assign w16170 = w13786 & w19524;
assign w16171 = ~w13584 & ~w16170;
assign w16172 = pi351 & ~w13584;
assign w16173 = w13502 & w13607;
assign w16174 = ~w16173 & w19896;
assign w16175 = w14528 & ~w16174;
assign w16176 = w13539 & w15281;
assign w16177 = ~w13844 & w19897;
assign w16178 = ~w16175 & w16177;
assign w16179 = (pi284 & w13584) | (pi284 & w13508) | (w13584 & w13508);
assign w16180 = (w16179 & ~w16168) | (w16179 & w19898) | (~w16168 & w19898);
assign w16181 = w16178 & ~w16180;
assign w16182 = (~pi284 & ~w16167) | (~pi284 & w20906) | (~w16167 & w20906);
assign w16183 = w16181 & ~w16182;
assign w16184 = ~w16158 & w16183;
assign w16185 = (pi193 & ~w16145) | (pi193 & w20907) | (~w16145 & w20907);
assign w16186 = w16184 & ~w16185;
assign w16187 = ~pi210 & pi385;
assign w16188 = pi210 & ~pi385;
assign w16189 = ~w16187 & ~w16188;
assign w16190 = (w16189 & ~w16184) | (w16189 & w20908) | (~w16184 & w20908);
assign w16191 = w16184 & w20909;
assign w16192 = ~w16190 & ~w16191;
assign w16193 = ~pi208 & ~w16192;
assign w16194 = pi208 & w16192;
assign w16195 = ~w16193 & ~w16194;
assign w16196 = w16129 & ~w16195;
assign w16197 = ~w16129 & w16195;
assign w16198 = pi532 & pi559;
assign w16199 = ~w16196 & ~w16197;
assign w16200 = ~pi532 & w16199;
assign w16201 = ~w16198 & ~w16200;
assign w16202 = pi532 & ~pi623;
assign w16203 = ~pi532 & ~w16195;
assign w16204 = ~w16202 & ~w16203;
assign w16205 = ~pi208 & w16186;
assign w16206 = pi208 & ~w16186;
assign w16207 = ~w16205 & ~w16206;
assign w16208 = ~pi209 & pi210;
assign w16209 = pi209 & ~pi210;
assign w16210 = ~w16208 & ~w16209;
assign w16211 = ~pi385 & ~w16210;
assign w16212 = pi385 & w16210;
assign w16213 = ~w16211 & ~w16212;
assign w16214 = ~w16207 & ~w16213;
assign w16215 = w16207 & w16213;
assign w16216 = pi532 & pi591;
assign w16217 = ~w16214 & ~w16215;
assign w16218 = ~pi532 & w16217;
assign w16219 = ~w16216 & ~w16218;
assign w16220 = pi532 & pi655;
assign w16221 = ~pi532 & ~w16192;
assign w16222 = ~w16220 & ~w16221;
assign w16223 = ~pi191 & w7034;
assign w16224 = pi191 & ~w7034;
assign w16225 = ~w16223 & ~w16224;
assign w16226 = ~pi321 & w4276;
assign w16227 = pi321 & ~w4276;
assign w16228 = ~w16226 & ~w16227;
assign w16229 = ~pi276 & w11044;
assign w16230 = pi276 & ~w11044;
assign w16231 = ~w16229 & ~w16230;
assign w16232 = w8340 & w19899;
assign w16233 = (pi150 & ~w8340) | (pi150 & w19900) | (~w8340 & w19900);
assign w16234 = ~w16232 & ~w16233;
assign w16235 = ~pi215 & ~w14869;
assign w16236 = pi215 & w14869;
assign w16237 = pi532 & pi547;
assign w16238 = ~w16235 & ~w16236;
assign w16239 = ~pi532 & w16238;
assign w16240 = ~w16237 & ~w16239;
assign w16241 = w9700 & w19901;
assign w16242 = (pi190 & ~w9700) | (pi190 & w19902) | (~w9700 & w19902);
assign w16243 = ~w16241 & ~w16242;
assign w16244 = ~pi217 & pi371;
assign w16245 = pi217 & ~pi371;
assign w16246 = ~w16244 & ~w16245;
assign w16247 = ~pi346 & ~w16246;
assign w16248 = pi346 & w16246;
assign w16249 = ~w16247 & ~w16248;
assign w16250 = ~w13186 & ~w13210;
assign w16251 = (pi231 & ~w13237) | (pi231 & w13236) | (~w13237 & w13236);
assign w16252 = w16250 & w16251;
assign w16253 = ~w13204 & w13705;
assign w16254 = ~w16252 & ~w16253;
assign w16255 = ~w13181 & ~w14942;
assign w16256 = (~w14924 & ~w16255) | (~w14924 & w19903) | (~w16255 & w19903);
assign w16257 = (~pi285 & w16254) | (~pi285 & w19904) | (w16254 & w19904);
assign w16258 = (pi285 & w13690) | (pi285 & w13741) | (w13690 & w13741);
assign w16259 = w14955 & ~w15625;
assign w16260 = ~w13253 & ~w13315;
assign w16261 = (w13294 & ~w16260) | (w13294 & w19905) | (~w16260 & w19905);
assign w16262 = ~pi215 & w14895;
assign w16263 = ~w14958 & ~w16262;
assign w16264 = ~w16261 & w16263;
assign w16265 = ~w15619 & w16264;
assign w16266 = ~w16257 & w16265;
assign w16267 = (pi234 & ~w16266) | (pi234 & w19906) | (~w16266 & w19906);
assign w16268 = pi270 & w14956;
assign w16269 = ~w13680 & ~w16268;
assign w16270 = w15605 & w16269;
assign w16271 = ~w15609 & ~w16270;
assign w16272 = ~w13731 & ~w14889;
assign w16273 = pi231 & ~w16272;
assign w16274 = ~pi231 & ~w13180;
assign w16275 = ~w13243 & ~w13248;
assign w16276 = w16274 & ~w16275;
assign w16277 = ~w15459 & ~w16276;
assign w16278 = ~w16273 & w16277;
assign w16279 = ~pi234 & ~w16278;
assign w16280 = pi233 & w13200;
assign w16281 = ~w13704 & ~w16280;
assign w16282 = w13198 & w13715;
assign w16283 = w16281 & ~w16282;
assign w16284 = pi231 & ~w16283;
assign w16285 = ~w16279 & ~w16284;
assign w16286 = (pi285 & ~w16285) | (pi285 & w19907) | (~w16285 & w19907);
assign w16287 = w13180 & w13296;
assign w16288 = ~w13226 & ~w16287;
assign w16289 = w13194 & w13679;
assign w16290 = ~w13221 & ~w13757;
assign w16291 = w13679 & w19908;
assign w16292 = w16290 & ~w16291;
assign w16293 = ~pi285 & ~w16288;
assign w16294 = w16292 & ~w16293;
assign w16295 = ~w13703 & w19909;
assign w16296 = ~pi231 & ~w16295;
assign w16297 = (w13294 & w13277) | (w13294 & w19910) | (w13277 & w19910);
assign w16298 = ~pi215 & ~w13248;
assign w16299 = w13687 & w16298;
assign w16300 = ~w15453 & ~w16299;
assign w16301 = ~w15419 & ~w16297;
assign w16302 = w16300 & w16301;
assign w16303 = ~w16296 & w16302;
assign w16304 = ~w13230 & ~w14961;
assign w16305 = w13265 & ~w16304;
assign w16306 = ~w13298 & ~w16305;
assign w16307 = (w16306 & w16303) | (w16306 & w19911) | (w16303 & w19911);
assign w16308 = ~pi234 & ~w16294;
assign w16309 = w16307 & ~w16308;
assign w16310 = ~w16267 & w16309;
assign w16311 = w16310 & w19912;
assign w16312 = (~w16249 & ~w16310) | (~w16249 & w19913) | (~w16310 & w19913);
assign w16313 = pi532 & pi583;
assign w16314 = ~w16311 & ~w16312;
assign w16315 = ~pi532 & w16314;
assign w16316 = ~w16313 & ~w16315;
assign w16317 = ~w14377 & w15903;
assign w16318 = ~w15549 & ~w16317;
assign w16319 = ~w14295 & ~w14637;
assign w16320 = ~pi138 & ~w16319;
assign w16321 = ~w14453 & ~w14624;
assign w16322 = ~w14327 & ~w16320;
assign w16323 = w16322 & w19914;
assign w16324 = ~pi302 & ~w16323;
assign w16325 = ~pi185 & pi207;
assign w16326 = w14233 & w16325;
assign w16327 = (pi302 & w14653) | (pi302 & w19915) | (w14653 & w19915);
assign w16328 = ~w14268 & ~w14316;
assign w16329 = (w14210 & ~w16328) | (w14210 & w16729) | (~w16328 & w16729);
assign w16330 = ~pi138 & w14624;
assign w16331 = pi147 & w14193;
assign w16332 = ~w14438 & ~w16331;
assign w16333 = w14304 & ~w16332;
assign w16334 = ~w14648 & ~w15886;
assign w16335 = ~w16330 & w16334;
assign w16336 = w16335 & w19916;
assign w16337 = ~w16329 & w16336;
assign w16338 = ~w16324 & w16337;
assign w16339 = ~w14290 & ~w15511;
assign w16340 = pi207 & w16339;
assign w16341 = pi147 & w14270;
assign w16342 = ~w14241 & ~w16341;
assign w16343 = w14615 & w16342;
assign w16344 = ~w16340 & ~w16343;
assign w16345 = (pi302 & w16344) | (pi302 & w19917) | (w16344 & w19917);
assign w16346 = pi207 & ~w15874;
assign w16347 = ~w14339 & ~w16346;
assign w16348 = w14284 & w14329;
assign w16349 = ~w14386 & ~w16348;
assign w16350 = (~w14257 & w16349) | (~w14257 & w19918) | (w16349 & w19918);
assign w16351 = ~w16347 & w16350;
assign w16352 = ~w16345 & w16351;
assign w16353 = ~pi139 & ~w16352;
assign w16354 = ~w15517 & w19919;
assign w16355 = ~pi207 & ~w16354;
assign w16356 = (w14210 & w14427) | (w14210 & w19920) | (w14427 & w19920);
assign w16357 = ~w14193 & w14205;
assign w16358 = ~w14240 & w16357;
assign w16359 = ~w15501 & ~w16358;
assign w16360 = w14232 & w14239;
assign w16361 = w16359 & w19921;
assign w16362 = ~w16355 & w16361;
assign w16363 = ~pi302 & ~w16362;
assign w16364 = ~w14413 & w19922;
assign w16365 = ~pi207 & ~w16364;
assign w16366 = w14210 & w14630;
assign w16367 = (pi302 & w16365) | (pi302 & w19923) | (w16365 & w19923);
assign w16368 = ~w14294 & ~w14324;
assign w16369 = pi302 & ~w16368;
assign w16370 = ~w14390 & ~w15886;
assign w16371 = ~w16369 & w16370;
assign w16372 = ~w16363 & ~w16367;
assign w16373 = (~w14442 & w16371) | (~w14442 & w19924) | (w16371 & w19924);
assign w16374 = w16372 & w16373;
assign w16375 = ~w16353 & w16374;
assign w16376 = ~pi218 & pi349;
assign w16377 = pi218 & ~pi349;
assign w16378 = ~w16376 & ~w16377;
assign w16379 = ~pi350 & ~w16378;
assign w16380 = pi350 & w16378;
assign w16381 = ~w16379 & ~w16380;
assign w16382 = w16375 & w19925;
assign w16383 = (~w16381 & ~w16375) | (~w16381 & w19926) | (~w16375 & w19926);
assign w16384 = pi532 & pi567;
assign w16385 = ~w16382 & ~w16383;
assign w16386 = ~pi532 & w16385;
assign w16387 = ~w16384 & ~w16386;
assign w16388 = ~w13195 & ~w13199;
assign w16389 = ~pi231 & ~w16388;
assign w16390 = ~w14972 & ~w16389;
assign w16391 = ~w13317 & ~w13664;
assign w16392 = ~w13256 & ~w14903;
assign w16393 = (~pi231 & w13703) | (~pi231 & w19927) | (w13703 & w19927);
assign w16394 = ~w13254 & ~w13725;
assign w16395 = pi231 & ~w16394;
assign w16396 = w13190 & ~w13281;
assign w16397 = w14894 & w16396;
assign w16398 = ~w15657 & ~w16397;
assign w16399 = ~pi234 & w16398;
assign w16400 = ~w16395 & w16399;
assign w16401 = (~pi285 & ~w16391) | (~pi285 & w19928) | (~w16391 & w19928);
assign w16402 = w16400 & w20910;
assign w16403 = (pi285 & ~w16390) | (pi285 & w19929) | (~w16390 & w19929);
assign w16404 = w16402 & ~w16403;
assign w16405 = pi231 & ~w13230;
assign w16406 = ~w13714 & ~w16405;
assign w16407 = w13210 & ~w15594;
assign w16408 = ~pi285 & ~w13755;
assign w16409 = ~w16407 & w16408;
assign w16410 = ~w16406 & w16409;
assign w16411 = ~w13679 & w15624;
assign w16412 = ~pi231 & w16411;
assign w16413 = w16410 & ~w16412;
assign w16414 = ~w13282 & ~w13290;
assign w16415 = ~w13730 & ~w14889;
assign w16416 = w16414 & w16415;
assign w16417 = pi231 & ~w16416;
assign w16418 = (pi285 & ~w13679) | (pi285 & w19930) | (~w13679 & w19930);
assign w16419 = ~w14893 & w16418;
assign w16420 = ~w16417 & w16419;
assign w16421 = ~w16413 & ~w16420;
assign w16422 = w13197 & w13295;
assign w16423 = ~w14908 & ~w16422;
assign w16424 = w13190 & w14962;
assign w16425 = w16423 & ~w16424;
assign w16426 = ~w13220 & ~w14923;
assign w16427 = w13265 & ~w16426;
assign w16428 = (pi234 & ~w13186) | (pi234 & w19931) | (~w13186 & w19931);
assign w16429 = ~w16427 & w16428;
assign w16430 = w16425 & w16429;
assign w16431 = ~w16421 & w16430;
assign w16432 = ~w14923 & ~w14961;
assign w16433 = w16432 & w19932;
assign w16434 = ~w13695 & ~w13721;
assign w16435 = (w16434 & w16433) | (w16434 & w19933) | (w16433 & w19933);
assign w16436 = w13213 & ~w13255;
assign w16437 = (pi175 & ~w14932) | (pi175 & w19934) | (~w14932 & w19934);
assign w16438 = (pi285 & w16437) | (pi285 & w19935) | (w16437 & w19935);
assign w16439 = ~w16435 & w16438;
assign w16440 = ~w13226 & ~w16397;
assign w16441 = (~pi285 & ~w16440) | (~pi285 & w19936) | (~w16440 & w19936);
assign w16442 = w13198 & w13290;
assign w16443 = ~w13678 & ~w16442;
assign w16444 = ~w16289 & w19937;
assign w16445 = w13303 & ~w16444;
assign w16446 = ~pi231 & ~w16443;
assign w16447 = ~w16445 & ~w16446;
assign w16448 = ~w16441 & w16447;
assign w16449 = ~w16439 & w16448;
assign w16450 = (w19938 & w20911) | (w19938 & w20912) | (w20911 & w20912);
assign w16451 = (~w19938 & w20913) | (~w19938 & w20914) | (w20913 & w20914);
assign w16452 = ~w16450 & ~w16451;
assign w16453 = ~pi219 & pi375;
assign w16454 = pi219 & ~pi375;
assign w16455 = ~w16453 & ~w16454;
assign w16456 = ~w16452 & w16455;
assign w16457 = w16452 & ~w16455;
assign w16458 = ~w16456 & ~w16457;
assign w16459 = pi532 & ~pi588;
assign w16460 = ~pi532 & ~w16458;
assign w16461 = ~w16459 & ~w16460;
assign w16462 = ~w13277 & ~w14907;
assign w16463 = w14968 & w16462;
assign w16464 = ~w14973 & w15427;
assign w16465 = ~w13731 & w16464;
assign w16466 = ~w16463 & ~w16465;
assign w16467 = w13225 & w13303;
assign w16468 = (~pi215 & w16467) | (~pi215 & w19939) | (w16467 & w19939);
assign w16469 = pi234 & ~w16468;
assign w16470 = ~w16466 & w16469;
assign w16471 = ~w13716 & ~w14902;
assign w16472 = ~pi231 & ~w16471;
assign w16473 = w13183 & ~w13740;
assign w16474 = ~w16472 & ~w16473;
assign w16475 = ~w13265 & ~w13664;
assign w16476 = ~w13717 & ~w16475;
assign w16477 = w13190 & w15601;
assign w16478 = w15601 & w19940;
assign w16479 = ~w16262 & ~w16478;
assign w16480 = ~w16476 & w16479;
assign w16481 = ~pi234 & w16480;
assign w16482 = w13201 & w13236;
assign w16483 = ~w15461 & ~w16482;
assign w16484 = ~w13664 & w16483;
assign w16485 = w13186 & w13190;
assign w16486 = w16484 & ~w16485;
assign w16487 = ~w16466 & w19941;
assign w16488 = w16481 & w16486;
assign w16489 = ~w16487 & ~w16488;
assign w16490 = ~w13297 & ~w14942;
assign w16491 = ~pi175 & ~w16490;
assign w16492 = ~w13721 & ~w13755;
assign w16493 = ~w13196 & w16492;
assign w16494 = ~w16491 & w16493;
assign w16495 = ~w13703 & ~w15635;
assign w16496 = ~w16477 & w16495;
assign w16497 = w13193 & ~w16262;
assign w16498 = w16496 & w16497;
assign w16499 = pi231 & ~w16494;
assign w16500 = w16498 & ~w16499;
assign w16501 = ~w13306 & ~w13756;
assign w16502 = w13237 & w15594;
assign w16503 = w16501 & ~w16502;
assign w16504 = w13212 & ~w13292;
assign w16505 = w16503 & ~w16504;
assign w16506 = ~w13221 & ~w13297;
assign w16507 = ~w15595 & w16506;
assign w16508 = ~pi231 & ~w16507;
assign w16509 = w13214 & w13265;
assign w16510 = ~w16509 & w19942;
assign w16511 = ~w16508 & w16510;
assign w16512 = w16470 & w16505;
assign w16513 = w16481 & w16511;
assign w16514 = w13296 & w14913;
assign w16515 = ~w14916 & w16418;
assign w16516 = ~w13205 & w16274;
assign w16517 = w16515 & ~w16516;
assign w16518 = ~w14971 & ~w15434;
assign w16519 = ~w16514 & w16518;
assign w16520 = w16517 & w16519;
assign w16521 = ~w16489 & w16500;
assign w16522 = (w16520 & w16512) | (w16520 & w19943) | (w16512 & w19943);
assign w16523 = ~w16521 & ~w16522;
assign w16524 = ~pi231 & w13736;
assign w16525 = (pi175 & w16524) | (pi175 & w19944) | (w16524 & w19944);
assign w16526 = ~pi220 & pi356;
assign w16527 = pi220 & ~pi356;
assign w16528 = ~w16526 & ~w16527;
assign w16529 = ~pi357 & ~w16528;
assign w16530 = pi357 & w16528;
assign w16531 = ~w16529 & ~w16530;
assign w16532 = ~w16523 & w19945;
assign w16533 = (~w16531 & w16523) | (~w16531 & w19946) | (w16523 & w19946);
assign w16534 = pi532 & pi585;
assign w16535 = ~w16532 & ~w16533;
assign w16536 = ~pi532 & w16535;
assign w16537 = ~w16534 & ~w16536;
assign w16538 = ~pi221 & pi255;
assign w16539 = pi221 & ~pi255;
assign w16540 = ~w16538 & ~w16539;
assign w16541 = ~pi384 & ~w16540;
assign w16542 = pi384 & w16540;
assign w16543 = ~w16541 & ~w16542;
assign w16544 = ~w16015 & w16543;
assign w16545 = w16015 & ~w16543;
assign w16546 = pi532 & pi593;
assign w16547 = ~w16544 & ~w16545;
assign w16548 = ~pi532 & w16547;
assign w16549 = ~w16546 & ~w16548;
assign w16550 = w14779 & w19947;
assign w16551 = (pi222 & ~w14779) | (pi222 & w19948) | (~w14779 & w19948);
assign w16552 = ~w16550 & ~w16551;
assign w16553 = pi532 & ~pi639;
assign w16554 = ~pi532 & ~w16552;
assign w16555 = ~w16553 & ~w16554;
assign w16556 = ~pi223 & w15834;
assign w16557 = pi223 & ~w15834;
assign w16558 = ~w16556 & ~w16557;
assign w16559 = pi532 & ~pi642;
assign w16560 = ~pi532 & ~w16558;
assign w16561 = ~w16559 & ~w16560;
assign w16562 = ~pi224 & w15157;
assign w16563 = pi224 & ~w15157;
assign w16564 = ~w16562 & ~w16563;
assign w16565 = pi532 & ~pi644;
assign w16566 = ~pi532 & ~w16564;
assign w16567 = ~w16565 & ~w16566;
assign w16568 = ~w15065 & w19949;
assign w16569 = (pi225 & w15065) | (pi225 & w19950) | (w15065 & w19950);
assign w16570 = ~w16568 & ~w16569;
assign w16571 = pi532 & ~pi637;
assign w16572 = ~pi532 & ~w16570;
assign w16573 = ~w16571 & ~w16572;
assign w16574 = pi226 & ~w16558;
assign w16575 = ~pi226 & w16558;
assign w16576 = pi532 & pi610;
assign w16577 = ~w16574 & ~w16575;
assign w16578 = ~pi532 & w16577;
assign w16579 = ~w16576 & ~w16578;
assign w16580 = pi227 & w14863;
assign w16581 = ~pi227 & ~w14863;
assign w16582 = pi532 & pi611;
assign w16583 = ~w16580 & ~w16581;
assign w16584 = ~pi532 & w16583;
assign w16585 = ~w16582 & ~w16584;
assign w16586 = ~pi228 & ~w16564;
assign w16587 = pi228 & w16564;
assign w16588 = pi532 & pi612;
assign w16589 = ~w16586 & ~w16587;
assign w16590 = ~pi532 & w16589;
assign w16591 = ~w16588 & ~w16590;
assign w16592 = ~pi229 & ~w16552;
assign w16593 = pi229 & w16552;
assign w16594 = pi532 & pi607;
assign w16595 = ~w16592 & ~w16593;
assign w16596 = ~pi532 & w16595;
assign w16597 = ~w16594 & ~w16596;
assign w16598 = ~pi230 & ~w16570;
assign w16599 = pi230 & w16570;
assign w16600 = pi532 & pi605;
assign w16601 = ~w16598 & ~w16599;
assign w16602 = ~pi532 & w16601;
assign w16603 = ~w16600 & ~w16602;
assign w16604 = ~pi231 & w14687;
assign w16605 = pi231 & ~w14687;
assign w16606 = ~w16604 & ~w16605;
assign w16607 = w14779 & w19951;
assign w16608 = (w16606 & ~w14779) | (w16606 & w19952) | (~w14779 & w19952);
assign w16609 = pi532 & pi543;
assign w16610 = ~w16607 & ~w16608;
assign w16611 = ~pi532 & w16610;
assign w16612 = ~w16609 & ~w16611;
assign w16613 = ~pi226 & pi232;
assign w16614 = pi226 & ~pi232;
assign w16615 = ~w16613 & ~w16614;
assign w16616 = w15767 & w16615;
assign w16617 = ~w15767 & ~w16615;
assign w16618 = ~w16616 & ~w16617;
assign w16619 = ~w15834 & ~w16618;
assign w16620 = w15834 & w16618;
assign w16621 = pi532 & pi546;
assign w16622 = ~w16619 & ~w16620;
assign w16623 = ~pi532 & w16622;
assign w16624 = ~w16621 & ~w16623;
assign w16625 = ~pi233 & w15079;
assign w16626 = pi233 & ~w15079;
assign w16627 = ~w16625 & ~w16626;
assign w16628 = w15157 & ~w16627;
assign w16629 = ~w15157 & w16627;
assign w16630 = pi532 & pi548;
assign w16631 = ~w16628 & ~w16629;
assign w16632 = ~pi532 & w16631;
assign w16633 = ~w16630 & ~w16632;
assign w16634 = ~pi234 & w14992;
assign w16635 = pi234 & ~w14992;
assign w16636 = ~w16634 & ~w16635;
assign w16637 = ~w15065 & w19953;
assign w16638 = (w16636 & w15065) | (w16636 & w19954) | (w15065 & w19954);
assign w16639 = pi532 & pi541;
assign w16640 = ~w16637 & ~w16638;
assign w16641 = ~pi532 & w16640;
assign w16642 = ~w16639 & ~w16641;
assign w16643 = w11418 & w19955;
assign w16644 = (pi129 & ~w11418) | (pi129 & w19956) | (~w11418 & w19956);
assign w16645 = ~w16643 & ~w16644;
assign w16646 = w5071 & w19957;
assign w16647 = (pi121 & ~w5071) | (pi121 & w19958) | (~w5071 & w19958);
assign w16648 = ~w16646 & ~w16647;
assign w16649 = ~w8073 & w19959;
assign w16650 = (pi179 & w8073) | (pi179 & w19960) | (w8073 & w19960);
assign w16651 = ~w16649 & ~w16650;
assign w16652 = w3101 & w19961;
assign w16653 = (pi280 & ~w3101) | (pi280 & w19962) | (~w3101 & w19962);
assign w16654 = ~w16652 & ~w16653;
assign w16655 = w6622 & w19963;
assign w16656 = (pi225 & ~w6622) | (pi225 & w19964) | (~w6622 & w19964);
assign w16657 = ~w16655 & ~w16656;
assign w16658 = ~w9372 & w19965;
assign w16659 = (pi226 & w9372) | (pi226 & w19966) | (w9372 & w19966);
assign w16660 = ~w16658 & ~w16659;
assign w16661 = ~pi232 & w10775;
assign w16662 = pi232 & ~w10775;
assign w16663 = ~w16661 & ~w16662;
assign w16664 = w6173 & w19967;
assign w16665 = (pi130 & ~w6173) | (pi130 & w19968) | (~w6173 & w19968);
assign w16666 = ~w16664 & ~w16665;
assign w16667 = w3769 & w19969;
assign w16668 = (pi132 & ~w3769) | (pi132 & w19970) | (~w3769 & w19970);
assign w16669 = ~w16667 & ~w16668;
assign w16670 = w143 & w19971;
assign w16671 = (pi156 & ~w143) | (pi156 & w19972) | (~w143 & w19972);
assign w16672 = ~w16670 & ~w16671;
assign w16673 = w5328 & w19973;
assign w16674 = (pi151 & ~w5328) | (pi151 & w19974) | (~w5328 & w19974);
assign w16675 = ~w16673 & ~w16674;
assign w16676 = ~w8431 & w19975;
assign w16677 = (pi228 & w8431) | (pi228 & w19976) | (w8431 & w19976);
assign w16678 = ~w16676 & ~w16677;
assign w16679 = ~pi229 & w9551;
assign w16680 = pi229 & ~w9551;
assign w16681 = ~w16679 & ~w16680;
assign w16682 = ~pi319 & w6869;
assign w16683 = pi319 & ~w6869;
assign w16684 = ~w16682 & ~w16683;
assign w16685 = ~pi153 & w11527;
assign w16686 = pi153 & ~w11527;
assign w16687 = ~w16685 & ~w16686;
assign w16688 = ~pi146 & w11884;
assign w16689 = pi146 & ~w11884;
assign w16690 = ~w16688 & ~w16689;
assign w16691 = ~pi256 & w10526;
assign w16692 = pi256 & ~w10526;
assign w16693 = ~w16691 & ~w16692;
assign w16694 = ~pi227 & w11750;
assign w16695 = pi227 & ~w11750;
assign w16696 = ~w16694 & ~w16695;
assign w16697 = ~pi303 & w9891;
assign w16698 = pi303 & ~w9891;
assign w16699 = ~w16697 & ~w16698;
assign w16700 = ~pi255 & w10014;
assign w16701 = pi255 & ~w10014;
assign w16702 = ~w16700 & ~w16701;
assign w16703 = ~pi384 & w16012;
assign w16704 = pi384 & ~w16012;
assign w16705 = ~w16703 & ~w16704;
assign w16706 = pi255 & ~w16705;
assign w16707 = ~pi255 & w16705;
assign w16708 = pi532 & pi657;
assign w16709 = ~w16706 & ~w16707;
assign w16710 = ~pi532 & w16709;
assign w16711 = ~w16708 & ~w16710;
assign w16712 = pi532 & pi643;
assign w16713 = ~pi532 & w14863;
assign w16714 = ~w16712 & ~w16713;
assign w16715 = (~w14226 & ~w16332) | (~w14226 & w19977) | (~w16332 & w19977);
assign w16716 = (pi207 & w14231) | (pi207 & w19978) | (w14231 & w19978);
assign w16717 = ~w14207 & w14291;
assign w16718 = ~w16716 & w16717;
assign w16719 = ~pi207 & ~w16715;
assign w16720 = w16718 & ~w16719;
assign w16721 = w14292 & w19639;
assign w16722 = ~w14427 & ~w16721;
assign w16723 = ~w14232 & w14316;
assign w16724 = w14251 & w14590;
assign w16725 = ~w16723 & ~w16724;
assign w16726 = ~w16330 & w16725;
assign w16727 = (~pi302 & ~w16726) | (~pi302 & w19979) | (~w16726 & w19979);
assign w16728 = ~w14328 & ~w15885;
assign w16729 = w14210 & w14405;
assign w16730 = w16728 & ~w16729;
assign w16731 = (w14232 & w14234) | (w14232 & w19980) | (w14234 & w19980);
assign w16732 = ~w14398 & ~w16731;
assign w16733 = w16730 & w16732;
assign w16734 = ~w16727 & w16733;
assign w16735 = pi302 & ~w16720;
assign w16736 = w16734 & ~w16735;
assign w16737 = ~w14391 & ~w15887;
assign w16738 = (pi207 & ~w16737) | (pi207 & w19981) | (~w16737 & w19981);
assign w16739 = w14209 & w14284;
assign w16740 = w14190 & w14194;
assign w16741 = w14197 & ~w16325;
assign w16742 = pi166 & w16740;
assign w16743 = ~w16741 & ~w16742;
assign w16744 = ~w14630 & ~w16739;
assign w16745 = ~pi302 & w16744;
assign w16746 = w16743 & w16745;
assign w16747 = ~w14413 & w19982;
assign w16748 = ~w16738 & w16747;
assign w16749 = ~w16746 & ~w16748;
assign w16750 = ~w14637 & ~w15525;
assign w16751 = w14193 & ~w16750;
assign w16752 = ~w14405 & ~w15512;
assign w16753 = ~w14620 & w16752;
assign w16754 = pi207 & ~w14204;
assign w16755 = (~w16754 & ~w16753) | (~w16754 & w19983) | (~w16753 & w19983);
assign w16756 = ~w16751 & ~w16755;
assign w16757 = ~w16749 & w16756;
assign w16758 = pi139 & ~w16757;
assign w16759 = ~w14190 & ~w14209;
assign w16760 = w15525 & w16759;
assign w16761 = ~w14207 & ~w16740;
assign w16762 = ~pi207 & ~w16761;
assign w16763 = w14240 & w14601;
assign w16764 = (pi302 & ~w14637) | (pi302 & w19785) | (~w14637 & w19785);
assign w16765 = ~w16762 & ~w16763;
assign w16766 = (pi207 & w16760) | (pi207 & w19984) | (w16760 & w19984);
assign w16767 = w16765 & w20915;
assign w16768 = ~w14364 & ~w14606;
assign w16769 = ~w14279 & w16768;
assign w16770 = ~pi207 & ~w16769;
assign w16771 = ~w14285 & w14373;
assign w16772 = ~w16770 & w16771;
assign w16773 = ~w14243 & ~w14317;
assign w16774 = ~pi138 & w14448;
assign w16775 = (w16774 & ~w16773) | (w16774 & w19985) | (~w16773 & w19985);
assign w16776 = w14249 & w16326;
assign w16777 = ~w14455 & ~w16776;
assign w16778 = ~w16775 & w16777;
assign w16779 = (w16778 & w16767) | (w16778 & w19986) | (w16767 & w19986);
assign w16780 = ~w16758 & w16779;
assign w16781 = ~pi139 & ~w16736;
assign w16782 = w16780 & ~w16781;
assign w16783 = ~pi376 & w16782;
assign w16784 = pi376 & ~w16782;
assign w16785 = ~w16783 & ~w16784;
assign w16786 = ~pi257 & pi373;
assign w16787 = pi257 & ~pi373;
assign w16788 = ~w16786 & ~w16787;
assign w16789 = ~w16785 & w16788;
assign w16790 = w16785 & ~w16788;
assign w16791 = ~w16789 & ~w16790;
assign w16792 = pi532 & ~pi566;
assign w16793 = ~pi532 & ~w16791;
assign w16794 = ~w16792 & ~w16793;
assign w16795 = ~w14200 & w14213;
assign w16796 = ~w14438 & ~w16795;
assign w16797 = pi207 & ~w14390;
assign w16798 = w15531 & w16796;
assign w16799 = ~w16797 & ~w16798;
assign w16800 = w14377 & ~w16325;
assign w16801 = (~pi302 & w16799) | (~pi302 & w19987) | (w16799 & w19987);
assign w16802 = ~w14251 & ~w14438;
assign w16803 = w15881 & w16802;
assign w16804 = pi207 & ~w16803;
assign w16805 = ~w14591 & ~w15874;
assign w16806 = (pi302 & w16804) | (pi302 & w19988) | (w16804 & w19988);
assign w16807 = ~pi185 & w14292;
assign w16808 = ~w14195 & ~w16807;
assign w16809 = w14232 & ~w16808;
assign w16810 = w14436 & w15875;
assign w16811 = ~w14451 & ~w16810;
assign w16812 = ~w14216 & ~w14612;
assign w16813 = ~w16809 & w16811;
assign w16814 = ~w16801 & ~w16806;
assign w16815 = w14210 & w14305;
assign w16816 = ~w15925 & ~w16815;
assign w16817 = ~w14325 & ~w14606;
assign w16818 = ~pi302 & w16817;
assign w16819 = w16816 & w16818;
assign w16820 = ~w14283 & ~w14364;
assign w16821 = ~pi207 & ~w16820;
assign w16822 = ~w14661 & ~w15526;
assign w16823 = pi302 & ~w15512;
assign w16824 = w16822 & w16823;
assign w16825 = ~w16821 & w16824;
assign w16826 = ~w16819 & ~w16825;
assign w16827 = ~pi207 & ~w14278;
assign w16828 = ~w15517 & w16827;
assign w16829 = w14336 & ~w14413;
assign w16830 = ~w14214 & w14436;
assign w16831 = w14592 & w16830;
assign w16832 = ~w16776 & ~w16831;
assign w16833 = (w16832 & w16829) | (w16832 & w19990) | (w16829 & w19990);
assign w16834 = w14194 & ~w14200;
assign w16835 = (pi138 & ~w14631) | (pi138 & w19991) | (~w14631 & w19991);
assign w16836 = ~pi207 & ~w16835;
assign w16837 = ~w14337 & ~w16807;
assign w16838 = (~pi138 & ~w16837) | (~pi138 & w19992) | (~w16837 & w19992);
assign w16839 = ~w14253 & ~w14289;
assign w16840 = pi207 & w16839;
assign w16841 = ~w16838 & w16840;
assign w16842 = w14249 & w14325;
assign w16843 = ~w16831 & ~w16842;
assign w16844 = w16843 & w19993;
assign w16845 = (w14448 & w15874) | (w14448 & w19994) | (w15874 & w19994);
assign w16846 = ~pi129 & w14264;
assign w16847 = ~w14218 & ~w16846;
assign w16848 = ~pi207 & ~w16847;
assign w16849 = ~w16845 & ~w16848;
assign w16850 = ~pi302 & ~w16844;
assign w16851 = w16849 & ~w16850;
assign w16852 = ~w16836 & ~w16841;
assign w16853 = pi302 & w16852;
assign w16854 = w16851 & ~w16853;
assign w16855 = (~pi139 & w16826) | (~pi139 & w19995) | (w16826 & w19995);
assign w16856 = w16854 & ~w16855;
assign w16857 = w16856 & w19996;
assign w16858 = (pi370 & ~w16856) | (pi370 & w19997) | (~w16856 & w19997);
assign w16859 = ~w16857 & ~w16858;
assign w16860 = ~pi258 & pi348;
assign w16861 = pi258 & ~pi348;
assign w16862 = ~w16860 & ~w16861;
assign w16863 = ~w16859 & w16862;
assign w16864 = w16859 & ~w16862;
assign w16865 = ~w16863 & ~w16864;
assign w16866 = pi532 & ~pi572;
assign w16867 = ~pi532 & ~w16865;
assign w16868 = ~w16866 & ~w16867;
assign w16869 = ~pi157 & w11133;
assign w16870 = pi157 & ~w11133;
assign w16871 = ~w16869 & ~w16870;
assign w16872 = ~pi160 & w2849;
assign w16873 = pi160 & ~w2849;
assign w16874 = ~w16872 & ~w16873;
assign w16875 = w4984 & w19998;
assign w16876 = (pi193 & ~w4984) | (pi193 & w19999) | (~w4984 & w19999);
assign w16877 = ~w16875 & ~w16876;
assign w16878 = ~pi170 & w10983;
assign w16879 = pi170 & ~w10983;
assign w16880 = ~w16878 & ~w16879;
assign w16881 = w7655 & w20000;
assign w16882 = (pi142 & ~w7655) | (pi142 & w20001) | (~w7655 & w20001);
assign w16883 = ~w16881 & ~w16882;
assign w16884 = w807 & w20002;
assign w16885 = (pi143 & ~w807) | (pi143 & w20003) | (~w807 & w20003);
assign w16886 = ~w16884 & ~w16885;
assign w16887 = ~pi178 & w9783;
assign w16888 = pi178 & ~w9783;
assign w16889 = ~w16887 & ~w16888;
assign w16890 = ~pi180 & w8809;
assign w16891 = pi180 & ~w8809;
assign w16892 = ~w16890 & ~w16891;
assign w16893 = ~pi267 & pi303;
assign w16894 = pi267 & ~pi303;
assign w16895 = ~w16893 & ~w16894;
assign w16896 = ~pi389 & ~w16895;
assign w16897 = pi389 & w16895;
assign w16898 = ~w16896 & ~w16897;
assign w16899 = (~w16169 & ~w16139) | (~w16169 & w20004) | (~w16139 & w20004);
assign w16900 = (pi351 & w13781) | (pi351 & w20005) | (w13781 & w20005);
assign w16901 = w13499 & ~w13581;
assign w16902 = ~w16900 & w16901;
assign w16903 = ~pi351 & ~w16899;
assign w16904 = w16902 & ~w16903;
assign w16905 = pi284 & ~w16904;
assign w16906 = (~pi351 & w14476) | (~pi351 & w20006) | (w14476 & w20006);
assign w16907 = ~w13854 & ~w15953;
assign w16908 = w16907 & w20007;
assign w16909 = (~pi284 & ~w16908) | (~pi284 & w20008) | (~w16908 & w20008);
assign w16910 = ~pi132 & w13591;
assign w16911 = ~w15954 & ~w16910;
assign w16912 = ~w13837 & w16911;
assign w16913 = ~w13543 & w15282;
assign w16914 = w16912 & w16913;
assign w16915 = ~w16905 & w20009;
assign w16916 = ~pi193 & ~w16915;
assign w16917 = pi157 & w14496;
assign w16918 = ~w13485 & ~w14080;
assign w16919 = ~w16917 & w16918;
assign w16920 = ~pi284 & w16919;
assign w16921 = (w13482 & w16130) | (w13482 & w20010) | (w16130 & w20010);
assign w16922 = w16920 & ~w16921;
assign w16923 = ~w13777 & ~w14107;
assign w16924 = (pi351 & ~w16923) | (pi351 & w20011) | (~w16923 & w20011);
assign w16925 = w16168 & ~w16924;
assign w16926 = pi284 & w16925;
assign w16927 = ~w16922 & ~w16926;
assign w16928 = ~w13515 & ~w13539;
assign w16929 = w13550 & ~w16928;
assign w16930 = ~w13787 & ~w14117;
assign w16931 = ~w14517 & w16009;
assign w16932 = (~w16172 & ~w16931) | (~w16172 & w20012) | (~w16931 & w20012);
assign w16933 = (pi193 & w16927) | (pi193 & w20013) | (w16927 & w20013);
assign w16934 = ~w14105 & ~w15307;
assign w16935 = (~pi351 & ~w16934) | (~pi351 & w20014) | (~w16934 & w20014);
assign w16936 = ~w13486 & ~w13818;
assign w16937 = (~pi284 & w16935) | (~pi284 & w20015) | (w16935 & w20015);
assign w16938 = (w14528 & ~w14494) | (w14528 & w20016) | (~w14494 & w20016);
assign w16939 = ~w16917 & w20017;
assign w16940 = w13510 & ~w14100;
assign w16941 = w16939 & ~w16940;
assign w16942 = ~w13566 & ~w14133;
assign w16943 = ~w13473 & w16942;
assign w16944 = w13850 & ~w16943;
assign w16945 = ~w13858 & ~w15326;
assign w16946 = ~w16944 & w16945;
assign w16947 = w13508 & ~w16941;
assign w16948 = w16946 & ~w16947;
assign w16949 = w16948 & w20018;
assign w16950 = ~w16933 & w16949;
assign w16951 = ~w16916 & w16950;
assign w16952 = ~pi268 & w16951;
assign w16953 = pi268 & ~w16951;
assign w16954 = ~w16952 & ~w16953;
assign w16955 = ~w16898 & ~w16954;
assign w16956 = w16898 & w16954;
assign w16957 = pi532 & pi590;
assign w16958 = ~w16955 & ~w16956;
assign w16959 = ~pi532 & w16958;
assign w16960 = ~w16957 & ~w16959;
assign w16961 = ~pi268 & pi303;
assign w16962 = pi268 & ~pi303;
assign w16963 = ~w16961 & ~w16962;
assign w16964 = ~pi389 & w16951;
assign w16965 = pi389 & ~w16951;
assign w16966 = ~w16964 & ~w16965;
assign w16967 = ~w16963 & ~w16966;
assign w16968 = w16963 & w16966;
assign w16969 = pi532 & pi622;
assign w16970 = ~w16967 & ~w16968;
assign w16971 = ~pi532 & w16970;
assign w16972 = ~w16969 & ~w16971;
assign w16973 = ~w15254 & w20019;
assign w16974 = (pi269 & w15254) | (pi269 & w20020) | (w15254 & w20020);
assign w16975 = ~w16973 & ~w16974;
assign w16976 = pi532 & ~pi641;
assign w16977 = ~pi532 & ~w16975;
assign w16978 = ~w16976 & ~w16977;
assign w16979 = ~pi270 & ~w15181;
assign w16980 = pi270 & w15181;
assign w16981 = ~w16979 & ~w16980;
assign w16982 = w15257 & ~w16981;
assign w16983 = ~w15257 & w16981;
assign w16984 = pi532 & pi545;
assign w16985 = ~w16982 & ~w16983;
assign w16986 = ~pi532 & w16985;
assign w16987 = ~w16984 & ~w16986;
assign w16988 = w15480 & w20021;
assign w16989 = (pi271 & ~w15480) | (pi271 & w20022) | (~w15480 & w20022);
assign w16990 = ~w16988 & ~w16989;
assign w16991 = pi532 & ~pi651;
assign w16992 = ~pi532 & ~w16990;
assign w16993 = ~w16991 & ~w16992;
assign w16994 = ~pi272 & w15556;
assign w16995 = pi272 & ~w15556;
assign w16996 = ~w16994 & ~w16995;
assign w16997 = pi532 & ~pi635;
assign w16998 = ~pi532 & ~w16996;
assign w16999 = ~w16997 & ~w16998;
assign w17000 = ~pi273 & ~w16990;
assign w17001 = pi273 & w16990;
assign w17002 = pi532 & pi619;
assign w17003 = ~w17000 & ~w17001;
assign w17004 = ~pi532 & w17003;
assign w17005 = ~w17002 & ~w17004;
assign w17006 = ~pi274 & ~w16996;
assign w17007 = pi274 & w16996;
assign w17008 = pi532 & pi603;
assign w17009 = ~w17006 & ~w17007;
assign w17010 = ~pi532 & w17009;
assign w17011 = ~w17008 & ~w17010;
assign w17012 = ~pi275 & w15417;
assign w17013 = pi275 & ~w15417;
assign w17014 = ~w17012 & ~w17013;
assign w17015 = w15480 & w20023;
assign w17016 = (w17014 & ~w15480) | (w17014 & w20024) | (~w15480 & w20024);
assign w17017 = pi532 & pi555;
assign w17018 = ~w17015 & ~w17016;
assign w17019 = ~pi532 & w17018;
assign w17020 = ~w17017 & ~w17019;
assign w17021 = ~pi276 & w15492;
assign w17022 = pi276 & ~w15492;
assign w17023 = ~w17021 & ~w17022;
assign w17024 = w15556 & ~w17023;
assign w17025 = ~w15556 & w17023;
assign w17026 = pi532 & pi539;
assign w17027 = ~w17024 & ~w17025;
assign w17028 = ~pi532 & w17027;
assign w17029 = ~w17026 & ~w17028;
assign w17030 = ~pi164 & w1206;
assign w17031 = pi164 & ~w1206;
assign w17032 = ~w17030 & ~w17031;
assign w17033 = ~w15641 & w20025;
assign w17034 = (pi278 & w15641) | (pi278 & w20026) | (w15641 & w20026);
assign w17035 = ~w17033 & ~w17034;
assign w17036 = pi532 & ~pi646;
assign w17037 = ~pi532 & ~w17035;
assign w17038 = ~w17036 & ~w17037;
assign w17039 = w1935 & w20027;
assign w17040 = (pi162 & ~w1935) | (pi162 & w20028) | (~w1935 & w20028);
assign w17041 = ~w17039 & ~w17040;
assign w17042 = ~pi280 & w15731;
assign w17043 = pi280 & ~w15731;
assign w17044 = ~w17042 & ~w17043;
assign w17045 = pi532 & ~pi638;
assign w17046 = ~pi532 & ~w17044;
assign w17047 = ~w17045 & ~w17046;
assign w17048 = ~pi281 & ~w17035;
assign w17049 = pi281 & w17035;
assign w17050 = pi532 & pi614;
assign w17051 = ~w17048 & ~w17049;
assign w17052 = ~pi532 & w17051;
assign w17053 = ~w17050 & ~w17052;
assign w17054 = ~pi133 & w7302;
assign w17055 = pi133 & ~w7302;
assign w17056 = ~w17054 & ~w17055;
assign w17057 = ~pi283 & ~w17044;
assign w17058 = pi283 & w17044;
assign w17059 = pi532 & pi606;
assign w17060 = ~w17057 & ~w17058;
assign w17061 = ~pi532 & w17060;
assign w17062 = ~w17059 & ~w17061;
assign w17063 = ~pi284 & w15592;
assign w17064 = pi284 & ~w15592;
assign w17065 = ~w17063 & ~w17064;
assign w17066 = ~w15641 & w20029;
assign w17067 = (w17065 & w15641) | (w17065 & w20030) | (w15641 & w20030);
assign w17068 = pi532 & pi550;
assign w17069 = ~w17066 & ~w17067;
assign w17070 = ~pi532 & w17069;
assign w17071 = ~w17068 & ~w17070;
assign w17072 = ~pi285 & w15737;
assign w17073 = pi285 & ~w15737;
assign w17074 = ~w17072 & ~w17073;
assign w17075 = w15731 & ~w17074;
assign w17076 = ~w15731 & w17074;
assign w17077 = pi532 & pi542;
assign w17078 = ~w17075 & ~w17076;
assign w17079 = ~pi532 & w17078;
assign w17080 = ~w17077 & ~w17079;
assign w17081 = w9234 & w20031;
assign w17082 = (pi149 & ~w9234) | (pi149 & w20032) | (~w9234 & w20032);
assign w17083 = ~w17081 & ~w17082;
assign w17084 = ~pi131 & w8992;
assign w17085 = pi131 & ~w8992;
assign w17086 = ~w17084 & ~w17085;
assign w17087 = ~pi139 & w4828;
assign w17088 = pi139 & ~w4828;
assign w17089 = ~w17087 & ~w17088;
assign w17090 = w8532 & w20033;
assign w17091 = (pi172 & ~w8532) | (pi172 & w20034) | (~w8532 & w20034);
assign w17092 = ~w17090 & ~w17091;
assign w17093 = w6003 & w20035;
assign w17094 = (pi134 & ~w6003) | (pi134 & w20036) | (~w6003 & w20036);
assign w17095 = ~w17093 & ~w17094;
assign w17096 = w2196 & w20037;
assign w17097 = (pi283 & ~w2196) | (pi283 & w20038) | (~w2196 & w20038);
assign w17098 = ~w17096 & ~w17097;
assign w17099 = ~pi222 & w6098;
assign w17100 = pi222 & ~w6098;
assign w17101 = ~w17099 & ~w17100;
assign w17102 = w12018 & w20039;
assign w17103 = (pi346 & ~w12018) | (pi346 & w20040) | (~w12018 & w20040);
assign w17104 = ~w17102 & ~w17103;
assign w17105 = ~pi147 & w10908;
assign w17106 = pi147 & ~w10908;
assign w17107 = ~w17105 & ~w17106;
assign w17108 = w3515 & w20041;
assign w17109 = (pi354 & ~w3515) | (pi354 & w20042) | (~w3515 & w20042);
assign w17110 = ~w17108 & ~w17109;
assign w17111 = ~pi351 & w4357;
assign w17112 = pi351 & ~w4357;
assign w17113 = ~w17111 & ~w17112;
assign w17114 = ~pi371 & w10600;
assign w17115 = pi371 & ~w10600;
assign w17116 = ~w17114 & ~w17115;
assign w17117 = w8149 & w20043;
assign w17118 = (pi267 & ~w8149) | (pi267 & w20044) | (~w8149 & w20044);
assign w17119 = ~w17117 & ~w17118;
assign w17120 = ~pi268 & w9471;
assign w17121 = pi268 & ~w9471;
assign w17122 = ~w17120 & ~w17121;
assign w17123 = ~w504 & w20045;
assign w17124 = (pi221 & w504) | (pi221 & w20046) | (w504 & w20046);
assign w17125 = ~w17123 & ~w17124;
assign w17126 = ~pi301 & ~w16975;
assign w17127 = pi301 & w16975;
assign w17128 = pi532 & pi609;
assign w17129 = ~w17126 & ~w17127;
assign w17130 = ~pi532 & w17129;
assign w17131 = ~w17128 & ~w17130;
assign w17132 = ~pi268 & pi302;
assign w17133 = pi268 & ~pi302;
assign w17134 = ~w17132 & ~w17133;
assign w17135 = w16895 & w17134;
assign w17136 = ~w16895 & ~w17134;
assign w17137 = ~w17135 & ~w17136;
assign w17138 = w16966 & ~w17137;
assign w17139 = ~w16966 & w17137;
assign w17140 = pi532 & pi558;
assign w17141 = ~w17138 & ~w17139;
assign w17142 = ~pi532 & w17141;
assign w17143 = ~w17140 & ~w17142;
assign w17144 = ~pi303 & ~w16966;
assign w17145 = pi303 & w16966;
assign w17146 = pi532 & pi654;
assign w17147 = ~w17144 & ~w17145;
assign w17148 = ~pi532 & w17147;
assign w17149 = ~w17146 & ~w17148;
assign w17150 = ~pi174 & w1367;
assign w17151 = pi174 & ~w1367;
assign w17152 = ~w17150 & ~w17151;
assign w17153 = w7991 & w20047;
assign w17154 = (pi372 & ~w7991) | (pi372 & w20048) | (~w7991 & w20048);
assign w17155 = ~w17153 & ~w17154;
assign w17156 = w4747 & w20049;
assign w17157 = (pi342 & ~w4747) | (pi342 & w20050) | (~w4747 & w20050);
assign w17158 = ~w17156 & ~w17157;
assign w17159 = w7512 & w20051;
assign w17160 = (pi169 & ~w7512) | (pi169 & w20052) | (~w7512 & w20052);
assign w17161 = ~w17159 & ~w17160;
assign w17162 = ~pi183 & w901;
assign w17163 = pi183 & ~w901;
assign w17164 = ~w17162 & ~w17163;
assign w17165 = w1525 & w20053;
assign w17166 = (pi257 & ~w1525) | (pi257 & w20054) | (~w1525 & w20054);
assign w17167 = ~w17165 & ~w17166;
assign w17168 = w700 & w20055;
assign w17169 = (pi258 & ~w700) | (pi258 & w20056) | (~w700 & w20056);
assign w17170 = ~w17168 & ~w17169;
assign w17171 = ~w8898 & w20057;
assign w17172 = (pi320 & w8898) | (pi320 & w20058) | (w8898 & w20058);
assign w17173 = ~w17171 & ~w17172;
assign w17174 = w11809 & w20059;
assign w17175 = (pi274 & ~w11809) | (pi274 & w20060) | (~w11809 & w20060);
assign w17176 = ~w17174 & ~w17175;
assign w17177 = w5777 & w20061;
assign w17178 = (pi348 & ~w5777) | (pi348 & w20062) | (~w5777 & w20062);
assign w17179 = ~w17177 & ~w17178;
assign w17180 = ~pi217 & w5393;
assign w17181 = pi217 & ~w5393;
assign w17182 = ~w17180 & ~w17181;
assign w17183 = w5150 & w20063;
assign w17184 = (pi136 & ~w5150) | (pi136 & w20064) | (~w5150 & w20064);
assign w17185 = ~w17183 & ~w17184;
assign w17186 = w9068 & w20065;
assign w17187 = (pi135 & ~w9068) | (pi135 & w20066) | (~w9068 & w20066);
assign w17188 = ~w17186 & ~w17187;
assign w17189 = w5646 & w20067;
assign w17190 = (pi155 & ~w5646) | (pi155 & w20068) | (~w5646 & w20068);
assign w17191 = ~w17189 & ~w17190;
assign w17192 = w5877 & w20069;
assign w17193 = (pi230 & ~w5877) | (pi230 & w20070) | (~w5877 & w20070);
assign w17194 = ~w17192 & ~w17193;
assign w17195 = ~pi319 & w15942;
assign w17196 = pi319 & ~w15942;
assign w17197 = ~w17195 & ~w17196;
assign w17198 = pi532 & ~pi633;
assign w17199 = ~pi532 & ~w17197;
assign w17200 = ~w17198 & ~w17199;
assign w17201 = ~pi320 & ~w17197;
assign w17202 = pi320 & w17197;
assign w17203 = pi532 & pi601;
assign w17204 = ~w17201 & ~w17202;
assign w17205 = ~pi532 & w17204;
assign w17206 = ~w17203 & ~w17205;
assign w17207 = ~pi321 & w15870;
assign w17208 = pi321 & ~w15870;
assign w17209 = ~w17207 & ~w17208;
assign w17210 = w15942 & ~w17209;
assign w17211 = ~w15942 & w17209;
assign w17212 = pi532 & pi537;
assign w17213 = ~w17210 & ~w17211;
assign w17214 = ~pi532 & w17213;
assign w17215 = ~w17212 & ~w17214;
assign w17216 = w7913 & w20071;
assign w17217 = (pi285 & ~w7913) | (pi285 & w20072) | (~w7913 & w20072);
assign w17218 = ~w17216 & ~w17217;
assign w17219 = ~w3619 & w20073;
assign w17220 = (pi166 & w3619) | (pi166 & w20074) | (w3619 & w20074);
assign w17221 = ~w17219 & ~w17220;
assign w17222 = ~pi272 & w12426;
assign w17223 = pi272 & ~w12426;
assign w17224 = ~w17222 & ~w17223;
assign w17225 = ~w1127 & w20075;
assign w17226 = (pi219 & w1127) | (pi219 & w20076) | (w1127 & w20076);
assign w17227 = ~w17225 & ~w17226;
assign w17228 = ~pi168 & w7576;
assign w17229 = pi168 & ~w7576;
assign w17230 = ~w17228 & ~w17229;
assign w17231 = ~pi208 & w12100;
assign w17232 = pi208 & ~w12100;
assign w17233 = ~w17231 & ~w17232;
assign w17234 = ~w2708 & w20077;
assign w17235 = (pi353 & w2708) | (pi353 & w20078) | (w2708 & w20078);
assign w17236 = ~w17234 & ~w17235;
assign w17237 = w10837 & w20079;
assign w17238 = (pi275 & ~w10837) | (pi275 & w20080) | (~w10837 & w20080);
assign w17239 = ~w17237 & ~w17238;
assign w17240 = w6366 & w20081;
assign w17241 = (pi370 & ~w6366) | (pi370 & w20082) | (~w6366 & w20082);
assign w17242 = ~w17240 & ~w17241;
assign w17243 = ~pi233 & w7220;
assign w17244 = pi233 & ~w7220;
assign w17245 = ~w17243 & ~w17244;
assign w17246 = ~pi215 & w11195;
assign w17247 = pi215 & ~w11195;
assign w17248 = ~w17246 & ~w17247;
assign w17249 = ~pi184 & w8716;
assign w17250 = pi184 & ~w8716;
assign w17251 = ~w17249 & ~w17250;
assign w17252 = ~pi356 & w6711;
assign w17253 = pi356 & ~w6711;
assign w17254 = ~w17252 & ~w17253;
assign w17255 = ~pi350 & w9618;
assign w17256 = pi350 & ~w9618;
assign w17257 = ~w17255 & ~w17256;
assign w17258 = w4539 & w20083;
assign w17259 = (pi175 & ~w4539) | (pi175 & w20084) | (~w4539 & w20084);
assign w17260 = ~w17258 & ~w17259;
assign w17261 = ~pi218 & w5554;
assign w17262 = pi218 & ~w5554;
assign w17263 = ~w17261 & ~w17262;
assign w17264 = w3872 & w20085;
assign w17265 = (pi138 & ~w3872) | (pi138 & w20086) | (~w3872 & w20086);
assign w17266 = ~w17264 & ~w17265;
assign w17267 = ~pi352 & w7123;
assign w17268 = pi352 & ~w7123;
assign w17269 = ~w17267 & ~w17268;
assign w17270 = ~pi185 & w7755;
assign w17271 = pi185 & ~w7755;
assign w17272 = ~w17270 & ~w17271;
assign w17273 = ~pi302 & w11274;
assign w17274 = pi302 & ~w11274;
assign w17275 = ~w17273 & ~w17274;
assign w17276 = ~pi342 & ~w16865;
assign w17277 = pi342 & w16865;
assign w17278 = pi532 & pi540;
assign w17279 = ~w17276 & ~w17277;
assign w17280 = ~pi532 & w17279;
assign w17281 = ~w17278 & ~w17280;
assign w17282 = ~pi209 & w5482;
assign w17283 = pi209 & ~w5482;
assign w17284 = ~w17282 & ~w17283;
assign w17285 = ~pi210 & w12292;
assign w17286 = pi210 & ~w12292;
assign w17287 = ~w17285 & ~w17286;
assign w17288 = ~pi182 & w4641;
assign w17289 = pi182 & ~w4641;
assign w17290 = ~w17288 & ~w17289;
assign w17291 = w16310 & w20087;
assign w17292 = (pi371 & ~w16310) | (pi371 & w20088) | (~w16310 & w20088);
assign w17293 = ~w17291 & ~w17292;
assign w17294 = ~pi346 & ~w17293;
assign w17295 = pi346 & w17293;
assign w17296 = pi532 & pi615;
assign w17297 = ~w17294 & ~w17295;
assign w17298 = ~pi532 & w17297;
assign w17299 = ~w17296 & ~w17298;
assign w17300 = w2429 & w20089;
assign w17301 = (pi373 & ~w2429) | (pi373 & w20090) | (~w2429 & w20090);
assign w17302 = ~w17300 & ~w17301;
assign w17303 = pi348 & w16859;
assign w17304 = ~pi348 & ~w16859;
assign w17305 = pi532 & pi604;
assign w17306 = ~w17303 & ~w17304;
assign w17307 = ~pi532 & w17306;
assign w17308 = ~w17305 & ~w17307;
assign w17309 = w16375 & w20091;
assign w17310 = (pi349 & ~w16375) | (pi349 & w20092) | (~w16375 & w20092);
assign w17311 = ~w17309 & ~w17310;
assign w17312 = pi532 & ~pi631;
assign w17313 = ~pi532 & ~w17311;
assign w17314 = ~w17312 & ~w17313;
assign w17315 = ~pi350 & ~w17311;
assign w17316 = pi350 & w17311;
assign w17317 = pi532 & pi599;
assign w17318 = ~w17315 & ~w17316;
assign w17319 = ~pi532 & w17318;
assign w17320 = ~w17317 & ~w17319;
assign w17321 = ~pi351 & w16249;
assign w17322 = pi351 & ~w16249;
assign w17323 = ~w17321 & ~w17322;
assign w17324 = w16310 & w20093;
assign w17325 = (w17323 & ~w16310) | (w17323 & w20094) | (~w16310 & w20094);
assign w17326 = pi532 & pi551;
assign w17327 = ~w17324 & ~w17325;
assign w17328 = ~pi532 & w17327;
assign w17329 = ~w17326 & ~w17328;
assign w17330 = ~pi352 & w16381;
assign w17331 = pi352 & ~w16381;
assign w17332 = ~w17330 & ~w17331;
assign w17333 = w16375 & w20095;
assign w17334 = (w17332 & ~w16375) | (w17332 & w20096) | (~w16375 & w20096);
assign w17335 = pi532 & pi535;
assign w17336 = ~w17333 & ~w17334;
assign w17337 = ~pi532 & w17336;
assign w17338 = ~w17335 & ~w17337;
assign w17339 = pi532 & pi652;
assign w17340 = ~pi532 & w16452;
assign w17341 = ~w17339 & ~w17340;
assign w17342 = ~pi354 & ~w16458;
assign w17343 = pi354 & w16458;
assign w17344 = pi532 & pi556;
assign w17345 = ~w17342 & ~w17343;
assign w17346 = ~pi532 & w17345;
assign w17347 = ~w17344 & ~w17346;
assign w17348 = w10661 & w20097;
assign w17349 = (pi171 & ~w10661) | (pi171 & w20098) | (~w10661 & w20098);
assign w17350 = ~w17348 & ~w17349;
assign w17351 = ~w16523 & w20099;
assign w17352 = (pi356 & w16523) | (pi356 & w20100) | (w16523 & w20100);
assign w17353 = ~w17351 & ~w17352;
assign w17354 = pi532 & ~pi649;
assign w17355 = ~pi532 & ~w17353;
assign w17356 = ~w17354 & ~w17355;
assign w17357 = ~pi357 & ~w17353;
assign w17358 = pi357 & w17353;
assign w17359 = pi532 & pi617;
assign w17360 = ~w17357 & ~w17358;
assign w17361 = ~pi532 & w17360;
assign w17362 = ~w17359 & ~w17361;
assign w17363 = ~pi358 & w16531;
assign w17364 = pi358 & ~w16531;
assign w17365 = ~w17363 & ~w17364;
assign w17366 = ~w16523 & w20101;
assign w17367 = (w17365 & w16523) | (w17365 & w20102) | (w16523 & w20102);
assign w17368 = pi532 & pi553;
assign w17369 = ~w17366 & ~w17367;
assign w17370 = ~pi532 & w17369;
assign w17371 = ~w17368 & ~w17370;
assign w17372 = ~pi376 & w3353;
assign w17373 = pi376 & ~w3353;
assign w17374 = ~w17372 & ~w17373;
assign w17375 = ~w988 & w20103;
assign w17376 = (pi165 & w988) | (pi165 & w20104) | (w988 & w20104);
assign w17377 = ~w17375 & ~w17376;
assign w17378 = ~pi187 & w6948;
assign w17379 = pi187 & ~w6948;
assign w17380 = ~w17378 & ~w17379;
assign w17381 = ~pi278 & w3199;
assign w17382 = pi278 & ~w3199;
assign w17383 = ~w17381 & ~w17382;
assign w17384 = ~w2556 & w20105;
assign w17385 = (pi161 & w2556) | (pi161 & w20106) | (w2556 & w20106);
assign w17386 = ~w17384 & ~w17385;
assign w17387 = w10393 & w20107;
assign w17388 = (pi271 & ~w10393) | (pi271 & w20108) | (~w10393 & w20108);
assign w17389 = ~w17387 & ~w17388;
assign w17390 = w4439 & w20109;
assign w17391 = (pi207 & ~w4439) | (pi207 & w20110) | (~w4439 & w20110);
assign w17392 = ~w17390 & ~w17391;
assign w17393 = ~pi349 & w6530;
assign w17394 = pi349 & ~w6530;
assign w17395 = ~w17393 & ~w17394;
assign w17396 = ~pi220 & w402;
assign w17397 = pi220 & ~w402;
assign w17398 = ~w17396 & ~w17397;
assign w17399 = w8615 & w20111;
assign w17400 = (pi357 & ~w8615) | (pi357 & w20112) | (~w8615 & w20112);
assign w17401 = ~w17399 & ~w17400;
assign w17402 = ~w1649 & w20113;
assign w17403 = (pi163 & w1649) | (pi163 & w20114) | (w1649 & w20114);
assign w17404 = ~w17402 & ~w17403;
assign w17405 = pi532 & pi636;
assign w17406 = ~pi532 & w16859;
assign w17407 = ~w17405 & ~w17406;
assign w17408 = pi532 & ~pi647;
assign w17409 = ~pi532 & ~w17293;
assign w17410 = ~w17408 & ~w17409;
assign w17411 = ~pi372 & ~w16791;
assign w17412 = pi372 & w16791;
assign w17413 = pi532 & pi534;
assign w17414 = ~w17411 & ~w17412;
assign w17415 = ~pi532 & w17414;
assign w17416 = ~w17413 & ~w17415;
assign w17417 = pi373 & w16785;
assign w17418 = ~pi373 & ~w16785;
assign w17419 = pi532 & pi598;
assign w17420 = ~w17417 & ~w17418;
assign w17421 = ~pi532 & w17420;
assign w17422 = ~w17419 & ~w17421;
assign w17423 = ~pi358 & w3968;
assign w17424 = pi358 & ~w3968;
assign w17425 = ~w17423 & ~w17424;
assign w17426 = pi375 & w16452;
assign w17427 = ~pi375 & ~w16452;
assign w17428 = pi532 & pi620;
assign w17429 = ~w17426 & ~w17427;
assign w17430 = ~pi532 & w17429;
assign w17431 = ~w17428 & ~w17430;
assign w17432 = pi532 & pi630;
assign w17433 = ~pi532 & w16785;
assign w17434 = ~w17432 & ~w17433;
assign w17435 = w11699 & w20115;
assign w17436 = (pi273 & ~w11699) | (pi273 & w20116) | (~w11699 & w20116);
assign w17437 = ~w17435 & ~w17436;
assign w17438 = ~pi281 & w2286;
assign w17439 = pi281 & ~w2286;
assign w17440 = ~w17438 & ~w17439;
assign w17441 = ~pi181 & w6453;
assign w17442 = pi181 & ~w6453;
assign w17443 = ~w17441 & ~w17442;
assign w17444 = ~w1803 & w20117;
assign w17445 = (pi375 & w1803) | (pi375 & w20118) | (w1803 & w20118);
assign w17446 = ~w17444 & ~w17445;
assign w17447 = ~pi284 & w7845;
assign w17448 = pi284 & ~w7845;
assign w17449 = ~w17447 & ~w17448;
assign w17450 = w1438 & w20119;
assign w17451 = (pi173 & ~w1438) | (pi173 & w20120) | (~w1438 & w20120);
assign w17452 = ~w17450 & ~w17451;
assign w17453 = w4920 & w20121;
assign w17454 = (pi234 & ~w4920) | (pi234 & w20122) | (~w4920 & w20122);
assign w17455 = ~w17453 & ~w17454;
assign w17456 = pi487 & pi520;
assign w17457 = pi482 & w17456;
assign w17458 = (~pi396 & ~w17456) | (~pi396 & w17471) | (~w17456 & w17471);
assign w17459 = ~pi482 & ~w17456;
assign w17460 = ~w17457 & ~w17459;
assign w17461 = w17456 & w20123;
assign w17462 = ~pi487 & ~pi520;
assign w17463 = ~w17456 & ~w17462;
assign w17464 = ~w17460 & w20124;
assign w17465 = ~w17458 & w17464;
assign w17466 = (w17464 & w20125) | (w17464 & w20126) | (w20125 & w20126);
assign w17467 = ~pi396 & w17460;
assign w17468 = w17460 & w20127;
assign w17469 = ~w17465 & ~w17468;
assign w17470 = w17466 & ~w17469;
assign w17471 = ~pi396 & ~pi482;
assign w17472 = (pi520 & ~w17471) | (pi520 & w17456) | (~w17471 & w17456);
assign w17473 = w17466 & ~w17472;
assign w17474 = (~pi520 & ~w17471) | (~pi520 & w17462) | (~w17471 & w17462);
assign w17475 = ~pi520 & ~pi532;
assign w17476 = ~pi532 & w17464;
assign w17477 = (~w17475 & ~w17464) | (~w17475 & w20128) | (~w17464 & w20128);
assign w17478 = ~w17474 & ~w17477;
assign w17479 = ~pi393 & ~pi395;
assign w17480 = (pi387 & ~w17479) | (pi387 & w20129) | (~w17479 & w20129);
assign w17481 = ~pi532 & ~w17480;
assign w17482 = pi531 & ~w17481;
assign w17483 = ~w17469 & w17475;
assign w17484 = pi390 & ~w17479;
assign w17485 = w17479 & w20130;
assign w17486 = ~w17484 & ~w17485;
assign w17487 = pi531 & ~pi532;
assign w17488 = ~w17486 & w17487;
assign w17489 = ~pi532 & w17463;
assign w17490 = w17467 & w17489;
assign w17491 = pi520 & w17490;
assign w17492 = ~pi520 & w17490;
assign w17493 = ~pi387 & ~pi390;
assign w17494 = pi393 & pi395;
assign w17495 = ~pi532 & ~w17494;
assign w17496 = w17479 & ~w17493;
assign w17497 = w17495 & ~w17496;
assign w17498 = pi531 & ~w17497;
assign w17499 = ~pi532 & ~w17457;
assign w17500 = ~pi393 & w17493;
assign w17501 = (~pi395 & ~w17493) | (~pi395 & w20131) | (~w17493 & w20131);
assign w17502 = ~pi532 & ~w17501;
assign w17503 = pi531 & ~w17502;
assign w17504 = ~w17458 & ~w17461;
assign w17505 = ~pi532 & w17504;
assign w17506 = pi395 & ~pi532;
assign w17507 = w17500 & w17506;
assign w17508 = pi398 & ~pi532;
assign w17509 = pi532 & pi777;
assign w17510 = ~w17508 & ~w17509;
assign w17511 = pi399 & ~pi532;
assign w17512 = pi532 & pi772;
assign w17513 = ~w17511 & ~w17512;
assign w17514 = pi400 & ~pi532;
assign w17515 = pi532 & pi698;
assign w17516 = ~w17514 & ~w17515;
assign w17517 = pi401 & ~pi532;
assign w17518 = pi532 & pi675;
assign w17519 = ~w17517 & ~w17518;
assign w17520 = pi402 & ~pi532;
assign w17521 = pi532 & pi728;
assign w17522 = ~w17520 & ~w17521;
assign w17523 = pi403 & ~pi532;
assign w17524 = pi532 & pi708;
assign w17525 = ~w17523 & ~w17524;
assign w17526 = pi404 & ~pi532;
assign w17527 = pi532 & pi679;
assign w17528 = ~w17526 & ~w17527;
assign w17529 = pi405 & ~pi532;
assign w17530 = pi532 & pi661;
assign w17531 = ~w17529 & ~w17530;
assign w17532 = pi406 & ~pi532;
assign w17533 = pi532 & pi729;
assign w17534 = ~w17532 & ~w17533;
assign w17535 = pi407 & ~pi532;
assign w17536 = pi532 & pi710;
assign w17537 = ~w17535 & ~w17536;
assign w17538 = pi408 & ~pi532;
assign w17539 = pi532 & pi703;
assign w17540 = ~w17538 & ~w17539;
assign w17541 = pi409 & ~pi532;
assign w17542 = pi532 & pi788;
assign w17543 = ~w17541 & ~w17542;
assign w17544 = pi410 & ~pi532;
assign w17545 = pi532 & pi725;
assign w17546 = ~w17544 & ~w17545;
assign w17547 = pi411 & ~pi532;
assign w17548 = pi532 & pi715;
assign w17549 = ~w17547 & ~w17548;
assign w17550 = pi412 & ~pi532;
assign w17551 = pi532 & pi696;
assign w17552 = ~w17550 & ~w17551;
assign w17553 = pi413 & ~pi532;
assign w17554 = pi532 & pi667;
assign w17555 = ~w17553 & ~w17554;
assign w17556 = pi414 & ~pi532;
assign w17557 = pi532 & pi678;
assign w17558 = ~w17556 & ~w17557;
assign w17559 = pi415 & ~pi532;
assign w17560 = pi532 & pi769;
assign w17561 = ~w17559 & ~w17560;
assign w17562 = pi416 & ~pi532;
assign w17563 = pi532 & pi672;
assign w17564 = ~w17562 & ~w17563;
assign w17565 = pi417 & ~pi532;
assign w17566 = pi532 & pi784;
assign w17567 = ~w17565 & ~w17566;
assign w17568 = pi418 & ~pi532;
assign w17569 = pi532 & pi685;
assign w17570 = ~w17568 & ~w17569;
assign w17571 = pi419 & ~pi532;
assign w17572 = pi532 & pi687;
assign w17573 = ~w17571 & ~w17572;
assign w17574 = pi420 & ~pi532;
assign w17575 = pi532 & pi690;
assign w17576 = ~w17574 & ~w17575;
assign w17577 = pi421 & ~pi532;
assign w17578 = pi532 & pi707;
assign w17579 = ~w17577 & ~w17578;
assign w17580 = pi422 & ~pi532;
assign w17581 = pi532 & pi716;
assign w17582 = ~w17580 & ~w17581;
assign w17583 = pi423 & ~pi532;
assign w17584 = pi532 & pi722;
assign w17585 = ~w17583 & ~w17584;
assign w17586 = pi424 & ~pi532;
assign w17587 = pi532 & pi724;
assign w17588 = ~w17586 & ~w17587;
assign w17589 = pi425 & ~pi532;
assign w17590 = pi532 & pi739;
assign w17591 = ~w17589 & ~w17590;
assign w17592 = pi426 & ~pi532;
assign w17593 = pi532 & pi742;
assign w17594 = ~w17592 & ~w17593;
assign w17595 = pi427 & ~pi532;
assign w17596 = pi532 & pi747;
assign w17597 = ~w17595 & ~w17596;
assign w17598 = pi428 & ~pi532;
assign w17599 = pi532 & pi669;
assign w17600 = ~w17598 & ~w17599;
assign w17601 = pi429 & ~pi532;
assign w17602 = pi532 & pi760;
assign w17603 = ~w17601 & ~w17602;
assign w17604 = pi430 & ~pi532;
assign w17605 = pi532 & pi752;
assign w17606 = ~w17604 & ~w17605;
assign w17607 = pi431 & ~pi532;
assign w17608 = pi532 & pi700;
assign w17609 = ~w17607 & ~w17608;
assign w17610 = pi432 & ~pi532;
assign w17611 = pi532 & pi721;
assign w17612 = ~w17610 & ~w17611;
assign w17613 = pi433 & ~pi532;
assign w17614 = pi532 & pi764;
assign w17615 = ~w17613 & ~w17614;
assign w17616 = pi434 & ~pi532;
assign w17617 = pi532 & pi684;
assign w17618 = ~w17616 & ~w17617;
assign w17619 = pi435 & ~pi532;
assign w17620 = pi532 & pi719;
assign w17621 = ~w17619 & ~w17620;
assign w17622 = pi436 & ~pi532;
assign w17623 = pi532 & pi664;
assign w17624 = ~w17622 & ~w17623;
assign w17625 = pi437 & ~pi532;
assign w17626 = pi532 & pi779;
assign w17627 = ~w17625 & ~w17626;
assign w17628 = pi438 & ~pi532;
assign w17629 = pi532 & pi720;
assign w17630 = ~w17628 & ~w17629;
assign w17631 = pi439 & ~pi532;
assign w17632 = pi532 & pi757;
assign w17633 = ~w17631 & ~w17632;
assign w17634 = pi440 & ~pi532;
assign w17635 = pi532 & pi731;
assign w17636 = ~w17634 & ~w17635;
assign w17637 = pi441 & ~pi532;
assign w17638 = pi532 & pi712;
assign w17639 = ~w17637 & ~w17638;
assign w17640 = pi442 & ~pi532;
assign w17641 = pi532 & pi753;
assign w17642 = ~w17640 & ~w17641;
assign w17643 = pi443 & ~pi532;
assign w17644 = pi532 & pi768;
assign w17645 = ~w17643 & ~w17644;
assign w17646 = pi444 & ~pi532;
assign w17647 = pi532 & pi689;
assign w17648 = ~w17646 & ~w17647;
assign w17649 = pi445 & ~pi532;
assign w17650 = pi532 & pi738;
assign w17651 = ~w17649 & ~w17650;
assign w17652 = pi446 & ~pi532;
assign w17653 = pi532 & pi662;
assign w17654 = ~w17652 & ~w17653;
assign w17655 = pi447 & ~pi532;
assign w17656 = pi532 & pi680;
assign w17657 = ~w17655 & ~w17656;
assign w17658 = pi448 & ~pi532;
assign w17659 = pi532 & pi717;
assign w17660 = ~w17658 & ~w17659;
assign w17661 = pi449 & ~pi532;
assign w17662 = pi532 & pi751;
assign w17663 = ~w17661 & ~w17662;
assign w17664 = pi450 & ~pi532;
assign w17665 = pi532 & pi730;
assign w17666 = ~w17664 & ~w17665;
assign w17667 = pi451 & ~pi532;
assign w17668 = pi532 & pi673;
assign w17669 = ~w17667 & ~w17668;
assign w17670 = pi452 & ~pi532;
assign w17671 = pi532 & pi746;
assign w17672 = ~w17670 & ~w17671;
assign w17673 = pi453 & ~pi532;
assign w17674 = pi532 & pi741;
assign w17675 = ~w17673 & ~w17674;
assign w17676 = pi454 & ~pi532;
assign w17677 = pi532 & pi727;
assign w17678 = ~w17676 & ~w17677;
assign w17679 = pi455 & ~pi532;
assign w17680 = pi532 & pi670;
assign w17681 = ~w17679 & ~w17680;
assign w17682 = pi456 & ~pi532;
assign w17683 = pi532 & pi714;
assign w17684 = ~w17682 & ~w17683;
assign w17685 = pi457 & ~pi532;
assign w17686 = pi532 & pi706;
assign w17687 = ~w17685 & ~w17686;
assign w17688 = pi458 & ~pi532;
assign w17689 = pi532 & pi713;
assign w17690 = ~w17688 & ~w17689;
assign w17691 = pi459 & ~pi532;
assign w17692 = pi532 & pi758;
assign w17693 = ~w17691 & ~w17692;
assign w17694 = pi460 & ~pi532;
assign w17695 = pi532 & pi671;
assign w17696 = ~w17694 & ~w17695;
assign w17697 = pi461 & ~pi532;
assign w17698 = pi532 & pi695;
assign w17699 = ~w17697 & ~w17698;
assign w17700 = pi462 & ~pi532;
assign w17701 = pi532 & pi771;
assign w17702 = ~w17700 & ~w17701;
assign w17703 = pi463 & ~pi532;
assign w17704 = pi532 & pi691;
assign w17705 = ~w17703 & ~w17704;
assign w17706 = pi464 & ~pi532;
assign w17707 = pi532 & pi765;
assign w17708 = ~w17706 & ~w17707;
assign w17709 = pi465 & ~pi532;
assign w17710 = pi532 & pi726;
assign w17711 = ~w17709 & ~w17710;
assign w17712 = pi466 & ~pi532;
assign w17713 = pi532 & pi740;
assign w17714 = ~w17712 & ~w17713;
assign w17715 = pi467 & ~pi532;
assign w17716 = pi532 & pi668;
assign w17717 = ~w17715 & ~w17716;
assign w17718 = pi468 & ~pi532;
assign w17719 = pi532 & pi743;
assign w17720 = ~w17718 & ~w17719;
assign w17721 = pi469 & ~pi532;
assign w17722 = pi532 & pi787;
assign w17723 = ~w17721 & ~w17722;
assign w17724 = pi470 & ~pi532;
assign w17725 = pi532 & pi766;
assign w17726 = ~w17724 & ~w17725;
assign w17727 = pi471 & ~pi532;
assign w17728 = pi532 & pi674;
assign w17729 = ~w17727 & ~w17728;
assign w17730 = pi472 & ~pi532;
assign w17731 = pi532 & pi781;
assign w17732 = ~w17730 & ~w17731;
assign w17733 = pi473 & ~pi532;
assign w17734 = pi532 & pi745;
assign w17735 = ~w17733 & ~w17734;
assign w17736 = pi474 & ~pi532;
assign w17737 = pi532 & pi735;
assign w17738 = ~w17736 & ~w17737;
assign w17739 = pi475 & ~pi532;
assign w17740 = pi532 & pi677;
assign w17741 = ~w17739 & ~w17740;
assign w17742 = pi476 & ~pi532;
assign w17743 = pi532 & pi701;
assign w17744 = ~w17742 & ~w17743;
assign w17745 = pi477 & ~pi532;
assign w17746 = pi532 & pi676;
assign w17747 = ~w17745 & ~w17746;
assign w17748 = pi478 & ~pi532;
assign w17749 = pi532 & pi782;
assign w17750 = ~w17748 & ~w17749;
assign w17751 = pi479 & ~pi532;
assign w17752 = pi532 & pi702;
assign w17753 = ~w17751 & ~w17752;
assign w17754 = pi480 & ~pi532;
assign w17755 = pi532 & pi697;
assign w17756 = ~w17754 & ~w17755;
assign w17757 = pi481 & ~pi532;
assign w17758 = pi532 & pi681;
assign w17759 = ~w17757 & ~w17758;
assign w17760 = ~pi532 & w17460;
assign w17761 = pi483 & ~pi532;
assign w17762 = pi532 & pi693;
assign w17763 = ~w17761 & ~w17762;
assign w17764 = pi484 & ~pi532;
assign w17765 = pi532 & pi736;
assign w17766 = ~w17764 & ~w17765;
assign w17767 = pi485 & ~pi532;
assign w17768 = pi532 & pi749;
assign w17769 = ~w17767 & ~w17768;
assign w17770 = pi486 & ~pi532;
assign w17771 = pi532 & pi694;
assign w17772 = ~w17770 & ~w17771;
assign w17773 = pi488 & ~pi532;
assign w17774 = pi532 & pi786;
assign w17775 = ~w17773 & ~w17774;
assign w17776 = pi489 & ~pi532;
assign w17777 = pi532 & pi663;
assign w17778 = ~w17776 & ~w17777;
assign w17779 = pi490 & ~pi532;
assign w17780 = pi532 & pi705;
assign w17781 = ~w17779 & ~w17780;
assign w17782 = pi491 & ~pi532;
assign w17783 = pi532 & pi733;
assign w17784 = ~w17782 & ~w17783;
assign w17785 = pi492 & ~pi532;
assign w17786 = pi532 & pi762;
assign w17787 = ~w17785 & ~w17786;
assign w17788 = pi493 & ~pi532;
assign w17789 = pi532 & pi767;
assign w17790 = ~w17788 & ~w17789;
assign w17791 = pi494 & ~pi532;
assign w17792 = pi532 & pi665;
assign w17793 = ~w17791 & ~w17792;
assign w17794 = pi495 & ~pi532;
assign w17795 = pi532 & pi704;
assign w17796 = ~w17794 & ~w17795;
assign w17797 = pi496 & ~pi532;
assign w17798 = pi532 & pi773;
assign w17799 = ~w17797 & ~w17798;
assign w17800 = pi497 & ~pi532;
assign w17801 = pi532 & pi754;
assign w17802 = ~w17800 & ~w17801;
assign w17803 = pi498 & ~pi532;
assign w17804 = pi532 & pi734;
assign w17805 = ~w17803 & ~w17804;
assign w17806 = pi499 & ~pi532;
assign w17807 = pi532 & pi711;
assign w17808 = ~w17806 & ~w17807;
assign w17809 = pi500 & ~pi532;
assign w17810 = pi532 & pi761;
assign w17811 = ~w17809 & ~w17810;
assign w17812 = pi501 & ~pi532;
assign w17813 = pi532 & pi775;
assign w17814 = ~w17812 & ~w17813;
assign w17815 = pi502 & ~pi532;
assign w17816 = pi532 & pi686;
assign w17817 = ~w17815 & ~w17816;
assign w17818 = pi503 & ~pi532;
assign w17819 = pi532 & pi718;
assign w17820 = ~w17818 & ~w17819;
assign w17821 = pi504 & ~pi532;
assign w17822 = pi532 & pi756;
assign w17823 = ~w17821 & ~w17822;
assign w17824 = pi505 & ~pi532;
assign w17825 = pi532 & pi785;
assign w17826 = ~w17824 & ~w17825;
assign w17827 = pi506 & ~pi532;
assign w17828 = pi532 & pi776;
assign w17829 = ~w17827 & ~w17828;
assign w17830 = pi507 & ~pi532;
assign w17831 = pi532 & pi759;
assign w17832 = ~w17830 & ~w17831;
assign w17833 = pi508 & ~pi532;
assign w17834 = pi532 & pi692;
assign w17835 = ~w17833 & ~w17834;
assign w17836 = pi509 & ~pi532;
assign w17837 = pi532 & pi783;
assign w17838 = ~w17836 & ~w17837;
assign w17839 = pi510 & ~pi532;
assign w17840 = pi532 & pi780;
assign w17841 = ~w17839 & ~w17840;
assign w17842 = pi511 & ~pi532;
assign w17843 = pi532 & pi763;
assign w17844 = ~w17842 & ~w17843;
assign w17845 = pi512 & ~pi532;
assign w17846 = pi532 & pi737;
assign w17847 = ~w17845 & ~w17846;
assign w17848 = pi513 & ~pi532;
assign w17849 = pi532 & pi774;
assign w17850 = ~w17848 & ~w17849;
assign w17851 = pi514 & ~pi532;
assign w17852 = pi532 & pi755;
assign w17853 = ~w17851 & ~w17852;
assign w17854 = pi515 & ~pi532;
assign w17855 = pi532 & pi723;
assign w17856 = ~w17854 & ~w17855;
assign w17857 = pi516 & ~pi532;
assign w17858 = pi532 & pi709;
assign w17859 = ~w17857 & ~w17858;
assign w17860 = pi517 & ~pi532;
assign w17861 = pi532 & pi688;
assign w17862 = ~w17860 & ~w17861;
assign w17863 = pi518 & ~pi532;
assign w17864 = pi532 & pi770;
assign w17865 = ~w17863 & ~w17864;
assign w17866 = pi519 & ~pi532;
assign w17867 = pi532 & pi778;
assign w17868 = ~w17866 & ~w17867;
assign w17869 = pi521 & ~pi532;
assign w17870 = pi532 & pi682;
assign w17871 = ~w17869 & ~w17870;
assign w17872 = pi522 & ~pi532;
assign w17873 = pi532 & pi666;
assign w17874 = ~w17872 & ~w17873;
assign w17875 = pi523 & ~pi532;
assign w17876 = pi532 & pi683;
assign w17877 = ~w17875 & ~w17876;
assign w17878 = pi524 & ~pi532;
assign w17879 = pi532 & pi744;
assign w17880 = ~w17878 & ~w17879;
assign w17881 = pi525 & ~pi532;
assign w17882 = pi532 & pi699;
assign w17883 = ~w17881 & ~w17882;
assign w17884 = pi526 & ~pi532;
assign w17885 = pi532 & pi732;
assign w17886 = ~w17884 & ~w17885;
assign w17887 = pi527 & ~pi532;
assign w17888 = pi532 & pi750;
assign w17889 = ~w17887 & ~w17888;
assign w17890 = pi528 & ~pi532;
assign w17891 = pi532 & pi748;
assign w17892 = ~w17890 & ~w17891;
assign w17893 = pi107 & ~pi108;
assign w17894 = w29 & w20132;
assign w17895 = w33 & w36;
assign w17896 = w51 & w46;
assign w17897 = w2 & w18458;
assign w17898 = (~w59 & w234) | (~w59 & w20133) | (w234 & w20133);
assign w17899 = w73 & pi083;
assign w17900 = w25 & w70;
assign w17901 = (~w68 & w20134) | (~w68 & w20135) | (w20134 & w20135);
assign w17902 = pi014 & pi072;
assign w17903 = ~w124 & ~w125;
assign w17904 = (~w19 & w20136) | (~w19 & w20137) | (w20136 & w20137);
assign w17905 = w146 & pi083;
assign w17906 = ~pi072 & ~pi083;
assign w17907 = ~w161 & w20138;
assign w17908 = ~w174 & ~w171;
assign w17909 = w178 & w177;
assign w17910 = w149 & pi040;
assign w17911 = w187 & w78;
assign w17912 = w212 & ~pi083;
assign w17913 = (w190 & w88) | (w190 & w20139) | (w88 & w20139);
assign w17914 = w222 & w84;
assign w17915 = (~pi083 & ~w227) | (~pi083 & w20140) | (~w227 & w20140);
assign w17916 = w224 & pi040;
assign w17917 = w78 & pi108;
assign w17918 = ~w240 & ~w241;
assign w17919 = (~w198 & w20136) | (~w198 & w20141) | (w20136 & w20141);
assign w17920 = w186 & pi078;
assign w17921 = w278 & ~pi123;
assign w17922 = ~w256 & w17925;
assign w17923 = ~w270 & pi048;
assign w17924 = w310 & ~w316;
assign w17925 = pi111 & pi123;
assign w17926 = pi111 & pi027;
assign w17927 = pi123 & ~w362;
assign w17928 = pi027 & ~pi020;
assign w17929 = w347 & pi048;
assign w17930 = w380 & ~pi123;
assign w17931 = w383 & w285;
assign w17932 = ~w385 & ~w390;
assign w17933 = ~pi048 & w399;
assign w17934 = w400 & ~w401;
assign w17935 = pi054 & ~pi114;
assign w17936 = w467 & w479;
assign w17937 = pi054 & pi114;
assign w17938 = pi054 & pi013;
assign w17939 = pi114 & ~w496;
assign w17940 = ~pi054 & ~pi029;
assign w17941 = w501 & ~w473;
assign w17942 = pi054 & ~pi013;
assign w17943 = ~w513 & pi114;
assign w17944 = w477 & pi013;
assign w17945 = ~w514 & ~w518;
assign w17946 = w533 & ~pi114;
assign w17947 = ~w536 & pi001;
assign w17948 = ~w518 & w547;
assign w17949 = w567 & w20142;
assign w17950 = pi127 & ~pi126;
assign w17951 = w590 & ~pi104;
assign w17952 = w593 & ~pi127;
assign w17953 = w598 & w597;
assign w17954 = w608 & w604;
assign w17955 = w614 & w20143;
assign w17956 = ~pi126 & ~pi104;
assign w17957 = (~w616 & w17964) | (~w616 & w20144) | (w17964 & w20144);
assign w17958 = w584 & w617;
assign w17959 = w653 & pi104;
assign w17960 = w646 & pi126;
assign w17961 = w661 & ~pi069;
assign w17962 = ~w669 & ~w671;
assign w17963 = ~w675 & ~w676;
assign w17964 = ~pi104 & ~pi102;
assign w17965 = ~w695 & ~w673;
assign w17966 = (~w632 & w20145) | (~w632 & w20146) | (w20145 & w20146);
assign w17967 = w610 & ~pi012;
assign w17968 = ~pi126 & pi104;
assign w17969 = w719 & pi104;
assign w17970 = ~pi033 & ~pi104;
assign w17971 = w721 & pi102;
assign w17972 = w736 & w570;
assign w17973 = ~w740 & ~w742;
assign w17974 = (~w716 & w20145) | (~w716 & w20148) | (w20145 & w20148);
assign w17975 = w683 & w639;
assign w17976 = w765 & ~pi104;
assign w17977 = (w747 & w645) | (w747 & w20916) | (w645 & w20916);
assign w17978 = w741 & pi104;
assign w17979 = w779 & w622;
assign w17980 = w624 & ~pi104;
assign w17981 = w785 & pi102;
assign w17982 = (~w754 & w20917) | (~w754 & w20918) | (w20917 & w20918);
assign w17983 = w812 & w703;
assign w17984 = ~w566 & pi102;
assign w17985 = w708 & ~pi104;
assign w17986 = pi127 & ~pi012;
assign w17987 = pi102 & w869;
assign w17988 = ~w588 & pi102;
assign w17989 = ~w893 & ~w888;
assign w17990 = ~w907 & ~pi529;
assign w17991 = w922 & pi001;
assign w17992 = w938 & ~pi114;
assign w17993 = ~w448 & ~pi029;
assign w17994 = ~w956 & pi001;
assign w17995 = ~w475 & ~w515;
assign w17996 = ~w960 & w20149;
assign w17997 = w970 & pi114;
assign w17998 = w999 & pi013;
assign w17999 = w1005 & ~pi114;
assign w18000 = w1004 & ~pi001;
assign w18001 = w1036 & ~pi123;
assign w18002 = pi023 & ~pi093;
assign w18003 = pi027 & ~w1049;
assign w18004 = ~w1053 & pi020;
assign w18005 = ~pi111 & pi123;
assign w18006 = ~w1076 & ~pi048;
assign w18007 = ~w383 & ~pi020;
assign w18008 = ~w1077 & ~w1079;
assign w18009 = w1022 & pi093;
assign w18010 = w1103 & pi027;
assign w18011 = ~w1119 & ~w1120;
assign w18012 = w487 & pi007;
assign w18013 = w475 & pi001;
assign w18014 = w1139 & ~pi114;
assign w18015 = (~pi001 & w1137) | (~pi001 & w20150) | (w1137 & w20150);
assign w18016 = w434 & ~pi001;
assign w18017 = w403 & ~pi114;
assign w18018 = ~w1186 & ~w1185;
assign w18019 = w507 & w5474;
assign w18020 = ~w1189 & ~pi001;
assign w18021 = ~w1167 & w7344;
assign w18022 = w1159 & pi029;
assign w18023 = w326 & pi048;
assign w18024 = ~w1207 & ~w1082;
assign w18025 = w1049 & pi123;
assign w18026 = w1215 & ~pi048;
assign w18027 = ~pi111 & ~w259;
assign w18028 = ~w1243 & w1256;
assign w18029 = w1259 & w20151;
assign w18030 = ~w1266 & ~pi048;
assign w18031 = w324 & pi123;
assign w18032 = w1268 & pi048;
assign w18033 = w1273 & w1118;
assign w18034 = w1276 & ~w1275;
assign w18035 = w1289 & ~pi083;
assign w18036 = w1298 & ~pi083;
assign w18037 = w50 & w8;
assign w18038 = w164 & ~pi108;
assign w18039 = w1313 & ~w166;
assign w18040 = w1291 & ~pi040;
assign w18041 = w7 & w177;
assign w18042 = w1326 & ~pi040;
assign w18043 = ~w1321 & w20152;
assign w18044 = ~w42 & ~w4;
assign w18045 = ~w1343 & ~pi040;
assign w18046 = w16 & w20153;
assign w18047 = w1352 & w1348;
assign w18048 = w40 & pi083;
assign w18049 = w1317 & ~pi078;
assign w18050 = w257 & w318;
assign w18051 = w1229 & ~pi123;
assign w18052 = w281 & w343;
assign w18053 = w1381 & ~pi048;
assign w18054 = (~w1033 & w1420) | (~w1033 & w20154) | (w1420 & w20154);
assign w18055 = w274 & w383;
assign w18056 = w1081 & ~pi027;
assign w18057 = w1396 & w20155;
assign w18058 = ~w1395 & w20216;
assign w18059 = ~w1074 & ~w1064;
assign w18060 = ~w1414 & ~pi048;
assign w18061 = w364 & w20156;
assign w18062 = w1427 & w1426;
assign w18063 = ~w1419 & ~w1425;
assign w18064 = (~w1373 & w20157) | (~w1373 & w20158) | (w20157 & w20158);
assign w18065 = w1444 & ~pi104;
assign w18066 = w1454 & ~pi104;
assign w18067 = w579 & ~pi069;
assign w18068 = w1458 & pi102;
assign w18069 = w1446 & ~pi102;
assign w18070 = w566 & w20159;
assign w18071 = w1487 & ~pi102;
assign w18072 = ~w1482 & w20160;
assign w18073 = pi104 & ~w1503;
assign w18074 = pi104 & ~w1507;
assign w18075 = w567 & w20161;
assign w18076 = w794 & w597;
assign w18077 = ~w1522 & ~w1523;
assign w18078 = w1478 & ~pi012;
assign w18079 = ~w1526 & ~pi267;
assign w18080 = w1526 & pi267;
assign w18081 = pi117 & ~w1560;
assign w18082 = pi032 & ~pi105;
assign w18083 = w1573 & w20162;
assign w18084 = w1583 & w1577;
assign w18085 = (pi117 & ~w1610) | (pi117 & w20163) | (~w1610 & w20163);
assign w18086 = ~w1613 & w1647;
assign w18087 = w1654 & pi067;
assign w18088 = ~w1661 & pi002;
assign w18089 = ~w1673 & ~w1674;
assign w18090 = ~w1689 & ~w1676;
assign w18091 = w1710 & pi026;
assign w18092 = w1724 & ~pi115;
assign w18093 = ~w1730 & ~pi030;
assign w18094 = w1738 & ~pi026;
assign w18095 = w1695 & w20164;
assign w18096 = (~w1770 & w8982) | (~w1770 & w20165) | (w8982 & w20165);
assign w18097 = ~w1764 & pi115;
assign w18098 = ~w1717 & ~pi115;
assign w18099 = w1808 & pi008;
assign w18100 = ~pi059 & ~pi056;
assign w18101 = ~w1819 & ~w1806;
assign w18102 = w1816 & pi026;
assign w18103 = w1845 & pi117;
assign w18104 = w1847 & ~pi002;
assign w18105 = ~w1860 & pi117;
assign w18106 = ~pi064 & ~pi117;
assign w18107 = w1867 & pi002;
assign w18108 = ~w1871 & w1874;
assign w18109 = w1861 & pi036;
assign w18110 = ~pi117 & pi105;
assign w18111 = w1884 & w9060;
assign w18112 = w1902 & pi117;
assign w18113 = ~w1878 & pi117;
assign w18114 = w1909 & ~w1904;
assign w18115 = ~w1924 & pi002;
assign w18116 = ~pi117 & pi061;
assign w18117 = w1927 & ~pi032;
assign w18118 = ~w1883 & w9280;
assign w18119 = w1937 & pi115;
assign w18120 = w1701 & ~pi115;
assign w18121 = w1939 & ~pi026;
assign w18122 = w1767 & pi026;
assign w18123 = w1950 & ~pi115;
assign w18124 = ~w1972 & ~w1948;
assign w18125 = ~w1975 & ~pi026;
assign w18126 = pi095 & pi115;
assign w18127 = ~w1992 & ~w1993;
assign w18128 = w1723 & pi115;
assign w18129 = w2009 & w20166;
assign w18130 = ~w2016 & ~pi026;
assign w18131 = ~w2026 & pi026;
assign w18132 = w2028 & w1996;
assign w18133 = pi099 & ~pi115;
assign w18134 = w2050 & ~pi092;
assign w18135 = w2055 & ~pi089;
assign w18136 = w2075 & w5823;
assign w18137 = (~w2076 & w2162) | (~w2076 & w20167) | (w2162 & w20167);
assign w18138 = ~pi087 & ~pi092;
assign w18139 = w2104 & ~w2090;
assign w18140 = w2107 & w18891;
assign w18141 = ~w2129 & ~pi089;
assign w18142 = ~w2118 & w18978;
assign w18143 = ~w2160 & ~pi089;
assign w18144 = w2143 & w20168;
assign w18145 = w2187 & ~pi046;
assign w18146 = ~w2194 & ~w2161;
assign w18147 = ~w2106 & ~pi053;
assign w18148 = ~w2200 & ~w2199;
assign w18149 = w1966 & ~pi115;
assign w18150 = w1744 & w1773;
assign w18151 = w2211 & ~pi026;
assign w18152 = w1700 & w8537;
assign w18153 = w2237 & ~pi026;
assign w18154 = ~w2234 & w20169;
assign w18155 = ~w2258 & ~pi026;
assign w18156 = w1706 & w20170;
assign w18157 = w2262 & w2260;
assign w18158 = ~w2282 & ~w2259;
assign w18159 = w2292 & ~pi080;
assign w18160 = w2313 & ~pi080;
assign w18161 = w2319 & pi073;
assign w18162 = w2297 & ~pi073;
assign w18163 = w2363 & w2368;
assign w18164 = ~pi042 & ~pi080;
assign w18165 = w2367 & w20171;
assign w18166 = ~w2366 & w20332;
assign w18167 = ~w2394 & ~w2397;
assign w18168 = ~w2401 & ~pi073;
assign w18169 = ~pi075 & ~pi110;
assign w18170 = w2295 & w20172;
assign w18171 = w2404 & w20173;
assign w18172 = ~w2427 & ~w2402;
assign w18173 = w2356 & ~pi015;
assign w18174 = ~w2430 & ~pi268;
assign w18175 = w2430 & pi268;
assign w18176 = ~w2454 & w20174;
assign w18177 = ~w2489 & pi003;
assign w18178 = pi016 & pi041;
assign w18179 = w2496 & pi120;
assign w18180 = pi074 & pi041;
assign w18181 = (pi003 & w2521) | (pi003 & w20175) | (w2521 & w20175);
assign w18182 = ~pi041 & pi120;
assign w18183 = w2540 & ~pi120;
assign w18184 = w2537 & ~pi003;
assign w18185 = w2554 & ~w2525;
assign w18186 = w2499 & w2566;
assign w18187 = w2572 & pi074;
assign w18188 = (pi003 & w2581) | (pi003 & w5996) | (w2581 & w5996);
assign w18189 = w2601 & w20176;
assign w18190 = ~pi118 & w2599;
assign w18191 = ~w2604 & ~w2610;
assign w18192 = w2629 & w2636;
assign w18193 = w2680 & ~pi118;
assign w18194 = w2689 & ~pi034;
assign w18195 = w2670 & pi034;
assign w18196 = w2716 & ~pi034;
assign w18197 = (pi118 & ~w2711) | (pi118 & w3181) | (~w2711 & w3181);
assign w18198 = w2733 & ~pi118;
assign w18199 = w2739 & w20177;
assign w18200 = (w2738 & w3181) | (w2738 & w20178) | (w3181 & w20178);
assign w18201 = w2495 & pi120;
assign w18202 = w2751 & ~pi003;
assign w18203 = w2501 & ~pi120;
assign w18204 = w2772 & pi003;
assign w18205 = pi041 & ~pi074;
assign w18206 = ~w2758 & ~w2761;
assign w18207 = w2791 & w20179;
assign w18208 = w2470 & ~pi120;
assign w18209 = w2816 & pi120;
assign w18210 = w2821 & ~pi045;
assign w18211 = pi045 & ~pi120;
assign w18212 = ~w2841 & pi003;
assign w18213 = ~w2810 & ~pi044;
assign w18214 = ~pi066 & ~pi101;
assign w18215 = w2850 & pi118;
assign w18216 = w2852 & ~pi034;
assign w18217 = w2877 & pi034;
assign w18218 = w2884 & ~w2861;
assign w18219 = ~w2890 & ~w2892;
assign w18220 = w2668 & pi118;
assign w18221 = (~pi034 & ~w2902) | (~pi034 & w2895) | (~w2902 & w2895);
assign w18222 = ~w2599 & ~pi118;
assign w18223 = ~w2920 & ~pi034;
assign w18224 = w2927 & pi062;
assign w18225 = ~pi034 & ~w2936;
assign w18226 = ~w2913 & ~pi038;
assign w18227 = w2951 & ~pi116;
assign w18228 = w2956 & ~pi058;
assign w18229 = pi057 & ~pi011;
assign w18230 = ~pi097 & pi116;
assign w18231 = pi000 & ~pi116;
assign w18232 = (pi058 & w2991) | (pi058 & w20180) | (w2991 & w20180);
assign w18233 = w3000 & w2965;
assign w18234 = ~w3010 & ~pi060;
assign w18235 = w2969 & w3090;
assign w18236 = ~w3030 & ~pi058;
assign w18237 = ~w3020 & w20181;
assign w18238 = ~w3063 & ~pi058;
assign w18239 = w3081 & w20182;
assign w18240 = w3090 & ~pi057;
assign w18241 = w3099 & ~w3064;
assign w18242 = ~w3104 & ~w3103;
assign w18243 = w2666 & ~pi118;
assign w18244 = w3117 & ~pi034;
assign w18245 = w2644 & w18645;
assign w18246 = ~w3150 & ~pi034;
assign w18247 = ~w3144 & w18647;
assign w18248 = ~w3170 & ~pi034;
assign w18249 = w2664 & w20183;
assign w18250 = ~w3171 & ~w3180;
assign w18251 = w3205 & ~pi090;
assign w18252 = ~pi051 & pi019;
assign w18253 = ~w3210 & ~w3217;
assign w18254 = w3226 & w3250;
assign w18255 = w3257 & pi090;
assign w18256 = w3264 & w3262;
assign w18257 = (w3232 & w3321) | (w3232 & w20184) | (w3321 & w20184);
assign w18258 = w3244 & w3226;
assign w18259 = w3274 & ~pi088;
assign w18260 = ~pi112 & ~pi090;
assign w18261 = w3208 & pi088;
assign w18262 = w3298 & w3295;
assign w18263 = ~w3319 & ~pi088;
assign w18264 = ~w3327 & w3321;
assign w18265 = w3287 & w20185;
assign w18266 = pi070 & ~pi122;
assign w18267 = ~w3393 & w3759;
assign w18268 = ~w3390 & pi122;
assign w18269 = ~w3412 & pi122;
assign w18270 = w3477 & pi043;
assign w18271 = (~w3442 & w20186) | (~w3442 & w20187) | (w20186 & w20187);
assign w18272 = w3430 & pi017;
assign w18273 = ~w3537 & pi024;
assign w18274 = w3522 & w18392;
assign w18275 = (~w3542 & w3862) | (~w3542 & w20188) | (w3862 & w20188);
assign w18276 = w3585 & pi024;
assign w18277 = ~pi094 & pi091;
assign w18278 = ~w3594 & w20189;
assign w18279 = ~pi094 & pi004;
assign w18280 = w3603 & ~pi091;
assign w18281 = ~w3592 & ~w3601;
assign w18282 = w3520 & pi094;
assign w18283 = w3621 & ~pi005;
assign w18284 = w3634 & pi005;
assign w18285 = ~w3653 & ~w3649;
assign w18286 = w3676 & ~pi039;
assign w18287 = ~w3693 & ~w3690;
assign w18288 = w3697 & w3696;
assign w18289 = (~w3673 & w20190) | (~w3673 & w20191) | (w20190 & w20191);
assign w18290 = w3708 & w3404;
assign w18291 = (w3710 & w3756) | (w3710 & w20919) | (w3756 & w20919);
assign w18292 = w3373 & ~pi122;
assign w18293 = (~w3718 & w20186) | (~w3718 & w20920) | (w20186 & w20920);
assign w18294 = w3714 & w3418;
assign w18295 = pi076 & ~pi077;
assign w18296 = pi084 & pi091;
assign w18297 = w3784 & pi091;
assign w18298 = w3786 & pi024;
assign w18299 = w3805 & w3801;
assign w18300 = ~w3806 & ~w3807;
assign w18301 = (~w3782 & w20192) | (~w3782 & w20193) | (w20192 & w20193);
assign w18302 = w3648 & w4383;
assign w18303 = w3830 & ~pi091;
assign w18304 = (w3813 & w3858) | (w3813 & w20921) | (w3858 & w20921);
assign w18305 = w3840 & w3568;
assign w18306 = w3822 & ~pi004;
assign w18307 = (~w3819 & w11392) | (~w3819 & w20922) | (w11392 & w20922);
assign w18308 = ~w3887 & pi039;
assign w18309 = w3403 & w20194;
assign w18310 = w3894 & pi122;
assign w18311 = w3931 & pi017;
assign w18312 = w3891 & pi043;
assign w18313 = w3935 & ~pi122;
assign w18314 = ~w3464 & pi039;
assign w18315 = w3969 & w4044;
assign w18316 = w4011 & ~pi106;
assign w18317 = pi035 & pi065;
assign w18318 = ~w4053 & ~pi065;
assign w18319 = w4054 & ~w4062;
assign w18320 = ~w4003 & ~pi068;
assign w18321 = w4104 & w4116;
assign w18322 = w4033 & pi035;
assign w18323 = ~w4119 & ~w4030;
assign w18324 = ~pi124 & pi113;
assign w18325 = w4133 & pi096;
assign w18326 = w4160 & pi113;
assign w18327 = pi125 & pi010;
assign w18328 = pi009 & pi096;
assign w18329 = w4228 & ~pi113;
assign w18330 = ~w4138 & pi096;
assign w18331 = w4254 & ~pi113;
assign w18332 = ~pi124 & pi009;
assign w18333 = ~w3481 & ~w4300;
assign w18334 = (~w4301 & w20195) | (~w4301 & w20196) | (w20195 & w20196);
assign w18335 = ~w4305 & ~pi039;
assign w18336 = ~w4315 & w3756;
assign w18337 = w3761 & w3464;
assign w18338 = w4312 & pi017;
assign w18339 = ~pi122 & w4350;
assign w18340 = w4335 & w20197;
assign w18341 = ~pi091 & ~w3587;
assign w18342 = ~w4365 & pi024;
assign w18343 = ~pi091 & ~w3788;
assign w18344 = w3550 & ~pi091;
assign w18345 = pi091 & ~w4380;
assign w18346 = pi084 & ~pi005;
assign w18347 = w4381 & ~pi024;
assign w18348 = w3807 & w4393;
assign w18349 = w4396 & w3566;
assign w18350 = w4390 & pi018;
assign w18351 = ~w4416 & ~w4399;
assign w18352 = ~w4410 & w3862;
assign w18353 = ~w4424 & w4425;
assign w18354 = w4037 & w4086;
assign w18355 = (~w4449 & w7900) | (~w4449 & w20198) | (w7900 & w20198);
assign w18356 = pi037 & pi035;
assign w18357 = ~w4470 & ~w4466;
assign w18358 = w4474 & w4032;
assign w18359 = ~w4465 & ~pi065;
assign w18360 = (~w4455 & w20199) | (~w4455 & w20200) | (w20199 & w20200);
assign w18361 = w4484 & w4047;
assign w18362 = (w4488 & w7900) | (w4488 & w20923) | (w7900 & w20923);
assign w18363 = w4090 & ~pi106;
assign w18364 = (~w4494 & w7198) | (~w4494 & w20924) | (w7198 & w20924);
assign w18365 = w4520 & w4098;
assign w18366 = ~w4522 & ~w4524;
assign w18367 = ~w4531 & ~w4535;
assign w18368 = w4126 & w20201;
assign w18369 = w4234 & w4135;
assign w18370 = ~w4581 & ~w4578;
assign w18371 = (~w4547 & w4726) | (~w4547 & w20202) | (w4726 & w20202);
assign w18372 = w4583 & pi113;
assign w18373 = w4139 & ~pi113;
assign w18374 = (pi010 & ~w4613) | (pi010 & w20203) | (~w4613 & w20203);
assign w18375 = w4618 & w4150;
assign w18376 = w4241 & ~pi055;
assign w18377 = ~w4620 & ~w4623;
assign w18378 = (~w4632 & ~w4194) | (~w4632 & w20204) | (~w4194 & w20204);
assign w18379 = (~w4554 & w20205) | (~w4554 & w20206) | (w20205 & w20206);
assign w18380 = ~w4676 & ~pi096;
assign w18381 = (pi113 & ~w4665) | (pi113 & w20207) | (~w4665 & w20207);
assign w18382 = w4188 & w4626;
assign w18383 = w4144 & w4632;
assign w18384 = w4178 & ~pi113;
assign w18385 = ~w4718 & ~w4719;
assign w18386 = w4729 & w4726;
assign w18387 = ~w4715 & pi010;
assign w18388 = (w4667 & w20208) | (w4667 & w20209) | (w20208 & w20209);
assign w18389 = ~w4748 & ~pi191;
assign w18390 = (~w4689 & w20210) | (~w4689 & w20211) | (w20210 & w20211);
assign w18391 = ~w4753 & ~w3531;
assign w18392 = ~pi091 & pi004;
assign w18393 = w3539 & pi024;
assign w18394 = ~w4762 & w3822;
assign w18395 = w4777 & ~w4766;
assign w18396 = w4787 & w3862;
assign w18397 = w4378 & w20212;
assign w18398 = w3570 & pi004;
assign w18399 = ~w4818 & pi024;
assign w18400 = w3547 & ~pi004;
assign w18401 = ~w4786 & w11392;
assign w18402 = w4834 & pi106;
assign w18403 = w4836 & ~pi065;
assign w18404 = ~pi031 & ~pi100;
assign w18405 = ~w4853 & pi106;
assign w18406 = w4451 & pi065;
assign w18407 = w4854 & pi068;
assign w18408 = w3979 & ~pi106;
assign w18409 = pi031 & pi065;
assign w18410 = ~w4871 & w4890;
assign w18411 = w4463 & pi106;
assign w18412 = w3988 & pi065;
assign w18413 = (~pi065 & ~w4877) | (~pi065 & w4526) | (~w4877 & w4526);
assign w18414 = w4922 & pi122;
assign w18415 = w4924 & ~pi039;
assign w18416 = w3472 & ~pi122;
assign w18417 = w3761 & pi039;
assign w18418 = w4945 & ~w4937;
assign w18419 = ~w4935 & w20213;
assign w18420 = w3911 & w3759;
assign w18421 = ~w3693 & ~w4957;
assign w18422 = w3480 & w3756;
assign w18423 = w3464 & pi076;
assign w18424 = w3405 & w20214;
assign w18425 = w4968 & ~pi039;
assign w18426 = w3697 & w3394;
assign w18427 = w4972 & pi039;
assign w18428 = w3685 & w3459;
assign w18429 = ~w4752 & ~pi529;
assign w18430 = w294 & w17925;
assign w18431 = (~w5001 & w1416) | (~w5001 & w20215) | (w1416 & w20215);
assign w18432 = ~pi111 & ~w1040;
assign w18433 = w1396 & w1431;
assign w18434 = ~w5015 & ~pi048;
assign w18435 = (~w5006 & w20216) | (~w5006 & w20217) | (w20216 & w20217);
assign w18436 = w281 & w18005;
assign w18437 = w347 & ~pi123;
assign w18438 = (w5026 & w1416) | (w5026 & w20925) | (w1416 & w20925);
assign w18439 = w5028 & w353;
assign w18440 = w383 & pi093;
assign w18441 = ~w5060 & ~w5061;
assign w18442 = w396 & w1426;
assign w18443 = (~w5032 & w20157) | (~w5032 & w20926) | (w20157 & w20926);
assign w18444 = w971 & w5109;
assign w18445 = (w5083 & w5136) | (w5083 & w20218) | (w5136 & w20218);
assign w18446 = w5095 & w476;
assign w18447 = ~w5096 & ~w1184;
assign w18448 = w445 & w20927;
assign w18449 = (w5100 & w5136) | (w5100 & w20928) | (w5136 & w20928);
assign w18450 = w488 & ~pi114;
assign w18451 = (~w5106 & w7344) | (~w5106 & w20929) | (w7344 & w20929);
assign w18452 = w5101 & w479;
assign w18453 = (~w5080 & w20220) | (~w5080 & w20221) | (w20220 & w20221);
assign w18454 = ~w5161 & w5163;
assign w18455 = w5174 & ~pi083;
assign w18456 = w5197 & ~w5199;
assign w18457 = pi083 & ~w5233;
assign w18458 = pi107 & ~pi083;
assign w18459 = ~w26 & ~pi078;
assign w18460 = w5221 & w5238;
assign w18461 = w5218 & pi014;
assign w18462 = ~w5242 & ~w5187;
assign w18463 = (~pi083 & ~w14) | (~pi083 & w84) | (~w14 & w84);
assign w18464 = w5263 & ~w13;
assign w18465 = w40 & ~pi083;
assign w18466 = (~pi040 & ~w5285) | (~pi040 & w20222) | (~w5285 & w20222);
assign w18467 = w1289 & w46;
assign w18468 = (~w5284 & w20134) | (~w5284 & w20223) | (w20134 & w20223);
assign w18469 = ~w5311 & ~pi040;
assign w18470 = w1229 & w383;
assign w18471 = w5339 & pi048;
assign w18472 = (~w5336 & w20224) | (~w5336 & w20225) | (w20224 & w20225);
assign w18473 = w5359 & ~pi048;
assign w18474 = ~w5379 & w5378;
assign w18475 = ~w5348 & w5391;
assign w18476 = (w744 & w20226) | (w744 & w20227) | (w20226 & w20227);
assign w18477 = (~w744 & w20228) | (~w744 & w20229) | (w20228 & w20229);
assign w18478 = ~w5402 & ~pi529;
assign w18479 = ~w510 & ~w934;
assign w18480 = ~w5423 & ~pi001;
assign w18481 = w1185 & pi001;
assign w18482 = w1152 & w536;
assign w18483 = w993 & ~pi013;
assign w18484 = ~w5444 & ~pi001;
assign w18485 = w415 & ~pi114;
assign w18486 = pi098 & pi114;
assign w18487 = ~w5467 & w5468;
assign w18488 = ~w5446 & w5479;
assign w18489 = ~w5489 & w17964;
assign w18490 = pi104 & w5499;
assign w18491 = w1444 & w604;
assign w18492 = ~w607 & pi012;
assign w18493 = w5515 & ~w574;
assign w18494 = w584 & ~pi104;
assign w18495 = ~w5537 & ~pi102;
assign w18496 = w708 & pi102;
assign w18497 = (w612 & w20230) | (w612 & w20231) | (w20230 & w20231);
assign w18498 = (~w612 & w20232) | (~w612 & w20233) | (w20232 & w20233);
assign w18499 = w5579 & pi083;
assign w18500 = w80 & ~pi083;
assign w18501 = w5581 & ~pi040;
assign w18502 = w56 & ~pi083;
assign w18503 = w1289 & pi040;
assign w18504 = ~pi083 & ~w5593;
assign w18505 = ~w174 & ~w5610;
assign w18506 = ~w79 & ~w5614;
assign w18507 = ~w26 & ~pi083;
assign w18508 = w160 & pi083;
assign w18509 = w5632 & pi040;
assign w18510 = (pi078 & ~w5599) | (pi078 & w20234) | (~w5599 & w20234);
assign w18511 = ~w5672 & ~pi529;
assign w18512 = w2395 & ~pi080;
assign w18513 = w5693 & ~pi075;
assign w18514 = w5694 & ~pi073;
assign w18515 = w2405 & w2421;
assign w18516 = w2377 & pi073;
assign w18517 = w2299 & w20235;
assign w18518 = ~pi110 & ~pi080;
assign w18519 = (~w5708 & w8800) | (~w5708 & w20236) | (w8800 & w20236);
assign w18520 = w5722 & pi080;
assign w18521 = w5746 & ~pi080;
assign w18522 = w5748 & ~pi073;
assign w18523 = w2330 & w2415;
assign w18524 = ~w5749 & ~w5752;
assign w18525 = (~w5686 & w20237) | (~w5686 & w20238) | (w20237 & w20238);
assign w18526 = ~w5778 & ~pi190;
assign w18527 = (~w5705 & w20239) | (~w5705 & w20240) | (w20239 & w20240);
assign w18528 = w5786 & pi092;
assign w18529 = pi050 & ~pi092;
assign w18530 = w5788 & ~pi089;
assign w18531 = w5802 & pi046;
assign w18532 = w5806 & pi089;
assign w18533 = w5816 & ~w5807;
assign w18534 = ~w5801 & w19355;
assign w18535 = ~pi087 & pi050;
assign w18536 = ~w5827 & ~w5828;
assign w18537 = w2059 & w20241;
assign w18538 = w5844 & pi092;
assign w18539 = ~w5846 & w5857;
assign w18540 = w5814 & pi092;
assign w18541 = pi092 & w2051;
assign w18542 = w5861 & pi089;
assign w18543 = (~w5826 & w20242) | (~w5826 & w20243) | (w20242 & w20243);
assign w18544 = ~w745 & ~pi136;
assign w18545 = (~w744 & w20244) | (~w744 & w20245) | (w20244 & w20245);
assign w18546 = ~w5924 & w20179;
assign w18547 = w2523 & w5938;
assign w18548 = ~w5940 & ~w5937;
assign w18549 = w2568 & w9858;
assign w18550 = (w5944 & w5996) | (w5944 & w20930) | (w5996 & w20930);
assign w18551 = w2477 & ~pi120;
assign w18552 = (~w5953 & w10300) | (~w5953 & w20931) | (w10300 & w20931);
assign w18553 = w5974 & w2467;
assign w18554 = w5955 & ~pi016;
assign w18555 = pi081 & pi120;
assign w18556 = ~w5987 & ~w5989;
assign w18557 = (~w5922 & w20246) | (~w5922 & w20247) | (w20246 & w20247);
assign w18558 = pi116 & ~w6012;
assign w18559 = w6007 & w20248;
assign w18560 = ~pi000 & pi116;
assign w18561 = w3035 & w3090;
assign w18562 = w6038 & ~w6014;
assign w18563 = w3034 & pi058;
assign w18564 = w3060 & ~pi116;
assign w18565 = w2963 & w20249;
assign w18566 = ~pi000 & ~pi057;
assign w18567 = (w6066 & w10156) | (w6066 & w20250) | (w10156 & w20250);
assign w18568 = w3177 & pi118;
assign w18569 = w2653 & w18645;
assign w18570 = (~w6108 & w2895) | (~w6108 & w20251) | (w2895 & w20251);
assign w18571 = w2615 & ~pi118;
assign w18572 = w3168 & w3191;
assign w18573 = w6103 & pi034;
assign w18574 = w2719 & w18645;
assign w18575 = (w6124 & w3181) | (w6124 & w20252) | (w3181 & w20252);
assign w18576 = w6132 & ~pi034;
assign w18577 = (~w6130 & w20253) | (~w6130 & w20254) | (w20253 & w20254);
assign w18578 = w6126 & w2643;
assign w18579 = w2648 & pi119;
assign w18580 = w6122 & pi038;
assign w18581 = w3081 & w20255;
assign w18582 = ~w6183 & ~pi116;
assign w18583 = pi000 & ~pi058;
assign w18584 = w6188 & w3090;
assign w18585 = w3041 & w20256;
assign w18586 = w2962 & w18231;
assign w18587 = (~w6207 & w10156) | (~w6207 & w20932) | (w10156 & w20932);
assign w18588 = (pi116 & ~w6205) | (pi116 & w20257) | (~w6205 & w20257);
assign w18589 = ~w2950 & ~pi116;
assign w18590 = w6238 & pi011;
assign w18591 = pi000 & ~pi057;
assign w18592 = w6244 & pi058;
assign w18593 = w3300 & pi088;
assign w18594 = w6283 & w20258;
assign w18595 = ~pi086 & pi090;
assign w18596 = w6288 & w20259;
assign w18597 = w6286 & ~pi006;
assign w18598 = pi049 & pi112;
assign w18599 = w6316 & pi090;
assign w18600 = w3206 & pi051;
assign w18601 = w6338 & ~pi019;
assign w18602 = ~w6344 & ~w3239;
assign w18603 = w6356 & w6357;
assign w18604 = ~pi090 & ~pi088;
assign w18605 = ~w6361 & ~w6346;
assign w18606 = (~w6315 & w20260) | (~w6315 & w20261) | (w20260 & w20261);
assign w18607 = w3323 & pi090;
assign w18608 = w6370 & pi088;
assign w18609 = w3317 & w6274;
assign w18610 = ~w6393 & ~w6394;
assign w18611 = w6395 & ~w6376;
assign w18612 = w3229 & w20262;
assign w18613 = (w6400 & w3295) | (w6400 & w20263) | (w3295 & w20263);
assign w18614 = w6417 & ~pi090;
assign w18615 = (~w6407 & w20264) | (~w6407 & w20265) | (w20264 & w20265);
assign w18616 = w6429 & w3250;
assign w18617 = ~w6440 & pi088;
assign w18618 = w3275 & w6442;
assign w18619 = w3211 & w3228;
assign w18620 = ~w6458 & w18604;
assign w18621 = w3288 & ~w6301;
assign w18622 = w3205 & w6287;
assign w18623 = ~w3229 & pi006;
assign w18624 = ~w6513 & ~pi088;
assign w18625 = w3285 & pi088;
assign w18626 = w6307 & pi090;
assign w18627 = (w6298 & w20266) | (w6298 & w20267) | (w20266 & w20267);
assign w18628 = (~w6298 & w20268) | (~w6298 & w20269) | (w20268 & w20269);
assign w18629 = w6552 & pi116;
assign w18630 = w3076 & ~pi116;
assign w18631 = w2951 & pi058;
assign w18632 = ~pi116 & ~w6563;
assign w18633 = w6245 & w20270;
assign w18634 = ~w6575 & ~w6576;
assign w18635 = w3090 & pi022;
assign w18636 = (~pi058 & ~w3004) | (~pi058 & w3083) | (~w3004 & w3083);
assign w18637 = ~w6604 & pi058;
assign w18638 = pi097 & ~pi116;
assign w18639 = pi058 & w6618;
assign w18640 = (~w6558 & w20271) | (~w6558 & w20272) | (w20271 & w20272);
assign w18641 = w2613 & ~pi118;
assign w18642 = ~w2676 & ~pi038;
assign w18643 = ~w6655 & w6656;
assign w18644 = w6646 & w20273;
assign w18645 = ~pi103 & pi118;
assign w18646 = ~w6151 & w20274;
assign w18647 = pi034 & pi038;
assign w18648 = w6647 & pi066;
assign w18649 = ~pi034 & ~w6707;
assign w18650 = w3071 & w6015;
assign w18651 = ~w2965 & pi058;
assign w18652 = w6718 & w6722;
assign w18653 = w3060 & w20275;
assign w18654 = w3040 & ~pi116;
assign w18655 = ~pi011 & ~pi058;
assign w18656 = ~w6740 & w6742;
assign w18657 = ~w3060 & pi058;
assign w18658 = w3094 & w3076;
assign w18659 = pi116 & ~w6777;
assign w18660 = ~w3031 & ~pi060;
assign w18661 = w6764 & w6782;
assign w18662 = w6460 & pi088;
assign w18663 = ~pi090 & pi086;
assign w18664 = pi088 & pi006;
assign w18665 = w6420 & pi090;
assign w18666 = pi051 & ~pi006;
assign w18667 = w3203 & ~pi090;
assign w18668 = ~w6331 & w6382;
assign w18669 = w6802 & ~pi090;
assign w18670 = ~pi049 & pi088;
assign w18671 = w6849 & w6865;
assign w18672 = w6801 & pi090;
assign w18673 = w6886 & ~pi088;
assign w18674 = ~w6892 & ~w6896;
assign w18675 = w6808 & w18604;
assign w18676 = ~w6913 & w20264;
assign w18677 = ~w6930 & pi088;
assign w18678 = pi051 & ~pi090;
assign w18679 = w6934 & w6944;
assign w18680 = ~w6951 & ~pi529;
assign w18681 = ~pi025 & ~pi009;
assign w18682 = w6969 & pi113;
assign w18683 = w6971 & ~pi096;
assign w18684 = w4131 & pi096;
assign w18685 = w6978 & ~pi113;
assign w18686 = ~pi125 & ~pi055;
assign w18687 = ~w6977 & ~w6983;
assign w18688 = w4156 & ~w4555;
assign w18689 = w4195 & w20276;
assign w18690 = w4262 & w4726;
assign w18691 = w7012 & pi010;
assign w18692 = w4560 & pi113;
assign w18693 = ~w4236 & pi113;
assign w18694 = w7018 & ~w7014;
assign w18695 = w7024 & ~w7023;
assign w18696 = w7028 & w20277;
assign w18697 = ~w7037 & ~pi529;
assign w18698 = ~pi125 & pi096;
assign w18699 = ~pi025 & ~pi010;
assign w18700 = (~pi096 & ~w7060) | (~pi096 & w20278) | (~w7060 & w20278);
assign w18701 = w7080 & ~w4692;
assign w18702 = w4183 & ~pi113;
assign w18703 = ~w4137 & ~pi113;
assign w18704 = w7103 & ~w4254;
assign w18705 = w4213 & w20279;
assign w18706 = (w7108 & w20276) | (w7108 & w20280) | (w20276 & w20280);
assign w18707 = w4574 & pi113;
assign w18708 = w4837 & ~pi106;
assign w18709 = w4019 & w20281;
assign w18710 = w3977 & w4838;
assign w18711 = w4498 & w3973;
assign w18712 = (~w4862 & w20282) | (~w4862 & w20283) | (w20282 & w20283);
assign w18713 = ~w7159 & pi106;
assign w18714 = w4088 & w20284;
assign w18715 = w4041 & ~pi106;
assign w18716 = ~pi031 & ~pi128;
assign w18717 = w7173 & w4015;
assign w18718 = w7175 & ~pi068;
assign w18719 = w4106 & pi128;
assign w18720 = w7194 & w7198;
assign w18721 = ~w7201 & ~w7202;
assign w18722 = ~w7217 & ~w7177;
assign w18723 = ~w7144 & ~pi529;
assign w18724 = ~w294 & pi027;
assign w18725 = w7242 & pi123;
assign w18726 = ~w7258 & w7261;
assign w18727 = ~pi023 & ~pi048;
assign w18728 = w301 & ~w329;
assign w18729 = w285 & w318;
assign w18730 = w7273 & w1420;
assign w18731 = ~w7281 & pi020;
assign w18732 = w275 & w386;
assign w18733 = w5027 & w20285;
assign w18734 = w288 & w5058;
assign w18735 = ~w7262 & ~pi020;
assign w18736 = w7313 & w7311;
assign w18737 = w415 & w436;
assign w18738 = (~pi001 & w5118) | (~pi001 & w20286) | (w5118 & w20286);
assign w18739 = w7326 & ~pi114;
assign w18740 = w973 & pi114;
assign w18741 = w426 & w7311;
assign w18742 = w5074 & ~pi114;
assign w18743 = ~pi054 & ~w467;
assign w18744 = (~w7305 & w20220) | (~w7305 & w20287) | (w20220 & w20287);
assign w18745 = ~w7384 & w123;
assign w18746 = ~w7391 & ~w7403;
assign w18747 = ~w0 & pi040;
assign w18748 = w7415 & ~w7416;
assign w18749 = ~w22 & ~w166;
assign w18750 = w40 & w1348;
assign w18751 = w7430 & ~pi040;
assign w18752 = ~w7424 & w20288;
assign w18753 = w7470 & pi012;
assign w18754 = w7495 & ~pi102;
assign w18755 = ~w590 & ~w712;
assign w18756 = w812 & pi104;
assign w18757 = ~w7492 & w20289;
assign w18758 = ~w7517 & pi123;
assign w18759 = w5331 & ~pi123;
assign w18760 = ~pi123 & ~w312;
assign w18761 = ~w285 & pi048;
assign w18762 = w7541 & ~w7543;
assign w18763 = w379 & w314;
assign w18764 = ~w7558 & w20290;
assign w18765 = w1078 & pi048;
assign w18766 = w287 & w20291;
assign w18767 = w394 & pi048;
assign w18768 = ~w7252 & ~w7571;
assign w18769 = pi048 & w7572;
assign w18770 = ~w7382 & ~pi529;
assign w18771 = w572 & w689;
assign w18772 = w7600 & ~w7596;
assign w18773 = w598 & w639;
assign w18774 = ~w7614 & w7616;
assign w18775 = ~w594 & ~pi102;
assign w18776 = w880 & ~w7500;
assign w18777 = w584 & w703;
assign w18778 = w7453 & w7636;
assign w18779 = w580 & w20292;
assign w18780 = w5501 & w571;
assign w18781 = w608 & ~w585;
assign w18782 = w654 & w20293;
assign w18783 = ~w7619 & ~pi179;
assign w18784 = ~w7618 & w20294;
assign w18785 = ~w7661 & ~pi529;
assign w18786 = pi094 & pi091;
assign w18787 = pi094 & pi005;
assign w18788 = pi091 & ~w7707;
assign w18789 = ~w3777 & pi024;
assign w18790 = pi091 & ~w3830;
assign w18791 = w7730 & ~pi091;
assign w18792 = ~pi005 & pi024;
assign w18793 = ~w7734 & w7735;
assign w18794 = w7711 & pi005;
assign w18795 = w3761 & ~pi122;
assign w18796 = w3409 & w3418;
assign w18797 = w3474 & w3721;
assign w18798 = w7795 & ~w3684;
assign w18799 = w7778 & ~pi039;
assign w18800 = w3692 & w20295;
assign w18801 = w7808 & ~pi039;
assign w18802 = ~w7803 & w20190;
assign w18803 = ~w7822 & ~pi039;
assign w18804 = w3444 & w3692;
assign w18805 = w7825 & w7824;
assign w18806 = ~w7841 & ~w7823;
assign w18807 = w7799 & ~pi017;
assign w18808 = w4530 & ~pi106;
assign w18809 = w7852 & ~pi106;
assign w18810 = w7855 & pi065;
assign w18811 = w7847 & ~pi065;
assign w18812 = w3989 & w4032;
assign w18813 = w4474 & w20296;
assign w18814 = ~w7876 & w20199;
assign w18815 = ~w7894 & ~pi065;
assign w18816 = ~w7897 & w20297;
assign w18817 = w3994 & w20933;
assign w18818 = w7872 & ~pi068;
assign w18819 = pi125 & ~pi113;
assign w18820 = (pi096 & w7928) | (pi096 & w20298) | (w7928 & w20298);
assign w18821 = w4627 & ~pi113;
assign w18822 = w4663 & w4188;
assign w18823 = w7936 & ~pi096;
assign w18824 = (w7927 & w20299) | (w7927 & w20300) | (w20299 & w20300);
assign w18825 = w7096 & ~w4729;
assign w18826 = w4234 & w20301;
assign w18827 = w7950 & ~pi010;
assign w18828 = ~w7969 & ~pi096;
assign w18829 = w4163 & w20302;
assign w18830 = w7978 & w4738;
assign w18831 = (w7945 & w20303) | (w7945 & w20304) | (w20303 & w20304);
assign w18832 = (~w7945 & w20305) | (~w7945 & w20306) | (w20305 & w20306);
assign w18833 = w8011 & ~pi083;
assign w18834 = w69 & pi083;
assign w18835 = w8 & pi082;
assign w18836 = w7385 & w1348;
assign w18837 = w50 & w204;
assign w18838 = ~w8039 & w234;
assign w18839 = w173 & w9;
assign w18840 = ~w8061 & ~w81;
assign w18841 = w56 & w88;
assign w18842 = ~w8063 & w8069;
assign w18843 = w8071 & w20307;
assign w18844 = (pi142 & ~w8071) | (pi142 & w20308) | (~w8071 & w20308);
assign w18845 = ~w8080 & ~pi529;
assign w18846 = w1152 & ~w5109;
assign w18847 = w469 & w20309;
assign w18848 = w445 & w5109;
assign w18849 = w1013 & pi001;
assign w18850 = w7312 & w7311;
assign w18851 = w8104 & ~w8092;
assign w18852 = (~pi029 & ~w8096) | (~pi029 & w20310) | (~w8096 & w20310);
assign w18853 = w542 & w5136;
assign w18854 = w989 & pi001;
assign w18855 = ~w1154 & ~w942;
assign w18856 = w5101 & w20311;
assign w18857 = ~w927 & ~w917;
assign w18858 = ~w8131 & w7311;
assign w18859 = w425 & w446;
assign w18860 = w1163 & w8142;
assign w18861 = ~w5470 & w20312;
assign w18862 = ~w1526 & ~pi173;
assign w18863 = w1526 & pi173;
assign w18864 = w8156 & ~pi529;
assign w18865 = ~w4058 & ~w4087;
assign w18866 = ~w4851 & ~w4087;
assign w18867 = ~w8189 & ~w8191;
assign w18868 = w3989 & w4053;
assign w18869 = (~w8195 & w7896) | (~w8195 & w20313) | (w7896 & w20313);
assign w18870 = ~pi106 & ~w4056;
assign w18871 = (~w8207 & w4529) | (~w8207 & w20314) | (w4529 & w20314);
assign w18872 = ~w8217 & w8218;
assign w18873 = w566 & ~pi104;
assign w18874 = w8285 & ~pi102;
assign w18875 = ~w8291 & pi104;
assign w18876 = w614 & ~pi104;
assign w18877 = w1444 & pi102;
assign w18878 = w8299 & ~w8294;
assign w18879 = w8292 & pi012;
assign w18880 = w618 & ~pi104;
assign w18881 = w713 & pi104;
assign w18882 = ~w8330 & pi102;
assign w18883 = (w8303 & w20315) | (w8303 & w20316) | (w20315 & w20316);
assign w18884 = ~w8302 & ~pi164;
assign w18885 = (~w8301 & w20317) | (~w8301 & w20318) | (w20317 & w20318);
assign w18886 = ~w8344 & ~pi529;
assign w18887 = (w8301 & w20319) | (w8301 & w20320) | (w20319 & w20320);
assign w18888 = (~w8301 & w20321) | (~w8301 & w20322) | (w20321 & w20322);
assign w18889 = ~w8358 & ~pi529;
assign w18890 = (pi089 & w2144) | (pi089 & w19046) | (w2144 & w19046);
assign w18891 = ~pi087 & pi092;
assign w18892 = w8390 & ~pi089;
assign w18893 = w2052 & pi087;
assign w18894 = (~w8381 & w20323) | (~w8381 & w20324) | (w20323 & w20324);
assign w18895 = w8403 & ~pi089;
assign w18896 = w8417 & ~w8418;
assign w18897 = w8422 & pi092;
assign w18898 = ~w2108 & pi053;
assign w18899 = w2187 & w8438;
assign w18900 = w8440 & pi028;
assign w18901 = ~w8443 & ~w2086;
assign w18902 = ~w8445 & ~w8447;
assign w18903 = w2048 & w20325;
assign w18904 = (~w8457 & w2172) | (~w8457 & w20326) | (w2172 & w20326);
assign w18905 = w5864 & pi092;
assign w18906 = w8466 & ~pi089;
assign w18907 = ~w5827 & ~w8474;
assign w18908 = w8479 & pi092;
assign w18909 = ~w8483 & pi053;
assign w18910 = w2121 & w19043;
assign w18911 = (w8487 & w2172) | (w8487 & w20327) | (w2172 & w20327);
assign w18912 = w8501 & ~pi092;
assign w18913 = (~w8493 & w20242) | (~w8493 & w20328) | (w20242 & w20328);
assign w18914 = w8516 & w5823;
assign w18915 = ~w8518 & ~w8519;
assign w18916 = ~pi056 & pi008;
assign w18917 = pi099 & pi008;
assign w18918 = pi115 & ~w8558;
assign w18919 = w8545 & w8562;
assign w18920 = ~w1723 & pi026;
assign w18921 = w1976 & ~w8575;
assign w18922 = w8588 & pi030;
assign w18923 = w1718 & w1734;
assign w18924 = w1788 & w2265;
assign w18925 = w8538 & pi008;
assign w18926 = w8608 & w8614;
assign w18927 = ~w8668 & ~w8667;
assign w18928 = w8674 & ~pi002;
assign w18929 = w8702 & ~pi117;
assign w18930 = w8684 & pi067;
assign w18931 = w2346 & w20329;
assign w18932 = ~pi110 & pi080;
assign w18933 = w2367 & w8750;
assign w18934 = ~w8752 & ~w8753;
assign w18935 = (~w8724 & w2409) | (~w8724 & w20330) | (w2409 & w20330);
assign w18936 = w8757 & pi080;
assign w18937 = w8774 & ~pi080;
assign w18938 = w8759 & pi073;
assign w18939 = w8786 & pi080;
assign w18940 = w8788 & w2345;
assign w18941 = ~pi080 & ~pi075;
assign w18942 = w8732 & w20331;
assign w18943 = w8784 & ~pi015;
assign w18944 = (~w8730 & w20332) | (~w8730 & w20333) | (w20332 & w20333);
assign w18945 = w5716 & pi071;
assign w18946 = w8815 & pi080;
assign w18947 = w8829 & ~pi080;
assign w18948 = pi042 & pi073;
assign w18949 = ~w8820 & ~w8816;
assign w18950 = pi080 & ~w8864;
assign w18951 = w8866 & ~pi079;
assign w18952 = ~w8883 & w8880;
assign w18953 = ~w8843 & ~pi301;
assign w18954 = w8843 & pi301;
assign w18955 = w8722 & ~pi529;
assign w18956 = w2262 & pi115;
assign w18957 = ~w1992 & ~w8932;
assign w18958 = w2236 & w8537;
assign w18959 = w8926 & pi026;
assign w18960 = w1804 & w1771;
assign w18961 = w1715 & pi008;
assign w18962 = w8959 & ~w8954;
assign w18963 = w8547 & ~pi115;
assign w18964 = (~pi030 & ~w8968) | (~pi030 & w20334) | (~w8968 & w20334);
assign w18965 = w8947 & w1984;
assign w18966 = w8685 & pi117;
assign w18967 = w9002 & pi002;
assign w18968 = w1609 & w18110;
assign w18969 = w8688 & w8682;
assign w18970 = (~w8999 & w20336) | (~w8999 & w20337) | (w20336 & w20337);
assign w18971 = (pi002 & w1658) | (pi002 & w20934) | (w1658 & w20934);
assign w18972 = w8667 & ~pi117;
assign w18973 = (~w9026 & w9280) | (~w9026 & w20935) | (w9280 & w20935);
assign w18974 = w9045 & w1639;
assign w18975 = w9047 & pi002;
assign w18976 = pi046 & pi092;
assign w18977 = pi092 & ~w9076;
assign w18978 = pi089 & pi053;
assign w18979 = pi087 & pi092;
assign w18980 = ~w9109 & ~pi089;
assign w18981 = pi092 & ~w9113;
assign w18982 = ~w5848 & ~pi053;
assign w18983 = w2140 & w20338;
assign w18984 = w9134 & ~pi092;
assign w18985 = pi085 & pi089;
assign w18986 = ~w9139 & w9140;
assign w18987 = ~w5848 & ~pi089;
assign w18988 = w9106 & pi028;
assign w18989 = ~w8843 & ~pi184;
assign w18990 = w8843 & pi184;
assign w18991 = w9167 & ~pi115;
assign w18992 = w1759 & pi115;
assign w18993 = ~w9186 & pi115;
assign w18994 = w8573 & ~pi115;
assign w18995 = ~w9187 & w9191;
assign w18996 = ~w1736 & ~pi026;
assign w18997 = pi056 & pi026;
assign w18998 = w9201 & ~w1943;
assign w18999 = ~w2200 & ~w2000;
assign w19000 = w1720 & w1734;
assign w19001 = (~pi115 & w2001) | (~pi115 & w20339) | (w2001 & w20339);
assign w19002 = w9228 & pi026;
assign w19003 = (~pi002 & w9035) | (~pi002 & w20340) | (w9035 & w20340);
assign w19004 = w9246 & w9244;
assign w19005 = w1569 & w8631;
assign w19006 = (~w9239 & w20341) | (~w9239 & w20342) | (w20341 & w20342);
assign w19007 = w1607 & pi117;
assign w19008 = w8634 & w9244;
assign w19009 = ~w9268 & w9280;
assign w19010 = ~w9283 & ~w1545;
assign w19011 = w9018 & w1915;
assign w19012 = w2157 & ~w2085;
assign w19013 = w8421 & ~pi092;
assign w19014 = ~w9323 & ~w9321;
assign w19015 = w2099 & pi092;
assign w19016 = ~w9112 & w2177;
assign w19017 = w2060 & pi046;
assign w19018 = w5855 & w2162;
assign w19019 = w2138 & w20343;
assign w19020 = ~w9370 & ~w9354;
assign w19021 = w5810 & w2060;
assign w19022 = ~w9379 & ~w2143;
assign w19023 = w2060 & pi085;
assign w19024 = w9384 & pi089;
assign w19025 = w9391 & w20344;
assign w19026 = (pi178 & ~w9391) | (pi178 & w20345) | (~w9391 & w20345);
assign w19027 = w9399 & ~pi529;
assign w19028 = w1868 & ~w1927;
assign w19029 = w8693 & w20346;
assign w19030 = w1580 & w1927;
assign w19031 = w9421 & w9244;
assign w19032 = w1674 & pi002;
assign w19033 = ~w9426 & ~w9410;
assign w19034 = w1548 & w8682;
assign w19035 = w9436 & ~pi002;
assign w19036 = ~w9432 & w20347;
assign w19037 = ~w9450 & ~pi002;
assign w19038 = w1659 & w20348;
assign w19039 = w1545 & w20349;
assign w19040 = w8455 & ~pi281;
assign w19041 = ~w8455 & pi281;
assign w19042 = w9498 & ~pi089;
assign w19043 = ~pi085 & pi092;
assign w19044 = w2050 & w2187;
assign w19045 = ~w9508 & w18978;
assign w19046 = w2133 & pi089;
assign w19047 = w2075 & w2111;
assign w19048 = ~w8479 & ~w8433;
assign w19049 = ~w9529 & w8526;
assign w19050 = w8474 & pi092;
assign w19051 = ~w9528 & ~w9514;
assign w19052 = w2383 & ~w5706;
assign w19053 = w5753 & w2421;
assign w19054 = pi071 & pi015;
assign w19055 = (~pi073 & ~w9563) | (~pi073 & w20350) | (~w9563 & w20350);
assign w19056 = ~pi080 & ~w2305;
assign w19057 = w2347 & pi080;
assign w19058 = w2333 & ~pi080;
assign w19059 = w2347 & w2290;
assign w19060 = ~w9595 & w20351;
assign w19061 = w2316 & pi079;
assign w19062 = w5748 & pi080;
assign w19063 = w9610 & ~w9601;
assign w19064 = ~w9557 & ~pi529;
assign w19065 = w9633 & pi080;
assign w19066 = w9635 & ~pi073;
assign w19067 = ~w9645 & ~pi080;
assign w19068 = w2359 & pi073;
assign w19069 = ~w9655 & pi015;
assign w19070 = w8737 & pi080;
assign w19071 = w2421 & pi075;
assign w19072 = w9663 & ~w9658;
assign w19073 = w2337 & pi080;
assign w19074 = w5716 & w20352;
assign w19075 = ~w9666 & w9699;
assign w19076 = ~w9657 & ~pi162;
assign w19077 = w9657 & pi162;
assign w19078 = ~w9704 & ~pi529;
assign w19079 = ~w2314 & pi079;
assign w19080 = w2303 & w20353;
assign w19081 = ~w9736 & w9742;
assign w19082 = ~w2321 & ~pi073;
assign w19083 = w9756 & w2403;
assign w19084 = w2333 & w18941;
assign w19085 = ~w9759 & ~w9758;
assign w19086 = ~w9764 & pi015;
assign w19087 = w5753 & w8847;
assign w19088 = ~w9770 & w9772;
assign w19089 = w2405 & ~w2337;
assign w19090 = w2300 & w20354;
assign w19091 = ~w9743 & ~pi015;
assign w19092 = w9789 & ~pi529;
assign w19093 = ~w9657 & ~pi192;
assign w19094 = w9657 & pi192;
assign w19095 = ~w9800 & ~pi529;
assign w19096 = w2772 & ~pi120;
assign w19097 = w5917 & w5996;
assign w19098 = w2584 & pi003;
assign w19099 = w2449 & w2828;
assign w19100 = w9835 & w9832;
assign w19101 = w9842 & ~w9823;
assign w19102 = w2565 & pi003;
assign w19103 = w9847 & w5996;
assign w19104 = ~w2524 & ~w2776;
assign w19105 = w5950 & w20355;
assign w19106 = ~w9872 & ~pi003;
assign w19107 = w2541 & w5996;
assign w19108 = w2811 & w9832;
assign w19109 = ~w9873 & ~w9875;
assign w19110 = ~w6264 & ~pi278;
assign w19111 = w6264 & pi278;
assign w19112 = w2520 & w2467;
assign w19113 = w9957 & pi120;
assign w19114 = w9960 & ~w9943;
assign w19115 = ~w9876 & w9989;
assign w19116 = w9945 & pi074;
assign w19117 = w10002 & ~pi120;
assign w19118 = ~w2448 & pi003;
assign w19119 = ~w9996 & w10010;
assign w19120 = w10018 & ~pi118;
assign w19121 = ~w10020 & ~w2723;
assign w19122 = w2612 & w2719;
assign w19123 = ~w10032 & w10044;
assign w19124 = ~w2713 & ~pi034;
assign w19125 = w10059 & w3172;
assign w19126 = w2653 & w20356;
assign w19127 = ~w10062 & ~w10061;
assign w19128 = ~w10069 & pi038;
assign w19129 = w2676 & w3181;
assign w19130 = ~w10079 & ~w10082;
assign w19131 = w3174 & w10084;
assign w19132 = w2673 & w20357;
assign w19133 = w10093 & ~pi116;
assign w19134 = ~w10096 & ~w6240;
assign w19135 = w2958 & w3023;
assign w19136 = ~w3071 & ~pi060;
assign w19137 = w2966 & ~w2965;
assign w19138 = w10127 & ~pi058;
assign w19139 = w3066 & w3041;
assign w19140 = w10115 & w3065;
assign w19141 = w10146 & ~w10129;
assign w19142 = ~w10157 & ~w3081;
assign w19143 = w3076 & w3075;
assign w19144 = ~w10159 & ~w10160;
assign w19145 = w6941 & ~pi090;
assign w19146 = ~w10176 & ~w6351;
assign w19147 = w10194 & pi090;
assign w19148 = ~w10195 & w10200;
assign w19149 = ~pi112 & ~pi088;
assign w19150 = w3264 & w18663;
assign w19151 = w6432 & w3321;
assign w19152 = w3216 & w6817;
assign w19153 = w3246 & w3295;
assign w19154 = ~w3261 & ~w10238;
assign w19155 = w3324 & w10240;
assign w19156 = (~pi141 & w10203) | (~pi141 & w20358) | (w10203 & w20358);
assign w19157 = ~w10203 & w20359;
assign w19158 = ~w10017 & ~pi529;
assign w19159 = w2455 & w9850;
assign w19160 = w10270 & w9832;
assign w19161 = w2775 & w20360;
assign w19162 = w10280 & ~pi120;
assign w19163 = w2796 & w2821;
assign w19164 = ~w10282 & ~w10283;
assign w19165 = w10293 & pi003;
assign w19166 = ~w10322 & ~w2520;
assign w19167 = (~w10264 & w20361) | (~w10264 & w20362) | (w20361 & w20362);
assign w19168 = pi101 & pi118;
assign w19169 = ~w2643 & pi034;
assign w19170 = w10337 & w10345;
assign w19171 = ~w10349 & w20363;
assign w19172 = ~w2660 & pi034;
assign w19173 = w2855 & w6662;
assign w19174 = ~w10379 & ~pi034;
assign w19175 = pi103 & ~w2680;
assign w19176 = w2668 & w3172;
assign w19177 = (~pi038 & w10370) | (~pi038 & w20364) | (w10370 & w20364);
assign w19178 = (pi003 & w2763) | (pi003 & w20936) | (w2763 & w20936);
assign w19179 = pi120 & ~w5954;
assign w19180 = ~w2477 & ~w2547;
assign w19181 = pi045 & pi003;
assign w19182 = ~w10433 & w20365;
assign w19183 = w2524 & ~pi120;
assign w19184 = w10436 & ~pi003;
assign w19185 = w2478 & w9832;
assign w19186 = ~w10476 & pi116;
assign w19187 = pi116 & pi060;
assign w19188 = ~w10117 & w10156;
assign w19189 = ~w10483 & w18655;
assign w19190 = ~w2965 & ~pi060;
assign w19191 = (w10486 & w20366) | (w10486 & w20367) | (w20366 & w20367);
assign w19192 = ~pi116 & ~w6058;
assign w19193 = w10516 & ~pi058;
assign w19194 = w10504 & w10525;
assign w19195 = ~w3177 & ~w6165;
assign w19196 = ~w10562 & ~pi034;
assign w19197 = w3139 & w2648;
assign w19198 = w10563 & pi038;
assign w19199 = ~w10586 & w10587;
assign w19200 = ~w10588 & w10595;
assign w19201 = w6187 & pi116;
assign w19202 = ~w6575 & ~w6211;
assign w19203 = w10094 & w3094;
assign w19204 = w10614 & pi058;
assign w19205 = (~w10612 & w20271) | (~w10612 & w20369) | (w20271 & w20369);
assign w19206 = w3023 & w18560;
assign w19207 = (w10163 & w3075) | (w10163 & w20937) | (w3075 & w20937);
assign w19208 = w6769 & ~pi116;
assign w19209 = (~w10630 & w20720) | (~w10630 & w20938) | (w20720 & w20938);
assign w19210 = w10100 & w6015;
assign w19211 = w10648 & pi116;
assign w19212 = w3095 & w20370;
assign w19213 = ~w10654 & w10658;
assign w19214 = ~w10683 & ~pi529;
assign w19215 = w2743 & ~pi161;
assign w19216 = ~w2743 & pi161;
assign w19217 = ~w10459 & ~pi529;
assign w19218 = w4508 & ~pi106;
assign w19219 = w4833 & pi106;
assign w19220 = ~w4059 & ~pi065;
assign w19221 = w4043 & ~w4842;
assign w19222 = w10734 & w7896;
assign w19223 = w4044 & w20371;
assign w19224 = ~w10750 & ~w10749;
assign w19225 = ~w10755 & pi068;
assign w19226 = w3996 & w10759;
assign w19227 = w4486 & w7900;
assign w19228 = ~w8201 & ~w10764;
assign w19229 = w7173 & w10766;
assign w19230 = w4000 & w20372;
assign w19231 = ~w10720 & w7198;
assign w19232 = ~w3418 & pi039;
assign w19233 = ~w10794 & w20373;
assign w19234 = pi109 & ~pi122;
assign w19235 = ~pi109 & w7824;
assign w19236 = w10832 & ~w10830;
assign w19237 = ~w10803 & w20374;
assign w19238 = (pi024 & w4768) | (pi024 & w20939) | (w4768 & w20939);
assign w19239 = ~w3830 & ~w3610;
assign w19240 = ~w10843 & ~w10850;
assign w19241 = ~w3586 & pi024;
assign w19242 = w10870 & ~w10871;
assign w19243 = w4395 & ~pi091;
assign w19244 = w3530 & pi091;
assign w19245 = w3550 & w10858;
assign w19246 = w3778 & w3858;
assign w19247 = w10892 & ~pi024;
assign w19248 = ~w10886 & w20375;
assign w19249 = w10915 & ~pi113;
assign w19250 = ~w10917 & ~w4732;
assign w19251 = w10931 & pi113;
assign w19252 = w4180 & ~w6972;
assign w19253 = w10934 & w4738;
assign w19254 = w4183 & w20376;
assign w19255 = ~w10960 & ~w10959;
assign w19256 = ~w10965 & ~pi010;
assign w19257 = w4586 & w4136;
assign w19258 = w4197 & w4726;
assign w19259 = ~w7085 & ~w10978;
assign w19260 = ~w10984 & pi113;
assign w19261 = (~pi096 & w7113) | (~pi096 & w20377) | (w7113 & w20377);
assign w19262 = w4183 & w4738;
assign w19263 = w11029 & ~pi096;
assign w19264 = ~w11022 & w20378;
assign w19265 = w11060 & ~pi122;
assign w19266 = w3385 & pi122;
assign w19267 = ~w11079 & pi122;
assign w19268 = pi043 & pi039;
assign w19269 = ~w11098 & w11099;
assign w19270 = w3474 & w18266;
assign w19271 = ~w11110 & ~w11102;
assign w19272 = ~w11111 & pi017;
assign w19273 = w3443 & w3435;
assign w19274 = w3449 & w3756;
assign w19275 = ~w11152 & pi106;
assign w19276 = pi106 & pi068;
assign w19277 = (~pi065 & w8211) | (~pi065 & w20379) | (w8211 & w20379);
assign w19278 = pi128 & ~pi106;
assign w19279 = ~w11160 & ~w11161;
assign w19280 = w4000 & w20380;
assign w19281 = ~w4021 & ~pi068;
assign w19282 = (w11177 & w11165) | (w11177 & w20381) | (w11165 & w20381);
assign w19283 = (~pi106 & ~w4097) | (~pi106 & w20940) | (~w4097 & w20940);
assign w19284 = w7194 & ~pi106;
assign w19285 = w11184 & ~pi065;
assign w19286 = w11178 & w11194;
assign w19287 = w10867 & w3858;
assign w19288 = w11216 & w10858;
assign w19289 = w3789 & w3652;
assign w19290 = w3609 & w3547;
assign w19291 = w3649 & pi024;
assign w19292 = w11230 & ~w11213;
assign w19293 = w7744 & w3858;
assign w19294 = w3625 & pi024;
assign w19295 = w3783 & w20189;
assign w19296 = ~w4774 & ~w4396;
assign w19297 = ~w11255 & ~pi024;
assign w19298 = w3531 & w20382;
assign w19299 = w11271 & ~w11256;
assign w19300 = (w7945 & w20383) | (w7945 & w20384) | (w20383 & w20384);
assign w19301 = (~w7945 & w20385) | (~w7945 & w20386) | (w20385 & w20386);
assign w19302 = (w4689 & w20387) | (w4689 & w20388) | (w20387 & w20388);
assign w19303 = (~w4689 & w20389) | (~w4689 & w20390) | (w20389 & w20390);
assign w19304 = w11331 & ~pi529;
assign w19305 = w3570 & w3773;
assign w19306 = ~w11367 & ~w11366;
assign w19307 = w3645 & w20391;
assign w19308 = w3833 & ~pi091;
assign w19309 = ~pi094 & w3547;
assign w19310 = w3771 & ~pi091;
assign w19311 = w11387 & pi024;
assign w19312 = (w11392 & ~w11382) | (w11392 & w20392) | (~w11382 & w20392);
assign w19313 = w3602 & ~pi091;
assign w19314 = (~w11362 & w20192) | (~w11362 & w20393) | (w20192 & w20393);
assign w19315 = ~w11360 & ~pi529;
assign w19316 = ~w11440 & ~pi529;
assign w19317 = (~pi140 & w7618) | (~pi140 & w20394) | (w7618 & w20394);
assign w19318 = ~w7618 & w20395;
assign w19319 = ~w554 & ~pi529;
assign w19320 = ~w11472 & pi001;
assign w19321 = w927 & pi001;
assign w19322 = w11485 & ~w11487;
assign w19323 = ~w410 & ~w536;
assign w19324 = ~w11507 & w20396;
assign w19325 = w1152 & ~pi114;
assign w19326 = w11510 & ~pi001;
assign w19327 = pi007 & ~w938;
assign w19328 = w1132 & pi114;
assign w19329 = (~pi169 & w7618) | (~pi169 & w20397) | (w7618 & w20397);
assign w19330 = ~w7618 & w20398;
assign w19331 = ~w11553 & ~pi529;
assign w19332 = ~w7471 & ~pi152;
assign w19333 = w7471 & pi152;
assign w19334 = ~w11570 & ~pi529;
assign w19335 = ~w1526 & ~pi174;
assign w19336 = w1526 & pi174;
assign w19337 = w11593 & ~pi529;
assign w19338 = ~w11616 & ~pi529;
assign w19339 = (w8301 & w20399) | (w8301 & w20400) | (w20399 & w20400);
assign w19340 = (~w8301 & w20401) | (~w8301 & w20402) | (w20401 & w20402);
assign w19341 = ~w11627 & ~pi529;
assign w19342 = w1696 & w1766;
assign w19343 = w11642 & ~pi026;
assign w19344 = ~w11649 & ~pi115;
assign w19345 = ~w11656 & w1773;
assign w19346 = w11651 & ~pi030;
assign w19347 = w2262 & ~pi115;
assign w19348 = ~w11678 & w20403;
assign w19349 = w11685 & ~pi026;
assign w19350 = ~pi059 & ~w2260;
assign w19351 = w9134 & w20343;
assign w19352 = ~w2060 & ~pi053;
assign w19353 = (~pi089 & w11701) | (~pi089 & w20404) | (w11701 & w20404);
assign w19354 = ~w11727 & pi092;
assign w19355 = pi092 & pi053;
assign w19356 = (~pi089 & w9534) | (~pi089 & w20405) | (w9534 & w20405);
assign w19357 = ~w11740 & ~pi089;
assign w19358 = w2090 & w2172;
assign w19359 = w2099 & ~w5868;
assign w19360 = (~pi089 & ~w2127) | (~pi089 & w20406) | (~w2127 & w20406);
assign w19361 = w11734 & w11749;
assign w19362 = pi071 & pi073;
assign w19363 = ~w11770 & w20407;
assign w19364 = ~pi075 & pi073;
assign w19365 = w11786 & ~w11787;
assign w19366 = w2377 & ~pi080;
assign w19367 = w2336 & pi080;
assign w19368 = w11791 & ~pi073;
assign w19369 = ~w11775 & w20408;
assign w19370 = ~w11771 & ~pi146;
assign w19371 = (w11767 & w20409) | (w11767 & w20410) | (w20409 & w20410);
assign w19372 = ~w9316 & ~pi529;
assign w19373 = ~w8667 & ~w1581;
assign w19374 = ~w11828 & pi117;
assign w19375 = ~pi061 & pi002;
assign w19376 = w1859 & pi002;
assign w19377 = ~w11829 & ~w11833;
assign w19378 = w1555 & w1591;
assign w19379 = w1868 & ~pi117;
assign w19380 = ~w1566 & ~w1662;
assign w19381 = w11870 & ~pi002;
assign w19382 = ~w11860 & w20411;
assign w19383 = ~w11771 & ~pi273;
assign w19384 = (w11767 & w20412) | (w11767 & w20413) | (w20412 & w20413);
assign w19385 = w11896 & ~pi529;
assign w19386 = ~w8719 & ~pi529;
assign w19387 = ~w2430 & ~pi283;
assign w19388 = w2430 & pi283;
assign w19389 = w11947 & ~pi529;
assign w19390 = ~w1983 & ~w8575;
assign w19391 = ~w11971 & ~pi026;
assign w19392 = pi056 & pi115;
assign w19393 = pi115 & ~w11974;
assign w19394 = w2013 & w20414;
assign w19395 = w1966 & w1730;
assign w19396 = (pi030 & ~w11980) | (pi030 & w20415) | (~w11980 & w20415);
assign w19397 = ~pi115 & ~w1710;
assign w19398 = ~w11986 & pi026;
assign w19399 = pi026 & ~w8573;
assign w19400 = ~w12002 & w12003;
assign w19401 = w12000 & w20416;
assign w19402 = ~w12044 & w9060;
assign w19403 = pi117 & ~w9301;
assign w19404 = w9018 & w1577;
assign w19405 = (pi036 & ~w12058) | (pi036 & w20417) | (~w12058 & w20417);
assign w19406 = ~pi117 & ~w1560;
assign w19407 = ~w12065 & pi002;
assign w19408 = ~w12082 & ~w1858;
assign w19409 = ~w12078 & w1588;
assign w19410 = ~w12075 & ~w12060;
assign w19411 = ~w9657 & ~pi230;
assign w19412 = w9657 & pi230;
assign w19413 = ~w12127 & ~pi529;
assign w19414 = ~w12147 & ~pi529;
assign w19415 = (~pi148 & w10203) | (~pi148 & w20418) | (w10203 & w20418);
assign w19416 = ~w10203 & w20419;
assign w19417 = w10170 & ~pi167;
assign w19418 = ~w10170 & pi167;
assign w19419 = ~w12193 & ~pi529;
assign w19420 = (~pi223 & w10203) | (~pi223 & w20420) | (w10203 & w20420);
assign w19421 = ~w10203 & w20421;
assign w19422 = ~w12210 & ~pi529;
assign w19423 = ~w3012 & ~pi376;
assign w19424 = w3012 & pi376;
assign w19425 = w10005 & ~w5945;
assign w19426 = (w19425 & w20941) | (w19425 & w20942) | (w20941 & w20942);
assign w19427 = w10310 & pi003;
assign w19428 = (~w12241 & w20361) | (~w12241 & w20943) | (w20361 & w20943);
assign w19429 = w12261 & w20422;
assign w19430 = w2448 & pi120;
assign w19431 = w2461 & pi120;
assign w19432 = w12289 & ~w12285;
assign w19433 = ~w12252 & w12290;
assign w19434 = ~w10198 & w18604;
assign w19435 = ~w12370 & ~w12384;
assign w19436 = w6300 & w3286;
assign w19437 = w3300 & ~pi090;
assign w19438 = w12408 & ~pi088;
assign w19439 = pi112 & ~w3249;
assign w19440 = ~w12405 & w20423;
assign w19441 = ~w12444 & ~pi529;
assign w19442 = (w10625 & w20424) | (w10625 & w20425) | (w20424 & w20425);
assign w19443 = (~w10625 & w20426) | (~w10625 & w20427) | (w20426 & w20427);
assign w19444 = ~w12500 & ~pi529;
assign w19445 = ~w11301 & ~pi529;
assign w19446 = ~w12591 & ~pi529;
assign w19447 = ~w12608 & ~pi529;
assign w19448 = ~w7914 & ~pi372;
assign w19449 = w7914 & pi372;
assign w19450 = (w7945 & w20428) | (w7945 & w20429) | (w20428 & w20429);
assign w19451 = (~w7945 & w20430) | (~w7945 & w20431) | (w20430 & w20431);
assign w19452 = ~w12619 & ~pi529;
assign w19453 = ~w3516 & ~pi166;
assign w19454 = w3516 & pi166;
assign w19455 = ~w11443 & ~pi529;
assign w19456 = (~pi133 & w7618) | (~pi133 & w20432) | (w7618 & w20432);
assign w19457 = ~w7618 & w20433;
assign w19458 = (w612 & w20434) | (w612 & w20435) | (w20434 & w20435);
assign w19459 = (~w612 & w20436) | (~w612 & w20437) | (w20436 & w20437);
assign w19460 = w12781 & ~pi529;
assign w19461 = w1126 & ~pi165;
assign w19462 = ~w1126 & pi165;
assign w19463 = ~w11530 & ~pi529;
assign w19464 = w12812 & ~pi529;
assign w19465 = (~w11767 & w20438) | (~w11767 & w20439) | (w20438 & w20439);
assign w19466 = (w11767 & w20440) | (w11767 & w20441) | (w20440 & w20441);
assign w19467 = w12829 & ~pi529;
assign w19468 = ~w2197 & ~pi373;
assign w19469 = w2197 & pi373;
assign w19470 = w12858 & ~pi529;
assign w19471 = (w5705 & w20442) | (w5705 & w20443) | (w20442 & w20443);
assign w19472 = (~w5705 & w20444) | (~w5705 & w20445) | (w20444 & w20445);
assign w19473 = ~w12916 & ~pi529;
assign w19474 = (w6298 & w20446) | (w6298 & w20447) | (w20446 & w20447);
assign w19475 = (~w6298 & w20448) | (~w6298 & w20449) | (w20448 & w20449);
assign w19476 = w12971 & ~pi529;
assign w19477 = (~pi218 & w5275) | (~pi218 & w20450) | (w5275 & w20450);
assign w19478 = ~w5275 & w20451;
assign w19479 = ~w13056 & ~pi529;
assign w19480 = ~w11581 & ~pi529;
assign w19481 = ~w11941 & ~pi529;
assign w19482 = ~w13148 & ~pi529;
assign w19483 = ~w9918 & ~pi529;
assign w19484 = ~pi215 & ~pi285;
assign w19485 = ~w13188 & ~w13196;
assign w19486 = pi232 & ~pi231;
assign w19487 = pi270 & pi233;
assign w19488 = w13241 & w13236;
assign w19489 = w13248 & w19542;
assign w19490 = ~w13272 & ~w13264;
assign w19491 = ~pi232 & pi175;
assign w19492 = w13282 & ~pi231;
assign w19493 = (~pi234 & ~w13286) | (~pi234 & w20452) | (~w13286 & w20452);
assign w19494 = w13289 & w13190;
assign w19495 = ~pi270 & ~pi232;
assign w19496 = ~w13300 & pi285;
assign w19497 = w13294 & ~pi215;
assign w19498 = ~w13246 & pi234;
assign w19499 = ~w13324 & ~pi131;
assign w19500 = w13324 & pi131;
assign w19501 = ~w7471 & ~pi258;
assign w19502 = w7471 & pi258;
assign w19503 = w13375 & ~pi529;
assign w19504 = (~w11767 & w20453) | (~w11767 & w20454) | (w20453 & w20454);
assign w19505 = (w11767 & w20455) | (w11767 & w20456) | (w20455 & w20456);
assign w19506 = w13413 & ~pi529;
assign w19507 = ~w13427 & ~pi529;
assign w19508 = (w5705 & w20457) | (w5705 & w20458) | (w20457 & w20458);
assign w19509 = (~w5705 & w20459) | (~w5705 & w20460) | (w20459 & w20460);
assign w19510 = pi157 & ~pi351;
assign w19511 = pi157 & pi132;
assign w19512 = ~w13483 & pi284;
assign w19513 = ~pi132 & ~pi157;
assign w19514 = w13484 & w20461;
assign w19515 = ~pi157 & pi358;
assign w19516 = w13509 & pi275;
assign w19517 = w13506 & w13508;
assign w19518 = w13521 & w20462;
assign w19519 = pi157 & pi358;
assign w19520 = pi358 & pi351;
assign w19521 = w13526 & w13508;
assign w19522 = w13502 & ~pi351;
assign w19523 = w13541 & pi358;
assign w19524 = pi358 & ~pi275;
assign w19525 = w13552 & ~w13551;
assign w19526 = w13472 & w19762;
assign w19527 = ~w13517 & ~w13566;
assign w19528 = ~pi358 & ~pi275;
assign w19529 = ~w13584 & ~w13585;
assign w19530 = ~pi157 & pi351;
assign w19531 = w13593 & ~pi132;
assign w19532 = pi157 & ~pi284;
assign w19533 = ~pi157 & ~pi358;
assign w19534 = w13615 & ~w13602;
assign w19535 = ~w13616 & ~pi193;
assign w19536 = ~w13617 & w20463;
assign w19537 = (pi388 & w13617) | (pi388 & w20464) | (w13617 & w20464);
assign w19538 = ~w13324 & ~pi130;
assign w19539 = w13324 & pi130;
assign w19540 = w13324 & ~w13654;
assign w19541 = ~w13324 & w13654;
assign w19542 = ~pi232 & pi231;
assign w19543 = pi270 & ~pi215;
assign w19544 = w13277 & ~pi175;
assign w19545 = w13237 & w13296;
assign w19546 = pi232 & ~pi175;
assign w19547 = ~pi232 & ~pi175;
assign w19548 = w13682 & ~w13672;
assign w19549 = ~w13691 & pi231;
assign w19550 = w13295 & w20465;
assign w19551 = w13195 & ~w13687;
assign w19552 = w13204 & ~pi285;
assign w19553 = ~w13727 & pi285;
assign w19554 = ~pi233 & pi285;
assign w19555 = ~pi233 & ~pi231;
assign w19556 = w13693 & w13760;
assign w19557 = w13758 & ~w13761;
assign w19558 = ~pi234 & w13762;
assign w19559 = (w13667 & w20466) | (w13667 & w20467) | (w20466 & w20467);
assign w19560 = ~w13765 & ~pi149;
assign w19561 = (~w13701 & w20468) | (~w13701 & w20469) | (w20468 & w20469);
assign w19562 = w13510 & w19530;
assign w19563 = ~w13779 & ~w13783;
assign w19564 = (w13776 & w14528) | (w13776 & w20470) | (w14528 & w20470);
assign w19565 = w13797 & ~pi351;
assign w19566 = ~w13795 & ~pi284;
assign w19567 = (~w13784 & w20471) | (~w13784 & w20472) | (w20471 & w20472);
assign w19568 = ~w13465 & ~pi351;
assign w19569 = (pi193 & w13836) | (pi193 & w20473) | (w13836 & w20473);
assign w19570 = w13585 & w13544;
assign w19571 = w13853 & w13855;
assign w19572 = w13541 & ~pi275;
assign w19573 = (w13806 & w20474) | (w13806 & w20475) | (w20474 & w20475);
assign w19574 = (~w13806 & w20476) | (~w13806 & w20477) | (w20476 & w20477);
assign w19575 = (w13806 & w20478) | (w13806 & w20479) | (w20478 & w20479);
assign w19576 = (~w13806 & w20480) | (~w13806 & w20481) | (w20480 & w20481);
assign w19577 = ~w13910 & ~w13913;
assign w19578 = ~w13935 & pi372;
assign w19579 = pi170 & pi352;
assign w19580 = w13948 & w13965;
assign w19581 = pi321 & pi191;
assign w19582 = ~pi170 & pi321;
assign w19583 = w13988 & w14040;
assign w19584 = ~pi321 & ~pi276;
assign w19585 = ~w13905 & pi372;
assign w19586 = w13997 & ~w14000;
assign w19587 = ~w14007 & ~pi352;
assign w19588 = w13973 & ~w13915;
assign w19589 = w14024 & pi352;
assign w19590 = w13994 & w13938;
assign w19591 = w14031 & w20482;
assign w19592 = w14043 & w14045;
assign w19593 = w14014 & ~pi276;
assign w19594 = ~w14046 & w14050;
assign w19595 = w14052 & w13903;
assign w19596 = ~w14052 & ~w13903;
assign w19597 = ~w14071 & ~w13545;
assign w19598 = ~w13470 & ~pi193;
assign w19599 = w14089 & ~w14087;
assign w19600 = w13563 & pi351;
assign w19601 = ~w13483 & ~pi284;
assign w19602 = w13528 & ~pi351;
assign w19603 = w14094 & ~w14103;
assign w19604 = ~w13491 & w14108;
assign w19605 = w13497 & ~w13555;
assign w19606 = ~w14110 & ~w14113;
assign w19607 = pi157 & ~pi132;
assign w19608 = ~w14075 & ~w14079;
assign w19609 = pi354 & ~pi351;
assign w19610 = ~w13502 & pi284;
assign w19611 = w13579 & pi351;
assign w19612 = w14123 & pi275;
assign w19613 = ~w13617 & w20483;
assign w19614 = (pi144 & w13617) | (pi144 & w20484) | (w13617 & w20484);
assign w19615 = w14197 & ~pi207;
assign w19616 = w14222 & ~w14199;
assign w19617 = ~pi185 & ~pi147;
assign w19618 = ~pi147 & pi185;
assign w19619 = pi129 & pi185;
assign w19620 = ~pi129 & ~pi185;
assign w19621 = ~w14258 & ~w14259;
assign w19622 = ~w14223 & w20485;
assign w19623 = ~w14193 & ~pi302;
assign w19624 = pi138 & pi302;
assign w19625 = w14280 & ~w14285;
assign w19626 = pi185 & ~pi129;
assign w19627 = pi185 & ~pi207;
assign w19628 = ~w14294 & w14296;
assign w19629 = ~pi207 & pi129;
assign w19630 = ~w14327 & ~w14332;
assign w19631 = ~w14333 & ~pi302;
assign w19632 = w14215 & w20486;
assign w19633 = ~w14335 & w14347;
assign w19634 = (w14263 & w20487) | (w14263 & w20488) | (w20487 & w20488);
assign w19635 = (~w14263 & w20489) | (~w14263 & w20490) | (w20489 & w20490);
assign w19636 = ~w14205 & ~pi302;
assign w19637 = pi166 & ~pi207;
assign w19638 = ~pi129 & pi139;
assign w19639 = ~pi129 & pi207;
assign w19640 = ~w14425 & ~pi207;
assign w19641 = ~w14190 & ~pi139;
assign w19642 = w14438 & w14436;
assign w19643 = w14440 & pi302;
assign w19644 = ~pi207 & ~pi302;
assign w19645 = w14452 & w14453;
assign w19646 = w14459 & w20491;
assign w19647 = (~w14363 & ~w14459) | (~w14363 & w20492) | (~w14459 & w20492);
assign w19648 = ~w13606 & w20493;
assign w19649 = ~w13585 & ~w13796;
assign w19650 = ~w14475 & ~w14488;
assign w19651 = pi351 & ~w14514;
assign w19652 = w14515 & ~pi193;
assign w19653 = ~w14523 & ~pi284;
assign w19654 = pi358 & ~w13792;
assign w19655 = w13502 & w13508;
assign w19656 = (w13701 & w20494) | (w13701 & w20495) | (w20494 & w20495);
assign w19657 = (~w13701 & w20496) | (~w13701 & w20497) | (w20496 & w20497);
assign w19658 = ~pi129 & ~pi138;
assign w19659 = w14589 & ~w14603;
assign w19660 = pi147 & pi185;
assign w19661 = pi129 & ~pi138;
assign w19662 = w14604 & pi139;
assign w19663 = w14292 & w14209;
assign w19664 = w14264 & w19644;
assign w19665 = ~w14627 & pi302;
assign w19666 = w14230 & pi207;
assign w19667 = ~w14667 & pi302;
assign w19668 = w14647 & ~pi139;
assign w19669 = ~w14623 & ~pi190;
assign w19670 = w14623 & pi190;
assign w19671 = w14014 & ~w13916;
assign w19672 = ~pi170 & ~pi182;
assign w19673 = pi352 & ~w13980;
assign w19674 = w13979 & ~w13935;
assign w19675 = ~w13980 & ~pi372;
assign w19676 = ~w14729 & ~w14730;
assign w19677 = pi170 & pi321;
assign w19678 = ~pi342 & pi321;
assign w19679 = w14009 & w14014;
assign w19680 = w13977 & pi372;
assign w19681 = w14771 & w14778;
assign w19682 = (w14687 & w14713) | (w14687 & w20498) | (w14713 & w20498);
assign w19683 = ~w14713 & w20499;
assign w19684 = ~pi276 & pi372;
assign w19685 = ~w14801 & w14802;
assign w19686 = ~w14806 & ~pi352;
assign w19687 = w14809 & pi352;
assign w19688 = ~w13994 & ~w14816;
assign w19689 = w14702 & ~pi352;
assign w19690 = w14836 & w20500;
assign w19691 = ~w14734 & ~w13977;
assign w19692 = ~w13975 & ~w13942;
assign w19693 = ~w14030 & pi372;
assign w19694 = ~pi352 & w14854;
assign w19695 = w14856 & ~w13976;
assign w19696 = w14855 & w14858;
assign w19697 = w14859 & ~pi256;
assign w19698 = ~w14859 & pi256;
assign w19699 = ~pi270 & ~w14890;
assign w19700 = w13315 & pi285;
assign w19701 = pi232 & pi231;
assign w19702 = ~pi231 & ~pi285;
assign w19703 = (~pi234 & ~w13294) | (~pi234 & w20501) | (~w13294 & w20501);
assign w19704 = (w14943 & w20502) | (w14943 & w20503) | (w20502 & w20503);
assign w19705 = pi233 & ~pi231;
assign w19706 = ~w13243 & ~pi231;
assign w19707 = w14958 & ~w14955;
assign w19708 = w13236 & ~pi232;
assign w19709 = ~w14972 & pi285;
assign w19710 = ~w14977 & w20504;
assign w19711 = (pi192 & w14977) | (pi192 & w20505) | (w14977 & w20505);
assign w19712 = ~w13910 & ~w14809;
assign w19713 = w13906 & pi352;
assign w19714 = ~w14040 & ~pi191;
assign w19715 = w14752 & ~w15014;
assign w19716 = w15016 & w15019;
assign w19717 = w13959 & pi352;
assign w19718 = w14703 & w13938;
assign w19719 = w13905 & ~pi352;
assign w19720 = w15057 & ~pi342;
assign w19721 = pi170 & pi372;
assign w19722 = w14790 & pi276;
assign w19723 = ~w15067 & w14992;
assign w19724 = w15067 & ~w14992;
assign w19725 = ~pi182 & pi372;
assign w19726 = ~pi321 & ~pi352;
assign w19727 = w15093 & w15109;
assign w19728 = ~pi170 & pi352;
assign w19729 = ~w15116 & ~pi372;
assign w19730 = w15112 & ~w15117;
assign w19731 = w15014 & w14014;
assign w19732 = ~w15122 & ~w15120;
assign w19733 = w15133 & pi182;
assign w19734 = ~w14703 & ~w15084;
assign w19735 = w14014 & w15138;
assign w19736 = w15147 & w14035;
assign w19737 = ~pi352 & ~pi170;
assign w19738 = (w15156 & w15146) | (w15156 & w20506) | (w15146 & w20506);
assign w19739 = w13765 & ~w15169;
assign w19740 = (w13701 & w20507) | (w13701 & w20508) | (w20507 & w20508);
assign w19741 = w13952 & w14040;
assign w19742 = pi276 & pi321;
assign w19743 = pi276 & ~pi191;
assign w19744 = ~w15204 & w15205;
assign w19745 = w15195 & w15199;
assign w19746 = ~w14023 & ~pi352;
assign w19747 = ~pi276 & ~pi372;
assign w19748 = pi352 & ~w14719;
assign w19749 = w15195 & w15232;
assign w19750 = w14031 & ~pi352;
assign w19751 = ~w15185 & ~pi301;
assign w19752 = w15185 & pi301;
assign w19753 = ~w13554 & pi284;
assign w19754 = w13459 & w19859;
assign w19755 = ~w15279 & w15286;
assign w19756 = w15290 & ~w13563;
assign w19757 = ~w15298 & pi193;
assign w19758 = w13474 & pi354;
assign w19759 = pi132 & w15303;
assign w19760 = w15300 & w13562;
assign w19761 = ~pi132 & ~pi284;
assign w19762 = pi275 & pi351;
assign w19763 = ~w15329 & ~pi193;
assign w19764 = w13581 & w13850;
assign w19765 = w15306 & pi284;
assign w19766 = ~w15344 & ~w15299;
assign w19767 = (w14263 & w20509) | (w14263 & w20510) | (w20509 & w20510);
assign w19768 = (~w14263 & w20511) | (~w14263 & w20512) | (w20511 & w20512);
assign w19769 = w13693 & ~w13294;
assign w19770 = ~w13249 & pi231;
assign w19771 = (~pi285 & w15423) | (~pi285 & w20513) | (w15423 & w20513);
assign w19772 = w15422 & ~pi234;
assign w19773 = ~w13180 & pi285;
assign w19774 = ~w13221 & ~pi285;
assign w19775 = ~w13221 & ~w13315;
assign w19776 = ~w19555 & pi285;
assign w19777 = ~pi231 & w15473;
assign w19778 = w13199 & w13236;
assign w19779 = ~w13264 & ~w14973;
assign w19780 = ~w15443 & w20514;
assign w19781 = ~w15440 & w15417;
assign w19782 = w15440 & ~w15417;
assign w19783 = w14214 & pi147;
assign w19784 = w14201 & pi207;
assign w19785 = ~w14436 & pi302;
assign w19786 = ~w14257 & ~pi302;
assign w19787 = ~w15495 & w20515;
assign w19788 = ~w15515 & ~w14339;
assign w19789 = w14249 & w14200;
assign w19790 = w15523 & ~pi139;
assign w19791 = w15549 & ~w14404;
assign w19792 = w15516 & pi302;
assign w19793 = ~w15555 & ~w15510;
assign w19794 = (~w14263 & w20516) | (~w14263 & w20517) | (w20516 & w20517);
assign w19795 = (w14263 & w20518) | (w14263 & w20519) | (w20518 & w20519);
assign w19796 = w14052 & ~pi171;
assign w19797 = ~w14052 & pi171;
assign w19798 = ~w13695 & pi285;
assign w19799 = ~w15611 & ~w15609;
assign w19800 = ~w13249 & pi234;
assign w19801 = w13315 & ~pi231;
assign w19802 = ~w13740 & ~w14956;
assign w19803 = w13224 & w13236;
assign w19804 = ~w13676 & pi285;
assign w19805 = ~pi285 & ~w15618;
assign w19806 = w14890 & pi231;
assign w19807 = (~pi234 & ~w13221) | (~pi234 & w20520) | (~w13221 & w20520);
assign w19808 = ~w13199 & ~w14903;
assign w19809 = ~w15643 & w20521;
assign w19810 = ~w14957 & ~w13204;
assign w19811 = w15653 & w15659;
assign w19812 = w15660 & w15592;
assign w19813 = ~w15660 & ~w15592;
assign w19814 = ~w14822 & ~w14787;
assign w19815 = w13933 & w13965;
assign w19816 = ~w14734 & ~pi352;
assign w19817 = ~w15678 & ~pi372;
assign w19818 = w14014 & pi321;
assign w19819 = w13911 & w14040;
assign w19820 = ~w15182 & ~w15000;
assign w19821 = ~w15713 & ~pi372;
assign w19822 = w15183 & w14774;
assign w19823 = w13917 & w20522;
assign w19824 = w15014 & w15149;
assign w19825 = w14052 & ~w15746;
assign w19826 = ~w14052 & w15746;
assign w19827 = (w10279 & w20523) | (w10279 & w20524) | (w20523 & w20524);
assign w19828 = (~w10279 & w20525) | (~w10279 & w20526) | (w20525 & w20526);
assign w19829 = w13946 & w14030;
assign w19830 = ~pi342 & ~pi372;
assign w19831 = w15781 & w15783;
assign w19832 = w15770 & ~w15784;
assign w19833 = w15790 & ~w14800;
assign w19834 = ~w15791 & ~pi191;
assign w19835 = ~w14008 & ~pi372;
assign w19836 = w14023 & w19721;
assign w19837 = w13979 & pi276;
assign w19838 = ~w14023 & pi372;
assign w19839 = ~w15826 & ~w15825;
assign w19840 = w15832 & ~w15792;
assign w19841 = w14459 & w20527;
assign w19842 = (pi181 & ~w14459) | (pi181 & w20528) | (~w14459 & w20528);
assign w19843 = w14459 & w20529;
assign w19844 = (w15858 & ~w14459) | (w15858 & w20530) | (~w14459 & w20530);
assign w19845 = w15871 & ~pi207;
assign w19846 = ~w15881 & w20531;
assign w19847 = pi185 & pi207;
assign w19848 = w14318 & ~w15903;
assign w19849 = ~w14225 & pi139;
assign w19850 = w14441 & ~pi207;
assign w19851 = w15929 & ~pi302;
assign w19852 = w14193 & ~pi207;
assign w19853 = ~pi129 & ~pi139;
assign w19854 = ~w15896 & ~w15900;
assign w19855 = ~w14470 & w15950;
assign w19856 = pi354 & ~pi284;
assign w19857 = ~w15954 & w15959;
assign w19858 = ~w13465 & ~pi284;
assign w19859 = pi358 & ~pi351;
assign w19860 = pi157 & pi351;
assign w19861 = w14107 & ~pi351;
assign w19862 = pi351 & ~w16002;
assign w19863 = pi275 & ~pi193;
assign w19864 = ~w16004 & w16005;
assign w19865 = ~w15969 & ~w16011;
assign w19866 = (~pi144 & w9258) | (~pi144 & w20532) | (w9258 & w20532);
assign w19867 = ~w9258 & w20533;
assign w19868 = ~w14623 & ~pi187;
assign w19869 = w14623 & pi187;
assign w19870 = (w7325 & w20534) | (w7325 & w20535) | (w20534 & w20535);
assign w19871 = (~w7325 & w20536) | (~w7325 & w20537) | (w20536 & w20537);
assign w19872 = ~w14977 & w20538;
assign w19873 = (pi189 & w14977) | (pi189 & w20539) | (w14977 & w20539);
assign w19874 = w14623 & ~w16063;
assign w19875 = ~w14623 & w16063;
assign w19876 = (~w16081 & w14977) | (~w16081 & w20540) | (w14977 & w20540);
assign w19877 = ~w14977 & w20541;
assign w19878 = ~w10245 & ~pi167;
assign w19879 = ~w10203 & w20542;
assign w19880 = ~w247 & ~pi137;
assign w19881 = w247 & pi137;
assign w19882 = w10170 & ~pi223;
assign w19883 = ~w10170 & pi223;
assign w19884 = ~w6264 & ~pi224;
assign w19885 = w6264 & pi224;
assign w19886 = ~w14470 & ~w15992;
assign w19887 = w16133 & ~w13517;
assign w19888 = ~pi358 & pi351;
assign w19889 = w16135 & pi284;
assign w19890 = w13787 & w13541;
assign w19891 = ~w16143 & ~w16136;
assign w19892 = w16148 & ~w14517;
assign w19893 = w13481 & w19519;
assign w19894 = w14501 & w20543;
assign w19895 = w13464 & w13541;
assign w19896 = ~w13516 & ~w13780;
assign w19897 = ~w16176 & ~w15283;
assign w19898 = ~w16171 & w16179;
assign w19899 = (w8301 & w20544) | (w8301 & w20545) | (w20544 & w20545);
assign w19900 = (~w8301 & w20546) | (~w8301 & w20547) | (w20546 & w20547);
assign w19901 = ~w9657 & ~pi190;
assign w19902 = w9657 & pi190;
assign w19903 = pi175 & ~w14924;
assign w19904 = w16256 & ~pi285;
assign w19905 = w15610 & w13294;
assign w19906 = ~w16259 & w20548;
assign w19907 = w16271 & pi285;
assign w19908 = w13194 & pi231;
assign w19909 = ~w13241 & ~w14961;
assign w19910 = w13182 & w13294;
assign w19911 = ~w16305 & w20549;
assign w19912 = ~w16286 & w16249;
assign w19913 = w16286 & ~w16249;
assign w19914 = w16321 & ~w16318;
assign w19915 = w16326 & pi302;
assign w19916 = ~w16333 & ~w16327;
assign w19917 = w15512 & pi302;
assign w19918 = pi302 & ~w14257;
assign w19919 = ~w14392 & ~w14337;
assign w19920 = w14205 & w14210;
assign w19921 = ~w16360 & ~w16356;
assign w19922 = ~w14253 & ~w14227;
assign w19923 = (pi302 & w16366) | (pi302 & w20550) | (w16366 & w20550);
assign w19924 = ~pi207 & ~w14442;
assign w19925 = (w16381 & w16338) | (w16381 & w20551) | (w16338 & w20551);
assign w19926 = ~w16338 & w20552;
assign w19927 = w15470 & ~pi231;
assign w19928 = ~w16392 & ~pi285;
assign w19929 = (pi285 & w15423) | (pi285 & w20553) | (w15423 & w20553);
assign w19930 = ~w13194 & pi285;
assign w19931 = ~w13236 & pi234;
assign w19932 = ~w13665 & ~pi175;
assign w19933 = w13294 & w16434;
assign w19934 = w16436 & pi175;
assign w19935 = pi231 & pi285;
assign w19936 = w15433 & w19702;
assign w19937 = ~w13676 & ~w13250;
assign w19938 = w16431 & w16449;
assign w19939 = w13294 & w20554;
assign w19940 = w13190 & pi233;
assign w19941 = w16469 & w16474;
assign w19942 = ~w14925 & ~w13282;
assign w19943 = w16513 & w16520;
assign w19944 = w16482 & pi175;
assign w19945 = ~w16525 & w16531;
assign w19946 = w16525 & ~w16531;
assign w19947 = (~pi222 & w14713) | (~pi222 & w20555) | (w14713 & w20555);
assign w19948 = ~w14713 & w20556;
assign w19949 = ~w15067 & ~pi225;
assign w19950 = w15067 & pi225;
assign w19951 = (~w16606 & w14713) | (~w16606 & w20557) | (w14713 & w20557);
assign w19952 = ~w14713 & w20558;
assign w19953 = ~w15067 & ~w16636;
assign w19954 = w15067 & w16636;
assign w19955 = (w11374 & w20559) | (w11374 & w20560) | (w20559 & w20560);
assign w19956 = (~w11374 & w20561) | (~w11374 & w20562) | (w20561 & w20562);
assign w19957 = (w5024 & w20563) | (w5024 & w20564) | (w20563 & w20564);
assign w19958 = (~w5024 & w20565) | (~w5024 & w20566) | (w20565 & w20566);
assign w19959 = w8071 & w20567;
assign w19960 = (pi179 & ~w8071) | (pi179 & w20568) | (~w8071 & w20568);
assign w19961 = ~w3012 & ~pi280;
assign w19962 = w3012 & pi280;
assign w19963 = (w6574 & w20569) | (w6574 & w20570) | (w20569 & w20570);
assign w19964 = (~w6574 & w20571) | (~w6574 & w20572) | (w20571 & w20572);
assign w19965 = w9391 & w20573;
assign w19966 = (pi226 & ~w9391) | (pi226 & w20574) | (~w9391 & w20574);
assign w19967 = ~w6174 & ~pi130;
assign w19968 = w6174 & pi130;
assign w19969 = (w3706 & w20575) | (w3706 & w20576) | (w20575 & w20576);
assign w19970 = (~w3706 & w20577) | (~w3706 & w20578) | (w20577 & w20578);
assign w19971 = (w55 & w20579) | (w55 & w20580) | (w20579 & w20580);
assign w19972 = (~w55 & w20581) | (~w55 & w20582) | (w20581 & w20582);
assign w19973 = (~pi151 & w5275) | (~pi151 & w20583) | (w5275 & w20583);
assign w19974 = ~w5275 & w20584;
assign w19975 = w8455 & ~pi228;
assign w19976 = ~w8455 & pi228;
assign w19977 = ~w14303 & ~w14226;
assign w19978 = w14208 & w19847;
assign w19979 = ~w16722 & w20585;
assign w19980 = w14240 & w14232;
assign w19981 = w14252 & w16325;
assign w19982 = ~w14253 & pi302;
assign w19983 = ~w15897 & ~w16754;
assign w19984 = w15898 & pi207;
assign w19985 = w14611 & w16774;
assign w19986 = w16772 & w16778;
assign w19987 = (~pi302 & w16800) | (~pi302 & w20586) | (w16800 & w20586);
assign w19988 = ~w16805 & pi302;
assign w19989 = (pi139 & ~w16813) | (pi139 & w20587) | (~w16813 & w20587);
assign w19990 = w16828 & w16832;
assign w19991 = w16834 & pi138;
assign w19992 = w14318 & ~pi138;
assign w19993 = ~w14344 & ~w14386;
assign w19994 = w14207 & w14448;
assign w19995 = ~w16833 & ~pi139;
assign w19996 = (w16814 & w20588) | (w16814 & w20589) | (w20588 & w20589);
assign w19997 = (~w16814 & w20590) | (~w16814 & w20591) | (w20590 & w20591);
assign w19998 = ~w4948 & ~pi193;
assign w19999 = (~w4947 & w20592) | (~w4947 & w20593) | (w20592 & w20593);
assign w20000 = (~pi142 & w7618) | (~pi142 & w20594) | (w7618 & w20594);
assign w20001 = ~w7618 & w20595;
assign w20002 = (w744 & w20596) | (w744 & w20597) | (w20596 & w20597);
assign w20003 = (~w744 & w20598) | (~w744 & w20599) | (w20598 & w20599);
assign w20004 = ~w13505 & ~w16169;
assign w20005 = w13470 & w19520;
assign w20006 = w13556 & ~pi351;
assign w20007 = ~w13859 & ~w16140;
assign w20008 = w16906 & ~pi284;
assign w20009 = ~w16909 & w16914;
assign w20010 = w14525 & w13482;
assign w20011 = w15956 & pi351;
assign w20012 = ~w16930 & ~w16172;
assign w20013 = (pi193 & w16932) | (pi193 & w20600) | (w16932 & w20600);
assign w20014 = w13490 & ~pi351;
assign w20015 = ~w16936 & ~pi284;
assign w20016 = w14501 & w14528;
assign w20017 = ~w14470 & ~w13581;
assign w20018 = ~w16937 & ~w16938;
assign w20019 = ~w15185 & ~pi269;
assign w20020 = w15185 & pi269;
assign w20021 = ~w15440 & ~pi271;
assign w20022 = w15440 & pi271;
assign w20023 = ~w15440 & ~w17014;
assign w20024 = w15440 & w17014;
assign w20025 = w15660 & ~pi278;
assign w20026 = ~w15660 & pi278;
assign w20027 = (w1876 & w20601) | (w1876 & w20602) | (w20601 & w20602);
assign w20028 = (~w1876 & w20603) | (~w1876 & w20604) | (w20603 & w20604);
assign w20029 = w15660 & ~w17065;
assign w20030 = ~w15660 & w17065;
assign w20031 = (~pi149 & w9194) | (~pi149 & w20605) | (w9194 & w20605);
assign w20032 = ~w9194 & w20606;
assign w20033 = ~w8485 & ~pi172;
assign w20034 = w8485 & pi172;
assign w20035 = (w5942 & w20607) | (w5942 & w20608) | (w20607 & w20608);
assign w20036 = (~w5942 & w20609) | (~w5942 & w20610) | (w20609 & w20610);
assign w20037 = ~w2197 & ~pi283;
assign w20038 = w2197 & pi283;
assign w20039 = (w11981 & w20611) | (w11981 & w20612) | (w20611 & w20612);
assign w20040 = (~w11981 & w20613) | (~w11981 & w20614) | (w20613 & w20614);
assign w20041 = ~w3516 & ~pi354;
assign w20042 = w3516 & pi354;
assign w20043 = (w8106 & w20615) | (w8106 & w20616) | (w20615 & w20616);
assign w20044 = (~w8106 & w20617) | (~w8106 & w20618) | (w20617 & w20618);
assign w20045 = ~w550 & ~pi221;
assign w20046 = w550 & pi221;
assign w20047 = (w7945 & w20619) | (w7945 & w20620) | (w20619 & w20620);
assign w20048 = (~w7945 & w20621) | (~w7945 & w20622) | (w20621 & w20622);
assign w20049 = (w4689 & w20623) | (w4689 & w20624) | (w20623 & w20624);
assign w20050 = (~w4689 & w20625) | (~w4689 & w20626) | (w20625 & w20626);
assign w20051 = ~w7471 & ~pi169;
assign w20052 = w7471 & pi169;
assign w20053 = ~w1526 & ~pi257;
assign w20054 = w1526 & pi257;
assign w20055 = (w612 & w20627) | (w612 & w20628) | (w20627 & w20628);
assign w20056 = (~w612 & w20629) | (~w612 & w20630) | (w20629 & w20630);
assign w20057 = ~w8843 & ~pi320;
assign w20058 = w8843 & pi320;
assign w20059 = (~w11767 & w20631) | (~w11767 & w20632) | (w20631 & w20632);
assign w20060 = (w11767 & w20633) | (w11767 & w20634) | (w20633 & w20634);
assign w20061 = (w5705 & w20635) | (w5705 & w20636) | (w20635 & w20636);
assign w20062 = (~w5705 & w20637) | (~w5705 & w20638) | (w20637 & w20638);
assign w20063 = (w5098 & w20639) | (w5098 & w20640) | (w20639 & w20640);
assign w20064 = (~w5098 & w20641) | (~w5098 & w20642) | (w20641 & w20642);
assign w20065 = (w9016 & w20643) | (w9016 & w20644) | (w20643 & w20644);
assign w20066 = (~w9016 & w20645) | (~w9016 & w20646) | (w20645 & w20646);
assign w20067 = (w5601 & w20647) | (w5601 & w20648) | (w20647 & w20648);
assign w20068 = (~w5601 & w20649) | (~w5601 & w20650) | (w20649 & w20650);
assign w20069 = (w5818 & w20651) | (w5818 & w20652) | (w20651 & w20652);
assign w20070 = (~w5818 & w20653) | (~w5818 & w20654) | (w20653 & w20654);
assign w20071 = ~w7914 & ~pi285;
assign w20072 = w7914 & pi285;
assign w20073 = w3658 & w20655;
assign w20074 = (pi166 & ~w3658) | (pi166 & w20656) | (~w3658 & w20656);
assign w20075 = w1126 & ~pi219;
assign w20076 = ~w1126 & pi219;
assign w20077 = w2743 & ~pi353;
assign w20078 = ~w2743 & pi353;
assign w20079 = (~w10791 & w20657) | (~w10791 & w20658) | (w20657 & w20658);
assign w20080 = (w10791 & w20659) | (w10791 & w20660) | (w20659 & w20660);
assign w20081 = (w6298 & w20661) | (w6298 & w20662) | (w20661 & w20662);
assign w20082 = (~w6298 & w20663) | (~w6298 & w20664) | (w20663 & w20664);
assign w20083 = (w4482 & w20665) | (w4482 & w20666) | (w20665 & w20666);
assign w20084 = (~w4482 & w20667) | (~w4482 & w20668) | (w20667 & w20668);
assign w20085 = (w3809 & w20669) | (w3809 & w20670) | (w20669 & w20670);
assign w20086 = (~w3809 & w20671) | (~w3809 & w20672) | (w20671 & w20672);
assign w20087 = ~w16286 & ~pi371;
assign w20088 = w16286 & pi371;
assign w20089 = ~w2430 & ~pi373;
assign w20090 = w2430 & pi373;
assign w20091 = (~pi349 & w16338) | (~pi349 & w20673) | (w16338 & w20673);
assign w20092 = ~w16338 & w20674;
assign w20093 = ~w16286 & ~w17323;
assign w20094 = w16286 & w17323;
assign w20095 = (~w17332 & w16338) | (~w17332 & w20675) | (w16338 & w20675);
assign w20096 = ~w16338 & w20676;
assign w20097 = ~w10626 & ~pi171;
assign w20098 = (~w10625 & w20677) | (~w10625 & w20678) | (w20677 & w20678);
assign w20099 = ~w16525 & ~pi356;
assign w20100 = w16525 & pi356;
assign w20101 = ~w16525 & ~w17365;
assign w20102 = w16525 & w17365;
assign w20103 = w1020 & ~pi165;
assign w20104 = ~w1020 & pi165;
assign w20105 = w2595 & ~pi161;
assign w20106 = ~w2595 & pi161;
assign w20107 = (~w10347 & w20679) | (~w10347 & w20680) | (w20679 & w20680);
assign w20108 = (w10347 & w20681) | (w10347 & w20682) | (w20681 & w20682);
assign w20109 = w4438 & ~pi207;
assign w20110 = ~w4438 & pi207;
assign w20111 = w8616 & ~pi357;
assign w20112 = ~w8616 & pi357;
assign w20113 = w1691 & ~pi163;
assign w20114 = ~w1691 & pi163;
assign w20115 = (w11660 & w20683) | (w11660 & w20684) | (w20683 & w20684);
assign w20116 = (~w11660 & w20685) | (~w11660 & w20686) | (w20685 & w20686);
assign w20117 = ~w1840 & ~pi375;
assign w20118 = w1840 & pi375;
assign w20119 = (w1390 & w20687) | (w1390 & w20688) | (w20687 & w20688);
assign w20120 = (~w1390 & w20689) | (~w1390 & w20690) | (w20689 & w20690);
assign w20121 = (w4869 & w20691) | (w4869 & w20692) | (w20691 & w20692);
assign w20122 = (~w4869 & w20693) | (~w4869 & w20694) | (w20693 & w20694);
assign w20123 = pi482 & pi396;
assign w20124 = ~w17461 & ~w17463;
assign w20125 = ~pi532 & pi520;
assign w20126 = (~pi532 & ~w17458) | (~pi532 & w20125) | (~w17458 & w20125);
assign w20127 = ~pi396 & ~w17463;
assign w20128 = pi532 & ~w17475;
assign w20129 = pi390 & pi387;
assign w20130 = ~pi390 & pi387;
assign w20131 = pi393 & ~pi395;
assign w20132 = w0 & ~pi083;
assign w20133 = ~pi040 & w17897;
assign w20134 = pi078 & ~pi040;
assign w20135 = pi078 & w17898;
assign w20136 = ~pi078 & pi040;
assign w20137 = w13 & w20136;
assign w20138 = ~w158 & ~pi040;
assign w20139 = pi040 & w17911;
assign w20140 = ~w202 & ~pi083;
assign w20141 = ~pi078 & w17913;
assign w20142 = ~pi069 & pi102;
assign w20143 = pi127 & ~pi104;
assign w20144 = ~pi102 & w17955;
assign w20145 = pi012 & ~pi102;
assign w20146 = pi012 & w17957;
assign w20147 = ~w703 & ~pi102;
assign w20148 = ~w706 & w20695;
assign w20149 = w958 & ~pi001;
assign w20150 = w934 & ~pi001;
assign w20151 = w258 & ~pi123;
assign w20152 = pi040 & pi078;
assign w20153 = pi107 & w88;
assign w20154 = pi048 & w18050;
assign w20155 = ~w304 & ~pi048;
assign w20156 = ~pi027 & w1416;
assign w20157 = ~pi020 & pi048;
assign w20158 = ~pi020 & w18054;
assign w20159 = pi063 & pi104;
assign w20160 = pi102 & pi012;
assign w20161 = ~pi069 & w645;
assign w20162 = w1552 & ~pi117;
assign w20163 = w1611 & pi117;
assign w20164 = pi059 & ~pi115;
assign w20165 = ~pi026 & w18095;
assign w20166 = w1719 & ~pi115;
assign w20167 = pi089 & w18136;
assign w20168 = ~pi028 & w2172;
assign w20169 = pi026 & pi030;
assign w20170 = ~pi008 & w2265;
assign w20171 = ~w2368 & ~pi073;
assign w20172 = pi075 & w2409;
assign w20173 = ~w2347 & w2403;
assign w20174 = w2453 & ~pi003;
assign w20175 = w2524 & pi003;
assign w20176 = pi103 & ~pi118;
assign w20177 = w2676 & pi118;
assign w20178 = pi034 & w18199;
assign w20179 = ~pi120 & ~pi003;
assign w20180 = w2993 & pi058;
assign w20181 = pi058 & pi060;
assign w20182 = ~pi011 & w3075;
assign w20183 = w2613 & w3181;
assign w20184 = pi088 & w18254;
assign w20185 = w3207 & w3295;
assign w20186 = ~pi017 & pi039;
assign w20187 = w3440 & w20186;
assign w20188 = ~pi024 & w18274;
assign w20189 = w3593 & ~pi024;
assign w20190 = pi017 & pi039;
assign w20191 = ~w3664 & w20696;
assign w20192 = pi018 & ~pi024;
assign w20193 = ~w3772 & w20697;
assign w20194 = ~pi043 & ~pi039;
assign w20195 = pi039 & w3674;
assign w20196 = (pi039 & w3674) | (pi039 & w7824) | (w3674 & w7824);
assign w20197 = ~w3474 & ~pi039;
assign w20198 = pi065 & w18354;
assign w20199 = pi068 & pi065;
assign w20200 = pi068 & w18355;
assign w20201 = pi025 & pi113;
assign w20202 = pi096 & w18368;
assign w20203 = w4614 & pi010;
assign w20204 = ~w4631 & ~w4632;
assign w20205 = ~pi010 & pi096;
assign w20206 = ~pi010 & w18371;
assign w20207 = w4666 & pi113;
assign w20208 = ~pi010 & pi113;
assign w20209 = ~pi010 & w18381;
assign w20210 = pi191 & ~pi010;
assign w20211 = pi191 & w18388;
assign w20212 = ~w3620 & ~pi091;
assign w20213 = pi122 & pi017;
assign w20214 = ~w3701 & ~pi122;
assign w20215 = pi048 & w18430;
assign w20216 = pi020 & pi048;
assign w20217 = pi020 & w18431;
assign w20218 = pi001 & w18444;
assign w20219 = ~w436 & ~pi001;
assign w20220 = pi029 & ~pi001;
assign w20221 = ~w5078 & w20698;
assign w20222 = w5277 & ~pi040;
assign w20223 = pi078 & w18466;
assign w20224 = pi020 & ~pi048;
assign w20225 = ~w5330 & w20699;
assign w20226 = ~pi121 & ~pi012;
assign w20227 = (w716 & w20700) | (w716 & w20701) | (w20700 & w20701);
assign w20228 = pi121 & pi012;
assign w20229 = (~w716 & w20702) | (~w716 & w20703) | (w20702 & w20703);
assign w20230 = ~pi150 & pi012;
assign w20231 = (~pi150 & ~w610) | (~pi150 & w20230) | (~w610 & w20230);
assign w20232 = pi150 & ~pi012;
assign w20233 = w610 & w20232;
assign w20234 = w1330 & pi078;
assign w20235 = pi075 & ~pi080;
assign w20236 = ~pi073 & w18517;
assign w20237 = ~pi015 & pi073;
assign w20238 = w2377 & w20237;
assign w20239 = pi190 & ~pi015;
assign w20240 = (~w5686 & w20704) | (~w5686 & w20705) | (w20704 & w20705);
assign w20241 = w2187 & pi089;
assign w20242 = ~pi053 & pi089;
assign w20243 = ~pi053 & w18537;
assign w20244 = pi136 & pi012;
assign w20245 = (~w716 & w20706) | (~w716 & w20707) | (w20706 & w20707);
assign w20246 = pi044 & pi003;
assign w20247 = ~w5916 & w20708;
assign w20248 = w2958 & pi058;
assign w20249 = w2978 & ~pi116;
assign w20250 = ~pi058 & w18565;
assign w20251 = ~pi034 & w18569;
assign w20252 = pi034 & w18574;
assign w20253 = ~pi038 & pi034;
assign w20254 = ~pi038 & w18575;
assign w20255 = ~pi011 & pi058;
assign w20256 = pi097 & ~pi058;
assign w20257 = w6204 & pi116;
assign w20258 = w3258 & ~pi090;
assign w20259 = w3207 & ~pi088;
assign w20260 = pi006 & ~pi088;
assign w20261 = ~w6304 & w20709;
assign w20262 = ~pi051 & pi090;
assign w20263 = pi088 & w18612;
assign w20264 = ~pi006 & pi088;
assign w20265 = ~pi006 & w18613;
assign w20266 = ~pi187 & pi006;
assign w20267 = (~pi187 & ~w6286) | (~pi187 & w20266) | (~w6286 & w20266);
assign w20268 = pi187 & ~pi006;
assign w20269 = w6286 & w20268;
assign w20270 = w6015 & ~pi058;
assign w20271 = pi060 & ~pi058;
assign w20272 = pi060 & w18633;
assign w20273 = w2669 & pi034;
assign w20274 = ~w2625 & w3172;
assign w20275 = ~pi000 & pi022;
assign w20276 = ~pi113 & ~pi096;
assign w20277 = w4124 & pi096;
assign w20278 = w7028 & ~pi096;
assign w20279 = w4197 & ~pi113;
assign w20280 = ~pi096 & w18705;
assign w20281 = w4018 & pi065;
assign w20282 = ~pi065 & w4838;
assign w20283 = ~pi065 & w18710;
assign w20284 = w4015 & ~pi065;
assign w20285 = w264 & pi048;
assign w20286 = w506 & ~pi001;
assign w20287 = pi029 & w18738;
assign w20288 = ~w7423 & ~pi078;
assign w20289 = ~w7490 & ~pi012;
assign w20290 = ~w7556 & ~pi020;
assign w20291 = w1063 & pi123;
assign w20292 = w579 & ~pi104;
assign w20293 = w755 & pi102;
assign w20294 = ~pi012 & pi179;
assign w20295 = pi109 & pi122;
assign w20296 = ~w4047 & ~pi065;
assign w20297 = w4467 & w7896;
assign w20298 = w4719 & pi096;
assign w20299 = pi010 & pi096;
assign w20300 = pi010 & w18820;
assign w20301 = ~w4181 & ~pi096;
assign w20302 = ~pi009 & w4726;
assign w20303 = ~pi302 & ~pi010;
assign w20304 = ~pi302 & ~w18824;
assign w20305 = pi302 & pi010;
assign w20306 = pi302 & w18824;
assign w20307 = (~pi142 & w8059) | (~pi142 & w20710) | (w8059 & w20710);
assign w20308 = ~w8059 & w20711;
assign w20309 = w428 & ~pi001;
assign w20310 = (~pi029 & w1186) | (~pi029 & w20712) | (w1186 & w20712);
assign w20311 = ~pi013 & ~pi001;
assign w20312 = w455 & w20713;
assign w20313 = pi065 & w18868;
assign w20314 = w8206 & w4529;
assign w20315 = ~pi012 & ~pi102;
assign w20316 = w856 & w20714;
assign w20317 = pi164 & pi012;
assign w20318 = w8292 & w20317;
assign w20319 = ~pi154 & ~pi012;
assign w20320 = (~pi154 & ~w8292) | (~pi154 & w20319) | (~w8292 & w20319);
assign w20321 = pi154 & pi012;
assign w20322 = w8292 & w20321;
assign w20323 = ~w8391 & ~pi089;
assign w20324 = ~w8391 & ~w18890;
assign w20325 = pi050 & pi092;
assign w20326 = pi089 & w18903;
assign w20327 = pi089 & w18910;
assign w20328 = ~pi053 & w18911;
assign w20329 = pi110 & pi080;
assign w20330 = pi073 & w18931;
assign w20331 = w18941 & pi073;
assign w20332 = pi015 & pi073;
assign w20333 = pi015 & w18935;
assign w20334 = ~w8965 & w20715;
assign w20335 = ~w8631 & ~pi002;
assign w20336 = pi036 & ~pi002;
assign w20337 = ~w8994 & w20716;
assign w20338 = w2048 & pi089;
assign w20339 = w2241 & ~pi115;
assign w20340 = w1664 & ~pi002;
assign w20341 = ~w9248 & pi002;
assign w20342 = ~w9248 & ~w19003;
assign w20343 = ~pi085 & ~pi092;
assign w20344 = (~pi178 & w9376) | (~pi178 & w20717) | (w9376 & w20717);
assign w20345 = ~w9376 & w20718;
assign w20346 = w1677 & ~pi002;
assign w20347 = pi002 & pi036;
assign w20348 = w1677 & w9244;
assign w20349 = ~pi067 & w9051;
assign w20350 = w8876 & ~pi073;
assign w20351 = w9596 & ~w2295;
assign w20352 = w2333 & pi073;
assign w20353 = w2381 & pi080;
assign w20354 = w8750 & pi073;
assign w20355 = ~pi074 & ~pi003;
assign w20356 = ~pi103 & ~pi118;
assign w20357 = w2660 & w6164;
assign w20358 = pi006 & ~pi141;
assign w20359 = ~pi006 & pi141;
assign w20360 = ~w2828 & ~pi003;
assign w20361 = pi044 & ~pi003;
assign w20362 = pi044 & w19161;
assign w20363 = (pi038 & ~w10350) | (pi038 & w20719) | (~w10350 & w20719);
assign w20364 = w10367 & ~pi038;
assign w20365 = ~w10431 & ~pi044;
assign w20366 = (w10501 & w20720) | (w10501 & w20721) | (w20720 & w20721);
assign w20367 = w10503 & ~w19189;
assign w20368 = ~w3041 & ~pi058;
assign w20369 = ~w10607 & w20722;
assign w20370 = w3041 & pi058;
assign w20371 = ~pi128 & ~pi106;
assign w20372 = w3982 & w4529;
assign w20373 = (pi017 & ~w10792) | (pi017 & w20213) | (~w10792 & w20213);
assign w20374 = ~w10801 & ~pi017;
assign w20375 = ~w10885 & ~pi018;
assign w20376 = ~pi125 & ~pi113;
assign w20377 = w4198 & ~pi096;
assign w20378 = ~w11020 & pi010;
assign w20379 = w4056 & ~pi065;
assign w20380 = w3982 & pi065;
assign w20381 = (w11175 & w7198) | (w11175 & w20723) | (w7198 & w20723);
assign w20382 = ~pi005 & w3858;
assign w20383 = ~pi284 & ~pi010;
assign w20384 = ~pi284 & ~w18824;
assign w20385 = pi284 & pi010;
assign w20386 = pi284 & w18824;
assign w20387 = ~pi233 & pi010;
assign w20388 = ~pi233 & ~w18388;
assign w20389 = pi233 & ~pi010;
assign w20390 = pi233 & w18388;
assign w20391 = ~w3547 & ~pi024;
assign w20392 = w3645 & w20724;
assign w20393 = pi018 & w19307;
assign w20394 = pi012 & ~pi140;
assign w20395 = ~pi012 & pi140;
assign w20396 = ~w11505 & ~pi029;
assign w20397 = pi012 & ~pi169;
assign w20398 = ~pi012 & pi169;
assign w20399 = ~pi155 & ~pi012;
assign w20400 = (~pi155 & ~w8292) | (~pi155 & w20399) | (~w8292 & w20399);
assign w20401 = pi155 & pi012;
assign w20402 = w8292 & w20401;
assign w20403 = (pi030 & ~w11676) | (pi030 & w20725) | (~w11676 & w20725);
assign w20404 = w11702 & ~pi089;
assign w20405 = w8458 & ~pi089;
assign w20406 = ~w2111 & ~pi089;
assign w20407 = (pi015 & ~w11768) | (pi015 & w20726) | (~w11768 & w20726);
assign w20408 = ~w11777 & ~pi015;
assign w20409 = pi146 & pi015;
assign w20410 = ~w11770 & w20727;
assign w20411 = ~w11862 & ~pi036;
assign w20412 = pi273 & pi015;
assign w20413 = ~w11770 & w20728;
assign w20414 = w1752 & pi026;
assign w20415 = w11977 & pi030;
assign w20416 = ~w1744 & ~pi026;
assign w20417 = w12056 & pi036;
assign w20418 = pi006 & ~pi148;
assign w20419 = ~pi006 & pi148;
assign w20420 = pi006 & ~pi223;
assign w20421 = ~pi006 & pi223;
assign w20422 = w2480 & ~pi003;
assign w20423 = ~w12404 & ~pi006;
assign w20424 = ~pi181 & ~pi060;
assign w20425 = (w10612 & w20729) | (w10612 & w20730) | (w20729 & w20730);
assign w20426 = pi181 & pi060;
assign w20427 = (~w10612 & w20731) | (~w10612 & w20732) | (w20731 & w20732);
assign w20428 = ~pi285 & ~pi010;
assign w20429 = ~pi285 & ~w18824;
assign w20430 = pi285 & pi010;
assign w20431 = pi285 & w18824;
assign w20432 = pi012 & ~pi133;
assign w20433 = ~pi012 & pi133;
assign w20434 = ~pi156 & pi012;
assign w20435 = (~pi156 & ~w610) | (~pi156 & w20434) | (~w610 & w20434);
assign w20436 = pi156 & ~pi012;
assign w20437 = w610 & w20436;
assign w20438 = ~pi227 & ~pi015;
assign w20439 = (~pi227 & w11770) | (~pi227 & w20733) | (w11770 & w20733);
assign w20440 = pi227 & pi015;
assign w20441 = ~w11770 & w20734;
assign w20442 = ~pi163 & pi015;
assign w20443 = (w5686 & w20735) | (w5686 & w20736) | (w20735 & w20736);
assign w20444 = pi163 & ~pi015;
assign w20445 = (~w5686 & w20737) | (~w5686 & w20738) | (w20737 & w20738);
assign w20446 = ~pi224 & pi006;
assign w20447 = (~pi224 & ~w6286) | (~pi224 & w20446) | (~w6286 & w20446);
assign w20448 = pi224 & ~pi006;
assign w20449 = w6286 & w20448;
assign w20450 = pi078 & ~pi218;
assign w20451 = ~pi078 & pi218;
assign w20452 = ~w13278 & w20502;
assign w20453 = ~pi348 & ~pi015;
assign w20454 = (~pi348 & w11770) | (~pi348 & w20739) | (w11770 & w20739);
assign w20455 = pi348 & pi015;
assign w20456 = ~w11770 & w20740;
assign w20457 = ~pi228 & pi015;
assign w20458 = (w5686 & w20741) | (w5686 & w20742) | (w20741 & w20742);
assign w20459 = pi228 & ~pi015;
assign w20460 = (~w5686 & w20743) | (~w5686 & w20744) | (w20743 & w20744);
assign w20461 = ~pi358 & ~pi351;
assign w20462 = ~w13522 & ~w13501;
assign w20463 = w13549 & ~pi388;
assign w20464 = ~w13549 & pi388;
assign w20465 = w13182 & ~pi285;
assign w20466 = ~pi234 & ~pi285;
assign w20467 = ~pi234 & w19550;
assign w20468 = pi149 & ~pi234;
assign w20469 = pi149 & w19559;
assign w20470 = pi284 & w19562;
assign w20471 = ~pi193 & pi284;
assign w20472 = ~pi193 & w19564;
assign w20473 = ~w13838 & pi193;
assign w20474 = ~pi386 & pi193;
assign w20475 = ~pi386 & ~w19567;
assign w20476 = pi386 & ~pi193;
assign w20477 = pi386 & w19567;
assign w20478 = ~pi135 & pi193;
assign w20479 = ~pi135 & ~w19567;
assign w20480 = pi135 & ~pi193;
assign w20481 = pi135 & w19567;
assign w20482 = w14030 & pi372;
assign w20483 = w13549 & ~pi144;
assign w20484 = ~w13549 & pi144;
assign w20485 = pi302 & ~pi139;
assign w20486 = w14232 & pi302;
assign w20487 = ~pi178 & pi139;
assign w20488 = (~pi178 & w14223) | (~pi178 & w20745) | (w14223 & w20745);
assign w20489 = pi178 & ~pi139;
assign w20490 = ~w14223 & w20746;
assign w20491 = ~w14447 & w14363;
assign w20492 = w14447 & ~w14363;
assign w20493 = ~pi351 & ~pi284;
assign w20494 = ~pi148 & pi234;
assign w20495 = ~pi148 & ~w19559;
assign w20496 = pi148 & ~pi234;
assign w20497 = pi148 & w19559;
assign w20498 = ~w14692 & w20747;
assign w20499 = (~w14687 & w14692) | (~w14687 & w20748) | (w14692 & w20748);
assign w20500 = ~w13908 & pi191;
assign w20501 = pi270 & ~pi234;
assign w20502 = pi231 & ~pi234;
assign w20503 = pi231 & w19703;
assign w20504 = (~pi192 & w14952) | (~pi192 & w20749) | (w14952 & w20749);
assign w20505 = ~w14952 & w20750;
assign w20506 = w15145 & w15156;
assign w20507 = w15169 & pi234;
assign w20508 = w15169 & ~w19559;
assign w20509 = ~pi167 & pi139;
assign w20510 = (~pi167 & w14223) | (~pi167 & w20751) | (w14223 & w20751);
assign w20511 = pi167 & ~pi139;
assign w20512 = ~w14223 & w20752;
assign w20513 = w15433 & ~pi285;
assign w20514 = (pi234 & ~w15441) | (pi234 & w20753) | (~w15441 & w20753);
assign w20515 = ~w15497 & pi139;
assign w20516 = ~w15568 & ~pi139;
assign w20517 = ~w14223 & w20754;
assign w20518 = w15568 & pi139;
assign w20519 = w15568 & ~w19622;
assign w20520 = ~w13190 & ~pi234;
assign w20521 = w15424 & pi285;
assign w20522 = ~w14008 & w14743;
assign w20523 = ~pi141 & ~pi044;
assign w20524 = ~pi141 & ~w19167;
assign w20525 = pi141 & pi044;
assign w20526 = pi141 & w19167;
assign w20527 = ~w14447 & ~pi181;
assign w20528 = w14447 & pi181;
assign w20529 = ~w14447 & ~w15858;
assign w20530 = w14447 & w15858;
assign w20531 = pi129 & pi207;
assign w20532 = ~pi036 & ~pi144;
assign w20533 = pi036 & pi144;
assign w20534 = ~pi140 & ~pi029;
assign w20535 = ~pi140 & ~w18744;
assign w20536 = pi140 & pi029;
assign w20537 = pi140 & w18744;
assign w20538 = ~w14954 & ~pi189;
assign w20539 = w14954 & pi189;
assign w20540 = w14954 & ~w16081;
assign w20541 = ~w14954 & w16081;
assign w20542 = ~pi006 & pi167;
assign w20543 = ~pi354 & ~pi351;
assign w20544 = ~pi150 & ~pi012;
assign w20545 = ~pi150 & ~w18879;
assign w20546 = pi150 & pi012;
assign w20547 = pi150 & w18879;
assign w20548 = w16258 & pi234;
assign w20549 = ~w13298 & pi285;
assign w20550 = w14204 & pi302;
assign w20551 = ~pi139 & w16381;
assign w20552 = pi139 & ~w16381;
assign w20553 = w15459 & pi285;
assign w20554 = ~pi270 & ~pi215;
assign w20555 = w14699 & ~pi222;
assign w20556 = ~w14699 & pi222;
assign w20557 = w14699 & ~w16606;
assign w20558 = ~w14699 & w16606;
assign w20559 = ~pi129 & ~pi018;
assign w20560 = ~pi129 & ~w19314;
assign w20561 = pi129 & pi018;
assign w20562 = pi129 & w19314;
assign w20563 = ~pi121 & ~pi020;
assign w20564 = ~pi121 & ~w18435;
assign w20565 = pi121 & pi020;
assign w20566 = pi121 & w18435;
assign w20567 = ~w8060 & ~pi179;
assign w20568 = w8060 & pi179;
assign w20569 = ~pi225 & ~pi060;
assign w20570 = ~pi225 & ~w18640;
assign w20571 = pi225 & pi060;
assign w20572 = pi225 & w18640;
assign w20573 = ~w9377 & ~pi226;
assign w20574 = w9377 & pi226;
assign w20575 = ~pi132 & ~pi017;
assign w20576 = ~pi132 & ~w18289;
assign w20577 = pi132 & pi017;
assign w20578 = pi132 & w18289;
assign w20579 = ~pi156 & pi078;
assign w20580 = ~pi156 & ~w17904;
assign w20581 = pi156 & ~pi078;
assign w20582 = pi156 & w17904;
assign w20583 = pi078 & ~pi151;
assign w20584 = ~pi078 & pi151;
assign w20585 = pi138 & ~pi302;
assign w20586 = w15882 & ~pi302;
assign w20587 = ~w16812 & pi139;
assign w20588 = ~pi370 & ~pi139;
assign w20589 = ~pi370 & ~w19989;
assign w20590 = pi370 & pi139;
assign w20591 = pi370 & w19989;
assign w20592 = pi193 & pi017;
assign w20593 = pi193 & w18419;
assign w20594 = pi012 & ~pi142;
assign w20595 = ~pi012 & pi142;
assign w20596 = ~pi143 & ~pi012;
assign w20597 = ~pi143 & ~w17974;
assign w20598 = pi143 & pi012;
assign w20599 = pi143 & w17974;
assign w20600 = w16929 & pi193;
assign w20601 = ~pi162 & ~pi036;
assign w20602 = ~pi162 & ~w18109;
assign w20603 = pi162 & pi036;
assign w20604 = pi162 & w18109;
assign w20605 = pi030 & ~pi149;
assign w20606 = ~pi030 & pi149;
assign w20607 = ~pi134 & ~pi044;
assign w20608 = ~pi134 & ~w18557;
assign w20609 = pi134 & pi044;
assign w20610 = pi134 & w18557;
assign w20611 = ~pi346 & ~pi030;
assign w20612 = ~pi346 & ~w19396;
assign w20613 = pi346 & pi030;
assign w20614 = pi346 & w19396;
assign w20615 = ~pi267 & pi029;
assign w20616 = ~pi267 & ~w18852;
assign w20617 = pi267 & ~pi029;
assign w20618 = pi267 & w18852;
assign w20619 = ~pi372 & ~pi010;
assign w20620 = ~pi372 & ~w18824;
assign w20621 = pi372 & pi010;
assign w20622 = pi372 & w18824;
assign w20623 = ~pi342 & pi010;
assign w20624 = ~pi342 & ~w18388;
assign w20625 = pi342 & ~pi010;
assign w20626 = pi342 & w18388;
assign w20627 = ~pi258 & pi012;
assign w20628 = ~pi258 & ~w17967;
assign w20629 = pi258 & ~pi012;
assign w20630 = pi258 & w17967;
assign w20631 = ~pi274 & ~pi015;
assign w20632 = ~pi274 & ~w19363;
assign w20633 = pi274 & pi015;
assign w20634 = pi274 & w19363;
assign w20635 = ~pi348 & pi015;
assign w20636 = ~pi348 & ~w18525;
assign w20637 = pi348 & ~pi015;
assign w20638 = pi348 & w18525;
assign w20639 = ~pi136 & ~pi029;
assign w20640 = ~pi136 & ~w18453;
assign w20641 = pi136 & pi029;
assign w20642 = pi136 & w18453;
assign w20643 = ~pi135 & ~pi036;
assign w20644 = ~pi135 & ~w18970;
assign w20645 = pi135 & pi036;
assign w20646 = pi135 & w18970;
assign w20647 = ~pi155 & ~pi078;
assign w20648 = ~pi155 & ~w18510;
assign w20649 = pi155 & pi078;
assign w20650 = pi155 & w18510;
assign w20651 = ~pi230 & ~pi053;
assign w20652 = ~pi230 & ~w18534;
assign w20653 = pi230 & pi053;
assign w20654 = pi230 & w18534;
assign w20655 = ~w3637 & ~pi166;
assign w20656 = w3637 & pi166;
assign w20657 = ~pi275 & ~pi017;
assign w20658 = ~pi275 & ~w19233;
assign w20659 = pi275 & pi017;
assign w20660 = pi275 & w19233;
assign w20661 = ~pi370 & pi006;
assign w20662 = ~pi370 & ~w18597;
assign w20663 = pi370 & ~pi006;
assign w20664 = pi370 & w18597;
assign w20665 = ~pi175 & ~pi068;
assign w20666 = ~pi175 & ~w18360;
assign w20667 = pi175 & pi068;
assign w20668 = pi175 & w18360;
assign w20669 = ~pi138 & ~pi018;
assign w20670 = ~pi138 & ~w18301;
assign w20671 = pi138 & pi018;
assign w20672 = pi138 & w18301;
assign w20673 = ~pi139 & ~pi349;
assign w20674 = pi139 & pi349;
assign w20675 = ~pi139 & ~w17332;
assign w20676 = pi139 & w17332;
assign w20677 = pi171 & pi060;
assign w20678 = pi171 & w19205;
assign w20679 = ~pi271 & ~pi038;
assign w20680 = ~pi271 & ~w19171;
assign w20681 = pi271 & pi038;
assign w20682 = pi271 & w19171;
assign w20683 = ~pi273 & pi030;
assign w20684 = ~pi273 & ~w19346;
assign w20685 = pi273 & ~pi030;
assign w20686 = pi273 & w19346;
assign w20687 = ~pi173 & pi020;
assign w20688 = ~pi173 & ~w18064;
assign w20689 = pi173 & ~pi020;
assign w20690 = pi173 & w18064;
assign w20691 = ~pi234 & ~pi068;
assign w20692 = ~pi234 & ~w18407;
assign w20693 = pi234 & pi068;
assign w20694 = pi234 & w18407;
assign w20695 = w20147 & pi012;
assign w20696 = w7824 & pi017;
assign w20697 = w3862 & pi018;
assign w20698 = w20219 & pi029;
assign w20699 = w5058 & pi020;
assign w20700 = ~pi121 & ~w20145;
assign w20701 = ~pi121 & ~w20148;
assign w20702 = pi121 & w20145;
assign w20703 = pi121 & w20148;
assign w20704 = pi190 & w20237;
assign w20705 = pi190 & w20238;
assign w20706 = pi136 & w20145;
assign w20707 = pi136 & w20148;
assign w20708 = w5996 & pi044;
assign w20709 = w18604 & pi006;
assign w20710 = pi040 & ~pi142;
assign w20711 = ~pi040 & pi142;
assign w20712 = w498 & ~pi029;
assign w20713 = pi007 & ~pi001;
assign w20714 = w17964 & ~pi012;
assign w20715 = pi115 & ~pi030;
assign w20716 = w20335 & pi036;
assign w20717 = pi089 & ~pi178;
assign w20718 = ~pi089 & pi178;
assign w20719 = pi118 & pi038;
assign w20720 = pi058 & ~pi060;
assign w20721 = pi058 & w19190;
assign w20722 = w20368 & pi060;
assign w20723 = pi065 & w19281;
assign w20724 = w3560 & w11392;
assign w20725 = pi115 & pi030;
assign w20726 = pi080 & pi015;
assign w20727 = w20407 & pi146;
assign w20728 = w20407 & pi273;
assign w20729 = ~pi181 & ~w20271;
assign w20730 = ~pi181 & ~w20369;
assign w20731 = pi181 & w20271;
assign w20732 = pi181 & w20369;
assign w20733 = ~w20407 & ~pi227;
assign w20734 = w20407 & pi227;
assign w20735 = ~pi163 & ~w20237;
assign w20736 = ~pi163 & ~w20238;
assign w20737 = pi163 & w20237;
assign w20738 = pi163 & w20238;
assign w20739 = ~w20407 & ~pi348;
assign w20740 = w20407 & pi348;
assign w20741 = ~pi228 & ~w20237;
assign w20742 = ~pi228 & ~w20238;
assign w20743 = pi228 & w20237;
assign w20744 = pi228 & w20238;
assign w20745 = ~w20485 & ~pi178;
assign w20746 = w20485 & pi178;
assign w20747 = w14698 & w14687;
assign w20748 = ~w14698 & ~w14687;
assign w20749 = w14953 & ~pi192;
assign w20750 = ~w14953 & pi192;
assign w20751 = ~w20485 & ~pi167;
assign w20752 = w20485 & pi167;
assign w20753 = w13669 & pi234;
assign w20754 = w20485 & ~w15568;
assign w20755 = ~w101 & ~w144;
assign w20756 = w1078 & ~pi123;
assign w20757 = w1068 & pi048;
assign w20758 = w1156 & ~w1157;
assign w20759 = w499 & ~pi114;
assign w20760 = w1199 & ~pi001;
assign w20761 = w1199 & ~w18019;
assign w20762 = w1301 & pi040;
assign w20763 = ~w1705 & pi115;
assign w20764 = w2544 & w2499;
assign w20765 = ~w2908 & pi034;
assign w20766 = ~pi018 & ~w3616;
assign w20767 = ~w4343 & ~pi017;
assign w20768 = w4517 & pi106;
assign w20769 = w4518 & pi065;
assign w20770 = w4616 & pi113;
assign w20771 = w4617 & pi096;
assign w20772 = w4630 & pi009;
assign w20773 = w18379 | ~pi010;
assign w20774 = (~pi010 & w18379) | (~pi010 & ~w4582) | (w18379 & ~w4582);
assign w20775 = ~w4640 & ~pi138;
assign w20776 = w4640 & pi138;
assign w20777 = w3558 & pi091;
assign w20778 = w4754 & ~pi024;
assign w20779 = w4760 & pi018;
assign w20780 = ~w5315 & w5316;
assign w20781 = w5428 & pi029;
assign w20782 = w5721 & pi015;
assign w20783 = w18543 | ~pi053;
assign w20784 = (~pi053 & w18543) | (~pi053 & w5843) | (w18543 & w5843);
assign w20785 = ~w6080 & w6081;
assign w20786 = w6138 & ~pi118;
assign w20787 = ~pi086 & ~pi090;
assign w20788 = ~w6386 & ~pi088;
assign w20789 = w6396 & pi006;
assign w20790 = w6651 & ~pi034;
assign w20791 = w18649 & ~w6707;
assign w20792 = (~w6707 & w18649) | (~w6707 & ~w6699) | (w18649 & ~w6699);
assign w20793 = w3207 & ~pi090;
assign w20794 = w6371 & pi088;
assign w20795 = ~w6898 & w6905;
assign w20796 = ~w6906 & pi006;
assign w20797 = ~w7025 & ~pi096;
assign w20798 = ~w7025 & ~w18696;
assign w20799 = w7178 & ~pi035;
assign w20800 = pi065 & ~w4098;
assign w20801 = w7148 & pi068;
assign w20802 = ~w7631 & ~w7637;
assign w20803 = ~w7638 & pi012;
assign w20804 = ~w7658 & ~w901;
assign w20805 = w7658 & w901;
assign w20806 = ~w7219 & ~pi358;
assign w20807 = w7219 & pi358;
assign w20808 = w7737 & ~w7753;
assign w20809 = w7791 & pi039;
assign w20810 = ~w8054 & ~w8055;
assign w20811 = w8056 & w8072;
assign w20812 = w8056 & w18843;
assign w20813 = w18844 & pi142;
assign w20814 = (pi142 & w18844) | (pi142 & ~w8056) | (w18844 & ~w8056);
assign w20815 = ~pi106 & ~w7194;
assign w20816 = w8197 & ~pi068;
assign w20817 = ~w4640 & ~pi132;
assign w20818 = w4640 & pi132;
assign w20819 = w8395 & ~pi092;
assign w20820 = pi087 & pi046;
assign w20821 = w8513 & pi092;
assign w20822 = w8514 & pi089;
assign w20823 = w18944 | pi015;
assign w20824 = (pi015 & w18944) | (pi015 & ~w8754) | (w18944 & ~w8754);
assign w20825 = w1665 & ~pi061;
assign w20826 = w9142 & ~w9146;
assign w20827 = w2157 & ~pi092;
assign w20828 = ~w19033 & ~pi036;
assign w20829 = ~w9540 & w9541;
assign w20830 = ~w9542 & ~w8519;
assign w20831 = pi073 & w2295;
assign w20832 = pi073 & ~w19060;
assign w20833 = ~w9599 & w9615;
assign w20834 = w9721 & pi073;
assign w20835 = ~w10224 & ~w10225;
assign w20836 = ~w10226 & pi006;
assign w20837 = ~pi003 & w5954;
assign w20838 = ~pi003 & ~w19179;
assign w20839 = w10480 & ~w10481;
assign w20840 = ~pi272 & w10525;
assign w20841 = ~pi272 & w10482;
assign w20842 = pi272 & ~w10525;
assign w20843 = pi272 & ~w10482;
assign w20844 = ~w10532 & ~pi529;
assign w20845 = w10583 & ~pi034;
assign w20846 = ~w6397 & ~pi130;
assign w20847 = w6397 & pi130;
assign w20848 = w10819 & ~pi039;
assign w20849 = w11156 & ~w11158;
assign w20850 = ~pi275 & w11194;
assign w20851 = ~pi275 & w11159;
assign w20852 = pi275 & ~w11194;
assign w20853 = pi275 & ~w11159;
assign w20854 = w11201 & ~pi529;
assign w20855 = w11394 & ~w11419;
assign w20856 = ~w488 & ~w7362;
assign w20857 = ~w11474 & pi114;
assign w20858 = w11475 & pi029;
assign w20859 = ~w11539 & ~pi529;
assign w20860 = ~w1723 & ~pi115;
assign w20861 = ~w11711 & w11713;
assign w20862 = w11836 & ~w11842;
assign w20863 = ~w11843 & pi036;
assign w20864 = w1665 & pi002;
assign w20865 = ~pi274 & w11749;
assign w20866 = ~pi274 & w11716;
assign w20867 = pi274 & ~w11749;
assign w20868 = pi274 & ~w11716;
assign w20869 = ~w11916 & ~pi529;
assign w20870 = ~w11991 & ~pi030;
assign w20871 = ~w8808 & ~pi131;
assign w20872 = w8808 & pi131;
assign w20873 = pi002 & w9301;
assign w20874 = pi002 & ~w19403;
assign w20875 = ~w12087 & w12088;
assign w20876 = ~w8808 & ~pi135;
assign w20877 = w8808 & pi135;
assign w20878 = w12173 & ~pi529;
assign w20879 = ~w6397 & ~pi134;
assign w20880 = w6397 & pi134;
assign w20881 = w12746 & ~pi529;
assign w20882 = ~w1366 & ~pi257;
assign w20883 = w1366 & pi257;
assign w20884 = w9147 & ~pi357;
assign w20885 = ~w9147 & pi357;
assign w20886 = w9550 & ~pi350;
assign w20887 = ~w9550 & pi350;
assign w20888 = ~w12905 & ~pi529;
assign w20889 = w9616 & ~pi229;
assign w20890 = ~w9616 & pi229;
assign w20891 = w12936 & ~pi529;
assign w20892 = ~pi276 & w11194;
assign w20893 = ~pi276 & w11159;
assign w20894 = pi276 & ~w11194;
assign w20895 = pi276 & ~w11159;
assign w20896 = w13039 & ~pi529;
assign w20897 = w9616 & ~pi346;
assign w20898 = ~w9616 & pi346;
assign w20899 = w13137 & ~pi529;
assign w20900 = w13450 & ~pi529;
assign w20901 = ~pi232 & ~pi231;
assign w20902 = w14205 & pi207;
assign w20903 = w13593 & w15973;
assign w20904 = w16001 & w16006;
assign w20905 = w16131 & ~pi284;
assign w20906 = w16160 & ~pi284;
assign w20907 = w16134 & pi193;
assign w20908 = w16185 & w16189;
assign w20909 = ~w16185 & ~w16189;
assign w20910 = ~w16393 & ~w16401;
assign w20911 = ~pi353 & w16449;
assign w20912 = ~pi353 & w16404;
assign w20913 = pi353 & ~w16449;
assign w20914 = pi353 & ~w16404;
assign w20915 = w16764 & ~w16766;
assign w20916 = pi102 & w17975;
assign w20917 = ~pi012 & pi102;
assign w20918 = ~pi012 & w17977;
assign w20919 = pi039 & w18290;
assign w20920 = ~pi017 & w18291;
assign w20921 = pi024 & w18302;
assign w20922 = ~pi018 & w18304;
assign w20923 = pi065 & w18361;
assign w20924 = ~pi068 & w18362;
assign w20925 = pi048 & w18436;
assign w20926 = ~pi020 & w18438;
assign w20927 = ~pi054 & pi114;
assign w20928 = pi001 & w18448;
assign w20929 = ~pi029 & w18449;
assign w20930 = pi003 & w18549;
assign w20931 = ~pi044 & w18550;
assign w20932 = ~pi058 & w18586;
assign w20933 = pi031 & w7900;
assign w20934 = w1919 & pi002;
assign w20935 = ~pi036 & w18971;
assign w20936 = w2533 & pi003;
assign w20937 = pi058 & w19206;
assign w20938 = ~pi060 & w19207;
assign w20939 = w4767 & pi024;
assign w20940 = ~w4498 & ~pi106;
assign w20941 = ~pi003 & ~w5945;
assign w20942 = ~pi003 & w9876;
assign w20943 = pi044 & w19426;
assign w20944 = pi065 & ~w19283;
assign w20945 = pi065 & w8201;
assign w20946 = ~w11182 & w11193;
assign one = 1;
assign po000 = pi397;// level 0
assign po001 = pi211;// level 0
assign po002 = pi305;// level 0
assign po003 = pi339;// level 0
assign po004 = pi345;// level 0
assign po005 = pi212;// level 0
assign po006 = pi262;// level 0
assign po007 = pi213;// level 0
assign po008 = pi306;// level 0
assign po009 = pi383;// level 0
assign po010 = pi322;// level 0
assign po011 = pi206;// level 0
assign po012 = pi336;// level 0
assign po013 = pi158;// level 0
assign po014 = pi241;// level 0
assign po015 = pi332;// level 0
assign po016 = pi331;// level 0
assign po017 = pi261;// level 0
assign po018 = pi381;// level 0
assign po019 = pi296;// level 0
assign po020 = pi243;// level 0
assign po021 = pi374;// level 0
assign po022 = pi259;// level 0
assign po023 = pi329;// level 0
assign po024 = pi295;// level 0
assign po025 = pi288;// level 0
assign po026 = pi341;// level 0
assign po027 = pi365;// level 0
assign po028 = pi338;// level 0
assign po029 = pi340;// level 0
assign po030 = pi235;// level 0
assign po031 = pi294;// level 0
assign po032 = pi323;// level 0
assign po033 = pi214;// level 0
assign po034 = pi309;// level 0
assign po035 = pi337;// level 0
assign po036 = pi264;// level 0
assign po037 = pi308;// level 0
assign po038 = pi263;// level 0
assign po039 = pi307;// level 0
assign po040 = pi310;// level 0
assign po041 = pi317;// level 0
assign po042 = pi304;// level 0
assign po043 = pi245;// level 0
assign po044 = pi196;// level 0
assign po045 = pi177;// level 0
assign po046 = pi237;// level 0
assign po047 = pi204;// level 0
assign po048 = pi244;// level 0
assign po049 = pi201;// level 0
assign po050 = pi382;// level 0
assign po051 = pi314;// level 0
assign po052 = pi236;// level 0
assign po053 = pi367;// level 0
assign po054 = pi282;// level 0
assign po055 = pi326;// level 0
assign po056 = pi325;// level 0
assign po057 = pi277;// level 0
assign po058 = pi298;// level 0
assign po059 = pi343;// level 0
assign po060 = pi315;// level 0
assign po061 = pi300;// level 0
assign po062 = pi188;// level 0
assign po063 = pi249;// level 0
assign po064 = pi360;// level 0
assign po065 = pi216;// level 0
assign po066 = pi347;// level 0
assign po067 = pi335;// level 0
assign po068 = pi266;// level 0
assign po069 = pi311;// level 0
assign po070 = pi265;// level 0
assign po071 = pi312;// level 0
assign po072 = pi313;// level 0
assign po073 = pi318;// level 0
assign po074 = pi291;// level 0
assign po075 = pi247;// level 0
assign po076 = pi289;// level 0
assign po077 = pi199;// level 0
assign po078 = pi240;// level 0
assign po079 = pi252;// level 0
assign po080 = pi246;// level 0
assign po081 = pi202;// level 0
assign po082 = pi378;// level 0
assign po083 = pi293;// level 0
assign po084 = pi287;// level 0
assign po085 = pi368;// level 0
assign po086 = pi286;// level 0
assign po087 = pi377;// level 0
assign po088 = pi380;// level 0
assign po089 = pi279;// level 0
assign po090 = pi299;// level 0
assign po091 = pi327;// level 0
assign po092 = pi316;// level 0
assign po093 = pi333;// level 0
assign po094 = pi186;// level 0
assign po095 = pi250;// level 0
assign po096 = pi369;// level 0
assign po097 = pi361;// level 0
assign po098 = pi359;// level 0
assign po099 = pi366;// level 0
assign po100 = pi379;// level 0
assign po101 = pi248;// level 0
assign po102 = pi194;// level 0
assign po103 = pi324;// level 0
assign po104 = pi330;// level 0
assign po105 = pi239;// level 0
assign po106 = pi238;// level 0
assign po107 = pi292;// level 0
assign po108 = pi355;// level 0
assign po109 = pi195;// level 0
assign po110 = pi197;// level 0
assign po111 = pi251;// level 0
assign po112 = pi200;// level 0
assign po113 = pi203;// level 0
assign po114 = pi362;// level 0
assign po115 = pi297;// level 0
assign po116 = pi242;// level 0
assign po117 = pi334;// level 0
assign po118 = pi198;// level 0
assign po119 = pi364;// level 0
assign po120 = pi328;// level 0
assign po121 = pi260;// level 0
assign po122 = pi253;// level 0
assign po123 = pi344;// level 0
assign po124 = pi290;// level 0
assign po125 = pi254;// level 0
assign po126 = pi176;// level 0
assign po127 = pi205;// level 0
assign po128 = pi363;// level 0
assign po129 = pi530;// level 0
assign po130 = w915;// level 18
assign po131 = ~w1542;// level 18
assign po132 = ~w2446;// level 18
assign po133 = ~w3368;// level 18
assign po134 = w4291;// level 18
assign po135 = w4656;// level 18
assign po136 = ~w4999;// level 17
assign po137 = w5261;// level 18
assign po138 = w5416;// level 18
assign po139 = w5572;// level 18
assign po140 = one;// level 0
assign po141 = w5657;// level 16
assign po142 = pi529;// level 0
assign po143 = ~w5660;// level 2
assign po144 = w5680;// level 18
assign po145 = ~w5887;// level 16
assign po146 = w5890;// level 2
assign po147 = w5914;// level 18
assign po148 = w6545;// level 18
assign po149 = w6633;// level 16
assign po150 = ~w6636;// level 2
assign po151 = w6884;// level 18
assign po152 = ~w6968;// level 17
assign po153 = ~w7048;// level 17
assign po154 = w7141;// level 18
assign po155 = ~w7237;// level 17
assign po156 = w7590;// level 17
assign po157 = ~w7669;// level 18
assign po158 = w7770;// level 18
assign po159 = ~w8007;// level 18
assign po160 = ~w8088;// level 18
assign po161 = ~w8173;// level 18
assign po162 = w8259;// level 18
assign po163 = w8283;// level 18
assign po164 = ~w8355;// level 17
assign po165 = ~w8375;// level 17
assign po166 = w8913;// level 18
assign po167 = ~w9166;// level 18
assign po168 = ~w9407;// level 18
assign po169 = ~w9495;// level 18
assign po170 = w9632;// level 18
assign po171 = ~w9715;// level 17
assign po172 = ~w9797;// level 18
assign po173 = ~w9817;// level 17
assign po174 = ~w9915;// level 18
assign po175 = ~w9939;// level 18
assign po176 = w10260;// level 17
assign po177 = ~w10540;// level 17
assign po178 = w10680;// level 18
assign po179 = ~w10694;// level 17
assign po180 = w10711;// level 17
assign po181 = w11059;// level 18
assign po182 = w11209;// level 17
assign po183 = ~w11298;// level 18
assign po184 = w11322;// level 18
assign po185 = w11339;// level 17
assign po186 = w11357;// level 18
assign po187 = w11437;// level 17
assign po188 = w11454;// level 17
assign po189 = ~w11471;// level 17
assign po190 = ~w11547;// level 17
assign po191 = w11561;// level 18
assign po192 = ~w11578;// level 17
assign po193 = ~w11601;// level 18
assign po194 = w11624;// level 18
assign po195 = w11641;// level 17
assign po196 = ~w11824;// level 17
assign po197 = w11904;// level 18
assign po198 = ~w11924;// level 17
assign po199 = w11938;// level 18
assign po200 = ~w11964;// level 18
assign po201 = ~w12043;// level 18
assign po202 = ~w12124;// level 18
assign po203 = w12141;// level 17
assign po204 = w12164;// level 18
assign po205 = w12181;// level 17
assign po206 = ~w12201;// level 18
assign po207 = ~w12218;// level 18
assign po208 = ~w12236;// level 18
assign po209 = w12316;// level 18
assign po210 = w12337;// level 18
assign po211 = w12361;// level 18
assign po212 = w12441;// level 18
assign po213 = w12455;// level 17
assign po214 = w12476;// level 18
assign po215 = w12497;// level 18
assign po216 = w12514;// level 18
assign po217 = w12532;// level 18
assign po218 = w12550;// level 18
assign po219 = ~w12564;// level 17
assign po220 = w12582;// level 18
assign po221 = ~w12599;// level 18
assign po222 = ~w12616;// level 18
assign po223 = ~w12640;// level 18
assign po224 = ~w12658;// level 18
assign po225 = ~w12676;// level 18
assign po226 = w12690;// level 17
assign po227 = w12708;// level 18
assign po228 = w12723;// level 18
assign po229 = w12737;// level 17
assign po230 = w12754;// level 17
assign po231 = ~w12772;// level 18
assign po232 = w12789;// level 17
assign po233 = w12803;// level 17
assign po234 = w12820;// level 18
assign po235 = w12837;// level 17
assign po236 = ~w12855;// level 18
assign po237 = ~w12872;// level 18
assign po238 = w12896;// level 18
assign po239 = ~w12913;// level 17
assign po240 = ~w12927;// level 17
assign po241 = w12944;// level 17
assign po242 = w12962;// level 18
assign po243 = w12979;// level 17
assign po244 = w12994;// level 18
assign po245 = w13012;// level 18
assign po246 = w13030;// level 18
assign po247 = w13047;// level 17
assign po248 = ~w13064;// level 17
assign po249 = w13078;// level 17
assign po250 = w13096;// level 18
assign po251 = w13114;// level 18
assign po252 = ~w13128;// level 17
assign po253 = w13145;// level 17
assign po254 = w13159;// level 18
assign po255 = w13176;// level 17
assign po256 = ~w13333;// level 15
assign po257 = w13348;// level 18
assign po258 = w13366;// level 18
assign po259 = w13383;// level 17
assign po260 = w13404;// level 18
assign po261 = w13421;// level 17
assign po262 = w13441;// level 18
assign po263 = w13458;// level 17
assign po264 = ~w13636;// level 16
assign po265 = w13642;// level 13
assign po266 = ~w13648;// level 15
assign po267 = ~w13660;// level 13
assign po268 = ~w13774;// level 16
assign po269 = ~w13873;// level 15
assign po270 = ~w13882;// level 15
assign po271 = ~w13897;// level 15
assign po272 = ~w14058;// level 13
assign po273 = ~w14070;// level 15
assign po274 = ~w14168;// level 16
assign po275 = ~w14180;// level 16
assign po276 = w14186;// level 16
assign po277 = ~w14357;// level 16
assign po278 = ~w14466;// level 13
assign po279 = w14469;// level 16
assign po280 = pi532;// level 0
assign po281 = pi626;// level 0
assign po282 = ~w14547;// level 16
assign po283 = ~w14556;// level 16
assign po284 = ~w14571;// level 16
assign po285 = w14577;// level 14
assign po286 = ~w14583;// level 16
assign po287 = ~w14681;// level 15
assign po288 = ~w14785;// level 13
assign po289 = w14872;// level 15
assign po290 = ~w14884;// level 16
assign po291 = ~w14986;// level 15
assign po292 = ~w15073;// level 14
assign po293 = ~w15163;// level 14
assign po294 = ~w15175;// level 14
assign po295 = w15178;// level 12
assign po296 = ~w15263;// level 16
assign po297 = w15269;// level 16
assign po298 = ~w15354;// level 16
assign po299 = w15357;// level 16
assign po300 = pi621;// level 0
assign po301 = ~w15366;// level 16
assign po302 = ~w15378;// level 16
assign po303 = ~w15393;// level 16
assign po304 = ~w15405;// level 16
assign po305 = w15411;// level 14
assign po306 = ~w15486;// level 13
assign po307 = ~w15562;// level 14
assign po308 = ~w15574;// level 14
assign po309 = w15580;// level 13
assign po310 = ~w15586;// level 15
assign po311 = ~w15666;// level 13
assign po312 = ~w15743;// level 14
assign po313 = ~w15752;// level 13
assign po314 = w15755;// level 12
assign po315 = w15758;// level 12
assign po316 = ~w15764;// level 16
assign po317 = ~w15843;// level 16
assign po318 = ~w15852;// level 15
assign po319 = w15855;// level 13
assign po320 = ~w15864;// level 13
assign po321 = ~w15948;// level 14
assign po322 = ~w16024;// level 16
assign po323 = ~w16033;// level 18
assign po324 = w16036;// level 12
assign po325 = w16042;// level 13
assign po326 = ~w16045;// level 12
assign po327 = w16051;// level 13
assign po328 = ~w16057;// level 15
assign po329 = ~w16069;// level 13
assign po330 = ~w16075;// level 15
assign po331 = ~w16087;// level 13
assign po332 = w16090;// level 12
assign po333 = w16093;// level 12
assign po334 = w16096;// level 11
assign po335 = w16099;// level 11
assign po336 = w16102;// level 12
assign po337 = w16105;// level 12
assign po338 = w16108;// level 11
assign po339 = w16111;// level 12
assign po340 = ~w16114;// level 12
assign po341 = w16117;// level 12
assign po342 = w16120;// level 12
assign po343 = w16123;// level 12
assign po344 = w16126;// level 12
assign po345 = ~w16201;// level 17
assign po346 = w16204;// level 15
assign po347 = ~w16219;// level 16
assign po348 = ~w16222;// level 13
assign po349 = w16225;// level 12
assign po350 = w16228;// level 12
assign po351 = w16231;// level 12
assign po352 = w16234;// level 11
assign po353 = ~w16240;// level 17
assign po354 = ~w16243;// level 11
assign po355 = ~w16316;// level 13
assign po356 = ~w16387;// level 14
assign po357 = w16461;// level 15
assign po358 = ~w16537;// level 14
assign po359 = ~w16549;// level 16
assign po360 = w16555;// level 13
assign po361 = w16561;// level 14
assign po362 = w16567;// level 14
assign po363 = w16573;// level 14
assign po364 = ~w16579;// level 16
assign po365 = ~w16585;// level 15
assign po366 = ~w16591;// level 16
assign po367 = ~w16597;// level 15
assign po368 = ~w16603;// level 16
assign po369 = ~w16612;// level 13
assign po370 = ~w16624;// level 14
assign po371 = ~w16633;// level 14
assign po372 = ~w16642;// level 14
assign po373 = w16645;// level 12
assign po374 = w16648;// level 11
assign po375 = w16651;// level 12
assign po376 = w16654;// level 11
assign po377 = w16657;// level 11
assign po378 = ~w16660;// level 11
assign po379 = w16663;// level 12
assign po380 = w16666;// level 11
assign po381 = w16669;// level 11
assign po382 = w16672;// level 12
assign po383 = w16675;// level 11
assign po384 = w16678;// level 11
assign po385 = w16681;// level 12
assign po386 = w16684;// level 12
assign po387 = w16687;// level 12
assign po388 = ~w16690;// level 12
assign po389 = w16693;// level 12
assign po390 = w16696;// level 12
assign po391 = w16699;// level 12
assign po392 = w16702;// level 12
assign po393 = ~w16711;// level 16
assign po394 = ~w16714;// level 13
assign po395 = w16794;// level 16
assign po396 = w16868;// level 15
assign po397 = w16871;// level 12
assign po398 = w16874;// level 12
assign po399 = w16877;// level 11
assign po400 = w16880;// level 12
assign po401 = w16883;// level 11
assign po402 = w16886;// level 11
assign po403 = ~w16889;// level 12
assign po404 = w16892;// level 12
assign po405 = ~w16960;// level 16
assign po406 = ~w16972;// level 16
assign po407 = w16978;// level 14
assign po408 = ~w16987;// level 16
assign po409 = w16993;// level 13
assign po410 = w16999;// level 14
assign po411 = ~w17005;// level 15
assign po412 = ~w17011;// level 16
assign po413 = ~w17020;// level 13
assign po414 = ~w17029;// level 14
assign po415 = w17032;// level 12
assign po416 = w17038;// level 13
assign po417 = w17041;// level 11
assign po418 = w17047;// level 14
assign po419 = ~w17053;// level 15
assign po420 = w17056;// level 12
assign po421 = ~w17062;// level 16
assign po422 = ~w17071;// level 13
assign po423 = ~w17080;// level 14
assign po424 = ~w17083;// level 12
assign po425 = ~w17086;// level 12
assign po426 = w17089;// level 12
assign po427 = w17092;// level 11
assign po428 = w17095;// level 11
assign po429 = w17098;// level 11
assign po430 = w17101;// level 12
assign po431 = w17104;// level 11
assign po432 = w17107;// level 12
assign po433 = w17110;// level 11
assign po434 = w17113;// level 12
assign po435 = w17116;// level 12
assign po436 = w17119;// level 11
assign po437 = ~w17122;// level 12
assign po438 = w17125;// level 11
assign po439 = ~w17131;// level 16
assign po440 = ~w17143;// level 16
assign po441 = ~w17149;// level 16
assign po442 = w17152;// level 12
assign po443 = w17155;// level 11
assign po444 = w17158;// level 11
assign po445 = w17161;// level 11
assign po446 = w17164;// level 12
assign po447 = w17167;// level 11
assign po448 = w17170;// level 11
assign po449 = w17173;// level 11
assign po450 = w17176;// level 11
assign po451 = w17179;// level 11
assign po452 = w17182;// level 12
assign po453 = w17185;// level 11
assign po454 = ~w17188;// level 11
assign po455 = w17191;// level 11
assign po456 = w17194;// level 11
assign po457 = w17200;// level 14
assign po458 = ~w17206;// level 16
assign po459 = ~w17215;// level 14
assign po460 = w17218;// level 11
assign po461 = w17221;// level 11
assign po462 = w17224;// level 12
assign po463 = w17227;// level 11
assign po464 = w17230;// level 12
assign po465 = ~w17233;// level 12
assign po466 = w17236;// level 11
assign po467 = w17239;// level 11
assign po468 = w17242;// level 11
assign po469 = w17245;// level 12
assign po470 = w17248;// level 12
assign po471 = ~w17251;// level 12
assign po472 = w17254;// level 12
assign po473 = w17257;// level 12
assign po474 = w17260;// level 11
assign po475 = w17263;// level 12
assign po476 = w17266;// level 11
assign po477 = w17269;// level 12
assign po478 = w17272;// level 12
assign po479 = w17275;// level 12
assign po480 = ~w17281;// level 17
assign po481 = w17284;// level 12
assign po482 = w17287;// level 12
assign po483 = w17290;// level 12
assign po484 = ~w17299;// level 15
assign po485 = w17302;// level 11
assign po486 = ~w17308;// level 15
assign po487 = w17314;// level 14
assign po488 = ~w17320;// level 16
assign po489 = ~w17329;// level 13
assign po490 = ~w17338;// level 14
assign po491 = ~w17341;// level 13
assign po492 = ~w17347;// level 17
assign po493 = w17350;// level 11
assign po494 = w17356;// level 14
assign po495 = ~w17362;// level 16
assign po496 = ~w17371;// level 14
assign po497 = w17374;// level 12
assign po498 = w17377;// level 11
assign po499 = w17380;// level 12
assign po500 = w17383;// level 12
assign po501 = w17386;// level 11
assign po502 = w17389;// level 11
assign po503 = w17392;// level 11
assign po504 = w17395;// level 12
assign po505 = w17398;// level 12
assign po506 = w17401;// level 11
assign po507 = ~w17404;// level 11
assign po508 = ~w17407;// level 13
assign po509 = w17410;// level 13
assign po510 = ~w17416;// level 18
assign po511 = ~w17422;// level 16
assign po512 = w17425;// level 12
assign po513 = ~w17431;// level 15
assign po514 = ~w17434;// level 14
assign po515 = w17437;// level 11
assign po516 = w17440;// level 12
assign po517 = w17443;// level 12
assign po518 = w17446;// level 11
assign po519 = w17449;// level 12
assign po520 = w17452;// level 11
assign po521 = w17455;// level 11
assign po522 = w17470;// level 7
assign po523 = w17473;// level 6
assign po524 = w17478;// level 6
assign po525 = w17482;// level 4
assign po526 = w17483;// level 7
assign po527 = w17476;// level 5
assign po528 = w17488;// level 4
assign po529 = w17491;// level 6
assign po530 = w17492;// level 6
assign po531 = w17498;// level 4
assign po532 = ~w17499;// level 3
assign po533 = w17503;// level 4
assign po534 = w17505;// level 4
assign po535 = w17507;// level 3
assign po536 = ~w17510;// level 2
assign po537 = ~w17513;// level 2
assign po538 = ~w17516;// level 2
assign po539 = ~w17519;// level 2
assign po540 = ~w17522;// level 2
assign po541 = ~w17525;// level 2
assign po542 = ~w17528;// level 2
assign po543 = ~w17531;// level 2
assign po544 = ~w17534;// level 2
assign po545 = ~w17537;// level 2
assign po546 = ~w17540;// level 2
assign po547 = ~w17543;// level 2
assign po548 = ~w17546;// level 2
assign po549 = ~w17549;// level 2
assign po550 = ~w17552;// level 2
assign po551 = ~w17555;// level 2
assign po552 = ~w17558;// level 2
assign po553 = ~w17561;// level 2
assign po554 = ~w17564;// level 2
assign po555 = ~w17567;// level 2
assign po556 = ~w17570;// level 2
assign po557 = ~w17573;// level 2
assign po558 = ~w17576;// level 2
assign po559 = ~w17579;// level 2
assign po560 = ~w17582;// level 2
assign po561 = ~w17585;// level 2
assign po562 = ~w17588;// level 2
assign po563 = ~w17591;// level 2
assign po564 = ~w17594;// level 2
assign po565 = ~w17597;// level 2
assign po566 = ~w17600;// level 2
assign po567 = ~w17603;// level 2
assign po568 = ~w17606;// level 2
assign po569 = ~w17609;// level 2
assign po570 = ~w17612;// level 2
assign po571 = ~w17615;// level 2
assign po572 = ~w17618;// level 2
assign po573 = ~w17621;// level 2
assign po574 = ~w17624;// level 2
assign po575 = ~w17627;// level 2
assign po576 = ~w17630;// level 2
assign po577 = ~w17633;// level 2
assign po578 = ~w17636;// level 2
assign po579 = ~w17639;// level 2
assign po580 = ~w17642;// level 2
assign po581 = ~w17645;// level 2
assign po582 = ~w17648;// level 2
assign po583 = ~w17651;// level 2
assign po584 = ~w17654;// level 2
assign po585 = ~w17657;// level 2
assign po586 = ~w17660;// level 2
assign po587 = ~w17663;// level 2
assign po588 = ~w17666;// level 2
assign po589 = ~w17669;// level 2
assign po590 = ~w17672;// level 2
assign po591 = ~w17675;// level 2
assign po592 = ~w17678;// level 2
assign po593 = ~w17681;// level 2
assign po594 = ~w17684;// level 2
assign po595 = ~w17687;// level 2
assign po596 = ~w17690;// level 2
assign po597 = ~w17693;// level 2
assign po598 = ~w17696;// level 2
assign po599 = ~w17699;// level 2
assign po600 = ~w17702;// level 2
assign po601 = ~w17705;// level 2
assign po602 = ~w17708;// level 2
assign po603 = ~w17711;// level 2
assign po604 = ~w17714;// level 2
assign po605 = ~w17717;// level 2
assign po606 = ~w17720;// level 2
assign po607 = ~w17723;// level 2
assign po608 = ~w17726;// level 2
assign po609 = ~w17729;// level 2
assign po610 = ~w17732;// level 2
assign po611 = ~w17735;// level 2
assign po612 = ~w17738;// level 2
assign po613 = ~w17741;// level 2
assign po614 = ~w17744;// level 2
assign po615 = ~w17747;// level 2
assign po616 = ~w17750;// level 2
assign po617 = ~w17753;// level 2
assign po618 = ~w17756;// level 2
assign po619 = ~w17759;// level 2
assign po620 = w17760;// level 4
assign po621 = ~w17763;// level 2
assign po622 = ~w17766;// level 2
assign po623 = ~w17769;// level 2
assign po624 = ~w17772;// level 2
assign po625 = w17489;// level 3
assign po626 = ~w17775;// level 2
assign po627 = ~w17778;// level 2
assign po628 = ~w17781;// level 2
assign po629 = ~w17784;// level 2
assign po630 = ~w17787;// level 2
assign po631 = ~w17790;// level 2
assign po632 = ~w17793;// level 2
assign po633 = ~w17796;// level 2
assign po634 = ~w17799;// level 2
assign po635 = ~w17802;// level 2
assign po636 = ~w17805;// level 2
assign po637 = ~w17808;// level 2
assign po638 = ~w17811;// level 2
assign po639 = ~w17814;// level 2
assign po640 = ~w17817;// level 2
assign po641 = ~w17820;// level 2
assign po642 = ~w17823;// level 2
assign po643 = ~w17826;// level 2
assign po644 = ~w17829;// level 2
assign po645 = ~w17832;// level 2
assign po646 = ~w17835;// level 2
assign po647 = ~w17838;// level 2
assign po648 = ~w17841;// level 2
assign po649 = ~w17844;// level 2
assign po650 = ~w17847;// level 2
assign po651 = ~w17850;// level 2
assign po652 = ~w17853;// level 2
assign po653 = ~w17856;// level 2
assign po654 = ~w17859;// level 2
assign po655 = ~w17862;// level 2
assign po656 = ~w17865;// level 2
assign po657 = ~w17868;// level 2
assign po658 = w17475;// level 1
assign po659 = ~w17871;// level 2
assign po660 = ~w17874;// level 2
assign po661 = ~w17877;// level 2
assign po662 = ~w17880;// level 2
assign po663 = ~w17883;// level 2
assign po664 = ~w17886;// level 2
assign po665 = ~w17889;// level 2
assign po666 = ~w17892;// level 2
assign po667 = pi532;// level 0
endmodule
