//Written by the Majority Logic Package Fri May  1 00:24:02 2015
module top (
            pi000, pi001, pi002, pi003, pi004, pi005, pi006, pi007, pi008, pi009, pi010, pi011, pi012, pi013, pi014, pi015, pi016, pi017, pi018, pi019, pi020, pi021, pi022, pi023, pi024, pi025, pi026, pi027, pi028, pi029, pi030, pi031, pi032, pi033, pi034, pi035, pi036, pi037, pi038, pi039, pi040, pi041, pi042, pi043, pi044, pi045, pi046, pi047, pi048, pi049, pi050, pi051, pi052, pi053, pi054, pi055, pi056, pi057, pi058, pi059, pi060, pi061, pi062, pi063, pi064, pi065, pi066, pi067, pi068, pi069, pi070, pi071, pi072, pi073, pi074, pi075, pi076, pi077, pi078, pi079, pi080, pi081, pi082, pi083, pi084, pi085, pi086, pi087, pi088, pi089, pi090, pi091, pi092, pi093, pi094, pi095, pi096, pi097, pi098, pi099, pi100, pi101, pi102, pi103, pi104, pi105, pi106, pi107, pi108, pi109, pi110, pi111, pi112, pi113, pi114, pi115, pi116, pi117, pi118, pi119, pi120, pi121, pi122, pi123, pi124, pi125, pi126, pi127, pi128, pi129, pi130, pi131, pi132, pi133, pi134, pi135, pi136, pi137, pi138, pi139, pi140, pi141, pi142, pi143, pi144, pi145, pi146, pi147, pi148, pi149, pi150, pi151, pi152, pi153, pi154, pi155, pi156, pi157, pi158, pi159, pi160, pi161, pi162, pi163, pi164, pi165, pi166, pi167, pi168, pi169, pi170, pi171, pi172, pi173, pi174, pi175, pi176, pi177, pi178, pi179, pi180, pi181, pi182, pi183, pi184, pi185, pi186, pi187, pi188, pi189, pi190, pi191, pi192, pi193, pi194, pi195, pi196, pi197, pi198, pi199, pi200, pi201, pi202, pi203, pi204, pi205, pi206, pi207, pi208, pi209, pi210, pi211, pi212, pi213, pi214, pi215, pi216, pi217, pi218, pi219, pi220, pi221, pi222, pi223, pi224, pi225, pi226, pi227, pi228, pi229, pi230, pi231, pi232, pi233, pi234, pi235, pi236, pi237, pi238, pi239, pi240, pi241, pi242, pi243, pi244, pi245, pi246, pi247, pi248, pi249, pi250, pi251, pi252, pi253, pi254, pi255, pi256, pi257, pi258, pi259, pi260, pi261, pi262, pi263, pi264, pi265, pi266, pi267, pi268, pi269, pi270, pi271, pi272, pi273, pi274, pi275, pi276, pi277, pi278, pi279, pi280, pi281, pi282, pi283, pi284, pi285, pi286, pi287, pi288, pi289, pi290, pi291, pi292, pi293, pi294, pi295, pi296, pi297, pi298, pi299, pi300, pi301, pi302, pi303, pi304, pi305, pi306, pi307, pi308, pi309, pi310, pi311, pi312, pi313, pi314, pi315, pi316, pi317, pi318, pi319, pi320, pi321, pi322, pi323, pi324, pi325, pi326, pi327, pi328, pi329, pi330, pi331, pi332, pi333, pi334, pi335, pi336, pi337, pi338, pi339, pi340, pi341, pi342, pi343, pi344, pi345, pi346, pi347, pi348, pi349, pi350, pi351, pi352, pi353, 
            po000, po001, po002, po003, po004, po005, po006, po007, po008, po009, po010, po011, po012, po013, po014, po015, po016, po017, po018, po019, po020, po021, po022, po023, po024, po025, po026, po027, po028, po029, po030, po031, po032, po033, po034, po035, po036, po037, po038, po039, po040, po041, po042, po043, po044, po045, po046, po047, po048, po049, po050, po051, po052, po053, po054, po055, po056, po057, po058, po059, po060, po061, po062, po063, po064, po065, po066, po067, po068, po069, po070, po071, po072, po073, po074, po075, po076, po077, po078, po079, po080, po081, po082, po083, po084, po085, po086, po087, po088, po089, po090, po091, po092, po093, po094, po095, po096, po097, po098, po099, po100, po101, po102, po103, po104, po105, po106, po107, po108, po109, po110, po111, po112, po113, po114, po115, po116, po117, po118, po119, po120, po121, po122, po123, po124, po125, po126, po127, po128, po129, po130, po131, po132, po133, po134, po135, po136, po137, po138, po139, po140, po141, po142, po143, po144, po145, po146, po147, po148, po149, po150, po151, po152, po153, po154, po155, po156, po157, po158, po159, po160, po161, po162, po163, po164, po165, po166, po167, po168, po169, po170, po171, po172, po173, po174, po175, po176, po177, po178, po179, po180, po181, po182, po183, po184, po185, po186, po187, po188, po189, po190, po191, po192, po193, po194, po195, po196, po197, po198, po199, po200, po201, po202, po203, po204, po205, po206, po207, po208, po209, po210, po211, po212, po213, po214, po215, po216, po217, po218, po219, po220, po221, po222, po223, po224, po225, po226, po227, po228, po229, po230, po231, po232, po233, po234, po235, po236, po237, po238, po239, po240, po241, po242, po243, po244, po245, po246, po247, po248, po249, po250, po251, po252, po253, po254, po255, po256, po257, po258, po259, po260, po261, po262, po263, po264, po265, po266, po267, po268, po269, po270, po271, po272, po273, po274, po275, po276, po277, po278, po279, po280, po281, po282, po283, po284, po285, po286, po287, po288);
input pi000, pi001, pi002, pi003, pi004, pi005, pi006, pi007, pi008, pi009, pi010, pi011, pi012, pi013, pi014, pi015, pi016, pi017, pi018, pi019, pi020, pi021, pi022, pi023, pi024, pi025, pi026, pi027, pi028, pi029, pi030, pi031, pi032, pi033, pi034, pi035, pi036, pi037, pi038, pi039, pi040, pi041, pi042, pi043, pi044, pi045, pi046, pi047, pi048, pi049, pi050, pi051, pi052, pi053, pi054, pi055, pi056, pi057, pi058, pi059, pi060, pi061, pi062, pi063, pi064, pi065, pi066, pi067, pi068, pi069, pi070, pi071, pi072, pi073, pi074, pi075, pi076, pi077, pi078, pi079, pi080, pi081, pi082, pi083, pi084, pi085, pi086, pi087, pi088, pi089, pi090, pi091, pi092, pi093, pi094, pi095, pi096, pi097, pi098, pi099, pi100, pi101, pi102, pi103, pi104, pi105, pi106, pi107, pi108, pi109, pi110, pi111, pi112, pi113, pi114, pi115, pi116, pi117, pi118, pi119, pi120, pi121, pi122, pi123, pi124, pi125, pi126, pi127, pi128, pi129, pi130, pi131, pi132, pi133, pi134, pi135, pi136, pi137, pi138, pi139, pi140, pi141, pi142, pi143, pi144, pi145, pi146, pi147, pi148, pi149, pi150, pi151, pi152, pi153, pi154, pi155, pi156, pi157, pi158, pi159, pi160, pi161, pi162, pi163, pi164, pi165, pi166, pi167, pi168, pi169, pi170, pi171, pi172, pi173, pi174, pi175, pi176, pi177, pi178, pi179, pi180, pi181, pi182, pi183, pi184, pi185, pi186, pi187, pi188, pi189, pi190, pi191, pi192, pi193, pi194, pi195, pi196, pi197, pi198, pi199, pi200, pi201, pi202, pi203, pi204, pi205, pi206, pi207, pi208, pi209, pi210, pi211, pi212, pi213, pi214, pi215, pi216, pi217, pi218, pi219, pi220, pi221, pi222, pi223, pi224, pi225, pi226, pi227, pi228, pi229, pi230, pi231, pi232, pi233, pi234, pi235, pi236, pi237, pi238, pi239, pi240, pi241, pi242, pi243, pi244, pi245, pi246, pi247, pi248, pi249, pi250, pi251, pi252, pi253, pi254, pi255, pi256, pi257, pi258, pi259, pi260, pi261, pi262, pi263, pi264, pi265, pi266, pi267, pi268, pi269, pi270, pi271, pi272, pi273, pi274, pi275, pi276, pi277, pi278, pi279, pi280, pi281, pi282, pi283, pi284, pi285, pi286, pi287, pi288, pi289, pi290, pi291, pi292, pi293, pi294, pi295, pi296, pi297, pi298, pi299, pi300, pi301, pi302, pi303, pi304, pi305, pi306, pi307, pi308, pi309, pi310, pi311, pi312, pi313, pi314, pi315, pi316, pi317, pi318, pi319, pi320, pi321, pi322, pi323, pi324, pi325, pi326, pi327, pi328, pi329, pi330, pi331, pi332, pi333, pi334, pi335, pi336, pi337, pi338, pi339, pi340, pi341, pi342, pi343, pi344, pi345, pi346, pi347, pi348, pi349, pi350, pi351, pi352, pi353;
output po000, po001, po002, po003, po004, po005, po006, po007, po008, po009, po010, po011, po012, po013, po014, po015, po016, po017, po018, po019, po020, po021, po022, po023, po024, po025, po026, po027, po028, po029, po030, po031, po032, po033, po034, po035, po036, po037, po038, po039, po040, po041, po042, po043, po044, po045, po046, po047, po048, po049, po050, po051, po052, po053, po054, po055, po056, po057, po058, po059, po060, po061, po062, po063, po064, po065, po066, po067, po068, po069, po070, po071, po072, po073, po074, po075, po076, po077, po078, po079, po080, po081, po082, po083, po084, po085, po086, po087, po088, po089, po090, po091, po092, po093, po094, po095, po096, po097, po098, po099, po100, po101, po102, po103, po104, po105, po106, po107, po108, po109, po110, po111, po112, po113, po114, po115, po116, po117, po118, po119, po120, po121, po122, po123, po124, po125, po126, po127, po128, po129, po130, po131, po132, po133, po134, po135, po136, po137, po138, po139, po140, po141, po142, po143, po144, po145, po146, po147, po148, po149, po150, po151, po152, po153, po154, po155, po156, po157, po158, po159, po160, po161, po162, po163, po164, po165, po166, po167, po168, po169, po170, po171, po172, po173, po174, po175, po176, po177, po178, po179, po180, po181, po182, po183, po184, po185, po186, po187, po188, po189, po190, po191, po192, po193, po194, po195, po196, po197, po198, po199, po200, po201, po202, po203, po204, po205, po206, po207, po208, po209, po210, po211, po212, po213, po214, po215, po216, po217, po218, po219, po220, po221, po222, po223, po224, po225, po226, po227, po228, po229, po230, po231, po232, po233, po234, po235, po236, po237, po238, po239, po240, po241, po242, po243, po244, po245, po246, po247, po248, po249, po250, po251, po252, po253, po254, po255, po256, po257, po258, po259, po260, po261, po262, po263, po264, po265, po266, po267, po268, po269, po270, po271, po272, po273, po274, po275, po276, po277, po278, po279, po280, po281, po282, po283, po284, po285, po286, po287, po288;
wire one, w0, w1, w2, w3, w4, w5, w6, w7, w8, w9, w10, w11, w12, w13, w14, w15, w16, w17, w18, w19, w20, w21, w22, w23, w24, w25, w26, w27, w28, w29, w30, w31, w32, w33, w34, w35, w36, w37, w38, w39, w40, w41, w42, w43, w44, w45, w46, w47, w48, w49, w50, w51, w52, w53, w54, w55, w56, w57, w58, w59, w60, w61, w62, w63, w64, w65, w66, w67, w68, w69, w70, w71, w72, w73, w74, w75, w76, w77, w78, w79, w80, w81, w82, w83, w84, w85, w86, w87, w88, w89, w90, w91, w92, w93, w94, w95, w96, w97, w98, w99, w100, w101, w102, w103, w104, w105, w106, w107, w108, w109, w110, w111, w112, w113, w114, w115, w116, w117, w118, w119, w120, w121, w122, w123, w124, w125, w126, w127, w128, w129, w130, w131, w132, w133, w134, w135, w136, w137, w138, w139, w140, w141, w142, w143, w144, w145, w146, w147, w148, w149, w150, w151, w152, w153, w154, w155, w156, w157, w158, w159, w160, w161, w162, w163, w164, w165, w166, w167, w168, w169, w170, w171, w172, w173, w174, w175, w176, w177, w178, w179, w180, w181, w182, w183, w184, w185, w186, w187, w188, w189, w190, w191, w192, w193, w194, w195, w196, w197, w198, w199, w200, w201, w202, w203, w204, w205, w206, w207, w208, w209, w210, w211, w212, w213, w214, w215, w216, w217, w218, w219, w220, w221, w222, w223, w224, w225, w226, w227, w228, w229, w230, w231, w232, w233, w234, w235, w236, w237, w238, w239, w240, w241, w242, w243, w244, w245, w246, w247, w248, w249, w250, w251, w252, w253, w254, w255, w256, w257, w258, w259, w260, w261, w262, w263, w264, w265, w266, w267, w268, w269, w270, w271, w272, w273, w274, w275, w276, w277, w278, w279, w280, w281, w282, w283, w284, w285, w286, w287, w288, w289, w290, w291, w292, w293, w294, w295, w296, w297, w298, w299, w300, w301, w302, w303, w304, w305, w306, w307, w308, w309, w310, w311, w312, w313, w314, w315, w316, w317, w318, w319, w320, w321, w322, w323, w324, w325, w326, w327, w328, w329, w330, w331, w332, w333, w334, w335, w336, w337, w338, w339, w340, w341, w342, w343, w344, w345, w346, w347, w348, w349, w350, w351, w352, w353, w354, w355, w356, w357, w358, w359, w360, w361, w362, w363, w364, w365, w366, w367, w368, w369, w370, w371, w372, w373, w374, w375, w376, w377, w378, w379, w380, w381, w382, w383, w384, w385, w386, w387, w388, w389, w390, w391, w392, w393, w394, w395, w396, w397, w398, w399, w400, w401, w402, w403, w404, w405, w406, w407, w408, w409, w410, w411, w412, w413, w414, w415, w416, w417, w418, w419, w420, w421, w422, w423, w424, w425, w426, w427, w428, w429, w430, w431, w432, w433, w434, w435, w436, w437, w438, w439, w440, w441, w442, w443, w444, w445, w446, w447, w448, w449, w450, w451, w452, w453, w454, w455, w456, w457, w458, w459, w460, w461, w462, w463, w464, w465, w466, w467, w468, w469, w470, w471, w472, w473, w474, w475, w476, w477, w478, w479, w480, w481, w482, w483, w484, w485, w486, w487, w488, w489, w490, w491, w492, w493, w494, w495, w496, w497, w498, w499, w500, w501, w502, w503, w504, w505, w506, w507, w508, w509, w510, w511, w512, w513, w514, w515, w516, w517, w518, w519, w520, w521, w522, w523, w524, w525, w526, w527, w528, w529, w530, w531, w532, w533, w534, w535, w536, w537, w538, w539, w540, w541, w542, w543, w544, w545, w546, w547, w548, w549, w550, w551, w552, w553, w554, w555, w556, w557, w558, w559, w560, w561, w562, w563, w564, w565, w566, w567, w568, w569, w570, w571, w572, w573, w574, w575, w576, w577, w578, w579, w580, w581, w582, w583, w584, w585, w586, w587, w588, w589, w590, w591, w592, w593, w594, w595, w596, w597, w598, w599, w600, w601, w602, w603, w604, w605, w606, w607, w608, w609, w610, w611, w612, w613, w614, w615, w616, w617, w618, w619, w620, w621, w622, w623, w624, w625, w626, w627, w628, w629, w630, w631, w632, w633, w634, w635, w636, w637, w638, w639, w640, w641, w642, w643, w644, w645, w646, w647, w648, w649, w650, w651, w652, w653, w654, w655, w656, w657, w658, w659, w660, w661, w662, w663, w664, w665, w666, w667, w668, w669, w670, w671, w672, w673, w674, w675, w676, w677, w678, w679, w680, w681, w682, w683, w684, w685, w686, w687, w688, w689, w690, w691, w692, w693, w694, w695, w696, w697, w698, w699, w700, w701, w702, w703, w704, w705, w706, w707, w708, w709, w710, w711, w712, w713, w714, w715, w716, w717, w718, w719, w720, w721, w722, w723, w724, w725, w726, w727, w728, w729, w730, w731, w732, w733, w734, w735, w736, w737, w738, w739, w740, w741, w742, w743, w744, w745, w746, w747, w748, w749, w750, w751, w752, w753, w754, w755, w756, w757, w758, w759, w760, w761, w762, w763, w764, w765, w766, w767, w768, w769, w770, w771, w772, w773, w774, w775, w776, w777, w778, w779, w780, w781, w782, w783, w784, w785, w786, w787, w788, w789, w790, w791, w792, w793, w794, w795, w796, w797, w798, w799, w800, w801, w802, w803, w804, w805, w806, w807, w808, w809, w810, w811, w812, w813, w814, w815, w816, w817, w818, w819, w820, w821, w822, w823, w824, w825, w826, w827, w828, w829, w830, w831, w832, w833, w834, w835, w836, w837, w838, w839, w840, w841, w842, w843, w844, w845, w846, w847, w848, w849, w850, w851, w852, w853, w854, w855, w856, w857, w858, w859, w860, w861, w862, w863, w864, w865, w866, w867, w868, w869, w870, w871, w872, w873, w874, w875, w876, w877, w878, w879, w880, w881, w882, w883, w884, w885, w886, w887, w888, w889, w890, w891, w892, w893, w894, w895, w896, w897, w898, w899, w900, w901, w902, w903, w904, w905, w906, w907, w908, w909, w910, w911, w912, w913, w914, w915, w916, w917, w918, w919, w920, w921, w922, w923, w924, w925, w926, w927, w928, w929, w930, w931, w932, w933, w934, w935, w936, w937, w938, w939, w940, w941, w942, w943, w944, w945, w946, w947, w948, w949, w950, w951, w952, w953, w954, w955, w956, w957, w958, w959, w960, w961, w962, w963, w964, w965, w966, w967, w968, w969, w970, w971, w972, w973, w974, w975, w976, w977, w978, w979, w980, w981, w982, w983, w984, w985, w986, w987, w988, w989, w990, w991, w992, w993, w994, w995, w996, w997, w998, w999, w1000, w1001, w1002, w1003, w1004, w1005, w1006, w1007, w1008, w1009, w1010, w1011, w1012, w1013, w1014, w1015, w1016, w1017, w1018, w1019, w1020, w1021, w1022, w1023, w1024, w1025, w1026, w1027, w1028, w1029, w1030, w1031, w1032, w1033, w1034, w1035, w1036, w1037, w1038, w1039, w1040, w1041, w1042, w1043, w1044, w1045, w1046, w1047, w1048, w1049, w1050, w1051, w1052, w1053, w1054, w1055, w1056, w1057, w1058, w1059, w1060, w1061, w1062, w1063, w1064, w1065, w1066, w1067, w1068, w1069, w1070, w1071, w1072, w1073, w1074, w1075, w1076, w1077, w1078, w1079, w1080, w1081, w1082, w1083, w1084, w1085, w1086, w1087, w1088, w1089, w1090, w1091, w1092, w1093, w1094, w1095, w1096, w1097, w1098, w1099, w1100, w1101, w1102, w1103, w1104, w1105, w1106, w1107, w1108, w1109, w1110, w1111, w1112, w1113, w1114, w1115, w1116, w1117, w1118, w1119, w1120, w1121, w1122, w1123, w1124, w1125, w1126, w1127, w1128, w1129, w1130, w1131, w1132, w1133, w1134, w1135, w1136, w1137, w1138, w1139, w1140, w1141, w1142, w1143, w1144, w1145, w1146, w1147, w1148, w1149, w1150, w1151, w1152, w1153, w1154, w1155, w1156, w1157, w1158, w1159, w1160, w1161, w1162, w1163, w1164, w1165, w1166, w1167, w1168, w1169, w1170, w1171, w1172, w1173, w1174, w1175, w1176, w1177, w1178, w1179, w1180, w1181, w1182, w1183, w1184, w1185, w1186, w1187, w1188, w1189, w1190, w1191, w1192, w1193, w1194, w1195, w1196, w1197, w1198, w1199, w1200, w1201, w1202, w1203, w1204, w1205, w1206, w1207, w1208, w1209, w1210, w1211, w1212, w1213, w1214, w1215, w1216, w1217, w1218, w1219, w1220, w1221, w1222, w1223, w1224, w1225, w1226, w1227, w1228, w1229, w1230, w1231, w1232, w1233, w1234, w1235, w1236, w1237, w1238, w1239, w1240, w1241, w1242, w1243, w1244, w1245, w1246, w1247, w1248, w1249, w1250, w1251, w1252, w1253, w1254, w1255, w1256, w1257, w1258, w1259, w1260, w1261, w1262, w1263, w1264, w1265, w1266, w1267, w1268, w1269, w1270, w1271, w1272, w1273, w1274, w1275, w1276, w1277, w1278, w1279, w1280, w1281, w1282, w1283, w1284, w1285, w1286, w1287, w1288, w1289, w1290, w1291, w1292, w1293, w1294, w1295, w1296, w1297, w1298, w1299, w1300, w1301, w1302, w1303, w1304, w1305, w1306, w1307, w1308, w1309, w1310, w1311, w1312, w1313, w1314, w1315, w1316, w1317, w1318, w1319, w1320, w1321, w1322, w1323, w1324, w1325, w1326, w1327, w1328, w1329, w1330, w1331, w1332, w1333, w1334, w1335, w1336, w1337, w1338, w1339, w1340, w1341, w1342, w1343, w1344, w1345, w1346, w1347, w1348, w1349, w1350, w1351, w1352, w1353, w1354, w1355, w1356, w1357, w1358, w1359, w1360, w1361, w1362, w1363, w1364, w1365, w1366, w1367, w1368, w1369, w1370, w1371, w1372, w1373, w1374, w1375, w1376, w1377, w1378, w1379, w1380, w1381, w1382, w1383, w1384, w1385, w1386, w1387, w1388, w1389, w1390, w1391, w1392, w1393, w1394, w1395, w1396, w1397, w1398, w1399, w1400, w1401, w1402, w1403, w1404, w1405, w1406, w1407, w1408, w1409, w1410, w1411, w1412, w1413, w1414, w1415, w1416, w1417, w1418, w1419, w1420, w1421, w1422, w1423, w1424, w1425, w1426, w1427, w1428, w1429, w1430, w1431, w1432, w1433, w1434, w1435, w1436, w1437, w1438, w1439, w1440, w1441, w1442, w1443, w1444, w1445, w1446, w1447, w1448, w1449, w1450, w1451, w1452, w1453, w1454, w1455, w1456, w1457, w1458, w1459, w1460, w1461, w1462, w1463, w1464, w1465, w1466, w1467, w1468, w1469, w1470, w1471, w1472, w1473, w1474, w1475, w1476, w1477, w1478, w1479, w1480, w1481, w1482, w1483, w1484, w1485, w1486, w1487, w1488, w1489, w1490, w1491, w1492, w1493, w1494, w1495, w1496, w1497, w1498, w1499, w1500, w1501, w1502, w1503, w1504, w1505, w1506, w1507, w1508, w1509, w1510, w1511, w1512, w1513, w1514, w1515, w1516, w1517, w1518, w1519, w1520, w1521, w1522, w1523, w1524, w1525, w1526, w1527, w1528, w1529, w1530, w1531, w1532, w1533, w1534, w1535, w1536, w1537, w1538, w1539, w1540, w1541, w1542, w1543, w1544, w1545, w1546, w1547, w1548, w1549, w1550, w1551, w1552, w1553, w1554, w1555, w1556, w1557, w1558, w1559, w1560, w1561, w1562, w1563, w1564, w1565, w1566, w1567, w1568, w1569, w1570, w1571, w1572, w1573, w1574, w1575, w1576, w1577, w1578, w1579, w1580, w1581, w1582, w1583, w1584, w1585, w1586, w1587, w1588, w1589, w1590, w1591, w1592, w1593, w1594, w1595, w1596, w1597, w1598, w1599, w1600, w1601, w1602, w1603, w1604, w1605, w1606, w1607, w1608, w1609, w1610, w1611, w1612, w1613, w1614, w1615, w1616, w1617, w1618, w1619, w1620, w1621, w1622, w1623, w1624, w1625, w1626, w1627, w1628, w1629, w1630, w1631, w1632, w1633, w1634, w1635, w1636, w1637, w1638, w1639, w1640, w1641, w1642, w1643, w1644, w1645, w1646, w1647, w1648, w1649, w1650, w1651, w1652, w1653, w1654, w1655, w1656, w1657, w1658, w1659, w1660, w1661, w1662, w1663, w1664, w1665, w1666, w1667, w1668, w1669, w1670, w1671, w1672, w1673, w1674, w1675, w1676, w1677, w1678, w1679, w1680, w1681, w1682, w1683, w1684, w1685, w1686, w1687, w1688, w1689, w1690, w1691, w1692, w1693, w1694, w1695, w1696, w1697, w1698, w1699, w1700, w1701, w1702, w1703, w1704, w1705, w1706, w1707, w1708, w1709, w1710, w1711, w1712, w1713, w1714, w1715, w1716, w1717, w1718, w1719, w1720, w1721, w1722, w1723, w1724, w1725, w1726, w1727, w1728, w1729, w1730, w1731, w1732, w1733, w1734, w1735, w1736, w1737, w1738, w1739, w1740, w1741, w1742, w1743, w1744, w1745, w1746, w1747, w1748, w1749, w1750, w1751, w1752, w1753, w1754, w1755, w1756, w1757, w1758, w1759, w1760, w1761, w1762, w1763, w1764, w1765, w1766, w1767, w1768, w1769, w1770, w1771, w1772, w1773, w1774, w1775, w1776, w1777, w1778, w1779, w1780, w1781, w1782, w1783, w1784, w1785, w1786, w1787, w1788, w1789, w1790, w1791, w1792, w1793, w1794, w1795, w1796, w1797, w1798, w1799, w1800, w1801, w1802, w1803, w1804, w1805, w1806, w1807, w1808, w1809, w1810, w1811, w1812, w1813, w1814, w1815, w1816, w1817, w1818, w1819, w1820, w1821, w1822, w1823, w1824, w1825, w1826, w1827, w1828, w1829, w1830, w1831, w1832, w1833, w1834, w1835, w1836, w1837, w1838, w1839, w1840, w1841, w1842, w1843, w1844, w1845, w1846, w1847, w1848, w1849, w1850, w1851, w1852, w1853, w1854, w1855, w1856, w1857, w1858, w1859, w1860, w1861, w1862, w1863, w1864, w1865, w1866, w1867, w1868, w1869, w1870, w1871, w1872, w1873, w1874, w1875, w1876, w1877, w1878, w1879, w1880, w1881, w1882, w1883, w1884, w1885, w1886, w1887, w1888, w1889, w1890, w1891, w1892, w1893, w1894, w1895, w1896, w1897, w1898, w1899, w1900, w1901, w1902, w1903, w1904, w1905, w1906, w1907, w1908, w1909, w1910, w1911, w1912, w1913, w1914, w1915, w1916, w1917, w1918, w1919, w1920, w1921, w1922, w1923, w1924, w1925, w1926, w1927, w1928, w1929, w1930, w1931, w1932, w1933, w1934, w1935, w1936, w1937, w1938, w1939, w1940, w1941, w1942, w1943, w1944, w1945, w1946, w1947, w1948, w1949, w1950, w1951, w1952, w1953, w1954, w1955, w1956, w1957, w1958, w1959, w1960, w1961, w1962, w1963, w1964, w1965, w1966, w1967, w1968, w1969, w1970, w1971, w1972, w1973, w1974, w1975, w1976, w1977, w1978, w1979, w1980, w1981, w1982, w1983, w1984, w1985, w1986, w1987, w1988, w1989, w1990, w1991, w1992, w1993, w1994, w1995, w1996, w1997, w1998, w1999, w2000, w2001, w2002, w2003, w2004, w2005, w2006, w2007, w2008, w2009, w2010, w2011, w2012, w2013, w2014, w2015, w2016, w2017, w2018, w2019, w2020, w2021, w2022, w2023, w2024, w2025, w2026, w2027, w2028, w2029, w2030, w2031, w2032, w2033, w2034, w2035, w2036, w2037, w2038, w2039, w2040, w2041, w2042, w2043, w2044, w2045, w2046, w2047, w2048, w2049, w2050, w2051, w2052, w2053, w2054, w2055, w2056, w2057, w2058, w2059, w2060, w2061, w2062, w2063, w2064, w2065, w2066, w2067, w2068, w2069, w2070, w2071, w2072, w2073, w2074, w2075, w2076, w2077, w2078, w2079, w2080, w2081, w2082, w2083, w2084, w2085, w2086, w2087, w2088, w2089, w2090, w2091, w2092, w2093, w2094, w2095, w2096, w2097, w2098, w2099, w2100, w2101, w2102, w2103, w2104, w2105, w2106, w2107, w2108, w2109, w2110, w2111, w2112, w2113, w2114, w2115, w2116, w2117, w2118, w2119, w2120, w2121, w2122, w2123, w2124, w2125, w2126, w2127, w2128, w2129, w2130, w2131, w2132, w2133, w2134, w2135, w2136, w2137, w2138, w2139, w2140, w2141, w2142, w2143, w2144, w2145, w2146, w2147, w2148, w2149, w2150, w2151, w2152, w2153, w2154, w2155, w2156, w2157, w2158, w2159, w2160, w2161, w2162, w2163, w2164, w2165, w2166, w2167, w2168, w2169, w2170, w2171, w2172, w2173, w2174, w2175, w2176, w2177, w2178, w2179, w2180, w2181, w2182, w2183, w2184, w2185, w2186, w2187, w2188, w2189, w2190, w2191, w2192, w2193, w2194, w2195, w2196, w2197, w2198, w2199, w2200, w2201, w2202, w2203, w2204, w2205, w2206, w2207, w2208, w2209, w2210, w2211, w2212, w2213, w2214, w2215, w2216, w2217, w2218, w2219, w2220, w2221, w2222, w2223, w2224, w2225, w2226, w2227, w2228, w2229, w2230, w2231, w2232, w2233, w2234, w2235, w2236, w2237, w2238, w2239, w2240, w2241, w2242, w2243, w2244, w2245, w2246, w2247, w2248, w2249, w2250, w2251, w2252, w2253, w2254, w2255, w2256, w2257, w2258, w2259, w2260, w2261, w2262, w2263, w2264, w2265, w2266, w2267, w2268, w2269, w2270, w2271, w2272, w2273, w2274, w2275, w2276, w2277, w2278, w2279, w2280, w2281, w2282, w2283, w2284, w2285, w2286, w2287, w2288, w2289, w2290, w2291, w2292, w2293, w2294, w2295, w2296, w2297, w2298, w2299, w2300, w2301, w2302, w2303, w2304, w2305, w2306, w2307, w2308, w2309, w2310, w2311, w2312, w2313, w2314, w2315, w2316, w2317, w2318, w2319, w2320, w2321, w2322, w2323, w2324, w2325, w2326, w2327, w2328, w2329, w2330, w2331, w2332, w2333, w2334, w2335, w2336, w2337, w2338, w2339, w2340, w2341, w2342, w2343, w2344, w2345, w2346, w2347, w2348, w2349, w2350, w2351, w2352, w2353, w2354, w2355, w2356, w2357, w2358, w2359, w2360, w2361, w2362, w2363, w2364, w2365, w2366, w2367, w2368, w2369, w2370, w2371, w2372, w2373, w2374, w2375, w2376, w2377, w2378, w2379, w2380, w2381, w2382, w2383, w2384, w2385, w2386, w2387, w2388, w2389, w2390, w2391, w2392, w2393, w2394, w2395, w2396, w2397, w2398, w2399, w2400, w2401, w2402, w2403, w2404, w2405, w2406, w2407, w2408, w2409, w2410, w2411, w2412, w2413, w2414, w2415, w2416, w2417, w2418, w2419, w2420, w2421, w2422, w2423, w2424, w2425, w2426, w2427, w2428, w2429, w2430, w2431, w2432, w2433, w2434, w2435, w2436, w2437, w2438, w2439, w2440, w2441, w2442, w2443, w2444, w2445, w2446, w2447, w2448, w2449, w2450, w2451, w2452, w2453, w2454, w2455, w2456, w2457, w2458, w2459, w2460, w2461, w2462, w2463, w2464, w2465, w2466, w2467, w2468, w2469, w2470, w2471, w2472, w2473, w2474, w2475, w2476, w2477, w2478, w2479, w2480, w2481, w2482, w2483, w2484, w2485, w2486, w2487, w2488, w2489, w2490, w2491, w2492, w2493, w2494, w2495, w2496, w2497, w2498, w2499, w2500, w2501, w2502, w2503, w2504, w2505, w2506, w2507, w2508, w2509, w2510, w2511, w2512, w2513, w2514, w2515, w2516, w2517, w2518, w2519, w2520, w2521, w2522, w2523, w2524, w2525, w2526, w2527, w2528, w2529, w2530, w2531, w2532, w2533, w2534, w2535, w2536, w2537, w2538, w2539, w2540, w2541, w2542, w2543, w2544, w2545, w2546, w2547, w2548, w2549, w2550, w2551, w2552, w2553, w2554, w2555, w2556, w2557, w2558, w2559, w2560, w2561, w2562, w2563, w2564, w2565, w2566, w2567, w2568, w2569, w2570, w2571, w2572, w2573, w2574, w2575, w2576, w2577, w2578, w2579, w2580, w2581, w2582, w2583, w2584, w2585, w2586, w2587, w2588, w2589, w2590, w2591, w2592, w2593, w2594, w2595, w2596, w2597, w2598, w2599, w2600, w2601, w2602, w2603, w2604, w2605, w2606, w2607, w2608, w2609, w2610, w2611, w2612, w2613, w2614, w2615, w2616, w2617, w2618, w2619, w2620, w2621, w2622, w2623, w2624, w2625, w2626, w2627, w2628, w2629, w2630, w2631, w2632, w2633, w2634, w2635, w2636, w2637, w2638, w2639, w2640, w2641, w2642, w2643, w2644, w2645, w2646, w2647, w2648, w2649, w2650, w2651, w2652, w2653, w2654, w2655, w2656, w2657, w2658, w2659, w2660, w2661, w2662, w2663, w2664, w2665, w2666, w2667, w2668, w2669, w2670, w2671, w2672, w2673, w2674, w2675, w2676, w2677, w2678, w2679, w2680, w2681, w2682, w2683, w2684, w2685, w2686, w2687, w2688, w2689, w2690, w2691, w2692, w2693, w2694, w2695, w2696, w2697, w2698, w2699, w2700, w2701, w2702, w2703, w2704, w2705, w2706, w2707, w2708, w2709, w2710, w2711, w2712, w2713, w2714, w2715, w2716, w2717, w2718, w2719, w2720, w2721, w2722, w2723, w2724, w2725, w2726, w2727, w2728, w2729, w2730, w2731, w2732, w2733, w2734, w2735, w2736, w2737, w2738, w2739, w2740, w2741, w2742, w2743, w2744, w2745, w2746, w2747, w2748, w2749, w2750, w2751, w2752, w2753, w2754, w2755, w2756, w2757, w2758, w2759, w2760, w2761, w2762, w2763, w2764, w2765, w2766, w2767, w2768, w2769, w2770, w2771, w2772, w2773, w2774, w2775, w2776, w2777, w2778, w2779, w2780, w2781, w2782, w2783, w2784, w2785, w2786, w2787, w2788, w2789, w2790, w2791, w2792, w2793, w2794, w2795, w2796, w2797, w2798, w2799, w2800, w2801, w2802, w2803, w2804, w2805, w2806, w2807, w2808, w2809, w2810, w2811, w2812, w2813, w2814, w2815, w2816, w2817, w2818, w2819, w2820, w2821, w2822, w2823, w2824, w2825, w2826, w2827, w2828, w2829, w2830, w2831, w2832, w2833, w2834, w2835, w2836, w2837, w2838, w2839, w2840, w2841, w2842, w2843, w2844, w2845, w2846, w2847, w2848, w2849, w2850, w2851, w2852, w2853, w2854, w2855, w2856, w2857, w2858, w2859, w2860, w2861, w2862, w2863, w2864, w2865, w2866, w2867, w2868, w2869, w2870, w2871, w2872, w2873, w2874, w2875, w2876, w2877, w2878, w2879, w2880, w2881, w2882, w2883, w2884, w2885, w2886, w2887, w2888, w2889, w2890, w2891, w2892, w2893, w2894, w2895, w2896, w2897, w2898, w2899, w2900, w2901, w2902, w2903, w2904, w2905, w2906, w2907, w2908, w2909, w2910, w2911, w2912, w2913, w2914, w2915, w2916, w2917, w2918, w2919, w2920, w2921, w2922, w2923, w2924, w2925, w2926, w2927, w2928, w2929, w2930, w2931, w2932, w2933, w2934, w2935, w2936, w2937, w2938, w2939, w2940, w2941, w2942, w2943, w2944, w2945, w2946, w2947, w2948, w2949, w2950, w2951, w2952, w2953, w2954, w2955, w2956, w2957, w2958, w2959, w2960, w2961, w2962, w2963, w2964, w2965, w2966, w2967, w2968, w2969, w2970, w2971, w2972, w2973, w2974, w2975, w2976, w2977, w2978, w2979, w2980, w2981, w2982, w2983, w2984, w2985, w2986, w2987, w2988, w2989, w2990, w2991, w2992, w2993, w2994, w2995, w2996, w2997, w2998, w2999, w3000, w3001, w3002, w3003, w3004, w3005, w3006, w3007, w3008, w3009, w3010, w3011, w3012, w3013, w3014, w3015, w3016, w3017, w3018, w3019, w3020, w3021, w3022, w3023, w3024, w3025, w3026, w3027, w3028, w3029, w3030, w3031, w3032, w3033, w3034, w3035, w3036, w3037, w3038, w3039, w3040, w3041, w3042, w3043, w3044, w3045, w3046, w3047, w3048, w3049, w3050, w3051, w3052, w3053, w3054, w3055, w3056, w3057, w3058, w3059, w3060, w3061, w3062, w3063, w3064, w3065, w3066, w3067, w3068, w3069, w3070, w3071, w3072, w3073, w3074, w3075, w3076, w3077, w3078, w3079, w3080, w3081, w3082, w3083, w3084, w3085, w3086, w3087, w3088, w3089, w3090, w3091, w3092, w3093, w3094, w3095, w3096, w3097, w3098, w3099, w3100, w3101, w3102, w3103, w3104, w3105, w3106, w3107, w3108, w3109, w3110, w3111, w3112, w3113, w3114, w3115, w3116, w3117, w3118, w3119, w3120, w3121, w3122, w3123, w3124, w3125, w3126, w3127, w3128, w3129, w3130, w3131, w3132, w3133, w3134, w3135, w3136, w3137, w3138, w3139, w3140, w3141, w3142, w3143, w3144, w3145, w3146, w3147, w3148, w3149, w3150, w3151, w3152, w3153, w3154, w3155, w3156, w3157, w3158, w3159, w3160, w3161, w3162, w3163, w3164, w3165, w3166, w3167, w3168, w3169, w3170, w3171, w3172, w3173, w3174, w3175, w3176, w3177, w3178, w3179, w3180, w3181, w3182, w3183, w3184, w3185, w3186, w3187, w3188, w3189, w3190, w3191, w3192, w3193, w3194, w3195, w3196, w3197, w3198, w3199, w3200, w3201, w3202, w3203, w3204, w3205, w3206, w3207, w3208, w3209, w3210, w3211, w3212, w3213, w3214, w3215, w3216, w3217, w3218, w3219, w3220, w3221, w3222, w3223, w3224, w3225, w3226, w3227, w3228, w3229, w3230, w3231, w3232, w3233, w3234, w3235, w3236, w3237, w3238, w3239, w3240, w3241, w3242, w3243, w3244, w3245, w3246, w3247, w3248, w3249, w3250, w3251, w3252, w3253, w3254, w3255, w3256, w3257, w3258, w3259, w3260, w3261, w3262, w3263, w3264, w3265, w3266, w3267, w3268, w3269, w3270, w3271, w3272, w3273, w3274, w3275, w3276, w3277, w3278, w3279, w3280, w3281, w3282, w3283, w3284, w3285, w3286, w3287, w3288, w3289, w3290, w3291, w3292, w3293, w3294, w3295, w3296, w3297, w3298, w3299, w3300, w3301, w3302, w3303, w3304, w3305, w3306, w3307, w3308, w3309, w3310, w3311, w3312, w3313, w3314, w3315, w3316, w3317, w3318, w3319, w3320, w3321, w3322, w3323, w3324, w3325, w3326, w3327, w3328, w3329, w3330, w3331, w3332, w3333, w3334, w3335, w3336, w3337, w3338, w3339, w3340, w3341, w3342, w3343, w3344, w3345, w3346, w3347, w3348, w3349, w3350, w3351, w3352, w3353, w3354, w3355, w3356, w3357, w3358, w3359, w3360, w3361, w3362, w3363, w3364, w3365, w3366, w3367, w3368, w3369, w3370, w3371, w3372, w3373, w3374, w3375, w3376, w3377, w3378, w3379, w3380, w3381, w3382, w3383, w3384, w3385, w3386, w3387, w3388, w3389, w3390, w3391, w3392, w3393, w3394, w3395, w3396, w3397, w3398, w3399, w3400, w3401, w3402, w3403, w3404, w3405, w3406, w3407, w3408, w3409, w3410, w3411, w3412, w3413, w3414, w3415, w3416, w3417, w3418, w3419, w3420, w3421, w3422, w3423, w3424, w3425, w3426, w3427, w3428, w3429, w3430, w3431, w3432, w3433, w3434, w3435, w3436, w3437, w3438, w3439, w3440, w3441, w3442, w3443, w3444, w3445, w3446, w3447, w3448, w3449, w3450, w3451, w3452, w3453, w3454, w3455, w3456, w3457, w3458, w3459, w3460, w3461, w3462, w3463, w3464, w3465, w3466, w3467, w3468, w3469, w3470, w3471, w3472, w3473, w3474, w3475, w3476, w3477, w3478, w3479, w3480, w3481, w3482, w3483, w3484, w3485, w3486, w3487, w3488, w3489, w3490, w3491, w3492, w3493, w3494, w3495, w3496, w3497, w3498, w3499, w3500, w3501, w3502, w3503, w3504, w3505, w3506, w3507, w3508, w3509, w3510, w3511, w3512, w3513, w3514, w3515, w3516, w3517, w3518, w3519, w3520, w3521, w3522, w3523, w3524, w3525, w3526, w3527, w3528, w3529, w3530, w3531, w3532, w3533, w3534, w3535, w3536, w3537, w3538, w3539, w3540, w3541, w3542, w3543, w3544, w3545, w3546, w3547, w3548, w3549, w3550, w3551, w3552, w3553, w3554, w3555, w3556, w3557, w3558, w3559, w3560, w3561, w3562, w3563, w3564, w3565, w3566, w3567, w3568, w3569, w3570, w3571, w3572, w3573, w3574, w3575, w3576, w3577, w3578, w3579, w3580, w3581, w3582, w3583, w3584, w3585, w3586, w3587, w3588, w3589, w3590, w3591, w3592, w3593, w3594, w3595, w3596, w3597, w3598, w3599, w3600, w3601, w3602, w3603, w3604, w3605, w3606, w3607, w3608, w3609, w3610, w3611, w3612, w3613, w3614, w3615, w3616, w3617, w3618, w3619, w3620, w3621, w3622, w3623, w3624, w3625, w3626, w3627, w3628, w3629, w3630, w3631, w3632, w3633, w3634, w3635, w3636, w3637, w3638, w3639, w3640, w3641, w3642, w3643, w3644, w3645, w3646, w3647, w3648, w3649, w3650, w3651, w3652, w3653, w3654, w3655, w3656, w3657, w3658, w3659, w3660, w3661, w3662, w3663, w3664, w3665, w3666, w3667, w3668, w3669, w3670, w3671, w3672, w3673, w3674, w3675, w3676, w3677, w3678, w3679, w3680, w3681, w3682, w3683, w3684, w3685, w3686, w3687, w3688, w3689, w3690, w3691, w3692, w3693, w3694, w3695, w3696, w3697, w3698, w3699, w3700, w3701, w3702, w3703, w3704, w3705, w3706, w3707, w3708, w3709, w3710, w3711, w3712, w3713, w3714, w3715, w3716, w3717, w3718, w3719, w3720, w3721, w3722, w3723, w3724, w3725, w3726, w3727, w3728, w3729, w3730, w3731, w3732, w3733, w3734, w3735, w3736, w3737, w3738, w3739, w3740, w3741, w3742, w3743, w3744, w3745, w3746, w3747, w3748, w3749, w3750, w3751, w3752, w3753, w3754, w3755, w3756, w3757, w3758, w3759, w3760, w3761, w3762, w3763, w3764, w3765, w3766, w3767, w3768, w3769, w3770, w3771, w3772, w3773, w3774, w3775, w3776, w3777, w3778, w3779, w3780, w3781, w3782, w3783, w3784, w3785, w3786, w3787, w3788, w3789, w3790, w3791, w3792, w3793, w3794, w3795, w3796, w3797, w3798, w3799, w3800, w3801, w3802, w3803, w3804, w3805, w3806, w3807, w3808, w3809, w3810, w3811, w3812, w3813, w3814, w3815, w3816, w3817, w3818, w3819, w3820, w3821, w3822, w3823, w3824, w3825, w3826, w3827, w3828, w3829, w3830, w3831, w3832, w3833, w3834, w3835, w3836, w3837, w3838, w3839, w3840, w3841, w3842, w3843, w3844, w3845, w3846, w3847, w3848, w3849, w3850, w3851, w3852, w3853, w3854, w3855, w3856, w3857, w3858, w3859, w3860, w3861, w3862, w3863, w3864, w3865, w3866, w3867, w3868, w3869, w3870, w3871, w3872, w3873, w3874, w3875, w3876, w3877, w3878, w3879, w3880, w3881, w3882, w3883, w3884, w3885, w3886, w3887, w3888, w3889, w3890, w3891, w3892, w3893, w3894, w3895, w3896, w3897, w3898, w3899, w3900, w3901, w3902, w3903, w3904, w3905, w3906, w3907, w3908, w3909, w3910, w3911, w3912, w3913, w3914, w3915, w3916, w3917, w3918, w3919, w3920, w3921, w3922, w3923, w3924, w3925, w3926, w3927, w3928, w3929, w3930, w3931, w3932, w3933, w3934, w3935, w3936, w3937, w3938, w3939, w3940, w3941, w3942, w3943, w3944, w3945, w3946, w3947, w3948, w3949, w3950, w3951, w3952, w3953, w3954, w3955, w3956, w3957, w3958, w3959, w3960, w3961, w3962, w3963, w3964, w3965, w3966, w3967, w3968, w3969, w3970, w3971, w3972, w3973, w3974, w3975, w3976, w3977, w3978, w3979, w3980, w3981, w3982, w3983, w3984, w3985, w3986, w3987, w3988, w3989, w3990, w3991, w3992, w3993, w3994, w3995, w3996, w3997, w3998, w3999, w4000, w4001, w4002, w4003, w4004, w4005, w4006, w4007, w4008, w4009, w4010, w4011, w4012, w4013, w4014, w4015, w4016, w4017, w4018, w4019, w4020, w4021, w4022, w4023, w4024, w4025, w4026, w4027, w4028, w4029, w4030, w4031, w4032, w4033, w4034, w4035, w4036, w4037, w4038, w4039, w4040, w4041, w4042, w4043, w4044, w4045, w4046, w4047, w4048, w4049, w4050, w4051, w4052, w4053, w4054, w4055, w4056, w4057, w4058, w4059, w4060, w4061, w4062, w4063, w4064, w4065, w4066, w4067, w4068, w4069, w4070, w4071, w4072, w4073, w4074, w4075, w4076, w4077, w4078, w4079, w4080, w4081, w4082, w4083, w4084, w4085, w4086, w4087, w4088, w4089, w4090, w4091, w4092, w4093, w4094, w4095, w4096, w4097, w4098, w4099, w4100, w4101, w4102, w4103, w4104, w4105, w4106, w4107, w4108, w4109, w4110, w4111, w4112, w4113, w4114, w4115, w4116, w4117, w4118, w4119, w4120, w4121, w4122, w4123, w4124, w4125, w4126, w4127, w4128, w4129, w4130, w4131, w4132, w4133, w4134, w4135, w4136, w4137, w4138, w4139, w4140, w4141, w4142, w4143, w4144, w4145, w4146, w4147, w4148, w4149, w4150, w4151, w4152, w4153, w4154, w4155, w4156, w4157, w4158, w4159, w4160, w4161, w4162, w4163, w4164, w4165, w4166, w4167, w4168, w4169, w4170, w4171, w4172, w4173, w4174, w4175, w4176, w4177, w4178, w4179, w4180, w4181, w4182, w4183, w4184, w4185, w4186, w4187, w4188, w4189, w4190, w4191, w4192, w4193, w4194, w4195, w4196, w4197, w4198, w4199, w4200, w4201, w4202, w4203, w4204, w4205, w4206, w4207, w4208, w4209, w4210, w4211, w4212, w4213, w4214, w4215, w4216, w4217, w4218, w4219, w4220, w4221, w4222, w4223, w4224, w4225, w4226, w4227, w4228, w4229, w4230, w4231, w4232, w4233, w4234, w4235, w4236, w4237, w4238, w4239, w4240, w4241, w4242, w4243, w4244, w4245, w4246, w4247, w4248, w4249, w4250, w4251, w4252, w4253, w4254, w4255, w4256, w4257, w4258, w4259, w4260, w4261, w4262, w4263, w4264, w4265, w4266, w4267, w4268, w4269, w4270, w4271, w4272, w4273, w4274, w4275, w4276, w4277, w4278, w4279, w4280, w4281, w4282, w4283, w4284, w4285, w4286, w4287, w4288, w4289, w4290, w4291, w4292, w4293, w4294, w4295, w4296, w4297, w4298, w4299, w4300, w4301, w4302, w4303, w4304, w4305, w4306, w4307, w4308, w4309, w4310, w4311, w4312, w4313, w4314, w4315, w4316, w4317, w4318, w4319, w4320, w4321, w4322, w4323, w4324, w4325, w4326, w4327, w4328, w4329, w4330, w4331, w4332, w4333, w4334, w4335, w4336, w4337, w4338, w4339, w4340, w4341, w4342, w4343, w4344, w4345, w4346, w4347, w4348, w4349, w4350, w4351, w4352, w4353, w4354, w4355, w4356, w4357, w4358, w4359, w4360, w4361, w4362, w4363, w4364, w4365, w4366, w4367, w4368, w4369, w4370, w4371, w4372, w4373, w4374, w4375, w4376, w4377, w4378, w4379, w4380, w4381, w4382, w4383, w4384, w4385, w4386, w4387, w4388, w4389, w4390, w4391, w4392, w4393, w4394, w4395, w4396, w4397, w4398, w4399, w4400, w4401, w4402, w4403, w4404, w4405, w4406, w4407, w4408, w4409, w4410, w4411, w4412, w4413, w4414, w4415, w4416, w4417, w4418, w4419, w4420, w4421, w4422, w4423, w4424, w4425, w4426, w4427, w4428, w4429, w4430, w4431, w4432, w4433, w4434, w4435, w4436, w4437, w4438, w4439, w4440, w4441, w4442, w4443, w4444, w4445, w4446, w4447, w4448, w4449, w4450, w4451, w4452, w4453, w4454, w4455, w4456, w4457, w4458, w4459, w4460, w4461, w4462, w4463, w4464, w4465, w4466, w4467, w4468, w4469, w4470, w4471, w4472, w4473, w4474, w4475, w4476, w4477, w4478, w4479, w4480, w4481, w4482, w4483, w4484, w4485, w4486, w4487, w4488, w4489, w4490, w4491, w4492, w4493, w4494, w4495, w4496, w4497, w4498, w4499, w4500, w4501, w4502, w4503, w4504, w4505, w4506, w4507, w4508, w4509, w4510, w4511, w4512, w4513, w4514, w4515, w4516, w4517, w4518, w4519, w4520, w4521, w4522, w4523, w4524, w4525, w4526, w4527, w4528, w4529, w4530, w4531, w4532, w4533, w4534, w4535, w4536, w4537, w4538, w4539, w4540, w4541, w4542, w4543, w4544, w4545, w4546, w4547, w4548, w4549, w4550, w4551, w4552, w4553, w4554, w4555, w4556, w4557, w4558, w4559, w4560, w4561, w4562, w4563, w4564, w4565, w4566, w4567, w4568, w4569, w4570, w4571, w4572, w4573, w4574, w4575, w4576, w4577, w4578, w4579, w4580, w4581, w4582, w4583, w4584, w4585, w4586, w4587, w4588, w4589, w4590, w4591, w4592, w4593, w4594, w4595, w4596, w4597, w4598, w4599, w4600, w4601, w4602, w4603, w4604, w4605, w4606, w4607, w4608, w4609, w4610, w4611, w4612, w4613, w4614, w4615, w4616, w4617, w4618, w4619, w4620, w4621, w4622, w4623, w4624, w4625, w4626, w4627, w4628, w4629, w4630, w4631, w4632, w4633, w4634, w4635, w4636, w4637, w4638, w4639, w4640, w4641, w4642, w4643, w4644, w4645, w4646, w4647, w4648, w4649, w4650, w4651, w4652, w4653, w4654, w4655, w4656, w4657, w4658, w4659, w4660, w4661, w4662, w4663, w4664, w4665, w4666, w4667, w4668, w4669, w4670, w4671, w4672, w4673, w4674, w4675, w4676, w4677, w4678, w4679, w4680, w4681, w4682, w4683, w4684, w4685, w4686, w4687, w4688, w4689, w4690, w4691, w4692, w4693, w4694, w4695, w4696, w4697, w4698, w4699, w4700, w4701, w4702, w4703, w4704, w4705, w4706, w4707, w4708, w4709, w4710, w4711, w4712, w4713, w4714, w4715, w4716, w4717, w4718, w4719, w4720, w4721, w4722, w4723, w4724, w4725, w4726, w4727, w4728, w4729, w4730, w4731, w4732, w4733, w4734, w4735, w4736, w4737, w4738, w4739, w4740, w4741, w4742, w4743, w4744, w4745, w4746, w4747, w4748, w4749, w4750, w4751, w4752, w4753, w4754, w4755, w4756, w4757, w4758, w4759, w4760, w4761, w4762, w4763, w4764, w4765, w4766, w4767, w4768, w4769, w4770, w4771, w4772, w4773, w4774, w4775, w4776, w4777, w4778, w4779, w4780, w4781, w4782, w4783, w4784, w4785, w4786, w4787, w4788, w4789, w4790, w4791, w4792, w4793, w4794, w4795, w4796, w4797, w4798, w4799, w4800, w4801, w4802, w4803, w4804, w4805, w4806, w4807, w4808, w4809, w4810, w4811, w4812, w4813, w4814, w4815, w4816, w4817, w4818, w4819, w4820, w4821, w4822, w4823, w4824, w4825, w4826, w4827, w4828, w4829, w4830, w4831, w4832, w4833, w4834, w4835, w4836, w4837, w4838, w4839, w4840, w4841, w4842, w4843, w4844, w4845, w4846, w4847, w4848, w4849, w4850, w4851, w4852, w4853, w4854, w4855, w4856, w4857, w4858, w4859, w4860, w4861, w4862, w4863, w4864, w4865, w4866, w4867, w4868, w4869, w4870, w4871, w4872, w4873, w4874, w4875, w4876, w4877, w4878, w4879, w4880, w4881, w4882, w4883, w4884, w4885, w4886, w4887, w4888, w4889, w4890, w4891, w4892, w4893, w4894, w4895, w4896, w4897, w4898, w4899, w4900, w4901, w4902, w4903, w4904, w4905, w4906, w4907, w4908, w4909, w4910, w4911, w4912, w4913, w4914, w4915, w4916, w4917, w4918, w4919, w4920, w4921, w4922, w4923, w4924, w4925, w4926, w4927, w4928, w4929, w4930, w4931, w4932, w4933, w4934, w4935, w4936, w4937, w4938, w4939, w4940, w4941, w4942, w4943, w4944, w4945, w4946, w4947, w4948, w4949, w4950, w4951, w4952, w4953, w4954, w4955, w4956, w4957, w4958, w4959, w4960, w4961, w4962, w4963, w4964, w4965, w4966, w4967, w4968, w4969, w4970, w4971, w4972, w4973, w4974, w4975, w4976, w4977, w4978, w4979, w4980, w4981, w4982, w4983, w4984, w4985, w4986, w4987, w4988, w4989, w4990, w4991, w4992, w4993, w4994, w4995, w4996, w4997, w4998, w4999, w5000, w5001, w5002, w5003, w5004, w5005, w5006, w5007, w5008, w5009, w5010, w5011, w5012, w5013, w5014, w5015, w5016, w5017, w5018, w5019, w5020, w5021, w5022, w5023, w5024, w5025, w5026, w5027, w5028, w5029, w5030, w5031, w5032, w5033, w5034, w5035, w5036, w5037, w5038, w5039, w5040, w5041, w5042, w5043, w5044, w5045, w5046, w5047, w5048, w5049, w5050, w5051, w5052, w5053, w5054, w5055, w5056, w5057, w5058, w5059, w5060, w5061, w5062, w5063, w5064, w5065, w5066, w5067, w5068, w5069, w5070, w5071, w5072, w5073, w5074, w5075, w5076, w5077, w5078, w5079, w5080, w5081, w5082, w5083, w5084, w5085, w5086, w5087, w5088, w5089, w5090, w5091, w5092, w5093, w5094, w5095, w5096, w5097, w5098, w5099, w5100, w5101, w5102, w5103, w5104, w5105, w5106, w5107, w5108, w5109, w5110, w5111, w5112, w5113, w5114, w5115, w5116, w5117, w5118, w5119, w5120, w5121, w5122, w5123, w5124, w5125, w5126, w5127, w5128, w5129, w5130, w5131, w5132, w5133, w5134, w5135, w5136, w5137, w5138, w5139, w5140, w5141, w5142, w5143, w5144, w5145, w5146, w5147, w5148, w5149, w5150, w5151, w5152, w5153, w5154, w5155, w5156, w5157, w5158, w5159, w5160, w5161, w5162, w5163, w5164, w5165, w5166, w5167, w5168, w5169, w5170, w5171, w5172, w5173, w5174, w5175, w5176, w5177, w5178, w5179, w5180, w5181, w5182, w5183, w5184, w5185, w5186, w5187, w5188, w5189, w5190, w5191, w5192, w5193, w5194, w5195, w5196, w5197, w5198, w5199, w5200, w5201, w5202, w5203, w5204, w5205, w5206, w5207, w5208, w5209, w5210, w5211, w5212, w5213, w5214, w5215, w5216, w5217, w5218, w5219, w5220, w5221, w5222, w5223, w5224, w5225, w5226, w5227, w5228, w5229, w5230, w5231, w5232, w5233, w5234, w5235, w5236, w5237, w5238, w5239, w5240, w5241, w5242, w5243, w5244, w5245, w5246, w5247, w5248, w5249, w5250, w5251, w5252, w5253, w5254, w5255, w5256, w5257, w5258, w5259, w5260, w5261, w5262, w5263, w5264, w5265, w5266, w5267, w5268, w5269, w5270, w5271, w5272, w5273, w5274, w5275, w5276, w5277, w5278, w5279, w5280, w5281, w5282, w5283, w5284, w5285, w5286, w5287, w5288, w5289, w5290, w5291, w5292, w5293, w5294, w5295, w5296, w5297, w5298, w5299, w5300, w5301, w5302, w5303, w5304, w5305, w5306, w5307, w5308, w5309, w5310, w5311, w5312, w5313, w5314, w5315, w5316, w5317, w5318, w5319, w5320, w5321, w5322, w5323, w5324, w5325, w5326, w5327, w5328, w5329, w5330, w5331, w5332, w5333, w5334, w5335, w5336, w5337, w5338, w5339, w5340, w5341, w5342, w5343, w5344, w5345, w5346, w5347, w5348, w5349, w5350, w5351, w5352, w5353, w5354, w5355, w5356, w5357, w5358, w5359, w5360, w5361, w5362, w5363, w5364, w5365, w5366, w5367, w5368, w5369, w5370, w5371, w5372, w5373, w5374, w5375, w5376, w5377, w5378, w5379, w5380, w5381, w5382, w5383, w5384, w5385, w5386, w5387, w5388, w5389, w5390, w5391, w5392, w5393, w5394, w5395, w5396, w5397, w5398, w5399, w5400, w5401, w5402, w5403, w5404, w5405, w5406, w5407, w5408, w5409, w5410, w5411, w5412, w5413, w5414, w5415, w5416, w5417, w5418, w5419, w5420, w5421, w5422, w5423, w5424, w5425, w5426, w5427, w5428, w5429, w5430, w5431, w5432, w5433, w5434, w5435, w5436, w5437, w5438, w5439, w5440, w5441, w5442, w5443, w5444, w5445, w5446, w5447, w5448, w5449, w5450, w5451, w5452, w5453, w5454, w5455, w5456, w5457, w5458, w5459, w5460, w5461, w5462, w5463, w5464, w5465, w5466, w5467, w5468, w5469, w5470, w5471, w5472, w5473, w5474, w5475, w5476, w5477, w5478, w5479, w5480, w5481, w5482, w5483, w5484, w5485, w5486, w5487, w5488, w5489, w5490, w5491, w5492, w5493, w5494, w5495, w5496, w5497, w5498, w5499, w5500, w5501, w5502, w5503, w5504, w5505, w5506, w5507, w5508, w5509, w5510, w5511, w5512, w5513, w5514, w5515, w5516, w5517, w5518, w5519, w5520, w5521, w5522, w5523, w5524, w5525, w5526, w5527, w5528, w5529, w5530, w5531, w5532, w5533, w5534, w5535, w5536, w5537, w5538, w5539, w5540, w5541, w5542, w5543, w5544, w5545, w5546, w5547, w5548, w5549, w5550, w5551, w5552, w5553, w5554, w5555, w5556, w5557, w5558, w5559, w5560, w5561, w5562, w5563, w5564, w5565, w5566, w5567, w5568, w5569, w5570, w5571, w5572, w5573, w5574, w5575, w5576, w5577, w5578, w5579, w5580, w5581, w5582, w5583, w5584, w5585, w5586, w5587, w5588, w5589, w5590, w5591, w5592, w5593, w5594, w5595, w5596, w5597, w5598, w5599, w5600, w5601, w5602, w5603, w5604, w5605, w5606, w5607, w5608, w5609, w5610, w5611, w5612, w5613, w5614, w5615, w5616, w5617, w5618, w5619, w5620, w5621, w5622, w5623, w5624, w5625, w5626, w5627, w5628, w5629, w5630, w5631, w5632, w5633, w5634, w5635, w5636, w5637, w5638, w5639, w5640, w5641, w5642, w5643, w5644, w5645, w5646, w5647, w5648, w5649, w5650, w5651, w5652, w5653, w5654, w5655, w5656, w5657, w5658, w5659, w5660, w5661, w5662, w5663, w5664, w5665, w5666, w5667, w5668, w5669, w5670, w5671, w5672, w5673, w5674, w5675, w5676, w5677, w5678, w5679, w5680, w5681, w5682, w5683, w5684, w5685, w5686, w5687, w5688, w5689, w5690, w5691, w5692, w5693, w5694, w5695, w5696, w5697, w5698, w5699, w5700, w5701, w5702, w5703, w5704, w5705, w5706, w5707, w5708, w5709, w5710, w5711, w5712, w5713, w5714, w5715, w5716, w5717, w5718, w5719, w5720, w5721, w5722, w5723, w5724, w5725, w5726, w5727, w5728, w5729, w5730, w5731, w5732, w5733, w5734, w5735, w5736, w5737, w5738, w5739, w5740, w5741, w5742, w5743, w5744, w5745, w5746, w5747, w5748, w5749, w5750, w5751, w5752, w5753, w5754, w5755, w5756, w5757, w5758, w5759, w5760, w5761, w5762, w5763, w5764, w5765, w5766, w5767, w5768, w5769, w5770, w5771, w5772, w5773, w5774, w5775, w5776, w5777, w5778, w5779, w5780, w5781, w5782, w5783, w5784, w5785, w5786, w5787, w5788, w5789, w5790, w5791, w5792, w5793, w5794, w5795, w5796, w5797, w5798, w5799, w5800, w5801, w5802, w5803, w5804, w5805, w5806, w5807, w5808, w5809, w5810, w5811, w5812, w5813, w5814, w5815, w5816, w5817, w5818, w5819, w5820, w5821, w5822, w5823, w5824, w5825, w5826, w5827, w5828, w5829, w5830, w5831, w5832, w5833, w5834, w5835, w5836, w5837, w5838, w5839, w5840, w5841, w5842, w5843, w5844, w5845, w5846, w5847, w5848, w5849, w5850, w5851, w5852, w5853, w5854, w5855, w5856, w5857, w5858, w5859, w5860, w5861, w5862, w5863, w5864, w5865, w5866, w5867, w5868, w5869, w5870, w5871, w5872, w5873, w5874, w5875, w5876, w5877, w5878, w5879, w5880, w5881, w5882, w5883, w5884, w5885, w5886, w5887, w5888, w5889, w5890, w5891, w5892, w5893, w5894, w5895, w5896, w5897, w5898, w5899, w5900, w5901, w5902, w5903, w5904, w5905, w5906, w5907, w5908, w5909, w5910, w5911, w5912, w5913, w5914, w5915, w5916, w5917, w5918, w5919, w5920, w5921, w5922, w5923, w5924, w5925, w5926, w5927, w5928, w5929, w5930, w5931, w5932, w5933, w5934, w5935, w5936, w5937, w5938, w5939, w5940, w5941, w5942, w5943, w5944, w5945, w5946, w5947, w5948, w5949, w5950, w5951, w5952, w5953, w5954, w5955, w5956, w5957, w5958, w5959, w5960, w5961, w5962, w5963, w5964, w5965, w5966, w5967, w5968, w5969, w5970, w5971, w5972, w5973, w5974, w5975, w5976, w5977, w5978, w5979, w5980, w5981, w5982, w5983, w5984, w5985, w5986, w5987, w5988, w5989, w5990, w5991, w5992, w5993, w5994, w5995, w5996, w5997, w5998, w5999, w6000, w6001, w6002, w6003, w6004, w6005, w6006, w6007, w6008, w6009, w6010, w6011, w6012, w6013, w6014, w6015, w6016, w6017, w6018, w6019, w6020, w6021, w6022, w6023, w6024, w6025, w6026, w6027, w6028, w6029, w6030, w6031, w6032, w6033, w6034, w6035, w6036, w6037, w6038, w6039, w6040, w6041, w6042, w6043, w6044, w6045, w6046, w6047, w6048, w6049, w6050, w6051, w6052, w6053, w6054, w6055, w6056, w6057, w6058, w6059, w6060, w6061, w6062, w6063, w6064, w6065, w6066, w6067, w6068, w6069, w6070, w6071, w6072, w6073, w6074, w6075, w6076, w6077, w6078, w6079, w6080, w6081, w6082, w6083, w6084, w6085, w6086, w6087, w6088, w6089, w6090, w6091, w6092, w6093, w6094, w6095, w6096, w6097, w6098, w6099, w6100, w6101, w6102, w6103, w6104, w6105, w6106, w6107, w6108, w6109, w6110, w6111, w6112, w6113, w6114, w6115, w6116, w6117, w6118, w6119, w6120, w6121, w6122, w6123, w6124, w6125, w6126, w6127, w6128, w6129, w6130, w6131, w6132, w6133, w6134, w6135, w6136, w6137, w6138, w6139, w6140, w6141, w6142, w6143, w6144, w6145, w6146, w6147, w6148, w6149, w6150, w6151, w6152, w6153, w6154, w6155, w6156, w6157, w6158, w6159, w6160, w6161, w6162, w6163, w6164, w6165, w6166, w6167, w6168, w6169, w6170, w6171, w6172, w6173, w6174, w6175, w6176, w6177, w6178, w6179, w6180, w6181, w6182, w6183, w6184, w6185, w6186, w6187, w6188, w6189, w6190, w6191, w6192, w6193, w6194, w6195, w6196, w6197, w6198, w6199, w6200, w6201, w6202, w6203, w6204, w6205, w6206, w6207, w6208, w6209, w6210, w6211, w6212, w6213, w6214, w6215, w6216, w6217, w6218, w6219, w6220, w6221, w6222, w6223, w6224, w6225, w6226, w6227, w6228, w6229, w6230, w6231, w6232, w6233, w6234, w6235, w6236, w6237, w6238, w6239, w6240, w6241, w6242, w6243, w6244, w6245, w6246, w6247, w6248, w6249, w6250, w6251, w6252, w6253, w6254, w6255, w6256, w6257, w6258, w6259, w6260, w6261, w6262, w6263, w6264, w6265, w6266, w6267, w6268, w6269, w6270, w6271, w6272, w6273, w6274, w6275, w6276, w6277, w6278, w6279, w6280, w6281, w6282, w6283, w6284, w6285, w6286, w6287, w6288, w6289, w6290, w6291, w6292, w6293, w6294, w6295, w6296, w6297, w6298, w6299, w6300, w6301, w6302, w6303, w6304, w6305, w6306, w6307, w6308, w6309, w6310, w6311, w6312, w6313, w6314, w6315, w6316, w6317, w6318, w6319, w6320, w6321, w6322, w6323, w6324, w6325, w6326, w6327, w6328, w6329, w6330, w6331, w6332, w6333, w6334, w6335, w6336, w6337, w6338, w6339, w6340, w6341, w6342, w6343, w6344, w6345, w6346, w6347, w6348, w6349, w6350, w6351, w6352, w6353, w6354, w6355, w6356, w6357, w6358, w6359, w6360, w6361, w6362, w6363, w6364, w6365, w6366, w6367, w6368, w6369, w6370, w6371, w6372, w6373, w6374, w6375, w6376, w6377, w6378, w6379, w6380, w6381, w6382, w6383, w6384, w6385, w6386, w6387, w6388, w6389, w6390, w6391, w6392, w6393, w6394, w6395, w6396, w6397, w6398, w6399, w6400, w6401, w6402, w6403, w6404, w6405, w6406, w6407, w6408, w6409, w6410, w6411, w6412, w6413, w6414, w6415, w6416, w6417, w6418, w6419, w6420, w6421, w6422, w6423, w6424, w6425, w6426, w6427, w6428, w6429, w6430, w6431, w6432, w6433, w6434, w6435, w6436, w6437, w6438, w6439, w6440, w6441, w6442, w6443, w6444, w6445, w6446, w6447, w6448, w6449, w6450, w6451, w6452, w6453, w6454, w6455, w6456, w6457, w6458, w6459, w6460, w6461, w6462, w6463, w6464, w6465, w6466, w6467, w6468, w6469, w6470, w6471, w6472, w6473, w6474, w6475, w6476, w6477, w6478, w6479, w6480, w6481, w6482, w6483, w6484, w6485, w6486, w6487, w6488, w6489, w6490, w6491, w6492, w6493, w6494, w6495, w6496, w6497, w6498, w6499, w6500, w6501, w6502, w6503, w6504, w6505, w6506, w6507, w6508, w6509, w6510, w6511, w6512, w6513, w6514, w6515, w6516, w6517, w6518, w6519, w6520, w6521, w6522, w6523, w6524, w6525, w6526, w6527, w6528, w6529, w6530, w6531, w6532, w6533, w6534, w6535, w6536, w6537, w6538, w6539, w6540, w6541, w6542, w6543, w6544, w6545, w6546, w6547, w6548, w6549, w6550, w6551, w6552, w6553, w6554, w6555, w6556, w6557, w6558, w6559, w6560, w6561, w6562, w6563, w6564, w6565, w6566, w6567, w6568, w6569, w6570, w6571, w6572, w6573, w6574, w6575, w6576, w6577, w6578, w6579, w6580, w6581, w6582, w6583, w6584, w6585, w6586, w6587, w6588, w6589, w6590, w6591, w6592, w6593, w6594, w6595, w6596, w6597, w6598, w6599, w6600, w6601, w6602, w6603, w6604, w6605, w6606, w6607, w6608, w6609, w6610, w6611, w6612, w6613, w6614, w6615, w6616, w6617, w6618, w6619, w6620, w6621, w6622, w6623, w6624, w6625, w6626, w6627, w6628, w6629, w6630, w6631, w6632, w6633, w6634, w6635, w6636, w6637, w6638, w6639, w6640, w6641, w6642, w6643, w6644, w6645, w6646, w6647, w6648, w6649, w6650, w6651, w6652, w6653, w6654, w6655, w6656, w6657, w6658, w6659, w6660, w6661, w6662, w6663, w6664, w6665, w6666, w6667, w6668, w6669, w6670, w6671, w6672, w6673, w6674, w6675, w6676, w6677, w6678, w6679, w6680, w6681, w6682, w6683, w6684, w6685, w6686, w6687, w6688, w6689, w6690, w6691, w6692, w6693, w6694, w6695, w6696, w6697, w6698, w6699, w6700, w6701, w6702, w6703, w6704, w6705, w6706, w6707, w6708, w6709, w6710, w6711, w6712, w6713, w6714, w6715, w6716, w6717, w6718, w6719, w6720, w6721, w6722, w6723, w6724, w6725, w6726, w6727, w6728, w6729, w6730, w6731, w6732, w6733, w6734, w6735, w6736, w6737, w6738, w6739, w6740, w6741, w6742, w6743, w6744, w6745, w6746, w6747, w6748, w6749, w6750, w6751, w6752, w6753, w6754, w6755, w6756, w6757, w6758, w6759, w6760, w6761, w6762, w6763, w6764, w6765, w6766, w6767, w6768, w6769, w6770, w6771, w6772, w6773, w6774, w6775, w6776, w6777, w6778, w6779, w6780, w6781, w6782, w6783, w6784, w6785, w6786, w6787, w6788, w6789, w6790, w6791, w6792, w6793, w6794, w6795, w6796, w6797, w6798, w6799, w6800, w6801, w6802, w6803, w6804, w6805, w6806, w6807, w6808, w6809, w6810, w6811, w6812, w6813, w6814, w6815, w6816, w6817, w6818, w6819, w6820, w6821, w6822, w6823, w6824, w6825, w6826, w6827, w6828, w6829, w6830, w6831, w6832, w6833, w6834, w6835, w6836, w6837, w6838, w6839, w6840, w6841, w6842, w6843, w6844, w6845, w6846, w6847, w6848, w6849, w6850, w6851, w6852, w6853, w6854, w6855, w6856, w6857, w6858, w6859, w6860, w6861, w6862, w6863, w6864, w6865, w6866, w6867, w6868, w6869, w6870, w6871, w6872, w6873, w6874, w6875, w6876, w6877, w6878, w6879, w6880, w6881, w6882, w6883, w6884, w6885, w6886, w6887, w6888, w6889, w6890, w6891, w6892, w6893, w6894, w6895, w6896, w6897, w6898, w6899, w6900, w6901, w6902, w6903, w6904, w6905, w6906, w6907, w6908, w6909, w6910, w6911, w6912, w6913, w6914, w6915, w6916, w6917, w6918, w6919, w6920, w6921, w6922, w6923, w6924, w6925, w6926, w6927, w6928, w6929, w6930, w6931, w6932, w6933, w6934, w6935, w6936, w6937, w6938, w6939, w6940, w6941, w6942, w6943, w6944, w6945, w6946, w6947, w6948, w6949, w6950, w6951, w6952, w6953, w6954, w6955, w6956, w6957, w6958, w6959, w6960, w6961, w6962, w6963, w6964, w6965, w6966, w6967, w6968, w6969, w6970, w6971, w6972, w6973, w6974, w6975, w6976, w6977, w6978, w6979, w6980, w6981, w6982, w6983, w6984, w6985, w6986, w6987, w6988, w6989, w6990, w6991, w6992, w6993, w6994, w6995, w6996, w6997, w6998, w6999, w7000, w7001, w7002, w7003, w7004, w7005, w7006, w7007, w7008, w7009, w7010, w7011, w7012, w7013, w7014, w7015, w7016, w7017, w7018, w7019, w7020, w7021, w7022, w7023, w7024, w7025, w7026, w7027, w7028, w7029, w7030, w7031, w7032, w7033, w7034, w7035, w7036, w7037, w7038, w7039, w7040, w7041, w7042, w7043, w7044, w7045, w7046, w7047, w7048, w7049, w7050, w7051, w7052, w7053, w7054, w7055, w7056, w7057, w7058, w7059, w7060, w7061, w7062, w7063, w7064, w7065, w7066, w7067, w7068, w7069, w7070, w7071, w7072, w7073, w7074, w7075, w7076, w7077, w7078, w7079, w7080, w7081, w7082, w7083, w7084, w7085, w7086, w7087, w7088, w7089, w7090, w7091, w7092, w7093, w7094, w7095, w7096, w7097, w7098, w7099, w7100, w7101, w7102, w7103, w7104, w7105, w7106, w7107, w7108, w7109, w7110, w7111, w7112, w7113, w7114, w7115, w7116, w7117, w7118, w7119, w7120, w7121, w7122, w7123, w7124, w7125, w7126, w7127, w7128, w7129, w7130, w7131, w7132, w7133, w7134, w7135, w7136, w7137, w7138, w7139, w7140, w7141, w7142, w7143, w7144, w7145, w7146, w7147, w7148, w7149, w7150, w7151, w7152, w7153, w7154, w7155, w7156, w7157, w7158, w7159, w7160, w7161, w7162, w7163, w7164, w7165, w7166, w7167, w7168, w7169, w7170, w7171, w7172, w7173, w7174, w7175, w7176, w7177, w7178, w7179, w7180, w7181, w7182, w7183, w7184, w7185, w7186, w7187, w7188, w7189, w7190, w7191, w7192, w7193, w7194, w7195, w7196, w7197, w7198, w7199, w7200, w7201, w7202, w7203, w7204, w7205, w7206, w7207, w7208, w7209, w7210, w7211, w7212, w7213, w7214, w7215, w7216, w7217, w7218, w7219, w7220, w7221, w7222, w7223, w7224, w7225, w7226, w7227, w7228, w7229, w7230, w7231, w7232, w7233, w7234, w7235, w7236, w7237, w7238, w7239, w7240, w7241, w7242, w7243, w7244, w7245, w7246, w7247, w7248, w7249, w7250, w7251, w7252, w7253, w7254, w7255, w7256, w7257, w7258, w7259, w7260, w7261, w7262, w7263, w7264, w7265, w7266, w7267, w7268, w7269, w7270, w7271, w7272, w7273, w7274, w7275, w7276, w7277, w7278, w7279, w7280, w7281, w7282, w7283, w7284, w7285, w7286, w7287, w7288, w7289, w7290, w7291, w7292, w7293, w7294, w7295, w7296, w7297, w7298, w7299, w7300, w7301, w7302, w7303, w7304, w7305, w7306, w7307, w7308, w7309, w7310, w7311, w7312, w7313, w7314, w7315, w7316, w7317, w7318, w7319, w7320, w7321, w7322, w7323, w7324, w7325, w7326, w7327, w7328, w7329, w7330, w7331, w7332, w7333, w7334, w7335, w7336, w7337, w7338, w7339, w7340, w7341, w7342, w7343, w7344, w7345, w7346, w7347, w7348, w7349, w7350, w7351, w7352, w7353, w7354, w7355, w7356, w7357, w7358, w7359, w7360, w7361, w7362, w7363, w7364, w7365, w7366, w7367, w7368, w7369, w7370, w7371, w7372, w7373, w7374, w7375, w7376, w7377, w7378, w7379, w7380, w7381, w7382, w7383, w7384, w7385, w7386, w7387, w7388, w7389, w7390, w7391, w7392, w7393, w7394, w7395, w7396, w7397, w7398, w7399, w7400, w7401, w7402, w7403, w7404, w7405, w7406, w7407, w7408, w7409, w7410, w7411, w7412, w7413, w7414, w7415, w7416, w7417, w7418, w7419, w7420, w7421, w7422, w7423, w7424, w7425, w7426, w7427, w7428, w7429, w7430, w7431, w7432, w7433, w7434, w7435, w7436, w7437, w7438, w7439, w7440, w7441, w7442, w7443, w7444, w7445, w7446, w7447, w7448, w7449, w7450, w7451, w7452, w7453, w7454, w7455, w7456, w7457, w7458, w7459, w7460, w7461, w7462, w7463, w7464, w7465, w7466, w7467, w7468, w7469, w7470, w7471, w7472, w7473, w7474, w7475, w7476, w7477, w7478, w7479, w7480, w7481, w7482, w7483, w7484, w7485, w7486, w7487, w7488, w7489, w7490, w7491, w7492, w7493, w7494, w7495, w7496, w7497, w7498, w7499, w7500, w7501, w7502, w7503, w7504, w7505, w7506, w7507, w7508, w7509, w7510, w7511, w7512, w7513, w7514, w7515, w7516, w7517, w7518, w7519, w7520, w7521, w7522, w7523, w7524, w7525, w7526, w7527, w7528, w7529, w7530, w7531, w7532, w7533, w7534, w7535, w7536, w7537, w7538, w7539, w7540, w7541, w7542, w7543, w7544, w7545, w7546, w7547, w7548, w7549, w7550, w7551, w7552, w7553, w7554, w7555, w7556, w7557, w7558, w7559, w7560, w7561, w7562, w7563, w7564, w7565, w7566, w7567, w7568, w7569, w7570, w7571, w7572, w7573, w7574, w7575, w7576, w7577, w7578, w7579, w7580, w7581, w7582, w7583, w7584, w7585, w7586, w7587, w7588, w7589, w7590, w7591, w7592, w7593, w7594, w7595, w7596, w7597, w7598, w7599, w7600, w7601, w7602, w7603, w7604, w7605, w7606, w7607, w7608, w7609, w7610, w7611, w7612, w7613, w7614, w7615, w7616, w7617, w7618, w7619, w7620, w7621, w7622, w7623, w7624, w7625, w7626, w7627, w7628, w7629, w7630, w7631, w7632, w7633, w7634, w7635, w7636, w7637, w7638, w7639, w7640, w7641, w7642, w7643, w7644, w7645, w7646, w7647, w7648, w7649, w7650, w7651, w7652, w7653, w7654, w7655, w7656, w7657, w7658, w7659, w7660, w7661, w7662, w7663, w7664, w7665, w7666, w7667, w7668, w7669, w7670, w7671, w7672, w7673, w7674, w7675, w7676, w7677, w7678, w7679, w7680, w7681, w7682, w7683, w7684, w7685, w7686, w7687, w7688, w7689, w7690, w7691, w7692, w7693, w7694, w7695, w7696, w7697, w7698, w7699, w7700, w7701, w7702, w7703, w7704, w7705, w7706, w7707, w7708, w7709, w7710, w7711, w7712, w7713, w7714, w7715, w7716, w7717, w7718, w7719, w7720, w7721, w7722, w7723, w7724, w7725, w7726, w7727, w7728, w7729, w7730, w7731, w7732, w7733, w7734, w7735, w7736, w7737, w7738, w7739, w7740, w7741, w7742, w7743, w7744, w7745, w7746, w7747, w7748, w7749, w7750, w7751, w7752, w7753, w7754, w7755, w7756, w7757, w7758, w7759, w7760, w7761, w7762, w7763, w7764, w7765, w7766, w7767, w7768, w7769, w7770, w7771, w7772, w7773, w7774, w7775, w7776, w7777, w7778, w7779, w7780, w7781, w7782, w7783, w7784, w7785, w7786, w7787, w7788, w7789, w7790, w7791, w7792, w7793, w7794, w7795, w7796, w7797, w7798, w7799, w7800, w7801, w7802, w7803, w7804, w7805, w7806, w7807, w7808, w7809, w7810, w7811, w7812, w7813, w7814, w7815, w7816, w7817, w7818, w7819, w7820, w7821, w7822, w7823, w7824, w7825, w7826, w7827, w7828, w7829, w7830, w7831, w7832, w7833, w7834, w7835, w7836, w7837, w7838, w7839, w7840, w7841, w7842, w7843, w7844, w7845, w7846, w7847, w7848, w7849, w7850, w7851, w7852, w7853, w7854, w7855, w7856, w7857, w7858, w7859, w7860, w7861, w7862, w7863, w7864, w7865, w7866, w7867, w7868, w7869, w7870, w7871, w7872, w7873, w7874, w7875, w7876, w7877, w7878, w7879, w7880, w7881, w7882, w7883, w7884, w7885, w7886, w7887, w7888, w7889, w7890, w7891, w7892, w7893, w7894, w7895, w7896, w7897, w7898, w7899, w7900, w7901, w7902, w7903, w7904, w7905, w7906, w7907, w7908, w7909, w7910, w7911, w7912, w7913, w7914, w7915, w7916, w7917, w7918, w7919, w7920, w7921, w7922, w7923, w7924, w7925, w7926, w7927, w7928, w7929, w7930, w7931, w7932, w7933, w7934, w7935, w7936, w7937, w7938, w7939, w7940, w7941, w7942, w7943, w7944, w7945, w7946, w7947, w7948, w7949, w7950, w7951, w7952, w7953, w7954, w7955, w7956, w7957, w7958, w7959, w7960, w7961, w7962, w7963, w7964, w7965, w7966, w7967, w7968, w7969, w7970, w7971, w7972, w7973, w7974, w7975, w7976, w7977, w7978, w7979, w7980, w7981, w7982, w7983, w7984, w7985, w7986, w7987, w7988, w7989, w7990, w7991, w7992, w7993, w7994, w7995, w7996, w7997, w7998, w7999, w8000, w8001, w8002, w8003, w8004, w8005, w8006, w8007, w8008, w8009, w8010, w8011, w8012, w8013, w8014, w8015, w8016, w8017, w8018, w8019, w8020, w8021, w8022, w8023, w8024, w8025, w8026, w8027, w8028, w8029, w8030, w8031, w8032, w8033, w8034, w8035, w8036, w8037, w8038, w8039, w8040, w8041, w8042, w8043, w8044, w8045, w8046, w8047, w8048, w8049, w8050, w8051, w8052, w8053, w8054, w8055, w8056, w8057, w8058, w8059, w8060, w8061, w8062, w8063, w8064, w8065, w8066, w8067, w8068, w8069, w8070, w8071, w8072, w8073, w8074, w8075, w8076, w8077, w8078, w8079, w8080, w8081, w8082, w8083, w8084, w8085, w8086, w8087, w8088, w8089, w8090, w8091, w8092, w8093, w8094, w8095, w8096, w8097, w8098, w8099, w8100, w8101, w8102, w8103, w8104, w8105, w8106, w8107, w8108, w8109, w8110, w8111, w8112, w8113, w8114, w8115, w8116, w8117, w8118, w8119, w8120, w8121, w8122, w8123, w8124, w8125, w8126, w8127, w8128, w8129, w8130, w8131, w8132, w8133, w8134, w8135, w8136, w8137, w8138, w8139, w8140, w8141, w8142, w8143, w8144, w8145, w8146, w8147, w8148, w8149, w8150, w8151, w8152, w8153, w8154, w8155, w8156, w8157, w8158, w8159, w8160, w8161, w8162, w8163, w8164, w8165, w8166, w8167, w8168, w8169, w8170, w8171, w8172, w8173, w8174, w8175, w8176, w8177, w8178, w8179, w8180, w8181, w8182, w8183, w8184, w8185, w8186, w8187, w8188, w8189, w8190, w8191, w8192, w8193, w8194, w8195, w8196, w8197, w8198, w8199, w8200, w8201, w8202, w8203, w8204, w8205, w8206, w8207, w8208, w8209, w8210, w8211, w8212, w8213, w8214, w8215, w8216, w8217, w8218, w8219, w8220, w8221, w8222, w8223, w8224, w8225, w8226, w8227, w8228, w8229, w8230, w8231, w8232, w8233, w8234, w8235, w8236, w8237, w8238, w8239, w8240, w8241, w8242, w8243, w8244, w8245, w8246, w8247, w8248, w8249, w8250, w8251, w8252, w8253, w8254, w8255, w8256, w8257, w8258, w8259, w8260, w8261, w8262, w8263, w8264, w8265, w8266, w8267, w8268, w8269, w8270, w8271, w8272, w8273, w8274, w8275, w8276, w8277, w8278, w8279, w8280, w8281, w8282, w8283, w8284, w8285, w8286, w8287, w8288, w8289, w8290, w8291, w8292, w8293, w8294, w8295, w8296, w8297, w8298, w8299, w8300, w8301, w8302, w8303, w8304, w8305, w8306, w8307, w8308, w8309, w8310, w8311, w8312, w8313, w8314, w8315, w8316, w8317, w8318, w8319, w8320, w8321, w8322, w8323, w8324, w8325, w8326, w8327, w8328, w8329, w8330, w8331, w8332, w8333, w8334, w8335, w8336, w8337, w8338, w8339, w8340, w8341, w8342, w8343, w8344, w8345, w8346, w8347, w8348, w8349, w8350, w8351, w8352, w8353, w8354, w8355, w8356, w8357, w8358, w8359, w8360, w8361, w8362, w8363, w8364, w8365, w8366, w8367, w8368, w8369, w8370, w8371, w8372, w8373, w8374, w8375, w8376, w8377, w8378, w8379, w8380, w8381, w8382, w8383, w8384, w8385, w8386, w8387, w8388, w8389, w8390, w8391, w8392, w8393, w8394, w8395, w8396, w8397, w8398, w8399, w8400, w8401, w8402, w8403, w8404, w8405, w8406, w8407, w8408, w8409, w8410, w8411, w8412, w8413, w8414, w8415, w8416, w8417, w8418, w8419, w8420, w8421, w8422, w8423, w8424, w8425, w8426, w8427, w8428, w8429, w8430, w8431, w8432, w8433, w8434, w8435, w8436, w8437, w8438, w8439, w8440, w8441, w8442, w8443, w8444, w8445, w8446, w8447, w8448, w8449, w8450, w8451, w8452, w8453, w8454, w8455, w8456, w8457, w8458, w8459, w8460, w8461, w8462, w8463, w8464, w8465, w8466, w8467, w8468, w8469, w8470, w8471, w8472, w8473, w8474, w8475, w8476, w8477, w8478, w8479, w8480, w8481, w8482, w8483, w8484, w8485, w8486, w8487, w8488, w8489, w8490, w8491, w8492, w8493, w8494, w8495, w8496, w8497, w8498, w8499, w8500, w8501, w8502, w8503, w8504, w8505, w8506, w8507, w8508, w8509, w8510, w8511, w8512, w8513, w8514, w8515, w8516, w8517, w8518, w8519, w8520, w8521, w8522, w8523, w8524, w8525, w8526, w8527, w8528, w8529, w8530, w8531, w8532, w8533, w8534, w8535, w8536, w8537, w8538, w8539, w8540, w8541, w8542, w8543, w8544, w8545, w8546, w8547, w8548, w8549, w8550, w8551, w8552, w8553, w8554, w8555, w8556, w8557, w8558, w8559, w8560, w8561, w8562, w8563, w8564, w8565, w8566, w8567, w8568, w8569, w8570, w8571, w8572, w8573, w8574, w8575, w8576, w8577, w8578, w8579, w8580, w8581, w8582, w8583, w8584, w8585, w8586, w8587, w8588, w8589, w8590, w8591, w8592, w8593, w8594, w8595, w8596, w8597, w8598, w8599, w8600, w8601, w8602, w8603, w8604, w8605, w8606, w8607, w8608, w8609, w8610, w8611, w8612, w8613, w8614, w8615, w8616, w8617, w8618, w8619, w8620, w8621, w8622, w8623, w8624, w8625, w8626, w8627, w8628, w8629, w8630, w8631, w8632, w8633, w8634, w8635, w8636, w8637, w8638, w8639, w8640, w8641, w8642, w8643, w8644, w8645, w8646, w8647, w8648, w8649, w8650, w8651, w8652, w8653, w8654, w8655, w8656, w8657, w8658, w8659, w8660, w8661, w8662, w8663, w8664, w8665, w8666, w8667, w8668, w8669, w8670, w8671, w8672, w8673, w8674, w8675, w8676, w8677, w8678, w8679, w8680, w8681, w8682, w8683, w8684, w8685, w8686, w8687, w8688, w8689, w8690, w8691, w8692, w8693, w8694, w8695, w8696, w8697, w8698, w8699, w8700, w8701, w8702, w8703, w8704, w8705, w8706, w8707, w8708, w8709, w8710, w8711, w8712, w8713, w8714, w8715, w8716, w8717, w8718, w8719, w8720, w8721, w8722, w8723, w8724, w8725, w8726, w8727, w8728, w8729, w8730, w8731, w8732, w8733, w8734, w8735, w8736, w8737, w8738, w8739, w8740, w8741, w8742, w8743, w8744, w8745, w8746, w8747, w8748, w8749, w8750, w8751, w8752, w8753, w8754, w8755, w8756, w8757, w8758, w8759, w8760, w8761, w8762, w8763, w8764, w8765, w8766, w8767, w8768, w8769, w8770, w8771, w8772, w8773, w8774, w8775, w8776, w8777, w8778, w8779, w8780, w8781, w8782, w8783, w8784, w8785, w8786, w8787, w8788, w8789, w8790, w8791, w8792, w8793, w8794, w8795, w8796, w8797, w8798, w8799, w8800, w8801, w8802, w8803, w8804, w8805, w8806, w8807, w8808, w8809, w8810, w8811, w8812, w8813, w8814, w8815, w8816, w8817, w8818, w8819, w8820, w8821, w8822, w8823, w8824, w8825, w8826, w8827, w8828, w8829, w8830, w8831, w8832, w8833, w8834, w8835, w8836, w8837, w8838, w8839, w8840, w8841, w8842, w8843, w8844, w8845, w8846, w8847, w8848, w8849, w8850, w8851, w8852, w8853, w8854, w8855, w8856, w8857, w8858, w8859, w8860, w8861, w8862, w8863, w8864, w8865, w8866, w8867, w8868, w8869, w8870, w8871, w8872, w8873, w8874, w8875, w8876, w8877, w8878, w8879, w8880, w8881, w8882, w8883, w8884, w8885, w8886, w8887, w8888, w8889, w8890, w8891, w8892, w8893, w8894, w8895, w8896, w8897, w8898, w8899, w8900, w8901, w8902, w8903, w8904, w8905, w8906, w8907, w8908, w8909, w8910, w8911, w8912, w8913, w8914, w8915, w8916, w8917, w8918, w8919, w8920, w8921, w8922, w8923, w8924, w8925, w8926, w8927, w8928, w8929, w8930, w8931, w8932, w8933, w8934, w8935, w8936, w8937, w8938, w8939, w8940, w8941, w8942, w8943, w8944, w8945, w8946, w8947, w8948, w8949, w8950, w8951, w8952, w8953, w8954, w8955, w8956, w8957, w8958, w8959, w8960, w8961, w8962, w8963, w8964, w8965, w8966, w8967, w8968, w8969, w8970, w8971, w8972, w8973, w8974, w8975, w8976, w8977, w8978, w8979, w8980, w8981, w8982, w8983, w8984, w8985, w8986, w8987, w8988, w8989, w8990, w8991, w8992, w8993, w8994, w8995, w8996, w8997, w8998, w8999, w9000, w9001, w9002, w9003, w9004, w9005, w9006, w9007, w9008, w9009, w9010, w9011, w9012, w9013, w9014, w9015, w9016, w9017, w9018, w9019, w9020, w9021, w9022, w9023, w9024, w9025, w9026, w9027, w9028, w9029, w9030, w9031, w9032, w9033, w9034, w9035, w9036, w9037, w9038, w9039, w9040, w9041, w9042, w9043, w9044, w9045, w9046, w9047, w9048, w9049, w9050, w9051, w9052, w9053, w9054, w9055, w9056, w9057, w9058, w9059, w9060, w9061, w9062, w9063, w9064, w9065, w9066, w9067, w9068, w9069, w9070, w9071, w9072, w9073, w9074, w9075, w9076, w9077, w9078, w9079, w9080, w9081, w9082, w9083, w9084, w9085, w9086, w9087, w9088, w9089, w9090, w9091, w9092, w9093, w9094, w9095, w9096, w9097, w9098, w9099, w9100, w9101, w9102, w9103, w9104, w9105, w9106, w9107, w9108, w9109, w9110, w9111, w9112, w9113, w9114, w9115, w9116, w9117, w9118, w9119, w9120, w9121, w9122, w9123, w9124, w9125, w9126, w9127, w9128, w9129, w9130, w9131, w9132, w9133, w9134, w9135, w9136, w9137, w9138, w9139, w9140, w9141, w9142, w9143, w9144, w9145, w9146, w9147, w9148, w9149, w9150, w9151, w9152, w9153, w9154, w9155, w9156, w9157, w9158, w9159, w9160, w9161, w9162, w9163, w9164, w9165, w9166, w9167, w9168, w9169, w9170, w9171, w9172, w9173, w9174, w9175, w9176, w9177, w9178, w9179, w9180, w9181, w9182, w9183, w9184, w9185, w9186, w9187, w9188, w9189, w9190, w9191, w9192, w9193, w9194, w9195, w9196, w9197, w9198, w9199, w9200, w9201, w9202, w9203, w9204, w9205, w9206, w9207, w9208, w9209, w9210, w9211, w9212, w9213, w9214, w9215, w9216, w9217, w9218, w9219, w9220, w9221, w9222, w9223, w9224, w9225, w9226, w9227, w9228, w9229, w9230, w9231, w9232, w9233, w9234, w9235, w9236, w9237, w9238, w9239, w9240, w9241, w9242, w9243, w9244, w9245, w9246, w9247, w9248, w9249, w9250, w9251, w9252, w9253, w9254, w9255, w9256, w9257, w9258, w9259, w9260, w9261, w9262, w9263, w9264, w9265, w9266, w9267, w9268, w9269, w9270, w9271, w9272, w9273, w9274, w9275, w9276, w9277, w9278, w9279, w9280, w9281, w9282, w9283, w9284, w9285, w9286, w9287, w9288, w9289, w9290, w9291, w9292, w9293, w9294, w9295, w9296, w9297, w9298, w9299, w9300, w9301, w9302, w9303, w9304, w9305, w9306, w9307, w9308, w9309, w9310, w9311, w9312, w9313, w9314, w9315, w9316, w9317, w9318, w9319, w9320, w9321, w9322, w9323, w9324, w9325, w9326, w9327, w9328, w9329, w9330, w9331, w9332, w9333, w9334, w9335, w9336, w9337, w9338, w9339, w9340, w9341, w9342, w9343, w9344, w9345, w9346, w9347, w9348, w9349, w9350, w9351, w9352, w9353, w9354, w9355, w9356, w9357, w9358, w9359, w9360, w9361, w9362, w9363, w9364, w9365, w9366, w9367, w9368, w9369, w9370, w9371, w9372, w9373, w9374, w9375, w9376, w9377, w9378, w9379, w9380, w9381, w9382, w9383, w9384, w9385, w9386, w9387, w9388, w9389, w9390, w9391, w9392, w9393, w9394, w9395, w9396, w9397, w9398, w9399, w9400, w9401, w9402, w9403, w9404, w9405, w9406, w9407, w9408, w9409, w9410, w9411, w9412, w9413, w9414, w9415, w9416, w9417, w9418, w9419, w9420, w9421, w9422, w9423, w9424, w9425, w9426, w9427, w9428, w9429, w9430, w9431, w9432, w9433, w9434, w9435, w9436, w9437, w9438, w9439, w9440, w9441, w9442, w9443, w9444, w9445, w9446, w9447, w9448, w9449, w9450, w9451, w9452, w9453, w9454, w9455, w9456, w9457, w9458, w9459, w9460, w9461, w9462, w9463, w9464, w9465, w9466, w9467, w9468, w9469, w9470, w9471, w9472, w9473, w9474, w9475, w9476, w9477, w9478, w9479, w9480, w9481, w9482, w9483, w9484, w9485, w9486, w9487, w9488, w9489, w9490, w9491, w9492, w9493, w9494, w9495, w9496, w9497, w9498, w9499, w9500, w9501, w9502, w9503, w9504, w9505, w9506, w9507, w9508, w9509, w9510, w9511, w9512, w9513, w9514, w9515, w9516, w9517, w9518, w9519, w9520, w9521, w9522, w9523, w9524, w9525, w9526, w9527, w9528, w9529, w9530, w9531, w9532, w9533, w9534, w9535, w9536, w9537, w9538, w9539, w9540, w9541, w9542, w9543, w9544, w9545, w9546, w9547, w9548, w9549, w9550, w9551, w9552, w9553, w9554, w9555, w9556, w9557, w9558, w9559, w9560, w9561, w9562, w9563, w9564, w9565, w9566, w9567, w9568, w9569, w9570, w9571, w9572, w9573, w9574, w9575, w9576, w9577, w9578, w9579, w9580, w9581, w9582, w9583, w9584, w9585, w9586, w9587, w9588, w9589, w9590, w9591, w9592, w9593, w9594, w9595, w9596, w9597, w9598, w9599, w9600, w9601, w9602, w9603, w9604, w9605, w9606, w9607, w9608, w9609, w9610, w9611, w9612, w9613, w9614, w9615, w9616, w9617, w9618, w9619, w9620, w9621, w9622, w9623, w9624, w9625, w9626, w9627, w9628, w9629, w9630, w9631, w9632, w9633, w9634, w9635, w9636, w9637, w9638, w9639, w9640, w9641, w9642, w9643, w9644, w9645, w9646, w9647, w9648, w9649, w9650, w9651, w9652, w9653, w9654, w9655, w9656, w9657, w9658, w9659, w9660, w9661, w9662, w9663, w9664, w9665, w9666, w9667, w9668, w9669, w9670, w9671, w9672, w9673, w9674, w9675, w9676, w9677, w9678, w9679, w9680, w9681, w9682, w9683, w9684, w9685, w9686, w9687, w9688, w9689, w9690, w9691, w9692, w9693, w9694, w9695, w9696, w9697, w9698, w9699, w9700, w9701, w9702, w9703, w9704, w9705, w9706, w9707, w9708, w9709, w9710, w9711, w9712, w9713, w9714, w9715, w9716, w9717, w9718, w9719, w9720, w9721, w9722, w9723, w9724, w9725, w9726, w9727, w9728, w9729, w9730, w9731, w9732, w9733, w9734, w9735, w9736, w9737, w9738, w9739, w9740, w9741, w9742, w9743, w9744, w9745, w9746, w9747, w9748, w9749, w9750, w9751, w9752, w9753, w9754, w9755, w9756, w9757, w9758, w9759, w9760, w9761, w9762, w9763, w9764, w9765, w9766, w9767, w9768, w9769, w9770, w9771, w9772, w9773, w9774, w9775, w9776, w9777, w9778, w9779, w9780, w9781, w9782, w9783, w9784, w9785, w9786, w9787, w9788, w9789, w9790, w9791, w9792, w9793, w9794, w9795, w9796, w9797, w9798, w9799, w9800, w9801, w9802, w9803, w9804, w9805, w9806, w9807, w9808, w9809, w9810, w9811, w9812, w9813, w9814, w9815, w9816, w9817, w9818, w9819, w9820, w9821, w9822, w9823, w9824, w9825, w9826, w9827, w9828, w9829, w9830, w9831, w9832, w9833, w9834, w9835, w9836, w9837, w9838, w9839, w9840, w9841, w9842, w9843, w9844, w9845, w9846, w9847, w9848, w9849, w9850, w9851, w9852, w9853, w9854, w9855, w9856, w9857, w9858, w9859, w9860, w9861, w9862, w9863, w9864, w9865, w9866, w9867, w9868, w9869, w9870, w9871, w9872, w9873, w9874, w9875, w9876, w9877, w9878, w9879, w9880, w9881, w9882, w9883, w9884, w9885, w9886, w9887, w9888, w9889, w9890, w9891, w9892, w9893, w9894, w9895, w9896, w9897, w9898, w9899, w9900, w9901, w9902, w9903, w9904, w9905, w9906, w9907, w9908, w9909, w9910, w9911, w9912, w9913, w9914, w9915, w9916, w9917, w9918, w9919, w9920, w9921, w9922, w9923, w9924, w9925, w9926, w9927, w9928, w9929, w9930, w9931, w9932, w9933, w9934, w9935, w9936, w9937, w9938, w9939, w9940, w9941, w9942, w9943, w9944, w9945, w9946, w9947, w9948, w9949, w9950, w9951, w9952, w9953, w9954, w9955, w9956, w9957, w9958, w9959, w9960, w9961, w9962, w9963, w9964, w9965, w9966, w9967, w9968, w9969, w9970, w9971, w9972, w9973, w9974, w9975, w9976, w9977, w9978, w9979, w9980, w9981, w9982, w9983, w9984, w9985, w9986, w9987, w9988, w9989, w9990, w9991, w9992, w9993, w9994, w9995, w9996, w9997, w9998, w9999, w10000, w10001, w10002, w10003, w10004, w10005, w10006, w10007, w10008, w10009, w10010, w10011, w10012, w10013, w10014, w10015, w10016, w10017, w10018, w10019, w10020, w10021, w10022, w10023, w10024, w10025, w10026, w10027, w10028, w10029, w10030, w10031, w10032, w10033, w10034, w10035, w10036, w10037, w10038, w10039, w10040, w10041, w10042, w10043, w10044, w10045, w10046, w10047, w10048, w10049, w10050, w10051, w10052, w10053, w10054, w10055, w10056, w10057, w10058, w10059, w10060, w10061, w10062, w10063, w10064, w10065, w10066, w10067, w10068, w10069, w10070, w10071, w10072, w10073, w10074, w10075, w10076, w10077, w10078, w10079, w10080, w10081, w10082, w10083, w10084, w10085, w10086, w10087, w10088, w10089, w10090, w10091, w10092, w10093, w10094, w10095, w10096, w10097, w10098, w10099, w10100, w10101, w10102, w10103, w10104, w10105, w10106, w10107, w10108, w10109, w10110, w10111, w10112, w10113, w10114, w10115, w10116, w10117, w10118, w10119, w10120, w10121, w10122, w10123, w10124, w10125, w10126, w10127, w10128, w10129, w10130, w10131, w10132, w10133, w10134, w10135, w10136, w10137, w10138, w10139, w10140, w10141, w10142, w10143, w10144, w10145, w10146, w10147, w10148, w10149, w10150, w10151, w10152, w10153, w10154, w10155, w10156, w10157, w10158, w10159, w10160, w10161, w10162, w10163, w10164, w10165, w10166, w10167, w10168, w10169, w10170, w10171, w10172, w10173, w10174, w10175, w10176, w10177, w10178, w10179, w10180, w10181, w10182, w10183, w10184, w10185, w10186, w10187, w10188, w10189, w10190, w10191, w10192, w10193, w10194, w10195, w10196, w10197, w10198, w10199, w10200, w10201, w10202, w10203, w10204, w10205, w10206, w10207, w10208, w10209, w10210, w10211, w10212, w10213, w10214, w10215, w10216, w10217, w10218, w10219, w10220, w10221, w10222, w10223, w10224, w10225, w10226, w10227, w10228, w10229, w10230, w10231, w10232, w10233, w10234, w10235, w10236, w10237, w10238, w10239, w10240, w10241, w10242, w10243, w10244, w10245, w10246, w10247, w10248, w10249, w10250, w10251, w10252, w10253, w10254, w10255, w10256, w10257, w10258, w10259, w10260, w10261, w10262, w10263, w10264, w10265, w10266, w10267, w10268, w10269, w10270, w10271, w10272, w10273, w10274, w10275, w10276, w10277, w10278, w10279, w10280, w10281, w10282, w10283, w10284, w10285, w10286, w10287, w10288, w10289, w10290, w10291, w10292, w10293, w10294, w10295, w10296, w10297, w10298, w10299, w10300, w10301, w10302, w10303, w10304, w10305, w10306, w10307, w10308, w10309, w10310, w10311, w10312, w10313, w10314, w10315, w10316, w10317, w10318, w10319, w10320, w10321, w10322, w10323, w10324, w10325, w10326, w10327, w10328, w10329, w10330, w10331, w10332, w10333, w10334, w10335, w10336, w10337, w10338, w10339, w10340, w10341, w10342, w10343, w10344, w10345, w10346, w10347, w10348, w10349, w10350, w10351, w10352, w10353, w10354, w10355, w10356, w10357, w10358, w10359, w10360, w10361, w10362, w10363, w10364, w10365, w10366, w10367, w10368, w10369, w10370, w10371, w10372, w10373, w10374, w10375, w10376, w10377, w10378, w10379, w10380, w10381, w10382, w10383, w10384, w10385, w10386, w10387, w10388, w10389, w10390, w10391, w10392, w10393, w10394, w10395, w10396, w10397, w10398, w10399, w10400, w10401, w10402, w10403, w10404, w10405, w10406, w10407, w10408, w10409, w10410, w10411, w10412, w10413, w10414, w10415, w10416, w10417, w10418, w10419, w10420, w10421, w10422, w10423, w10424, w10425, w10426, w10427, w10428, w10429, w10430, w10431, w10432, w10433, w10434, w10435, w10436, w10437, w10438, w10439, w10440, w10441, w10442, w10443, w10444, w10445, w10446, w10447, w10448, w10449, w10450, w10451, w10452, w10453, w10454, w10455, w10456, w10457, w10458, w10459, w10460, w10461, w10462, w10463, w10464, w10465, w10466, w10467, w10468, w10469, w10470, w10471, w10472, w10473, w10474, w10475, w10476, w10477, w10478, w10479, w10480, w10481, w10482, w10483, w10484, w10485, w10486, w10487, w10488, w10489, w10490, w10491, w10492, w10493, w10494, w10495, w10496, w10497, w10498, w10499, w10500, w10501, w10502, w10503, w10504, w10505, w10506, w10507, w10508, w10509, w10510, w10511, w10512, w10513, w10514, w10515, w10516, w10517, w10518, w10519, w10520, w10521, w10522, w10523, w10524, w10525, w10526, w10527, w10528, w10529, w10530, w10531, w10532, w10533, w10534, w10535, w10536, w10537, w10538, w10539, w10540, w10541, w10542, w10543, w10544, w10545, w10546, w10547, w10548, w10549, w10550, w10551, w10552, w10553, w10554, w10555, w10556, w10557, w10558, w10559, w10560, w10561, w10562, w10563, w10564, w10565, w10566, w10567, w10568, w10569, w10570, w10571, w10572, w10573, w10574, w10575, w10576, w10577, w10578, w10579, w10580, w10581, w10582, w10583, w10584, w10585, w10586, w10587, w10588, w10589, w10590, w10591, w10592, w10593, w10594, w10595, w10596, w10597, w10598, w10599, w10600, w10601, w10602, w10603, w10604, w10605, w10606, w10607, w10608, w10609, w10610, w10611, w10612, w10613, w10614, w10615, w10616, w10617, w10618, w10619, w10620, w10621, w10622, w10623, w10624, w10625, w10626, w10627, w10628, w10629, w10630, w10631, w10632, w10633, w10634, w10635, w10636, w10637, w10638, w10639, w10640, w10641, w10642, w10643, w10644, w10645, w10646, w10647, w10648, w10649, w10650, w10651, w10652, w10653, w10654, w10655, w10656, w10657, w10658, w10659, w10660, w10661, w10662, w10663, w10664, w10665, w10666, w10667, w10668, w10669, w10670, w10671, w10672, w10673, w10674, w10675, w10676, w10677, w10678, w10679, w10680, w10681, w10682, w10683, w10684, w10685, w10686, w10687, w10688, w10689, w10690, w10691, w10692, w10693, w10694, w10695, w10696, w10697, w10698, w10699, w10700, w10701, w10702, w10703, w10704, w10705, w10706, w10707, w10708, w10709, w10710, w10711, w10712, w10713, w10714, w10715, w10716, w10717, w10718, w10719, w10720, w10721, w10722, w10723, w10724, w10725, w10726, w10727, w10728, w10729, w10730, w10731, w10732, w10733, w10734, w10735, w10736, w10737, w10738, w10739, w10740, w10741, w10742, w10743, w10744, w10745, w10746, w10747, w10748, w10749, w10750, w10751, w10752, w10753, w10754, w10755, w10756, w10757, w10758, w10759, w10760, w10761, w10762, w10763, w10764, w10765, w10766, w10767, w10768, w10769, w10770, w10771, w10772, w10773, w10774, w10775, w10776, w10777, w10778, w10779, w10780, w10781, w10782, w10783, w10784, w10785, w10786, w10787, w10788, w10789, w10790, w10791, w10792, w10793, w10794, w10795, w10796, w10797, w10798, w10799, w10800, w10801, w10802, w10803, w10804, w10805, w10806, w10807, w10808, w10809, w10810, w10811, w10812, w10813, w10814, w10815, w10816, w10817, w10818, w10819, w10820, w10821, w10822, w10823, w10824, w10825, w10826, w10827, w10828, w10829, w10830, w10831, w10832, w10833, w10834, w10835, w10836, w10837, w10838, w10839, w10840, w10841, w10842, w10843, w10844, w10845, w10846, w10847, w10848, w10849, w10850, w10851, w10852, w10853, w10854, w10855, w10856, w10857, w10858, w10859, w10860, w10861, w10862, w10863, w10864, w10865, w10866, w10867, w10868, w10869, w10870, w10871, w10872, w10873, w10874, w10875, w10876, w10877, w10878, w10879, w10880, w10881, w10882, w10883, w10884, w10885, w10886, w10887, w10888, w10889, w10890, w10891, w10892, w10893, w10894, w10895, w10896, w10897, w10898, w10899, w10900, w10901, w10902, w10903, w10904, w10905, w10906, w10907, w10908, w10909, w10910, w10911, w10912, w10913, w10914, w10915, w10916, w10917, w10918, w10919, w10920, w10921, w10922, w10923, w10924, w10925, w10926, w10927, w10928, w10929, w10930, w10931, w10932, w10933, w10934, w10935, w10936, w10937, w10938, w10939, w10940, w10941, w10942, w10943, w10944, w10945, w10946, w10947, w10948, w10949, w10950, w10951, w10952, w10953, w10954, w10955, w10956, w10957, w10958, w10959, w10960, w10961, w10962, w10963, w10964, w10965, w10966, w10967, w10968, w10969, w10970, w10971, w10972, w10973, w10974, w10975, w10976, w10977, w10978, w10979, w10980, w10981, w10982, w10983, w10984, w10985, w10986, w10987, w10988, w10989, w10990, w10991, w10992, w10993, w10994, w10995, w10996, w10997, w10998, w10999, w11000, w11001, w11002, w11003, w11004, w11005, w11006, w11007, w11008, w11009, w11010, w11011, w11012, w11013, w11014, w11015, w11016, w11017, w11018, w11019, w11020, w11021, w11022, w11023, w11024, w11025, w11026, w11027, w11028, w11029, w11030, w11031, w11032, w11033, w11034, w11035, w11036, w11037, w11038, w11039, w11040, w11041, w11042, w11043, w11044, w11045, w11046, w11047, w11048, w11049, w11050, w11051, w11052, w11053, w11054, w11055, w11056, w11057, w11058, w11059, w11060, w11061, w11062, w11063, w11064, w11065, w11066, w11067, w11068, w11069, w11070, w11071, w11072, w11073, w11074, w11075, w11076, w11077, w11078, w11079, w11080, w11081, w11082, w11083, w11084, w11085, w11086, w11087, w11088, w11089, w11090, w11091, w11092, w11093, w11094, w11095, w11096, w11097, w11098, w11099, w11100, w11101, w11102, w11103, w11104, w11105, w11106, w11107, w11108, w11109, w11110, w11111, w11112, w11113, w11114, w11115, w11116, w11117, w11118, w11119, w11120, w11121, w11122, w11123, w11124, w11125, w11126, w11127, w11128, w11129, w11130, w11131, w11132, w11133, w11134, w11135, w11136, w11137, w11138, w11139, w11140, w11141, w11142, w11143, w11144, w11145, w11146, w11147, w11148, w11149, w11150, w11151, w11152, w11153, w11154, w11155, w11156, w11157, w11158, w11159, w11160, w11161, w11162, w11163, w11164, w11165, w11166, w11167, w11168, w11169, w11170, w11171, w11172, w11173, w11174, w11175, w11176, w11177, w11178, w11179, w11180, w11181, w11182, w11183, w11184, w11185, w11186, w11187, w11188, w11189, w11190, w11191, w11192, w11193, w11194, w11195, w11196, w11197, w11198, w11199, w11200, w11201, w11202, w11203, w11204, w11205, w11206, w11207, w11208, w11209, w11210, w11211, w11212, w11213, w11214, w11215, w11216, w11217, w11218, w11219, w11220, w11221, w11222, w11223, w11224, w11225, w11226, w11227, w11228, w11229, w11230, w11231, w11232, w11233, w11234, w11235, w11236, w11237, w11238, w11239, w11240, w11241, w11242, w11243, w11244, w11245, w11246, w11247, w11248, w11249, w11250, w11251, w11252, w11253, w11254, w11255, w11256, w11257, w11258, w11259, w11260, w11261, w11262, w11263, w11264, w11265, w11266, w11267, w11268, w11269, w11270, w11271, w11272, w11273, w11274, w11275, w11276, w11277, w11278, w11279, w11280, w11281, w11282, w11283, w11284, w11285, w11286, w11287, w11288, w11289, w11290, w11291, w11292, w11293, w11294, w11295, w11296, w11297, w11298, w11299, w11300, w11301, w11302, w11303, w11304, w11305, w11306, w11307, w11308, w11309, w11310, w11311, w11312, w11313, w11314, w11315, w11316, w11317, w11318, w11319, w11320, w11321, w11322, w11323, w11324, w11325, w11326, w11327, w11328, w11329, w11330, w11331, w11332, w11333, w11334, w11335, w11336, w11337, w11338, w11339, w11340, w11341, w11342, w11343, w11344, w11345, w11346, w11347, w11348, w11349, w11350, w11351, w11352, w11353, w11354, w11355, w11356, w11357, w11358, w11359, w11360, w11361, w11362, w11363, w11364, w11365, w11366, w11367, w11368, w11369, w11370, w11371, w11372, w11373, w11374, w11375, w11376, w11377, w11378, w11379, w11380, w11381, w11382, w11383, w11384, w11385, w11386, w11387, w11388, w11389, w11390, w11391, w11392, w11393, w11394, w11395, w11396, w11397, w11398, w11399, w11400, w11401, w11402, w11403, w11404, w11405, w11406, w11407, w11408, w11409, w11410, w11411, w11412, w11413, w11414, w11415, w11416, w11417, w11418, w11419, w11420, w11421, w11422, w11423, w11424, w11425, w11426, w11427, w11428, w11429, w11430, w11431, w11432, w11433, w11434, w11435, w11436, w11437, w11438, w11439, w11440, w11441, w11442, w11443, w11444, w11445, w11446, w11447, w11448, w11449, w11450, w11451, w11452, w11453, w11454, w11455, w11456, w11457, w11458, w11459, w11460, w11461, w11462, w11463, w11464, w11465, w11466, w11467, w11468, w11469, w11470, w11471, w11472, w11473, w11474, w11475, w11476, w11477, w11478, w11479, w11480, w11481, w11482, w11483, w11484, w11485, w11486, w11487, w11488, w11489, w11490, w11491, w11492, w11493, w11494, w11495, w11496, w11497, w11498, w11499, w11500, w11501, w11502, w11503, w11504, w11505, w11506, w11507, w11508, w11509, w11510, w11511, w11512, w11513, w11514, w11515, w11516, w11517, w11518, w11519, w11520, w11521, w11522, w11523, w11524, w11525, w11526, w11527, w11528, w11529, w11530, w11531, w11532, w11533, w11534, w11535, w11536, w11537, w11538, w11539, w11540, w11541, w11542, w11543, w11544, w11545, w11546, w11547, w11548, w11549, w11550, w11551, w11552, w11553, w11554, w11555, w11556, w11557, w11558, w11559, w11560, w11561, w11562, w11563, w11564, w11565, w11566, w11567, w11568, w11569, w11570, w11571, w11572, w11573, w11574, w11575, w11576, w11577, w11578, w11579, w11580, w11581, w11582, w11583, w11584, w11585, w11586, w11587, w11588, w11589, w11590, w11591, w11592, w11593, w11594, w11595, w11596, w11597, w11598, w11599, w11600, w11601, w11602, w11603, w11604, w11605, w11606, w11607, w11608, w11609, w11610, w11611, w11612, w11613, w11614, w11615, w11616, w11617, w11618, w11619, w11620, w11621, w11622, w11623, w11624, w11625, w11626, w11627, w11628, w11629, w11630, w11631, w11632, w11633, w11634, w11635, w11636, w11637, w11638, w11639, w11640, w11641, w11642, w11643, w11644, w11645, w11646, w11647, w11648, w11649, w11650, w11651, w11652, w11653, w11654, w11655, w11656, w11657, w11658, w11659, w11660, w11661, w11662, w11663, w11664, w11665, w11666, w11667, w11668, w11669, w11670, w11671, w11672, w11673, w11674, w11675, w11676, w11677, w11678, w11679, w11680, w11681, w11682, w11683, w11684, w11685, w11686, w11687, w11688, w11689, w11690, w11691, w11692, w11693, w11694, w11695, w11696, w11697, w11698, w11699, w11700, w11701, w11702, w11703, w11704, w11705, w11706, w11707, w11708, w11709, w11710, w11711, w11712, w11713, w11714, w11715, w11716, w11717, w11718, w11719, w11720, w11721, w11722, w11723, w11724, w11725, w11726, w11727, w11728, w11729, w11730, w11731, w11732, w11733, w11734, w11735, w11736, w11737, w11738, w11739, w11740, w11741, w11742, w11743, w11744, w11745, w11746, w11747, w11748, w11749, w11750, w11751, w11752, w11753, w11754, w11755, w11756, w11757, w11758, w11759, w11760, w11761, w11762, w11763, w11764, w11765, w11766, w11767, w11768, w11769, w11770, w11771, w11772, w11773, w11774, w11775, w11776, w11777, w11778, w11779, w11780, w11781, w11782, w11783, w11784, w11785, w11786, w11787, w11788, w11789, w11790, w11791, w11792, w11793, w11794, w11795, w11796, w11797, w11798, w11799, w11800, w11801, w11802, w11803, w11804, w11805, w11806, w11807, w11808, w11809, w11810, w11811, w11812, w11813, w11814, w11815, w11816, w11817, w11818, w11819, w11820, w11821, w11822, w11823, w11824, w11825, w11826, w11827, w11828, w11829, w11830, w11831, w11832, w11833, w11834, w11835, w11836, w11837, w11838, w11839, w11840, w11841, w11842, w11843, w11844, w11845, w11846, w11847, w11848, w11849, w11850, w11851, w11852, w11853, w11854, w11855, w11856, w11857, w11858, w11859, w11860, w11861, w11862, w11863, w11864, w11865, w11866, w11867, w11868, w11869, w11870, w11871, w11872, w11873, w11874, w11875, w11876, w11877, w11878, w11879, w11880, w11881, w11882, w11883, w11884, w11885, w11886, w11887, w11888, w11889, w11890, w11891, w11892, w11893, w11894, w11895, w11896, w11897, w11898, w11899, w11900, w11901, w11902, w11903, w11904, w11905, w11906, w11907, w11908, w11909, w11910, w11911, w11912, w11913, w11914, w11915, w11916, w11917, w11918, w11919, w11920, w11921, w11922, w11923, w11924, w11925, w11926, w11927, w11928, w11929, w11930, w11931, w11932, w11933, w11934, w11935, w11936, w11937, w11938, w11939, w11940, w11941, w11942, w11943, w11944, w11945, w11946, w11947, w11948, w11949, w11950, w11951, w11952, w11953, w11954, w11955, w11956, w11957, w11958, w11959, w11960, w11961, w11962, w11963, w11964, w11965, w11966, w11967, w11968, w11969, w11970, w11971, w11972, w11973, w11974, w11975, w11976, w11977, w11978, w11979, w11980, w11981, w11982, w11983, w11984, w11985, w11986, w11987, w11988, w11989, w11990, w11991, w11992, w11993, w11994, w11995, w11996, w11997, w11998, w11999, w12000, w12001, w12002, w12003, w12004, w12005, w12006, w12007, w12008, w12009, w12010, w12011, w12012, w12013, w12014, w12015, w12016, w12017, w12018, w12019, w12020, w12021, w12022, w12023, w12024, w12025, w12026, w12027, w12028, w12029, w12030, w12031, w12032, w12033, w12034, w12035, w12036, w12037, w12038, w12039, w12040, w12041, w12042, w12043, w12044, w12045, w12046, w12047, w12048, w12049, w12050, w12051, w12052, w12053, w12054, w12055, w12056, w12057, w12058, w12059, w12060, w12061, w12062, w12063, w12064, w12065, w12066, w12067, w12068, w12069, w12070, w12071, w12072, w12073, w12074, w12075, w12076, w12077, w12078, w12079, w12080, w12081, w12082, w12083, w12084, w12085, w12086, w12087, w12088, w12089, w12090, w12091, w12092, w12093, w12094, w12095, w12096, w12097, w12098, w12099, w12100, w12101, w12102, w12103, w12104, w12105, w12106, w12107, w12108, w12109, w12110, w12111, w12112, w12113, w12114, w12115, w12116, w12117, w12118, w12119, w12120, w12121, w12122, w12123, w12124, w12125, w12126, w12127, w12128, w12129, w12130, w12131, w12132, w12133, w12134, w12135, w12136, w12137, w12138, w12139, w12140, w12141, w12142, w12143, w12144, w12145, w12146, w12147, w12148, w12149, w12150, w12151, w12152, w12153, w12154, w12155, w12156, w12157, w12158, w12159, w12160, w12161, w12162, w12163, w12164, w12165, w12166, w12167, w12168, w12169, w12170, w12171, w12172, w12173, w12174, w12175, w12176, w12177, w12178, w12179, w12180, w12181, w12182, w12183, w12184, w12185, w12186, w12187, w12188, w12189, w12190, w12191, w12192, w12193, w12194, w12195, w12196, w12197, w12198, w12199, w12200, w12201, w12202, w12203, w12204, w12205, w12206, w12207, w12208, w12209, w12210, w12211, w12212, w12213, w12214, w12215, w12216, w12217, w12218, w12219, w12220, w12221, w12222, w12223, w12224, w12225, w12226, w12227, w12228, w12229, w12230, w12231, w12232, w12233, w12234, w12235, w12236, w12237, w12238, w12239, w12240, w12241, w12242, w12243, w12244, w12245, w12246, w12247, w12248, w12249, w12250, w12251, w12252, w12253, w12254, w12255, w12256, w12257, w12258, w12259, w12260, w12261, w12262, w12263, w12264, w12265, w12266, w12267, w12268, w12269, w12270, w12271, w12272, w12273, w12274, w12275, w12276, w12277, w12278, w12279, w12280, w12281, w12282, w12283, w12284, w12285, w12286, w12287, w12288, w12289, w12290, w12291, w12292, w12293, w12294, w12295, w12296, w12297, w12298, w12299, w12300, w12301, w12302, w12303, w12304, w12305, w12306, w12307, w12308, w12309, w12310, w12311, w12312, w12313, w12314, w12315, w12316, w12317, w12318, w12319, w12320, w12321, w12322, w12323, w12324, w12325, w12326, w12327, w12328, w12329, w12330, w12331, w12332, w12333, w12334, w12335, w12336, w12337, w12338, w12339, w12340, w12341, w12342, w12343, w12344, w12345, w12346, w12347, w12348, w12349, w12350, w12351, w12352, w12353, w12354, w12355, w12356, w12357, w12358, w12359, w12360, w12361, w12362, w12363, w12364, w12365, w12366, w12367, w12368, w12369, w12370, w12371, w12372, w12373, w12374, w12375, w12376, w12377, w12378, w12379, w12380, w12381, w12382, w12383, w12384, w12385, w12386, w12387, w12388, w12389, w12390, w12391, w12392, w12393, w12394, w12395, w12396, w12397, w12398, w12399, w12400, w12401, w12402, w12403, w12404, w12405, w12406, w12407, w12408, w12409, w12410, w12411, w12412, w12413, w12414, w12415, w12416, w12417, w12418, w12419, w12420, w12421, w12422, w12423, w12424, w12425, w12426, w12427, w12428, w12429, w12430, w12431, w12432, w12433, w12434, w12435, w12436, w12437, w12438, w12439, w12440, w12441, w12442, w12443, w12444, w12445, w12446, w12447, w12448, w12449, w12450, w12451, w12452, w12453, w12454, w12455, w12456, w12457, w12458, w12459, w12460, w12461, w12462, w12463, w12464, w12465, w12466, w12467, w12468, w12469, w12470, w12471, w12472, w12473, w12474, w12475, w12476, w12477, w12478, w12479, w12480, w12481, w12482, w12483, w12484, w12485, w12486, w12487, w12488, w12489, w12490, w12491, w12492, w12493, w12494, w12495, w12496, w12497, w12498, w12499, w12500, w12501, w12502, w12503, w12504, w12505, w12506, w12507, w12508, w12509, w12510, w12511, w12512, w12513, w12514, w12515, w12516, w12517, w12518, w12519, w12520, w12521, w12522, w12523, w12524, w12525, w12526, w12527, w12528, w12529, w12530, w12531, w12532, w12533, w12534, w12535, w12536, w12537, w12538, w12539, w12540, w12541, w12542, w12543, w12544, w12545, w12546, w12547, w12548, w12549, w12550, w12551, w12552, w12553, w12554, w12555, w12556, w12557, w12558, w12559, w12560, w12561, w12562, w12563, w12564, w12565, w12566, w12567, w12568, w12569, w12570, w12571, w12572, w12573, w12574, w12575, w12576, w12577, w12578, w12579, w12580, w12581, w12582, w12583, w12584, w12585, w12586, w12587, w12588, w12589, w12590, w12591, w12592, w12593, w12594, w12595, w12596, w12597, w12598, w12599, w12600, w12601, w12602, w12603, w12604, w12605, w12606, w12607, w12608, w12609, w12610, w12611, w12612, w12613, w12614, w12615, w12616, w12617, w12618, w12619, w12620, w12621, w12622, w12623, w12624, w12625, w12626, w12627, w12628, w12629, w12630, w12631, w12632, w12633, w12634, w12635, w12636, w12637, w12638, w12639, w12640, w12641, w12642, w12643, w12644, w12645, w12646, w12647, w12648, w12649, w12650, w12651, w12652, w12653, w12654, w12655, w12656, w12657, w12658, w12659, w12660, w12661, w12662, w12663, w12664, w12665, w12666, w12667, w12668, w12669, w12670, w12671, w12672, w12673, w12674, w12675, w12676, w12677, w12678, w12679, w12680, w12681, w12682, w12683, w12684, w12685, w12686, w12687, w12688, w12689, w12690, w12691, w12692, w12693, w12694, w12695, w12696, w12697, w12698, w12699, w12700, w12701, w12702, w12703, w12704, w12705, w12706, w12707, w12708, w12709, w12710, w12711, w12712, w12713, w12714, w12715, w12716, w12717, w12718, w12719, w12720, w12721, w12722, w12723, w12724, w12725, w12726, w12727, w12728, w12729, w12730, w12731, w12732, w12733, w12734, w12735, w12736, w12737, w12738, w12739, w12740, w12741, w12742, w12743, w12744, w12745, w12746, w12747, w12748, w12749, w12750, w12751, w12752, w12753, w12754, w12755, w12756, w12757, w12758, w12759, w12760, w12761, w12762, w12763, w12764, w12765, w12766, w12767, w12768, w12769, w12770, w12771, w12772, w12773, w12774, w12775, w12776, w12777, w12778, w12779, w12780, w12781, w12782, w12783, w12784, w12785, w12786, w12787, w12788, w12789, w12790, w12791, w12792, w12793, w12794, w12795, w12796, w12797, w12798, w12799, w12800, w12801, w12802, w12803, w12804, w12805, w12806, w12807, w12808, w12809, w12810, w12811, w12812, w12813, w12814, w12815, w12816, w12817, w12818, w12819, w12820, w12821, w12822, w12823, w12824, w12825, w12826, w12827, w12828, w12829, w12830, w12831, w12832, w12833, w12834, w12835, w12836, w12837, w12838, w12839, w12840, w12841, w12842, w12843, w12844, w12845, w12846, w12847, w12848, w12849, w12850, w12851, w12852, w12853, w12854, w12855, w12856, w12857, w12858, w12859, w12860, w12861, w12862, w12863, w12864, w12865, w12866, w12867, w12868, w12869, w12870, w12871, w12872, w12873, w12874, w12875, w12876, w12877, w12878, w12879, w12880, w12881, w12882, w12883, w12884, w12885, w12886, w12887, w12888, w12889, w12890, w12891, w12892, w12893, w12894, w12895, w12896, w12897, w12898, w12899, w12900, w12901, w12902, w12903, w12904, w12905, w12906, w12907, w12908, w12909, w12910, w12911, w12912, w12913, w12914, w12915, w12916, w12917, w12918, w12919, w12920, w12921, w12922, w12923, w12924, w12925, w12926, w12927, w12928, w12929, w12930, w12931, w12932, w12933, w12934, w12935, w12936, w12937, w12938, w12939, w12940, w12941, w12942, w12943, w12944, w12945, w12946, w12947, w12948, w12949, w12950, w12951, w12952, w12953, w12954, w12955, w12956, w12957, w12958, w12959, w12960, w12961, w12962, w12963, w12964, w12965, w12966, w12967, w12968, w12969, w12970, w12971, w12972, w12973, w12974, w12975, w12976, w12977, w12978, w12979, w12980, w12981, w12982, w12983, w12984, w12985, w12986, w12987, w12988, w12989, w12990, w12991, w12992, w12993, w12994, w12995, w12996, w12997, w12998, w12999, w13000, w13001, w13002, w13003, w13004, w13005, w13006, w13007, w13008, w13009, w13010, w13011, w13012, w13013, w13014, w13015, w13016, w13017, w13018, w13019, w13020, w13021, w13022, w13023, w13024, w13025, w13026, w13027, w13028, w13029, w13030, w13031, w13032, w13033, w13034, w13035, w13036, w13037, w13038, w13039, w13040, w13041, w13042, w13043, w13044, w13045, w13046, w13047, w13048, w13049, w13050, w13051, w13052, w13053, w13054, w13055, w13056, w13057, w13058, w13059, w13060, w13061, w13062, w13063, w13064, w13065, w13066, w13067, w13068, w13069, w13070, w13071, w13072, w13073, w13074, w13075, w13076, w13077, w13078, w13079, w13080, w13081, w13082, w13083, w13084, w13085, w13086, w13087, w13088, w13089, w13090, w13091, w13092, w13093, w13094, w13095, w13096, w13097, w13098, w13099, w13100, w13101, w13102, w13103, w13104, w13105, w13106, w13107, w13108, w13109, w13110, w13111, w13112, w13113, w13114, w13115, w13116, w13117, w13118, w13119, w13120, w13121, w13122, w13123, w13124, w13125, w13126, w13127, w13128, w13129, w13130, w13131, w13132, w13133, w13134, w13135, w13136, w13137, w13138, w13139, w13140, w13141, w13142, w13143, w13144, w13145, w13146, w13147, w13148, w13149, w13150, w13151, w13152, w13153, w13154, w13155, w13156, w13157, w13158, w13159, w13160, w13161, w13162, w13163, w13164, w13165, w13166, w13167, w13168, w13169, w13170, w13171, w13172, w13173, w13174, w13175, w13176, w13177, w13178, w13179, w13180, w13181, w13182, w13183, w13184, w13185, w13186, w13187, w13188, w13189, w13190, w13191, w13192, w13193, w13194, w13195, w13196, w13197, w13198, w13199, w13200, w13201, w13202, w13203, w13204, w13205, w13206, w13207, w13208, w13209, w13210, w13211, w13212, w13213, w13214, w13215, w13216, w13217, w13218, w13219, w13220, w13221, w13222, w13223, w13224, w13225, w13226, w13227, w13228, w13229, w13230, w13231, w13232, w13233, w13234, w13235, w13236, w13237, w13238, w13239, w13240, w13241, w13242, w13243, w13244, w13245, w13246, w13247, w13248, w13249, w13250, w13251, w13252, w13253, w13254, w13255, w13256, w13257, w13258, w13259, w13260, w13261, w13262, w13263, w13264, w13265, w13266, w13267, w13268, w13269, w13270, w13271, w13272, w13273, w13274, w13275, w13276, w13277, w13278, w13279, w13280, w13281, w13282, w13283, w13284, w13285, w13286, w13287, w13288, w13289, w13290, w13291, w13292, w13293, w13294, w13295, w13296, w13297, w13298, w13299, w13300, w13301, w13302, w13303, w13304, w13305, w13306, w13307, w13308, w13309, w13310, w13311, w13312, w13313, w13314, w13315, w13316, w13317, w13318, w13319, w13320, w13321, w13322, w13323, w13324, w13325, w13326, w13327, w13328, w13329, w13330, w13331, w13332, w13333, w13334, w13335, w13336, w13337, w13338, w13339, w13340, w13341, w13342, w13343, w13344, w13345, w13346, w13347, w13348, w13349, w13350, w13351, w13352, w13353, w13354, w13355, w13356, w13357, w13358, w13359, w13360, w13361, w13362, w13363, w13364, w13365, w13366, w13367, w13368, w13369, w13370, w13371, w13372, w13373, w13374, w13375, w13376, w13377, w13378, w13379, w13380, w13381, w13382, w13383, w13384, w13385, w13386, w13387, w13388, w13389, w13390, w13391, w13392, w13393, w13394, w13395, w13396, w13397, w13398, w13399, w13400, w13401, w13402, w13403, w13404, w13405, w13406, w13407, w13408, w13409, w13410, w13411, w13412, w13413, w13414, w13415, w13416, w13417, w13418, w13419, w13420, w13421, w13422, w13423, w13424, w13425, w13426, w13427, w13428, w13429, w13430, w13431, w13432, w13433, w13434, w13435, w13436, w13437, w13438, w13439, w13440, w13441, w13442, w13443, w13444, w13445, w13446, w13447, w13448, w13449, w13450, w13451, w13452, w13453, w13454, w13455, w13456, w13457, w13458, w13459, w13460, w13461, w13462, w13463, w13464, w13465, w13466, w13467, w13468, w13469, w13470, w13471, w13472, w13473, w13474, w13475, w13476, w13477, w13478, w13479, w13480, w13481, w13482, w13483, w13484, w13485, w13486, w13487, w13488, w13489, w13490, w13491, w13492, w13493, w13494, w13495, w13496, w13497, w13498, w13499, w13500, w13501, w13502, w13503, w13504, w13505, w13506, w13507, w13508, w13509, w13510, w13511, w13512, w13513, w13514, w13515, w13516, w13517, w13518, w13519, w13520, w13521, w13522, w13523, w13524, w13525, w13526, w13527, w13528, w13529, w13530, w13531, w13532, w13533, w13534, w13535, w13536, w13537, w13538, w13539, w13540, w13541, w13542, w13543, w13544, w13545, w13546, w13547, w13548, w13549, w13550, w13551, w13552, w13553, w13554, w13555, w13556, w13557, w13558, w13559, w13560, w13561, w13562, w13563, w13564, w13565, w13566, w13567, w13568, w13569, w13570, w13571, w13572, w13573, w13574, w13575, w13576, w13577, w13578, w13579, w13580, w13581, w13582, w13583, w13584, w13585, w13586, w13587, w13588, w13589, w13590, w13591, w13592, w13593, w13594, w13595, w13596, w13597, w13598, w13599, w13600, w13601, w13602, w13603, w13604, w13605, w13606, w13607, w13608, w13609, w13610, w13611, w13612, w13613, w13614, w13615, w13616, w13617, w13618, w13619, w13620, w13621, w13622, w13623, w13624, w13625, w13626, w13627, w13628, w13629, w13630, w13631, w13632, w13633, w13634, w13635, w13636, w13637, w13638, w13639, w13640, w13641, w13642, w13643, w13644, w13645, w13646, w13647, w13648, w13649, w13650, w13651, w13652, w13653, w13654, w13655, w13656, w13657, w13658, w13659, w13660, w13661, w13662, w13663, w13664, w13665, w13666, w13667, w13668, w13669, w13670, w13671, w13672, w13673, w13674, w13675, w13676, w13677, w13678, w13679, w13680, w13681, w13682, w13683, w13684, w13685, w13686, w13687, w13688, w13689, w13690, w13691, w13692, w13693, w13694, w13695, w13696, w13697, w13698, w13699, w13700, w13701, w13702, w13703, w13704, w13705, w13706, w13707, w13708, w13709, w13710, w13711, w13712, w13713, w13714, w13715, w13716, w13717, w13718, w13719, w13720, w13721, w13722, w13723, w13724, w13725, w13726, w13727, w13728, w13729, w13730, w13731, w13732, w13733, w13734, w13735, w13736, w13737, w13738, w13739, w13740, w13741, w13742, w13743, w13744, w13745, w13746, w13747, w13748, w13749, w13750, w13751, w13752, w13753, w13754, w13755, w13756, w13757, w13758, w13759, w13760, w13761, w13762, w13763, w13764, w13765, w13766, w13767, w13768, w13769, w13770, w13771, w13772, w13773, w13774, w13775, w13776, w13777, w13778, w13779, w13780, w13781, w13782, w13783, w13784, w13785, w13786, w13787, w13788, w13789, w13790, w13791, w13792, w13793, w13794, w13795, w13796, w13797, w13798, w13799, w13800, w13801, w13802, w13803, w13804, w13805, w13806, w13807, w13808, w13809, w13810, w13811, w13812, w13813, w13814, w13815, w13816, w13817, w13818, w13819, w13820, w13821, w13822, w13823, w13824, w13825, w13826, w13827, w13828, w13829, w13830, w13831, w13832, w13833, w13834, w13835, w13836, w13837, w13838, w13839, w13840, w13841, w13842, w13843, w13844, w13845, w13846, w13847, w13848, w13849, w13850, w13851, w13852, w13853, w13854, w13855, w13856, w13857, w13858, w13859, w13860, w13861, w13862, w13863, w13864, w13865, w13866, w13867, w13868, w13869, w13870, w13871, w13872, w13873, w13874, w13875, w13876, w13877, w13878, w13879, w13880, w13881, w13882, w13883, w13884, w13885, w13886, w13887, w13888, w13889, w13890, w13891, w13892, w13893, w13894, w13895, w13896, w13897, w13898, w13899, w13900, w13901, w13902, w13903, w13904, w13905, w13906, w13907, w13908, w13909, w13910, w13911, w13912, w13913, w13914, w13915, w13916, w13917, w13918, w13919, w13920, w13921, w13922, w13923, w13924, w13925, w13926, w13927, w13928, w13929, w13930, w13931, w13932, w13933, w13934, w13935, w13936, w13937, w13938, w13939, w13940, w13941, w13942, w13943, w13944, w13945, w13946, w13947, w13948, w13949, w13950, w13951, w13952, w13953, w13954, w13955, w13956, w13957, w13958, w13959, w13960, w13961, w13962, w13963, w13964, w13965, w13966, w13967, w13968, w13969, w13970, w13971, w13972, w13973, w13974, w13975, w13976, w13977, w13978, w13979, w13980, w13981, w13982, w13983, w13984, w13985, w13986, w13987, w13988, w13989, w13990, w13991, w13992, w13993, w13994, w13995, w13996, w13997, w13998, w13999, w14000, w14001, w14002, w14003, w14004, w14005, w14006, w14007, w14008, w14009, w14010, w14011, w14012, w14013, w14014, w14015, w14016, w14017, w14018, w14019, w14020, w14021, w14022, w14023, w14024, w14025, w14026, w14027, w14028, w14029, w14030, w14031, w14032, w14033, w14034, w14035, w14036, w14037, w14038, w14039, w14040, w14041, w14042, w14043, w14044, w14045, w14046, w14047, w14048, w14049, w14050, w14051, w14052, w14053, w14054, w14055, w14056, w14057, w14058, w14059, w14060, w14061, w14062, w14063, w14064, w14065, w14066, w14067, w14068, w14069, w14070, w14071, w14072, w14073, w14074, w14075, w14076, w14077, w14078, w14079, w14080, w14081, w14082, w14083, w14084, w14085, w14086, w14087, w14088, w14089, w14090, w14091, w14092, w14093, w14094, w14095, w14096, w14097, w14098, w14099, w14100, w14101, w14102, w14103, w14104, w14105, w14106, w14107, w14108, w14109, w14110, w14111, w14112, w14113, w14114, w14115, w14116, w14117, w14118, w14119, w14120, w14121, w14122, w14123, w14124, w14125, w14126, w14127, w14128, w14129, w14130, w14131, w14132, w14133, w14134, w14135, w14136, w14137, w14138, w14139, w14140, w14141, w14142, w14143, w14144, w14145, w14146, w14147, w14148, w14149, w14150, w14151, w14152, w14153, w14154, w14155, w14156, w14157, w14158, w14159, w14160, w14161, w14162, w14163, w14164, w14165, w14166, w14167, w14168, w14169, w14170, w14171, w14172, w14173, w14174, w14175, w14176, w14177, w14178, w14179, w14180, w14181, w14182, w14183, w14184, w14185, w14186, w14187, w14188, w14189, w14190, w14191, w14192, w14193, w14194, w14195, w14196, w14197, w14198, w14199, w14200, w14201, w14202, w14203, w14204, w14205, w14206, w14207, w14208, w14209, w14210, w14211, w14212, w14213, w14214, w14215, w14216, w14217, w14218, w14219, w14220, w14221, w14222, w14223, w14224, w14225, w14226, w14227, w14228, w14229, w14230, w14231, w14232, w14233, w14234, w14235, w14236, w14237, w14238, w14239, w14240, w14241, w14242, w14243, w14244, w14245, w14246, w14247, w14248, w14249, w14250, w14251, w14252, w14253, w14254, w14255, w14256, w14257, w14258, w14259, w14260, w14261, w14262, w14263, w14264, w14265, w14266, w14267, w14268, w14269, w14270, w14271, w14272, w14273, w14274, w14275, w14276, w14277, w14278, w14279, w14280, w14281, w14282, w14283, w14284, w14285, w14286, w14287, w14288, w14289, w14290, w14291, w14292, w14293, w14294, w14295, w14296, w14297, w14298, w14299, w14300, w14301, w14302, w14303, w14304, w14305, w14306, w14307, w14308, w14309, w14310, w14311, w14312, w14313, w14314, w14315, w14316, w14317, w14318, w14319, w14320, w14321, w14322, w14323, w14324, w14325, w14326, w14327, w14328, w14329, w14330, w14331, w14332, w14333, w14334, w14335, w14336, w14337, w14338, w14339, w14340, w14341, w14342, w14343, w14344, w14345, w14346, w14347, w14348, w14349, w14350, w14351, w14352, w14353, w14354, w14355, w14356, w14357, w14358, w14359, w14360, w14361, w14362, w14363, w14364, w14365, w14366, w14367, w14368, w14369, w14370, w14371, w14372, w14373, w14374, w14375, w14376, w14377, w14378, w14379, w14380, w14381, w14382, w14383, w14384, w14385, w14386, w14387, w14388, w14389, w14390, w14391, w14392, w14393, w14394, w14395, w14396, w14397, w14398, w14399, w14400, w14401, w14402, w14403, w14404, w14405, w14406, w14407, w14408, w14409, w14410, w14411, w14412, w14413, w14414, w14415, w14416, w14417, w14418, w14419, w14420, w14421, w14422, w14423, w14424, w14425, w14426, w14427, w14428, w14429, w14430, w14431, w14432, w14433, w14434, w14435, w14436, w14437, w14438, w14439, w14440, w14441, w14442, w14443, w14444, w14445, w14446, w14447, w14448, w14449, w14450, w14451, w14452, w14453, w14454, w14455, w14456, w14457, w14458, w14459, w14460, w14461, w14462, w14463, w14464, w14465, w14466, w14467, w14468, w14469, w14470, w14471, w14472, w14473, w14474, w14475, w14476, w14477, w14478, w14479, w14480, w14481, w14482, w14483, w14484, w14485, w14486, w14487, w14488, w14489, w14490, w14491, w14492, w14493, w14494, w14495, w14496, w14497, w14498, w14499, w14500, w14501, w14502, w14503, w14504, w14505, w14506, w14507, w14508, w14509, w14510, w14511, w14512, w14513, w14514, w14515, w14516, w14517, w14518, w14519, w14520, w14521, w14522, w14523, w14524, w14525, w14526, w14527, w14528, w14529, w14530, w14531, w14532, w14533, w14534, w14535, w14536, w14537, w14538, w14539, w14540, w14541, w14542, w14543, w14544, w14545, w14546, w14547, w14548, w14549, w14550, w14551, w14552, w14553, w14554, w14555, w14556, w14557, w14558, w14559, w14560, w14561, w14562, w14563, w14564, w14565, w14566, w14567, w14568, w14569, w14570, w14571, w14572, w14573, w14574, w14575, w14576, w14577, w14578, w14579, w14580, w14581, w14582, w14583, w14584, w14585, w14586, w14587, w14588, w14589, w14590, w14591, w14592, w14593, w14594, w14595, w14596, w14597, w14598, w14599, w14600, w14601, w14602, w14603, w14604, w14605, w14606, w14607, w14608, w14609, w14610, w14611, w14612, w14613, w14614, w14615, w14616, w14617, w14618, w14619, w14620, w14621, w14622, w14623, w14624, w14625, w14626, w14627, w14628, w14629, w14630, w14631, w14632, w14633, w14634, w14635, w14636, w14637, w14638, w14639, w14640, w14641, w14642, w14643, w14644, w14645, w14646, w14647, w14648, w14649, w14650, w14651, w14652, w14653, w14654, w14655, w14656, w14657, w14658, w14659, w14660, w14661, w14662, w14663, w14664, w14665, w14666, w14667, w14668, w14669, w14670, w14671, w14672, w14673, w14674, w14675, w14676, w14677, w14678, w14679, w14680, w14681, w14682, w14683, w14684, w14685, w14686, w14687, w14688, w14689, w14690, w14691, w14692, w14693, w14694, w14695, w14696, w14697, w14698, w14699, w14700, w14701, w14702, w14703, w14704, w14705, w14706, w14707, w14708, w14709, w14710, w14711, w14712, w14713, w14714, w14715, w14716, w14717, w14718, w14719, w14720, w14721, w14722, w14723, w14724, w14725, w14726, w14727, w14728, w14729, w14730, w14731, w14732, w14733, w14734, w14735, w14736, w14737, w14738, w14739, w14740, w14741, w14742, w14743, w14744, w14745, w14746, w14747, w14748, w14749, w14750, w14751, w14752, w14753, w14754, w14755, w14756, w14757, w14758, w14759, w14760, w14761, w14762, w14763, w14764, w14765, w14766, w14767, w14768, w14769, w14770, w14771, w14772, w14773, w14774, w14775, w14776, w14777, w14778, w14779, w14780, w14781, w14782, w14783, w14784, w14785, w14786, w14787, w14788, w14789, w14790, w14791, w14792, w14793, w14794, w14795, w14796, w14797, w14798, w14799, w14800, w14801, w14802, w14803, w14804, w14805, w14806, w14807, w14808, w14809, w14810, w14811, w14812, w14813, w14814, w14815, w14816, w14817, w14818, w14819, w14820, w14821, w14822, w14823, w14824, w14825, w14826, w14827, w14828, w14829, w14830, w14831, w14832, w14833, w14834, w14835, w14836, w14837, w14838, w14839, w14840, w14841, w14842, w14843, w14844, w14845, w14846, w14847, w14848, w14849, w14850, w14851, w14852, w14853, w14854, w14855, w14856, w14857, w14858, w14859, w14860, w14861, w14862, w14863, w14864, w14865, w14866, w14867, w14868, w14869, w14870, w14871, w14872, w14873, w14874, w14875, w14876, w14877, w14878, w14879, w14880, w14881, w14882, w14883, w14884, w14885, w14886, w14887, w14888, w14889, w14890, w14891, w14892, w14893, w14894, w14895, w14896, w14897, w14898, w14899, w14900, w14901, w14902, w14903, w14904, w14905, w14906, w14907, w14908, w14909, w14910, w14911, w14912, w14913, w14914, w14915, w14916, w14917, w14918, w14919, w14920, w14921, w14922, w14923, w14924, w14925, w14926, w14927, w14928, w14929, w14930, w14931, w14932, w14933, w14934, w14935, w14936, w14937, w14938, w14939, w14940, w14941, w14942, w14943, w14944, w14945, w14946, w14947, w14948, w14949, w14950, w14951, w14952, w14953, w14954, w14955, w14956, w14957, w14958, w14959, w14960, w14961, w14962, w14963, w14964, w14965, w14966, w14967, w14968, w14969, w14970, w14971, w14972, w14973, w14974, w14975, w14976, w14977, w14978, w14979, w14980, w14981, w14982, w14983, w14984, w14985, w14986, w14987, w14988, w14989, w14990, w14991, w14992, w14993, w14994, w14995, w14996, w14997, w14998, w14999, w15000, w15001, w15002, w15003, w15004, w15005, w15006, w15007, w15008, w15009, w15010, w15011, w15012, w15013, w15014, w15015, w15016, w15017, w15018, w15019, w15020, w15021, w15022, w15023, w15024, w15025, w15026, w15027, w15028, w15029, w15030, w15031, w15032, w15033, w15034, w15035, w15036, w15037, w15038, w15039, w15040, w15041, w15042, w15043, w15044, w15045, w15046, w15047, w15048, w15049, w15050, w15051, w15052, w15053, w15054, w15055, w15056, w15057, w15058, w15059, w15060, w15061, w15062, w15063, w15064, w15065, w15066, w15067, w15068, w15069, w15070, w15071, w15072, w15073, w15074, w15075, w15076, w15077, w15078, w15079, w15080, w15081, w15082, w15083, w15084, w15085, w15086, w15087, w15088, w15089, w15090, w15091, w15092, w15093, w15094, w15095, w15096, w15097, w15098, w15099, w15100, w15101, w15102, w15103, w15104, w15105, w15106, w15107, w15108, w15109, w15110, w15111, w15112, w15113, w15114, w15115, w15116, w15117, w15118, w15119, w15120, w15121, w15122, w15123, w15124, w15125, w15126, w15127, w15128, w15129, w15130, w15131, w15132, w15133, w15134, w15135, w15136, w15137, w15138, w15139, w15140, w15141, w15142, w15143, w15144, w15145, w15146, w15147, w15148, w15149, w15150, w15151, w15152, w15153, w15154, w15155, w15156, w15157, w15158, w15159, w15160, w15161, w15162, w15163, w15164, w15165, w15166, w15167, w15168, w15169, w15170, w15171, w15172, w15173, w15174, w15175, w15176, w15177, w15178, w15179, w15180, w15181, w15182, w15183, w15184, w15185, w15186, w15187, w15188, w15189, w15190, w15191, w15192, w15193, w15194, w15195, w15196, w15197, w15198, w15199, w15200, w15201, w15202, w15203, w15204, w15205, w15206, w15207, w15208, w15209, w15210, w15211, w15212, w15213, w15214, w15215, w15216, w15217, w15218, w15219, w15220, w15221, w15222, w15223, w15224, w15225, w15226, w15227, w15228, w15229, w15230, w15231, w15232, w15233, w15234, w15235, w15236, w15237, w15238, w15239, w15240, w15241, w15242, w15243, w15244, w15245, w15246, w15247, w15248, w15249, w15250, w15251, w15252, w15253, w15254, w15255, w15256, w15257, w15258, w15259, w15260, w15261, w15262, w15263, w15264, w15265, w15266, w15267, w15268, w15269, w15270, w15271, w15272, w15273, w15274, w15275, w15276, w15277, w15278, w15279, w15280, w15281, w15282, w15283, w15284, w15285, w15286, w15287, w15288, w15289, w15290, w15291, w15292, w15293, w15294, w15295, w15296, w15297, w15298, w15299, w15300, w15301, w15302, w15303, w15304, w15305, w15306, w15307, w15308, w15309, w15310, w15311, w15312, w15313, w15314, w15315, w15316, w15317, w15318, w15319, w15320, w15321, w15322, w15323, w15324, w15325, w15326, w15327, w15328, w15329, w15330, w15331, w15332, w15333, w15334, w15335, w15336, w15337, w15338, w15339, w15340, w15341, w15342, w15343, w15344, w15345, w15346, w15347, w15348, w15349, w15350, w15351, w15352, w15353, w15354, w15355, w15356, w15357, w15358, w15359, w15360, w15361, w15362, w15363, w15364, w15365, w15366, w15367, w15368, w15369, w15370, w15371, w15372, w15373, w15374, w15375, w15376, w15377, w15378, w15379, w15380, w15381, w15382, w15383, w15384, w15385, w15386, w15387, w15388, w15389, w15390, w15391, w15392, w15393, w15394, w15395, w15396, w15397, w15398, w15399, w15400, w15401, w15402, w15403, w15404, w15405, w15406, w15407, w15408, w15409, w15410, w15411, w15412, w15413, w15414, w15415, w15416, w15417, w15418, w15419, w15420, w15421, w15422, w15423, w15424, w15425, w15426, w15427, w15428, w15429, w15430, w15431, w15432, w15433, w15434, w15435, w15436, w15437, w15438, w15439, w15440, w15441, w15442, w15443, w15444, w15445, w15446, w15447, w15448, w15449, w15450, w15451, w15452, w15453, w15454, w15455, w15456, w15457, w15458, w15459, w15460, w15461, w15462, w15463, w15464, w15465, w15466, w15467, w15468, w15469, w15470, w15471, w15472, w15473, w15474, w15475, w15476, w15477, w15478, w15479, w15480, w15481, w15482, w15483, w15484, w15485, w15486, w15487, w15488, w15489, w15490, w15491, w15492, w15493, w15494, w15495, w15496, w15497, w15498, w15499, w15500, w15501, w15502, w15503, w15504, w15505, w15506, w15507, w15508, w15509, w15510, w15511, w15512, w15513, w15514, w15515, w15516, w15517, w15518, w15519, w15520, w15521, w15522, w15523, w15524, w15525, w15526, w15527, w15528, w15529, w15530, w15531, w15532, w15533, w15534, w15535, w15536, w15537, w15538, w15539, w15540, w15541, w15542, w15543, w15544, w15545, w15546, w15547, w15548, w15549, w15550, w15551, w15552, w15553, w15554, w15555, w15556, w15557, w15558, w15559, w15560, w15561, w15562, w15563, w15564, w15565, w15566, w15567, w15568, w15569, w15570, w15571, w15572, w15573, w15574, w15575, w15576, w15577, w15578, w15579, w15580, w15581, w15582, w15583, w15584, w15585, w15586, w15587, w15588, w15589, w15590, w15591, w15592, w15593, w15594, w15595, w15596, w15597, w15598, w15599, w15600, w15601, w15602, w15603, w15604, w15605, w15606, w15607, w15608, w15609, w15610, w15611, w15612, w15613, w15614, w15615, w15616, w15617, w15618, w15619, w15620, w15621, w15622, w15623, w15624, w15625, w15626, w15627, w15628, w15629, w15630, w15631, w15632, w15633, w15634, w15635, w15636, w15637, w15638, w15639, w15640, w15641, w15642, w15643, w15644, w15645, w15646, w15647, w15648, w15649, w15650, w15651, w15652, w15653, w15654, w15655, w15656, w15657, w15658, w15659, w15660, w15661, w15662, w15663, w15664, w15665, w15666, w15667, w15668, w15669, w15670, w15671, w15672, w15673, w15674, w15675, w15676, w15677, w15678, w15679, w15680, w15681, w15682, w15683, w15684, w15685, w15686, w15687, w15688, w15689, w15690, w15691, w15692, w15693, w15694, w15695, w15696, w15697, w15698, w15699, w15700, w15701, w15702, w15703, w15704, w15705, w15706, w15707, w15708, w15709, w15710, w15711, w15712, w15713, w15714, w15715, w15716, w15717, w15718, w15719, w15720, w15721, w15722, w15723, w15724, w15725, w15726, w15727, w15728, w15729, w15730, w15731, w15732, w15733, w15734, w15735, w15736, w15737, w15738, w15739, w15740, w15741, w15742, w15743, w15744, w15745, w15746, w15747, w15748, w15749, w15750, w15751, w15752, w15753, w15754, w15755, w15756, w15757, w15758, w15759, w15760, w15761, w15762, w15763, w15764, w15765, w15766, w15767, w15768, w15769, w15770, w15771, w15772, w15773, w15774, w15775, w15776, w15777, w15778, w15779, w15780, w15781, w15782, w15783, w15784, w15785, w15786, w15787, w15788, w15789, w15790, w15791, w15792, w15793, w15794, w15795, w15796, w15797, w15798, w15799, w15800, w15801, w15802, w15803, w15804, w15805, w15806, w15807, w15808, w15809, w15810, w15811, w15812, w15813, w15814, w15815, w15816, w15817, w15818, w15819, w15820, w15821, w15822, w15823, w15824, w15825, w15826, w15827, w15828, w15829, w15830, w15831, w15832, w15833, w15834, w15835, w15836, w15837, w15838, w15839, w15840, w15841, w15842, w15843, w15844, w15845, w15846, w15847, w15848, w15849, w15850, w15851, w15852, w15853, w15854, w15855, w15856, w15857, w15858, w15859, w15860, w15861, w15862, w15863, w15864, w15865, w15866, w15867, w15868, w15869, w15870, w15871, w15872, w15873, w15874, w15875, w15876, w15877, w15878, w15879, w15880, w15881, w15882, w15883, w15884, w15885, w15886, w15887, w15888, w15889, w15890, w15891, w15892, w15893, w15894, w15895, w15896, w15897, w15898, w15899, w15900, w15901, w15902, w15903, w15904, w15905, w15906, w15907, w15908, w15909, w15910, w15911, w15912, w15913, w15914, w15915, w15916, w15917, w15918, w15919, w15920, w15921, w15922, w15923, w15924, w15925, w15926, w15927, w15928, w15929, w15930, w15931, w15932, w15933, w15934, w15935, w15936, w15937, w15938, w15939, w15940, w15941, w15942, w15943, w15944, w15945, w15946, w15947, w15948, w15949, w15950, w15951, w15952, w15953, w15954, w15955, w15956, w15957, w15958, w15959, w15960, w15961, w15962, w15963, w15964, w15965, w15966, w15967, w15968, w15969, w15970, w15971, w15972, w15973, w15974, w15975, w15976, w15977, w15978, w15979, w15980, w15981, w15982, w15983, w15984, w15985, w15986, w15987, w15988, w15989, w15990, w15991, w15992, w15993, w15994, w15995, w15996, w15997, w15998, w15999, w16000, w16001, w16002, w16003, w16004, w16005, w16006, w16007, w16008, w16009, w16010, w16011, w16012, w16013, w16014, w16015, w16016, w16017, w16018, w16019, w16020, w16021, w16022, w16023, w16024, w16025, w16026, w16027, w16028, w16029, w16030, w16031, w16032, w16033, w16034, w16035, w16036, w16037, w16038, w16039, w16040, w16041, w16042, w16043, w16044, w16045, w16046, w16047, w16048, w16049, w16050, w16051, w16052, w16053, w16054, w16055, w16056, w16057, w16058, w16059, w16060, w16061, w16062, w16063, w16064, w16065, w16066, w16067, w16068, w16069, w16070, w16071, w16072, w16073, w16074, w16075, w16076, w16077, w16078, w16079, w16080, w16081, w16082, w16083, w16084, w16085, w16086, w16087, w16088, w16089, w16090, w16091, w16092, w16093, w16094, w16095, w16096, w16097, w16098, w16099, w16100, w16101, w16102, w16103, w16104, w16105, w16106, w16107, w16108, w16109, w16110, w16111, w16112, w16113, w16114, w16115, w16116, w16117, w16118, w16119, w16120, w16121, w16122, w16123, w16124, w16125, w16126, w16127, w16128, w16129, w16130, w16131, w16132, w16133, w16134, w16135, w16136, w16137, w16138, w16139, w16140, w16141, w16142, w16143, w16144, w16145, w16146, w16147, w16148, w16149, w16150, w16151, w16152, w16153, w16154, w16155, w16156, w16157, w16158, w16159, w16160, w16161, w16162, w16163, w16164, w16165, w16166, w16167, w16168, w16169, w16170, w16171, w16172, w16173, w16174, w16175, w16176, w16177, w16178, w16179, w16180, w16181, w16182, w16183, w16184, w16185, w16186, w16187, w16188, w16189, w16190, w16191, w16192, w16193, w16194, w16195, w16196, w16197, w16198, w16199, w16200, w16201, w16202, w16203, w16204, w16205, w16206, w16207, w16208, w16209, w16210, w16211, w16212, w16213, w16214, w16215, w16216, w16217, w16218, w16219, w16220, w16221, w16222, w16223, w16224, w16225, w16226, w16227, w16228, w16229, w16230, w16231, w16232, w16233, w16234, w16235, w16236, w16237, w16238, w16239, w16240, w16241, w16242, w16243, w16244, w16245, w16246, w16247, w16248, w16249, w16250, w16251, w16252, w16253, w16254, w16255, w16256, w16257, w16258, w16259, w16260, w16261, w16262, w16263, w16264, w16265, w16266, w16267, w16268, w16269, w16270, w16271, w16272, w16273, w16274, w16275, w16276, w16277, w16278, w16279, w16280, w16281, w16282, w16283, w16284, w16285, w16286, w16287, w16288, w16289, w16290, w16291, w16292, w16293, w16294, w16295, w16296, w16297, w16298, w16299, w16300, w16301, w16302, w16303, w16304, w16305, w16306, w16307, w16308, w16309, w16310, w16311, w16312, w16313, w16314, w16315, w16316, w16317, w16318, w16319, w16320, w16321, w16322, w16323, w16324, w16325, w16326, w16327, w16328, w16329, w16330, w16331, w16332, w16333, w16334, w16335, w16336, w16337, w16338, w16339, w16340, w16341, w16342, w16343, w16344, w16345, w16346, w16347, w16348, w16349, w16350, w16351, w16352, w16353, w16354, w16355, w16356, w16357, w16358, w16359, w16360, w16361, w16362, w16363, w16364, w16365, w16366, w16367, w16368, w16369, w16370, w16371, w16372, w16373, w16374, w16375, w16376, w16377, w16378, w16379, w16380, w16381, w16382, w16383, w16384, w16385, w16386, w16387, w16388, w16389, w16390, w16391, w16392, w16393, w16394, w16395, w16396, w16397, w16398, w16399, w16400, w16401, w16402, w16403, w16404, w16405, w16406, w16407, w16408, w16409, w16410, w16411, w16412, w16413, w16414, w16415, w16416, w16417, w16418, w16419, w16420, w16421, w16422, w16423, w16424, w16425, w16426, w16427, w16428, w16429, w16430, w16431, w16432, w16433, w16434, w16435, w16436, w16437, w16438, w16439, w16440, w16441, w16442, w16443, w16444, w16445, w16446, w16447, w16448, w16449, w16450, w16451, w16452, w16453, w16454, w16455, w16456, w16457, w16458, w16459, w16460, w16461, w16462, w16463, w16464, w16465, w16466, w16467, w16468, w16469, w16470, w16471, w16472, w16473, w16474, w16475, w16476, w16477, w16478, w16479, w16480, w16481, w16482, w16483, w16484, w16485, w16486, w16487, w16488, w16489, w16490, w16491, w16492, w16493, w16494, w16495, w16496, w16497, w16498, w16499, w16500, w16501, w16502, w16503, w16504, w16505, w16506, w16507, w16508, w16509, w16510, w16511, w16512, w16513, w16514, w16515, w16516, w16517, w16518, w16519, w16520, w16521, w16522, w16523, w16524, w16525, w16526, w16527, w16528, w16529, w16530, w16531, w16532, w16533, w16534, w16535, w16536, w16537, w16538, w16539, w16540, w16541, w16542, w16543, w16544, w16545, w16546, w16547, w16548, w16549, w16550, w16551, w16552, w16553, w16554, w16555, w16556, w16557, w16558, w16559, w16560, w16561, w16562, w16563, w16564, w16565, w16566, w16567, w16568, w16569, w16570, w16571, w16572, w16573, w16574, w16575, w16576, w16577, w16578, w16579, w16580, w16581, w16582, w16583, w16584, w16585, w16586, w16587, w16588, w16589, w16590, w16591, w16592, w16593, w16594, w16595, w16596, w16597, w16598, w16599, w16600, w16601, w16602, w16603, w16604, w16605, w16606, w16607, w16608, w16609, w16610, w16611, w16612, w16613, w16614, w16615, w16616, w16617, w16618, w16619, w16620, w16621, w16622, w16623, w16624, w16625, w16626, w16627, w16628, w16629, w16630, w16631, w16632, w16633, w16634, w16635, w16636, w16637, w16638, w16639, w16640, w16641, w16642, w16643, w16644, w16645, w16646, w16647, w16648, w16649, w16650, w16651, w16652, w16653, w16654, w16655, w16656, w16657, w16658, w16659, w16660, w16661, w16662, w16663, w16664, w16665, w16666, w16667, w16668, w16669, w16670, w16671, w16672, w16673, w16674, w16675, w16676, w16677, w16678, w16679, w16680, w16681, w16682, w16683, w16684, w16685, w16686, w16687, w16688, w16689, w16690, w16691, w16692, w16693, w16694, w16695, w16696, w16697, w16698, w16699, w16700, w16701, w16702, w16703, w16704, w16705, w16706, w16707, w16708, w16709, w16710, w16711, w16712, w16713, w16714, w16715, w16716, w16717, w16718, w16719, w16720, w16721, w16722, w16723, w16724, w16725, w16726, w16727, w16728, w16729, w16730, w16731, w16732, w16733, w16734, w16735, w16736, w16737, w16738, w16739, w16740, w16741, w16742, w16743, w16744, w16745, w16746, w16747, w16748, w16749, w16750, w16751, w16752, w16753, w16754, w16755, w16756, w16757, w16758, w16759, w16760, w16761, w16762, w16763, w16764, w16765, w16766, w16767, w16768, w16769, w16770, w16771, w16772, w16773, w16774, w16775, w16776, w16777, w16778, w16779, w16780, w16781, w16782, w16783, w16784, w16785, w16786, w16787, w16788, w16789, w16790, w16791, w16792, w16793, w16794, w16795, w16796, w16797, w16798, w16799, w16800, w16801, w16802, w16803, w16804, w16805, w16806, w16807, w16808, w16809, w16810, w16811, w16812, w16813, w16814, w16815, w16816, w16817, w16818, w16819, w16820, w16821, w16822, w16823, w16824, w16825, w16826, w16827, w16828, w16829, w16830, w16831, w16832, w16833, w16834, w16835, w16836, w16837, w16838, w16839, w16840, w16841, w16842, w16843, w16844, w16845, w16846, w16847, w16848, w16849, w16850, w16851, w16852, w16853, w16854, w16855, w16856, w16857, w16858, w16859, w16860, w16861, w16862, w16863, w16864, w16865, w16866, w16867, w16868, w16869, w16870, w16871, w16872, w16873, w16874, w16875, w16876, w16877, w16878, w16879, w16880, w16881, w16882, w16883, w16884, w16885, w16886, w16887, w16888, w16889, w16890, w16891, w16892, w16893, w16894, w16895, w16896, w16897, w16898, w16899, w16900, w16901, w16902, w16903, w16904, w16905, w16906, w16907, w16908, w16909, w16910, w16911, w16912, w16913, w16914, w16915, w16916, w16917, w16918, w16919, w16920, w16921, w16922, w16923, w16924, w16925, w16926, w16927, w16928, w16929, w16930, w16931, w16932, w16933, w16934, w16935, w16936, w16937, w16938, w16939, w16940, w16941, w16942, w16943, w16944, w16945, w16946, w16947, w16948, w16949, w16950, w16951, w16952, w16953, w16954, w16955, w16956, w16957, w16958, w16959, w16960, w16961, w16962, w16963, w16964, w16965, w16966, w16967, w16968, w16969, w16970, w16971, w16972, w16973, w16974, w16975, w16976, w16977, w16978, w16979, w16980, w16981, w16982, w16983, w16984, w16985, w16986, w16987, w16988, w16989, w16990, w16991, w16992, w16993, w16994, w16995, w16996, w16997, w16998, w16999, w17000, w17001, w17002, w17003, w17004, w17005, w17006, w17007, w17008, w17009, w17010, w17011, w17012, w17013, w17014, w17015, w17016, w17017, w17018, w17019, w17020, w17021, w17022, w17023, w17024, w17025, w17026, w17027, w17028, w17029, w17030, w17031, w17032, w17033, w17034, w17035, w17036, w17037, w17038, w17039, w17040, w17041, w17042, w17043, w17044, w17045, w17046, w17047, w17048, w17049, w17050, w17051, w17052, w17053, w17054, w17055, w17056, w17057, w17058, w17059, w17060, w17061, w17062, w17063, w17064, w17065, w17066, w17067, w17068, w17069, w17070, w17071, w17072, w17073, w17074, w17075, w17076, w17077, w17078, w17079, w17080, w17081, w17082, w17083, w17084, w17085, w17086, w17087, w17088, w17089, w17090, w17091, w17092, w17093, w17094, w17095, w17096, w17097, w17098, w17099, w17100, w17101, w17102, w17103, w17104, w17105, w17106, w17107, w17108, w17109, w17110, w17111, w17112, w17113, w17114, w17115, w17116, w17117, w17118, w17119, w17120, w17121, w17122, w17123, w17124, w17125, w17126, w17127, w17128, w17129, w17130, w17131, w17132, w17133, w17134, w17135, w17136, w17137, w17138, w17139, w17140, w17141, w17142, w17143, w17144, w17145, w17146, w17147, w17148, w17149, w17150, w17151, w17152, w17153, w17154, w17155, w17156, w17157, w17158, w17159, w17160, w17161, w17162, w17163, w17164, w17165, w17166, w17167, w17168, w17169, w17170, w17171, w17172, w17173, w17174, w17175, w17176, w17177, w17178, w17179, w17180, w17181, w17182, w17183, w17184, w17185, w17186, w17187, w17188, w17189, w17190, w17191, w17192, w17193, w17194, w17195, w17196, w17197, w17198, w17199, w17200, w17201, w17202, w17203, w17204, w17205, w17206, w17207, w17208, w17209, w17210, w17211, w17212, w17213, w17214, w17215, w17216, w17217, w17218, w17219, w17220, w17221, w17222, w17223, w17224, w17225, w17226, w17227, w17228, w17229, w17230, w17231, w17232, w17233, w17234, w17235, w17236, w17237, w17238, w17239, w17240, w17241, w17242, w17243, w17244, w17245, w17246, w17247, w17248, w17249, w17250, w17251, w17252, w17253, w17254, w17255, w17256, w17257, w17258, w17259, w17260, w17261, w17262, w17263, w17264, w17265, w17266, w17267, w17268, w17269, w17270, w17271, w17272, w17273, w17274, w17275, w17276, w17277, w17278, w17279, w17280, w17281, w17282, w17283, w17284, w17285, w17286, w17287, w17288, w17289, w17290, w17291, w17292, w17293, w17294, w17295, w17296, w17297, w17298, w17299, w17300, w17301, w17302, w17303, w17304, w17305, w17306, w17307, w17308, w17309, w17310, w17311, w17312, w17313, w17314, w17315, w17316, w17317, w17318, w17319, w17320, w17321, w17322, w17323, w17324, w17325, w17326, w17327, w17328, w17329, w17330, w17331, w17332, w17333, w17334, w17335, w17336, w17337, w17338, w17339, w17340, w17341, w17342, w17343, w17344, w17345, w17346, w17347, w17348, w17349, w17350, w17351, w17352, w17353, w17354, w17355, w17356, w17357, w17358, w17359, w17360, w17361, w17362, w17363, w17364, w17365, w17366, w17367, w17368, w17369, w17370, w17371, w17372, w17373, w17374, w17375, w17376, w17377, w17378, w17379, w17380, w17381, w17382, w17383, w17384, w17385, w17386, w17387, w17388, w17389, w17390, w17391, w17392, w17393, w17394, w17395, w17396, w17397, w17398, w17399, w17400, w17401, w17402, w17403, w17404, w17405, w17406, w17407, w17408, w17409, w17410, w17411, w17412, w17413, w17414, w17415, w17416, w17417, w17418, w17419, w17420, w17421, w17422, w17423, w17424, w17425, w17426, w17427, w17428, w17429, w17430, w17431, w17432, w17433, w17434, w17435, w17436, w17437, w17438, w17439, w17440, w17441, w17442, w17443, w17444, w17445, w17446, w17447, w17448, w17449, w17450, w17451, w17452, w17453, w17454, w17455, w17456, w17457, w17458, w17459, w17460, w17461, w17462, w17463, w17464, w17465, w17466, w17467, w17468, w17469, w17470, w17471, w17472, w17473, w17474, w17475, w17476, w17477, w17478, w17479, w17480, w17481, w17482, w17483, w17484, w17485, w17486, w17487, w17488, w17489, w17490, w17491, w17492, w17493, w17494, w17495, w17496, w17497, w17498, w17499, w17500, w17501, w17502, w17503, w17504, w17505, w17506, w17507, w17508, w17509, w17510, w17511, w17512, w17513, w17514, w17515, w17516, w17517, w17518, w17519, w17520, w17521, w17522, w17523, w17524, w17525, w17526, w17527, w17528, w17529, w17530, w17531, w17532, w17533, w17534, w17535, w17536, w17537, w17538, w17539, w17540, w17541, w17542, w17543, w17544, w17545, w17546, w17547, w17548, w17549, w17550, w17551, w17552, w17553, w17554, w17555, w17556, w17557, w17558, w17559, w17560, w17561, w17562, w17563, w17564, w17565, w17566, w17567, w17568, w17569, w17570, w17571, w17572, w17573, w17574, w17575, w17576, w17577, w17578, w17579, w17580, w17581, w17582, w17583, w17584, w17585, w17586, w17587, w17588, w17589, w17590, w17591, w17592, w17593, w17594, w17595, w17596, w17597, w17598, w17599, w17600, w17601, w17602, w17603, w17604, w17605, w17606, w17607, w17608, w17609, w17610, w17611, w17612, w17613, w17614, w17615, w17616, w17617, w17618, w17619, w17620, w17621, w17622, w17623, w17624, w17625, w17626, w17627, w17628, w17629, w17630, w17631, w17632, w17633, w17634, w17635, w17636, w17637, w17638, w17639, w17640, w17641, w17642, w17643, w17644, w17645, w17646, w17647, w17648, w17649, w17650, w17651, w17652, w17653, w17654, w17655, w17656, w17657, w17658, w17659, w17660, w17661, w17662, w17663, w17664, w17665, w17666, w17667, w17668, w17669, w17670, w17671, w17672, w17673, w17674, w17675, w17676, w17677, w17678, w17679, w17680, w17681, w17682, w17683, w17684, w17685, w17686, w17687, w17688, w17689, w17690, w17691, w17692, w17693, w17694, w17695, w17696, w17697, w17698, w17699, w17700, w17701, w17702, w17703, w17704, w17705, w17706, w17707, w17708, w17709, w17710, w17711, w17712, w17713, w17714, w17715, w17716, w17717, w17718, w17719, w17720, w17721, w17722, w17723, w17724;
assign w0 = pi126 & ~pi352;
assign w1 = ~pi127 & pi353;
assign w2 = w0 & ~w1;
assign w3 = pi125 & ~pi351;
assign w4 = pi123 & ~pi349;
assign w5 = pi124 & ~pi350;
assign w6 = ~w4 & ~w5;
assign w7 = ~pi122 & pi348;
assign w8 = ~pi123 & pi349;
assign w9 = ~w7 & ~w8;
assign w10 = pi122 & ~pi348;
assign w11 = pi121 & ~pi347;
assign w12 = ~w10 & ~w11;
assign w13 = ~pi121 & pi347;
assign w14 = pi120 & ~pi346;
assign w15 = ~pi120 & pi346;
assign w16 = ~pi119 & pi345;
assign w17 = ~w15 & ~w16;
assign w18 = pi118 & ~pi344;
assign w19 = pi119 & ~pi345;
assign w20 = ~w18 & ~w19;
assign w21 = w17 & ~w20;
assign w22 = (~w13 & w21) | (~w13 & w16628) | (w21 & w16628);
assign w23 = (w9 & w22) | (w9 & w16629) | (w22 & w16629);
assign w24 = pi127 & ~pi353;
assign w25 = ~pi125 & pi351;
assign w26 = ~pi124 & pi350;
assign w27 = ~w3 & ~w24;
assign w28 = ~w25 & ~w26;
assign w29 = w27 & w28;
assign w30 = (w29 & w23) | (w29 & w16630) | (w23 & w16630);
assign w31 = ~pi126 & pi352;
assign w32 = ~w0 & ~w1;
assign w33 = ~w31 & w32;
assign w34 = (w33 & w30) | (w33 & w16631) | (w30 & w16631);
assign w35 = ~pi118 & pi344;
assign w36 = ~pi117 & pi343;
assign w37 = ~w13 & ~w14;
assign w38 = ~w35 & ~w36;
assign w39 = w37 & w38;
assign w40 = w6 & w9;
assign w41 = w12 & w17;
assign w42 = w20 & w41;
assign w43 = w39 & w40;
assign w44 = w29 & w33;
assign w45 = w43 & w44;
assign w46 = w42 & w45;
assign w47 = pi117 & ~pi343;
assign w48 = pi116 & ~pi342;
assign w49 = ~w47 & ~w48;
assign w50 = pi112 & ~pi338;
assign w51 = pi113 & ~pi339;
assign w52 = ~w50 & ~w51;
assign w53 = ~pi111 & pi337;
assign w54 = ~pi112 & pi338;
assign w55 = ~w53 & ~w54;
assign w56 = pi110 & ~pi336;
assign w57 = pi111 & ~pi337;
assign w58 = ~w56 & ~w57;
assign w59 = w55 & ~w58;
assign w60 = w52 & ~w59;
assign w61 = ~pi114 & pi340;
assign w62 = ~pi116 & pi342;
assign w63 = ~pi115 & pi341;
assign w64 = ~w62 & ~w63;
assign w65 = pi115 & ~pi341;
assign w66 = pi114 & ~pi340;
assign w67 = ~w65 & ~w66;
assign w68 = ~pi113 & pi339;
assign w69 = ~w61 & ~w68;
assign w70 = w49 & w69;
assign w71 = w64 & w67;
assign w72 = w70 & w71;
assign w73 = ~w60 & w72;
assign w74 = w64 & ~w67;
assign w75 = w49 & ~w74;
assign w76 = ~w73 & w75;
assign w77 = w46 & ~w76;
assign w78 = pi109 & ~pi335;
assign w79 = pi108 & ~pi334;
assign w80 = ~w78 & ~w79;
assign w81 = ~pi109 & pi335;
assign w82 = ~w80 & ~w81;
assign w83 = pi107 & ~pi333;
assign w84 = pi106 & ~pi332;
assign w85 = ~pi106 & pi332;
assign w86 = ~pi105 & pi331;
assign w87 = pi104 & ~pi330;
assign w88 = pi105 & ~pi331;
assign w89 = ~pi104 & pi330;
assign w90 = ~pi103 & pi329;
assign w91 = pi102 & ~pi328;
assign w92 = pi103 & ~pi329;
assign w93 = ~pi102 & pi328;
assign w94 = ~pi101 & pi327;
assign w95 = pi101 & ~pi327;
assign w96 = pi100 & ~pi326;
assign w97 = ~pi100 & pi326;
assign w98 = ~pi099 & pi325;
assign w99 = pi099 & ~pi325;
assign w100 = pi098 & ~pi324;
assign w101 = ~pi098 & pi324;
assign w102 = pi097 & ~pi323;
assign w103 = pi096 & ~pi322;
assign w104 = ~w102 & ~w103;
assign w105 = ~pi097 & pi323;
assign w106 = ~w101 & ~w105;
assign w107 = ~w104 & w106;
assign w108 = ~w99 & ~w100;
assign w109 = ~w97 & ~w98;
assign w110 = (w109 & w107) | (w109 & w16632) | (w107 & w16632);
assign w111 = ~w95 & ~w96;
assign w112 = ~w93 & ~w94;
assign w113 = ~w91 & ~w92;
assign w114 = w113 & w17620;
assign w115 = ~w89 & ~w90;
assign w116 = ~w87 & ~w88;
assign w117 = ~w85 & ~w86;
assign w118 = ~w83 & ~w84;
assign w119 = (w114 & w16637) | (w114 & w16638) | (w16637 & w16638);
assign w120 = ~pi107 & pi333;
assign w121 = ~pi108 & pi334;
assign w122 = ~w81 & ~w120;
assign w123 = ~w121 & w122;
assign w124 = w80 & w123;
assign w125 = (~w82 & w119) | (~w82 & w16639) | (w119 & w16639);
assign w126 = ~pi110 & pi336;
assign w127 = w52 & ~w126;
assign w128 = w55 & w58;
assign w129 = w127 & w128;
assign w130 = w72 & w129;
assign w131 = w46 & w130;
assign w132 = ~w125 & w131;
assign w133 = ~w24 & ~w77;
assign w134 = ~w34 & w133;
assign w135 = w134 & w16640;
assign w136 = ~pi160 & pi161;
assign w137 = w135 & w136;
assign w138 = ~pi160 & ~w137;
assign w139 = (pi162 & ~w135) | (pi162 & w16641) | (~w135 & w16641);
assign w140 = w135 & w16642;
assign w141 = ~w139 & ~w140;
assign w142 = (pi163 & ~w135) | (pi163 & w16643) | (~w135 & w16643);
assign w143 = w135 & w16644;
assign w144 = ~w142 & ~w143;
assign w145 = (pi164 & ~w135) | (pi164 & w16645) | (~w135 & w16645);
assign w146 = w135 & w16646;
assign w147 = ~w145 & ~w146;
assign w148 = (pi165 & ~w135) | (pi165 & w16647) | (~w135 & w16647);
assign w149 = w135 & w16648;
assign w150 = ~w148 & ~w149;
assign w151 = (pi166 & ~w135) | (pi166 & w16649) | (~w135 & w16649);
assign w152 = w135 & w16650;
assign w153 = ~w151 & ~w152;
assign w154 = (pi167 & ~w135) | (pi167 & w16651) | (~w135 & w16651);
assign w155 = w135 & w16652;
assign w156 = ~w154 & ~w155;
assign w157 = (pi168 & ~w135) | (pi168 & w16653) | (~w135 & w16653);
assign w158 = w135 & w16654;
assign w159 = ~w157 & ~w158;
assign w160 = (pi169 & ~w135) | (pi169 & w16655) | (~w135 & w16655);
assign w161 = w135 & w16656;
assign w162 = ~w160 & ~w161;
assign w163 = (pi170 & ~w135) | (pi170 & w16657) | (~w135 & w16657);
assign w164 = w135 & w16658;
assign w165 = ~w163 & ~w164;
assign w166 = (pi171 & ~w135) | (pi171 & w16659) | (~w135 & w16659);
assign w167 = w135 & w16660;
assign w168 = ~w166 & ~w167;
assign w169 = (pi172 & ~w135) | (pi172 & w16661) | (~w135 & w16661);
assign w170 = w135 & w16662;
assign w171 = ~w169 & ~w170;
assign w172 = (pi173 & ~w135) | (pi173 & w16663) | (~w135 & w16663);
assign w173 = w135 & w16664;
assign w174 = ~w172 & ~w173;
assign w175 = w135 & w16665;
assign w176 = (pi174 & ~w135) | (pi174 & w16666) | (~w135 & w16666);
assign w177 = ~w175 & ~w176;
assign w178 = (pi175 & ~w135) | (pi175 & w16667) | (~w135 & w16667);
assign w179 = w135 & w16668;
assign w180 = ~w178 & ~w179;
assign w181 = (pi176 & ~w135) | (pi176 & w16669) | (~w135 & w16669);
assign w182 = pi279 & w135;
assign w183 = w135 & w16670;
assign w184 = ~w181 & ~w183;
assign w185 = (pi177 & ~w135) | (pi177 & w16671) | (~w135 & w16671);
assign w186 = w135 & w16672;
assign w187 = ~w185 & ~w186;
assign w188 = (pi178 & ~w135) | (pi178 & w16673) | (~w135 & w16673);
assign w189 = pi281 & w135;
assign w190 = w135 & w16674;
assign w191 = ~w188 & ~w190;
assign w192 = (pi179 & ~w135) | (pi179 & w16675) | (~w135 & w16675);
assign w193 = pi282 & w135;
assign w194 = w135 & w16676;
assign w195 = ~w192 & ~w194;
assign w196 = (pi180 & ~w135) | (pi180 & w16677) | (~w135 & w16677);
assign w197 = w135 & w16678;
assign w198 = ~w196 & ~w197;
assign w199 = (pi181 & ~w135) | (pi181 & w16679) | (~w135 & w16679);
assign w200 = w135 & w16680;
assign w201 = ~w199 & ~w200;
assign w202 = (pi182 & ~w135) | (pi182 & w16681) | (~w135 & w16681);
assign w203 = pi285 & w135;
assign w204 = w135 & w16682;
assign w205 = ~w202 & ~w204;
assign w206 = (pi183 & ~w135) | (pi183 & w16683) | (~w135 & w16683);
assign w207 = pi286 & w135;
assign w208 = w135 & w16684;
assign w209 = ~w206 & ~w208;
assign w210 = (pi184 & ~w135) | (pi184 & w16685) | (~w135 & w16685);
assign w211 = pi287 & w135;
assign w212 = w135 & w16686;
assign w213 = ~w210 & ~w212;
assign w214 = (pi185 & ~w135) | (pi185 & w16687) | (~w135 & w16687);
assign w215 = w135 & w16688;
assign w216 = ~w214 & ~w215;
assign w217 = (pi186 & ~w135) | (pi186 & w16689) | (~w135 & w16689);
assign w218 = w135 & w16690;
assign w219 = ~w217 & ~w218;
assign w220 = (~pi187 & ~w135) | (~pi187 & w16691) | (~w135 & w16691);
assign w221 = w135 & w16692;
assign w222 = ~w220 & ~w221;
assign w223 = (pi188 & ~w135) | (pi188 & w16693) | (~w135 & w16693);
assign w224 = w135 & w16694;
assign w225 = ~w223 & ~w224;
assign w226 = (pi189 & ~w135) | (pi189 & w16695) | (~w135 & w16695);
assign w227 = w135 & w16696;
assign w228 = ~w226 & ~w227;
assign w229 = (pi190 & ~w135) | (pi190 & w16697) | (~w135 & w16697);
assign w230 = w135 & w16698;
assign w231 = ~w229 & ~w230;
assign w232 = (pi191 & ~w135) | (pi191 & w16699) | (~w135 & w16699);
assign w233 = w135 & w16700;
assign w234 = ~w232 & ~w233;
assign w235 = (pi192 & ~w135) | (pi192 & w16701) | (~w135 & w16701);
assign w236 = w135 & w16702;
assign w237 = ~w235 & ~w236;
assign w238 = (pi193 & ~w135) | (pi193 & w16703) | (~w135 & w16703);
assign w239 = w135 & w16704;
assign w240 = ~w238 & ~w239;
assign w241 = (pi194 & ~w135) | (pi194 & w16705) | (~w135 & w16705);
assign w242 = w135 & w16706;
assign w243 = ~w241 & ~w242;
assign w244 = (pi195 & ~w135) | (pi195 & w16707) | (~w135 & w16707);
assign w245 = pi323 & w135;
assign w246 = w135 & w16708;
assign w247 = ~w244 & ~w246;
assign w248 = (pi196 & ~w135) | (pi196 & w16709) | (~w135 & w16709);
assign w249 = w135 & w16710;
assign w250 = ~w248 & ~w249;
assign w251 = (pi197 & ~w135) | (pi197 & w16711) | (~w135 & w16711);
assign w252 = w135 & w16712;
assign w253 = ~w251 & ~w252;
assign w254 = (pi198 & ~w135) | (pi198 & w16713) | (~w135 & w16713);
assign w255 = w135 & w16714;
assign w256 = ~w254 & ~w255;
assign w257 = (pi199 & ~w135) | (pi199 & w16715) | (~w135 & w16715);
assign w258 = w135 & w16716;
assign w259 = ~w257 & ~w258;
assign w260 = (pi200 & ~w135) | (pi200 & w16717) | (~w135 & w16717);
assign w261 = w135 & w16718;
assign w262 = ~w260 & ~w261;
assign w263 = (pi201 & ~w135) | (pi201 & w16719) | (~w135 & w16719);
assign w264 = w135 & w16720;
assign w265 = ~w263 & ~w264;
assign w266 = (pi202 & ~w135) | (pi202 & w16721) | (~w135 & w16721);
assign w267 = w135 & w16722;
assign w268 = ~w266 & ~w267;
assign w269 = (pi203 & ~w135) | (pi203 & w16723) | (~w135 & w16723);
assign w270 = w135 & w16724;
assign w271 = ~w269 & ~w270;
assign w272 = (pi204 & ~w135) | (pi204 & w16725) | (~w135 & w16725);
assign w273 = w135 & w16726;
assign w274 = ~w272 & ~w273;
assign w275 = (pi205 & ~w135) | (pi205 & w16727) | (~w135 & w16727);
assign w276 = w135 & w16728;
assign w277 = ~w275 & ~w276;
assign w278 = (pi206 & ~w135) | (pi206 & w16729) | (~w135 & w16729);
assign w279 = pi324 & w135;
assign w280 = w135 & w16730;
assign w281 = ~w278 & ~w280;
assign w282 = (pi207 & ~w135) | (pi207 & w16731) | (~w135 & w16731);
assign w283 = w135 & w16732;
assign w284 = ~w282 & ~w283;
assign w285 = (pi208 & ~w135) | (pi208 & w16733) | (~w135 & w16733);
assign w286 = w135 & w16734;
assign w287 = ~w285 & ~w286;
assign w288 = (pi209 & ~w135) | (pi209 & w16735) | (~w135 & w16735);
assign w289 = w135 & w16736;
assign w290 = ~w288 & ~w289;
assign w291 = (pi210 & ~w135) | (pi210 & w16737) | (~w135 & w16737);
assign w292 = w135 & w16738;
assign w293 = ~w291 & ~w292;
assign w294 = (pi211 & ~w135) | (pi211 & w16739) | (~w135 & w16739);
assign w295 = w135 & w16740;
assign w296 = ~w294 & ~w295;
assign w297 = (pi212 & ~w135) | (pi212 & w16741) | (~w135 & w16741);
assign w298 = w135 & w16742;
assign w299 = ~w297 & ~w298;
assign w300 = (pi213 & ~w135) | (pi213 & w16743) | (~w135 & w16743);
assign w301 = w135 & w16744;
assign w302 = ~w300 & ~w301;
assign w303 = (pi214 & ~w135) | (pi214 & w16745) | (~w135 & w16745);
assign w304 = w135 & w16746;
assign w305 = ~w303 & ~w304;
assign w306 = (pi215 & ~w135) | (pi215 & w16747) | (~w135 & w16747);
assign w307 = w135 & w16748;
assign w308 = ~w306 & ~w307;
assign w309 = (pi216 & ~w135) | (pi216 & w16749) | (~w135 & w16749);
assign w310 = w135 & w16750;
assign w311 = ~w309 & ~w310;
assign w312 = (pi217 & ~w135) | (pi217 & w16751) | (~w135 & w16751);
assign w313 = pi325 & w135;
assign w314 = w135 & w16752;
assign w315 = ~w312 & ~w314;
assign w316 = (pi218 & ~w135) | (pi218 & w16753) | (~w135 & w16753);
assign w317 = w134 & w16754;
assign w318 = w136 & w317;
assign w319 = ~w316 & ~w318;
assign w320 = (pi219 & ~w135) | (pi219 & w16755) | (~w135 & w16755);
assign w321 = w135 & w16756;
assign w322 = ~w320 & ~w321;
assign w323 = (pi220 & ~w135) | (pi220 & w16757) | (~w135 & w16757);
assign w324 = w135 & w16758;
assign w325 = ~w323 & ~w324;
assign w326 = (pi221 & ~w135) | (pi221 & w16759) | (~w135 & w16759);
assign w327 = pi327 & w135;
assign w328 = w135 & w16760;
assign w329 = ~w326 & ~w328;
assign w330 = (pi222 & ~w135) | (pi222 & w16761) | (~w135 & w16761);
assign w331 = w135 & w16762;
assign w332 = ~w330 & ~w331;
assign w333 = (pi223 & ~w135) | (pi223 & w16763) | (~w135 & w16763);
assign w334 = pi329 & w135;
assign w335 = w135 & w16764;
assign w336 = ~w333 & ~w335;
assign w337 = (pi224 & ~w135) | (pi224 & w16765) | (~w135 & w16765);
assign w338 = pi330 & w135;
assign w339 = w135 & w16766;
assign w340 = ~w337 & ~w339;
assign w341 = (pi225 & ~w135) | (pi225 & w16767) | (~w135 & w16767);
assign w342 = w135 & w16768;
assign w343 = ~w341 & ~w342;
assign w344 = (pi226 & ~w135) | (pi226 & w16769) | (~w135 & w16769);
assign w345 = w135 & w16770;
assign w346 = ~w344 & ~w345;
assign w347 = (pi227 & ~w135) | (pi227 & w16771) | (~w135 & w16771);
assign w348 = pi320 & w135;
assign w349 = w135 & w16772;
assign w350 = ~w347 & ~w349;
assign w351 = (pi228 & ~w135) | (pi228 & w16773) | (~w135 & w16773);
assign w352 = w135 & w16774;
assign w353 = ~w351 & ~w352;
assign w354 = (pi229 & ~w135) | (pi229 & w16775) | (~w135 & w16775);
assign w355 = w135 & w16776;
assign w356 = ~w354 & ~w355;
assign w357 = (pi230 & ~w135) | (pi230 & w16777) | (~w135 & w16777);
assign w358 = w135 & w16778;
assign w359 = ~w357 & ~w358;
assign w360 = (pi231 & ~w135) | (pi231 & w16779) | (~w135 & w16779);
assign w361 = w135 & w16780;
assign w362 = ~w360 & ~w361;
assign w363 = (pi232 & ~w135) | (pi232 & w16781) | (~w135 & w16781);
assign w364 = w135 & w16782;
assign w365 = ~w363 & ~w364;
assign w366 = (pi233 & ~w135) | (pi233 & w16783) | (~w135 & w16783);
assign w367 = w135 & w16784;
assign w368 = ~w366 & ~w367;
assign w369 = (pi234 & ~w135) | (pi234 & w16785) | (~w135 & w16785);
assign w370 = w135 & w16786;
assign w371 = ~w369 & ~w370;
assign w372 = (pi235 & ~w135) | (pi235 & w16787) | (~w135 & w16787);
assign w373 = w135 & w16788;
assign w374 = ~w372 & ~w373;
assign w375 = (pi236 & ~w135) | (pi236 & w16789) | (~w135 & w16789);
assign w376 = w135 & w16790;
assign w377 = ~w375 & ~w376;
assign w378 = (pi237 & ~w135) | (pi237 & w16791) | (~w135 & w16791);
assign w379 = w135 & w16792;
assign w380 = ~w378 & ~w379;
assign w381 = (pi238 & ~w135) | (pi238 & w16793) | (~w135 & w16793);
assign w382 = pi319 & w135;
assign w383 = w135 & w16794;
assign w384 = ~w381 & ~w383;
assign w385 = (pi239 & ~w135) | (pi239 & w16795) | (~w135 & w16795);
assign w386 = w135 & w16796;
assign w387 = ~w385 & ~w386;
assign w388 = (pi240 & ~w135) | (pi240 & w16797) | (~w135 & w16797);
assign w389 = w135 & w16798;
assign w390 = ~w388 & ~w389;
assign w391 = (pi241 & ~w135) | (pi241 & w16799) | (~w135 & w16799);
assign w392 = w135 & w16800;
assign w393 = ~w391 & ~w392;
assign w394 = (pi242 & ~w135) | (pi242 & w16801) | (~w135 & w16801);
assign w395 = w135 & w16802;
assign w396 = ~w394 & ~w395;
assign w397 = (pi243 & ~w135) | (pi243 & w16803) | (~w135 & w16803);
assign w398 = w135 & w16804;
assign w399 = ~w397 & ~w398;
assign w400 = (pi244 & ~w135) | (pi244 & w16805) | (~w135 & w16805);
assign w401 = w135 & w16806;
assign w402 = ~w400 & ~w401;
assign w403 = (pi245 & ~w135) | (pi245 & w16807) | (~w135 & w16807);
assign w404 = w135 & w16808;
assign w405 = ~w403 & ~w404;
assign w406 = (pi246 & ~w135) | (pi246 & w16809) | (~w135 & w16809);
assign w407 = w135 & w16810;
assign w408 = ~w406 & ~w407;
assign w409 = (pi247 & ~w135) | (pi247 & w16811) | (~w135 & w16811);
assign w410 = w135 & w16812;
assign w411 = ~w409 & ~w410;
assign w412 = (pi248 & ~w135) | (pi248 & w16813) | (~w135 & w16813);
assign w413 = w135 & w16814;
assign w414 = ~w412 & ~w413;
assign w415 = (pi249 & ~w135) | (pi249 & w16815) | (~w135 & w16815);
assign w416 = w135 & w16816;
assign w417 = ~w415 & ~w416;
assign w418 = (pi250 & ~w135) | (pi250 & w16817) | (~w135 & w16817);
assign w419 = w135 & w16818;
assign w420 = ~w418 & ~w419;
assign w421 = (pi251 & ~w135) | (pi251 & w16819) | (~w135 & w16819);
assign w422 = w135 & w16820;
assign w423 = ~w421 & ~w422;
assign w424 = (pi252 & ~w135) | (pi252 & w16821) | (~w135 & w16821);
assign w425 = w135 & w16822;
assign w426 = ~w424 & ~w425;
assign w427 = (pi253 & ~w135) | (pi253 & w16823) | (~w135 & w16823);
assign w428 = w135 & w16824;
assign w429 = ~w427 & ~w428;
assign w430 = (pi254 & ~w135) | (pi254 & w16825) | (~w135 & w16825);
assign w431 = w135 & w16826;
assign w432 = ~w430 & ~w431;
assign w433 = (pi255 & ~w135) | (pi255 & w16827) | (~w135 & w16827);
assign w434 = w135 & w16828;
assign w435 = ~w433 & ~w434;
assign w436 = (pi256 & ~w135) | (pi256 & w16829) | (~w135 & w16829);
assign w437 = w135 & w16830;
assign w438 = ~w436 & ~w437;
assign w439 = (pi257 & ~w135) | (pi257 & w16831) | (~w135 & w16831);
assign w440 = w135 & w16832;
assign w441 = ~w439 & ~w440;
assign w442 = ~pi064 & ~pi161;
assign w443 = pi128 & ~pi258;
assign w444 = pi128 & pi322;
assign w445 = ~w443 & ~w444;
assign w446 = pi321 & ~w445;
assign w447 = ~w135 & w446;
assign w448 = pi128 & ~w135;
assign w449 = ~pi321 & ~pi322;
assign w450 = (pi258 & w135) | (pi258 & w16834) | (w135 & w16834);
assign w451 = pi161 & ~w447;
assign w452 = ~w450 & w451;
assign w453 = ~pi160 & ~w442;
assign w454 = ~w452 & w453;
assign w455 = ~pi065 & ~pi161;
assign w456 = pi128 & pi258;
assign w457 = pi323 & w456;
assign w458 = pi258 & pi259;
assign w459 = pi128 & ~pi129;
assign w460 = w458 & w459;
assign w461 = pi128 & pi259;
assign w462 = pi128 & pi129;
assign w463 = ~pi128 & ~pi129;
assign w464 = ~w462 & ~w463;
assign w465 = (~w461 & ~w464) | (~w461 & w16835) | (~w464 & w16835);
assign w466 = ~w460 & ~w465;
assign w467 = ~w465 & w16836;
assign w468 = w457 & ~w467;
assign w469 = ~w457 & w467;
assign w470 = ~w468 & ~w469;
assign w471 = pi259 & w470;
assign w472 = ~pi259 & ~w470;
assign w473 = ~w471 & ~w472;
assign w474 = ~w446 & ~w473;
assign w475 = w446 & w473;
assign w476 = ~w474 & ~w475;
assign w477 = pi128 & pi320;
assign w478 = (~w477 & ~w464) | (~w477 & w16837) | (~w464 & w16837);
assign w479 = pi320 & pi321;
assign w480 = w459 & w479;
assign w481 = ~w478 & ~w480;
assign w482 = ~w476 & w481;
assign w483 = w476 & ~w481;
assign w484 = ~w482 & ~w483;
assign w485 = ~w135 & w484;
assign w486 = (pi161 & ~w135) | (pi161 & w16838) | (~w135 & w16838);
assign w487 = ~w485 & w486;
assign w488 = ~pi160 & ~w455;
assign w489 = ~w487 & w488;
assign w490 = ~pi066 & ~pi161;
assign w491 = ~pi260 & w135;
assign w492 = ~pi128 & pi320;
assign w493 = pi128 & ~pi319;
assign w494 = ~w492 & ~w493;
assign w495 = ~pi130 & ~w463;
assign w496 = w494 & ~w495;
assign w497 = ~pi130 & ~w494;
assign w498 = pi321 & ~w496;
assign w499 = ~w497 & w498;
assign w500 = ~pi129 & pi320;
assign w501 = ~pi321 & ~w500;
assign w502 = pi128 & pi319;
assign w503 = ~w492 & ~w502;
assign w504 = w501 & ~w503;
assign w505 = pi130 & pi321;
assign w506 = w463 & w505;
assign w507 = ~pi321 & w493;
assign w508 = w500 & w507;
assign w509 = ~w504 & ~w506;
assign w510 = ~w508 & w509;
assign w511 = ~w499 & w510;
assign w512 = pi324 & w456;
assign w513 = pi130 & pi258;
assign w514 = ~pi128 & w513;
assign w515 = pi128 & ~pi260;
assign w516 = ~pi258 & pi259;
assign w517 = w515 & w516;
assign w518 = ~w514 & ~w517;
assign w519 = ~pi129 & ~w518;
assign w520 = pi129 & pi259;
assign w521 = pi128 & ~pi259;
assign w522 = ~w520 & ~w521;
assign w523 = ~pi258 & ~w515;
assign w524 = ~w522 & w523;
assign w525 = pi130 & pi260;
assign w526 = ~pi130 & ~pi260;
assign w527 = ~w525 & ~w526;
assign w528 = pi128 & ~w527;
assign w529 = pi129 & ~pi130;
assign w530 = ~pi259 & w529;
assign w531 = pi130 & pi259;
assign w532 = ~pi128 & ~w531;
assign w533 = ~w530 & w532;
assign w534 = (pi258 & w527) | (pi258 & w16839) | (w527 & w16839);
assign w535 = ~w533 & w534;
assign w536 = ~w519 & ~w524;
assign w537 = ~w535 & w536;
assign w538 = w536 & w16840;
assign w539 = ~w465 & w16842;
assign w540 = (w538 & w16843) | (w538 & w16844) | (w16843 & w16844);
assign w541 = pi322 & w456;
assign w542 = ~w539 & ~w541;
assign w543 = w542 & w17621;
assign w544 = pi324 & ~w537;
assign w545 = w536 & w16845;
assign w546 = (w541 & w537) | (w541 & w16846) | (w537 & w16846);
assign w547 = ~w545 & w546;
assign w548 = ~w547 & w16847;
assign w549 = ~w472 & w548;
assign w550 = w472 & ~w548;
assign w551 = ~w549 & ~w550;
assign w552 = pi260 & w551;
assign w553 = ~pi260 & ~w551;
assign w554 = ~w552 & ~w553;
assign w555 = w511 & w554;
assign w556 = ~w511 & ~w554;
assign w557 = ~w555 & ~w556;
assign w558 = (~w474 & ~w476) | (~w474 & w16848) | (~w476 & w16848);
assign w559 = ~w557 & ~w558;
assign w560 = (~w135 & ~w557) | (~w135 & w16849) | (~w557 & w16849);
assign w561 = ~w559 & w560;
assign w562 = (pi161 & w561) | (pi161 & w16850) | (w561 & w16850);
assign w563 = ~pi160 & ~w490;
assign w564 = ~w562 & w563;
assign w565 = ~pi067 & ~pi161;
assign w566 = (~w549 & ~w551) | (~w549 & w16851) | (~w551 & w16851);
assign w567 = pi325 & w456;
assign w568 = ~w465 & w16852;
assign w569 = (pi323 & ~w536) | (pi323 & w16853) | (~w536 & w16853);
assign w570 = ~w538 & w16854;
assign w571 = pi128 & pi261;
assign w572 = pi129 & pi260;
assign w573 = ~w461 & w572;
assign w574 = ~w571 & ~w573;
assign w575 = ~pi260 & ~w458;
assign w576 = pi129 & w571;
assign w577 = ~w575 & w576;
assign w578 = ~w574 & ~w577;
assign w579 = ~pi261 & ~w515;
assign w580 = pi258 & ~pi261;
assign w581 = ~pi260 & ~w580;
assign w582 = w520 & ~w579;
assign w583 = ~w581 & w582;
assign w584 = ~w578 & ~w583;
assign w585 = ~w456 & w520;
assign w586 = (w513 & w528) | (w513 & w15797) | (w528 & w15797);
assign w587 = ~w584 & w586;
assign w588 = w584 & ~w586;
assign w589 = ~w587 & ~w588;
assign w590 = pi131 & pi258;
assign w591 = w531 & ~w590;
assign w592 = ~w531 & w590;
assign w593 = ~w591 & ~w592;
assign w594 = ~w589 & w593;
assign w595 = w589 & ~w593;
assign w596 = ~w594 & ~w595;
assign w597 = ~pi128 & pi129;
assign w598 = w516 & w597;
assign w599 = pi259 & pi260;
assign w600 = ~pi259 & ~pi260;
assign w601 = ~w599 & ~w600;
assign w602 = pi258 & ~w601;
assign w603 = ~w601 & w16855;
assign w604 = ~pi129 & pi130;
assign w605 = ~w529 & ~w604;
assign w606 = pi258 & ~w605;
assign w607 = ~w575 & ~w599;
assign w608 = ~w606 & w607;
assign w609 = (pi128 & w608) | (pi128 & w16856) | (w608 & w16856);
assign w610 = (w604 & w602) | (w604 & w16857) | (w602 & w16857);
assign w611 = ~w598 & ~w610;
assign w612 = ~w609 & w611;
assign w613 = w596 & w612;
assign w614 = ~w596 & ~w612;
assign w615 = ~w613 & ~w614;
assign w616 = w570 & ~w615;
assign w617 = pi322 & ~w615;
assign w618 = (~w570 & w615) | (~w570 & w16858) | (w615 & w16858);
assign w619 = ~w616 & ~w618;
assign w620 = w569 & ~w619;
assign w621 = ~w569 & w619;
assign w622 = ~w620 & ~w621;
assign w623 = w536 & w16859;
assign w624 = (w512 & w539) | (w512 & w16860) | (w539 & w16860);
assign w625 = ~w623 & w624;
assign w626 = ~w622 & w625;
assign w627 = w622 & ~w625;
assign w628 = ~w626 & ~w627;
assign w629 = w568 & w628;
assign w630 = ~w568 & ~w628;
assign w631 = ~w629 & ~w630;
assign w632 = w567 & ~w631;
assign w633 = ~w567 & w631;
assign w634 = ~w632 & ~w633;
assign w635 = ~w566 & w634;
assign w636 = w566 & ~w634;
assign w637 = ~w635 & ~w636;
assign w638 = pi261 & w637;
assign w639 = ~pi261 & ~w637;
assign w640 = ~w638 & ~w639;
assign w641 = (~w556 & ~w557) | (~w556 & w16861) | (~w557 & w16861);
assign w642 = w640 & w641;
assign w643 = ~w640 & ~w641;
assign w644 = ~w642 & ~w643;
assign w645 = ~pi130 & ~w462;
assign w646 = pi129 & pi130;
assign w647 = ~pi320 & ~w646;
assign w648 = ~w645 & w647;
assign w649 = (pi131 & w648) | (pi131 & w16086) | (w648 & w16086);
assign w650 = (pi321 & w648) | (pi321 & w16543) | (w648 & w16543);
assign w651 = ~pi130 & w597;
assign w652 = pi130 & ~w597;
assign w653 = ~w651 & ~w652;
assign w654 = pi320 & ~pi321;
assign w655 = ~w653 & w654;
assign w656 = ~pi130 & pi321;
assign w657 = w502 & ~w656;
assign w658 = ~w501 & w657;
assign w659 = ~w655 & w17622;
assign w660 = w658 & w17623;
assign w661 = ~w659 & ~w660;
assign w662 = pi128 & pi318;
assign w663 = ~pi129 & pi319;
assign w664 = w662 & ~w663;
assign w665 = pi319 & w464;
assign w666 = w464 & w16862;
assign w667 = ~w664 & ~w666;
assign w668 = w661 & w667;
assign w669 = ~w661 & ~w667;
assign w670 = ~w668 & ~w669;
assign w671 = w644 & w670;
assign w672 = (~w135 & w644) | (~w135 & w16863) | (w644 & w16863);
assign w673 = ~w671 & w672;
assign w674 = (pi161 & ~w135) | (pi161 & w16864) | (~w135 & w16864);
assign w675 = ~w673 & w674;
assign w676 = ~pi160 & ~w565;
assign w677 = ~w675 & w676;
assign w678 = ~pi068 & ~pi161;
assign w679 = w661 & ~w663;
assign w680 = ~w661 & w663;
assign w681 = ~w679 & ~w680;
assign w682 = pi128 & w681;
assign w683 = pi319 & ~w653;
assign w684 = pi131 & pi132;
assign w685 = pi132 & w646;
assign w686 = (pi131 & w462) | (pi131 & w700) | (w462 & w700);
assign w687 = ~w685 & ~w686;
assign w688 = ~w684 & ~w687;
assign w689 = pi128 & pi131;
assign w690 = pi130 & ~pi131;
assign w691 = ~w689 & ~w690;
assign w692 = pi129 & ~w691;
assign w693 = ~pi130 & pi131;
assign w694 = pi132 & ~w693;
assign w695 = pi131 & ~pi132;
assign w696 = ~w694 & ~w695;
assign w697 = ~w692 & w696;
assign w698 = ~w688 & ~w697;
assign w699 = pi321 & w698;
assign w700 = pi130 & pi131;
assign w701 = pi129 & ~w700;
assign w702 = ~w691 & ~w701;
assign w703 = (w479 & w702) | (w479 & w16088) | (w702 & w16088);
assign w704 = ~w691 & w701;
assign w705 = ~pi128 & ~pi130;
assign w706 = pi129 & ~w705;
assign w707 = ~w690 & ~w693;
assign w708 = ~w706 & w707;
assign w709 = ~w704 & ~w708;
assign w710 = w703 & w709;
assign w711 = ~w703 & ~w709;
assign w712 = (pi320 & ~w709) | (pi320 & w16089) | (~w709 & w16089);
assign w713 = ~w711 & w712;
assign w714 = ~w699 & w713;
assign w715 = w699 & ~w713;
assign w716 = ~w714 & ~w715;
assign w717 = ~w659 & w665;
assign w718 = ~w660 & ~w717;
assign w719 = w716 & w718;
assign w720 = ~w716 & ~w718;
assign w721 = ~w719 & ~w720;
assign w722 = w683 & w721;
assign w723 = ~w683 & ~w721;
assign w724 = ~w722 & ~w723;
assign w725 = pi129 & ~w724;
assign w726 = ~pi129 & w724;
assign w727 = ~w725 & ~w726;
assign w728 = ~pi318 & ~w463;
assign w729 = (~w728 & ~w681) | (~w728 & w16865) | (~w681 & w16865);
assign w730 = ~w727 & w729;
assign w731 = w662 & ~w681;
assign w732 = ~pi318 & w724;
assign w733 = (w662 & ~w724) | (w662 & w16866) | (~w724 & w16866);
assign w734 = ~w732 & ~w733;
assign w735 = (~w731 & w724) | (~w731 & w16867) | (w724 & w16867);
assign w736 = ~w734 & w735;
assign w737 = ~w730 & ~w736;
assign w738 = pi128 & pi317;
assign w739 = w737 & ~w738;
assign w740 = ~w737 & w738;
assign w741 = ~w739 & ~w740;
assign w742 = pi326 & w456;
assign w743 = pi323 & ~w615;
assign w744 = pi132 & pi258;
assign w745 = pi259 & w590;
assign w746 = ~w596 & w745;
assign w747 = (w589 & w16868) | (w589 & w16869) | (w16868 & w16869);
assign w748 = (w747 & w596) | (w747 & w17582) | (w596 & w17582);
assign w749 = ~pi261 & ~w599;
assign w750 = ~w575 & ~w749;
assign w751 = w462 & w750;
assign w752 = pi129 & pi261;
assign w753 = pi128 & pi262;
assign w754 = ~w752 & ~w753;
assign w755 = w752 & w753;
assign w756 = ~w754 & ~w755;
assign w757 = w751 & ~w756;
assign w758 = ~w751 & w756;
assign w759 = ~w757 & ~w758;
assign w760 = w525 & ~w759;
assign w761 = ~w525 & w759;
assign w762 = ~w760 & ~w761;
assign w763 = (w531 & ~w584) | (w531 & w15800) | (~w584 & w15800);
assign w764 = ~w587 & ~w763;
assign w765 = w762 & ~w764;
assign w766 = ~w762 & w764;
assign w767 = ~w765 & ~w766;
assign w768 = ~w748 & ~w767;
assign w769 = w748 & w767;
assign w770 = ~w768 & ~w769;
assign w771 = ~w744 & ~w770;
assign w772 = w744 & w770;
assign w773 = ~w771 & ~w772;
assign w774 = pi129 & pi258;
assign w775 = ~w461 & w774;
assign w776 = w461 & ~w774;
assign w777 = ~w775 & ~w776;
assign w778 = w456 & w527;
assign w779 = pi260 & w443;
assign w780 = ~w514 & ~w779;
assign w781 = ~w520 & ~w780;
assign w782 = ~w513 & w585;
assign w783 = ~w779 & w782;
assign w784 = ~w778 & ~w781;
assign w785 = ~w783 & w784;
assign w786 = (~w777 & ~w784) | (~w777 & w16870) | (~w784 & w16870);
assign w787 = ~w596 & ~w786;
assign w788 = w612 & w785;
assign w789 = w596 & ~w788;
assign w790 = ~w787 & ~w789;
assign w791 = w773 & ~w790;
assign w792 = ~w773 & w790;
assign w793 = ~w791 & ~w792;
assign w794 = (w743 & w793) | (w743 & w16871) | (w793 & w16871);
assign w795 = ~w793 & w16872;
assign w796 = ~w794 & ~w795;
assign w797 = w569 & ~w618;
assign w798 = ~w616 & ~w797;
assign w799 = w796 & w798;
assign w800 = ~w796 & ~w798;
assign w801 = ~w799 & ~w800;
assign w802 = (~w626 & ~w628) | (~w626 & w16873) | (~w628 & w16873);
assign w803 = w544 & ~w802;
assign w804 = ~w544 & w802;
assign w805 = ~w803 & ~w804;
assign w806 = w801 & w805;
assign w807 = ~w801 & ~w805;
assign w808 = ~w806 & ~w807;
assign w809 = ~w465 & w16874;
assign w810 = w628 & w16876;
assign w811 = (w628 & w16877) | (w628 & w16878) | (w16877 & w16878);
assign w812 = ~w810 & w811;
assign w813 = ~w808 & w812;
assign w814 = w808 & ~w812;
assign w815 = ~w813 & ~w814;
assign w816 = w742 & ~w815;
assign w817 = ~w742 & w815;
assign w818 = ~w816 & ~w817;
assign w819 = (~w635 & ~w637) | (~w635 & w16879) | (~w637 & w16879);
assign w820 = ~w818 & ~w819;
assign w821 = w818 & w819;
assign w822 = ~w820 & ~w821;
assign w823 = pi262 & w822;
assign w824 = ~pi262 & ~w822;
assign w825 = ~w823 & ~w824;
assign w826 = (~w642 & ~w644) | (~w642 & w16880) | (~w644 & w16880);
assign w827 = w825 & ~w826;
assign w828 = ~w825 & w826;
assign w829 = ~w827 & ~w828;
assign w830 = ~w741 & w829;
assign w831 = (~w135 & w829) | (~w135 & w16881) | (w829 & w16881);
assign w832 = ~w830 & w831;
assign w833 = (pi161 & ~w135) | (pi161 & w16882) | (~w135 & w16882);
assign w834 = ~w832 & w833;
assign w835 = ~pi160 & ~w678;
assign w836 = ~w834 & w835;
assign w837 = ~pi069 & ~pi161;
assign w838 = pi128 & pi316;
assign w839 = pi129 & ~w737;
assign w840 = ~w462 & w737;
assign w841 = ~w839 & ~w840;
assign w842 = pi317 & ~w463;
assign w843 = ~w841 & w842;
assign w844 = pi318 & ~w653;
assign w845 = pi319 & w709;
assign w846 = pi132 & pi133;
assign w847 = ~w684 & ~w685;
assign w848 = pi133 & w686;
assign w849 = w847 & ~w848;
assign w850 = ~w846 & ~w849;
assign w851 = ~pi132 & ~pi133;
assign w852 = ~w846 & ~w851;
assign w853 = w847 & ~w852;
assign w854 = w687 & w853;
assign w855 = ~w850 & ~w854;
assign w856 = pi321 & w855;
assign w857 = ~w698 & w710;
assign w858 = w698 & w711;
assign w859 = ~w857 & ~w858;
assign w860 = pi320 & ~w859;
assign w861 = w856 & ~w860;
assign w862 = ~w856 & w857;
assign w863 = w711 & ~w855;
assign w864 = (w698 & w863) | (w698 & w16883) | (w863 & w16883);
assign w865 = ~w862 & ~w864;
assign w866 = pi320 & ~w865;
assign w867 = ~w861 & ~w866;
assign w868 = (~w720 & ~w721) | (~w720 & w16545) | (~w721 & w16545);
assign w869 = w867 & w868;
assign w870 = ~w867 & ~w868;
assign w871 = ~w869 & ~w870;
assign w872 = w845 & w871;
assign w873 = ~w845 & ~w871;
assign w874 = ~w872 & ~w873;
assign w875 = (w682 & ~w724) | (w682 & w16884) | (~w724 & w16884);
assign w876 = pi318 & ~w463;
assign w877 = (w876 & w724) | (w876 & w16885) | (w724 & w16885);
assign w878 = ~w875 & w877;
assign w879 = ~w874 & ~w878;
assign w880 = w874 & w878;
assign w881 = ~w879 & ~w880;
assign w882 = w844 & ~w881;
assign w883 = ~w844 & w881;
assign w884 = ~w882 & ~w883;
assign w885 = ~w843 & w884;
assign w886 = w843 & ~w884;
assign w887 = ~w885 & ~w886;
assign w888 = w838 & w887;
assign w889 = ~w838 & ~w887;
assign w890 = ~w888 & ~w889;
assign w891 = (~w820 & ~w822) | (~w820 & w16886) | (~w822 & w16886);
assign w892 = pi327 & w456;
assign w893 = ~w465 & w16887;
assign w894 = (~w803 & ~w801) | (~w803 & w16888) | (~w801 & w16888);
assign w895 = pi324 & ~w615;
assign w896 = pi133 & pi258;
assign w897 = pi132 & pi259;
assign w898 = pi131 & pi260;
assign w899 = ~w761 & ~w764;
assign w900 = ~w760 & ~w899;
assign w901 = w750 & w15801;
assign w902 = ~pi261 & w599;
assign w903 = pi262 & w462;
assign w904 = ~w902 & w903;
assign w905 = ~w901 & ~w904;
assign w906 = pi129 & pi262;
assign w907 = pi128 & pi263;
assign w908 = ~w906 & ~w907;
assign w909 = w906 & w907;
assign w910 = ~w908 & ~w909;
assign w911 = pi130 & w910;
assign w912 = ~w905 & w911;
assign w913 = (~w753 & ~w750) | (~w753 & w15802) | (~w750 & w15802);
assign w914 = ~w908 & w913;
assign w915 = w902 & w909;
assign w916 = ~w577 & ~w755;
assign w917 = ~w915 & w916;
assign w918 = (~w910 & ~w916) | (~w910 & w15803) | (~w916 & w15803);
assign w919 = (~pi130 & w918) | (~pi130 & w16889) | (w918 & w16889);
assign w920 = pi130 & pi261;
assign w921 = ~w910 & w920;
assign w922 = w913 & w921;
assign w923 = w910 & ~w920;
assign w924 = ~w921 & ~w923;
assign w925 = ~pi261 & ~pi262;
assign w926 = w462 & ~w925;
assign w927 = w750 & w926;
assign w928 = (~w752 & ~w750) | (~w752 & w16090) | (~w750 & w16090);
assign w929 = (~w915 & w924) | (~w915 & w16091) | (w924 & w16091);
assign w930 = ~w912 & ~w922;
assign w931 = w930 & w16890;
assign w932 = w900 & ~w931;
assign w933 = ~w900 & w931;
assign w934 = ~w932 & ~w933;
assign w935 = ~w898 & w934;
assign w936 = w898 & ~w934;
assign w937 = ~w935 & ~w936;
assign w938 = (~w746 & ~w748) | (~w746 & w15804) | (~w748 & w15804);
assign w939 = w937 & ~w938;
assign w940 = ~w937 & w938;
assign w941 = ~w939 & ~w940;
assign w942 = ~w897 & ~w941;
assign w943 = w897 & w941;
assign w944 = ~w942 & ~w943;
assign w945 = ~w773 & ~w789;
assign w946 = (~w787 & w773) | (~w787 & w16891) | (w773 & w16891);
assign w947 = w771 & ~w946;
assign w948 = ~w771 & w17624;
assign w949 = ~w947 & ~w948;
assign w950 = w944 & ~w949;
assign w951 = ~w944 & w949;
assign w952 = ~w950 & ~w951;
assign w953 = w896 & w952;
assign w954 = ~w896 & ~w952;
assign w955 = ~w953 & ~w954;
assign w956 = pi322 & ~w955;
assign w957 = pi323 & ~w793;
assign w958 = (~w957 & w796) | (~w957 & w16893) | (w796 & w16893);
assign w959 = w957 & w17625;
assign w960 = ~w958 & ~w959;
assign w961 = ~w956 & w960;
assign w962 = w956 & ~w960;
assign w963 = ~w961 & ~w962;
assign w964 = w895 & ~w963;
assign w965 = ~w895 & w963;
assign w966 = ~w964 & ~w965;
assign w967 = ~w894 & w966;
assign w968 = w894 & ~w966;
assign w969 = ~w967 & ~w968;
assign w970 = (~w466 & ~w628) | (~w466 & w16895) | (~w628 & w16895);
assign w971 = ~w465 & w16896;
assign w972 = w631 & w971;
assign w973 = (~w972 & ~w808) | (~w972 & w16897) | (~w808 & w16897);
assign w974 = (w808 & w16898) | (w808 & w16899) | (w16898 & w16899);
assign w975 = (pi325 & ~w973) | (pi325 & w16900) | (~w973 & w16900);
assign w976 = ~w974 & w975;
assign w977 = w969 & w976;
assign w978 = ~w969 & ~w976;
assign w979 = ~w977 & ~w978;
assign w980 = w816 & w979;
assign w981 = ~w816 & ~w979;
assign w982 = ~w980 & ~w981;
assign w983 = ~w893 & ~w982;
assign w984 = w893 & w982;
assign w985 = ~w983 & ~w984;
assign w986 = w892 & ~w985;
assign w987 = ~w892 & w985;
assign w988 = ~w986 & ~w987;
assign w989 = ~w891 & w988;
assign w990 = w891 & ~w988;
assign w991 = ~w989 & ~w990;
assign w992 = pi263 & w991;
assign w993 = ~pi263 & ~w991;
assign w994 = ~w992 & ~w993;
assign w995 = (~w827 & ~w829) | (~w827 & w16901) | (~w829 & w16901);
assign w996 = w994 & ~w995;
assign w997 = ~w994 & w995;
assign w998 = ~w996 & ~w997;
assign w999 = w890 & ~w998;
assign w1000 = (~w135 & ~w998) | (~w135 & w16902) | (~w998 & w16902);
assign w1001 = ~w999 & w1000;
assign w1002 = (pi161 & ~w135) | (pi161 & w16903) | (~w135 & w16903);
assign w1003 = ~w1001 & w1002;
assign w1004 = ~pi160 & ~w837;
assign w1005 = ~w1003 & w1004;
assign w1006 = ~pi070 & ~pi161;
assign w1007 = pi328 & w456;
assign w1008 = (pi326 & ~w536) | (pi326 & w16904) | (~w536 & w16904);
assign w1009 = pi325 & ~w615;
assign w1010 = (w808 & w16905) | (w808 & w16906) | (w16905 & w16906);
assign w1011 = ~w1009 & w17626;
assign w1012 = (w969 & w16908) | (w969 & w16909) | (w16908 & w16909);
assign w1013 = ~w1011 & ~w1012;
assign w1014 = pi324 & ~w793;
assign w1015 = (~w964 & ~w966) | (~w964 & w16910) | (~w966 & w16910);
assign w1016 = w1014 & ~w1015;
assign w1017 = ~w1014 & w1015;
assign w1018 = ~w1016 & ~w1017;
assign w1019 = (w772 & w941) | (w772 & w16092) | (w941 & w16092);
assign w1020 = ~w943 & ~w1019;
assign w1021 = pi132 & pi260;
assign w1022 = ~w918 & w16093;
assign w1023 = w929 & w1022;
assign w1024 = (pi261 & ~w462) | (pi261 & w16911) | (~w462 & w16911);
assign w1025 = (w1024 & ~w750) | (w1024 & w16912) | (~w750 & w16912);
assign w1026 = w911 & w1025;
assign w1027 = ~w917 & w921;
assign w1028 = ~w1026 & ~w1027;
assign w1029 = ~w760 & w1028;
assign w1030 = ~w899 & w1029;
assign w1031 = ~w1023 & ~w1030;
assign w1032 = pi131 & pi261;
assign w1033 = pi130 & pi262;
assign w1034 = ~w755 & ~w909;
assign w1035 = (~w908 & w927) | (~w908 & w15805) | (w927 & w15805);
assign w1036 = pi129 & pi263;
assign w1037 = pi128 & pi264;
assign w1038 = ~w1036 & ~w1037;
assign w1039 = w1036 & w1037;
assign w1040 = ~w1038 & ~w1039;
assign w1041 = w1035 & ~w1040;
assign w1042 = ~w1035 & w1040;
assign w1043 = ~w1041 & ~w1042;
assign w1044 = ~w1033 & w1043;
assign w1045 = w1033 & ~w1043;
assign w1046 = ~w1044 & ~w1045;
assign w1047 = w1032 & ~w1046;
assign w1048 = ~w1032 & w1046;
assign w1049 = ~w1047 & ~w1048;
assign w1050 = w1031 & w1049;
assign w1051 = ~w1031 & ~w1049;
assign w1052 = ~w1050 & ~w1051;
assign w1053 = ~w936 & w938;
assign w1054 = ~w935 & ~w1053;
assign w1055 = w1052 & ~w1054;
assign w1056 = ~w1052 & w1054;
assign w1057 = ~w1055 & ~w1056;
assign w1058 = ~w1021 & ~w1057;
assign w1059 = w1021 & w1052;
assign w1060 = w1054 & w1059;
assign w1061 = w1021 & ~w1052;
assign w1062 = ~w1054 & w1061;
assign w1063 = ~w1060 & ~w1062;
assign w1064 = ~w1058 & w1063;
assign w1065 = w1020 & ~w1064;
assign w1066 = ~w1020 & w1064;
assign w1067 = ~w1065 & ~w1066;
assign w1068 = pi259 & ~w744;
assign w1069 = ~w772 & ~w941;
assign w1070 = (pi258 & ~w770) | (pi258 & w16094) | (~w770 & w16094);
assign w1071 = w941 & ~w1070;
assign w1072 = ~w1069 & ~w1071;
assign w1073 = w1068 & w1072;
assign w1074 = (pi133 & w1072) | (pi133 & w16095) | (w1072 & w16095);
assign w1075 = ~w1073 & w1074;
assign w1076 = w1067 & w1075;
assign w1077 = ~w1067 & ~w1075;
assign w1078 = ~w1076 & ~w1077;
assign w1079 = pi134 & pi258;
assign w1080 = ~w1078 & ~w1079;
assign w1081 = w1078 & w1079;
assign w1082 = ~w1080 & ~w1081;
assign w1083 = w772 & w944;
assign w1084 = ~w772 & ~w944;
assign w1085 = ~w1083 & ~w1084;
assign w1086 = w896 & w1085;
assign w1087 = ~w896 & ~w1085;
assign w1088 = ~w1086 & ~w1087;
assign w1089 = w946 & w1088;
assign w1090 = ~w946 & ~w1088;
assign w1091 = ~w1089 & ~w1090;
assign w1092 = ~w1082 & ~w1091;
assign w1093 = ~w1082 & w1088;
assign w1094 = w1082 & ~w1088;
assign w1095 = ~w1093 & ~w1094;
assign w1096 = (w773 & w1088) | (w773 & w16913) | (w1088 & w16913);
assign w1097 = ~w1095 & w1096;
assign w1098 = (~w773 & ~w1088) | (~w773 & w16914) | (~w1088 & w16914);
assign w1099 = w1095 & w1098;
assign w1100 = (~w1092 & w1095) | (~w1092 & w16096) | (w1095 & w16096);
assign w1101 = ~w1099 & w1100;
assign w1102 = pi322 & w1101;
assign w1103 = ~w955 & w16915;
assign w1104 = (~w959 & w955) | (~w959 & w16916) | (w955 & w16916);
assign w1105 = ~w1103 & ~w1104;
assign w1106 = w1101 & w16917;
assign w1107 = (w1105 & ~w1101) | (w1105 & w16918) | (~w1101 & w16918);
assign w1108 = ~w1106 & ~w1107;
assign w1109 = w1018 & ~w1108;
assign w1110 = ~w1018 & w1108;
assign w1111 = ~w1109 & ~w1110;
assign w1112 = w1013 & w1111;
assign w1113 = ~w1013 & ~w1111;
assign w1114 = ~w1112 & ~w1113;
assign w1115 = w1008 & w1114;
assign w1116 = ~w1008 & ~w1114;
assign w1117 = ~w1115 & ~w1116;
assign w1118 = (~w980 & ~w982) | (~w980 & w16919) | (~w982 & w16919);
assign w1119 = ~w1117 & ~w1118;
assign w1120 = w1117 & w1118;
assign w1121 = ~w1119 & ~w1120;
assign w1122 = ~w465 & w16920;
assign w1123 = (~w1122 & ~w982) | (~w1122 & w16921) | (~w982 & w16921);
assign w1124 = w982 & w16922;
assign w1125 = pi327 & ~w1123;
assign w1126 = ~w1124 & w1125;
assign w1127 = w1121 & ~w1126;
assign w1128 = ~w1121 & w1126;
assign w1129 = ~w1127 & ~w1128;
assign w1130 = w1007 & w1129;
assign w1131 = ~w1007 & ~w1129;
assign w1132 = ~w1130 & ~w1131;
assign w1133 = (~w989 & ~w991) | (~w989 & w16923) | (~w991 & w16923);
assign w1134 = ~w1132 & ~w1133;
assign w1135 = w1132 & w1133;
assign w1136 = ~w1134 & ~w1135;
assign w1137 = pi264 & w1136;
assign w1138 = ~pi264 & ~w1136;
assign w1139 = ~w1137 & ~w1138;
assign w1140 = (~w890 & w994) | (~w890 & w16924) | (w994 & w16924);
assign w1141 = ~w996 & ~w1140;
assign w1142 = w1139 & ~w1141;
assign w1143 = ~w1139 & w1141;
assign w1144 = ~w1142 & ~w1143;
assign w1145 = pi128 & pi315;
assign w1146 = ~w737 & w16925;
assign w1147 = ~w886 & ~w1146;
assign w1148 = pi318 & w709;
assign w1149 = (~w844 & ~w874) | (~w844 & w16926) | (~w874 & w16926);
assign w1150 = ~w879 & ~w1149;
assign w1151 = pi319 & w698;
assign w1152 = pi320 & w855;
assign w1153 = ~w846 & w849;
assign w1154 = w849 & w16927;
assign w1155 = (pi134 & ~w849) | (pi134 & w16928) | (~w849 & w16928);
assign w1156 = ~w1154 & ~w1155;
assign w1157 = pi133 & w1156;
assign w1158 = ~pi133 & ~w1156;
assign w1159 = ~w1157 & ~w1158;
assign w1160 = (w710 & w856) | (w710 & w16546) | (w856 & w16546);
assign w1161 = (pi320 & w1160) | (pi320 & w15807) | (w1160 & w15807);
assign w1162 = w1159 & w1161;
assign w1163 = (w1160 & w1152) | (w1160 & w16097) | (w1152 & w16097);
assign w1164 = ~w1159 & ~w1163;
assign w1165 = (pi321 & w1163) | (pi321 & w16929) | (w1163 & w16929);
assign w1166 = ~w1161 & ~w1165;
assign w1167 = ~w1166 & w16930;
assign w1168 = (w1152 & w1166) | (w1152 & w16931) | (w1166 & w16931);
assign w1169 = ~w1167 & ~w1168;
assign w1170 = w1169 & w17627;
assign w1171 = (w871 & w16932) | (w871 & w16933) | (w16932 & w16933);
assign w1172 = ~w1170 & ~w1171;
assign w1173 = w1151 & ~w1172;
assign w1174 = ~w1151 & w1172;
assign w1175 = ~w1173 & ~w1174;
assign w1176 = ~w1150 & w1175;
assign w1177 = w1150 & ~w1175;
assign w1178 = ~w1176 & ~w1177;
assign w1179 = w1148 & w1178;
assign w1180 = ~w1148 & ~w1178;
assign w1181 = ~w1179 & ~w1180;
assign w1182 = ~w1147 & w1181;
assign w1183 = w1147 & ~w1181;
assign w1184 = ~w1182 & ~w1183;
assign w1185 = pi317 & ~w653;
assign w1186 = w1184 & w1185;
assign w1187 = ~w1184 & ~w1185;
assign w1188 = ~w1186 & ~w1187;
assign w1189 = (~pi129 & w887) | (~pi129 & w463) | (w887 & w463);
assign w1190 = (pi316 & w887) | (pi316 & w16934) | (w887 & w16934);
assign w1191 = ~w1189 & w1190;
assign w1192 = ~w1188 & ~w1191;
assign w1193 = w1188 & w1191;
assign w1194 = ~w1192 & ~w1193;
assign w1195 = ~w1145 & ~w1194;
assign w1196 = w1145 & w1194;
assign w1197 = ~w1195 & ~w1196;
assign w1198 = w1144 & ~w1197;
assign w1199 = (~w135 & w1144) | (~w135 & w16935) | (w1144 & w16935);
assign w1200 = ~w1198 & w1199;
assign w1201 = (pi161 & ~w135) | (pi161 & w16936) | (~w135 & w16936);
assign w1202 = ~w1200 & w1201;
assign w1203 = ~pi160 & ~w1006;
assign w1204 = ~w1202 & w1203;
assign w1205 = ~pi071 & ~pi161;
assign w1206 = pi128 & pi314;
assign w1207 = pi317 & w709;
assign w1208 = (~w1182 & ~w1184) | (~w1182 & w16937) | (~w1184 & w16937);
assign w1209 = pi318 & w698;
assign w1210 = w1148 & ~w1176;
assign w1211 = ~w1177 & ~w1210;
assign w1212 = pi319 & w855;
assign w1213 = w855 & w1159;
assign w1214 = pi134 & ~pi135;
assign w1215 = ~pi134 & pi135;
assign w1216 = ~w1214 & ~w1215;
assign w1217 = (~w1155 & ~w1156) | (~w1155 & w16938) | (~w1156 & w16938);
assign w1218 = w1216 & w1217;
assign w1219 = ~w1216 & ~w1217;
assign w1220 = ~w1218 & ~w1219;
assign w1221 = ~w1213 & ~w1220;
assign w1222 = ~w1162 & w1221;
assign w1223 = (pi320 & w1222) | (pi320 & w16939) | (w1222 & w16939);
assign w1224 = ~w1164 & w1223;
assign w1225 = ~w855 & w1159;
assign w1226 = ~w1163 & ~w1225;
assign w1227 = (pi320 & ~w1161) | (pi320 & w16940) | (~w1161 & w16940);
assign w1228 = ~w1226 & w1227;
assign w1229 = pi321 & w1220;
assign w1230 = ~w1228 & w1229;
assign w1231 = ~w1224 & ~w1230;
assign w1232 = w1151 & ~w1170;
assign w1233 = ~w1232 & w16941;
assign w1234 = (~w1231 & w1232) | (~w1231 & w16942) | (w1232 & w16942);
assign w1235 = ~w1233 & ~w1234;
assign w1236 = w1212 & ~w1235;
assign w1237 = ~w1212 & w1235;
assign w1238 = ~w1236 & ~w1237;
assign w1239 = w1211 & w1238;
assign w1240 = ~w1211 & ~w1238;
assign w1241 = ~w1239 & ~w1240;
assign w1242 = w1209 & w1241;
assign w1243 = ~w1209 & ~w1241;
assign w1244 = ~w1242 & ~w1243;
assign w1245 = w1208 & ~w1244;
assign w1246 = ~w1208 & w1244;
assign w1247 = ~w1245 & ~w1246;
assign w1248 = w1207 & w1247;
assign w1249 = ~w1207 & ~w1247;
assign w1250 = ~w1248 & ~w1249;
assign w1251 = w887 & w16943;
assign w1252 = (~w1251 & ~w1188) | (~w1251 & w16944) | (~w1188 & w16944);
assign w1253 = w1250 & ~w1252;
assign w1254 = ~w1250 & w1252;
assign w1255 = ~w1253 & ~w1254;
assign w1256 = pi316 & ~w653;
assign w1257 = w1255 & w1256;
assign w1258 = ~w1255 & ~w1256;
assign w1259 = ~w1257 & ~w1258;
assign w1260 = (~pi129 & w1194) | (~pi129 & w463) | (w1194 & w463);
assign w1261 = (pi315 & w1194) | (pi315 & w16945) | (w1194 & w16945);
assign w1262 = ~w1260 & w1261;
assign w1263 = ~w1259 & ~w1262;
assign w1264 = w1259 & w1262;
assign w1265 = ~w1263 & ~w1264;
assign w1266 = w1206 & ~w1265;
assign w1267 = ~w1206 & w1265;
assign w1268 = ~w1266 & ~w1267;
assign w1269 = pi329 & w456;
assign w1270 = ~w465 & w16946;
assign w1271 = (~w1270 & ~w1129) | (~w1270 & w16947) | (~w1129 & w16947);
assign w1272 = w1129 & w16948;
assign w1273 = ~w1271 & ~w1272;
assign w1274 = pi326 & ~w615;
assign w1275 = pi325 & ~w793;
assign w1276 = (w1111 & w16950) | (w1111 & w16951) | (w16950 & w16951);
assign w1277 = ~w1275 & w17628;
assign w1278 = ~w1276 & ~w1277;
assign w1279 = pi324 & ~w955;
assign w1280 = pi135 & pi258;
assign w1281 = (w1101 & w16952) | (w1101 & w16953) | (w16952 & w16953);
assign w1282 = pi134 & pi259;
assign w1283 = w1085 & w16098;
assign w1284 = ~w1076 & ~w1283;
assign w1285 = pi133 & pi260;
assign w1286 = ~w943 & w1063;
assign w1287 = ~w1019 & w1286;
assign w1288 = ~w1058 & ~w1287;
assign w1289 = pi131 & pi262;
assign w1290 = ~w1023 & ~w1044;
assign w1291 = ~w1030 & w1290;
assign w1292 = ~w1045 & ~w1291;
assign w1293 = pi130 & pi263;
assign w1294 = pi129 & pi264;
assign w1295 = pi128 & pi265;
assign w1296 = ~w1294 & ~w1295;
assign w1297 = w1294 & w1295;
assign w1298 = ~w1296 & ~w1297;
assign w1299 = (w1035 & w16099) | (w1035 & w16100) | (w16099 & w16100);
assign w1300 = w1298 & w17629;
assign w1301 = ~w1299 & ~w1300;
assign w1302 = w1293 & ~w1301;
assign w1303 = ~w1293 & w1301;
assign w1304 = ~w1302 & ~w1303;
assign w1305 = ~w1291 & w16101;
assign w1306 = (~w1304 & w1291) | (~w1304 & w16102) | (w1291 & w16102);
assign w1307 = ~w1305 & ~w1306;
assign w1308 = ~w1289 & w1307;
assign w1309 = w1289 & ~w1307;
assign w1310 = ~w1308 & ~w1309;
assign w1311 = w1032 & w1052;
assign w1312 = ~w1056 & w16103;
assign w1313 = (~w1310 & w1056) | (~w1310 & w16104) | (w1056 & w16104);
assign w1314 = ~w1312 & ~w1313;
assign w1315 = (w1314 & w1287) | (w1314 & w16105) | (w1287 & w16105);
assign w1316 = ~w1287 & w16106;
assign w1317 = ~w1315 & ~w1316;
assign w1318 = pi132 & pi261;
assign w1319 = w1317 & w1318;
assign w1320 = ~w1317 & ~w1318;
assign w1321 = ~w1319 & ~w1320;
assign w1322 = w1285 & w1321;
assign w1323 = ~w1285 & ~w1321;
assign w1324 = ~w1322 & ~w1323;
assign w1325 = w1284 & ~w1324;
assign w1326 = ~w1284 & w1324;
assign w1327 = ~w1325 & ~w1326;
assign w1328 = w1080 & ~w1327;
assign w1329 = ~w1080 & w1327;
assign w1330 = ~w1328 & ~w1329;
assign w1331 = w1282 & w1330;
assign w1332 = ~w1282 & ~w1330;
assign w1333 = ~w1331 & ~w1332;
assign w1334 = w1281 & ~w1333;
assign w1335 = ~w1281 & w1333;
assign w1336 = ~w1334 & ~w1335;
assign w1337 = w1280 & w1336;
assign w1338 = ~w1280 & ~w1336;
assign w1339 = ~w1337 & ~w1338;
assign w1340 = (~w1103 & ~w1101) | (~w1103 & w16954) | (~w1101 & w16954);
assign w1341 = w1102 & ~w1104;
assign w1342 = ~w1340 & ~w1341;
assign w1343 = w1339 & w16955;
assign w1344 = (~w1342 & ~w1339) | (~w1342 & w16956) | (~w1339 & w16956);
assign w1345 = ~w1343 & ~w1344;
assign w1346 = ~w1279 & ~w1345;
assign w1347 = w1279 & w1345;
assign w1348 = ~w1346 & ~w1347;
assign w1349 = (~w1016 & w1108) | (~w1016 & w16957) | (w1108 & w16957);
assign w1350 = w1348 & ~w1349;
assign w1351 = ~w1348 & w1349;
assign w1352 = ~w1350 & ~w1351;
assign w1353 = w1278 & ~w1352;
assign w1354 = ~w1278 & w1352;
assign w1355 = ~w1353 & ~w1354;
assign w1356 = ~w1274 & w1355;
assign w1357 = w1274 & ~w1355;
assign w1358 = ~w1356 & ~w1357;
assign w1359 = (~w1116 & ~w1117) | (~w1116 & w16958) | (~w1117 & w16958);
assign w1360 = w1358 & w1359;
assign w1361 = ~w1358 & ~w1359;
assign w1362 = ~w1360 & ~w1361;
assign w1363 = (pi327 & ~w536) | (pi327 & w16959) | (~w536 & w16959);
assign w1364 = w456 & w985;
assign w1365 = w1121 & ~w1364;
assign w1366 = (~w466 & w1121) | (~w466 & w16960) | (w1121 & w16960);
assign w1367 = pi327 & ~w1365;
assign w1368 = ~w1366 & w1367;
assign w1369 = (w1363 & ~w1367) | (w1363 & w16961) | (~w1367 & w16961);
assign w1370 = w1367 & w16962;
assign w1371 = ~w1369 & ~w1370;
assign w1372 = w1362 & ~w1371;
assign w1373 = ~w1362 & w1371;
assign w1374 = ~w1372 & ~w1373;
assign w1375 = w1273 & w1374;
assign w1376 = ~w1273 & ~w1374;
assign w1377 = ~w1375 & ~w1376;
assign w1378 = w1269 & w1377;
assign w1379 = ~w1269 & ~w1377;
assign w1380 = ~w1378 & ~w1379;
assign w1381 = (~w1134 & ~w1136) | (~w1134 & w16963) | (~w1136 & w16963);
assign w1382 = ~w1380 & ~w1381;
assign w1383 = w1380 & w1381;
assign w1384 = ~w1382 & ~w1383;
assign w1385 = pi265 & w1384;
assign w1386 = ~pi265 & ~w1384;
assign w1387 = ~w1385 & ~w1386;
assign w1388 = (~w1142 & ~w1144) | (~w1142 & w16964) | (~w1144 & w16964);
assign w1389 = w1387 & ~w1388;
assign w1390 = ~w1387 & w1388;
assign w1391 = ~w1389 & ~w1390;
assign w1392 = (w1268 & w1387) | (w1268 & w16965) | (w1387 & w16965);
assign w1393 = ~w1389 & w1392;
assign w1394 = (~w135 & w1391) | (~w135 & w16966) | (w1391 & w16966);
assign w1395 = ~w1393 & w1394;
assign w1396 = (pi161 & ~w135) | (pi161 & w16967) | (~w135 & w16967);
assign w1397 = ~w1395 & w1396;
assign w1398 = ~pi160 & ~w1205;
assign w1399 = ~w1397 & w1398;
assign w1400 = ~pi072 & ~pi161;
assign w1401 = pi128 & pi313;
assign w1402 = pi315 & ~w653;
assign w1403 = pi316 & w709;
assign w1404 = pi317 & w698;
assign w1405 = (~w1246 & ~w1247) | (~w1246 & w16968) | (~w1247 & w16968);
assign w1406 = pi318 & w855;
assign w1407 = pi319 & w1159;
assign w1408 = pi135 & ~pi136;
assign w1409 = ~pi135 & pi136;
assign w1410 = ~w1408 & ~w1409;
assign w1411 = (w849 & w16971) | (w849 & w16972) | (w16971 & w16972);
assign w1412 = (~pi134 & w1153) | (~pi134 & w16973) | (w1153 & w16973);
assign w1413 = (w1410 & w1412) | (w1410 & w16974) | (w1412 & w16974);
assign w1414 = pi134 & w1409;
assign w1415 = (~w1414 & w1153) | (~w1414 & w16975) | (w1153 & w16975);
assign w1416 = pi133 & ~w1415;
assign w1417 = pi134 & ~w1410;
assign w1418 = (w1417 & ~w849) | (w1417 & w16976) | (~w849 & w16976);
assign w1419 = ~w1416 & ~w1418;
assign w1420 = ~w1413 & w1419;
assign w1421 = w1419 & w16977;
assign w1422 = ~w1222 & w16978;
assign w1423 = ~w1220 & ~w1422;
assign w1424 = w1220 & ~w1223;
assign w1425 = ~w1423 & ~w1424;
assign w1426 = w1421 & ~w1425;
assign w1427 = ~w1421 & w1425;
assign w1428 = ~w1426 & ~w1427;
assign w1429 = w1212 & ~w1233;
assign w1430 = ~w1429 & w16979;
assign w1431 = (~w1428 & w1429) | (~w1428 & w16980) | (w1429 & w16980);
assign w1432 = ~w1430 & ~w1431;
assign w1433 = w1407 & ~w1432;
assign w1434 = ~w1407 & w1432;
assign w1435 = ~w1433 & ~w1434;
assign w1436 = (w1209 & ~w1211) | (w1209 & w16981) | (~w1211 & w16981);
assign w1437 = ~w1240 & ~w1436;
assign w1438 = w1435 & w1437;
assign w1439 = ~w1435 & ~w1437;
assign w1440 = ~w1438 & ~w1439;
assign w1441 = w1406 & w1440;
assign w1442 = ~w1406 & ~w1440;
assign w1443 = ~w1441 & ~w1442;
assign w1444 = w1405 & ~w1443;
assign w1445 = ~w1405 & w1443;
assign w1446 = ~w1444 & ~w1445;
assign w1447 = w1404 & w1446;
assign w1448 = ~w1404 & ~w1446;
assign w1449 = ~w1447 & ~w1448;
assign w1450 = (~w1253 & ~w1255) | (~w1253 & w16982) | (~w1255 & w16982);
assign w1451 = ~w1449 & w1450;
assign w1452 = w1449 & ~w1450;
assign w1453 = ~w1451 & ~w1452;
assign w1454 = w1403 & w1453;
assign w1455 = ~w1403 & ~w1453;
assign w1456 = ~w1454 & ~w1455;
assign w1457 = w1402 & w1456;
assign w1458 = ~w1402 & ~w1456;
assign w1459 = ~w1457 & ~w1458;
assign w1460 = w1194 & w16983;
assign w1461 = (~w1460 & ~w1259) | (~w1460 & w16984) | (~w1259 & w16984);
assign w1462 = w1459 & ~w1461;
assign w1463 = ~w1459 & w1461;
assign w1464 = ~w1462 & ~w1463;
assign w1465 = ~pi129 & w1265;
assign w1466 = pi314 & ~w463;
assign w1467 = (w1466 & w1265) | (w1466 & w16985) | (w1265 & w16985);
assign w1468 = ~w1465 & w1467;
assign w1469 = w1464 & ~w1468;
assign w1470 = ~w1464 & w1468;
assign w1471 = ~w1469 & ~w1470;
assign w1472 = w1401 & ~w1471;
assign w1473 = ~w1401 & w1471;
assign w1474 = ~w1472 & ~w1473;
assign w1475 = (~w1382 & ~w1384) | (~w1382 & w16986) | (~w1384 & w16986);
assign w1476 = pi330 & w456;
assign w1477 = ~w465 & w16987;
assign w1478 = (~w1477 & ~w1377) | (~w1477 & w16988) | (~w1377 & w16988);
assign w1479 = w1377 & w16989;
assign w1480 = ~w1478 & ~w1479;
assign w1481 = (pi328 & ~w536) | (pi328 & w16990) | (~w536 & w16990);
assign w1482 = pi327 & ~w615;
assign w1483 = w1362 & w1363;
assign w1484 = ~w1362 & ~w1363;
assign w1485 = ~w1483 & ~w1484;
assign w1486 = (~w1483 & ~w1485) | (~w1483 & w16991) | (~w1485 & w16991);
assign w1487 = w1482 & ~w1486;
assign w1488 = ~w1482 & w1486;
assign w1489 = ~w1487 & ~w1488;
assign w1490 = pi326 & ~w793;
assign w1491 = (~w1357 & ~w1358) | (~w1357 & w16992) | (~w1358 & w16992);
assign w1492 = w1490 & ~w1491;
assign w1493 = ~w1490 & w1491;
assign w1494 = ~w1492 & ~w1493;
assign w1495 = (~w1277 & w1352) | (~w1277 & w16993) | (w1352 & w16993);
assign w1496 = pi325 & ~w955;
assign w1497 = pi324 & w1101;
assign w1498 = (~w1347 & ~w1348) | (~w1347 & w16994) | (~w1348 & w16994);
assign w1499 = (~w1282 & ~w1078) | (~w1282 & w16995) | (~w1078 & w16995);
assign w1500 = w1078 & w16996;
assign w1501 = ~w1499 & ~w1500;
assign w1502 = w1327 & w1501;
assign w1503 = ~w1327 & ~w1501;
assign w1504 = ~w1502 & ~w1503;
assign w1505 = w1280 & w1504;
assign w1506 = ~w1280 & ~w1504;
assign w1507 = ~w1505 & ~w1506;
assign w1508 = w1281 & w1507;
assign w1509 = ~w1281 & ~w1507;
assign w1510 = ~w1508 & ~w1509;
assign w1511 = pi136 & pi258;
assign w1512 = pi135 & pi259;
assign w1513 = (~w1512 & ~w1504) | (~w1512 & w15809) | (~w1504 & w15809);
assign w1514 = w1504 & w15810;
assign w1515 = ~w1513 & ~w1514;
assign w1516 = (~w1500 & ~w1327) | (~w1500 & w15811) | (~w1327 & w15811);
assign w1517 = pi134 & pi260;
assign w1518 = pi133 & pi261;
assign w1519 = (w1318 & w1288) | (w1318 & w15812) | (w1288 & w15812);
assign w1520 = ~w1316 & ~w1519;
assign w1521 = ~w1056 & w15813;
assign w1522 = ~w1308 & ~w1521;
assign w1523 = pi132 & pi262;
assign w1524 = ~w1038 & ~w1296;
assign w1525 = pi130 & pi264;
assign w1526 = pi129 & pi265;
assign w1527 = pi128 & pi266;
assign w1528 = ~w1526 & ~w1527;
assign w1529 = w1526 & w1527;
assign w1530 = ~w1528 & ~w1529;
assign w1531 = w1525 & ~w1530;
assign w1532 = ~w1525 & w1530;
assign w1533 = ~w1531 & ~w1532;
assign w1534 = w17634 & w1533;
assign w1535 = ~w17634 & ~w1533;
assign w1536 = ~w1534 & ~w1535;
assign w1537 = pi131 & pi263;
assign w1538 = ~w1536 & w1537;
assign w1539 = w1536 & ~w1537;
assign w1540 = ~w1538 & ~w1539;
assign w1541 = ~w1293 & w17631;
assign w1542 = ~w1540 & w1541;
assign w1543 = ~pi131 & ~w1536;
assign w1544 = w1543 & w17632;
assign w1545 = ~pi263 & ~w1536;
assign w1546 = (w1291 & w16348) | (w1291 & w16349) | (w16348 & w16349);
assign w1547 = ~w1291 & w15816;
assign w1548 = ~pi131 & w1536;
assign w1549 = ~w1538 & ~w1548;
assign w1550 = w1547 & ~w1549;
assign w1551 = (w1291 & w16997) | (w1291 & w16998) | (w16997 & w16998);
assign w1552 = (w1291 & w16350) | (w1291 & w16351) | (w16350 & w16351);
assign w1553 = pi131 & ~w1552;
assign w1554 = w1551 & w1553;
assign w1555 = ~w1546 & ~w1550;
assign w1556 = ~w1542 & w1555;
assign w1557 = w1556 & w16352;
assign w1558 = w1523 & w1557;
assign w1559 = w1522 & w1558;
assign w1560 = w1523 & ~w1557;
assign w1561 = ~w1522 & w1560;
assign w1562 = ~w1559 & ~w1561;
assign w1563 = ~w1521 & w16999;
assign w1564 = (~w1523 & w1522) | (~w1523 & w16110) | (w1522 & w16110);
assign w1565 = ~w1563 & w1564;
assign w1566 = w1562 & ~w1565;
assign w1567 = w1520 & ~w1566;
assign w1568 = ~w1520 & w1566;
assign w1569 = ~w1567 & ~w1568;
assign w1570 = w1518 & w1569;
assign w1571 = ~w1518 & ~w1569;
assign w1572 = ~w1570 & ~w1571;
assign w1573 = (w1284 & ~w1321) | (w1284 & w15817) | (~w1321 & w15817);
assign w1574 = ~w1323 & ~w1573;
assign w1575 = w1572 & ~w1574;
assign w1576 = ~w1572 & w1574;
assign w1577 = ~w1575 & ~w1576;
assign w1578 = w1517 & ~w1577;
assign w1579 = ~w1517 & w1577;
assign w1580 = ~w1578 & ~w1579;
assign w1581 = w1516 & w1580;
assign w1582 = ~w1516 & ~w1580;
assign w1583 = ~w1581 & ~w1582;
assign w1584 = w1515 & ~w1583;
assign w1585 = ~w1515 & w1583;
assign w1586 = ~w1584 & ~w1585;
assign w1587 = w1511 & w1586;
assign w1588 = ~w1511 & ~w1586;
assign w1589 = ~w1587 & ~w1588;
assign w1590 = w1082 & ~w1510;
assign w1591 = (~w1507 & w1510) | (~w1507 & w17000) | (w1510 & w17000);
assign w1592 = w1589 & ~w1591;
assign w1593 = (w1101 & w17001) | (w1101 & w17002) | (w17001 & w17002);
assign w1594 = w1507 & ~w1593;
assign w1595 = (~w1594 & ~w1589) | (~w1594 & w16353) | (~w1589 & w16353);
assign w1596 = ~w1510 & w1595;
assign w1597 = (w1082 & ~w1589) | (w1082 & w16547) | (~w1589 & w16547);
assign w1598 = ~w1596 & w1597;
assign w1599 = ~w1508 & w1589;
assign w1600 = (~w1082 & w1589) | (~w1082 & w16548) | (w1589 & w16548);
assign w1601 = ~w1599 & w1600;
assign w1602 = ~w1598 & ~w1601;
assign w1603 = ~w1082 & w1510;
assign w1604 = (pi323 & w1510) | (pi323 & w17003) | (w1510 & w17003);
assign w1605 = ~w1603 & w1604;
assign w1606 = (~w1605 & ~w1602) | (~w1605 & w17004) | (~w1602 & w17004);
assign w1607 = w1602 & w17005;
assign w1608 = ~w1606 & ~w1607;
assign w1609 = (~w1341 & ~w1339) | (~w1341 & w17006) | (~w1339 & w17006);
assign w1610 = ~w1608 & w1609;
assign w1611 = w1608 & ~w1609;
assign w1612 = ~w1610 & ~w1611;
assign w1613 = w1498 & ~w1612;
assign w1614 = ~w1498 & w1612;
assign w1615 = ~w1613 & ~w1614;
assign w1616 = w1497 & ~w1615;
assign w1617 = ~w1497 & w1615;
assign w1618 = ~w1616 & ~w1617;
assign w1619 = w1496 & ~w1618;
assign w1620 = ~w1496 & w1618;
assign w1621 = ~w1619 & ~w1620;
assign w1622 = w1495 & w1621;
assign w1623 = ~w1495 & ~w1621;
assign w1624 = ~w1622 & ~w1623;
assign w1625 = ~w1494 & w1624;
assign w1626 = w1494 & ~w1624;
assign w1627 = ~w1625 & ~w1626;
assign w1628 = w1489 & ~w1627;
assign w1629 = ~w1489 & w1627;
assign w1630 = ~w1628 & ~w1629;
assign w1631 = ~w1368 & ~w1485;
assign w1632 = (~w1271 & ~w1485) | (~w1271 & w17007) | (~w1485 & w17007);
assign w1633 = ~w1631 & w1632;
assign w1634 = ~w1272 & ~w1633;
assign w1635 = ~w1630 & w1634;
assign w1636 = w1630 & ~w1634;
assign w1637 = ~w1635 & ~w1636;
assign w1638 = ~w1481 & w1637;
assign w1639 = w1481 & ~w1637;
assign w1640 = ~w1638 & ~w1639;
assign w1641 = w1480 & ~w1640;
assign w1642 = ~w1480 & w1640;
assign w1643 = ~w1641 & ~w1642;
assign w1644 = w1476 & w1643;
assign w1645 = ~w1476 & ~w1643;
assign w1646 = ~w1644 & ~w1645;
assign w1647 = ~w1475 & ~w1646;
assign w1648 = w1475 & w1646;
assign w1649 = ~w1647 & ~w1648;
assign w1650 = pi266 & w1649;
assign w1651 = ~pi266 & ~w1649;
assign w1652 = ~w1650 & ~w1651;
assign w1653 = ~w1389 & ~w1392;
assign w1654 = w1652 & ~w1653;
assign w1655 = ~w1652 & w1653;
assign w1656 = ~w1654 & ~w1655;
assign w1657 = ~w1474 & w1656;
assign w1658 = (~w135 & w1656) | (~w135 & w17008) | (w1656 & w17008);
assign w1659 = ~w1657 & w1658;
assign w1660 = (pi161 & ~w135) | (pi161 & w17009) | (~w135 & w17009);
assign w1661 = ~w1659 & w1660;
assign w1662 = ~pi160 & ~w1400;
assign w1663 = ~w1661 & w1662;
assign w1664 = ~pi073 & ~pi161;
assign w1665 = pi128 & pi312;
assign w1666 = (w1467 & w1464) | (w1467 & w17010) | (w1464 & w17010);
assign w1667 = pi314 & ~w653;
assign w1668 = pi315 & w709;
assign w1669 = pi316 & w698;
assign w1670 = pi317 & w855;
assign w1671 = (~w1445 & ~w1446) | (~w1445 & w17011) | (~w1446 & w17011);
assign w1672 = pi318 & w1159;
assign w1673 = pi319 & w1220;
assign w1674 = pi136 & pi137;
assign w1675 = ~pi137 & w1410;
assign w1676 = pi135 & pi137;
assign w1677 = (~w1676 & w1153) | (~w1676 & w17012) | (w1153 & w17012);
assign w1678 = pi134 & ~w1677;
assign w1679 = ~w1674 & w17633;
assign w1680 = pi134 & pi136;
assign w1681 = ~pi137 & w1680;
assign w1682 = (w849 & w17017) | (w849 & w17018) | (w17017 & w17018);
assign w1683 = pi133 & ~w1682;
assign w1684 = ~pi136 & ~pi137;
assign w1685 = pi137 & w1409;
assign w1686 = (~w1685 & ~w849) | (~w1685 & w17020) | (~w849 & w17020);
assign w1687 = ~pi134 & ~w1686;
assign w1688 = ~pi134 & w1684;
assign w1689 = (~w1688 & ~w849) | (~w1688 & w17022) | (~w849 & w17022);
assign w1690 = ~pi133 & ~w1689;
assign w1691 = ~w1687 & ~w1690;
assign w1692 = ~w1683 & w1691;
assign w1693 = ~w1679 & w1692;
assign w1694 = w1692 & w17023;
assign w1695 = (w1421 & w1422) | (w1421 & w17024) | (w1422 & w17024);
assign w1696 = (~w1420 & ~w1422) | (~w1420 & w17025) | (~w1422 & w17025);
assign w1697 = ~w1694 & ~w1695;
assign w1698 = ~w1696 & ~w1697;
assign w1699 = ~w1697 & w17026;
assign w1700 = (w1694 & ~w1699) | (w1694 & w17027) | (~w1699 & w17027);
assign w1701 = ~w1698 & w17026;
assign w1702 = ~w1700 & ~w1701;
assign w1703 = w1407 & ~w1430;
assign w1704 = ~w1703 & w17028;
assign w1705 = (~w1702 & w1703) | (~w1702 & w17029) | (w1703 & w17029);
assign w1706 = ~w1704 & ~w1705;
assign w1707 = w1673 & ~w1706;
assign w1708 = ~w1673 & w1706;
assign w1709 = ~w1707 & ~w1708;
assign w1710 = (w1406 & ~w1437) | (w1406 & w17030) | (~w1437 & w17030);
assign w1711 = ~w1439 & ~w1710;
assign w1712 = w1709 & w1711;
assign w1713 = ~w1709 & ~w1711;
assign w1714 = ~w1712 & ~w1713;
assign w1715 = w1672 & w1714;
assign w1716 = ~w1672 & ~w1714;
assign w1717 = ~w1715 & ~w1716;
assign w1718 = ~w1671 & w1717;
assign w1719 = w1671 & ~w1717;
assign w1720 = ~w1718 & ~w1719;
assign w1721 = w1670 & ~w1720;
assign w1722 = ~w1670 & w1720;
assign w1723 = ~w1721 & ~w1722;
assign w1724 = (~w1452 & ~w1453) | (~w1452 & w17031) | (~w1453 & w17031);
assign w1725 = w1723 & w1724;
assign w1726 = ~w1723 & ~w1724;
assign w1727 = ~w1725 & ~w1726;
assign w1728 = w1669 & w1727;
assign w1729 = ~w1669 & ~w1727;
assign w1730 = ~w1728 & ~w1729;
assign w1731 = w1668 & w1730;
assign w1732 = ~w1668 & ~w1730;
assign w1733 = ~w1731 & ~w1732;
assign w1734 = (~w1457 & ~w1459) | (~w1457 & w17032) | (~w1459 & w17032);
assign w1735 = w1733 & ~w1734;
assign w1736 = ~w1733 & w1734;
assign w1737 = ~w1735 & ~w1736;
assign w1738 = ~w1667 & ~w1737;
assign w1739 = w1667 & w1737;
assign w1740 = ~w1738 & ~w1739;
assign w1741 = w1666 & w1740;
assign w1742 = ~w1666 & ~w1740;
assign w1743 = ~w1741 & ~w1742;
assign w1744 = (~pi129 & ~w1471) | (~pi129 & w463) | (~w1471 & w463);
assign w1745 = (pi313 & ~w1471) | (pi313 & w17033) | (~w1471 & w17033);
assign w1746 = ~w1744 & w1745;
assign w1747 = ~w1743 & ~w1746;
assign w1748 = w1743 & w1746;
assign w1749 = ~w1747 & ~w1748;
assign w1750 = w1665 & w1749;
assign w1751 = ~w1665 & ~w1749;
assign w1752 = ~w1750 & ~w1751;
assign w1753 = pi331 & w456;
assign w1754 = pi328 & ~w615;
assign w1755 = (~w1635 & ~w1637) | (~w1635 & w17034) | (~w1637 & w17034);
assign w1756 = w1754 & w1755;
assign w1757 = ~w1754 & ~w1755;
assign w1758 = ~w1756 & ~w1757;
assign w1759 = pi327 & ~w793;
assign w1760 = (~w1487 & w1627) | (~w1487 & w17035) | (w1627 & w17035);
assign w1761 = ~w1759 & w1760;
assign w1762 = w1759 & ~w1760;
assign w1763 = ~w1761 & ~w1762;
assign w1764 = (~w1619 & ~w1621) | (~w1619 & w17036) | (~w1621 & w17036);
assign w1765 = pi325 & w1101;
assign w1766 = pi324 & w1339;
assign w1767 = (~w1613 & ~w1615) | (~w1613 & w17037) | (~w1615 & w17037);
assign w1768 = ~w1766 & ~w1767;
assign w1769 = w1766 & w1767;
assign w1770 = ~w1768 & ~w1769;
assign w1771 = pi323 & w1602;
assign w1772 = pi137 & pi258;
assign w1773 = pi136 & pi259;
assign w1774 = (~w1773 & ~w1586) | (~w1773 & w16111) | (~w1586 & w16111);
assign w1775 = w1586 & w16112;
assign w1776 = ~w1774 & ~w1775;
assign w1777 = (~w1514 & w1583) | (~w1514 & w16113) | (w1583 & w16113);
assign w1778 = ~w1571 & w1574;
assign w1779 = (~w1570 & ~w1574) | (~w1570 & w16114) | (~w1574 & w16114);
assign w1780 = pi133 & pi262;
assign w1781 = ~w1316 & w1562;
assign w1782 = (~w1565 & ~w1781) | (~w1565 & w15818) | (~w1781 & w15818);
assign w1783 = pi132 & pi263;
assign w1784 = pi131 & pi264;
assign w1785 = ~w1530 & w17634;
assign w1786 = (w1035 & w16354) | (w1035 & w16355) | (w16354 & w16355);
assign w1787 = ~w1785 & ~w1786;
assign w1788 = ~w1525 & ~w1787;
assign w1789 = w1525 & w1787;
assign w1790 = (w1292 & w16115) | (w1292 & w16116) | (w16115 & w16116);
assign w1791 = pi130 & pi265;
assign w1792 = pi129 & pi266;
assign w1793 = pi128 & pi267;
assign w1794 = ~w1792 & ~w1793;
assign w1795 = w1792 & w1793;
assign w1796 = ~w1794 & ~w1795;
assign w1797 = ~w1786 & w16549;
assign w1798 = (w1796 & w1786) | (w1796 & w16550) | (w1786 & w16550);
assign w1799 = ~w1797 & ~w1798;
assign w1800 = w1791 & w1799;
assign w1801 = ~w1791 & ~w1799;
assign w1802 = ~w1800 & ~w1801;
assign w1803 = ~w1790 & w16356;
assign w1804 = (~w1802 & w1790) | (~w1802 & w16357) | (w1790 & w16357);
assign w1805 = ~w1803 & ~w1804;
assign w1806 = ~w1784 & ~w1805;
assign w1807 = w1784 & w1805;
assign w1808 = ~w1806 & ~w1807;
assign w1809 = w1543 & w17635;
assign w1810 = ~w1545 & ~w1552;
assign w1811 = ~w1546 & ~w1810;
assign w1812 = (~w1292 & w16117) | (~w1292 & w16118) | (w16117 & w16118);
assign w1813 = ~w1308 & w15819;
assign w1814 = ~w1811 & w1813;
assign w1815 = ~w1536 & w17635;
assign w1816 = w1537 & ~w1551;
assign w1817 = ~w1815 & w1816;
assign w1818 = (~w1817 & w1521) | (~w1817 & w16119) | (w1521 & w16119);
assign w1819 = w1808 & ~w1818;
assign w1820 = ~w1808 & w1818;
assign w1821 = ~w1819 & ~w1820;
assign w1822 = w1783 & ~w1821;
assign w1823 = ~w1783 & w1821;
assign w1824 = ~w1822 & ~w1823;
assign w1825 = w1782 & ~w1824;
assign w1826 = ~w1782 & w1824;
assign w1827 = ~w1825 & ~w1826;
assign w1828 = ~w1780 & ~w1827;
assign w1829 = w1780 & w1827;
assign w1830 = ~w1828 & ~w1829;
assign w1831 = pi134 & pi261;
assign w1832 = w1830 & w1831;
assign w1833 = w1779 & w1832;
assign w1834 = ~w1830 & w1831;
assign w1835 = ~w1779 & w1834;
assign w1836 = ~w1833 & ~w1835;
assign w1837 = w1779 & w1830;
assign w1838 = (~w1831 & w1779) | (~w1831 & w15820) | (w1779 & w15820);
assign w1839 = ~w1837 & w1838;
assign w1840 = w1836 & ~w1839;
assign w1841 = ~w1516 & ~w1577;
assign w1842 = (w1517 & ~w1516) | (w1517 & w1578) | (~w1516 & w1578);
assign w1843 = ~w1841 & ~w1842;
assign w1844 = ~w1840 & w1843;
assign w1845 = w1840 & ~w1843;
assign w1846 = ~w1844 & ~w1845;
assign w1847 = w1777 & ~w1846;
assign w1848 = ~w1777 & w1846;
assign w1849 = ~w1847 & ~w1848;
assign w1850 = pi135 & pi260;
assign w1851 = ~w1849 & ~w1850;
assign w1852 = w1849 & w1850;
assign w1853 = ~w1851 & ~w1852;
assign w1854 = w1776 & w1853;
assign w1855 = ~w1776 & ~w1853;
assign w1856 = ~w1854 & ~w1855;
assign w1857 = w1772 & w1856;
assign w1858 = ~w1772 & ~w1856;
assign w1859 = ~w1857 & ~w1858;
assign w1860 = w1595 & ~w1859;
assign w1861 = ~w1595 & w1859;
assign w1862 = ~w1860 & ~w1861;
assign w1863 = w1589 & ~w1862;
assign w1864 = ~w1589 & w1862;
assign w1865 = ~w1863 & ~w1864;
assign w1866 = (~w1771 & w1865) | (~w1771 & w16551) | (w1865 & w16551);
assign w1867 = ~w1865 & w16552;
assign w1868 = ~w1866 & ~w1867;
assign w1869 = (~w1607 & ~w1608) | (~w1607 & w17038) | (~w1608 & w17038);
assign w1870 = w1868 & ~w1869;
assign w1871 = ~w1868 & w1869;
assign w1872 = ~w1870 & ~w1871;
assign w1873 = w1770 & w1872;
assign w1874 = ~w1770 & ~w1872;
assign w1875 = ~w1873 & ~w1874;
assign w1876 = ~w1765 & ~w1875;
assign w1877 = w1765 & w1875;
assign w1878 = ~w1876 & ~w1877;
assign w1879 = w1764 & w1878;
assign w1880 = ~w1764 & ~w1878;
assign w1881 = ~w1879 & ~w1880;
assign w1882 = pi326 & ~w955;
assign w1883 = (~w1493 & w1624) | (~w1493 & w17039) | (w1624 & w17039);
assign w1884 = w1882 & w1883;
assign w1885 = ~w1882 & ~w1883;
assign w1886 = ~w1884 & ~w1885;
assign w1887 = w1881 & w1886;
assign w1888 = ~w1881 & ~w1886;
assign w1889 = ~w1887 & ~w1888;
assign w1890 = ~w1763 & w1889;
assign w1891 = w1763 & ~w1889;
assign w1892 = ~w1890 & ~w1891;
assign w1893 = w1758 & w1892;
assign w1894 = ~w1758 & ~w1892;
assign w1895 = ~w1893 & ~w1894;
assign w1896 = (pi329 & ~w536) | (pi329 & w17040) | (~w536 & w17040);
assign w1897 = (w1640 & w17042) | (w1640 & w17043) | (w17042 & w17043);
assign w1898 = w1896 & w17636;
assign w1899 = ~w1897 & ~w1898;
assign w1900 = w1895 & ~w1899;
assign w1901 = ~w1895 & w1899;
assign w1902 = ~w1900 & ~w1901;
assign w1903 = ~w465 & w17044;
assign w1904 = (~w1903 & ~w1643) | (~w1903 & w17045) | (~w1643 & w17045);
assign w1905 = w971 & w1643;
assign w1906 = ~w1904 & ~w1905;
assign w1907 = w1902 & w1906;
assign w1908 = ~w1902 & ~w1906;
assign w1909 = ~w1907 & ~w1908;
assign w1910 = w1753 & ~w1909;
assign w1911 = ~w1753 & w1909;
assign w1912 = ~w1910 & ~w1911;
assign w1913 = (~w1647 & ~w1649) | (~w1647 & w17046) | (~w1649 & w17046);
assign w1914 = ~w1912 & ~w1913;
assign w1915 = w1912 & w1913;
assign w1916 = ~w1914 & ~w1915;
assign w1917 = pi267 & w1916;
assign w1918 = ~pi267 & ~w1916;
assign w1919 = ~w1917 & ~w1918;
assign w1920 = (~w1654 & ~w1656) | (~w1654 & w17047) | (~w1656 & w17047);
assign w1921 = w1919 & ~w1920;
assign w1922 = ~w1919 & w1920;
assign w1923 = ~w1921 & ~w1922;
assign w1924 = w1752 & ~w1923;
assign w1925 = (~w135 & ~w1923) | (~w135 & w17048) | (~w1923 & w17048);
assign w1926 = ~w1924 & w1925;
assign w1927 = (pi161 & ~w135) | (pi161 & w17049) | (~w135 & w17049);
assign w1928 = ~w1926 & w1927;
assign w1929 = ~pi160 & ~w1664;
assign w1930 = ~w1928 & w1929;
assign w1931 = ~pi074 & ~pi161;
assign w1932 = pi128 & pi311;
assign w1933 = pi312 & w464;
assign w1934 = pi313 & ~w653;
assign w1935 = pi315 & w698;
assign w1936 = pi316 & w855;
assign w1937 = pi318 & w1220;
assign w1938 = w1419 & w17050;
assign w1939 = (w1703 & w17051) | (w1703 & w17052) | (w17051 & w17052);
assign w1940 = ~w1705 & ~w1939;
assign w1941 = ~w1938 & w1940;
assign w1942 = w1938 & ~w1940;
assign w1943 = ~w1941 & ~w1942;
assign w1944 = ~pi135 & ~pi137;
assign w1945 = pi136 & ~w1944;
assign w1946 = pi135 & w17637;
assign w1947 = (pi133 & w1946) | (pi133 & w17053) | (w1946 & w17053);
assign w1948 = ~w1678 & w17054;
assign w1949 = ~pi138 & w1948;
assign w1950 = pi138 & ~w1948;
assign w1951 = ~w1949 & ~w1950;
assign w1952 = pi137 & w1951;
assign w1953 = ~pi137 & ~w1951;
assign w1954 = ~w1952 & ~w1953;
assign w1955 = pi321 & w1954;
assign w1956 = ~w1693 & ~w1699;
assign w1957 = (w1693 & w1698) | (w1693 & w17055) | (w1698 & w17055);
assign w1958 = ~w1956 & ~w1957;
assign w1959 = w1955 & ~w1958;
assign w1960 = ~w1955 & w1958;
assign w1961 = ~w1959 & ~w1960;
assign w1962 = w1943 & ~w1961;
assign w1963 = ~w1943 & w1961;
assign w1964 = ~w1962 & ~w1963;
assign w1965 = (w1672 & ~w1711) | (w1672 & w17056) | (~w1711 & w17056);
assign w1966 = ~w1713 & ~w1965;
assign w1967 = ~w1964 & w1966;
assign w1968 = w1964 & ~w1966;
assign w1969 = ~w1967 & ~w1968;
assign w1970 = w1937 & ~w1969;
assign w1971 = ~w1937 & w1969;
assign w1972 = ~w1970 & ~w1971;
assign w1973 = w1719 & w1972;
assign w1974 = ~w1722 & ~w1973;
assign w1975 = ~w1719 & ~w1972;
assign w1976 = (~w1159 & w1719) | (~w1159 & w17057) | (w1719 & w17057);
assign w1977 = pi317 & w1159;
assign w1978 = ~w1972 & w1977;
assign w1979 = ~w1718 & ~w1978;
assign w1980 = (~w1670 & ~w1972) | (~w1670 & w17058) | (~w1972 & w17058);
assign w1981 = w1979 & w1980;
assign w1982 = (~w1981 & ~w1974) | (~w1981 & w15822) | (~w1974 & w15822);
assign w1983 = w1718 & ~w1972;
assign w1984 = ~w1973 & ~w1983;
assign w1985 = w1977 & ~w1984;
assign w1986 = (w1213 & w1671) | (w1213 & w17059) | (w1671 & w17059);
assign w1987 = w1975 & w1986;
assign w1988 = ~w1985 & ~w1987;
assign w1989 = w1982 & w1988;
assign w1990 = w1726 & ~w1989;
assign w1991 = ~w1726 & w1989;
assign w1992 = ~w1728 & w1991;
assign w1993 = (w1936 & w1992) | (w1936 & w17060) | (w1992 & w17060);
assign w1994 = w698 & w1727;
assign w1995 = w1727 & w15823;
assign w1996 = ~w1669 & ~w1936;
assign w1997 = ~w1726 & w1996;
assign w1998 = (~w1989 & w1995) | (~w1989 & w17061) | (w1995 & w17061);
assign w1999 = (~w855 & w1989) | (~w855 & w17062) | (w1989 & w17062);
assign w2000 = ~w1992 & w1999;
assign w2001 = ~w1998 & ~w2000;
assign w2002 = ~w1993 & w2001;
assign w2003 = (~w1731 & ~w1733) | (~w1731 & w15824) | (~w1733 & w15824);
assign w2004 = w2002 & w2003;
assign w2005 = ~w2002 & ~w2003;
assign w2006 = ~w2004 & ~w2005;
assign w2007 = w1935 & ~w2006;
assign w2008 = ~w1935 & w2006;
assign w2009 = ~w2007 & ~w2008;
assign w2010 = (~w1739 & ~w1740) | (~w1739 & w17063) | (~w1740 & w17063);
assign w2011 = w2009 & w2010;
assign w2012 = ~w2009 & ~w2010;
assign w2013 = ~w2011 & ~w2012;
assign w2014 = pi314 & w709;
assign w2015 = w2013 & w2014;
assign w2016 = ~w2013 & ~w2014;
assign w2017 = ~w2015 & ~w2016;
assign w2018 = ~w1471 & w17064;
assign w2019 = (~w2018 & ~w1743) | (~w2018 & w17065) | (~w1743 & w17065);
assign w2020 = w2017 & ~w2019;
assign w2021 = ~w2017 & w2019;
assign w2022 = ~w2020 & ~w2021;
assign w2023 = ~w1934 & w2022;
assign w2024 = w1934 & ~w2022;
assign w2025 = ~w2023 & ~w2024;
assign w2026 = w1933 & ~w2025;
assign w2027 = ~w1933 & w2025;
assign w2028 = ~w2026 & ~w2027;
assign w2029 = w1750 & w2028;
assign w2030 = ~w1750 & ~w2028;
assign w2031 = ~w2029 & ~w2030;
assign w2032 = w1932 & w2031;
assign w2033 = ~w1932 & ~w2031;
assign w2034 = ~w2032 & ~w2033;
assign w2035 = (~w1914 & ~w1916) | (~w1914 & w17066) | (~w1916 & w17066);
assign w2036 = pi332 & w456;
assign w2037 = ~w465 & w17067;
assign w2038 = (~w2037 & w1909) | (~w2037 & w17068) | (w1909 & w17068);
assign w2039 = ~w1909 & w17069;
assign w2040 = ~w2038 & ~w2039;
assign w2041 = (~w1897 & w1895) | (~w1897 & w17070) | (w1895 & w17070);
assign w2042 = pi329 & ~w615;
assign w2043 = pi327 & ~w955;
assign w2044 = (~w1762 & w1889) | (~w1762 & w17071) | (w1889 & w17071);
assign w2045 = ~w2043 & w2044;
assign w2046 = w2043 & ~w2044;
assign w2047 = ~w2045 & ~w2046;
assign w2048 = pi326 & w1101;
assign w2049 = (~w1876 & ~w1878) | (~w1876 & w17072) | (~w1878 & w17072);
assign w2050 = pi325 & w1339;
assign w2051 = pi324 & w1602;
assign w2052 = (~w1769 & ~w1872) | (~w1769 & w17073) | (~w1872 & w17073);
assign w2053 = ~w2051 & w2052;
assign w2054 = w2051 & ~w2052;
assign w2055 = ~w2053 & ~w2054;
assign w2056 = pi323 & ~w1865;
assign w2057 = pi138 & pi258;
assign w2058 = pi137 & pi259;
assign w2059 = (~w2058 & ~w1856) | (~w2058 & w15825) | (~w1856 & w15825);
assign w2060 = w1856 & w15826;
assign w2061 = ~w2059 & ~w2060;
assign w2062 = pi135 & pi261;
assign w2063 = w1836 & ~w1841;
assign w2064 = (~w1839 & ~w2063) | (~w1839 & w15827) | (~w2063 & w15827);
assign w2065 = pi133 & pi263;
assign w2066 = (~w1783 & ~w1782) | (~w1783 & w16120) | (~w1782 & w16120);
assign w2067 = (~w15818 & w16121) | (~w15818 & w16122) | (w16121 & w16122);
assign w2068 = pi132 & pi264;
assign w2069 = (~w1799 & w1790) | (~w1799 & w15828) | (w1790 & w15828);
assign w2070 = (~w1791 & w1790) | (~w1791 & w16358) | (w1790 & w16358);
assign w2071 = ~w2069 & ~w2070;
assign w2072 = (~w1795 & w15830) | (~w1795 & w17638) | (w15830 & w17638);
assign w2073 = pi129 & pi267;
assign w2074 = pi128 & pi268;
assign w2075 = ~w2073 & ~w2074;
assign w2076 = pi129 & pi268;
assign w2077 = w1793 & w2076;
assign w2078 = ~w2075 & ~w2077;
assign w2079 = pi130 & pi266;
assign w2080 = w2078 & w2079;
assign w2081 = ~w2078 & ~w2079;
assign w2082 = ~w2080 & ~w2081;
assign w2083 = w2082 & w17639;
assign w2084 = ~w2078 & w17074;
assign w2085 = (w2084 & w1786) | (w2084 & w17075) | (w1786 & w17075);
assign w2086 = ~w1792 & ~w2078;
assign w2087 = ~w2082 & ~w2086;
assign w2088 = ~w2072 & w2087;
assign w2089 = ~w2083 & ~w2085;
assign w2090 = ~w2088 & w2089;
assign w2091 = (~w1790 & w16359) | (~w1790 & w16360) | (w16359 & w16360);
assign w2092 = (w1790 & w17076) | (w1790 & w17077) | (w17076 & w17077);
assign w2093 = (w2092 & w2071) | (w2092 & w17078) | (w2071 & w17078);
assign w2094 = pi131 & pi265;
assign w2095 = w2090 & w2094;
assign w2096 = ~w2090 & ~w2094;
assign w2097 = ~w2095 & ~w2096;
assign w2098 = (w1790 & w17079) | (w1790 & w17080) | (w17079 & w17080);
assign w2099 = (w1790 & w16555) | (w1790 & w16556) | (w16555 & w16556);
assign w2100 = ~pi265 & w2090;
assign w2101 = ~w1790 & w16557;
assign w2102 = ~w1790 & w17081;
assign w2103 = w700 & w2091;
assign w2104 = ~w2102 & w2103;
assign w2105 = ~w2099 & ~w2101;
assign w2106 = ~w2098 & w2105;
assign w2107 = ~w2104 & w2106;
assign w2108 = ~w2093 & w2107;
assign w2109 = (~w1807 & w1818) | (~w1807 & w16361) | (w1818 & w16361);
assign w2110 = w2108 & ~w2109;
assign w2111 = ~w2108 & w2109;
assign w2112 = ~w2110 & ~w2111;
assign w2113 = w2068 & ~w2112;
assign w2114 = ~w2068 & w2112;
assign w2115 = ~w2113 & ~w2114;
assign w2116 = ~w2066 & w16362;
assign w2117 = (~w2115 & w2066) | (~w2115 & w16363) | (w2066 & w16363);
assign w2118 = ~w2116 & ~w2117;
assign w2119 = ~w2065 & ~w2118;
assign w2120 = w2065 & w2118;
assign w2121 = ~w2119 & ~w2120;
assign w2122 = ~w1570 & ~w1829;
assign w2123 = ~w1778 & w2122;
assign w2124 = (~w1828 & ~w2122) | (~w1828 & w16364) | (~w2122 & w16364);
assign w2125 = pi134 & pi262;
assign w2126 = (w2125 & w2123) | (w2125 & w15831) | (w2123 & w15831);
assign w2127 = ~w2123 & w15832;
assign w2128 = ~w2126 & ~w2127;
assign w2129 = w2121 & w2128;
assign w2130 = ~w2121 & ~w2128;
assign w2131 = ~w2129 & ~w2130;
assign w2132 = w2064 & w2131;
assign w2133 = ~w2064 & ~w2131;
assign w2134 = ~w2132 & ~w2133;
assign w2135 = ~w2062 & w2134;
assign w2136 = w2062 & ~w2134;
assign w2137 = ~w2135 & ~w2136;
assign w2138 = (~w1850 & w1777) | (~w1850 & w15833) | (w1777 & w15833);
assign w2139 = ~w1847 & ~w2138;
assign w2140 = w2137 & ~w2139;
assign w2141 = ~w2137 & w2139;
assign w2142 = ~w2140 & ~w2141;
assign w2143 = pi136 & pi260;
assign w2144 = ~w1850 & ~w2143;
assign w2145 = (w1586 & w16365) | (w1586 & w16366) | (w16365 & w16366);
assign w2146 = (w2143 & w15834) | (w2143 & ~w1587) | (w15834 & ~w1587);
assign w2147 = pi135 & w17640;
assign w2148 = ~w2145 & ~w2147;
assign w2149 = w1849 & ~w2148;
assign w2150 = w1586 & w16367;
assign w2151 = w1851 & w2146;
assign w2152 = w2143 & w1774;
assign w2153 = ~w2150 & ~w2152;
assign w2154 = ~w2151 & w2153;
assign w2155 = ~w2149 & w2154;
assign w2156 = ~w2142 & ~w2155;
assign w2157 = w2142 & w2155;
assign w2158 = ~w2156 & ~w2157;
assign w2159 = w2061 & w2158;
assign w2160 = ~w2061 & ~w2158;
assign w2161 = ~w2159 & ~w2160;
assign w2162 = w2057 & w2161;
assign w2163 = ~w2057 & ~w2161;
assign w2164 = ~w2162 & ~w2163;
assign w2165 = ~w1592 & ~w1859;
assign w2166 = (w1859 & ~w1862) | (w1859 & w17082) | (~w1862 & w17082);
assign w2167 = (w1862 & w17083) | (w1862 & w17084) | (w17083 & w17084);
assign w2168 = w2164 & ~w2167;
assign w2169 = ~w2164 & w2167;
assign w2170 = ~w2168 & ~w2169;
assign w2171 = (~w2056 & w2170) | (~w2056 & w17085) | (w2170 & w17085);
assign w2172 = ~w2170 & w17086;
assign w2173 = ~w2171 & ~w2172;
assign w2174 = (~w1867 & ~w1868) | (~w1867 & w17087) | (~w1868 & w17087);
assign w2175 = ~w2173 & w2174;
assign w2176 = w2173 & ~w2174;
assign w2177 = ~w2175 & ~w2176;
assign w2178 = w2055 & w2177;
assign w2179 = ~w2055 & ~w2177;
assign w2180 = ~w2178 & ~w2179;
assign w2181 = w2050 & w2180;
assign w2182 = ~w2050 & ~w2180;
assign w2183 = ~w2181 & ~w2182;
assign w2184 = w2049 & ~w2183;
assign w2185 = ~w2049 & w2183;
assign w2186 = ~w2184 & ~w2185;
assign w2187 = (~w1885 & ~w1881) | (~w1885 & w17088) | (~w1881 & w17088);
assign w2188 = ~w2186 & w2187;
assign w2189 = w2186 & ~w2187;
assign w2190 = ~w2188 & ~w2189;
assign w2191 = w2048 & w2190;
assign w2192 = ~w2048 & ~w2190;
assign w2193 = ~w2191 & ~w2192;
assign w2194 = w2047 & w2193;
assign w2195 = ~w2047 & ~w2193;
assign w2196 = ~w2194 & ~w2195;
assign w2197 = pi328 & ~w793;
assign w2198 = (~w1756 & ~w1758) | (~w1756 & w17089) | (~w1758 & w17089);
assign w2199 = ~w2197 & w2198;
assign w2200 = w2197 & ~w2198;
assign w2201 = ~w2199 & ~w2200;
assign w2202 = w2196 & w2201;
assign w2203 = ~w2196 & ~w2201;
assign w2204 = ~w2202 & ~w2203;
assign w2205 = w2042 & w2204;
assign w2206 = ~w2042 & ~w2204;
assign w2207 = ~w2205 & ~w2206;
assign w2208 = w2041 & w2207;
assign w2209 = ~w2041 & ~w2207;
assign w2210 = ~w2208 & ~w2209;
assign w2211 = ~w537 & w2210;
assign w2212 = w537 & ~w2210;
assign w2213 = ~w2211 & ~w2212;
assign w2214 = (~w1904 & ~w1902) | (~w1904 & w17090) | (~w1902 & w17090);
assign w2215 = ~pi330 & ~w537;
assign w2216 = (w1902 & w17091) | (w1902 & w17092) | (w17091 & w17092);
assign w2217 = w2213 & ~w2216;
assign w2218 = ~w2213 & w2216;
assign w2219 = ~w2217 & ~w2218;
assign w2220 = w2040 & w2219;
assign w2221 = ~w2040 & ~w2219;
assign w2222 = ~w2220 & ~w2221;
assign w2223 = w2036 & w2222;
assign w2224 = ~w2036 & ~w2222;
assign w2225 = ~w2223 & ~w2224;
assign w2226 = ~w2035 & ~w2225;
assign w2227 = w2035 & w2225;
assign w2228 = ~w2226 & ~w2227;
assign w2229 = pi268 & w2228;
assign w2230 = ~pi268 & ~w2228;
assign w2231 = ~w2229 & ~w2230;
assign w2232 = (~w1752 & w1919) | (~w1752 & w17093) | (w1919 & w17093);
assign w2233 = ~w1921 & ~w2232;
assign w2234 = w2231 & ~w2233;
assign w2235 = ~w2231 & w2233;
assign w2236 = ~w2234 & ~w2235;
assign w2237 = w2034 & ~w2236;
assign w2238 = (~w135 & ~w2236) | (~w135 & w17094) | (~w2236 & w17094);
assign w2239 = ~w2237 & w2238;
assign w2240 = (pi161 & ~w135) | (pi161 & w17095) | (~w135 & w17095);
assign w2241 = ~w2239 & w2240;
assign w2242 = ~pi160 & ~w1931;
assign w2243 = ~w2241 & w2242;
assign w2244 = ~pi075 & ~pi161;
assign w2245 = pi333 & w456;
assign w2246 = (~w466 & ~w2222) | (~w466 & w16895) | (~w2222 & w16895);
assign w2247 = pi332 & ~w2246;
assign w2248 = w971 & w2222;
assign w2249 = w2247 & ~w2248;
assign w2250 = (pi331 & ~w536) | (pi331 & w17096) | (~w536 & w17096);
assign w2251 = ~w2250 & w17641;
assign w2252 = (w2219 & w17098) | (w2219 & w17099) | (w17098 & w17099);
assign w2253 = ~w2251 & ~w2252;
assign w2254 = pi329 & ~w793;
assign w2255 = (~w2205 & ~w2207) | (~w2205 & w17100) | (~w2207 & w17100);
assign w2256 = pi328 & ~w955;
assign w2257 = pi327 & w1101;
assign w2258 = (w2193 & w17102) | (w2193 & w17103) | (w17102 & w17103);
assign w2259 = ~w2257 & w17642;
assign w2260 = ~w2258 & ~w2259;
assign w2261 = pi326 & w1339;
assign w2262 = (~w2182 & ~w2183) | (~w2182 & w17104) | (~w2183 & w17104);
assign w2263 = pi325 & w1602;
assign w2264 = pi323 & ~w2170;
assign w2265 = pi138 & pi259;
assign w2266 = (~w2265 & ~w2161) | (~w2265 & w17105) | (~w2161 & w17105);
assign w2267 = w2161 & w17106;
assign w2268 = ~w2266 & ~w2267;
assign w2269 = pi137 & pi260;
assign w2270 = (w2269 & w2159) | (w2269 & w16368) | (w2159 & w16368);
assign w2271 = ~w2159 & w16369;
assign w2272 = ~w2270 & ~w2271;
assign w2273 = w2154 & w17107;
assign w2274 = ~w2156 & ~w2273;
assign w2275 = ~w2135 & ~w2140;
assign w2276 = pi134 & pi263;
assign w2277 = pi132 & pi265;
assign w2278 = ~w2067 & ~w2114;
assign w2279 = ~w2066 & w2278;
assign w2280 = (w2277 & w2279) | (w2277 & w15835) | (w2279 & w15835);
assign w2281 = ~w2279 & w15836;
assign w2282 = ~w2280 & ~w2281;
assign w2283 = pi131 & pi266;
assign w2284 = ~w2078 & w17639;
assign w2285 = (w1786 & w17108) | (w1786 & w17109) | (w17108 & w17109);
assign w2286 = ~w2284 & ~w2285;
assign w2287 = w2079 & w2286;
assign w2288 = ~w2079 & ~w2286;
assign w2289 = (~w1790 & w16370) | (~w1790 & w16371) | (w16370 & w16371);
assign w2290 = ~w2070 & w2289;
assign w2291 = pi130 & pi267;
assign w2292 = pi128 & pi269;
assign w2293 = ~w2076 & ~w2292;
assign w2294 = w2076 & w2292;
assign w2295 = ~w2293 & ~w2294;
assign w2296 = ~w2285 & w17110;
assign w2297 = (w2295 & w2285) | (w2295 & w17111) | (w2285 & w17111);
assign w2298 = ~w2296 & ~w2297;
assign w2299 = ~w2291 & ~w2298;
assign w2300 = ~w2074 & w17639;
assign w2301 = ~w2300 & w17112;
assign w2302 = (~w2295 & w2300) | (~w2295 & w17113) | (w2300 & w17113);
assign w2303 = w2291 & ~w2301;
assign w2304 = ~w2302 & w2303;
assign w2305 = ~w2299 & ~w2304;
assign w2306 = (w2305 & w2290) | (w2305 & w16558) | (w2290 & w16558);
assign w2307 = ~w2290 & w16559;
assign w2308 = ~w2306 & ~w2307;
assign w2309 = ~w2283 & ~w2308;
assign w2310 = w2283 & w2308;
assign w2311 = ~w2309 & ~w2310;
assign w2312 = ~w2090 & w17643;
assign w2313 = (~w2312 & w2071) | (~w2312 & w17116) | (w2071 & w17116);
assign w2314 = w2107 & ~w2313;
assign w2315 = (w1790 & w17117) | (w1790 & w17118) | (w17117 & w17118);
assign w2316 = w2094 & ~w2312;
assign w2317 = ~w2315 & w2316;
assign w2318 = (~w2317 & w2109) | (~w2317 & w15837) | (w2109 & w15837);
assign w2319 = w2311 & ~w2318;
assign w2320 = ~w2311 & w2318;
assign w2321 = ~w2319 & ~w2320;
assign w2322 = pi133 & pi264;
assign w2323 = w2321 & ~w2322;
assign w2324 = ~w2321 & w2322;
assign w2325 = ~w2323 & ~w2324;
assign w2326 = w2282 & w2325;
assign w2327 = ~w2282 & ~w2325;
assign w2328 = ~w2326 & ~w2327;
assign w2329 = (~w2119 & w2124) | (~w2119 & w16123) | (w2124 & w16123);
assign w2330 = ~w2328 & w2329;
assign w2331 = w2328 & ~w2329;
assign w2332 = ~w2330 & ~w2331;
assign w2333 = ~w2276 & ~w2332;
assign w2334 = w2276 & w2332;
assign w2335 = ~w2333 & ~w2334;
assign w2336 = w2125 & ~w2133;
assign w2337 = ~w2121 & ~w2124;
assign w2338 = w2121 & w2124;
assign w2339 = ~w2337 & ~w2338;
assign w2340 = w2064 & w2339;
assign w2341 = ~w2336 & w16372;
assign w2342 = (~w2335 & w2336) | (~w2335 & w16373) | (w2336 & w16373);
assign w2343 = ~w2341 & ~w2342;
assign w2344 = (w2343 & w2140) | (w2343 & w16374) | (w2140 & w16374);
assign w2345 = ~w2140 & w16375;
assign w2346 = ~w2344 & ~w2345;
assign w2347 = pi136 & pi261;
assign w2348 = pi135 & pi262;
assign w2349 = w2347 & ~w2348;
assign w2350 = ~w2347 & w2348;
assign w2351 = ~w2349 & ~w2350;
assign w2352 = w2346 & w2351;
assign w2353 = ~w2346 & ~w2351;
assign w2354 = ~w2352 & ~w2353;
assign w2355 = w2274 & ~w2354;
assign w2356 = ~w2274 & w2354;
assign w2357 = ~w2355 & ~w2356;
assign w2358 = w2272 & w2357;
assign w2359 = ~w2272 & ~w2357;
assign w2360 = ~w2358 & ~w2359;
assign w2361 = w2268 & w2360;
assign w2362 = ~w2268 & ~w2360;
assign w2363 = ~w2361 & ~w2362;
assign w2364 = pi139 & pi258;
assign w2365 = w2363 & ~w2364;
assign w2366 = ~w2363 & w2364;
assign w2367 = ~w2365 & ~w2366;
assign w2368 = ~w2164 & ~w2166;
assign w2369 = w2164 & ~w2165;
assign w2370 = ~w2368 & ~w2369;
assign w2371 = w2367 & ~w2370;
assign w2372 = ~w2367 & w2370;
assign w2373 = ~w2371 & ~w2372;
assign w2374 = (~w2264 & w2373) | (~w2264 & w17119) | (w2373 & w17119);
assign w2375 = ~w2373 & w17120;
assign w2376 = ~w2374 & ~w2375;
assign w2377 = (~w2172 & ~w2173) | (~w2172 & w17121) | (~w2173 & w17121);
assign w2378 = ~w2376 & w2377;
assign w2379 = w2376 & ~w2377;
assign w2380 = ~w2378 & ~w2379;
assign w2381 = pi324 & ~w1865;
assign w2382 = (~w2054 & ~w2055) | (~w2054 & w17122) | (~w2055 & w17122);
assign w2383 = ~w2381 & w2382;
assign w2384 = w2381 & ~w2382;
assign w2385 = ~w2383 & ~w2384;
assign w2386 = w2380 & w2385;
assign w2387 = ~w2380 & ~w2385;
assign w2388 = ~w2386 & ~w2387;
assign w2389 = w2263 & w2388;
assign w2390 = ~w2263 & ~w2388;
assign w2391 = ~w2389 & ~w2390;
assign w2392 = ~w2262 & ~w2391;
assign w2393 = w2262 & w2391;
assign w2394 = ~w2392 & ~w2393;
assign w2395 = (~w2188 & ~w2190) | (~w2188 & w17123) | (~w2190 & w17123);
assign w2396 = w2394 & ~w2395;
assign w2397 = ~w2394 & w2395;
assign w2398 = ~w2396 & ~w2397;
assign w2399 = w2261 & w2398;
assign w2400 = ~w2261 & ~w2398;
assign w2401 = ~w2399 & ~w2400;
assign w2402 = w2260 & w2401;
assign w2403 = ~w2260 & ~w2401;
assign w2404 = ~w2402 & ~w2403;
assign w2405 = ~w2256 & ~w2404;
assign w2406 = w2256 & w2404;
assign w2407 = ~w2405 & ~w2406;
assign w2408 = (~w2200 & ~w2196) | (~w2200 & w17124) | (~w2196 & w17124);
assign w2409 = w2407 & ~w2408;
assign w2410 = ~w2407 & w2408;
assign w2411 = ~w2409 & ~w2410;
assign w2412 = ~w2255 & w2411;
assign w2413 = w2255 & ~w2411;
assign w2414 = ~w2412 & ~w2413;
assign w2415 = w2254 & w2414;
assign w2416 = ~w2254 & ~w2414;
assign w2417 = ~w2415 & ~w2416;
assign w2418 = (~w2214 & ~w2210) | (~w2214 & w17125) | (~w2210 & w17125);
assign w2419 = (pi330 & w2210) | (pi330 & w17126) | (w2210 & w17126);
assign w2420 = ~w2418 & w2419;
assign w2421 = ~w615 & w2420;
assign w2422 = pi330 & ~w615;
assign w2423 = ~w2420 & ~w2422;
assign w2424 = ~w2421 & ~w2423;
assign w2425 = w2417 & w2424;
assign w2426 = ~w2417 & ~w2424;
assign w2427 = ~w2425 & ~w2426;
assign w2428 = w2253 & w2427;
assign w2429 = ~w2253 & ~w2427;
assign w2430 = ~w2428 & ~w2429;
assign w2431 = ~w2249 & w2430;
assign w2432 = w2249 & ~w2430;
assign w2433 = ~w2431 & ~w2432;
assign w2434 = w2245 & ~w2433;
assign w2435 = ~w2245 & w2433;
assign w2436 = ~w2434 & ~w2435;
assign w2437 = (~w2226 & ~w2228) | (~w2226 & w17127) | (~w2228 & w17127);
assign w2438 = ~w2436 & ~w2437;
assign w2439 = w2436 & w2437;
assign w2440 = ~w2438 & ~w2439;
assign w2441 = pi269 & w2440;
assign w2442 = ~pi269 & ~w2440;
assign w2443 = ~w2441 & ~w2442;
assign w2444 = (~w2034 & w2231) | (~w2034 & w17128) | (w2231 & w17128);
assign w2445 = ~w2234 & ~w2444;
assign w2446 = ~w2443 & w2445;
assign w2447 = w2443 & ~w2445;
assign w2448 = ~w2446 & ~w2447;
assign w2449 = pi128 & pi310;
assign w2450 = w2031 & w17129;
assign w2451 = pi311 & w464;
assign w2452 = (~w2451 & ~w2031) | (~w2451 & w17130) | (~w2031 & w17130);
assign w2453 = ~w2450 & ~w2452;
assign w2454 = pi312 & ~w653;
assign w2455 = (~w2026 & ~w2028) | (~w2026 & w17131) | (~w2028 & w17131);
assign w2456 = (~w2012 & ~w2013) | (~w2012 & w17132) | (~w2013 & w17132);
assign w2457 = pi315 & w855;
assign w2458 = (~w2004 & ~w2006) | (~w2004 & w17133) | (~w2006 & w17133);
assign w2459 = ~w2457 & ~w2458;
assign w2460 = w2457 & w2458;
assign w2461 = ~w2459 & ~w2460;
assign w2462 = pi316 & w1159;
assign w2463 = pi317 & w1220;
assign w2464 = w1419 & w17134;
assign w2465 = w1692 & w17135;
assign w2466 = (~w1942 & ~w1943) | (~w1942 & w17136) | (~w1943 & w17136);
assign w2467 = (w1698 & w17139) | (w1698 & w17140) | (w17139 & w17140);
assign w2468 = pi138 & ~pi139;
assign w2469 = ~pi138 & pi139;
assign w2470 = ~w2468 & ~w2469;
assign w2471 = ~w1952 & w17141;
assign w2472 = (w2470 & w1952) | (w2470 & w17142) | (w1952 & w17142);
assign w2473 = ~w2471 & ~w2472;
assign w2474 = pi321 & ~w2473;
assign w2475 = ~w2474 & w17644;
assign w2476 = w2467 & w2475;
assign w2477 = w1693 & ~w1699;
assign w2478 = ~w1697 & w17144;
assign w2479 = ~w2477 & ~w2478;
assign w2480 = (w2474 & ~w2479) | (w2474 & w17145) | (~w2479 & w17145);
assign w2481 = ~w2476 & ~w2480;
assign w2482 = w2466 & w2481;
assign w2483 = ~w2466 & ~w2481;
assign w2484 = ~w2482 & ~w2483;
assign w2485 = w2465 & ~w2484;
assign w2486 = ~w2465 & w2484;
assign w2487 = ~w2485 & ~w2486;
assign w2488 = (~w1967 & ~w1969) | (~w1967 & w15838) | (~w1969 & w15838);
assign w2489 = w2487 & ~w2488;
assign w2490 = ~w2487 & w2488;
assign w2491 = ~w2489 & ~w2490;
assign w2492 = w2464 & w2491;
assign w2493 = ~w2464 & ~w2491;
assign w2494 = ~w2492 & ~w2493;
assign w2495 = (w1979 & w1722) | (w1979 & w17146) | (w1722 & w17146);
assign w2496 = (~w2494 & ~w1982) | (~w2494 & w17147) | (~w1982 & w17147);
assign w2497 = w1982 & w17148;
assign w2498 = ~w2496 & ~w2497;
assign w2499 = w2463 & w2498;
assign w2500 = ~w2463 & ~w2498;
assign w2501 = ~w2499 & ~w2500;
assign w2502 = w2462 & w2501;
assign w2503 = ~w2462 & ~w2501;
assign w2504 = ~w2502 & ~w2503;
assign w2505 = (~w1936 & w1989) | (~w1936 & w17149) | (w1989 & w17149);
assign w2506 = w1991 & ~w1994;
assign w2507 = ~w1997 & ~w2505;
assign w2508 = ~w2506 & w2507;
assign w2509 = ~w2504 & ~w2508;
assign w2510 = w2504 & w2508;
assign w2511 = ~w2509 & ~w2510;
assign w2512 = ~w2461 & w2511;
assign w2513 = w2461 & ~w2511;
assign w2514 = ~w2512 & ~w2513;
assign w2515 = w2456 & w2514;
assign w2516 = ~w2456 & ~w2514;
assign w2517 = ~w2515 & ~w2516;
assign w2518 = pi314 & w698;
assign w2519 = ~w2517 & w2518;
assign w2520 = w2517 & ~w2518;
assign w2521 = ~w2519 & ~w2520;
assign w2522 = (w653 & ~w2017) | (w653 & w17150) | (~w2017 & w17150);
assign w2523 = ~w2021 & ~w2522;
assign w2524 = w709 & w2523;
assign w2525 = (pi313 & w2523) | (pi313 & w17151) | (w2523 & w17151);
assign w2526 = ~w2524 & w2525;
assign w2527 = w2521 & w2526;
assign w2528 = ~w2521 & ~w2526;
assign w2529 = ~w2527 & ~w2528;
assign w2530 = ~w2455 & ~w2529;
assign w2531 = w2455 & w2529;
assign w2532 = ~w2530 & ~w2531;
assign w2533 = w2454 & w2532;
assign w2534 = ~w2454 & ~w2532;
assign w2535 = ~w2533 & ~w2534;
assign w2536 = w2453 & w2535;
assign w2537 = ~w2453 & ~w2535;
assign w2538 = ~w2536 & ~w2537;
assign w2539 = w2449 & ~w2538;
assign w2540 = ~w2449 & w2538;
assign w2541 = ~w2539 & ~w2540;
assign w2542 = w2448 & w2541;
assign w2543 = (~w135 & w2448) | (~w135 & w17152) | (w2448 & w17152);
assign w2544 = ~w2542 & w2543;
assign w2545 = (pi161 & ~w135) | (pi161 & w17153) | (~w135 & w17153);
assign w2546 = ~w2544 & w2545;
assign w2547 = ~pi160 & ~w2244;
assign w2548 = ~w2546 & w2547;
assign w2549 = ~pi076 & ~pi161;
assign w2550 = (~w2438 & ~w2440) | (~w2438 & w17154) | (~w2440 & w17154);
assign w2551 = ~pi270 & w2550;
assign w2552 = pi270 & ~w2550;
assign w2553 = ~w2551 & ~w2552;
assign w2554 = pi334 & w456;
assign w2555 = ~w2433 & w17155;
assign w2556 = ~w465 & w17156;
assign w2557 = (~w2556 & w2433) | (~w2556 & w17157) | (w2433 & w17157);
assign w2558 = ~w2555 & ~w2557;
assign w2559 = pi331 & ~w615;
assign w2560 = ~w2559 & w17645;
assign w2561 = (w2427 & w17159) | (w2427 & w17160) | (w17159 & w17160);
assign w2562 = ~w2560 & ~w2561;
assign w2563 = pi329 & ~w955;
assign w2564 = pi327 & w1339;
assign w2565 = pi326 & w1602;
assign w2566 = (~w2396 & ~w2398) | (~w2396 & w17161) | (~w2398 & w17161);
assign w2567 = ~w2565 & w2566;
assign w2568 = w2565 & ~w2566;
assign w2569 = ~w2567 & ~w2568;
assign w2570 = (~w2389 & ~w2391) | (~w2389 & w17162) | (~w2391 & w17162);
assign w2571 = pi324 & ~w2170;
assign w2572 = (~w2384 & ~w2380) | (~w2384 & w17163) | (~w2380 & w17163);
assign w2573 = w2571 & ~w2572;
assign w2574 = ~w2571 & w2572;
assign w2575 = ~w2573 & ~w2574;
assign w2576 = pi323 & ~w2373;
assign w2577 = ~w2271 & ~w2357;
assign w2578 = ~w2270 & ~w2577;
assign w2579 = w2360 & w17164;
assign w2580 = ~w2266 & ~w2578;
assign w2581 = w2266 & w2578;
assign w2582 = ~w2580 & ~w2581;
assign w2583 = ~w2361 & w2582;
assign w2584 = ~w2579 & ~w2583;
assign w2585 = pi138 & pi260;
assign w2586 = pi137 & pi261;
assign w2587 = pi136 & pi262;
assign w2588 = pi135 & pi263;
assign w2589 = ~w2334 & ~w2340;
assign w2590 = (~w2333 & ~w2589) | (~w2333 & w15839) | (~w2589 & w15839);
assign w2591 = w2322 & w2328;
assign w2592 = ~w2330 & ~w2591;
assign w2593 = pi132 & pi266;
assign w2594 = (~w2310 & w2318) | (~w2310 & w16376) | (w2318 & w16376);
assign w2595 = pi131 & pi267;
assign w2596 = (pi130 & w2290) | (pi130 & w17165) | (w2290 & w17165);
assign w2597 = w2595 & ~w2596;
assign w2598 = pi130 & pi268;
assign w2599 = ~w2285 & w17168;
assign w2600 = pi129 & pi269;
assign w2601 = pi128 & pi270;
assign w2602 = ~w2600 & ~w2601;
assign w2603 = w2600 & w2601;
assign w2604 = ~w2602 & ~w2603;
assign w2605 = ~w2599 & w17169;
assign w2606 = (w2604 & w2599) | (w2604 & w17170) | (w2599 & w17170);
assign w2607 = ~w2605 & ~w2606;
assign w2608 = w2598 & ~w2607;
assign w2609 = ~w2598 & w2607;
assign w2610 = ~w2608 & ~w2609;
assign w2611 = (w2291 & w2290) | (w2291 & w17171) | (w2290 & w17171);
assign w2612 = (~w2610 & ~w2611) | (~w2610 & w17172) | (~w2611 & w17172);
assign w2613 = ~w2597 & ~w2612;
assign w2614 = (w2298 & w2290) | (w2298 & w17173) | (w2290 & w17173);
assign w2615 = ~w2596 & ~w2610;
assign w2616 = ~w2596 & w2619;
assign w2617 = ~w2614 & ~w2616;
assign w2618 = ~w2613 & w2617;
assign w2619 = w2595 & ~w2610;
assign w2620 = ~w2595 & w2610;
assign w2621 = ~w2619 & ~w2620;
assign w2622 = w2614 & ~w2621;
assign w2623 = w2611 & w17174;
assign w2624 = ~w2622 & ~w2623;
assign w2625 = ~w2618 & w2624;
assign w2626 = ~w2594 & w2625;
assign w2627 = w2594 & ~w2625;
assign w2628 = ~w2626 & ~w2627;
assign w2629 = ~w2593 & ~w2628;
assign w2630 = w2593 & w2628;
assign w2631 = ~w2629 & ~w2630;
assign w2632 = ~w2277 & ~w2321;
assign w2633 = (~w2632 & w2279) | (~w2632 & w16561) | (w2279 & w16561);
assign w2634 = w2631 & w2633;
assign w2635 = ~w2631 & ~w2633;
assign w2636 = ~w2634 & ~w2635;
assign w2637 = (w2636 & w2330) | (w2636 & w15841) | (w2330 & w15841);
assign w2638 = ~w2330 & w15842;
assign w2639 = ~w2637 & ~w2638;
assign w2640 = pi133 & pi265;
assign w2641 = pi134 & pi264;
assign w2642 = ~w2640 & w2641;
assign w2643 = w2640 & ~w2641;
assign w2644 = ~w2642 & ~w2643;
assign w2645 = w2639 & ~w2644;
assign w2646 = ~w2639 & w2644;
assign w2647 = ~w2645 & ~w2646;
assign w2648 = w2590 & w2647;
assign w2649 = ~w2590 & ~w2647;
assign w2650 = ~w2648 & ~w2649;
assign w2651 = w2588 & w2650;
assign w2652 = ~w2588 & ~w2650;
assign w2653 = ~w2651 & ~w2652;
assign w2654 = (~w2348 & ~w2275) | (~w2348 & w16124) | (~w2275 & w16124);
assign w2655 = ~w2344 & ~w2654;
assign w2656 = w2653 & ~w2655;
assign w2657 = ~w2653 & w2655;
assign w2658 = ~w2656 & ~w2657;
assign w2659 = ~w2587 & w2658;
assign w2660 = w2587 & ~w2658;
assign w2661 = ~w2659 & ~w2660;
assign w2662 = ~w2347 & w2354;
assign w2663 = ~w2355 & ~w2662;
assign w2664 = w2661 & w2663;
assign w2665 = ~w2661 & ~w2663;
assign w2666 = ~w2664 & ~w2665;
assign w2667 = w2586 & w2666;
assign w2668 = ~w2586 & ~w2666;
assign w2669 = ~w2667 & ~w2668;
assign w2670 = w2585 & ~w2669;
assign w2671 = ~w2585 & w2669;
assign w2672 = ~w2670 & ~w2671;
assign w2673 = w2584 & w2672;
assign w2674 = ~w2584 & ~w2672;
assign w2675 = ~w2673 & ~w2674;
assign w2676 = pi140 & pi258;
assign w2677 = pi139 & pi259;
assign w2678 = ~w2364 & ~w2676;
assign w2679 = ~w2677 & w2678;
assign w2680 = ~pi139 & pi140;
assign w2681 = pi140 & pi259;
assign w2682 = pi139 & pi140;
assign w2683 = ~w458 & ~w2682;
assign w2684 = ~w2681 & ~w2683;
assign w2685 = ~w516 & ~w2680;
assign w2686 = ~w2684 & w2685;
assign w2687 = ~w2679 & ~w2686;
assign w2688 = w2363 & w17175;
assign w2689 = (w2687 & ~w2363) | (w2687 & w17176) | (~w2363 & w17176);
assign w2690 = ~w2688 & ~w2689;
assign w2691 = w2367 & ~w2368;
assign w2692 = (~w2369 & ~w2367) | (~w2369 & w17177) | (~w2367 & w17177);
assign w2693 = w2690 & ~w2692;
assign w2694 = ~w2690 & w2692;
assign w2695 = ~w2693 & ~w2694;
assign w2696 = w2675 & w2695;
assign w2697 = ~w2675 & ~w2695;
assign w2698 = ~w2696 & ~w2697;
assign w2699 = pi322 & w2698;
assign w2700 = (~w2375 & ~w2376) | (~w2375 & w17178) | (~w2376 & w17178);
assign w2701 = w2699 & ~w2700;
assign w2702 = ~w2699 & w2700;
assign w2703 = ~w2701 & ~w2702;
assign w2704 = w2576 & w2703;
assign w2705 = ~w2576 & ~w2703;
assign w2706 = ~w2704 & ~w2705;
assign w2707 = w2575 & w2706;
assign w2708 = ~w2575 & ~w2706;
assign w2709 = ~w2707 & ~w2708;
assign w2710 = w2570 & ~w2709;
assign w2711 = ~w2570 & w2709;
assign w2712 = ~w2710 & ~w2711;
assign w2713 = pi325 & ~w1865;
assign w2714 = w2712 & w2713;
assign w2715 = ~w2712 & ~w2713;
assign w2716 = ~w2714 & ~w2715;
assign w2717 = w2569 & w2716;
assign w2718 = ~w2569 & ~w2716;
assign w2719 = ~w2717 & ~w2718;
assign w2720 = w2564 & w2719;
assign w2721 = ~w2564 & ~w2719;
assign w2722 = ~w2720 & ~w2721;
assign w2723 = (~w2258 & ~w2401) | (~w2258 & w17179) | (~w2401 & w17179);
assign w2724 = w2722 & ~w2723;
assign w2725 = ~w2722 & w2723;
assign w2726 = ~w2724 & ~w2725;
assign w2727 = pi328 & w1101;
assign w2728 = (~w2406 & ~w2407) | (~w2406 & w17180) | (~w2407 & w17180);
assign w2729 = w2727 & ~w2728;
assign w2730 = ~w2727 & w2728;
assign w2731 = ~w2729 & ~w2730;
assign w2732 = w2726 & ~w2731;
assign w2733 = ~w2726 & w2731;
assign w2734 = ~w2732 & ~w2733;
assign w2735 = w2563 & ~w2734;
assign w2736 = ~w2563 & w2734;
assign w2737 = ~w2735 & ~w2736;
assign w2738 = (~w2412 & ~w2414) | (~w2412 & w17181) | (~w2414 & w17181);
assign w2739 = ~w2737 & w2738;
assign w2740 = w2737 & ~w2738;
assign w2741 = ~w2739 & ~w2740;
assign w2742 = (w2417 & w17183) | (w2417 & w17184) | (w17183 & w17184);
assign w2743 = w793 & w17646;
assign w2744 = ~w2742 & ~w2743;
assign w2745 = pi330 & w2744;
assign w2746 = ~w2741 & ~w2745;
assign w2747 = w2741 & w2745;
assign w2748 = ~w2746 & ~w2747;
assign w2749 = w2562 & w2748;
assign w2750 = ~w2562 & ~w2748;
assign w2751 = ~w2749 & ~w2750;
assign w2752 = ~w2246 & w17185;
assign w2753 = (w2752 & w2430) | (w2752 & w17186) | (w2430 & w17186);
assign w2754 = (~w2246 & w2430) | (~w2246 & w17187) | (w2430 & w17187);
assign w2755 = w537 & ~w2754;
assign w2756 = pi332 & ~w2753;
assign w2757 = ~w2755 & w2756;
assign w2758 = w2751 & w2757;
assign w2759 = ~w2751 & ~w2757;
assign w2760 = ~w2758 & ~w2759;
assign w2761 = ~w2558 & w2760;
assign w2762 = w2558 & ~w2760;
assign w2763 = ~w2761 & ~w2762;
assign w2764 = ~w2554 & w2763;
assign w2765 = w2554 & ~w2763;
assign w2766 = ~w2764 & ~w2765;
assign w2767 = w2553 & w2766;
assign w2768 = ~w2553 & ~w2766;
assign w2769 = ~w2767 & ~w2768;
assign w2770 = (~w2447 & ~w2448) | (~w2447 & w17188) | (~w2448 & w17188);
assign w2771 = ~w2769 & ~w2770;
assign w2772 = w2769 & w2770;
assign w2773 = ~w2771 & ~w2772;
assign w2774 = pi128 & pi309;
assign w2775 = pi311 & ~w653;
assign w2776 = pi312 & w709;
assign w2777 = pi313 & w698;
assign w2778 = pi314 & w855;
assign w2779 = pi315 & w1159;
assign w2780 = pi316 & w1220;
assign w2781 = (~w2502 & ~w2504) | (~w2502 & w17189) | (~w2504 & w17189);
assign w2782 = w1419 & w17190;
assign w2783 = w1692 & w17191;
assign w2784 = (~w2490 & ~w2491) | (~w2490 & w17192) | (~w2491 & w17192);
assign w2785 = pi319 & w1954;
assign w2786 = pi320 & ~w2473;
assign w2787 = w2467 & ~w2475;
assign w2788 = pi139 & ~pi140;
assign w2789 = ~w2680 & ~w2788;
assign w2790 = (w1948 & w17194) | (w1948 & w17195) | (w17194 & w17195);
assign w2791 = ~pi137 & ~w2790;
assign w2792 = ~w1948 & w2788;
assign w2793 = (pi137 & ~w2468) | (pi137 & w17196) | (~w2468 & w17196);
assign w2794 = ~w2792 & w2793;
assign w2795 = ~w2791 & ~w2794;
assign w2796 = (~pi138 & w1948) | (~pi138 & w17197) | (w1948 & w17197);
assign w2797 = (~w2789 & ~w1948) | (~w2789 & w17198) | (~w1948 & w17198);
assign w2798 = ~w2796 & ~w2797;
assign w2799 = ~pi138 & ~w2789;
assign w2800 = ~w2798 & ~w2799;
assign w2801 = ~w2795 & ~w2800;
assign w2802 = pi321 & w2801;
assign w2803 = ~w2787 & ~w2802;
assign w2804 = w2787 & w2801;
assign w2805 = ~w2803 & ~w2804;
assign w2806 = w2786 & w2805;
assign w2807 = ~w2786 & ~w2805;
assign w2808 = ~w2806 & ~w2807;
assign w2809 = (~w2482 & ~w2484) | (~w2482 & w17199) | (~w2484 & w17199);
assign w2810 = ~w2808 & ~w2809;
assign w2811 = w2808 & w2809;
assign w2812 = ~w2810 & ~w2811;
assign w2813 = w2785 & ~w2812;
assign w2814 = ~w2785 & w2812;
assign w2815 = ~w2813 & ~w2814;
assign w2816 = w2784 & w2815;
assign w2817 = ~w2784 & ~w2815;
assign w2818 = ~w2816 & ~w2817;
assign w2819 = w2783 & w2818;
assign w2820 = ~w2783 & ~w2818;
assign w2821 = ~w2819 & ~w2820;
assign w2822 = (~w2497 & ~w2498) | (~w2497 & w17200) | (~w2498 & w17200);
assign w2823 = ~w2821 & w2822;
assign w2824 = w2821 & ~w2822;
assign w2825 = ~w2823 & ~w2824;
assign w2826 = w2782 & ~w2825;
assign w2827 = ~w2782 & w2825;
assign w2828 = ~w2826 & ~w2827;
assign w2829 = w2781 & w2828;
assign w2830 = ~w2781 & ~w2828;
assign w2831 = ~w2829 & ~w2830;
assign w2832 = w2780 & w2831;
assign w2833 = ~w2780 & ~w2831;
assign w2834 = ~w2832 & ~w2833;
assign w2835 = (~w2459 & ~w2461) | (~w2459 & w17201) | (~w2461 & w17201);
assign w2836 = ~w2834 & ~w2835;
assign w2837 = w2834 & w2835;
assign w2838 = ~w2836 & ~w2837;
assign w2839 = w2779 & w2838;
assign w2840 = ~w2779 & ~w2838;
assign w2841 = ~w2839 & ~w2840;
assign w2842 = w2778 & w2841;
assign w2843 = ~w2778 & ~w2841;
assign w2844 = ~w2842 & ~w2843;
assign w2845 = (~w2515 & ~w2517) | (~w2515 & w17202) | (~w2517 & w17202);
assign w2846 = w2844 & w2845;
assign w2847 = ~w2844 & ~w2845;
assign w2848 = ~w2846 & ~w2847;
assign w2849 = w2521 & ~w2524;
assign w2850 = w2525 & ~w2849;
assign w2851 = w2848 & w2850;
assign w2852 = ~w2848 & ~w2850;
assign w2853 = ~w2851 & ~w2852;
assign w2854 = w2777 & ~w2853;
assign w2855 = ~w2777 & w2853;
assign w2856 = ~w2854 & ~w2855;
assign w2857 = ~w2776 & w2856;
assign w2858 = w2776 & ~w2856;
assign w2859 = ~w2857 & ~w2858;
assign w2860 = (~w2530 & ~w2532) | (~w2530 & w17203) | (~w2532 & w17203);
assign w2861 = w2859 & ~w2860;
assign w2862 = ~w2859 & w2860;
assign w2863 = ~w2861 & ~w2862;
assign w2864 = (~w2450 & ~w2535) | (~w2450 & w17204) | (~w2535 & w17204);
assign w2865 = ~w2863 & w2864;
assign w2866 = w2863 & ~w2864;
assign w2867 = ~w2865 & ~w2866;
assign w2868 = w2775 & ~w2867;
assign w2869 = ~w2775 & w2867;
assign w2870 = ~w2868 & ~w2869;
assign w2871 = ~pi129 & w2538;
assign w2872 = (~w464 & ~w2538) | (~w464 & w17205) | (~w2538 & w17205);
assign w2873 = pi310 & ~w2871;
assign w2874 = ~w2872 & w2873;
assign w2875 = w2870 & w2874;
assign w2876 = ~w2870 & ~w2874;
assign w2877 = ~w2875 & ~w2876;
assign w2878 = ~w2774 & w2877;
assign w2879 = w2774 & ~w2877;
assign w2880 = ~w2878 & ~w2879;
assign w2881 = w2773 & ~w2880;
assign w2882 = (~w135 & w2773) | (~w135 & w17206) | (w2773 & w17206);
assign w2883 = ~w2881 & w2882;
assign w2884 = (pi161 & ~w135) | (pi161 & w17207) | (~w135 & w17207);
assign w2885 = ~w2883 & w2884;
assign w2886 = ~pi160 & ~w2549;
assign w2887 = ~w2885 & w2886;
assign w2888 = ~pi077 & ~pi161;
assign w2889 = pi128 & pi308;
assign w2890 = pi312 & w698;
assign w2891 = pi314 & w1159;
assign w2892 = (~w2842 & ~w2844) | (~w2842 & w17208) | (~w2844 & w17208);
assign w2893 = w2891 & ~w2892;
assign w2894 = ~w2891 & w2892;
assign w2895 = ~w2893 & ~w2894;
assign w2896 = pi315 & w1220;
assign w2897 = (~w2837 & ~w2838) | (~w2837 & w17209) | (~w2838 & w17209);
assign w2898 = ~w2896 & w2897;
assign w2899 = w2896 & ~w2897;
assign w2900 = ~w2898 & ~w2899;
assign w2901 = w1419 & w17210;
assign w2902 = w1692 & w17211;
assign w2903 = pi318 & w1954;
assign w2904 = (~w2817 & ~w2818) | (~w2817 & w17212) | (~w2818 & w17212);
assign w2905 = pi319 & ~w2473;
assign w2906 = pi320 & w2801;
assign w2907 = ~pi141 & w2789;
assign w2908 = pi140 & pi141;
assign w2909 = pi139 & pi141;
assign w2910 = (~w2909 & w1948) | (~w2909 & w17213) | (w1948 & w17213);
assign w2911 = ~w2910 & w17214;
assign w2912 = pi141 & w2680;
assign w2913 = ~pi140 & ~pi141;
assign w2914 = (~w2912 & ~w1948) | (~w2912 & w17215) | (~w1948 & w17215);
assign w2915 = ~pi138 & w2913;
assign w2916 = w1948 & w17216;
assign w2917 = (~pi137 & w2916) | (~pi137 & w17217) | (w2916 & w17217);
assign w2918 = pi138 & pi140;
assign w2919 = (pi141 & w1948) | (pi141 & w17218) | (w1948 & w17218);
assign w2920 = (pi137 & w2918) | (pi137 & w17219) | (w2918 & w17219);
assign w2921 = ~w2919 & w2920;
assign w2922 = (~w2907 & w2914) | (~w2907 & w17220) | (w2914 & w17220);
assign w2923 = ~w2921 & w2922;
assign w2924 = ~w2911 & ~w2917;
assign w2925 = w2923 & w2924;
assign w2926 = pi321 & w2925;
assign w2927 = (~w2804 & ~w2805) | (~w2804 & w17221) | (~w2805 & w17221);
assign w2928 = ~w2926 & w2927;
assign w2929 = w2926 & ~w2927;
assign w2930 = ~w2928 & ~w2929;
assign w2931 = w2906 & w2930;
assign w2932 = ~w2906 & ~w2930;
assign w2933 = ~w2931 & ~w2932;
assign w2934 = (~w2785 & ~w2809) | (~w2785 & w17222) | (~w2809 & w17222);
assign w2935 = ~w2810 & ~w2934;
assign w2936 = ~w2933 & ~w2935;
assign w2937 = w2933 & w2935;
assign w2938 = ~w2936 & ~w2937;
assign w2939 = w2905 & ~w2938;
assign w2940 = ~w2905 & w2938;
assign w2941 = ~w2939 & ~w2940;
assign w2942 = w2904 & w2941;
assign w2943 = ~w2904 & ~w2941;
assign w2944 = ~w2942 & ~w2943;
assign w2945 = w2903 & w2944;
assign w2946 = ~w2903 & ~w2944;
assign w2947 = ~w2945 & ~w2946;
assign w2948 = (~w2823 & ~w2825) | (~w2823 & w17223) | (~w2825 & w17223);
assign w2949 = w2947 & w2948;
assign w2950 = ~w2947 & ~w2948;
assign w2951 = ~w2949 & ~w2950;
assign w2952 = w2902 & ~w2951;
assign w2953 = ~w2902 & w2951;
assign w2954 = ~w2952 & ~w2953;
assign w2955 = (~w2830 & ~w2831) | (~w2830 & w17224) | (~w2831 & w17224);
assign w2956 = w2954 & w2955;
assign w2957 = ~w2954 & ~w2955;
assign w2958 = ~w2956 & ~w2957;
assign w2959 = w2901 & w2958;
assign w2960 = ~w2901 & ~w2958;
assign w2961 = ~w2959 & ~w2960;
assign w2962 = w2900 & w2961;
assign w2963 = ~w2900 & ~w2961;
assign w2964 = ~w2962 & ~w2963;
assign w2965 = w2895 & w2964;
assign w2966 = ~w2895 & ~w2964;
assign w2967 = ~w2965 & ~w2966;
assign w2968 = (~w2777 & ~w2848) | (~w2777 & w17225) | (~w2848 & w17225);
assign w2969 = ~w2852 & ~w2968;
assign w2970 = w855 & w2969;
assign w2971 = pi313 & w855;
assign w2972 = ~w2969 & ~w2971;
assign w2973 = ~w2970 & ~w2972;
assign w2974 = w2967 & w2973;
assign w2975 = ~w2967 & ~w2973;
assign w2976 = ~w2974 & ~w2975;
assign w2977 = w2890 & w2976;
assign w2978 = ~w2890 & ~w2976;
assign w2979 = ~w2977 & ~w2978;
assign w2980 = (~w2858 & ~w2859) | (~w2858 & w17226) | (~w2859 & w17226);
assign w2981 = w2979 & ~w2980;
assign w2982 = ~w2979 & w2980;
assign w2983 = ~w2981 & ~w2982;
assign w2984 = pi311 & w709;
assign w2985 = (~w2865 & ~w2867) | (~w2865 & w17227) | (~w2867 & w17227);
assign w2986 = w2984 & w2985;
assign w2987 = ~w2984 & ~w2985;
assign w2988 = ~w2986 & ~w2987;
assign w2989 = w2983 & ~w2988;
assign w2990 = ~w2983 & w2988;
assign w2991 = ~w2989 & ~w2990;
assign w2992 = (~w2872 & ~w2870) | (~w2872 & w17228) | (~w2870 & w17228);
assign w2993 = (pi310 & w2992) | (pi310 & w17229) | (w2992 & w17229);
assign w2994 = ~w17650 & w2993;
assign w2995 = ~w2991 & w2994;
assign w2996 = w2991 & ~w2994;
assign w2997 = ~w2995 & ~w2996;
assign w2998 = ~pi129 & ~w2877;
assign w2999 = pi309 & w464;
assign w3000 = (~w2999 & w2877) | (~w2999 & w17230) | (w2877 & w17230);
assign w3001 = ~w2998 & ~w3000;
assign w3002 = w2997 & ~w3001;
assign w3003 = ~w2997 & w3001;
assign w3004 = ~w3002 & ~w3003;
assign w3005 = ~w2889 & w3004;
assign w3006 = w2889 & ~w3004;
assign w3007 = ~w3005 & ~w3006;
assign w3008 = pi335 & w456;
assign w3009 = (pi333 & ~w536) | (pi333 & w17231) | (~w536 & w17231);
assign w3010 = (~w2557 & w2760) | (~w2557 & w17232) | (w2760 & w17232);
assign w3011 = ~w3009 & ~w3010;
assign w3012 = (w2760 & w17233) | (w2760 & w17234) | (w17233 & w17234);
assign w3013 = ~w3011 & ~w3012;
assign w3014 = pi332 & ~w615;
assign w3015 = (w3014 & w2758) | (w3014 & w17235) | (w2758 & w17235);
assign w3016 = ~w2758 & w17236;
assign w3017 = ~w3015 & ~w3016;
assign w3018 = (~w2561 & ~w2748) | (~w2561 & w17237) | (~w2748 & w17237);
assign w3019 = (~w2735 & ~w2737) | (~w2735 & w17238) | (~w2737 & w17238);
assign w3020 = ~w3018 & w3019;
assign w3021 = w3018 & ~w3019;
assign w3022 = ~w3020 & ~w3021;
assign w3023 = pi331 & ~w793;
assign w3024 = pi328 & w1339;
assign w3025 = (~w3024 & w2733) | (~w3024 & w17239) | (w2733 & w17239);
assign w3026 = ~w2733 & w17240;
assign w3027 = ~w3025 & ~w3026;
assign w3028 = (~w2720 & ~w2722) | (~w2720 & w17241) | (~w2722 & w17241);
assign w3029 = pi327 & w1602;
assign w3030 = w3028 & ~w3029;
assign w3031 = ~w3028 & w3029;
assign w3032 = ~w3030 & ~w3031;
assign w3033 = (~w2568 & ~w2569) | (~w2568 & w17242) | (~w2569 & w17242);
assign w3034 = pi326 & ~w1865;
assign w3035 = (~w2711 & ~w2712) | (~w2711 & w17243) | (~w2712 & w17243);
assign w3036 = pi325 & ~w2170;
assign w3037 = ~w3035 & w3036;
assign w3038 = w3035 & ~w3036;
assign w3039 = ~w3037 & ~w3038;
assign w3040 = (~w2573 & ~w2706) | (~w2573 & w17244) | (~w2706 & w17244);
assign w3041 = pi323 & w2698;
assign w3042 = (~w2366 & ~w2675) | (~w2366 & w16377) | (~w2675 & w16377);
assign w3043 = ~w2675 & ~w2677;
assign w3044 = (pi139 & w2675) | (pi139 & w16378) | (w2675 & w16378);
assign w3045 = ~w3042 & w3044;
assign w3046 = pi137 & pi262;
assign w3047 = (~w2660 & ~w2663) | (~w2660 & w16125) | (~w2663 & w16125);
assign w3048 = ~w2344 & ~w2652;
assign w3049 = (~w2651 & ~w3048) | (~w2651 & w16126) | (~w3048 & w16126);
assign w3050 = (~w2641 & ~w2590) | (~w2641 & w16379) | (~w2590 & w16379);
assign w3051 = ~w2639 & ~w2640;
assign w3052 = w2639 & w2640;
assign w3053 = ~w3051 & ~w3052;
assign w3054 = ~w2590 & ~w3053;
assign w3055 = pi134 & pi265;
assign w3056 = ~w2629 & w2633;
assign w3057 = pi131 & pi268;
assign w3058 = pi130 & pi269;
assign w3059 = ~w2293 & ~w2602;
assign w3060 = pi129 & pi270;
assign w3061 = pi128 & pi271;
assign w3062 = ~w3060 & ~w3061;
assign w3063 = w3060 & w3061;
assign w3064 = ~w3062 & ~w3063;
assign w3065 = ~w3064 & w17724;
assign w3066 = ~w2602 & ~w3063;
assign w3067 = (w2285 & w17250) | (w2285 & w17251) | (w17250 & w17251);
assign w3068 = ~w3065 & ~w3067;
assign w3069 = w3058 & w3068;
assign w3070 = ~w3058 & ~w3068;
assign w3071 = ~w3069 & ~w3070;
assign w3072 = ~w2304 & ~w2608;
assign w3073 = (w2290 & w17254) | (w2290 & w17255) | (w17254 & w17255);
assign w3074 = w3071 & w3073;
assign w3075 = ~w3071 & ~w3073;
assign w3076 = ~w3074 & ~w3075;
assign w3077 = ~w3057 & ~w3076;
assign w3078 = w3057 & w3076;
assign w3079 = ~w3077 & ~w3078;
assign w3080 = (w2290 & w17256) | (w2290 & w17257) | (w17256 & w17257);
assign w3081 = ~w2615 & ~w3080;
assign w3082 = ~w2611 & ~w2614;
assign w3083 = w2610 & w3082;
assign w3084 = (~w2595 & w3082) | (~w2595 & w2620) | (w3082 & w2620);
assign w3085 = ~w3083 & w3084;
assign w3086 = (~w3081 & w2594) | (~w3081 & w17258) | (w2594 & w17258);
assign w3087 = w3079 & ~w3086;
assign w3088 = (w2594 & w17259) | (w2594 & w17260) | (w17259 & w17260);
assign w3089 = ~w3087 & ~w3088;
assign w3090 = (w2633 & w17261) | (w2633 & w17262) | (w17261 & w17262);
assign w3091 = ~w2630 & ~w3089;
assign w3092 = (w3091 & ~w2633) | (w3091 & w17263) | (~w2633 & w17263);
assign w3093 = ~w3090 & ~w3092;
assign w3094 = pi133 & pi266;
assign w3095 = pi132 & pi267;
assign w3096 = w3094 & ~w3095;
assign w3097 = ~w3094 & w3095;
assign w3098 = ~w3096 & ~w3097;
assign w3099 = w3093 & w3098;
assign w3100 = ~w3093 & ~w3098;
assign w3101 = ~w3099 & ~w3100;
assign w3102 = w2636 & w2640;
assign w3103 = ~w2636 & ~w2640;
assign w3104 = (~w2592 & w17264) | (~w2592 & w17265) | (w17264 & w17265);
assign w3105 = (w2592 & w17266) | (w2592 & w17267) | (w17266 & w17267);
assign w3106 = ~w3104 & ~w3105;
assign w3107 = ~w3055 & ~w3106;
assign w3108 = w3055 & w3106;
assign w3109 = ~w3107 & ~w3108;
assign w3110 = (w3109 & w3050) | (w3109 & w16127) | (w3050 & w16127);
assign w3111 = ~w3050 & w16128;
assign w3112 = ~w3110 & ~w3111;
assign w3113 = (w16126 & w16562) | (w16126 & w16563) | (w16562 & w16563);
assign w3114 = (~w16126 & w16564) | (~w16126 & w16565) | (w16564 & w16565);
assign w3115 = ~w3113 & ~w3114;
assign w3116 = pi136 & pi263;
assign w3117 = pi135 & pi264;
assign w3118 = w3116 & ~w3117;
assign w3119 = ~w3116 & w3117;
assign w3120 = ~w3118 & ~w3119;
assign w3121 = w3115 & w3120;
assign w3122 = ~w3115 & ~w3120;
assign w3123 = ~w3121 & ~w3122;
assign w3124 = w3047 & w3123;
assign w3125 = ~w3047 & ~w3123;
assign w3126 = ~w3124 & ~w3125;
assign w3127 = ~w3046 & ~w3126;
assign w3128 = w3046 & w3126;
assign w3129 = ~w3127 & ~w3128;
assign w3130 = (~w2578 & w2666) | (~w2578 & w16381) | (w2666 & w16381);
assign w3131 = ~w2667 & ~w3130;
assign w3132 = w3129 & w3131;
assign w3133 = ~w3129 & ~w3131;
assign w3134 = ~w3132 & ~w3133;
assign w3135 = w2585 & w17647;
assign w3136 = (w2360 & w17268) | (w2360 & w17269) | (w17268 & w17269);
assign w3137 = ~w2578 & w2669;
assign w3138 = w2578 & ~w2669;
assign w3139 = ~w3137 & ~w3138;
assign w3140 = (~w3135 & ~w3139) | (~w3135 & w15845) | (~w3139 & w15845);
assign w3141 = w3134 & w3140;
assign w3142 = ~w3134 & ~w3140;
assign w3143 = ~w3141 & ~w3142;
assign w3144 = pi139 & pi260;
assign w3145 = pi138 & pi261;
assign w3146 = w3144 & ~w3145;
assign w3147 = ~w3144 & w3145;
assign w3148 = ~w3146 & ~w3147;
assign w3149 = w3143 & w3148;
assign w3150 = ~w3143 & ~w3148;
assign w3151 = ~w3149 & ~w3150;
assign w3152 = ~w3045 & w3151;
assign w3153 = w3045 & ~w3151;
assign w3154 = ~w3152 & ~w3153;
assign w3155 = ~pi139 & ~w2675;
assign w3156 = ~w3044 & ~w3155;
assign w3157 = (~w2363 & ~w2675) | (~w2363 & w16566) | (~w2675 & w16566);
assign w3158 = ~w3156 & w3157;
assign w3159 = w2675 & w2677;
assign w3160 = ~w3043 & ~w3159;
assign w3161 = ~w3158 & w15847;
assign w3162 = (~w2681 & w3158) | (~w2681 & w15848) | (w3158 & w15848);
assign w3163 = ~w3161 & ~w3162;
assign w3164 = ~w3154 & ~w3163;
assign w3165 = w3154 & w3163;
assign w3166 = ~w3164 & ~w3165;
assign w3167 = pi141 & pi258;
assign w3168 = w3166 & w3167;
assign w3169 = ~w3166 & ~w3167;
assign w3170 = ~w3168 & ~w3169;
assign w3171 = ~w2367 & ~w2369;
assign w3172 = w2363 & w2686;
assign w3173 = (~w2679 & w2363) | (~w2679 & w17270) | (w2363 & w17270);
assign w3174 = ~w3172 & w3173;
assign w3175 = w2675 & w3174;
assign w3176 = ~w2675 & ~w3174;
assign w3177 = ~w3175 & ~w3176;
assign w3178 = ~w3171 & w3177;
assign w3179 = ~w2691 & ~w3177;
assign w3180 = ~w3178 & ~w3179;
assign w3181 = w3170 & ~w3180;
assign w3182 = ~w3170 & w3180;
assign w3183 = ~w3181 & ~w3182;
assign w3184 = pi322 & ~w3183;
assign w3185 = (~w2701 & ~w2703) | (~w2701 & w17271) | (~w2703 & w17271);
assign w3186 = (w3185 & w3183) | (w3185 & w17272) | (w3183 & w17272);
assign w3187 = ~w3183 & w17273;
assign w3188 = ~w3186 & ~w3187;
assign w3189 = ~w3041 & ~w3188;
assign w3190 = w3041 & w3188;
assign w3191 = ~w3189 & ~w3190;
assign w3192 = ~w3040 & w3191;
assign w3193 = w3040 & ~w3191;
assign w3194 = ~w3192 & ~w3193;
assign w3195 = pi324 & ~w2373;
assign w3196 = ~w3194 & w3195;
assign w3197 = w3194 & ~w3195;
assign w3198 = ~w3196 & ~w3197;
assign w3199 = w3039 & ~w3198;
assign w3200 = ~w3039 & w3198;
assign w3201 = ~w3199 & ~w3200;
assign w3202 = w3034 & w3201;
assign w3203 = ~w3034 & ~w3201;
assign w3204 = ~w3202 & ~w3203;
assign w3205 = w3033 & ~w3204;
assign w3206 = ~w3033 & w3204;
assign w3207 = ~w3205 & ~w3206;
assign w3208 = w3032 & w3207;
assign w3209 = ~w3032 & ~w3207;
assign w3210 = ~w3208 & ~w3209;
assign w3211 = ~w3027 & ~w3210;
assign w3212 = w3027 & w3210;
assign w3213 = ~w3211 & ~w3212;
assign w3214 = ~w3023 & w3213;
assign w3215 = w3023 & ~w3213;
assign w3216 = ~w3214 & ~w3215;
assign w3217 = w3022 & w3216;
assign w3218 = ~w3022 & ~w3216;
assign w3219 = ~w3217 & ~w3218;
assign w3220 = pi329 & w1101;
assign w3221 = w2741 & w2744;
assign w3222 = (~w15849 & ~w2741) | (~w15849 & w17274) | (~w2741 & w17274);
assign w3223 = (w2741 & w17275) | (w2741 & w17276) | (w17275 & w17276);
assign w3224 = (pi330 & w2742) | (pi330 & w17277) | (w2742 & w17277);
assign w3225 = ~w2747 & ~w3224;
assign w3226 = ~w3223 & ~w3225;
assign w3227 = (w3220 & w3225) | (w3220 & w15850) | (w3225 & w15850);
assign w3228 = ~w3225 & w15851;
assign w3229 = ~w3227 & ~w3228;
assign w3230 = w3219 & w3229;
assign w3231 = ~w3219 & ~w3229;
assign w3232 = ~w3230 & ~w3231;
assign w3233 = w3017 & w3232;
assign w3234 = ~w3017 & ~w3232;
assign w3235 = ~w3233 & ~w3234;
assign w3236 = w3013 & ~w3235;
assign w3237 = ~w3013 & w3235;
assign w3238 = ~w3236 & ~w3237;
assign w3239 = ~w466 & ~w3238;
assign w3240 = w466 & w3238;
assign w3241 = ~w3239 & ~w3240;
assign w3242 = ~w465 & w17278;
assign w3243 = (~w3242 & w2763) | (~w3242 & w17279) | (w2763 & w17279);
assign w3244 = w3241 & ~w3243;
assign w3245 = ~w3241 & w3243;
assign w3246 = ~w3244 & ~w3245;
assign w3247 = w3008 & w3246;
assign w3248 = ~w3008 & ~w3246;
assign w3249 = ~w3247 & ~w3248;
assign w3250 = ~w2551 & ~w2767;
assign w3251 = ~w3249 & w3250;
assign w3252 = w3249 & ~w3250;
assign w3253 = ~w3251 & ~w3252;
assign w3254 = pi271 & w3253;
assign w3255 = ~pi271 & ~w3253;
assign w3256 = ~w3254 & ~w3255;
assign w3257 = (~w2771 & ~w2773) | (~w2771 & w17280) | (~w2773 & w17280);
assign w3258 = w3256 & ~w3257;
assign w3259 = ~w3256 & w3257;
assign w3260 = ~w3258 & ~w3259;
assign w3261 = ~w3007 & w3260;
assign w3262 = (~w135 & w3260) | (~w135 & w17281) | (w3260 & w17281);
assign w3263 = ~w3261 & w3262;
assign w3264 = (pi161 & ~w135) | (pi161 & w17282) | (~w135 & w17282);
assign w3265 = ~w3263 & w3264;
assign w3266 = ~pi160 & ~w2888;
assign w3267 = ~w3265 & w3266;
assign w3268 = ~pi078 & ~pi161;
assign w3269 = pi128 & pi307;
assign w3270 = pi308 & w464;
assign w3271 = (~w3270 & w3004) | (~w3270 & w17283) | (w3004 & w17283);
assign w3272 = ~w3004 & w17284;
assign w3273 = ~w3271 & ~w3272;
assign w3274 = pi310 & w709;
assign w3275 = pi311 & w698;
assign w3276 = (~w2977 & ~w2979) | (~w2977 & w17285) | (~w2979 & w17285);
assign w3277 = pi312 & w855;
assign w3278 = pi313 & w1159;
assign w3279 = pi314 & w1220;
assign w3280 = w1419 & w17286;
assign w3281 = ~w3280 & w17648;
assign w3282 = (w2900 & w17287) | (w2900 & w17288) | (w17287 & w17288);
assign w3283 = ~w3281 & ~w3282;
assign w3284 = w1692 & w17289;
assign w3285 = (~w2957 & ~w2958) | (~w2957 & w15853) | (~w2958 & w15853);
assign w3286 = pi318 & ~w2473;
assign w3287 = pi319 & w2801;
assign w3288 = (~w2905 & ~w2935) | (~w2905 & w15854) | (~w2935 & w15854);
assign w3289 = ~w2936 & ~w3288;
assign w3290 = ~w3287 & ~w3289;
assign w3291 = w3287 & w3289;
assign w3292 = ~w3290 & ~w3291;
assign w3293 = pi320 & w2925;
assign w3294 = (~w2918 & w1948) | (~w2918 & w17290) | (w1948 & w17290);
assign w3295 = pi137 & ~w3294;
assign w3296 = ~w2682 & ~w2908;
assign w3297 = (w3296 & w2910) | (w3296 & w17291) | (w2910 & w17291);
assign w3298 = ~w3295 & w3297;
assign w3299 = ~pi142 & w3298;
assign w3300 = pi142 & ~w3298;
assign w3301 = ~w3299 & ~w3300;
assign w3302 = pi141 & w3301;
assign w3303 = ~pi141 & ~w3301;
assign w3304 = ~w3302 & ~w3303;
assign w3305 = pi321 & w3304;
assign w3306 = (~w2929 & ~w2930) | (~w2929 & w17292) | (~w2930 & w17292);
assign w3307 = ~w3305 & w3306;
assign w3308 = w3305 & ~w3306;
assign w3309 = ~w3307 & ~w3308;
assign w3310 = w3293 & w3309;
assign w3311 = ~w3293 & ~w3309;
assign w3312 = ~w3310 & ~w3311;
assign w3313 = w3292 & w3312;
assign w3314 = ~w3292 & ~w3312;
assign w3315 = ~w3313 & ~w3314;
assign w3316 = ~w3315 & w17649;
assign w3317 = (w2944 & w17293) | (w2944 & w17294) | (w17293 & w17294);
assign w3318 = ~w3316 & ~w3317;
assign w3319 = w3286 & ~w3318;
assign w3320 = ~w3286 & w3318;
assign w3321 = ~w3319 & ~w3320;
assign w3322 = ~w2949 & ~w3321;
assign w3323 = pi317 & w1954;
assign w3324 = (~w2902 & ~w1954) | (~w2902 & w17295) | (~w1954 & w17295);
assign w3325 = (~w1693 & ~w2948) | (~w1693 & w17296) | (~w2948 & w17296);
assign w3326 = (w1954 & w2948) | (w1954 & w17297) | (w2948 & w17297);
assign w3327 = ~w3325 & w3326;
assign w3328 = ~w3324 & ~w3327;
assign w3329 = w3322 & ~w3328;
assign w3330 = ~w2950 & w3321;
assign w3331 = ~w3325 & w3330;
assign w3332 = (w3323 & w2949) | (w3323 & w17298) | (w2949 & w17298);
assign w3333 = ~w3331 & w3332;
assign w3334 = w2950 & ~w3321;
assign w3335 = ~w3330 & ~w3334;
assign w3336 = (~w1954 & ~w2951) | (~w1954 & w17299) | (~w2951 & w17299);
assign w3337 = ~w3335 & w3336;
assign w3338 = ~w3329 & ~w3333;
assign w3339 = ~w3337 & w3338;
assign w3340 = w3285 & w3339;
assign w3341 = ~w3285 & ~w3339;
assign w3342 = ~w3340 & ~w3341;
assign w3343 = w3284 & ~w3342;
assign w3344 = ~w3284 & w3342;
assign w3345 = ~w3343 & ~w3344;
assign w3346 = w3283 & ~w3345;
assign w3347 = ~w3283 & w3345;
assign w3348 = ~w3346 & ~w3347;
assign w3349 = w3279 & w3348;
assign w3350 = ~w3279 & ~w3348;
assign w3351 = ~w3349 & ~w3350;
assign w3352 = (~w2893 & ~w2895) | (~w2893 & w17300) | (~w2895 & w17300);
assign w3353 = w3351 & ~w3352;
assign w3354 = ~w3351 & w3352;
assign w3355 = ~w3353 & ~w3354;
assign w3356 = (~w2970 & ~w2973) | (~w2970 & w17301) | (~w2973 & w17301);
assign w3357 = w3355 & ~w3356;
assign w3358 = ~w3355 & w3356;
assign w3359 = ~w3357 & ~w3358;
assign w3360 = w3278 & w3359;
assign w3361 = ~w3278 & ~w3359;
assign w3362 = ~w3360 & ~w3361;
assign w3363 = ~w3277 & ~w3362;
assign w3364 = w3277 & w3362;
assign w3365 = ~w3363 & ~w3364;
assign w3366 = w3276 & ~w3365;
assign w3367 = ~w3276 & w3365;
assign w3368 = ~w3366 & ~w3367;
assign w3369 = (~w2987 & ~w2988) | (~w2987 & w17302) | (~w2988 & w17302);
assign w3370 = w3368 & w3369;
assign w3371 = ~w3368 & ~w3369;
assign w3372 = ~w3370 & ~w3371;
assign w3373 = w3275 & w3372;
assign w3374 = ~w3275 & ~w3372;
assign w3375 = ~w3373 & ~w3374;
assign w3376 = w3274 & w3375;
assign w3377 = ~w3274 & ~w3375;
assign w3378 = ~w3376 & ~w3377;
assign w3379 = pi310 & w17650;
assign w3380 = ~w2995 & ~w3379;
assign w3381 = w3378 & ~w3380;
assign w3382 = ~w3378 & w3380;
assign w3383 = ~w3381 & ~w3382;
assign w3384 = w597 & ~w2997;
assign w3385 = ~w2997 & ~w2998;
assign w3386 = (pi128 & ~w2877) | (pi128 & w459) | (~w2877 & w459);
assign w3387 = ~w3385 & w3386;
assign w3388 = ~w3387 & w17303;
assign w3389 = (pi130 & w3387) | (pi130 & w17304) | (w3387 & w17304);
assign w3390 = pi309 & ~w3388;
assign w3391 = ~w3389 & w3390;
assign w3392 = w3383 & w3391;
assign w3393 = ~w3383 & ~w3391;
assign w3394 = ~w3392 & ~w3393;
assign w3395 = ~w3273 & ~w3394;
assign w3396 = w3273 & w3394;
assign w3397 = ~w3395 & ~w3396;
assign w3398 = w3269 & w3397;
assign w3399 = ~w3269 & ~w3397;
assign w3400 = ~w3398 & ~w3399;
assign w3401 = (~w3251 & ~w3253) | (~w3251 & w17305) | (~w3253 & w17305);
assign w3402 = pi336 & w456;
assign w3403 = ~w465 & w17306;
assign w3404 = w456 & ~w2763;
assign w3405 = (~w3404 & ~w3238) | (~w3404 & w15856) | (~w3238 & w15856);
assign w3406 = ~w3239 & ~w3405;
assign w3407 = (pi334 & w3406) | (pi334 & w17307) | (w3406 & w17307);
assign w3408 = ~w537 & w3406;
assign w3409 = w3407 & ~w3408;
assign w3410 = pi333 & ~w615;
assign w3411 = (w3235 & w17309) | (w3235 & w17310) | (w17309 & w17310);
assign w3412 = w3410 & w17651;
assign w3413 = ~w3411 & ~w3412;
assign w3414 = pi332 & ~w793;
assign w3415 = w3414 & w17652;
assign w3416 = (w3232 & w17312) | (w3232 & w17313) | (w17312 & w17313);
assign w3417 = ~w3415 & ~w3416;
assign w3418 = pi331 & ~w955;
assign w3419 = w3019 & ~w3213;
assign w3420 = ~w3019 & w3213;
assign w3421 = ~w3419 & ~w3420;
assign w3422 = ~w3222 & w3224;
assign w3423 = (w3220 & w3222) | (w3220 & w17314) | (w3222 & w17314);
assign w3424 = pi330 & w1101;
assign w3425 = (~w3424 & w2747) | (~w3424 & w17315) | (w2747 & w17315);
assign w3426 = ~w3423 & ~w3425;
assign w3427 = w1101 & w17316;
assign w3428 = w3421 & w17317;
assign w3429 = ~w1101 & w3422;
assign w3430 = ~w2747 & w17318;
assign w3431 = w1101 & w17319;
assign w3432 = ~w3223 & w3431;
assign w3433 = ~w3421 & w3432;
assign w3434 = ~w3429 & ~w3430;
assign w3435 = ~w3433 & w3434;
assign w3436 = ~w3428 & w3435;
assign w3437 = pi328 & w1602;
assign w3438 = pi327 & ~w1865;
assign w3439 = (w3207 & w17321) | (w3207 & w17322) | (w17321 & w17322);
assign w3440 = ~w3438 & w17653;
assign w3441 = ~w3439 & ~w3440;
assign w3442 = (~w3202 & ~w3204) | (~w3202 & w17323) | (~w3204 & w17323);
assign w3443 = pi326 & ~w2170;
assign w3444 = w3442 & ~w3443;
assign w3445 = ~w3442 & w3443;
assign w3446 = ~w3444 & ~w3445;
assign w3447 = (~w3037 & w3198) | (~w3037 & w17324) | (w3198 & w17324);
assign w3448 = pi325 & ~w2373;
assign w3449 = pi323 & ~w3183;
assign w3450 = pi142 & pi258;
assign w3451 = pi141 & pi259;
assign w3452 = (~w3451 & ~w3166) | (~w3451 & w16567) | (~w3166 & w16567);
assign w3453 = w3166 & w16568;
assign w3454 = ~w3452 & ~w3453;
assign w3455 = ~w3161 & ~w3165;
assign w3456 = pi139 & pi261;
assign w3457 = pi138 & pi262;
assign w3458 = (~w3127 & ~w3129) | (~w3127 & w16382) | (~w3129 & w16382);
assign w3459 = w3116 & w3123;
assign w3460 = ~w3125 & ~w3459;
assign w3461 = (~w3117 & w3049) | (~w3117 & w15857) | (w3049 & w15857);
assign w3462 = ~w3113 & ~w3461;
assign w3463 = pi135 & pi265;
assign w3464 = (~w3107 & w2590) | (~w3107 & w16383) | (w2590 & w16383);
assign w3465 = ~w3050 & w3464;
assign w3466 = ~w3108 & ~w3465;
assign w3467 = pi134 & pi266;
assign w3468 = pi133 & pi267;
assign w3469 = (w3095 & w3056) | (w3095 & w16384) | (w3056 & w16384);
assign w3470 = pi132 & pi268;
assign w3471 = pi131 & pi269;
assign w3472 = pi130 & pi270;
assign w3473 = pi129 & pi271;
assign w3474 = pi128 & pi272;
assign w3475 = (~w3063 & w15858) | (~w3063 & w17724) | (w15858 & w17724);
assign w3476 = w3474 & ~w3475;
assign w3477 = ~w3474 & w17654;
assign w3478 = ~w3476 & w17325;
assign w3479 = (~w3473 & w3476) | (~w3473 & w17326) | (w3476 & w17326);
assign w3480 = ~w3478 & ~w3479;
assign w3481 = w3472 & w3480;
assign w3482 = ~w3472 & ~w3480;
assign w3483 = ~w3481 & ~w3482;
assign w3484 = (w3073 & w17328) | (w3073 & w17329) | (w17328 & w17329);
assign w3485 = ~w3483 & w17655;
assign w3486 = ~w3484 & ~w3485;
assign w3487 = w3471 & w3486;
assign w3488 = ~w3471 & ~w3486;
assign w3489 = ~w3487 & ~w3488;
assign w3490 = w3489 & w17656;
assign w3491 = (w3086 & w17330) | (w3086 & w17331) | (w17330 & w17331);
assign w3492 = ~w3490 & ~w3491;
assign w3493 = ~w3470 & ~w3492;
assign w3494 = w3470 & w3492;
assign w3495 = ~w3493 & ~w3494;
assign w3496 = ~w3469 & w17332;
assign w3497 = (~w3495 & w3469) | (~w3495 & w17333) | (w3469 & w17333);
assign w3498 = ~w3496 & ~w3497;
assign w3499 = w3468 & ~w3498;
assign w3500 = ~w3468 & w3498;
assign w3501 = ~w3499 & ~w3500;
assign w3502 = w3094 & w3101;
assign w3503 = ~w3104 & ~w3502;
assign w3504 = ~w3501 & ~w3503;
assign w3505 = w3501 & w3503;
assign w3506 = ~w3504 & ~w3505;
assign w3507 = ~w3467 & w3506;
assign w3508 = w3467 & ~w3506;
assign w3509 = ~w3507 & ~w3508;
assign w3510 = w3466 & ~w3509;
assign w3511 = ~w3466 & w3509;
assign w3512 = ~w3510 & ~w3511;
assign w3513 = ~w3463 & ~w3512;
assign w3514 = w3463 & w3512;
assign w3515 = ~w3513 & ~w3514;
assign w3516 = w3462 & w3515;
assign w3517 = ~w3462 & ~w3515;
assign w3518 = ~w3516 & ~w3517;
assign w3519 = ~w3125 & w16569;
assign w3520 = (~w3518 & w3125) | (~w3518 & w16570) | (w3125 & w16570);
assign w3521 = ~w3519 & ~w3520;
assign w3522 = pi137 & pi263;
assign w3523 = pi136 & pi264;
assign w3524 = w3522 & ~w3523;
assign w3525 = ~w3522 & w3523;
assign w3526 = ~w3524 & ~w3525;
assign w3527 = w3521 & w3526;
assign w3528 = ~w3521 & ~w3526;
assign w3529 = ~w3527 & ~w3528;
assign w3530 = w3458 & ~w3529;
assign w3531 = ~w3458 & w3529;
assign w3532 = ~w3530 & ~w3531;
assign w3533 = w3457 & ~w3532;
assign w3534 = ~w3457 & w3532;
assign w3535 = ~w3533 & ~w3534;
assign w3536 = ~w3141 & w3145;
assign w3537 = ~w3142 & ~w3536;
assign w3538 = w3535 & ~w3537;
assign w3539 = ~w3535 & w3537;
assign w3540 = ~w3538 & ~w3539;
assign w3541 = ~w3456 & ~w3540;
assign w3542 = w3456 & w3540;
assign w3543 = ~w3541 & ~w3542;
assign w3544 = pi140 & pi260;
assign w3545 = w3144 & w3151;
assign w3546 = ~w3153 & ~w3545;
assign w3547 = w3544 & ~w3546;
assign w3548 = ~w3544 & w3546;
assign w3549 = ~w3547 & ~w3548;
assign w3550 = w3543 & w3549;
assign w3551 = ~w3543 & ~w3549;
assign w3552 = ~w3550 & ~w3551;
assign w3553 = ~w3455 & w3552;
assign w3554 = w3455 & ~w3552;
assign w3555 = ~w3553 & ~w3554;
assign w3556 = w3454 & w3555;
assign w3557 = ~w3454 & ~w3555;
assign w3558 = ~w3556 & ~w3557;
assign w3559 = w3450 & w3558;
assign w3560 = ~w3450 & ~w3558;
assign w3561 = ~w3559 & ~w3560;
assign w3562 = ~w3170 & ~w3178;
assign w3563 = w3561 & w3562;
assign w3564 = w3170 & ~w3179;
assign w3565 = ~w3561 & w3564;
assign w3566 = (~w3562 & ~w3561) | (~w3562 & w16385) | (~w3561 & w16385);
assign w3567 = ~w3565 & w3566;
assign w3568 = ~w3563 & ~w3567;
assign w3569 = (pi322 & w3567) | (pi322 & w16571) | (w3567 & w16571);
assign w3570 = ~w3449 & ~w3569;
assign w3571 = (pi323 & w3567) | (pi323 & w16572) | (w3567 & w16572);
assign w3572 = w3184 & w3571;
assign w3573 = ~w3570 & ~w3572;
assign w3574 = (~w3187 & ~w3188) | (~w3187 & w17334) | (~w3188 & w17334);
assign w3575 = ~w3573 & w3574;
assign w3576 = w3573 & ~w3574;
assign w3577 = ~w3575 & ~w3576;
assign w3578 = pi324 & w2698;
assign w3579 = (~w3193 & ~w3194) | (~w3193 & w17335) | (~w3194 & w17335);
assign w3580 = w3578 & w3579;
assign w3581 = ~w3578 & ~w3579;
assign w3582 = ~w3580 & ~w3581;
assign w3583 = w3577 & ~w3582;
assign w3584 = ~w3577 & w3582;
assign w3585 = ~w3583 & ~w3584;
assign w3586 = w3448 & ~w3585;
assign w3587 = ~w3448 & w3585;
assign w3588 = ~w3586 & ~w3587;
assign w3589 = w3447 & ~w3588;
assign w3590 = ~w3447 & w3588;
assign w3591 = ~w3589 & ~w3590;
assign w3592 = ~w3446 & w3591;
assign w3593 = w3446 & ~w3591;
assign w3594 = ~w3592 & ~w3593;
assign w3595 = ~w3441 & w3594;
assign w3596 = w3441 & ~w3594;
assign w3597 = ~w3595 & ~w3596;
assign w3598 = ~w3437 & ~w3597;
assign w3599 = w3437 & w3597;
assign w3600 = ~w3598 & ~w3599;
assign w3601 = (~w3026 & ~w3210) | (~w3026 & w17336) | (~w3210 & w17336);
assign w3602 = w3600 & ~w3601;
assign w3603 = ~w3600 & w3601;
assign w3604 = ~w3602 & ~w3603;
assign w3605 = pi329 & w1339;
assign w3606 = (~w3220 & ~w3213) | (~w3220 & w17337) | (~w3213 & w17337);
assign w3607 = ~w3419 & ~w3606;
assign w3608 = ~w3605 & ~w3607;
assign w3609 = w3605 & w3607;
assign w3610 = ~w3608 & ~w3609;
assign w3611 = w3604 & ~w3610;
assign w3612 = ~w3604 & w3610;
assign w3613 = ~w3611 & ~w3612;
assign w3614 = w3436 & w3613;
assign w3615 = ~w3436 & ~w3613;
assign w3616 = ~w3614 & ~w3615;
assign w3617 = ~w3018 & w3023;
assign w3618 = w3018 & ~w3023;
assign w3619 = w3229 & w3421;
assign w3620 = ~w3229 & ~w3421;
assign w3621 = ~w3619 & ~w3620;
assign w3622 = (~w3617 & w3621) | (~w3617 & w17338) | (w3621 & w17338);
assign w3623 = w3616 & ~w3622;
assign w3624 = ~w3616 & w3622;
assign w3625 = ~w3623 & ~w3624;
assign w3626 = w3418 & w3625;
assign w3627 = ~w3418 & ~w3625;
assign w3628 = ~w3626 & ~w3627;
assign w3629 = w3417 & ~w3628;
assign w3630 = ~w3417 & w3628;
assign w3631 = ~w3629 & ~w3630;
assign w3632 = w3413 & ~w3631;
assign w3633 = ~w3413 & w3631;
assign w3634 = ~w3632 & ~w3633;
assign w3635 = ~w3409 & w3634;
assign w3636 = w3409 & ~w3634;
assign w3637 = ~w3635 & ~w3636;
assign w3638 = w3247 & ~w3637;
assign w3639 = ~w3247 & w3637;
assign w3640 = ~w3638 & ~w3639;
assign w3641 = w3403 & w3640;
assign w3642 = ~w3403 & ~w3640;
assign w3643 = ~w3641 & ~w3642;
assign w3644 = w3402 & w3643;
assign w3645 = ~w3402 & ~w3643;
assign w3646 = ~w3644 & ~w3645;
assign w3647 = pi272 & ~w3646;
assign w3648 = ~pi272 & w3646;
assign w3649 = ~w3647 & ~w3648;
assign w3650 = w3401 & ~w3649;
assign w3651 = ~w3401 & w3649;
assign w3652 = ~w3650 & ~w3651;
assign w3653 = ~w3400 & w3652;
assign w3654 = w3400 & ~w3652;
assign w3655 = ~w3653 & ~w3654;
assign w3656 = (~w3258 & ~w3260) | (~w3258 & w17339) | (~w3260 & w17339);
assign w3657 = w3655 & ~w3656;
assign w3658 = (~w135 & w3655) | (~w135 & w17340) | (w3655 & w17340);
assign w3659 = ~w3657 & w3658;
assign w3660 = (pi161 & ~w135) | (pi161 & w17341) | (~w135 & w17341);
assign w3661 = ~w3659 & w3660;
assign w3662 = ~pi160 & ~w3268;
assign w3663 = ~w3661 & w3662;
assign w3664 = ~pi079 & ~pi161;
assign w3665 = pi128 & pi306;
assign w3666 = pi307 & w464;
assign w3667 = (~w3666 & ~w3397) | (~w3666 & w17342) | (~w3397 & w17342);
assign w3668 = w3397 & w17343;
assign w3669 = ~w3667 & ~w3668;
assign w3670 = pi308 & ~w653;
assign w3671 = ~w3670 & w17657;
assign w3672 = (w3394 & w17345) | (w3394 & w17346) | (w17345 & w17346);
assign w3673 = ~w3671 & ~w3672;
assign w3674 = pi309 & w709;
assign w3675 = pi310 & w698;
assign w3676 = (~w3376 & ~w3378) | (~w3376 & w17347) | (~w3378 & w17347);
assign w3677 = w3675 & ~w3676;
assign w3678 = ~w3675 & w3676;
assign w3679 = ~w3677 & ~w3678;
assign w3680 = (~w3370 & ~w3372) | (~w3370 & w17348) | (~w3372 & w17348);
assign w3681 = pi311 & w855;
assign w3682 = (~w3364 & ~w3365) | (~w3364 & w17349) | (~w3365 & w17349);
assign w3683 = pi312 & w1159;
assign w3684 = ~w3682 & w3683;
assign w3685 = w3682 & ~w3683;
assign w3686 = ~w3684 & ~w3685;
assign w3687 = w1419 & w17350;
assign w3688 = (~w3349 & ~w3351) | (~w3349 & w17351) | (~w3351 & w17351);
assign w3689 = w3687 & ~w3688;
assign w3690 = ~w3687 & w3688;
assign w3691 = ~w3689 & ~w3690;
assign w3692 = w1692 & w17352;
assign w3693 = (~w3282 & ~w3283) | (~w3282 & w17353) | (~w3283 & w17353);
assign w3694 = ~w3692 & w3693;
assign w3695 = w3692 & ~w3693;
assign w3696 = ~w3694 & ~w3695;
assign w3697 = pi316 & w1954;
assign w3698 = pi317 & ~w2473;
assign w3699 = pi318 & w2801;
assign w3700 = (~w3316 & ~w3318) | (~w3316 & w17354) | (~w3318 & w17354);
assign w3701 = pi319 & w2925;
assign w3702 = (~w3291 & ~w3292) | (~w3291 & w17355) | (~w3292 & w17355);
assign w3703 = pi320 & w3304;
assign w3704 = pi142 & ~pi143;
assign w3705 = ~pi142 & pi143;
assign w3706 = ~w3704 & ~w3705;
assign w3707 = (~w3300 & ~w3301) | (~w3300 & w17356) | (~w3301 & w17356);
assign w3708 = w3706 & w3707;
assign w3709 = ~w3706 & ~w3707;
assign w3710 = ~w3708 & ~w3709;
assign w3711 = pi321 & w3710;
assign w3712 = (~w3308 & ~w3309) | (~w3308 & w17357) | (~w3309 & w17357);
assign w3713 = ~w3711 & w3712;
assign w3714 = w3711 & ~w3712;
assign w3715 = ~w3713 & ~w3714;
assign w3716 = w3703 & w3715;
assign w3717 = ~w3703 & ~w3715;
assign w3718 = ~w3716 & ~w3717;
assign w3719 = w3702 & ~w3718;
assign w3720 = ~w3702 & w3718;
assign w3721 = ~w3719 & ~w3720;
assign w3722 = w3701 & w3721;
assign w3723 = ~w3701 & ~w3721;
assign w3724 = ~w3722 & ~w3723;
assign w3725 = ~w3700 & ~w3724;
assign w3726 = w3700 & w3724;
assign w3727 = ~w3725 & ~w3726;
assign w3728 = w3699 & ~w3727;
assign w3729 = ~w3699 & w3727;
assign w3730 = ~w3728 & ~w3729;
assign w3731 = w3698 & ~w3730;
assign w3732 = ~w3698 & w3730;
assign w3733 = ~w3731 & ~w3732;
assign w3734 = w3321 & ~w3327;
assign w3735 = (~w3324 & w2948) | (~w3324 & w17359) | (w2948 & w17359);
assign w3736 = w2949 & ~w3321;
assign w3737 = (~w3736 & w3734) | (~w3736 & w17360) | (w3734 & w17360);
assign w3738 = w3733 & ~w3737;
assign w3739 = ~w3733 & w3737;
assign w3740 = ~w3738 & ~w3739;
assign w3741 = (~w3340 & ~w3342) | (~w3340 & w17361) | (~w3342 & w17361);
assign w3742 = w3740 & w3741;
assign w3743 = ~w3740 & ~w3741;
assign w3744 = ~w3742 & ~w3743;
assign w3745 = w3697 & w3744;
assign w3746 = ~w3697 & ~w3744;
assign w3747 = ~w3745 & ~w3746;
assign w3748 = ~w3696 & ~w3747;
assign w3749 = w3696 & w3747;
assign w3750 = ~w3748 & ~w3749;
assign w3751 = w3691 & w3750;
assign w3752 = ~w3691 & ~w3750;
assign w3753 = ~w3751 & ~w3752;
assign w3754 = pi313 & w1220;
assign w3755 = ~w3753 & ~w3754;
assign w3756 = w3753 & w3754;
assign w3757 = ~w3755 & ~w3756;
assign w3758 = (~w3357 & ~w3359) | (~w3357 & w17362) | (~w3359 & w17362);
assign w3759 = ~w3757 & w3758;
assign w3760 = w3757 & ~w3758;
assign w3761 = ~w3759 & ~w3760;
assign w3762 = w3686 & w3761;
assign w3763 = ~w3686 & ~w3761;
assign w3764 = ~w3762 & ~w3763;
assign w3765 = ~w3681 & ~w3764;
assign w3766 = w3681 & w3764;
assign w3767 = ~w3765 & ~w3766;
assign w3768 = w3680 & ~w3767;
assign w3769 = ~w3680 & w3767;
assign w3770 = ~w3768 & ~w3769;
assign w3771 = w3679 & ~w3770;
assign w3772 = ~w3679 & w3770;
assign w3773 = ~w3771 & ~w3772;
assign w3774 = ~w3674 & w3773;
assign w3775 = w3674 & ~w3773;
assign w3776 = ~w3774 & ~w3775;
assign w3777 = ~w653 & ~w3000;
assign w3778 = (w3777 & w2997) | (w3777 & w17363) | (w2997 & w17363);
assign w3779 = ~w3392 & ~w3778;
assign w3780 = ~w3776 & w3779;
assign w3781 = w3776 & ~w3779;
assign w3782 = ~w3780 & ~w3781;
assign w3783 = ~w3673 & w3782;
assign w3784 = w3673 & ~w3782;
assign w3785 = ~w3783 & ~w3784;
assign w3786 = w3669 & ~w3785;
assign w3787 = ~w3669 & w3785;
assign w3788 = ~w3786 & ~w3787;
assign w3789 = w3665 & w3788;
assign w3790 = ~w3665 & ~w3788;
assign w3791 = ~w3789 & ~w3790;
assign w3792 = pi337 & w456;
assign w3793 = ~w465 & w17364;
assign w3794 = (~w3793 & ~w3643) | (~w3793 & w17365) | (~w3643 & w17365);
assign w3795 = w3643 & w17366;
assign w3796 = ~w3794 & ~w3795;
assign w3797 = (pi335 & ~w536) | (pi335 & w17367) | (~w536 & w17367);
assign w3798 = (~w3638 & ~w3640) | (~w3638 & w17368) | (~w3640 & w17368);
assign w3799 = w3797 & ~w3798;
assign w3800 = ~w3797 & w3798;
assign w3801 = ~w3799 & ~w3800;
assign w3802 = pi334 & ~w615;
assign w3803 = ~w3802 & w17658;
assign w3804 = (w3634 & w17370) | (w3634 & w17371) | (w17370 & w17371);
assign w3805 = ~w3803 & ~w3804;
assign w3806 = pi333 & ~w793;
assign w3807 = w3806 & w17659;
assign w3808 = (w3631 & w17373) | (w3631 & w17374) | (w17373 & w17374);
assign w3809 = ~w3807 & ~w3808;
assign w3810 = pi332 & ~w955;
assign w3811 = ~w3810 & w17660;
assign w3812 = (w3628 & w17376) | (w3628 & w17377) | (w17376 & w17377);
assign w3813 = ~w3811 & ~w3812;
assign w3814 = pi330 & w1339;
assign w3815 = (~w3422 & ~w3621) | (~w3422 & w17378) | (~w3621 & w17378);
assign w3816 = ~w3613 & w17379;
assign w3817 = (w3814 & w3613) | (w3814 & w17380) | (w3613 & w17380);
assign w3818 = ~w3424 & ~w3817;
assign w3819 = w1101 & w1339;
assign w3820 = (w3819 & ~w3613) | (w3819 & w17381) | (~w3613 & w17381);
assign w3821 = w3613 & w17382;
assign w3822 = ~w3820 & ~w3821;
assign w3823 = ~w3818 & w3822;
assign w3824 = ~w3816 & ~w3823;
assign w3825 = pi329 & w1602;
assign w3826 = (w3604 & w17384) | (w3604 & w17385) | (w17384 & w17385);
assign w3827 = ~w3825 & w17661;
assign w3828 = ~w3826 & ~w3827;
assign w3829 = pi328 & ~w1865;
assign w3830 = (~w3599 & ~w3600) | (~w3599 & w17386) | (~w3600 & w17386);
assign w3831 = w3829 & ~w3830;
assign w3832 = ~w3829 & w3830;
assign w3833 = ~w3831 & ~w3832;
assign w3834 = pi327 & ~w2170;
assign w3835 = (w3594 & w17388) | (w3594 & w17389) | (w17388 & w17389);
assign w3836 = w3834 & w17662;
assign w3837 = ~w3835 & ~w3836;
assign w3838 = pi325 & w2698;
assign w3839 = pi324 & ~w3183;
assign w3840 = (w3577 & w17391) | (w3577 & w17392) | (w17391 & w17392);
assign w3841 = ~w3839 & w17663;
assign w3842 = ~w3840 & ~w3841;
assign w3843 = pi143 & pi258;
assign w3844 = pi142 & pi259;
assign w3845 = (~w3844 & ~w3558) | (~w3844 & w16573) | (~w3558 & w16573);
assign w3846 = w3558 & w16574;
assign w3847 = ~w3845 & ~w3846;
assign w3848 = pi140 & pi261;
assign w3849 = (~w3533 & ~w3535) | (~w3533 & w15860) | (~w3535 & w15860);
assign w3850 = pi137 & pi264;
assign w3851 = pi136 & pi265;
assign w3852 = ~w3113 & ~w3513;
assign w3853 = (~w3514 & ~w3852) | (~w3514 & w15861) | (~w3852 & w15861);
assign w3854 = pi135 & pi266;
assign w3855 = pi134 & pi267;
assign w3856 = (~w3500 & ~w3503) | (~w3500 & w16575) | (~w3503 & w16575);
assign w3857 = (~w3493 & w3469) | (~w3493 & w17393) | (w3469 & w17393);
assign w3858 = (~w3469 & w17394) | (~w3469 & w17395) | (w17394 & w17395);
assign w3859 = pi131 & pi270;
assign w3860 = ~w3481 & ~w3484;
assign w3861 = pi129 & pi272;
assign w3862 = pi128 & pi273;
assign w3863 = ~w3861 & ~w3862;
assign w3864 = pi129 & pi273;
assign w3865 = w3474 & w3864;
assign w3866 = ~w3863 & ~w3865;
assign w3867 = pi130 & w3866;
assign w3868 = w529 & ~w3866;
assign w3869 = ~w3867 & ~w3868;
assign w3870 = pi271 & ~w3869;
assign w3871 = (w3870 & w3478) | (w3870 & w17396) | (w3478 & w17396);
assign w3872 = pi130 & pi271;
assign w3873 = ~w3866 & ~w3872;
assign w3874 = w3477 & ~w3867;
assign w3875 = (~w3473 & w3869) | (~w3473 & w17397) | (w3869 & w17397);
assign w3876 = (w3875 & w3475) | (w3875 & w17398) | (w3475 & w17398);
assign w3877 = ~w3874 & ~w3876;
assign w3878 = ~w3475 & w17399;
assign w3879 = (~w3878 & w3877) | (~w3878 & w17400) | (w3877 & w17400);
assign w3880 = ~w3871 & w3879;
assign w3881 = ~w3860 & w3880;
assign w3882 = w3860 & ~w3880;
assign w3883 = ~w3881 & ~w3882;
assign w3884 = w3859 & ~w3883;
assign w3885 = ~w3859 & w3883;
assign w3886 = ~w3884 & ~w3885;
assign w3887 = ~w3490 & w17401;
assign w3888 = (w3886 & w3490) | (w3886 & w17402) | (w3490 & w17402);
assign w3889 = ~w3887 & ~w3888;
assign w3890 = ~w3858 & w3889;
assign w3891 = ~w3494 & ~w3889;
assign w3892 = ~w3857 & w3891;
assign w3893 = ~w3890 & ~w3892;
assign w3894 = pi133 & pi268;
assign w3895 = pi132 & pi269;
assign w3896 = w3894 & ~w3895;
assign w3897 = ~w3894 & w3895;
assign w3898 = ~w3896 & ~w3897;
assign w3899 = w3893 & w3898;
assign w3900 = ~w3893 & ~w3898;
assign w3901 = ~w3899 & ~w3900;
assign w3902 = w3856 & ~w3901;
assign w3903 = ~w3856 & w3901;
assign w3904 = ~w3902 & ~w3903;
assign w3905 = ~w3855 & ~w3904;
assign w3906 = w3855 & w3904;
assign w3907 = ~w3905 & ~w3906;
assign w3908 = (~w3508 & w3466) | (~w3508 & w16129) | (w3466 & w16129);
assign w3909 = w3907 & ~w3908;
assign w3910 = ~w3907 & w3908;
assign w3911 = ~w3909 & ~w3910;
assign w3912 = w3854 & w3911;
assign w3913 = ~w3854 & ~w3911;
assign w3914 = ~w3912 & ~w3913;
assign w3915 = ~w3853 & w3914;
assign w3916 = w3853 & ~w3914;
assign w3917 = ~w3915 & ~w3916;
assign w3918 = ~w3851 & ~w3917;
assign w3919 = w3851 & w3917;
assign w3920 = ~w3918 & ~w3919;
assign w3921 = w3518 & w3523;
assign w3922 = ~w3518 & ~w3523;
assign w3923 = (~w3921 & w3460) | (~w3921 & w15863) | (w3460 & w15863);
assign w3924 = w3920 & ~w3923;
assign w3925 = ~w3920 & w3923;
assign w3926 = ~w3924 & ~w3925;
assign w3927 = ~w3850 & ~w3926;
assign w3928 = w3850 & w3926;
assign w3929 = ~w3927 & ~w3928;
assign w3930 = (w3522 & ~w3529) | (w3522 & w16386) | (~w3529 & w16386);
assign w3931 = ~w3521 & ~w3523;
assign w3932 = w3521 & w3523;
assign w3933 = ~w3931 & ~w3932;
assign w3934 = w3458 & ~w3933;
assign w3935 = ~w3930 & ~w3934;
assign w3936 = w3929 & ~w3935;
assign w3937 = ~w3929 & w3935;
assign w3938 = ~w3936 & ~w3937;
assign w3939 = w3849 & ~w3938;
assign w3940 = ~w3849 & w3938;
assign w3941 = ~w3939 & ~w3940;
assign w3942 = pi139 & pi262;
assign w3943 = pi138 & pi263;
assign w3944 = w3942 & ~w3943;
assign w3945 = ~w3942 & w3943;
assign w3946 = ~w3944 & ~w3945;
assign w3947 = w3941 & w3946;
assign w3948 = ~w3941 & ~w3946;
assign w3949 = ~w3947 & ~w3948;
assign w3950 = ~w3541 & ~w3546;
assign w3951 = ~w3542 & ~w3950;
assign w3952 = ~w3949 & ~w3951;
assign w3953 = w3949 & w3951;
assign w3954 = ~w3952 & ~w3953;
assign w3955 = ~w3848 & ~w3954;
assign w3956 = w3848 & w3954;
assign w3957 = ~w3955 & ~w3956;
assign w3958 = w3544 & ~w3552;
assign w3959 = ~w3553 & ~w3958;
assign w3960 = ~w3957 & ~w3959;
assign w3961 = w3957 & w3959;
assign w3962 = ~w3960 & ~w3961;
assign w3963 = pi141 & pi260;
assign w3964 = (w3555 & w16576) | (w3555 & w16577) | (w16576 & w16577);
assign w3965 = (~w3555 & w16578) | (~w3555 & w16579) | (w16578 & w16579);
assign w3966 = ~w3964 & ~w3965;
assign w3967 = w3962 & ~w3966;
assign w3968 = ~w3962 & w3966;
assign w3969 = ~w3967 & ~w3968;
assign w3970 = w3847 & w3969;
assign w3971 = ~w3847 & ~w3969;
assign w3972 = ~w3970 & ~w3971;
assign w3973 = w3843 & w3972;
assign w3974 = ~w3843 & ~w3972;
assign w3975 = ~w3973 & ~w3974;
assign w3976 = ~w3563 & ~w3565;
assign w3977 = w3975 & ~w3976;
assign w3978 = ~w3975 & w3976;
assign w3979 = ~w3977 & ~w3978;
assign w3980 = (~w3571 & ~w3979) | (~w3571 & w17403) | (~w3979 & w17403);
assign w3981 = w3979 & w17404;
assign w3982 = ~w3980 & ~w3981;
assign w3983 = (~w3572 & ~w3573) | (~w3572 & w17405) | (~w3573 & w17405);
assign w3984 = ~w3982 & w3983;
assign w3985 = w3982 & ~w3983;
assign w3986 = ~w3984 & ~w3985;
assign w3987 = w3842 & w3986;
assign w3988 = ~w3842 & ~w3986;
assign w3989 = ~w3987 & ~w3988;
assign w3990 = w3838 & w3989;
assign w3991 = ~w3838 & ~w3989;
assign w3992 = ~w3990 & ~w3991;
assign w3993 = (~w3586 & ~w3588) | (~w3586 & w17406) | (~w3588 & w17406);
assign w3994 = w3992 & ~w3993;
assign w3995 = ~w3992 & w3993;
assign w3996 = ~w3994 & ~w3995;
assign w3997 = pi326 & ~w2373;
assign w3998 = (w3591 & w17408) | (w3591 & w17409) | (w17408 & w17409);
assign w3999 = ~w3997 & w17664;
assign w4000 = ~w3998 & ~w3999;
assign w4001 = ~w3996 & ~w4000;
assign w4002 = w3996 & w4000;
assign w4003 = ~w4001 & ~w4002;
assign w4004 = w3837 & w4003;
assign w4005 = ~w3837 & ~w4003;
assign w4006 = ~w4004 & ~w4005;
assign w4007 = w3833 & ~w4006;
assign w4008 = ~w3833 & w4006;
assign w4009 = ~w4007 & ~w4008;
assign w4010 = w3828 & w4009;
assign w4011 = ~w3828 & ~w4009;
assign w4012 = ~w4010 & ~w4011;
assign w4013 = ~w3824 & ~w4012;
assign w4014 = w3824 & w4012;
assign w4015 = ~w4013 & ~w4014;
assign w4016 = pi331 & w1101;
assign w4017 = (~w3623 & ~w3625) | (~w3623 & w17410) | (~w3625 & w17410);
assign w4018 = w4016 & ~w4017;
assign w4019 = ~w4016 & w4017;
assign w4020 = ~w4018 & ~w4019;
assign w4021 = w4015 & w4020;
assign w4022 = ~w4015 & ~w4020;
assign w4023 = ~w4021 & ~w4022;
assign w4024 = w3813 & ~w4023;
assign w4025 = ~w3813 & w4023;
assign w4026 = ~w4024 & ~w4025;
assign w4027 = w3809 & ~w4026;
assign w4028 = ~w3809 & w4026;
assign w4029 = ~w4027 & ~w4028;
assign w4030 = w3805 & w4029;
assign w4031 = ~w3805 & ~w4029;
assign w4032 = ~w4030 & ~w4031;
assign w4033 = w3801 & w4032;
assign w4034 = ~w3801 & ~w4032;
assign w4035 = ~w4033 & ~w4034;
assign w4036 = w3796 & w4035;
assign w4037 = ~w3796 & ~w4035;
assign w4038 = ~w4036 & ~w4037;
assign w4039 = w3792 & w4038;
assign w4040 = ~w3792 & ~w4038;
assign w4041 = ~w4039 & ~w4040;
assign w4042 = (~w3647 & ~w3649) | (~w3647 & w17411) | (~w3649 & w17411);
assign w4043 = ~w4041 & ~w4042;
assign w4044 = w4041 & w4042;
assign w4045 = ~w4043 & ~w4044;
assign w4046 = pi273 & w4045;
assign w4047 = ~pi273 & ~w4045;
assign w4048 = ~w4046 & ~w4047;
assign w4049 = (~w3656 & w3652) | (~w3656 & w17412) | (w3652 & w17412);
assign w4050 = ~w3653 & ~w4049;
assign w4051 = w4048 & ~w4050;
assign w4052 = ~w4048 & w4050;
assign w4053 = ~w4051 & ~w4052;
assign w4054 = w3791 & ~w4053;
assign w4055 = (~w135 & ~w4053) | (~w135 & w17413) | (~w4053 & w17413);
assign w4056 = ~w4054 & w4055;
assign w4057 = (pi161 & ~w135) | (pi161 & w17414) | (~w135 & w17414);
assign w4058 = ~w4056 & w4057;
assign w4059 = ~pi160 & ~w3664;
assign w4060 = ~w4058 & w4059;
assign w4061 = ~pi080 & ~pi161;
assign w4062 = (~w4043 & ~w4045) | (~w4043 & w17415) | (~w4045 & w17415);
assign w4063 = pi274 & ~w4062;
assign w4064 = ~pi274 & w4062;
assign w4065 = ~w4063 & ~w4064;
assign w4066 = pi338 & w456;
assign w4067 = (pi336 & ~w536) | (pi336 & w17416) | (~w536 & w17416);
assign w4068 = (~w3795 & ~w4035) | (~w3795 & w17417) | (~w4035 & w17417);
assign w4069 = ~w4067 & w4068;
assign w4070 = ~w537 & ~w4068;
assign w4071 = ~w4069 & ~w4070;
assign w4072 = pi335 & ~w615;
assign w4073 = (~w3799 & ~w3801) | (~w3799 & w17418) | (~w3801 & w17418);
assign w4074 = w4072 & ~w4073;
assign w4075 = ~w4072 & w4073;
assign w4076 = ~w4074 & ~w4075;
assign w4077 = (~w3807 & w4026) | (~w3807 & w17419) | (w4026 & w17419);
assign w4078 = pi333 & ~w955;
assign w4079 = ~w4077 & w4078;
assign w4080 = w4077 & ~w4078;
assign w4081 = ~w4079 & ~w4080;
assign w4082 = pi332 & w1101;
assign w4083 = (~w3811 & w4023) | (~w3811 & w17420) | (w4023 & w17420);
assign w4084 = w4082 & w4083;
assign w4085 = ~w4082 & ~w4083;
assign w4086 = ~w4084 & ~w4085;
assign w4087 = pi329 & ~w1865;
assign w4088 = (~w3827 & ~w4009) | (~w3827 & w17421) | (~w4009 & w17421);
assign w4089 = w4087 & w4088;
assign w4090 = ~w4087 & ~w4088;
assign w4091 = ~w4089 & ~w4090;
assign w4092 = pi328 & ~w2170;
assign w4093 = (~w3832 & ~w3833) | (~w3832 & w17422) | (~w3833 & w17422);
assign w4094 = w4092 & w4093;
assign w4095 = ~w4092 & ~w4093;
assign w4096 = ~w4094 & ~w4095;
assign w4097 = pi327 & ~w2373;
assign w4098 = ~w4097 & w17665;
assign w4099 = (w4003 & w17424) | (w4003 & w17425) | (w17424 & w17425);
assign w4100 = ~w4098 & ~w4099;
assign w4101 = (~w3998 & ~w3996) | (~w3998 & w17426) | (~w3996 & w17426);
assign w4102 = pi326 & w2698;
assign w4103 = pi325 & ~w3183;
assign w4104 = pi323 & w3979;
assign w4105 = (~w3846 & ~w3969) | (~w3846 & w17427) | (~w3969 & w17427);
assign w4106 = pi141 & pi261;
assign w4107 = (~w3955 & ~w3957) | (~w3955 & w16387) | (~w3957 & w16387);
assign w4108 = pi139 & pi263;
assign w4109 = (~w3943 & w3849) | (~w3943 & w16388) | (w3849 & w16388);
assign w4110 = ~w3939 & ~w4109;
assign w4111 = pi138 & pi264;
assign w4112 = ~w3928 & ~w3934;
assign w4113 = (~w3927 & ~w4112) | (~w3927 & w16389) | (~w4112 & w16389);
assign w4114 = pi135 & pi267;
assign w4115 = pi134 & pi268;
assign w4116 = pi133 & pi269;
assign w4117 = pi132 & pi270;
assign w4118 = pi131 & pi271;
assign w4119 = pi130 & pi272;
assign w4120 = ~pi271 & ~pi273;
assign w4121 = w3861 & ~w4120;
assign w4122 = ~w4121 & w17654;
assign w4123 = pi271 & w3862;
assign w4124 = ~w3474 & ~w4123;
assign w4125 = pi128 & pi274;
assign w4126 = ~w3864 & ~w4125;
assign w4127 = w3864 & w4125;
assign w4128 = ~w4126 & ~w4127;
assign w4129 = ~w4122 & w17428;
assign w4130 = (w4128 & w4122) | (w4128 & w17429) | (w4122 & w17429);
assign w4131 = ~w4129 & ~w4130;
assign w4132 = w4119 & ~w4131;
assign w4133 = ~w4119 & w4131;
assign w4134 = ~w4132 & ~w4133;
assign w4135 = ~w3478 & w17430;
assign w4136 = (w3866 & w3478) | (w3866 & w17431) | (w3478 & w17431);
assign w4137 = ~w4135 & ~w4136;
assign w4138 = ~w3872 & ~w4137;
assign w4139 = w3872 & w4137;
assign w4140 = (~w4138 & ~w3860) | (~w4138 & w17432) | (~w3860 & w17432);
assign w4141 = w4134 & w4140;
assign w4142 = (w3860 & w17433) | (w3860 & w17434) | (w17433 & w17434);
assign w4143 = ~w4141 & w17435;
assign w4144 = (~w4118 & w4141) | (~w4118 & w17436) | (w4141 & w17436);
assign w4145 = ~w4143 & ~w4144;
assign w4146 = ~w3884 & ~w3888;
assign w4147 = ~w4145 & w4146;
assign w4148 = w4145 & ~w4146;
assign w4149 = ~w4147 & ~w4148;
assign w4150 = w4117 & w4149;
assign w4151 = ~w4117 & ~w4149;
assign w4152 = ~w4150 & ~w4151;
assign w4153 = (w3895 & w3857) | (w3895 & w15865) | (w3857 & w15865);
assign w4154 = ~w3890 & ~w4153;
assign w4155 = w4152 & w4154;
assign w4156 = ~w4152 & ~w4154;
assign w4157 = ~w4155 & ~w4156;
assign w4158 = ~w4116 & w4157;
assign w4159 = w4116 & ~w4157;
assign w4160 = ~w4158 & ~w4159;
assign w4161 = w3894 & w3901;
assign w4162 = ~w3902 & ~w4161;
assign w4163 = w4160 & ~w4162;
assign w4164 = ~w4160 & w4162;
assign w4165 = ~w4163 & ~w4164;
assign w4166 = w4115 & w4165;
assign w4167 = ~w4115 & ~w4165;
assign w4168 = ~w4166 & ~w4167;
assign w4169 = (~w3906 & w3908) | (~w3906 & w16580) | (w3908 & w16580);
assign w4170 = w4168 & ~w4169;
assign w4171 = ~w4168 & w4169;
assign w4172 = ~w4170 & ~w4171;
assign w4173 = ~w4114 & ~w4172;
assign w4174 = w4114 & w4172;
assign w4175 = ~w4173 & ~w4174;
assign w4176 = (~w3912 & w3853) | (~w3912 & w17437) | (w3853 & w17437);
assign w4177 = ~w4175 & w4176;
assign w4178 = w4175 & ~w4176;
assign w4179 = ~w4177 & ~w4178;
assign w4180 = ~w3919 & w17666;
assign w4181 = w4179 & w17667;
assign w4182 = ~w4180 & ~w4181;
assign w4183 = pi137 & pi265;
assign w4184 = pi136 & pi266;
assign w4185 = w4183 & ~w4184;
assign w4186 = ~w4183 & w4184;
assign w4187 = ~w4185 & ~w4186;
assign w4188 = w4182 & w4187;
assign w4189 = ~w4182 & ~w4187;
assign w4190 = ~w4188 & ~w4189;
assign w4191 = w4113 & ~w4190;
assign w4192 = ~w4113 & w4190;
assign w4193 = ~w4191 & ~w4192;
assign w4194 = w4111 & w4193;
assign w4195 = ~w4111 & ~w4193;
assign w4196 = ~w4194 & ~w4195;
assign w4197 = w4110 & w4196;
assign w4198 = ~w4110 & ~w4196;
assign w4199 = ~w4197 & ~w4198;
assign w4200 = ~w4108 & ~w4199;
assign w4201 = w4108 & w4199;
assign w4202 = ~w4200 & ~w4201;
assign w4203 = pi140 & pi262;
assign w4204 = w3942 & w3949;
assign w4205 = ~w3952 & ~w4204;
assign w4206 = w4203 & ~w4205;
assign w4207 = ~w4203 & w4205;
assign w4208 = ~w4206 & ~w4207;
assign w4209 = w4202 & w4208;
assign w4210 = ~w4202 & ~w4208;
assign w4211 = ~w4209 & ~w4210;
assign w4212 = w4107 & w4211;
assign w4213 = ~w4107 & ~w4211;
assign w4214 = ~w4212 & ~w4213;
assign w4215 = ~w4106 & ~w4214;
assign w4216 = w4106 & w4214;
assign w4217 = ~w4215 & ~w4216;
assign w4218 = (~w3964 & w3962) | (~w3964 & w17438) | (w3962 & w17438);
assign w4219 = ~w4217 & w4218;
assign w4220 = w4217 & ~w4218;
assign w4221 = ~w4219 & ~w4220;
assign w4222 = w4105 & ~w4221;
assign w4223 = pi142 & pi260;
assign w4224 = (~w4223 & ~w4221) | (~w4223 & w16390) | (~w4221 & w16390);
assign w4225 = ~w4222 & w4224;
assign w4226 = ~w4221 & w16391;
assign w4227 = ~w4105 & w4223;
assign w4228 = w4221 & w4227;
assign w4229 = ~w4226 & ~w4228;
assign w4230 = ~w4225 & w4229;
assign w4231 = pi144 & pi258;
assign w4232 = pi143 & pi259;
assign w4233 = (~w4232 & ~w3972) | (~w4232 & w16582) | (~w3972 & w16582);
assign w4234 = w3972 & w16583;
assign w4235 = ~w4233 & ~w4234;
assign w4236 = ~w4231 & w4235;
assign w4237 = w4231 & ~w4235;
assign w4238 = ~w4236 & ~w4237;
assign w4239 = w4230 & w4238;
assign w4240 = ~w4230 & ~w4238;
assign w4241 = ~w4239 & ~w4240;
assign w4242 = w3561 & ~w3562;
assign w4243 = (~w3564 & ~w3561) | (~w3564 & w17439) | (~w3561 & w17439);
assign w4244 = w3561 & w3975;
assign w4245 = (~w3565 & w3975) | (~w3565 & w17440) | (w3975 & w17440);
assign w4246 = ~w4244 & w4245;
assign w4247 = w4241 & w4246;
assign w4248 = (pi322 & w4241) | (pi322 & w16584) | (w4241 & w16584);
assign w4249 = ~w4247 & w4248;
assign w4250 = ~w4104 & ~w4249;
assign w4251 = w4104 & w4249;
assign w4252 = ~w4250 & ~w4251;
assign w4253 = (~w3981 & ~w3982) | (~w3981 & w17441) | (~w3982 & w17441);
assign w4254 = ~w4252 & w4253;
assign w4255 = w4252 & ~w4253;
assign w4256 = ~w4254 & ~w4255;
assign w4257 = (pi324 & w3567) | (pi324 & w17442) | (w3567 & w17442);
assign w4258 = ~w4257 & w17668;
assign w4259 = (w3986 & w17444) | (w3986 & w17445) | (w17444 & w17445);
assign w4260 = ~w4258 & ~w4259;
assign w4261 = w4256 & w4260;
assign w4262 = ~w4256 & ~w4260;
assign w4263 = ~w4261 & ~w4262;
assign w4264 = w4103 & w4263;
assign w4265 = ~w4103 & ~w4263;
assign w4266 = ~w4264 & ~w4265;
assign w4267 = (~w3990 & ~w3992) | (~w3990 & w17446) | (~w3992 & w17446);
assign w4268 = w4266 & ~w4267;
assign w4269 = ~w4266 & w4267;
assign w4270 = ~w4268 & ~w4269;
assign w4271 = w4102 & w4270;
assign w4272 = ~w4102 & ~w4270;
assign w4273 = ~w4271 & ~w4272;
assign w4274 = w4101 & ~w4273;
assign w4275 = ~w4101 & w4273;
assign w4276 = ~w4274 & ~w4275;
assign w4277 = w4100 & w4276;
assign w4278 = ~w4100 & ~w4276;
assign w4279 = ~w4277 & ~w4278;
assign w4280 = w4096 & w4279;
assign w4281 = ~w4096 & ~w4279;
assign w4282 = ~w4280 & ~w4281;
assign w4283 = w4091 & ~w4282;
assign w4284 = ~w4091 & w4282;
assign w4285 = ~w4283 & ~w4284;
assign w4286 = w3814 & ~w3823;
assign w4287 = (w1602 & w4013) | (w1602 & w17447) | (w4013 & w17447);
assign w4288 = ~w4013 & w17448;
assign w4289 = pi330 & ~w4287;
assign w4290 = ~w4288 & w4289;
assign w4291 = ~w4285 & w4290;
assign w4292 = w4285 & ~w4290;
assign w4293 = ~w4291 & ~w4292;
assign w4294 = pi331 & w1339;
assign w4295 = (~w4018 & ~w4020) | (~w4018 & w17449) | (~w4020 & w17449);
assign w4296 = ~w4294 & w4295;
assign w4297 = w4294 & ~w4295;
assign w4298 = ~w4296 & ~w4297;
assign w4299 = ~w4293 & ~w4298;
assign w4300 = w4293 & w4298;
assign w4301 = ~w4299 & ~w4300;
assign w4302 = w4086 & w4301;
assign w4303 = ~w4086 & ~w4301;
assign w4304 = ~w4302 & ~w4303;
assign w4305 = w4081 & w4304;
assign w4306 = ~w4081 & ~w4304;
assign w4307 = ~w4305 & ~w4306;
assign w4308 = pi334 & ~w793;
assign w4309 = (~w3804 & ~w4029) | (~w3804 & w17450) | (~w4029 & w17450);
assign w4310 = ~w4308 & w4309;
assign w4311 = w4308 & ~w4309;
assign w4312 = ~w4310 & ~w4311;
assign w4313 = ~w4307 & ~w4312;
assign w4314 = w4307 & w4312;
assign w4315 = ~w4313 & ~w4314;
assign w4316 = ~w4076 & w4315;
assign w4317 = w4076 & ~w4315;
assign w4318 = ~w4316 & ~w4317;
assign w4319 = w4071 & ~w4318;
assign w4320 = ~w4071 & w4318;
assign w4321 = ~w4319 & ~w4320;
assign w4322 = ~w465 & w17451;
assign w4323 = (~w4322 & ~w4038) | (~w4322 & w17452) | (~w4038 & w17452);
assign w4324 = w4038 & w17453;
assign w4325 = ~w4323 & ~w4324;
assign w4326 = w4321 & w4325;
assign w4327 = ~w4321 & ~w4325;
assign w4328 = ~w4326 & ~w4327;
assign w4329 = w4066 & ~w4328;
assign w4330 = ~w4066 & w4328;
assign w4331 = ~w4329 & ~w4330;
assign w4332 = w4065 & w4331;
assign w4333 = ~w4065 & ~w4331;
assign w4334 = ~w4332 & ~w4333;
assign w4335 = (~w3791 & w4048) | (~w3791 & w17454) | (w4048 & w17454);
assign w4336 = ~w4051 & ~w4335;
assign w4337 = w4334 & ~w4336;
assign w4338 = ~w4334 & w4336;
assign w4339 = ~w4337 & ~w4338;
assign w4340 = pi128 & pi305;
assign w4341 = pi306 & w464;
assign w4342 = pi307 & ~w653;
assign w4343 = pi308 & w709;
assign w4344 = pi309 & w698;
assign w4345 = (~w3775 & ~w3776) | (~w3775 & w17455) | (~w3776 & w17455);
assign w4346 = pi310 & w855;
assign w4347 = (~w3678 & ~w3679) | (~w3678 & w17456) | (~w3679 & w17456);
assign w4348 = pi311 & w1159;
assign w4349 = pi312 & w1220;
assign w4350 = w1692 & w17457;
assign w4351 = pi315 & w1954;
assign w4352 = (~w3695 & ~w3696) | (~w3695 & w17458) | (~w3696 & w17458);
assign w4353 = ~w4351 & w4352;
assign w4354 = w4351 & ~w4352;
assign w4355 = ~w4353 & ~w4354;
assign w4356 = pi316 & ~w2473;
assign w4357 = pi317 & w2801;
assign w4358 = (~w3731 & ~w3733) | (~w3731 & w17459) | (~w3733 & w17459);
assign w4359 = w4357 & ~w4358;
assign w4360 = ~w4357 & w4358;
assign w4361 = ~w4359 & ~w4360;
assign w4362 = pi318 & w2925;
assign w4363 = (~w3699 & ~w3700) | (~w3699 & w17460) | (~w3700 & w17460);
assign w4364 = ~w3725 & ~w4363;
assign w4365 = pi319 & w3304;
assign w4366 = (~w3720 & ~w3721) | (~w3720 & w17461) | (~w3721 & w17461);
assign w4367 = pi320 & w3710;
assign w4368 = ~pi143 & pi144;
assign w4369 = pi143 & ~pi144;
assign w4370 = ~w4368 & ~w4369;
assign w4371 = (w3298 & w17463) | (w3298 & w17464) | (w17463 & w17464);
assign w4372 = ~pi141 & ~w4371;
assign w4373 = ~w3298 & w4369;
assign w4374 = (pi141 & ~w3704) | (pi141 & w17465) | (~w3704 & w17465);
assign w4375 = ~w4373 & w4374;
assign w4376 = ~w4372 & ~w4375;
assign w4377 = (~pi142 & w3298) | (~pi142 & w17466) | (w3298 & w17466);
assign w4378 = (~w4370 & ~w3298) | (~w4370 & w17467) | (~w3298 & w17467);
assign w4379 = ~w4377 & ~w4378;
assign w4380 = ~pi142 & ~w4370;
assign w4381 = ~w4379 & ~w4380;
assign w4382 = ~w4376 & ~w4381;
assign w4383 = pi321 & w4382;
assign w4384 = (~w3714 & ~w3715) | (~w3714 & w17468) | (~w3715 & w17468);
assign w4385 = ~w4383 & w4384;
assign w4386 = w4383 & ~w4384;
assign w4387 = ~w4385 & ~w4386;
assign w4388 = w4367 & w4387;
assign w4389 = ~w4367 & ~w4387;
assign w4390 = ~w4388 & ~w4389;
assign w4391 = w4366 & ~w4390;
assign w4392 = ~w4366 & w4390;
assign w4393 = ~w4391 & ~w4392;
assign w4394 = w4365 & w4393;
assign w4395 = ~w4365 & ~w4393;
assign w4396 = ~w4394 & ~w4395;
assign w4397 = ~w4364 & ~w4396;
assign w4398 = w4364 & w4396;
assign w4399 = ~w4397 & ~w4398;
assign w4400 = w4362 & ~w4399;
assign w4401 = ~w4362 & w4399;
assign w4402 = ~w4400 & ~w4401;
assign w4403 = ~w4361 & w4402;
assign w4404 = w4361 & ~w4402;
assign w4405 = ~w4403 & ~w4404;
assign w4406 = ~w4356 & ~w4405;
assign w4407 = w4356 & w4405;
assign w4408 = ~w4406 & ~w4407;
assign w4409 = (~w3697 & ~w3741) | (~w3697 & w17469) | (~w3741 & w17469);
assign w4410 = ~w3743 & ~w4409;
assign w4411 = w4408 & w4410;
assign w4412 = ~w4408 & ~w4410;
assign w4413 = ~w4411 & ~w4412;
assign w4414 = w4355 & w4413;
assign w4415 = ~w4355 & ~w4413;
assign w4416 = ~w4414 & ~w4415;
assign w4417 = w4350 & w4416;
assign w4418 = ~w4350 & ~w4416;
assign w4419 = ~w4417 & ~w4418;
assign w4420 = (~w3689 & ~w3691) | (~w3689 & w17470) | (~w3691 & w17470);
assign w4421 = w4419 & ~w4420;
assign w4422 = ~w4419 & w4420;
assign w4423 = ~w4421 & ~w4422;
assign w4424 = w1419 & w17471;
assign w4425 = (~w3756 & ~w3757) | (~w3756 & w17472) | (~w3757 & w17472);
assign w4426 = ~w4424 & w4425;
assign w4427 = w4424 & ~w4425;
assign w4428 = ~w4426 & ~w4427;
assign w4429 = w4423 & w4428;
assign w4430 = ~w4423 & ~w4428;
assign w4431 = ~w4429 & ~w4430;
assign w4432 = ~w4349 & ~w4431;
assign w4433 = w4349 & w4431;
assign w4434 = ~w4432 & ~w4433;
assign w4435 = (~w3684 & ~w3686) | (~w3684 & w17473) | (~w3686 & w17473);
assign w4436 = w4434 & w4435;
assign w4437 = ~w4434 & ~w4435;
assign w4438 = ~w4436 & ~w4437;
assign w4439 = (~w3766 & ~w3767) | (~w3766 & w17474) | (~w3767 & w17474);
assign w4440 = w4438 & w4439;
assign w4441 = ~w4438 & ~w4439;
assign w4442 = ~w4440 & ~w4441;
assign w4443 = w4348 & ~w4442;
assign w4444 = ~w4348 & w4442;
assign w4445 = ~w4443 & ~w4444;
assign w4446 = w4347 & ~w4445;
assign w4447 = ~w4347 & w4445;
assign w4448 = ~w4446 & ~w4447;
assign w4449 = ~w4346 & ~w4448;
assign w4450 = w4346 & w4448;
assign w4451 = ~w4449 & ~w4450;
assign w4452 = ~w4345 & w4451;
assign w4453 = w4345 & ~w4451;
assign w4454 = ~w4452 & ~w4453;
assign w4455 = w4344 & w4454;
assign w4456 = ~w4344 & ~w4454;
assign w4457 = ~w4455 & ~w4456;
assign w4458 = w4343 & w4457;
assign w4459 = ~w4343 & ~w4457;
assign w4460 = ~w4458 & ~w4459;
assign w4461 = (~w3671 & w3782) | (~w3671 & w17475) | (w3782 & w17475);
assign w4462 = w4460 & ~w4461;
assign w4463 = ~w4460 & w4461;
assign w4464 = ~w4462 & ~w4463;
assign w4465 = (~w3668 & w3785) | (~w3668 & w17476) | (w3785 & w17476);
assign w4466 = ~w4464 & ~w4465;
assign w4467 = w4464 & w4465;
assign w4468 = ~w4466 & ~w4467;
assign w4469 = w4342 & w4468;
assign w4470 = ~w4342 & ~w4468;
assign w4471 = ~w4469 & ~w4470;
assign w4472 = w4341 & w4471;
assign w4473 = ~w4341 & ~w4471;
assign w4474 = ~w4472 & ~w4473;
assign w4475 = w3789 & ~w4474;
assign w4476 = ~w3789 & w4474;
assign w4477 = ~w4475 & ~w4476;
assign w4478 = w4340 & w4477;
assign w4479 = ~w4340 & ~w4477;
assign w4480 = ~w4478 & ~w4479;
assign w4481 = ~w4339 & w4480;
assign w4482 = w4339 & ~w4480;
assign w4483 = ~w4481 & ~w4482;
assign w4484 = ~w135 & ~w4483;
assign w4485 = (pi161 & ~w135) | (pi161 & w17477) | (~w135 & w17477);
assign w4486 = ~w4484 & w4485;
assign w4487 = ~pi160 & ~w4061;
assign w4488 = ~w4486 & w4487;
assign w4489 = ~pi081 & ~pi161;
assign w4490 = pi128 & pi304;
assign w4491 = pi129 & ~pi305;
assign w4492 = (~w4491 & ~w4477) | (~w4491 & w17478) | (~w4477 & w17478);
assign w4493 = pi306 & ~w653;
assign w4494 = (~w3789 & ~w4471) | (~w3789 & w17479) | (~w4471 & w17479);
assign w4495 = ~w4473 & ~w4494;
assign w4496 = ~w4493 & ~w4495;
assign w4497 = w4493 & w4495;
assign w4498 = ~w4496 & ~w4497;
assign w4499 = pi307 & w709;
assign w4500 = (~w4466 & ~w4468) | (~w4466 & w17480) | (~w4468 & w17480);
assign w4501 = pi308 & w698;
assign w4502 = (~w4459 & ~w4460) | (~w4459 & w17481) | (~w4460 & w17481);
assign w4503 = w4501 & w4502;
assign w4504 = ~w4501 & ~w4502;
assign w4505 = ~w4503 & ~w4504;
assign w4506 = pi309 & w855;
assign w4507 = pi311 & w1220;
assign w4508 = (~w4432 & ~w4434) | (~w4432 & w17482) | (~w4434 & w17482);
assign w4509 = w1419 & w17483;
assign w4510 = w1692 & w17484;
assign w4511 = pi314 & w1954;
assign w4512 = pi315 & ~w2473;
assign w4513 = pi316 & w2801;
assign w4514 = pi317 & w2925;
assign w4515 = pi318 & w3304;
assign w4516 = (~w4362 & ~w4364) | (~w4362 & w17485) | (~w4364 & w17485);
assign w4517 = ~w4397 & ~w4516;
assign w4518 = pi319 & w3710;
assign w4519 = pi320 & w4382;
assign w4520 = ~pi145 & w4370;
assign w4521 = pi142 & pi144;
assign w4522 = pi145 & w4521;
assign w4523 = pi143 & pi145;
assign w4524 = (~w4523 & w3298) | (~w4523 & w17486) | (w3298 & w17486);
assign w4525 = pi142 & ~w4524;
assign w4526 = ~pi144 & ~pi145;
assign w4527 = pi145 & w4368;
assign w4528 = (~w4527 & ~w3298) | (~w4527 & w17487) | (~w3298 & w17487);
assign w4529 = ~pi142 & ~w4528;
assign w4530 = ~w4525 & ~w4529;
assign w4531 = ~w4522 & ~w4530;
assign w4532 = ~pi142 & w4526;
assign w4533 = (~w4532 & ~w3298) | (~w4532 & w17488) | (~w3298 & w17488);
assign w4534 = (pi145 & w3298) | (pi145 & w17489) | (w3298 & w17489);
assign w4535 = (pi141 & w4521) | (pi141 & w17490) | (w4521 & w17490);
assign w4536 = ~w4534 & w4535;
assign w4537 = (~w4520 & w4533) | (~w4520 & w17491) | (w4533 & w17491);
assign w4538 = ~w4536 & w4537;
assign w4539 = ~w4531 & w4538;
assign w4540 = ~w4531 & w17492;
assign w4541 = (~w4386 & ~w4387) | (~w4386 & w17493) | (~w4387 & w17493);
assign w4542 = ~w4540 & w4541;
assign w4543 = w4540 & ~w4541;
assign w4544 = ~w4542 & ~w4543;
assign w4545 = w4519 & w4544;
assign w4546 = ~w4519 & ~w4544;
assign w4547 = ~w4545 & ~w4546;
assign w4548 = (~w4392 & ~w4393) | (~w4392 & w17494) | (~w4393 & w17494);
assign w4549 = ~w4547 & w4548;
assign w4550 = w4547 & ~w4548;
assign w4551 = ~w4549 & ~w4550;
assign w4552 = w4518 & w4551;
assign w4553 = ~w4518 & ~w4551;
assign w4554 = ~w4552 & ~w4553;
assign w4555 = ~w4517 & ~w4554;
assign w4556 = w4517 & w4554;
assign w4557 = ~w4555 & ~w4556;
assign w4558 = w4515 & ~w4557;
assign w4559 = ~w4515 & w4557;
assign w4560 = ~w4558 & ~w4559;
assign w4561 = w4514 & ~w4560;
assign w4562 = ~w4514 & w4560;
assign w4563 = ~w4561 & ~w4562;
assign w4564 = (~w4359 & ~w4361) | (~w4359 & w17495) | (~w4361 & w17495);
assign w4565 = ~w4563 & w4564;
assign w4566 = w4563 & ~w4564;
assign w4567 = ~w4565 & ~w4566;
assign w4568 = ~w4411 & w17496;
assign w4569 = (w4567 & w4411) | (w4567 & w17497) | (w4411 & w17497);
assign w4570 = ~w4568 & ~w4569;
assign w4571 = w4513 & ~w4570;
assign w4572 = ~w4513 & w4570;
assign w4573 = ~w4571 & ~w4572;
assign w4574 = w4512 & ~w4573;
assign w4575 = ~w4512 & w4573;
assign w4576 = ~w4574 & ~w4575;
assign w4577 = (~w4354 & ~w4355) | (~w4354 & w17498) | (~w4355 & w17498);
assign w4578 = w4576 & ~w4577;
assign w4579 = ~w4576 & w4577;
assign w4580 = ~w4578 & ~w4579;
assign w4581 = w4511 & w4580;
assign w4582 = ~w4511 & ~w4580;
assign w4583 = ~w4581 & ~w4582;
assign w4584 = (~w4417 & ~w4419) | (~w4417 & w17499) | (~w4419 & w17499);
assign w4585 = w4583 & w4584;
assign w4586 = ~w4583 & ~w4584;
assign w4587 = ~w4585 & ~w4586;
assign w4588 = ~w4510 & w4587;
assign w4589 = w4510 & ~w4587;
assign w4590 = ~w4588 & ~w4589;
assign w4591 = (~w4427 & ~w4428) | (~w4427 & w17500) | (~w4428 & w17500);
assign w4592 = ~w4590 & w4591;
assign w4593 = w4590 & ~w4591;
assign w4594 = ~w4592 & ~w4593;
assign w4595 = w4509 & w4594;
assign w4596 = ~w4509 & ~w4594;
assign w4597 = ~w4595 & ~w4596;
assign w4598 = w4508 & w4597;
assign w4599 = ~w4508 & ~w4597;
assign w4600 = ~w4598 & ~w4599;
assign w4601 = w4507 & w4600;
assign w4602 = ~w4507 & ~w4600;
assign w4603 = ~w4601 & ~w4602;
assign w4604 = (~w4440 & ~w4442) | (~w4440 & w17501) | (~w4442 & w17501);
assign w4605 = w4603 & w4604;
assign w4606 = ~w4603 & ~w4604;
assign w4607 = ~w4605 & ~w4606;
assign w4608 = ~w1159 & w4346;
assign w4609 = (w4608 & w4347) | (w4608 & w17502) | (w4347 & w17502);
assign w4610 = ~w4607 & w4609;
assign w4611 = pi310 & w1159;
assign w4612 = ~w4607 & ~w4611;
assign w4613 = w4607 & w4611;
assign w4614 = ~w4612 & ~w4613;
assign w4615 = w4347 & ~w4614;
assign w4616 = w1213 & ~w4347;
assign w4617 = w4607 & w4616;
assign w4618 = (~w4445 & w4615) | (~w4445 & w17503) | (w4615 & w17503);
assign w4619 = w1159 & w4607;
assign w4620 = w855 & w4347;
assign w4621 = w4619 & ~w4620;
assign w4622 = w4347 & ~w4619;
assign w4623 = (w4445 & w4607) | (w4445 & w17504) | (w4607 & w17504);
assign w4624 = ~w4621 & w4623;
assign w4625 = ~w4622 & w4624;
assign w4626 = (~w4346 & ~w4347) | (~w4346 & w17505) | (~w4347 & w17505);
assign w4627 = w4614 & w4626;
assign w4628 = ~w4625 & ~w4627;
assign w4629 = ~w4610 & ~w4618;
assign w4630 = w4628 & w4629;
assign w4631 = w4506 & ~w4630;
assign w4632 = ~w4506 & w4630;
assign w4633 = ~w4631 & ~w4632;
assign w4634 = (~w4452 & ~w4454) | (~w4452 & w17506) | (~w4454 & w17506);
assign w4635 = ~w4633 & w4634;
assign w4636 = w4633 & ~w4634;
assign w4637 = ~w4635 & ~w4636;
assign w4638 = w4505 & w4637;
assign w4639 = ~w4505 & ~w4637;
assign w4640 = ~w4638 & ~w4639;
assign w4641 = w4500 & ~w4640;
assign w4642 = ~w4500 & w4640;
assign w4643 = ~w4641 & ~w4642;
assign w4644 = w4499 & ~w4643;
assign w4645 = ~w4499 & w4643;
assign w4646 = ~w4644 & ~w4645;
assign w4647 = w4498 & ~w4646;
assign w4648 = ~w4498 & w4646;
assign w4649 = ~w4647 & ~w4648;
assign w4650 = pi129 & ~w4649;
assign w4651 = ~pi129 & w4649;
assign w4652 = ~w4650 & ~w4651;
assign w4653 = w4492 & w4652;
assign w4654 = ~w4492 & ~w4652;
assign w4655 = ~w4653 & ~w4654;
assign w4656 = w4490 & w4655;
assign w4657 = ~w4490 & ~w4655;
assign w4658 = ~w4656 & ~w4657;
assign w4659 = pi339 & w456;
assign w4660 = pi336 & ~w615;
assign w4661 = ~w4070 & ~w4319;
assign w4662 = pi335 & ~w793;
assign w4663 = ~w4074 & ~w4315;
assign w4664 = ~w4663 & w17507;
assign w4665 = (~w4662 & w4663) | (~w4662 & w17508) | (w4663 & w17508);
assign w4666 = ~w4664 & ~w4665;
assign w4667 = (w955 & ~w4309) | (w955 & w17509) | (~w4309 & w17509);
assign w4668 = pi334 & ~w955;
assign w4669 = (w4309 & w17511) | (w4309 & w17512) | (w17511 & w17512);
assign w4670 = ~w4667 & ~w4669;
assign w4671 = w4077 & ~w4304;
assign w4672 = ~w4077 & w4304;
assign w4673 = ~w4671 & ~w4672;
assign w4674 = ~w4670 & w4673;
assign w4675 = (~w4668 & w4309) | (~w4668 & w17513) | (w4309 & w17513);
assign w4676 = (~w955 & ~w4309) | (~w955 & w17514) | (~w4309 & w17514);
assign w4677 = ~w4675 & ~w4676;
assign w4678 = (w4309 & w17515) | (w4309 & w17516) | (w17515 & w17516);
assign w4679 = (~w4677 & w4673) | (~w4677 & w17517) | (w4673 & w17517);
assign w4680 = ~w4674 & w4679;
assign w4681 = pi333 & w1101;
assign w4682 = pi332 & w1339;
assign w4683 = (~w4084 & ~w4301) | (~w4084 & w17518) | (~w4301 & w17518);
assign w4684 = ~w4682 & w4683;
assign w4685 = w4682 & ~w4683;
assign w4686 = ~w4684 & ~w4685;
assign w4687 = pi331 & w1602;
assign w4688 = (~w4297 & ~w4293) | (~w4297 & w17519) | (~w4293 & w17519);
assign w4689 = w4687 & ~w4688;
assign w4690 = ~w4687 & w4688;
assign w4691 = ~w4689 & ~w4690;
assign w4692 = pi328 & ~w2373;
assign w4693 = (w4279 & w17521) | (w4279 & w17522) | (w17521 & w17522);
assign w4694 = ~w4692 & w17669;
assign w4695 = ~w4693 & ~w4694;
assign w4696 = pi327 & w2698;
assign w4697 = (w4276 & w17524) | (w4276 & w17525) | (w17524 & w17525);
assign w4698 = ~w4696 & w17670;
assign w4699 = ~w4697 & ~w4698;
assign w4700 = (~w4264 & ~w4266) | (~w4264 & w17526) | (~w4266 & w17526);
assign w4701 = (~w4251 & ~w4252) | (~w4251 & w17527) | (~w4252 & w17527);
assign w4702 = (~w4242 & ~w3975) | (~w4242 & w17528) | (~w3975 & w17528);
assign w4703 = ~w4241 & w4702;
assign w4704 = w4241 & ~w4702;
assign w4705 = ~w4703 & ~w4704;
assign w4706 = w3975 & ~w4705;
assign w4707 = ~w3975 & w4705;
assign w4708 = ~w4706 & ~w4707;
assign w4709 = pi323 & ~w4708;
assign w4710 = pi144 & pi259;
assign w4711 = (~w4710 & w4241) | (~w4710 & w16585) | (w4241 & w16585);
assign w4712 = ~w4241 & w16586;
assign w4713 = ~w4711 & ~w4712;
assign w4714 = (~w4234 & ~w4221) | (~w4234 & w16587) | (~w4221 & w16587);
assign w4715 = ~w4226 & w4714;
assign w4716 = ~w4225 & w4715;
assign w4717 = ~w4222 & ~w4224;
assign w4718 = ~w4233 & ~w4717;
assign w4719 = ~w4716 & w4718;
assign w4720 = ~w4233 & ~w4714;
assign w4721 = w4717 & ~w4720;
assign w4722 = ~w4719 & ~w4721;
assign w4723 = pi143 & pi260;
assign w4724 = pi140 & pi263;
assign w4725 = ~w3939 & ~w4195;
assign w4726 = (~w4194 & ~w4725) | (~w4194 & w15867) | (~w4725 & w15867);
assign w4727 = w4183 & w4190;
assign w4728 = ~w4191 & ~w4727;
assign w4729 = pi137 & pi266;
assign w4730 = ~w4181 & ~w4184;
assign w4731 = ~w4180 & ~w4730;
assign w4732 = pi136 & pi267;
assign w4733 = pi135 & pi268;
assign w4734 = (~w4174 & w4176) | (~w4174 & w16588) | (w4176 & w16588);
assign w4735 = pi134 & pi269;
assign w4736 = pi133 & pi270;
assign w4737 = pi131 & pi272;
assign w4738 = pi130 & pi273;
assign w4739 = pi129 & pi274;
assign w4740 = pi128 & pi275;
assign w4741 = ~w4739 & ~w4740;
assign w4742 = w4739 & w4740;
assign w4743 = ~w4741 & ~w4742;
assign w4744 = ~w4743 & w17671;
assign w4745 = (w4122 & w17531) | (w4122 & w17532) | (w17531 & w17532);
assign w4746 = ~w4744 & ~w4745;
assign w4747 = ~w4738 & w4746;
assign w4748 = w4738 & ~w4746;
assign w4749 = ~w4747 & ~w4748;
assign w4750 = (w4140 & w17534) | (w4140 & w17535) | (w17534 & w17535);
assign w4751 = ~w4749 & w17672;
assign w4752 = ~w4750 & ~w4751;
assign w4753 = ~w4737 & ~w4752;
assign w4754 = w4737 & w4752;
assign w4755 = ~w4753 & ~w4754;
assign w4756 = w4755 & w17673;
assign w4757 = (w4146 & w17537) | (w4146 & w17538) | (w17537 & w17538);
assign w4758 = ~w4756 & ~w4757;
assign w4759 = (w4154 & w17539) | (w4154 & w17540) | (w17539 & w17540);
assign w4760 = (w15870 & ~w4154) | (w15870 & w17541) | (~w4154 & w17541);
assign w4761 = ~w4759 & ~w4760;
assign w4762 = pi132 & pi271;
assign w4763 = ~w4761 & w4762;
assign w4764 = w4761 & ~w4762;
assign w4765 = ~w4763 & ~w4764;
assign w4766 = ~w4736 & w4765;
assign w4767 = w4736 & ~w4765;
assign w4768 = ~w4766 & ~w4767;
assign w4769 = (~w4159 & w4162) | (~w4159 & w15871) | (w4162 & w15871);
assign w4770 = w4768 & w4769;
assign w4771 = ~w4768 & ~w4769;
assign w4772 = ~w4770 & ~w4771;
assign w4773 = ~w4735 & w4772;
assign w4774 = w4735 & ~w4772;
assign w4775 = ~w4773 & ~w4774;
assign w4776 = ~w4166 & ~w4170;
assign w4777 = w4775 & w4776;
assign w4778 = ~w4775 & ~w4776;
assign w4779 = ~w4777 & ~w4778;
assign w4780 = (w15868 & w16130) | (w15868 & w16131) | (w16130 & w16131);
assign w4781 = ~w4779 & w17674;
assign w4782 = ~w4780 & ~w4781;
assign w4783 = w4733 & w4782;
assign w4784 = ~w4733 & ~w4782;
assign w4785 = ~w4783 & ~w4784;
assign w4786 = ~w4732 & ~w4785;
assign w4787 = w4732 & w4785;
assign w4788 = ~w4786 & ~w4787;
assign w4789 = w4731 & ~w4788;
assign w4790 = ~w4731 & w4788;
assign w4791 = ~w4789 & ~w4790;
assign w4792 = w4729 & ~w4791;
assign w4793 = ~w4729 & w4791;
assign w4794 = ~w4792 & ~w4793;
assign w4795 = w4728 & ~w4794;
assign w4796 = ~w4728 & w4794;
assign w4797 = ~w4795 & ~w4796;
assign w4798 = w4726 & ~w4797;
assign w4799 = ~w4726 & w4797;
assign w4800 = ~w4798 & ~w4799;
assign w4801 = pi139 & pi264;
assign w4802 = pi138 & pi265;
assign w4803 = w4801 & ~w4802;
assign w4804 = ~w4801 & w4802;
assign w4805 = ~w4803 & ~w4804;
assign w4806 = w4800 & w4805;
assign w4807 = ~w4800 & ~w4805;
assign w4808 = ~w4806 & ~w4807;
assign w4809 = (~w4201 & w4205) | (~w4201 & w16392) | (w4205 & w16392);
assign w4810 = w4808 & w4809;
assign w4811 = ~w4808 & ~w4809;
assign w4812 = ~w4810 & ~w4811;
assign w4813 = w4724 & w4812;
assign w4814 = ~w4724 & ~w4812;
assign w4815 = ~w4813 & ~w4814;
assign w4816 = w4203 & ~w4211;
assign w4817 = ~w4212 & ~w4816;
assign w4818 = w4815 & ~w4817;
assign w4819 = ~w4815 & w4817;
assign w4820 = ~w4818 & ~w4819;
assign w4821 = (w4218 & ~w4214) | (w4218 & w17542) | (~w4214 & w17542);
assign w4822 = ~w4215 & ~w4821;
assign w4823 = w4820 & w4822;
assign w4824 = ~w4820 & ~w4822;
assign w4825 = ~w4823 & ~w4824;
assign w4826 = pi142 & pi261;
assign w4827 = pi141 & pi262;
assign w4828 = w4826 & ~w4827;
assign w4829 = ~w4826 & w4827;
assign w4830 = ~w4828 & ~w4829;
assign w4831 = w4825 & w4830;
assign w4832 = ~w4825 & ~w4830;
assign w4833 = ~w4831 & ~w4832;
assign w4834 = w4723 & ~w4833;
assign w4835 = ~w4723 & w4833;
assign w4836 = ~w4834 & ~w4835;
assign w4837 = w4722 & w4836;
assign w4838 = ~w4722 & ~w4836;
assign w4839 = ~w4837 & ~w4838;
assign w4840 = w4713 & w4839;
assign w4841 = ~w4713 & ~w4839;
assign w4842 = ~w4840 & ~w4841;
assign w4843 = (~w3975 & ~w4241) | (~w3975 & w16132) | (~w4241 & w16132);
assign w4844 = ~w4703 & ~w4843;
assign w4845 = pi145 & pi258;
assign w4846 = ~w4241 & w4845;
assign w4847 = w4241 & ~w4845;
assign w4848 = ~w4846 & ~w4847;
assign w4849 = w4844 & ~w4848;
assign w4850 = ~w4844 & w4848;
assign w4851 = ~w4849 & ~w4850;
assign w4852 = w4842 & w4851;
assign w4853 = ~w4842 & ~w4851;
assign w4854 = ~w4852 & ~w4853;
assign w4855 = ~w4854 & w16133;
assign w4856 = (~w4709 & w4854) | (~w4709 & w16134) | (w4854 & w16134);
assign w4857 = ~w4855 & ~w4856;
assign w4858 = w4701 & ~w4857;
assign w4859 = ~w4701 & w4857;
assign w4860 = ~w4858 & ~w4859;
assign w4861 = (~w4259 & ~w4256) | (~w4259 & w17543) | (~w4256 & w17543);
assign w4862 = w4860 & ~w4861;
assign w4863 = ~w4860 & w4861;
assign w4864 = ~w4862 & ~w4863;
assign w4865 = pi324 & w3979;
assign w4866 = (pi325 & w3567) | (pi325 & w17544) | (w3567 & w17544);
assign w4867 = w3979 & w17545;
assign w4868 = (w4866 & ~w3979) | (w4866 & w17546) | (~w3979 & w17546);
assign w4869 = ~w4867 & ~w4868;
assign w4870 = w4864 & w4869;
assign w4871 = ~w4864 & ~w4869;
assign w4872 = ~w4870 & ~w4871;
assign w4873 = w4700 & w4872;
assign w4874 = ~w4700 & ~w4872;
assign w4875 = ~w4873 & ~w4874;
assign w4876 = pi326 & ~w3183;
assign w4877 = (~w4273 & w16135) | (~w4273 & w16136) | (w16135 & w16136);
assign w4878 = (w4273 & w16137) | (w4273 & w16138) | (w16137 & w16138);
assign w4879 = ~w4877 & ~w4878;
assign w4880 = w4875 & ~w4879;
assign w4881 = ~w4875 & w4879;
assign w4882 = ~w4880 & ~w4881;
assign w4883 = w4699 & ~w4882;
assign w4884 = ~w4699 & w4882;
assign w4885 = ~w4883 & ~w4884;
assign w4886 = ~w4695 & ~w4885;
assign w4887 = w4695 & w4885;
assign w4888 = ~w4886 & ~w4887;
assign w4889 = pi329 & ~w2170;
assign w4890 = (w4282 & w17547) | (w4282 & w17548) | (w17547 & w17548);
assign w4891 = ~w4889 & w17675;
assign w4892 = ~w4890 & ~w4891;
assign w4893 = w4888 & w4892;
assign w4894 = ~w4888 & ~w4892;
assign w4895 = ~w4893 & ~w4894;
assign w4896 = pi330 & ~w1865;
assign w4897 = ~w4288 & w4896;
assign w4898 = (w4897 & ~w4285) | (w4897 & w17549) | (~w4285 & w17549);
assign w4899 = ~w4287 & ~w4896;
assign w4900 = (w4899 & w4285) | (w4899 & w17550) | (w4285 & w17550);
assign w4901 = ~w4898 & ~w4900;
assign w4902 = w4895 & w4901;
assign w4903 = ~w4895 & ~w4901;
assign w4904 = ~w4902 & ~w4903;
assign w4905 = ~w4691 & ~w4904;
assign w4906 = w4691 & w4904;
assign w4907 = ~w4905 & ~w4906;
assign w4908 = w4686 & w4907;
assign w4909 = ~w4686 & ~w4907;
assign w4910 = ~w4908 & ~w4909;
assign w4911 = w4681 & w4910;
assign w4912 = ~w4681 & ~w4910;
assign w4913 = ~w4911 & ~w4912;
assign w4914 = (~w4079 & ~w4304) | (~w4079 & w17551) | (~w4304 & w17551);
assign w4915 = ~w4913 & w4914;
assign w4916 = w4913 & ~w4914;
assign w4917 = ~w4915 & ~w4916;
assign w4918 = w4680 & w4917;
assign w4919 = ~w4680 & ~w4917;
assign w4920 = ~w4918 & ~w4919;
assign w4921 = ~w4666 & w4920;
assign w4922 = w4666 & ~w4920;
assign w4923 = ~w4921 & ~w4922;
assign w4924 = ~w4661 & w4923;
assign w4925 = w4661 & ~w4923;
assign w4926 = ~w4924 & ~w4925;
assign w4927 = w4660 & w4926;
assign w4928 = ~w4660 & ~w4926;
assign w4929 = ~w4927 & ~w4928;
assign w4930 = (pi337 & ~w536) | (pi337 & w17552) | (~w536 & w17552);
assign w4931 = (~w4324 & ~w4321) | (~w4324 & w16140) | (~w4321 & w16140);
assign w4932 = ~w4930 & w4931;
assign w4933 = w4930 & ~w4931;
assign w4934 = ~w4932 & ~w4933;
assign w4935 = w4929 & w4934;
assign w4936 = ~w4929 & ~w4934;
assign w4937 = ~w4935 & ~w4936;
assign w4938 = (~w466 & ~w4328) | (~w466 & w16895) | (~w4328 & w16895);
assign w4939 = w971 & w4328;
assign w4940 = (pi338 & ~w4328) | (pi338 & w17553) | (~w4328 & w17553);
assign w4941 = ~w4938 & w4940;
assign w4942 = w4937 & ~w4941;
assign w4943 = ~w4937 & w4941;
assign w4944 = ~w4942 & ~w4943;
assign w4945 = w4659 & ~w4944;
assign w4946 = ~w4659 & w4944;
assign w4947 = ~w4945 & ~w4946;
assign w4948 = ~w4063 & ~w4332;
assign w4949 = ~w4947 & ~w4948;
assign w4950 = w4947 & w4948;
assign w4951 = ~w4949 & ~w4950;
assign w4952 = pi275 & w4951;
assign w4953 = ~pi275 & ~w4951;
assign w4954 = ~w4952 & ~w4953;
assign w4955 = (~w4338 & ~w4339) | (~w4338 & w17554) | (~w4339 & w17554);
assign w4956 = w4954 & w4955;
assign w4957 = ~w4954 & ~w4955;
assign w4958 = ~w4956 & ~w4957;
assign w4959 = (~w4658 & w4954) | (~w4658 & w17555) | (w4954 & w17555);
assign w4960 = ~w4956 & w4959;
assign w4961 = (~w135 & w4958) | (~w135 & w17556) | (w4958 & w17556);
assign w4962 = ~w4960 & w4961;
assign w4963 = (pi161 & ~w135) | (pi161 & w17557) | (~w135 & w17557);
assign w4964 = ~w4962 & w4963;
assign w4965 = ~pi160 & ~w4489;
assign w4966 = ~w4964 & w4965;
assign w4967 = ~pi082 & ~pi161;
assign w4968 = pi276 & w135;
assign w4969 = ~w4956 & ~w4959;
assign w4970 = pi340 & w456;
assign w4971 = ~w4944 & w17558;
assign w4972 = ~w465 & w17559;
assign w4973 = (~w4972 & w4944) | (~w4972 & w17560) | (w4944 & w17560);
assign w4974 = ~w4971 & ~w4973;
assign w4975 = (~w4939 & ~w4937) | (~w4939 & w16141) | (~w4937 & w16141);
assign w4976 = (w4937 & w17563) | (w4937 & w17564) | (w17563 & w17564);
assign w4977 = ~w537 & ~w4975;
assign w4978 = w4976 & ~w4977;
assign w4979 = pi337 & ~w615;
assign w4980 = (w4929 & w16142) | (w4929 & w16143) | (w16142 & w16143);
assign w4981 = (~w4929 & w16144) | (~w4929 & w16145) | (w16144 & w16145);
assign w4982 = ~w4980 & ~w4981;
assign w4983 = pi336 & ~w793;
assign w4984 = (w4926 & w16146) | (w4926 & w16147) | (w16146 & w16147);
assign w4985 = (~w4926 & w16148) | (~w4926 & w16149) | (w16148 & w16149);
assign w4986 = ~w4984 & ~w4985;
assign w4987 = pi335 & ~w955;
assign w4988 = pi334 & w1101;
assign w4989 = (~w4311 & ~w4307) | (~w4311 & w17565) | (~w4307 & w17565);
assign w4990 = w4668 & ~w4989;
assign w4991 = ~w4668 & w4989;
assign w4992 = (w4917 & w16150) | (w4917 & w16151) | (w16150 & w16151);
assign w4993 = ~w4988 & w17676;
assign w4994 = ~w4992 & ~w4993;
assign w4995 = pi333 & w1339;
assign w4996 = (~w4913 & w16152) | (~w4913 & w16153) | (w16152 & w16153);
assign w4997 = (w4913 & w16154) | (w4913 & w16155) | (w16154 & w16155);
assign w4998 = ~w4996 & ~w4997;
assign w4999 = pi332 & w1602;
assign w5000 = ~w4908 & w16156;
assign w5001 = (w4999 & w4908) | (w4999 & w16157) | (w4908 & w16157);
assign w5002 = ~w5000 & ~w5001;
assign w5003 = pi331 & ~w1865;
assign w5004 = (~w4689 & ~w4691) | (~w4689 & w16158) | (~w4691 & w16158);
assign w5005 = w5003 & ~w5004;
assign w5006 = ~w5003 & w5004;
assign w5007 = ~w5005 & ~w5006;
assign w5008 = ~w2170 & w17677;
assign w5009 = ~w4898 & w17678;
assign w5010 = pi330 & ~w5009;
assign w5011 = ~w5008 & w5010;
assign w5012 = pi329 & ~w2373;
assign w5013 = (w5012 & w4893) | (w5012 & w17567) | (w4893 & w17567);
assign w5014 = ~w4893 & w17568;
assign w5015 = ~w5013 & ~w5014;
assign w5016 = pi327 & ~w3183;
assign w5017 = w4866 & w4872;
assign w5018 = ~w4874 & ~w5017;
assign w5019 = pi325 & w3979;
assign w5020 = w5018 & ~w5019;
assign w5021 = ~w5018 & w5019;
assign w5022 = ~w5020 & ~w5021;
assign w5023 = (pi326 & w3567) | (pi326 & w17569) | (w3567 & w17569);
assign w5024 = (~w4865 & ~w4860) | (~w4865 & w17570) | (~w4860 & w17570);
assign w5025 = ~w4863 & ~w5024;
assign w5026 = w5023 & ~w5025;
assign w5027 = ~w5023 & w5025;
assign w5028 = ~w5026 & ~w5027;
assign w5029 = w5022 & w5028;
assign w5030 = ~w5022 & ~w5028;
assign w5031 = ~w5029 & ~w5030;
assign w5032 = ~w4877 & ~w4881;
assign w5033 = w4842 & ~w4845;
assign w5034 = ~w4842 & w4845;
assign w5035 = ~w5033 & ~w5034;
assign w5036 = (w4844 & w4842) | (w4844 & w17571) | (w4842 & w17571);
assign w5037 = ~w5036 & w17679;
assign w5038 = ~w5033 & ~w5037;
assign w5039 = w5033 & w17679;
assign w5040 = ~w5038 & ~w5039;
assign w5041 = pi146 & pi258;
assign w5042 = pi145 & pi259;
assign w5043 = pi144 & pi260;
assign w5044 = (~w4839 & w16393) | (~w4839 & w16394) | (w16393 & w16394);
assign w5045 = (w15875 & w4839) | (w15875 & w16395) | (w4839 & w16395);
assign w5046 = ~w5044 & ~w5045;
assign w5047 = pi143 & pi261;
assign w5048 = pi142 & pi262;
assign w5049 = pi141 & pi263;
assign w5050 = (~w4813 & w4817) | (~w4813 & w16396) | (w4817 & w16396);
assign w5051 = pi139 & pi265;
assign w5052 = pi138 & pi266;
assign w5053 = pi136 & pi268;
assign w5054 = pi135 & pi269;
assign w5055 = pi134 & pi270;
assign w5056 = pi133 & pi271;
assign w5057 = pi132 & pi272;
assign w5058 = pi131 & pi273;
assign w5059 = pi130 & pi274;
assign w5060 = pi129 & pi275;
assign w5061 = pi128 & pi276;
assign w5062 = ~w5060 & ~w5061;
assign w5063 = w5060 & w5061;
assign w5064 = ~w5062 & ~w5063;
assign w5065 = (w16160 & w3478) | (w16160 & w17572) | (w3478 & w17572);
assign w5066 = ~w3865 & ~w4127;
assign w5067 = ~w4742 & w5066;
assign w5068 = (~w4741 & w5065) | (~w4741 & w17573) | (w5065 & w17573);
assign w5069 = w5064 & ~w5068;
assign w5070 = (w5065 & w17574) | (w5065 & w17575) | (w17574 & w17575);
assign w5071 = (w5059 & w5069) | (w5059 & w17576) | (w5069 & w17576);
assign w5072 = ~w5069 & w17577;
assign w5073 = ~w5071 & ~w5072;
assign w5074 = (~w4748 & w16161) | (~w4748 & w17672) | (w16161 & w17672);
assign w5075 = ~w5073 & w5074;
assign w5076 = (w4140 & w17580) | (w4140 & w17581) | (w17580 & w17581);
assign w5077 = ~w5075 & ~w5076;
assign w5078 = ~w5058 & ~w5077;
assign w5079 = w5058 & w5077;
assign w5080 = ~w5078 & ~w5079;
assign w5081 = ~w4754 & ~w4756;
assign w5082 = ~w5080 & w5081;
assign w5083 = w5080 & ~w5081;
assign w5084 = ~w5082 & ~w5083;
assign w5085 = ~w5057 & ~w5084;
assign w5086 = w5057 & w5084;
assign w5087 = ~w5085 & ~w5086;
assign w5088 = ~w4760 & ~w4762;
assign w5089 = ~w4759 & ~w5088;
assign w5090 = ~w5087 & w5089;
assign w5091 = w5087 & ~w5089;
assign w5092 = ~w5090 & ~w5091;
assign w5093 = ~w4766 & ~w4769;
assign w5094 = ~w5093 & w16162;
assign w5095 = (~w5092 & w5093) | (~w5092 & w16163) | (w5093 & w16163);
assign w5096 = ~w5094 & ~w5095;
assign w5097 = w5056 & ~w5096;
assign w5098 = ~w5056 & w5096;
assign w5099 = ~w5097 & ~w5098;
assign w5100 = (~w4774 & w4776) | (~w4774 & w15876) | (w4776 & w15876);
assign w5101 = ~w5099 & ~w5100;
assign w5102 = w5099 & w5100;
assign w5103 = ~w5101 & ~w5102;
assign w5104 = w5055 & w5103;
assign w5105 = ~w5055 & ~w5103;
assign w5106 = ~w5104 & ~w5105;
assign w5107 = ~w5054 & ~w5106;
assign w5108 = w5054 & w5106;
assign w5109 = ~w5107 & ~w5108;
assign w5110 = (~w4781 & ~w4782) | (~w4781 & w15877) | (~w4782 & w15877);
assign w5111 = ~w5109 & w5110;
assign w5112 = w5109 & ~w5110;
assign w5113 = ~w5111 & ~w5112;
assign w5114 = w5053 & w5113;
assign w5115 = ~w5053 & ~w5113;
assign w5116 = ~w5114 & ~w5115;
assign w5117 = pi137 & pi267;
assign w5118 = ~w4731 & ~w4787;
assign w5119 = (~w4786 & w4731) | (~w4786 & w16164) | (w4731 & w16164);
assign w5120 = (w5117 & w5118) | (w5117 & w15878) | (w5118 & w15878);
assign w5121 = ~w5118 & w15879;
assign w5122 = ~w5120 & ~w5121;
assign w5123 = w5116 & w5122;
assign w5124 = ~w5116 & ~w5122;
assign w5125 = ~w5123 & ~w5124;
assign w5126 = (~w4793 & ~w4728) | (~w4793 & w17583) | (~w4728 & w17583);
assign w5127 = w5125 & w5126;
assign w5128 = ~w5125 & ~w5126;
assign w5129 = ~w5127 & ~w5128;
assign w5130 = w5052 & ~w5129;
assign w5131 = ~w5052 & w5129;
assign w5132 = ~w5130 & ~w5131;
assign w5133 = (~w4802 & w4726) | (~w4802 & w17584) | (w4726 & w17584);
assign w5134 = ~w4798 & ~w5133;
assign w5135 = w5132 & w5134;
assign w5136 = ~w5132 & ~w5134;
assign w5137 = ~w5135 & ~w5136;
assign w5138 = ~w5051 & ~w5137;
assign w5139 = w5051 & w5137;
assign w5140 = ~w5138 & ~w5139;
assign w5141 = pi140 & pi264;
assign w5142 = w4801 & w4808;
assign w5143 = ~w4811 & ~w5142;
assign w5144 = w5141 & ~w5143;
assign w5145 = ~w5141 & w5143;
assign w5146 = ~w5144 & ~w5145;
assign w5147 = w5140 & w5146;
assign w5148 = ~w5140 & ~w5146;
assign w5149 = ~w5147 & ~w5148;
assign w5150 = ~w5050 & w5149;
assign w5151 = w5050 & ~w5149;
assign w5152 = ~w5150 & ~w5151;
assign w5153 = w5049 & w5152;
assign w5154 = ~w5049 & ~w5152;
assign w5155 = ~w5153 & ~w5154;
assign w5156 = (~w4827 & ~w4822) | (~w4827 & w15880) | (~w4822 & w15880);
assign w5157 = ~w4824 & ~w5156;
assign w5158 = w5155 & ~w5157;
assign w5159 = ~w5155 & w5157;
assign w5160 = ~w5158 & ~w5159;
assign w5161 = ~w5048 & w5160;
assign w5162 = w5048 & ~w5160;
assign w5163 = ~w5161 & ~w5162;
assign w5164 = ~w4717 & ~w4833;
assign w5165 = ~w4826 & w4833;
assign w5166 = ~w5164 & ~w5165;
assign w5167 = w5163 & w5166;
assign w5168 = ~w5163 & ~w5166;
assign w5169 = ~w5167 & ~w5168;
assign w5170 = w5047 & w5169;
assign w5171 = ~w5047 & ~w5169;
assign w5172 = ~w5170 & ~w5171;
assign w5173 = ~w4233 & ~w4716;
assign w5174 = ~w4723 & ~w5173;
assign w5175 = w4723 & w5173;
assign w5176 = w4717 & w4833;
assign w5177 = ~w5164 & ~w5176;
assign w5178 = ~w5175 & w5177;
assign w5179 = ~w5174 & ~w5178;
assign w5180 = ~w5172 & w5179;
assign w5181 = w5172 & ~w5179;
assign w5182 = ~w5180 & ~w5181;
assign w5183 = w5046 & w5182;
assign w5184 = ~w5046 & ~w5182;
assign w5185 = ~w5183 & ~w5184;
assign w5186 = ~w5042 & w5185;
assign w5187 = w5042 & ~w5185;
assign w5188 = ~w5186 & ~w5187;
assign w5189 = w5041 & w5188;
assign w5190 = ~w5041 & ~w5188;
assign w5191 = ~w5189 & ~w5190;
assign w5192 = w5040 & w5191;
assign w5193 = ~w5040 & ~w5191;
assign w5194 = ~w5192 & ~w5193;
assign w5195 = ~w4855 & ~w4859;
assign w5196 = w5194 & w15881;
assign w5197 = (w5195 & ~w5194) | (w5195 & w15882) | (~w5194 & w15882);
assign w5198 = ~w5196 & ~w5197;
assign w5199 = pi323 & ~w4854;
assign w5200 = pi324 & ~w4708;
assign w5201 = ~w5199 & w5200;
assign w5202 = w5199 & ~w5200;
assign w5203 = ~w5201 & ~w5202;
assign w5204 = w5198 & w5203;
assign w5205 = ~w5198 & ~w5203;
assign w5206 = ~w5204 & ~w5205;
assign w5207 = w5032 & ~w5206;
assign w5208 = ~w5032 & w5206;
assign w5209 = ~w5207 & ~w5208;
assign w5210 = w5031 & w5209;
assign w5211 = ~w5031 & ~w5209;
assign w5212 = ~w5210 & ~w5211;
assign w5213 = w5016 & ~w5212;
assign w5214 = ~w5016 & w5212;
assign w5215 = ~w5213 & ~w5214;
assign w5216 = ~w4697 & ~w4883;
assign w5217 = w5215 & ~w5216;
assign w5218 = ~w5215 & w5216;
assign w5219 = ~w5217 & ~w5218;
assign w5220 = pi328 & w2698;
assign w5221 = ~w4693 & ~w4887;
assign w5222 = w5220 & ~w5221;
assign w5223 = ~w5220 & w5221;
assign w5224 = ~w5222 & ~w5223;
assign w5225 = w5219 & w5224;
assign w5226 = ~w5219 & ~w5224;
assign w5227 = ~w5225 & ~w5226;
assign w5228 = ~w5015 & ~w5227;
assign w5229 = w5015 & w5227;
assign w5230 = ~w5228 & ~w5229;
assign w5231 = w5011 & w5230;
assign w5232 = ~w5011 & ~w5230;
assign w5233 = ~w5231 & ~w5232;
assign w5234 = w5007 & w5233;
assign w5235 = ~w5007 & ~w5233;
assign w5236 = ~w5234 & ~w5235;
assign w5237 = ~w5002 & w5236;
assign w5238 = w5002 & ~w5236;
assign w5239 = ~w5237 & ~w5238;
assign w5240 = w4998 & ~w5239;
assign w5241 = ~w4998 & w5239;
assign w5242 = ~w5240 & ~w5241;
assign w5243 = ~w4994 & w5242;
assign w5244 = w4994 & ~w5242;
assign w5245 = ~w5243 & ~w5244;
assign w5246 = ~w4664 & ~w4922;
assign w5247 = w5245 & w5246;
assign w5248 = ~w5245 & ~w5246;
assign w5249 = ~w5247 & ~w5248;
assign w5250 = w4987 & w5249;
assign w5251 = ~w4987 & ~w5249;
assign w5252 = ~w5250 & ~w5251;
assign w5253 = w4986 & w5252;
assign w5254 = ~w4986 & ~w5252;
assign w5255 = ~w5253 & ~w5254;
assign w5256 = w4982 & w5255;
assign w5257 = ~w4982 & ~w5255;
assign w5258 = ~w5256 & ~w5257;
assign w5259 = ~w4978 & w5258;
assign w5260 = w4978 & ~w5258;
assign w5261 = ~w5259 & ~w5260;
assign w5262 = w4974 & ~w5261;
assign w5263 = ~w4974 & w5261;
assign w5264 = ~w5262 & ~w5263;
assign w5265 = w4970 & w5264;
assign w5266 = ~w4970 & ~w5264;
assign w5267 = ~w5265 & ~w5266;
assign w5268 = ~w4949 & ~w4952;
assign w5269 = ~w5267 & ~w5268;
assign w5270 = w5267 & w5268;
assign w5271 = ~w5269 & ~w5270;
assign w5272 = pi276 & w5271;
assign w5273 = ~pi276 & ~w5271;
assign w5274 = ~w5272 & ~w5273;
assign w5275 = pi128 & pi303;
assign w5276 = pi304 & w464;
assign w5277 = ~w4656 & ~w5276;
assign w5278 = ~pi129 & w4656;
assign w5279 = ~w5277 & ~w5278;
assign w5280 = pi306 & w709;
assign w5281 = pi307 & w698;
assign w5282 = pi308 & w855;
assign w5283 = pi309 & w1159;
assign w5284 = pi310 & w1220;
assign w5285 = pi311 & w1420;
assign w5286 = pi312 & w1693;
assign w5287 = pi313 & w1954;
assign w5288 = (w5287 & w4593) | (w5287 & w16165) | (w4593 & w16165);
assign w5289 = ~w4593 & w16166;
assign w5290 = ~w5288 & ~w5289;
assign w5291 = pi314 & ~w2473;
assign w5292 = pi315 & w2801;
assign w5293 = (~w4574 & w4577) | (~w4574 & w16167) | (w4577 & w16167);
assign w5294 = ~w5292 & w5293;
assign w5295 = w5292 & ~w5293;
assign w5296 = ~w5294 & ~w5295;
assign w5297 = pi316 & w2925;
assign w5298 = pi317 & w3304;
assign w5299 = pi318 & w3710;
assign w5300 = pi319 & w4382;
assign w5301 = (~w4518 & w4548) | (~w4518 & w15883) | (w4548 & w15883);
assign w5302 = ~w4549 & ~w5301;
assign w5303 = pi320 & w4539;
assign w5304 = ~pi143 & ~pi145;
assign w5305 = pi144 & ~w5304;
assign w5306 = ~w3298 & w4523;
assign w5307 = ~w4521 & ~w5306;
assign w5308 = pi141 & ~w5307;
assign w5309 = ~w4525 & ~w5305;
assign w5310 = ~w5308 & w5309;
assign w5311 = ~pi146 & w5310;
assign w5312 = pi146 & ~w5310;
assign w5313 = ~w5311 & ~w5312;
assign w5314 = pi145 & w5313;
assign w5315 = ~pi145 & ~w5313;
assign w5316 = ~w5314 & ~w5315;
assign w5317 = pi321 & w5316;
assign w5318 = (~w4543 & ~w4544) | (~w4543 & w16168) | (~w4544 & w16168);
assign w5319 = ~w5317 & w5318;
assign w5320 = w5317 & ~w5318;
assign w5321 = ~w5319 & ~w5320;
assign w5322 = w5303 & w5321;
assign w5323 = ~w5303 & ~w5321;
assign w5324 = ~w5322 & ~w5323;
assign w5325 = w5302 & w5324;
assign w5326 = ~w5302 & ~w5324;
assign w5327 = ~w5325 & ~w5326;
assign w5328 = w5300 & ~w5327;
assign w5329 = ~w5300 & w5327;
assign w5330 = ~w5328 & ~w5329;
assign w5331 = w5299 & ~w5330;
assign w5332 = ~w5299 & w5330;
assign w5333 = ~w5331 & ~w5332;
assign w5334 = ~w4555 & ~w4559;
assign w5335 = w5333 & w5334;
assign w5336 = ~w5333 & ~w5334;
assign w5337 = ~w5335 & ~w5336;
assign w5338 = w5298 & w5337;
assign w5339 = ~w5298 & ~w5337;
assign w5340 = ~w5338 & ~w5339;
assign w5341 = ~w4561 & ~w4566;
assign w5342 = w5340 & w5341;
assign w5343 = ~w5340 & ~w5341;
assign w5344 = ~w5342 & ~w5343;
assign w5345 = w4568 & w5344;
assign w5346 = w4569 & ~w5344;
assign w5347 = ~w5345 & ~w5346;
assign w5348 = w5297 & ~w5347;
assign w5349 = ~w4568 & ~w5344;
assign w5350 = w2801 & w2925;
assign w5351 = ~w4569 & w5350;
assign w5352 = w5349 & w5351;
assign w5353 = w5297 & ~w5344;
assign w5354 = ~w5297 & w5344;
assign w5355 = ~w4513 & ~w4569;
assign w5356 = ~w5353 & w5355;
assign w5357 = ~w5354 & w5356;
assign w5358 = ~w2925 & ~w5345;
assign w5359 = ~w5349 & w5358;
assign w5360 = ~w4572 & w5359;
assign w5361 = ~w5348 & ~w5352;
assign w5362 = ~w5357 & w5361;
assign w5363 = ~w5360 & w5362;
assign w5364 = ~w5296 & w5363;
assign w5365 = w5296 & ~w5363;
assign w5366 = ~w5364 & ~w5365;
assign w5367 = w5291 & w5366;
assign w5368 = ~w5291 & ~w5366;
assign w5369 = ~w5367 & ~w5368;
assign w5370 = ~w4582 & ~w4585;
assign w5371 = ~w5369 & w5370;
assign w5372 = w5369 & ~w5370;
assign w5373 = ~w5371 & ~w5372;
assign w5374 = w5290 & ~w5373;
assign w5375 = ~w5290 & w5373;
assign w5376 = ~w5374 & ~w5375;
assign w5377 = ~w5286 & ~w5376;
assign w5378 = w5286 & w5376;
assign w5379 = ~w5377 & ~w5378;
assign w5380 = ~w4595 & ~w4598;
assign w5381 = w5379 & w5380;
assign w5382 = ~w5379 & ~w5380;
assign w5383 = ~w5381 & ~w5382;
assign w5384 = ~w4601 & ~w4605;
assign w5385 = ~w5383 & ~w5384;
assign w5386 = w5383 & w5384;
assign w5387 = ~w5385 & ~w5386;
assign w5388 = w5285 & w5387;
assign w5389 = ~w5285 & ~w5387;
assign w5390 = ~w5388 & ~w5389;
assign w5391 = w5284 & w5390;
assign w5392 = ~w5284 & ~w5390;
assign w5393 = ~w5391 & ~w5392;
assign w5394 = ~w4612 & w17680;
assign w5395 = ~w5393 & ~w5394;
assign w5396 = w5393 & w5394;
assign w5397 = ~w5395 & ~w5396;
assign w5398 = (~w4631 & ~w4633) | (~w4631 & w16169) | (~w4633 & w16169);
assign w5399 = ~w5397 & w5398;
assign w5400 = w5397 & ~w5398;
assign w5401 = ~w5399 & ~w5400;
assign w5402 = w5283 & w5401;
assign w5403 = ~w5283 & ~w5401;
assign w5404 = ~w5402 & ~w5403;
assign w5405 = w5282 & w5404;
assign w5406 = ~w5282 & ~w5404;
assign w5407 = ~w5405 & ~w5406;
assign w5408 = ~w4503 & ~w4638;
assign w5409 = w5407 & ~w5408;
assign w5410 = ~w5407 & w5408;
assign w5411 = ~w5409 & ~w5410;
assign w5412 = (~w4641 & ~w4643) | (~w4641 & w16170) | (~w4643 & w16170);
assign w5413 = w5411 & w5412;
assign w5414 = ~w5411 & ~w5412;
assign w5415 = ~w5413 & ~w5414;
assign w5416 = w5281 & ~w5415;
assign w5417 = ~w5281 & w5415;
assign w5418 = ~w5416 & ~w5417;
assign w5419 = w5280 & ~w5418;
assign w5420 = ~w5280 & w5418;
assign w5421 = ~w5419 & ~w5420;
assign w5422 = ~w4497 & ~w4647;
assign w5423 = w5421 & ~w5422;
assign w5424 = ~w5421 & w5422;
assign w5425 = ~w5423 & ~w5424;
assign w5426 = pi128 & w605;
assign w5427 = ~w4652 & w5426;
assign w5428 = w651 & ~w4649;
assign w5429 = w4340 & ~w4477;
assign w5430 = ~w4650 & w5429;
assign w5431 = pi128 & w4651;
assign w5432 = ~w5430 & ~w5431;
assign w5433 = pi130 & ~w4650;
assign w5434 = w5432 & w5433;
assign w5435 = ~w5427 & ~w5428;
assign w5436 = ~w5434 & w5435;
assign w5437 = pi305 & ~w5436;
assign w5438 = pi305 & w651;
assign w5439 = ~w652 & ~w5438;
assign w5440 = w5430 & w5439;
assign w5441 = ~w5437 & ~w5440;
assign w5442 = w5425 & ~w5441;
assign w5443 = ~w5425 & w5441;
assign w5444 = ~w5442 & ~w5443;
assign w5445 = w5279 & w5444;
assign w5446 = ~w5279 & ~w5444;
assign w5447 = ~w5445 & ~w5446;
assign w5448 = w5275 & w5447;
assign w5449 = ~w5275 & ~w5447;
assign w5450 = ~w5448 & ~w5449;
assign w5451 = w5274 & ~w5450;
assign w5452 = ~w5274 & w5450;
assign w5453 = ~w5451 & ~w5452;
assign w5454 = w4969 & ~w5453;
assign w5455 = ~w4969 & ~w5452;
assign w5456 = ~w5451 & w5455;
assign w5457 = ~w135 & ~w5454;
assign w5458 = ~w5456 & w5457;
assign w5459 = pi161 & ~w4968;
assign w5460 = ~w5458 & w5459;
assign w5461 = ~pi160 & ~w4967;
assign w5462 = ~w5460 & w5461;
assign w5463 = ~pi083 & ~pi161;
assign w5464 = pi277 & w135;
assign w5465 = pi341 & w456;
assign w5466 = pi340 & w466;
assign w5467 = ~w5265 & ~w5466;
assign w5468 = w466 & w5265;
assign w5469 = ~w5467 & ~w5468;
assign w5470 = ~w4977 & ~w5258;
assign w5471 = w4976 & ~w5470;
assign w5472 = ~w615 & w5471;
assign w5473 = pi338 & ~w615;
assign w5474 = ~w5471 & ~w5473;
assign w5475 = ~w5472 & ~w5474;
assign w5476 = pi337 & ~w793;
assign w5477 = ~w4980 & ~w5256;
assign w5478 = ~w5476 & w5477;
assign w5479 = w5476 & ~w5477;
assign w5480 = ~w5478 & ~w5479;
assign w5481 = pi335 & w1101;
assign w5482 = pi334 & w1339;
assign w5483 = ~w4993 & ~w5244;
assign w5484 = ~w5482 & ~w5483;
assign w5485 = w5482 & w5483;
assign w5486 = ~w5484 & ~w5485;
assign w5487 = pi333 & w1602;
assign w5488 = ~w4997 & ~w5240;
assign w5489 = w5487 & ~w5488;
assign w5490 = ~w5487 & w5488;
assign w5491 = ~w5489 & ~w5490;
assign w5492 = pi331 & ~w2170;
assign w5493 = ~w5005 & ~w5234;
assign w5494 = ~w5492 & w5493;
assign w5495 = w5492 & ~w5493;
assign w5496 = ~w5494 & ~w5495;
assign w5497 = ~w5008 & ~w5230;
assign w5498 = ~w2373 & ~w5009;
assign w5499 = ~w5497 & w5498;
assign w5500 = pi330 & ~w2373;
assign w5501 = w5010 & w5230;
assign w5502 = ~w5008 & ~w5500;
assign w5503 = ~w5501 & w5502;
assign w5504 = ~w5499 & ~w5503;
assign w5505 = (~w5213 & ~w5215) | (~w5213 & w17585) | (~w5215 & w17585);
assign w5506 = pi327 & ~w3568;
assign w5507 = ~w5505 & w5506;
assign w5508 = w5505 & ~w5506;
assign w5509 = ~w5507 & ~w5508;
assign w5510 = pi326 & w3979;
assign w5511 = ~w5023 & ~w5032;
assign w5512 = w5023 & w5032;
assign w5513 = w5025 & ~w5206;
assign w5514 = ~w5025 & w5206;
assign w5515 = ~w5513 & ~w5514;
assign w5516 = w5022 & ~w5515;
assign w5517 = ~w5022 & w5515;
assign w5518 = ~w5512 & ~w5516;
assign w5519 = ~w5517 & w5518;
assign w5520 = ~w5511 & ~w5519;
assign w5521 = ~w5510 & ~w5520;
assign w5522 = w5510 & w5520;
assign w5523 = ~w5521 & ~w5522;
assign w5524 = pi325 & ~w4708;
assign w5525 = pi145 & ~w4842;
assign w5526 = w5041 & ~w5525;
assign w5527 = w5038 & ~w5041;
assign w5528 = ~w5188 & ~w5526;
assign w5529 = ~w5527 & w5528;
assign w5530 = ~w5038 & w5041;
assign w5531 = ~pi146 & ~w4842;
assign w5532 = w4845 & w5531;
assign w5533 = ~w5530 & ~w5532;
assign w5534 = w5188 & ~w5533;
assign w5535 = ~w5039 & ~w5529;
assign w5536 = ~w5534 & w5535;
assign w5537 = (w5034 & ~w5185) | (w5034 & w16171) | (~w5185 & w16171);
assign w5538 = ~w5187 & ~w5537;
assign w5539 = ~w5536 & w5538;
assign w5540 = w5536 & ~w5538;
assign w5541 = ~w5539 & ~w5540;
assign w5542 = pi147 & pi258;
assign w5543 = (~w5045 & ~w5182) | (~w5045 & w15885) | (~w5182 & w15885);
assign w5544 = pi143 & pi262;
assign w5545 = (~w5162 & ~w5163) | (~w5162 & w15886) | (~w5163 & w15886);
assign w5546 = pi140 & pi265;
assign w5547 = pi137 & pi268;
assign w5548 = (~w5115 & w5119) | (~w5115 & w16589) | (w5119 & w16589);
assign w5549 = pi134 & pi271;
assign w5550 = pi133 & pi272;
assign w5551 = pi131 & pi274;
assign w5552 = pi130 & pi275;
assign w5553 = pi129 & pi276;
assign w5554 = pi128 & pi277;
assign w5555 = ~w5062 & ~w5069;
assign w5556 = w5554 & w5555;
assign w5557 = ~w5554 & ~w5555;
assign w5558 = ~w5556 & ~w5557;
assign w5559 = w5553 & ~w5558;
assign w5560 = ~w5553 & w5558;
assign w5561 = ~w5559 & ~w5560;
assign w5562 = w5552 & ~w5561;
assign w5563 = ~w5552 & w5561;
assign w5564 = ~w5562 & ~w5563;
assign w5565 = ~w5071 & ~w5076;
assign w5566 = w5564 & ~w5565;
assign w5567 = ~w5564 & w5565;
assign w5568 = ~w5566 & ~w5567;
assign w5569 = ~w5551 & ~w5568;
assign w5570 = w5551 & w5568;
assign w5571 = ~w5569 & ~w5570;
assign w5572 = ~w5079 & ~w5083;
assign w5573 = w5571 & w5572;
assign w5574 = ~w5571 & ~w5572;
assign w5575 = ~w5573 & ~w5574;
assign w5576 = ~w5085 & ~w5091;
assign w5577 = (w5575 & w5091) | (w5575 & w16172) | (w5091 & w16172);
assign w5578 = ~w5091 & w16173;
assign w5579 = ~w5577 & ~w5578;
assign w5580 = pi132 & pi273;
assign w5581 = ~w5579 & w5580;
assign w5582 = w5579 & ~w5580;
assign w5583 = ~w5581 & ~w5582;
assign w5584 = w5550 & ~w5583;
assign w5585 = ~w5550 & w5583;
assign w5586 = ~w5584 & ~w5585;
assign w5587 = w5056 & ~w5094;
assign w5588 = ~w5095 & ~w5587;
assign w5589 = w5586 & ~w5588;
assign w5590 = ~w5586 & w5588;
assign w5591 = ~w5589 & ~w5590;
assign w5592 = w5549 & w5591;
assign w5593 = ~w5549 & ~w5591;
assign w5594 = ~w5592 & ~w5593;
assign w5595 = (w5055 & ~w5100) | (w5055 & w16174) | (~w5100 & w16174);
assign w5596 = ~w5101 & ~w5595;
assign w5597 = w5594 & ~w5596;
assign w5598 = ~w5594 & w5596;
assign w5599 = ~w5597 & ~w5598;
assign w5600 = ~w5108 & w5110;
assign w5601 = (~w5107 & ~w5110) | (~w5107 & w16590) | (~w5110 & w16590);
assign w5602 = (~w5599 & w5600) | (~w5599 & w16175) | (w5600 & w16175);
assign w5603 = w5599 & w5601;
assign w5604 = ~w5602 & ~w5603;
assign w5605 = pi136 & pi269;
assign w5606 = pi135 & pi270;
assign w5607 = w5605 & ~w5606;
assign w5608 = ~w5605 & w5606;
assign w5609 = ~w5607 & ~w5608;
assign w5610 = w5604 & w5609;
assign w5611 = ~w5604 & ~w5609;
assign w5612 = ~w5610 & ~w5611;
assign w5613 = w5548 & w5612;
assign w5614 = ~w5548 & ~w5612;
assign w5615 = ~w5613 & ~w5614;
assign w5616 = ~w5547 & w5615;
assign w5617 = w5547 & ~w5615;
assign w5618 = ~w5616 & ~w5617;
assign w5619 = ~w5117 & w5125;
assign w5620 = ~w5128 & ~w5619;
assign w5621 = w5618 & w5620;
assign w5622 = ~w5618 & ~w5620;
assign w5623 = ~w5621 & ~w5622;
assign w5624 = ~w5135 & w15887;
assign w5625 = (w5623 & w5135) | (w5623 & w15888) | (w5135 & w15888);
assign w5626 = ~w5624 & ~w5625;
assign w5627 = pi139 & pi266;
assign w5628 = pi138 & pi267;
assign w5629 = w5627 & ~w5628;
assign w5630 = ~w5627 & w5628;
assign w5631 = ~w5629 & ~w5630;
assign w5632 = w5626 & w5631;
assign w5633 = ~w5626 & ~w5631;
assign w5634 = ~w5632 & ~w5633;
assign w5635 = (~w5138 & ~w5143) | (~w5138 & w17586) | (~w5143 & w17586);
assign w5636 = ~w5634 & w5635;
assign w5637 = w5634 & ~w5635;
assign w5638 = ~w5636 & ~w5637;
assign w5639 = ~w5546 & ~w5638;
assign w5640 = w5546 & w5638;
assign w5641 = ~w5639 & ~w5640;
assign w5642 = w5141 & ~w5149;
assign w5643 = ~w5150 & ~w5642;
assign w5644 = ~w5641 & ~w5643;
assign w5645 = w5641 & w5643;
assign w5646 = ~w5644 & ~w5645;
assign w5647 = (~w5154 & ~w5155) | (~w5154 & w15889) | (~w5155 & w15889);
assign w5648 = (~w15889 & w16397) | (~w15889 & w16398) | (w16397 & w16398);
assign w5649 = (w15889 & w16399) | (w15889 & w16400) | (w16399 & w16400);
assign w5650 = ~w5648 & ~w5649;
assign w5651 = pi142 & pi263;
assign w5652 = pi141 & pi264;
assign w5653 = w5651 & ~w5652;
assign w5654 = ~w5651 & w5652;
assign w5655 = ~w5653 & ~w5654;
assign w5656 = w5650 & w5655;
assign w5657 = ~w5650 & ~w5655;
assign w5658 = ~w5656 & ~w5657;
assign w5659 = ~w5545 & w5658;
assign w5660 = w5545 & ~w5658;
assign w5661 = ~w5659 & ~w5660;
assign w5662 = w5544 & ~w5661;
assign w5663 = ~w5544 & w5661;
assign w5664 = ~w5662 & ~w5663;
assign w5665 = ~w5170 & ~w5179;
assign w5666 = ~w5171 & ~w5665;
assign w5667 = w5664 & w5666;
assign w5668 = ~w5664 & ~w5666;
assign w5669 = ~w5667 & ~w5668;
assign w5670 = w5543 & w5669;
assign w5671 = ~w5543 & ~w5669;
assign w5672 = ~w5670 & ~w5671;
assign w5673 = pi145 & pi260;
assign w5674 = pi144 & pi261;
assign w5675 = w5673 & ~w5674;
assign w5676 = ~w5673 & w5674;
assign w5677 = ~w5675 & ~w5676;
assign w5678 = w5672 & w5677;
assign w5679 = ~w5672 & ~w5677;
assign w5680 = ~w5678 & ~w5679;
assign w5681 = w5542 & ~w5680;
assign w5682 = ~w5542 & w5680;
assign w5683 = ~w5681 & ~w5682;
assign w5684 = pi145 & w4842;
assign w5685 = ~w5185 & w5684;
assign w5686 = w5185 & ~w5684;
assign w5687 = ~w5685 & ~w5686;
assign w5688 = pi259 & ~w5687;
assign w5689 = ~w5034 & w5185;
assign w5690 = pi258 & ~pi259;
assign w5691 = ~w5525 & w5690;
assign w5692 = ~w5185 & ~w5691;
assign w5693 = ~w5689 & ~w5692;
assign w5694 = ~w516 & ~w5693;
assign w5695 = ~w5688 & w5694;
assign w5696 = ~w5042 & w5526;
assign w5697 = ~w5042 & ~w5532;
assign w5698 = pi146 & w4842;
assign w5699 = ~w5531 & ~w5698;
assign w5700 = w458 & ~w5699;
assign w5701 = ~w5697 & ~w5700;
assign w5702 = ~w5696 & ~w5701;
assign w5703 = w5185 & w5702;
assign w5704 = ~w5185 & ~w5702;
assign w5705 = ~w5703 & ~w5704;
assign w5706 = ~w5695 & w16591;
assign w5707 = (w5705 & w5695) | (w5705 & w16592) | (w5695 & w16592);
assign w5708 = ~w5706 & ~w5707;
assign w5709 = w5683 & ~w5708;
assign w5710 = ~w5683 & w5708;
assign w5711 = ~w5709 & ~w5710;
assign w5712 = w5541 & w5711;
assign w5713 = ~w5541 & ~w5711;
assign w5714 = ~w5712 & ~w5713;
assign w5715 = pi322 & w5714;
assign w5716 = pi323 & w5194;
assign w5717 = (~w5199 & ~w5194) | (~w5199 & w16593) | (~w5194 & w16593);
assign w5718 = ~w5197 & ~w5717;
assign w5719 = w5716 & w5718;
assign w5720 = ~w5716 & ~w5718;
assign w5721 = ~w5719 & ~w5720;
assign w5722 = w5715 & w5721;
assign w5723 = ~w5715 & ~w5721;
assign w5724 = ~w5722 & ~w5723;
assign w5725 = pi324 & ~w4854;
assign w5726 = w5200 & w5206;
assign w5727 = ~w5513 & ~w5726;
assign w5728 = w5725 & ~w5727;
assign w5729 = ~w5725 & w5727;
assign w5730 = ~w5728 & ~w5729;
assign w5731 = w5724 & w5730;
assign w5732 = ~w5724 & ~w5730;
assign w5733 = ~w5731 & ~w5732;
assign w5734 = ~w5020 & ~w5516;
assign w5735 = w5733 & ~w5734;
assign w5736 = ~w5733 & w5734;
assign w5737 = ~w5735 & ~w5736;
assign w5738 = w5524 & ~w5737;
assign w5739 = ~w5524 & w5737;
assign w5740 = ~w5738 & ~w5739;
assign w5741 = w5523 & w5740;
assign w5742 = ~w5523 & ~w5740;
assign w5743 = ~w5741 & ~w5742;
assign w5744 = w5509 & w5743;
assign w5745 = ~w5509 & ~w5743;
assign w5746 = ~w5744 & ~w5745;
assign w5747 = pi328 & ~w3183;
assign w5748 = ~w5222 & ~w5225;
assign w5749 = w5747 & ~w5748;
assign w5750 = ~w5747 & w5748;
assign w5751 = ~w5749 & ~w5750;
assign w5752 = w5746 & w5751;
assign w5753 = ~w5746 & ~w5751;
assign w5754 = ~w5752 & ~w5753;
assign w5755 = ~w5013 & ~w5229;
assign w5756 = pi329 & w2698;
assign w5757 = w5755 & ~w5756;
assign w5758 = ~w5755 & w5756;
assign w5759 = ~w5757 & ~w5758;
assign w5760 = w5754 & w5759;
assign w5761 = ~w5754 & ~w5759;
assign w5762 = ~w5760 & ~w5761;
assign w5763 = w5504 & w5762;
assign w5764 = ~w5504 & ~w5762;
assign w5765 = ~w5763 & ~w5764;
assign w5766 = w5496 & w5765;
assign w5767 = ~w5496 & ~w5765;
assign w5768 = ~w5766 & ~w5767;
assign w5769 = pi332 & ~w1865;
assign w5770 = ~w5000 & ~w5238;
assign w5771 = w5769 & w5770;
assign w5772 = ~w5769 & ~w5770;
assign w5773 = ~w5771 & ~w5772;
assign w5774 = w5768 & ~w5773;
assign w5775 = ~w5768 & w5773;
assign w5776 = ~w5774 & ~w5775;
assign w5777 = w5491 & ~w5776;
assign w5778 = ~w5491 & w5776;
assign w5779 = ~w5777 & ~w5778;
assign w5780 = w5486 & w5779;
assign w5781 = ~w5486 & ~w5779;
assign w5782 = ~w5780 & ~w5781;
assign w5783 = ~w5248 & ~w5250;
assign w5784 = ~w5782 & w5783;
assign w5785 = w5782 & ~w5783;
assign w5786 = ~w5784 & ~w5785;
assign w5787 = ~w5481 & w5786;
assign w5788 = w5481 & ~w5786;
assign w5789 = ~w5787 & ~w5788;
assign w5790 = pi336 & ~w955;
assign w5791 = ~w4984 & ~w5253;
assign w5792 = w5790 & ~w5791;
assign w5793 = ~w5790 & w5791;
assign w5794 = ~w5792 & ~w5793;
assign w5795 = w5789 & ~w5794;
assign w5796 = ~w5789 & w5794;
assign w5797 = ~w5795 & ~w5796;
assign w5798 = w5480 & w5797;
assign w5799 = ~w5480 & ~w5797;
assign w5800 = ~w5798 & ~w5799;
assign w5801 = w5475 & w5800;
assign w5802 = ~w5475 & ~w5800;
assign w5803 = ~w5801 & ~w5802;
assign w5804 = pi339 & ~w537;
assign w5805 = ~w4971 & ~w5262;
assign w5806 = w5804 & ~w5805;
assign w5807 = ~w5804 & w5805;
assign w5808 = ~w5806 & ~w5807;
assign w5809 = ~w5803 & ~w5808;
assign w5810 = w5803 & w5808;
assign w5811 = ~w5809 & ~w5810;
assign w5812 = w5469 & w5811;
assign w5813 = ~w5469 & ~w5811;
assign w5814 = ~w5812 & ~w5813;
assign w5815 = w5465 & w5814;
assign w5816 = ~w5465 & ~w5814;
assign w5817 = ~w5815 & ~w5816;
assign w5818 = ~w5269 & ~w5272;
assign w5819 = ~w5817 & ~w5818;
assign w5820 = w5817 & w5818;
assign w5821 = ~w5819 & ~w5820;
assign w5822 = pi277 & w5821;
assign w5823 = ~pi277 & ~w5821;
assign w5824 = ~w5822 & ~w5823;
assign w5825 = ~pi129 & w5448;
assign w5826 = pi303 & w464;
assign w5827 = ~w5448 & ~w5826;
assign w5828 = ~w5825 & ~w5827;
assign w5829 = pi304 & ~w653;
assign w5830 = pi305 & w709;
assign w5831 = pi306 & w698;
assign w5832 = ~w5419 & ~w5423;
assign w5833 = ~w5831 & w5832;
assign w5834 = w5831 & ~w5832;
assign w5835 = ~w5833 & ~w5834;
assign w5836 = pi307 & w855;
assign w5837 = pi308 & w1159;
assign w5838 = pi309 & w1220;
assign w5839 = pi310 & w1420;
assign w5840 = (~w5391 & ~w5393) | (~w5391 & w16176) | (~w5393 & w16176);
assign w5841 = w5839 & ~w5840;
assign w5842 = ~w5839 & w5840;
assign w5843 = ~w5841 & ~w5842;
assign w5844 = pi311 & w1693;
assign w5845 = pi312 & w1954;
assign w5846 = ~w5377 & ~w5381;
assign w5847 = pi313 & ~w2473;
assign w5848 = pi314 & w2801;
assign w5849 = pi315 & w2925;
assign w5850 = pi316 & w3304;
assign w5851 = ~w5339 & ~w5342;
assign w5852 = ~w5331 & ~w5335;
assign w5853 = ~w4382 & w5325;
assign w5854 = pi319 & w4539;
assign w5855 = pi320 & w5316;
assign w5856 = ~pi147 & w5310;
assign w5857 = pi147 & ~w5310;
assign w5858 = ~w5856 & ~w5857;
assign w5859 = ~w5311 & ~w5314;
assign w5860 = w5858 & w5859;
assign w5861 = ~w5858 & ~w5859;
assign w5862 = ~w5860 & ~w5861;
assign w5863 = pi321 & w5862;
assign w5864 = ~w5320 & ~w5322;
assign w5865 = ~w5863 & w5864;
assign w5866 = w5863 & ~w5864;
assign w5867 = ~w5865 & ~w5866;
assign w5868 = w5855 & w5867;
assign w5869 = ~w5855 & ~w5867;
assign w5870 = ~w5868 & ~w5869;
assign w5871 = w5854 & w5870;
assign w5872 = ~w5854 & ~w5870;
assign w5873 = ~w5871 & ~w5872;
assign w5874 = w4382 & w5326;
assign w5875 = ~w5873 & ~w5874;
assign w5876 = pi318 & ~w5875;
assign w5877 = ~w5853 & ~w5876;
assign w5878 = ~pi319 & ~w5325;
assign w5879 = ~w5326 & ~w5853;
assign w5880 = ~w5878 & w5879;
assign w5881 = w5873 & ~w5880;
assign w5882 = ~w5877 & ~w5881;
assign w5883 = ~w5300 & ~w5325;
assign w5884 = pi318 & w4382;
assign w5885 = ~w5873 & ~w5884;
assign w5886 = w5873 & w5884;
assign w5887 = ~w5885 & ~w5886;
assign w5888 = w5883 & w5887;
assign w5889 = ~w5326 & ~w5883;
assign w5890 = w5873 & w5889;
assign w5891 = ~w5873 & ~w5889;
assign w5892 = ~w5890 & ~w5891;
assign w5893 = ~pi318 & ~w5329;
assign w5894 = w5892 & w5893;
assign w5895 = ~w5882 & ~w5888;
assign w5896 = ~w5894 & w5895;
assign w5897 = ~w5852 & w5896;
assign w5898 = w5852 & ~w5896;
assign w5899 = ~w5897 & ~w5898;
assign w5900 = w5851 & ~w5899;
assign w5901 = ~w5851 & w5899;
assign w5902 = ~w5900 & ~w5901;
assign w5903 = pi317 & w3710;
assign w5904 = ~w5902 & w5903;
assign w5905 = w5902 & ~w5903;
assign w5906 = ~w5904 & ~w5905;
assign w5907 = (w5362 & w16177) | (w5362 & w16178) | (w16177 & w16178);
assign w5908 = ~w5906 & w5907;
assign w5909 = w5906 & ~w5907;
assign w5910 = ~w5908 & ~w5909;
assign w5911 = w5850 & w5910;
assign w5912 = ~w5850 & ~w5910;
assign w5913 = ~w5911 & ~w5912;
assign w5914 = w5849 & w5913;
assign w5915 = ~w5849 & ~w5913;
assign w5916 = ~w5914 & ~w5915;
assign w5917 = ~w5295 & ~w5365;
assign w5918 = w5916 & w5917;
assign w5919 = ~w5916 & ~w5917;
assign w5920 = ~w5918 & ~w5919;
assign w5921 = w5848 & ~w5920;
assign w5922 = ~w5848 & w5920;
assign w5923 = ~w5921 & ~w5922;
assign w5924 = ~w5368 & ~w5372;
assign w5925 = w5923 & w5924;
assign w5926 = ~w5923 & ~w5924;
assign w5927 = ~w5925 & ~w5926;
assign w5928 = ~w5847 & ~w5927;
assign w5929 = w5847 & w5927;
assign w5930 = ~w5928 & ~w5929;
assign w5931 = ~w5288 & ~w5374;
assign w5932 = ~w5930 & w5931;
assign w5933 = w5930 & ~w5931;
assign w5934 = ~w5932 & ~w5933;
assign w5935 = w5846 & w5934;
assign w5936 = ~w5846 & ~w5934;
assign w5937 = ~w5935 & ~w5936;
assign w5938 = w5845 & w5937;
assign w5939 = ~w5845 & ~w5937;
assign w5940 = ~w5938 & ~w5939;
assign w5941 = w5844 & w5940;
assign w5942 = ~w5844 & ~w5940;
assign w5943 = ~w5941 & ~w5942;
assign w5944 = ~w5385 & ~w5388;
assign w5945 = w5943 & ~w5944;
assign w5946 = ~w5943 & w5944;
assign w5947 = ~w5945 & ~w5946;
assign w5948 = w5843 & ~w5947;
assign w5949 = ~w5843 & w5947;
assign w5950 = ~w5948 & ~w5949;
assign w5951 = ~w5838 & w5950;
assign w5952 = w5838 & ~w5950;
assign w5953 = ~w5951 & ~w5952;
assign w5954 = ~w5400 & ~w5402;
assign w5955 = w5953 & ~w5954;
assign w5956 = ~w5953 & w5954;
assign w5957 = ~w5955 & ~w5956;
assign w5958 = w5837 & w5957;
assign w5959 = ~w5837 & ~w5957;
assign w5960 = ~w5958 & ~w5959;
assign w5961 = ~w5405 & ~w5409;
assign w5962 = w5960 & w5961;
assign w5963 = ~w5960 & ~w5961;
assign w5964 = ~w5962 & ~w5963;
assign w5965 = w5836 & ~w5964;
assign w5966 = ~w5836 & w5964;
assign w5967 = ~w5965 & ~w5966;
assign w5968 = ~w5414 & ~w5417;
assign w5969 = w5967 & w5968;
assign w5970 = ~w5967 & ~w5968;
assign w5971 = ~w5969 & ~w5970;
assign w5972 = w5835 & w5971;
assign w5973 = ~w5835 & ~w5971;
assign w5974 = ~w5972 & ~w5973;
assign w5975 = ~w5830 & ~w5974;
assign w5976 = w5830 & w5974;
assign w5977 = ~w5975 & ~w5976;
assign w5978 = pi130 & pi305;
assign w5979 = ~w5432 & w5978;
assign w5980 = w4649 & w5438;
assign w5981 = ~w5979 & ~w5980;
assign w5982 = ~w5442 & w5981;
assign w5983 = ~w5977 & w5982;
assign w5984 = w5977 & ~w5982;
assign w5985 = ~w5983 & ~w5984;
assign w5986 = ~w5278 & ~w5445;
assign w5987 = w5985 & ~w5986;
assign w5988 = ~w5985 & w5986;
assign w5989 = ~w5987 & ~w5988;
assign w5990 = w5829 & w5989;
assign w5991 = ~w5829 & ~w5989;
assign w5992 = ~w5990 & ~w5991;
assign w5993 = w5828 & w5992;
assign w5994 = ~w5828 & ~w5992;
assign w5995 = ~w5993 & ~w5994;
assign w5996 = pi128 & pi302;
assign w5997 = w5995 & w5996;
assign w5998 = ~w5995 & ~w5996;
assign w5999 = ~w5997 & ~w5998;
assign w6000 = ~w5451 & ~w5455;
assign w6001 = ~w5999 & ~w6000;
assign w6002 = w5999 & w6000;
assign w6003 = ~w6001 & ~w6002;
assign w6004 = ~w5824 & ~w6003;
assign w6005 = w5824 & w6003;
assign w6006 = ~w135 & ~w6004;
assign w6007 = ~w6005 & w6006;
assign w6008 = pi161 & ~w5464;
assign w6009 = ~w6007 & w6008;
assign w6010 = ~pi160 & ~w5463;
assign w6011 = ~w6009 & w6010;
assign w6012 = ~pi084 & ~pi161;
assign w6013 = pi278 & w135;
assign w6014 = pi342 & w456;
assign w6015 = pi341 & w466;
assign w6016 = ~w5815 & ~w6015;
assign w6017 = w466 & w5815;
assign w6018 = ~w6016 & ~w6017;
assign w6019 = pi340 & ~w537;
assign w6020 = ~w5468 & ~w5812;
assign w6021 = ~w5806 & ~w5810;
assign w6022 = pi339 & ~w615;
assign w6023 = ~w6021 & w6022;
assign w6024 = w6021 & ~w6022;
assign w6025 = ~w6023 & ~w6024;
assign w6026 = ~w5472 & ~w5801;
assign w6027 = pi338 & ~w793;
assign w6028 = ~w6026 & w6027;
assign w6029 = w6026 & ~w6027;
assign w6030 = ~w6028 & ~w6029;
assign w6031 = pi336 & w1101;
assign w6032 = ~w5792 & w6031;
assign w6033 = pi335 & w6032;
assign w6034 = ~w5481 & ~w6031;
assign w6035 = ~w5793 & w6034;
assign w6036 = ~w6033 & ~w6035;
assign w6037 = w5786 & ~w6036;
assign w6038 = ~w5792 & ~w6031;
assign w6039 = ~w5793 & w6031;
assign w6040 = ~w6038 & ~w6039;
assign w6041 = ~pi335 & ~w5786;
assign w6042 = w6032 & w6041;
assign w6043 = ~w6040 & ~w6042;
assign w6044 = ~w6037 & w6043;
assign w6045 = pi335 & w1339;
assign w6046 = ~w6044 & w6045;
assign w6047 = w6044 & ~w6045;
assign w6048 = ~w6046 & ~w6047;
assign w6049 = (~w5784 & ~w5786) | (~w5784 & w16594) | (~w5786 & w16594);
assign w6050 = (~w5479 & ~w5797) | (~w5479 & w16595) | (~w5797 & w16595);
assign w6051 = (w5797 & w17587) | (w5797 & w17588) | (w17587 & w17588);
assign w6052 = ~w6049 & w6050;
assign w6053 = ~w6051 & ~w6052;
assign w6054 = w6048 & w6053;
assign w6055 = ~w6048 & ~w6053;
assign w6056 = ~w6054 & ~w6055;
assign w6057 = pi337 & ~w955;
assign w6058 = pi334 & w1602;
assign w6059 = (w5779 & w17589) | (w5779 & w17590) | (w17589 & w17590);
assign w6060 = ~w6058 & w17681;
assign w6061 = ~w6059 & ~w6060;
assign w6062 = pi333 & ~w1865;
assign w6063 = w6062 & w17682;
assign w6064 = (w5776 & w17591) | (w5776 & w17592) | (w17591 & w17592);
assign w6065 = ~w6063 & ~w6064;
assign w6066 = pi332 & ~w2170;
assign w6067 = (~w5772 & w5768) | (~w5772 & w16179) | (w5768 & w16179);
assign w6068 = (w5768 & w16598) | (w5768 & w16599) | (w16598 & w16599);
assign w6069 = w6066 & ~w6067;
assign w6070 = ~w6068 & ~w6069;
assign w6071 = pi328 & ~w3568;
assign w6072 = ~w6071 & w17683;
assign w6073 = (w5746 & w16600) | (w5746 & w16601) | (w16600 & w16601);
assign w6074 = ~w6072 & ~w6073;
assign w6075 = pi327 & w3979;
assign w6076 = ~w6075 & w17684;
assign w6077 = (w5743 & w16602) | (w5743 & w16603) | (w16602 & w16603);
assign w6078 = ~w6076 & ~w6077;
assign w6079 = ~w5522 & ~w5741;
assign w6080 = pi324 & w5194;
assign w6081 = (w5538 & w5695) | (w5538 & w15890) | (w5695 & w15890);
assign w6082 = ~w5695 & w15891;
assign w6083 = ~w6081 & ~w6082;
assign w6084 = w5681 & ~w6083;
assign w6085 = w5542 & w5680;
assign w6086 = w6083 & w6085;
assign w6087 = ~w6084 & ~w6086;
assign w6088 = w5683 & w6083;
assign w6089 = ~w5683 & ~w6083;
assign w6090 = ~w6088 & ~w6089;
assign w6091 = w6087 & ~w6090;
assign w6092 = ~w5536 & ~w6090;
assign w6093 = (~w5705 & ~w6090) | (~w5705 & w16182) | (~w6090 & w16182);
assign w6094 = ~w6092 & ~w6093;
assign w6095 = w6091 & ~w6094;
assign w6096 = ~w6091 & w6094;
assign w6097 = ~w6095 & ~w6096;
assign w6098 = ~pi259 & ~w5693;
assign w6099 = pi146 & pi260;
assign w6100 = w6098 & w6099;
assign w6101 = ~w5538 & w5680;
assign w6102 = pi146 & w458;
assign w6103 = w5687 & w6102;
assign w6104 = (~w6103 & w5680) | (~w6103 & w16604) | (w5680 & w16604);
assign w6105 = (w6099 & ~w5680) | (w6099 & w16183) | (~w5680 & w16183);
assign w6106 = (~w6100 & ~w6104) | (~w6100 & w16184) | (~w6104 & w16184);
assign w6107 = pi146 & ~pi260;
assign w6108 = ~w6098 & w6107;
assign w6109 = (w6108 & ~w6104) | (w6108 & w16185) | (~w6104 & w16185);
assign w6110 = w6106 & ~w6109;
assign w6111 = pi145 & pi261;
assign w6112 = pi144 & pi262;
assign w6113 = (~w5663 & w5666) | (~w5663 & w15892) | (w5666 & w15892);
assign w6114 = (w15892 & w16401) | (w15892 & w16402) | (w16401 & w16402);
assign w6115 = (~w15892 & w16403) | (~w15892 & w16404) | (w16403 & w16404);
assign w6116 = ~w6114 & ~w6115;
assign w6117 = pi141 & pi265;
assign w6118 = (~w5639 & ~w5643) | (~w5639 & w17593) | (~w5643 & w17593);
assign w6119 = pi139 & pi267;
assign w6120 = pi138 & pi268;
assign w6121 = ~w5617 & ~w5621;
assign w6122 = pi136 & pi270;
assign w6123 = pi135 & pi271;
assign w6124 = pi134 & pi272;
assign w6125 = ~w5592 & w5596;
assign w6126 = pi133 & pi273;
assign w6127 = pi132 & pi274;
assign w6128 = pi131 & pi275;
assign w6129 = ~w5562 & ~w5566;
assign w6130 = pi130 & pi276;
assign w6131 = pi129 & ~w5557;
assign w6132 = ~pi130 & ~w6131;
assign w6133 = ~pi276 & ~w5556;
assign w6134 = ~w6132 & ~w6133;
assign w6135 = pi128 & pi278;
assign w6136 = pi129 & pi277;
assign w6137 = ~w6135 & w6136;
assign w6138 = w6135 & ~w6136;
assign w6139 = ~w6137 & ~w6138;
assign w6140 = ~w6134 & ~w6139;
assign w6141 = ~w646 & ~w6132;
assign w6142 = pi276 & ~w6141;
assign w6143 = ~w6133 & w6139;
assign w6144 = ~w6142 & w6143;
assign w6145 = ~w6130 & ~w6140;
assign w6146 = ~w6144 & w6145;
assign w6147 = w6131 & ~w6139;
assign w6148 = ~w6131 & w6139;
assign w6149 = w6130 & ~w6147;
assign w6150 = ~w6148 & w6149;
assign w6151 = ~w6146 & ~w6150;
assign w6152 = ~w6129 & ~w6151;
assign w6153 = w6129 & w6151;
assign w6154 = ~w6152 & ~w6153;
assign w6155 = ~w6128 & w6154;
assign w6156 = w6128 & ~w6154;
assign w6157 = ~w6155 & ~w6156;
assign w6158 = ~w5569 & ~w5573;
assign w6159 = w6157 & ~w6158;
assign w6160 = ~w6157 & w6158;
assign w6161 = ~w6159 & ~w6160;
assign w6162 = ~w6127 & w6161;
assign w6163 = w6127 & ~w6161;
assign w6164 = ~w6162 & ~w6163;
assign w6165 = (~w5577 & ~w5579) | (~w5577 & w15893) | (~w5579 & w15893);
assign w6166 = ~w6164 & ~w6165;
assign w6167 = w6164 & w6165;
assign w6168 = ~w6166 & ~w6167;
assign w6169 = w6126 & w6168;
assign w6170 = ~w6126 & ~w6168;
assign w6171 = ~w6169 & ~w6170;
assign w6172 = ~w5585 & ~w5588;
assign w6173 = ~w5584 & ~w6172;
assign w6174 = w6171 & ~w6173;
assign w6175 = ~w6171 & w6173;
assign w6176 = ~w6174 & ~w6175;
assign w6177 = ~w6125 & w15894;
assign w6178 = (~w6176 & w6125) | (~w6176 & w15895) | (w6125 & w15895);
assign w6179 = ~w6177 & ~w6178;
assign w6180 = w6124 & w6179;
assign w6181 = ~w6124 & ~w6179;
assign w6182 = ~w6180 & ~w6181;
assign w6183 = ~w6123 & ~w6182;
assign w6184 = w6123 & w6182;
assign w6185 = ~w6183 & ~w6184;
assign w6186 = (~w5606 & ~w5601) | (~w5606 & w15896) | (~w5601 & w15896);
assign w6187 = ~w5602 & ~w6186;
assign w6188 = w6185 & ~w6187;
assign w6189 = ~w6185 & w6187;
assign w6190 = ~w6188 & ~w6189;
assign w6191 = w6122 & ~w6190;
assign w6192 = ~w6122 & w6190;
assign w6193 = ~w6191 & ~w6192;
assign w6194 = pi137 & pi269;
assign w6195 = ~w5605 & w5612;
assign w6196 = ~w5614 & ~w6195;
assign w6197 = w6194 & ~w6196;
assign w6198 = ~w6194 & w6196;
assign w6199 = ~w6197 & ~w6198;
assign w6200 = w6193 & ~w6199;
assign w6201 = ~w6193 & w6199;
assign w6202 = ~w6200 & ~w6201;
assign w6203 = ~w6121 & ~w6202;
assign w6204 = w6121 & w6202;
assign w6205 = ~w6203 & ~w6204;
assign w6206 = w6120 & ~w6205;
assign w6207 = ~w6120 & w6205;
assign w6208 = ~w6206 & ~w6207;
assign w6209 = ~w5625 & ~w5628;
assign w6210 = ~w5624 & ~w6209;
assign w6211 = w6208 & ~w6210;
assign w6212 = ~w6208 & w6210;
assign w6213 = ~w6211 & ~w6212;
assign w6214 = ~w6119 & w6213;
assign w6215 = w6119 & ~w6213;
assign w6216 = ~w6214 & ~w6215;
assign w6217 = pi140 & pi266;
assign w6218 = w5627 & w5634;
assign w6219 = ~w5636 & ~w6218;
assign w6220 = w6217 & ~w6219;
assign w6221 = ~w6217 & w6219;
assign w6222 = ~w6220 & ~w6221;
assign w6223 = w6216 & ~w6222;
assign w6224 = ~w6216 & w6222;
assign w6225 = ~w6223 & ~w6224;
assign w6226 = w6118 & ~w6225;
assign w6227 = ~w6118 & w6225;
assign w6228 = ~w6226 & ~w6227;
assign w6229 = w6117 & w6228;
assign w6230 = ~w6117 & ~w6228;
assign w6231 = ~w6229 & ~w6230;
assign w6232 = (~w5652 & ~w5647) | (~w5652 & w15897) | (~w5647 & w15897);
assign w6233 = ~w5648 & ~w6232;
assign w6234 = w6231 & w6233;
assign w6235 = ~w6231 & ~w6233;
assign w6236 = ~w6234 & ~w6235;
assign w6237 = ~w5651 & w5658;
assign w6238 = ~w5660 & ~w6237;
assign w6239 = ~w5660 & w16605;
assign w6240 = (~w6236 & w5660) | (~w6236 & w16606) | (w5660 & w16606);
assign w6241 = ~w6239 & ~w6240;
assign w6242 = pi142 & pi264;
assign w6243 = pi143 & pi263;
assign w6244 = ~w6242 & w6243;
assign w6245 = w6242 & ~w6243;
assign w6246 = ~w6244 & ~w6245;
assign w6247 = w6241 & w6246;
assign w6248 = ~w6241 & ~w6246;
assign w6249 = ~w6247 & ~w6248;
assign w6250 = ~w6116 & ~w6249;
assign w6251 = w6116 & w6249;
assign w6252 = ~w6250 & ~w6251;
assign w6253 = (~w5674 & ~w5669) | (~w5674 & w16405) | (~w5669 & w16405);
assign w6254 = ~w5671 & ~w6253;
assign w6255 = w6252 & w6254;
assign w6256 = ~w6252 & ~w6254;
assign w6257 = ~w6255 & ~w6256;
assign w6258 = w6111 & w6257;
assign w6259 = ~w6111 & ~w6257;
assign w6260 = ~w6258 & ~w6259;
assign w6261 = ~w5672 & ~w5674;
assign w6262 = w5672 & w5674;
assign w6263 = ~w6261 & ~w6262;
assign w6264 = (~w5538 & w6263) | (~w5538 & w16186) | (w6263 & w16186);
assign w6265 = w5673 & w6263;
assign w6266 = ~w6264 & ~w6265;
assign w6267 = w6260 & ~w6266;
assign w6268 = ~w6260 & w6266;
assign w6269 = ~w6267 & ~w6268;
assign w6270 = w6110 & ~w6269;
assign w6271 = ~w6110 & w6269;
assign w6272 = ~w6270 & ~w6271;
assign w6273 = pi148 & pi258;
assign w6274 = pi147 & pi259;
assign w6275 = w6273 & ~w6274;
assign w6276 = ~w6273 & w6274;
assign w6277 = ~w6275 & ~w6276;
assign w6278 = ~w6272 & w6277;
assign w6279 = w6272 & ~w6277;
assign w6280 = ~w6278 & ~w6279;
assign w6281 = w6097 & w6280;
assign w6282 = ~w6097 & ~w6280;
assign w6283 = ~w6281 & ~w6282;
assign w6284 = pi322 & w6283;
assign w6285 = pi323 & w5714;
assign w6286 = (~w5719 & ~w5715) | (~w5719 & w15898) | (~w5715 & w15898);
assign w6287 = w6285 & ~w6286;
assign w6288 = ~w6285 & w6286;
assign w6289 = ~w6287 & ~w6288;
assign w6290 = w6284 & w6289;
assign w6291 = ~w6284 & ~w6289;
assign w6292 = ~w6290 & ~w6291;
assign w6293 = w6080 & w6292;
assign w6294 = ~w6080 & ~w6292;
assign w6295 = ~w6293 & ~w6294;
assign w6296 = ~w5728 & ~w5731;
assign w6297 = ~w6295 & w6296;
assign w6298 = w6295 & ~w6296;
assign w6299 = ~w6297 & ~w6298;
assign w6300 = pi325 & ~w4854;
assign w6301 = ~w5516 & w16406;
assign w6302 = (~w5524 & w5516) | (~w5524 & w16407) | (w5516 & w16407);
assign w6303 = ~w6300 & w17685;
assign w6304 = (w5733 & w16408) | (w5733 & w16409) | (w16408 & w16409);
assign w6305 = ~w6303 & ~w6304;
assign w6306 = pi326 & ~w4708;
assign w6307 = w6305 & ~w6306;
assign w6308 = ~w6305 & w6306;
assign w6309 = ~w6307 & ~w6308;
assign w6310 = w6299 & w6309;
assign w6311 = ~w6299 & ~w6309;
assign w6312 = ~w6310 & ~w6311;
assign w6313 = w6079 & ~w6312;
assign w6314 = ~w6079 & w6312;
assign w6315 = ~w6313 & ~w6314;
assign w6316 = w6078 & w6315;
assign w6317 = ~w6078 & ~w6315;
assign w6318 = ~w6316 & ~w6317;
assign w6319 = w6074 & w6318;
assign w6320 = ~w6074 & ~w6318;
assign w6321 = ~w6319 & ~w6320;
assign w6322 = ~w5758 & ~w5760;
assign w6323 = w6321 & w6322;
assign w6324 = ~w6321 & ~w6322;
assign w6325 = ~w6323 & ~w6324;
assign w6326 = pi330 & w2698;
assign w6327 = pi330 & w5499;
assign w6328 = (w5762 & w16410) | (w5762 & w16411) | (w16410 & w16411);
assign w6329 = ~w6326 & w17686;
assign w6330 = ~w6328 & ~w6329;
assign w6331 = w6325 & w6330;
assign w6332 = ~w6325 & ~w6330;
assign w6333 = ~w6331 & ~w6332;
assign w6334 = ~w5495 & ~w5766;
assign w6335 = pi331 & ~w2373;
assign w6336 = pi329 & ~w3183;
assign w6337 = w6335 & ~w6336;
assign w6338 = ~w6335 & w6336;
assign w6339 = ~w6337 & ~w6338;
assign w6340 = (w15901 & ~w5765) | (w15901 & w16412) | (~w5765 & w16412);
assign w6341 = (w5765 & w16413) | (w5765 & w16414) | (w16413 & w16414);
assign w6342 = ~w6340 & ~w6341;
assign w6343 = w6333 & w6342;
assign w6344 = ~w6333 & ~w6342;
assign w6345 = ~w6343 & ~w6344;
assign w6346 = w6070 & w6345;
assign w6347 = ~w6070 & ~w6345;
assign w6348 = ~w6346 & ~w6347;
assign w6349 = w6065 & w6348;
assign w6350 = ~w6065 & ~w6348;
assign w6351 = ~w6349 & ~w6350;
assign w6352 = ~w6061 & ~w6351;
assign w6353 = w6061 & w6351;
assign w6354 = ~w6352 & ~w6353;
assign w6355 = ~w6057 & w6354;
assign w6356 = w6057 & ~w6354;
assign w6357 = ~w6355 & ~w6356;
assign w6358 = w6056 & w6357;
assign w6359 = ~w6056 & ~w6357;
assign w6360 = ~w6358 & ~w6359;
assign w6361 = w6030 & w6360;
assign w6362 = ~w6030 & ~w6360;
assign w6363 = ~w6361 & ~w6362;
assign w6364 = w6025 & ~w6363;
assign w6365 = ~w6025 & w6363;
assign w6366 = ~w6364 & ~w6365;
assign w6367 = ~w6020 & w6366;
assign w6368 = w6020 & ~w6366;
assign w6369 = ~w6367 & ~w6368;
assign w6370 = ~w6019 & w6369;
assign w6371 = w6019 & ~w6369;
assign w6372 = ~w6370 & ~w6371;
assign w6373 = w6018 & ~w6372;
assign w6374 = ~w6018 & w6372;
assign w6375 = ~w6373 & ~w6374;
assign w6376 = w6014 & w6375;
assign w6377 = ~w6014 & ~w6375;
assign w6378 = ~w6376 & ~w6377;
assign w6379 = ~w5819 & ~w5822;
assign w6380 = ~w6378 & ~w6379;
assign w6381 = w6378 & w6379;
assign w6382 = ~w6380 & ~w6381;
assign w6383 = pi278 & w6382;
assign w6384 = ~pi278 & ~w6382;
assign w6385 = ~w6383 & ~w6384;
assign w6386 = ~w6001 & ~w6005;
assign w6387 = ~w6385 & w6386;
assign w6388 = w6385 & ~w6386;
assign w6389 = ~w6387 & ~w6388;
assign w6390 = pi128 & pi301;
assign w6391 = pi302 & w464;
assign w6392 = ~w5997 & ~w6391;
assign w6393 = ~pi129 & w5997;
assign w6394 = ~w6392 & ~w6393;
assign w6395 = pi303 & ~w653;
assign w6396 = pi304 & w709;
assign w6397 = pi305 & w698;
assign w6398 = (~w5976 & ~w5977) | (~w5976 & w15903) | (~w5977 & w15903);
assign w6399 = pi306 & w855;
assign w6400 = pi307 & w1159;
assign w6401 = pi308 & w1220;
assign w6402 = (~w5952 & w5954) | (~w5952 & w16415) | (w5954 & w16415);
assign w6403 = pi309 & w1420;
assign w6404 = pi310 & w1693;
assign w6405 = pi311 & w1954;
assign w6406 = pi312 & ~w2473;
assign w6407 = pi314 & w2925;
assign w6408 = pi315 & w3304;
assign w6409 = (~w6408 & w5918) | (~w6408 & w15904) | (w5918 & w15904);
assign w6410 = ~w5918 & w15905;
assign w6411 = ~w6409 & ~w6410;
assign w6412 = pi316 & w3710;
assign w6413 = (w5892 & w5335) | (w5892 & w16416) | (w5335 & w16416);
assign w6414 = ~w5335 & w16417;
assign w6415 = pi319 & w5316;
assign w6416 = ~w5871 & ~w5890;
assign w6417 = pi320 & w5862;
assign w6418 = pi146 & pi148;
assign w6419 = ~pi147 & w6418;
assign w6420 = ~pi148 & w5857;
assign w6421 = pi145 & ~w6419;
assign w6422 = ~w6420 & w6421;
assign w6423 = ~pi147 & ~pi148;
assign w6424 = w5310 & w6423;
assign w6425 = pi147 & pi148;
assign w6426 = ~pi146 & w6425;
assign w6427 = ~pi145 & ~w6426;
assign w6428 = ~w6424 & w6427;
assign w6429 = ~w6422 & ~w6428;
assign w6430 = pi146 & ~w5856;
assign w6431 = ~w6423 & ~w6425;
assign w6432 = pi148 & ~w5310;
assign w6433 = ~w6431 & ~w6432;
assign w6434 = ~w6430 & ~w6433;
assign w6435 = pi146 & ~w6431;
assign w6436 = ~w6434 & ~w6435;
assign w6437 = ~w6429 & ~w6436;
assign w6438 = pi321 & w6437;
assign w6439 = ~w5855 & ~w5866;
assign w6440 = ~w5865 & ~w6439;
assign w6441 = ~w6438 & ~w6440;
assign w6442 = w6438 & w6440;
assign w6443 = ~w6441 & ~w6442;
assign w6444 = w6417 & ~w6443;
assign w6445 = ~w6417 & w6443;
assign w6446 = ~w6444 & ~w6445;
assign w6447 = ~w6416 & ~w6446;
assign w6448 = w6416 & w6446;
assign w6449 = ~w6447 & ~w6448;
assign w6450 = w6415 & w6449;
assign w6451 = ~w6415 & ~w6449;
assign w6452 = ~w6450 & ~w6451;
assign w6453 = ~w6414 & w6452;
assign w6454 = w4382 & w4539;
assign w6455 = ~w6413 & ~w6454;
assign w6456 = w6453 & ~w6455;
assign w6457 = ~w6413 & w6456;
assign w6458 = w6414 & ~w6452;
assign w6459 = ~w5884 & ~w6413;
assign w6460 = ~w6414 & w6459;
assign w6461 = (~w4539 & ~w6452) | (~w4539 & w16418) | (~w6452 & w16418);
assign w6462 = ~w6458 & w6461;
assign w6463 = ~w6460 & w6462;
assign w6464 = pi318 & w4539;
assign w6465 = w6452 & w6464;
assign w6466 = ~w6452 & ~w6464;
assign w6467 = w6459 & ~w6465;
assign w6468 = ~w6466 & w6467;
assign w6469 = ~w6463 & ~w6468;
assign w6470 = (w6464 & w6456) | (w6464 & w16419) | (w6456 & w16419);
assign w6471 = ~w6457 & ~w6470;
assign w6472 = w6469 & w6471;
assign w6473 = ~w5901 & ~w6472;
assign w6474 = w3710 & w6473;
assign w6475 = w4382 & w6474;
assign w6476 = pi317 & w4382;
assign w6477 = ~w6472 & w6476;
assign w6478 = w6472 & ~w6476;
assign w6479 = ~w5903 & ~w6477;
assign w6480 = ~w6478 & w6479;
assign w6481 = ~w6475 & ~w6480;
assign w6482 = ~w5900 & ~w6481;
assign w6483 = w5901 & w6472;
assign w6484 = ~w6473 & ~w6483;
assign w6485 = ~w4382 & ~w5905;
assign w6486 = w6484 & w6485;
assign w6487 = ~w5902 & w6476;
assign w6488 = ~w6484 & w6487;
assign w6489 = ~w6486 & ~w6488;
assign w6490 = ~w6482 & w6489;
assign w6491 = ~w6412 & w6490;
assign w6492 = w6412 & ~w6490;
assign w6493 = ~w6491 & ~w6492;
assign w6494 = ~w5908 & ~w5911;
assign w6495 = ~w6493 & ~w6494;
assign w6496 = w6493 & w6494;
assign w6497 = ~w6495 & ~w6496;
assign w6498 = w6411 & w6497;
assign w6499 = ~w6411 & ~w6497;
assign w6500 = ~w6498 & ~w6499;
assign w6501 = w6407 & ~w6500;
assign w6502 = ~w6407 & w6500;
assign w6503 = ~w6501 & ~w6502;
assign w6504 = ~w5921 & ~w5925;
assign w6505 = w6503 & ~w6504;
assign w6506 = ~w6503 & w6504;
assign w6507 = ~w6505 & ~w6506;
assign w6508 = pi313 & w2801;
assign w6509 = w6507 & w6508;
assign w6510 = ~w6507 & ~w6508;
assign w6511 = ~w6509 & ~w6510;
assign w6512 = w2473 & ~w5927;
assign w6513 = ~w5931 & ~w6512;
assign w6514 = ~w5929 & ~w6513;
assign w6515 = w6511 & w6514;
assign w6516 = ~w6511 & ~w6514;
assign w6517 = ~w6515 & ~w6516;
assign w6518 = ~w6406 & w6517;
assign w6519 = w6406 & ~w6517;
assign w6520 = ~w6518 & ~w6519;
assign w6521 = (~w5935 & ~w5937) | (~w5935 & w15906) | (~w5937 & w15906);
assign w6522 = w6520 & w6521;
assign w6523 = ~w6520 & ~w6521;
assign w6524 = ~w6522 & ~w6523;
assign w6525 = (~w5941 & ~w5943) | (~w5941 & w15907) | (~w5943 & w15907);
assign w6526 = w6524 & w6525;
assign w6527 = ~w6524 & ~w6525;
assign w6528 = ~w6526 & ~w6527;
assign w6529 = w6405 & ~w6528;
assign w6530 = ~w6405 & w6528;
assign w6531 = ~w6529 & ~w6530;
assign w6532 = (~w5842 & ~w5843) | (~w5842 & w15908) | (~w5843 & w15908);
assign w6533 = ~w6531 & w6532;
assign w6534 = w6531 & ~w6532;
assign w6535 = ~w6533 & ~w6534;
assign w6536 = w6404 & w6535;
assign w6537 = ~w6404 & ~w6535;
assign w6538 = ~w6536 & ~w6537;
assign w6539 = w6403 & w6538;
assign w6540 = ~w6403 & ~w6538;
assign w6541 = ~w6539 & ~w6540;
assign w6542 = w6402 & ~w6541;
assign w6543 = ~w6402 & w6541;
assign w6544 = ~w6542 & ~w6543;
assign w6545 = w6401 & w6544;
assign w6546 = ~w6401 & ~w6544;
assign w6547 = ~w6545 & ~w6546;
assign w6548 = ~w5959 & ~w5962;
assign w6549 = ~w6547 & w6548;
assign w6550 = w6547 & ~w6548;
assign w6551 = ~w6549 & ~w6550;
assign w6552 = (~w6551 & w5969) | (~w6551 & w16420) | (w5969 & w16420);
assign w6553 = ~w5969 & w16421;
assign w6554 = ~w6552 & ~w6553;
assign w6555 = w6400 & w6554;
assign w6556 = ~w6400 & ~w6554;
assign w6557 = ~w6555 & ~w6556;
assign w6558 = (w5835 & w16422) | (w5835 & w16423) | (w16422 & w16423);
assign w6559 = ~w6557 & w17687;
assign w6560 = ~w6558 & ~w6559;
assign w6561 = w6399 & ~w6560;
assign w6562 = ~w6399 & w6560;
assign w6563 = ~w6561 & ~w6562;
assign w6564 = ~w6398 & ~w6563;
assign w6565 = w6398 & w6563;
assign w6566 = ~w6564 & ~w6565;
assign w6567 = w6397 & w6566;
assign w6568 = ~w6397 & ~w6566;
assign w6569 = ~w6567 & ~w6568;
assign w6570 = w6396 & w6569;
assign w6571 = ~w6396 & ~w6569;
assign w6572 = ~w6570 & ~w6571;
assign w6573 = ~w5987 & ~w5990;
assign w6574 = ~w6572 & w6573;
assign w6575 = w6572 & ~w6573;
assign w6576 = ~w6574 & ~w6575;
assign w6577 = ~w5825 & ~w5993;
assign w6578 = w6576 & ~w6577;
assign w6579 = ~w6576 & w6577;
assign w6580 = ~w6578 & ~w6579;
assign w6581 = w6395 & ~w6580;
assign w6582 = ~w6395 & w6580;
assign w6583 = ~w6581 & ~w6582;
assign w6584 = w6394 & ~w6583;
assign w6585 = ~w6394 & w6583;
assign w6586 = ~w6584 & ~w6585;
assign w6587 = w6390 & ~w6586;
assign w6588 = ~w6390 & w6586;
assign w6589 = ~w6587 & ~w6588;
assign w6590 = ~w6389 & w6589;
assign w6591 = w6389 & ~w6589;
assign w6592 = ~w6590 & ~w6591;
assign w6593 = ~w135 & ~w6592;
assign w6594 = pi161 & ~w6013;
assign w6595 = ~w6593 & w6594;
assign w6596 = ~pi160 & ~w6012;
assign w6597 = ~w6595 & w6596;
assign w6598 = ~pi085 & ~pi161;
assign w6599 = pi128 & pi300;
assign w6600 = pi129 & ~pi301;
assign w6601 = ~w6587 & ~w6600;
assign w6602 = pi302 & ~w653;
assign w6603 = ~w6393 & ~w6584;
assign w6604 = ~w6602 & w6603;
assign w6605 = w6602 & ~w6603;
assign w6606 = ~w6604 & ~w6605;
assign w6607 = pi303 & w709;
assign w6608 = (~w6570 & ~w6572) | (~w6570 & w16424) | (~w6572 & w16424);
assign w6609 = pi304 & w698;
assign w6610 = ~w6608 & w6609;
assign w6611 = w6608 & ~w6609;
assign w6612 = ~w6610 & ~w6611;
assign w6613 = pi305 & w855;
assign w6614 = pi307 & w1220;
assign w6615 = pi308 & w1420;
assign w6616 = (~w6615 & w6550) | (~w6615 & w16425) | (w6550 & w16425);
assign w6617 = ~w6550 & w16426;
assign w6618 = ~w6616 & ~w6617;
assign w6619 = pi309 & w1693;
assign w6620 = pi311 & ~w2473;
assign w6621 = pi312 & w2801;
assign w6622 = (~w6621 & w6522) | (~w6621 & w16427) | (w6522 & w16427);
assign w6623 = ~w6522 & w16428;
assign w6624 = ~w6622 & ~w6623;
assign w6625 = pi314 & w3304;
assign w6626 = ~w6501 & ~w6505;
assign w6627 = w6625 & ~w6626;
assign w6628 = ~w6625 & w6626;
assign w6629 = ~w6627 & ~w6628;
assign w6630 = pi315 & w3710;
assign w6631 = pi316 & w4382;
assign w6632 = pi317 & w4539;
assign w6633 = pi318 & w5316;
assign w6634 = pi319 & w5862;
assign w6635 = pi320 & w6437;
assign w6636 = pi148 & pi149;
assign w6637 = ~pi146 & ~pi148;
assign w6638 = ~w5314 & w6637;
assign w6639 = w6431 & ~w6638;
assign w6640 = ~pi149 & ~w6639;
assign w6641 = pi149 & w5857;
assign w6642 = ~w6418 & ~w6641;
assign w6643 = pi145 & ~w6642;
assign w6644 = pi147 & pi149;
assign w6645 = ~w6432 & ~w6644;
assign w6646 = pi146 & ~w6645;
assign w6647 = ~w6643 & ~w6646;
assign w6648 = ~w6640 & w6647;
assign w6649 = ~w6636 & ~w6648;
assign w6650 = pi149 & w6437;
assign w6651 = w6639 & w6650;
assign w6652 = ~w6649 & ~w6651;
assign w6653 = pi321 & w6652;
assign w6654 = ~w6417 & ~w6442;
assign w6655 = ~w6441 & ~w6654;
assign w6656 = ~w6653 & ~w6655;
assign w6657 = w6653 & w6655;
assign w6658 = ~w6656 & ~w6657;
assign w6659 = w6635 & ~w6658;
assign w6660 = ~w6635 & w6658;
assign w6661 = ~w6659 & ~w6660;
assign w6662 = w6634 & ~w6661;
assign w6663 = ~w6634 & w6661;
assign w6664 = ~w6662 & ~w6663;
assign w6665 = pi319 & ~w6448;
assign w6666 = w6664 & w6665;
assign w6667 = ~w6664 & ~w6665;
assign w6668 = w6633 & ~w6666;
assign w6669 = ~w6667 & w6668;
assign w6670 = ~w6447 & ~w6450;
assign w6671 = ~w6664 & ~w6670;
assign w6672 = ~w6662 & w6670;
assign w6673 = ~w6663 & w6672;
assign w6674 = ~w6633 & ~w6671;
assign w6675 = ~w6673 & w6674;
assign w6676 = ~w6669 & ~w6675;
assign w6677 = ~w6458 & ~w6466;
assign w6678 = w6469 & w6677;
assign w6679 = ~w6676 & ~w6678;
assign w6680 = w6676 & w6678;
assign w6681 = ~w6679 & ~w6680;
assign w6682 = w6632 & w6681;
assign w6683 = ~w6632 & ~w6681;
assign w6684 = ~w6682 & ~w6683;
assign w6685 = w5900 & ~w6478;
assign w6686 = w3710 & ~w5901;
assign w6687 = w6472 & ~w6686;
assign w6688 = w4382 & ~w6687;
assign w6689 = ~w6474 & ~w6688;
assign w6690 = pi317 & ~w6689;
assign w6691 = ~w6685 & ~w6690;
assign w6692 = w6684 & ~w6691;
assign w6693 = ~w6684 & w6691;
assign w6694 = ~w6692 & ~w6693;
assign w6695 = ~w6491 & ~w6496;
assign w6696 = ~w6694 & ~w6695;
assign w6697 = w6694 & w6695;
assign w6698 = ~w6696 & ~w6697;
assign w6699 = w6631 & w6698;
assign w6700 = ~w6631 & ~w6698;
assign w6701 = ~w6699 & ~w6700;
assign w6702 = w6630 & w6701;
assign w6703 = ~w6630 & ~w6701;
assign w6704 = ~w6702 & ~w6703;
assign w6705 = ~w6409 & ~w6498;
assign w6706 = w6704 & ~w6705;
assign w6707 = ~w6704 & w6705;
assign w6708 = ~w6706 & ~w6707;
assign w6709 = w6629 & ~w6708;
assign w6710 = ~w6629 & w6708;
assign w6711 = ~w6709 & ~w6710;
assign w6712 = pi313 & w2925;
assign w6713 = w6711 & w6712;
assign w6714 = ~w6711 & ~w6712;
assign w6715 = ~w6713 & ~w6714;
assign w6716 = ~w6510 & ~w6515;
assign w6717 = w6715 & w6716;
assign w6718 = ~w6715 & ~w6716;
assign w6719 = ~w6717 & ~w6718;
assign w6720 = ~w6624 & ~w6719;
assign w6721 = w6624 & w6719;
assign w6722 = ~w6720 & ~w6721;
assign w6723 = w6620 & w6722;
assign w6724 = ~w6620 & ~w6722;
assign w6725 = ~w6723 & ~w6724;
assign w6726 = (~w6526 & ~w6528) | (~w6526 & w16429) | (~w6528 & w16429);
assign w6727 = w6725 & w6726;
assign w6728 = ~w6725 & ~w6726;
assign w6729 = ~w6727 & ~w6728;
assign w6730 = ~w6534 & ~w6729;
assign w6731 = ~w6533 & w6729;
assign w6732 = pi310 & ~w6730;
assign w6733 = ~w6731 & w6732;
assign w6734 = ~w6534 & w6729;
assign w6735 = w1693 & ~w6533;
assign w6736 = w6734 & w6735;
assign w6737 = ~w6733 & ~w6736;
assign w6738 = w1954 & ~w6737;
assign w6739 = ~w6404 & ~w6533;
assign w6740 = pi310 & w1954;
assign w6741 = ~w6729 & ~w6740;
assign w6742 = w6729 & w6740;
assign w6743 = w6739 & ~w6741;
assign w6744 = ~w6742 & w6743;
assign w6745 = (~w6729 & w6739) | (~w6729 & w16430) | (w6739 & w16430);
assign w6746 = ~w1954 & ~w6734;
assign w6747 = ~w6745 & w6746;
assign w6748 = ~w6744 & ~w6747;
assign w6749 = ~w6738 & w6748;
assign w6750 = ~w6619 & w6749;
assign w6751 = w6619 & ~w6749;
assign w6752 = ~w6750 & ~w6751;
assign w6753 = ~w6539 & ~w6543;
assign w6754 = ~w6752 & ~w6753;
assign w6755 = w6752 & w6753;
assign w6756 = ~w6754 & ~w6755;
assign w6757 = w6618 & ~w6756;
assign w6758 = ~w6618 & w6756;
assign w6759 = ~w6757 & ~w6758;
assign w6760 = w6614 & w6759;
assign w6761 = ~w6614 & ~w6759;
assign w6762 = ~w6760 & ~w6761;
assign w6763 = ~w6552 & ~w6555;
assign w6764 = w6762 & ~w6763;
assign w6765 = ~w6762 & w6763;
assign w6766 = ~w6764 & ~w6765;
assign w6767 = ~w6558 & ~w6766;
assign w6768 = w855 & ~w6559;
assign w6769 = w6767 & ~w6768;
assign w6770 = w1159 & ~w6769;
assign w6771 = ~w6559 & w6766;
assign w6772 = pi306 & ~w6771;
assign w6773 = ~w6767 & ~w6772;
assign w6774 = w6770 & ~w6773;
assign w6775 = w6559 & ~w6766;
assign w6776 = ~w6399 & ~w6558;
assign w6777 = w6771 & ~w6776;
assign w6778 = ~w6775 & ~w6777;
assign w6779 = ~w1159 & ~w6778;
assign w6780 = pi306 & w1159;
assign w6781 = ~w6766 & w6780;
assign w6782 = w6766 & ~w6780;
assign w6783 = w6776 & ~w6781;
assign w6784 = ~w6782 & w6783;
assign w6785 = ~w6774 & ~w6784;
assign w6786 = ~w6779 & w6785;
assign w6787 = w6613 & w6786;
assign w6788 = ~w6613 & ~w6786;
assign w6789 = ~w6787 & ~w6788;
assign w6790 = ~w6564 & ~w6567;
assign w6791 = w6789 & ~w6790;
assign w6792 = ~w6789 & w6790;
assign w6793 = ~w6791 & ~w6792;
assign w6794 = w6612 & w6793;
assign w6795 = ~w6612 & ~w6793;
assign w6796 = ~w6794 & ~w6795;
assign w6797 = (~w6579 & ~w6580) | (~w6579 & w16431) | (~w6580 & w16431);
assign w6798 = w6796 & w6797;
assign w6799 = ~w6796 & ~w6797;
assign w6800 = ~w6798 & ~w6799;
assign w6801 = w6607 & ~w6800;
assign w6802 = ~w6607 & w6800;
assign w6803 = ~w6801 & ~w6802;
assign w6804 = w6606 & w6803;
assign w6805 = ~w6606 & ~w6803;
assign w6806 = ~w6804 & ~w6805;
assign w6807 = pi129 & w6806;
assign w6808 = ~pi129 & ~w6806;
assign w6809 = ~w6807 & ~w6808;
assign w6810 = w6601 & ~w6809;
assign w6811 = ~w6601 & w6809;
assign w6812 = ~w6810 & ~w6811;
assign w6813 = w6599 & ~w6812;
assign w6814 = ~w6599 & w6812;
assign w6815 = ~w6813 & ~w6814;
assign w6816 = ~w6387 & ~w6591;
assign w6817 = w6815 & ~w6816;
assign w6818 = ~w6815 & w6816;
assign w6819 = ~w6817 & ~w6818;
assign w6820 = pi343 & w456;
assign w6821 = pi342 & w466;
assign w6822 = ~w6376 & ~w6821;
assign w6823 = w466 & w6376;
assign w6824 = ~w6822 & ~w6823;
assign w6825 = pi341 & ~w537;
assign w6826 = w6825 & w17688;
assign w6827 = (w6372 & w16432) | (w6372 & w16433) | (w16432 & w16433);
assign w6828 = ~w6826 & ~w6827;
assign w6829 = pi340 & ~w615;
assign w6830 = (w6369 & w16434) | (w6369 & w16435) | (w16434 & w16435);
assign w6831 = w537 & ~w6367;
assign w6832 = ~w6368 & w6829;
assign w6833 = ~w6831 & w6832;
assign w6834 = ~w6830 & ~w6833;
assign w6835 = pi339 & ~w793;
assign w6836 = ~w6023 & ~w6364;
assign w6837 = ~w6835 & w6836;
assign w6838 = w6835 & ~w6836;
assign w6839 = ~w6837 & ~w6838;
assign w6840 = w793 & w6026;
assign w6841 = (~w6840 & ~w6360) | (~w6840 & w16436) | (~w6360 & w16436);
assign w6842 = w955 & ~w6841;
assign w6843 = pi338 & ~w6842;
assign w6844 = ~w955 & w6841;
assign w6845 = w6843 & ~w6844;
assign w6846 = pi336 & w1339;
assign w6847 = w6049 & w6354;
assign w6848 = ~w6049 & ~w6354;
assign w6849 = ~w6847 & ~w6848;
assign w6850 = w6045 & w6849;
assign w6851 = ~w6045 & ~w6849;
assign w6852 = ~w6850 & ~w6851;
assign w6853 = w5789 & ~w5792;
assign w6854 = w6039 & ~w6853;
assign w6855 = ~w5796 & w6038;
assign w6856 = (~w6855 & w6852) | (~w6855 & w17594) | (w6852 & w17594);
assign w6857 = ~w6846 & ~w6856;
assign w6858 = w6846 & w6856;
assign w6859 = ~w6857 & ~w6858;
assign w6860 = (~w6847 & ~w6849) | (~w6847 & w17595) | (~w6849 & w17595);
assign w6861 = pi335 & w1602;
assign w6862 = w6860 & ~w6861;
assign w6863 = ~w6860 & w6861;
assign w6864 = ~w6862 & ~w6863;
assign w6865 = pi334 & ~w1865;
assign w6866 = ~w6059 & ~w6353;
assign w6867 = w6067 & ~w6345;
assign w6868 = (~w2170 & ~w6345) | (~w2170 & w15911) | (~w6345 & w15911);
assign w6869 = ~w6867 & ~w6868;
assign w6870 = w2373 & w6869;
assign w6871 = ~w2373 & ~w6869;
assign w6872 = ~w6870 & ~w6871;
assign w6873 = pi332 & w6872;
assign w6874 = pi331 & w2698;
assign w6875 = (~w6063 & ~w6065) | (~w6063 & w15912) | (~w6065 & w15912);
assign w6876 = w6874 & ~w6875;
assign w6877 = ~w6063 & w17689;
assign w6878 = ~w6876 & ~w6877;
assign w6879 = w6873 & w6878;
assign w6880 = ~w6873 & ~w6878;
assign w6881 = ~w6879 & ~w6880;
assign w6882 = pi329 & ~w3568;
assign w6883 = (~w6336 & w6321) | (~w6336 & w17596) | (w6321 & w17596);
assign w6884 = ~w6323 & ~w6883;
assign w6885 = w6882 & w6884;
assign w6886 = ~w6882 & ~w6884;
assign w6887 = ~w6885 & ~w6886;
assign w6888 = pi328 & w3979;
assign w6889 = (~w6076 & ~w6315) | (~w6076 & w16608) | (~w6315 & w16608);
assign w6890 = pi327 & ~w4708;
assign w6891 = pi326 & ~w4854;
assign w6892 = (~w6303 & w6299) | (~w6303 & w15913) | (w6299 & w15913);
assign w6893 = (w6299 & w17597) | (w6299 & w17598) | (w17597 & w17598);
assign w6894 = w6891 & ~w6892;
assign w6895 = ~w6893 & ~w6894;
assign w6896 = ~w6890 & w6895;
assign w6897 = w6890 & ~w6895;
assign w6898 = ~w6896 & ~w6897;
assign w6899 = w6889 & w6898;
assign w6900 = ~w6889 & ~w6898;
assign w6901 = ~w6899 & ~w6900;
assign w6902 = ~w6306 & w6312;
assign w6903 = ~w6313 & ~w6902;
assign w6904 = pi324 & w5714;
assign w6905 = (w6295 & w17599) | (w6295 & w17600) | (w17599 & w17600);
assign w6906 = ~w6904 & w17690;
assign w6907 = ~w6905 & ~w6906;
assign w6908 = pi323 & w6283;
assign w6909 = ~w6087 & w6274;
assign w6910 = w6087 & ~w6274;
assign w6911 = ~w6909 & ~w6910;
assign w6912 = w6272 & w6911;
assign w6913 = ~w6272 & ~w6911;
assign w6914 = ~w6912 & ~w6913;
assign w6915 = w6273 & w6914;
assign w6916 = ~w6273 & ~w6914;
assign w6917 = ~w6915 & ~w6916;
assign w6918 = ~w6090 & ~w6094;
assign w6919 = w6917 & ~w6918;
assign w6920 = w6090 & ~w6093;
assign w6921 = ~w6917 & ~w6920;
assign w6922 = ~w6919 & ~w6921;
assign w6923 = pi146 & pi261;
assign w6924 = (~w6258 & ~w6260) | (~w6258 & w16187) | (~w6260 & w16187);
assign w6925 = pi143 & pi264;
assign w6926 = (~w6242 & ~w6238) | (~w6242 & w15915) | (~w6238 & w15915);
assign w6927 = ~w6240 & ~w6926;
assign w6928 = pi140 & pi267;
assign w6929 = pi137 & pi270;
assign w6930 = pi134 & pi273;
assign w6931 = pi133 & pi274;
assign w6932 = pi132 & pi275;
assign w6933 = pi131 & pi276;
assign w6934 = ~w6146 & ~w6153;
assign w6935 = pi129 & pi278;
assign w6936 = pi128 & pi279;
assign w6937 = ~w6935 & ~w6936;
assign w6938 = w6935 & w6936;
assign w6939 = ~w6937 & ~w6938;
assign w6940 = w6131 & ~w6133;
assign w6941 = ~w6135 & ~w6940;
assign w6942 = w6135 & w6940;
assign w6943 = (~w6136 & ~w6940) | (~w6136 & w16437) | (~w6940 & w16437);
assign w6944 = ~w6941 & ~w6943;
assign w6945 = w6939 & ~w6944;
assign w6946 = pi129 & ~w6939;
assign w6947 = ~w6941 & w6946;
assign w6948 = ~w6945 & ~w6947;
assign w6949 = ~pi130 & w6948;
assign w6950 = ~w6939 & w6942;
assign w6951 = ~pi277 & ~w6950;
assign w6952 = ~w6945 & w6951;
assign w6953 = ~w6949 & ~w6952;
assign w6954 = pi130 & pi277;
assign w6955 = ~w6948 & w6954;
assign w6956 = w6953 & ~w6955;
assign w6957 = w6934 & ~w6956;
assign w6958 = ~w6934 & w6956;
assign w6959 = ~w6957 & ~w6958;
assign w6960 = w6933 & ~w6959;
assign w6961 = ~w6933 & w6959;
assign w6962 = ~w6960 & ~w6961;
assign w6963 = ~w6155 & ~w6159;
assign w6964 = w6962 & ~w6963;
assign w6965 = ~w6962 & w6963;
assign w6966 = ~w6964 & ~w6965;
assign w6967 = w6932 & ~w6966;
assign w6968 = ~w6932 & w6966;
assign w6969 = ~w6967 & ~w6968;
assign w6970 = ~w6163 & ~w6167;
assign w6971 = ~w6969 & w6970;
assign w6972 = w6969 & ~w6970;
assign w6973 = ~w6971 & ~w6972;
assign w6974 = (~w6169 & w6173) | (~w6169 & w15917) | (w6173 & w15917);
assign w6975 = w6973 & ~w6974;
assign w6976 = ~w6973 & w6974;
assign w6977 = ~w6975 & ~w6976;
assign w6978 = w6931 & ~w6977;
assign w6979 = ~w6931 & w6977;
assign w6980 = ~w6978 & ~w6979;
assign w6981 = ~w6930 & w6980;
assign w6982 = w6930 & ~w6980;
assign w6983 = ~w6981 & ~w6982;
assign w6984 = (~w6177 & ~w6179) | (~w6177 & w16438) | (~w6179 & w16438);
assign w6985 = w6983 & ~w6984;
assign w6986 = ~w6983 & w6984;
assign w6987 = ~w6985 & ~w6986;
assign w6988 = (~w6183 & w6187) | (~w6183 & w16188) | (w6187 & w16188);
assign w6989 = w6987 & w6988;
assign w6990 = ~w6987 & ~w6988;
assign w6991 = ~w6989 & ~w6990;
assign w6992 = pi136 & pi271;
assign w6993 = pi135 & pi272;
assign w6994 = w6992 & ~w6993;
assign w6995 = ~w6992 & w6993;
assign w6996 = ~w6994 & ~w6995;
assign w6997 = w6991 & w6996;
assign w6998 = ~w6991 & ~w6996;
assign w6999 = ~w6997 & ~w6998;
assign w7000 = ~w6192 & w6196;
assign w7001 = ~w6191 & ~w7000;
assign w7002 = ~w6999 & w7001;
assign w7003 = w6999 & ~w7001;
assign w7004 = ~w7002 & ~w7003;
assign w7005 = ~w6929 & w7004;
assign w7006 = w6929 & ~w7004;
assign w7007 = ~w7005 & ~w7006;
assign w7008 = ~w6194 & ~w6202;
assign w7009 = ~w6204 & ~w7008;
assign w7010 = w7007 & w7009;
assign w7011 = ~w7007 & ~w7009;
assign w7012 = ~w7010 & ~w7011;
assign w7013 = (~w7012 & w6211) | (~w7012 & w15918) | (w6211 & w15918);
assign w7014 = ~w6211 & w15919;
assign w7015 = ~w7013 & ~w7014;
assign w7016 = pi139 & pi268;
assign w7017 = pi138 & pi269;
assign w7018 = w7016 & ~w7017;
assign w7019 = ~w7016 & w7017;
assign w7020 = ~w7018 & ~w7019;
assign w7021 = w7015 & w7020;
assign w7022 = ~w7015 & ~w7020;
assign w7023 = ~w7021 & ~w7022;
assign w7024 = ~w6215 & w6219;
assign w7025 = ~w6214 & ~w7024;
assign w7026 = w7023 & w7025;
assign w7027 = ~w7023 & ~w7025;
assign w7028 = ~w7026 & ~w7027;
assign w7029 = ~w6928 & w7028;
assign w7030 = w6928 & ~w7028;
assign w7031 = ~w7029 & ~w7030;
assign w7032 = w6217 & w6225;
assign w7033 = ~w6226 & ~w7032;
assign w7034 = w7031 & ~w7033;
assign w7035 = ~w7031 & w7033;
assign w7036 = ~w7034 & ~w7035;
assign w7037 = (w15916 & w16439) | (w15916 & w16440) | (w16439 & w16440);
assign w7038 = (~w15916 & w16441) | (~w15916 & w16442) | (w16441 & w16442);
assign w7039 = ~w7037 & ~w7038;
assign w7040 = pi142 & pi265;
assign w7041 = pi141 & pi266;
assign w7042 = w7040 & ~w7041;
assign w7043 = ~w7040 & w7041;
assign w7044 = ~w7042 & ~w7043;
assign w7045 = w7039 & w7044;
assign w7046 = ~w7039 & ~w7044;
assign w7047 = ~w7045 & ~w7046;
assign w7048 = w6927 & ~w7047;
assign w7049 = ~w6927 & w7047;
assign w7050 = ~w7048 & ~w7049;
assign w7051 = w6925 & w7050;
assign w7052 = ~w6925 & ~w7050;
assign w7053 = ~w7051 & ~w7052;
assign w7054 = w6113 & ~w6249;
assign w7055 = w6243 & w6249;
assign w7056 = ~w7054 & ~w7055;
assign w7057 = w7053 & ~w7056;
assign w7058 = ~w7053 & w7056;
assign w7059 = ~w7057 & ~w7058;
assign w7060 = w6112 & ~w6252;
assign w7061 = ~w6255 & ~w7060;
assign w7062 = ~w7059 & w7061;
assign w7063 = w7059 & ~w7061;
assign w7064 = ~w7062 & ~w7063;
assign w7065 = pi145 & pi262;
assign w7066 = pi144 & pi263;
assign w7067 = w7065 & ~w7066;
assign w7068 = ~w7065 & w7066;
assign w7069 = ~w7067 & ~w7068;
assign w7070 = w7064 & w7069;
assign w7071 = ~w7064 & ~w7069;
assign w7072 = ~w7070 & ~w7071;
assign w7073 = ~w6924 & ~w7072;
assign w7074 = w6924 & w7072;
assign w7075 = ~w7073 & ~w7074;
assign w7076 = ~w6923 & ~w7075;
assign w7077 = w6923 & w7075;
assign w7078 = ~w7076 & ~w7077;
assign w7079 = w6099 & w6106;
assign w7080 = ~w6271 & ~w7079;
assign w7081 = w7078 & ~w7080;
assign w7082 = ~w7078 & w7080;
assign w7083 = ~w7081 & ~w7082;
assign w7084 = ~w6909 & ~w6912;
assign w7085 = w7083 & ~w7084;
assign w7086 = ~w7083 & w7084;
assign w7087 = ~w7085 & ~w7086;
assign w7088 = pi148 & pi259;
assign w7089 = (~w7088 & ~w6914) | (~w7088 & w15920) | (~w6914 & w15920);
assign w7090 = pi147 & w6087;
assign w7091 = ~w6272 & ~w7090;
assign w7092 = pi148 & w458;
assign w7093 = (w7092 & ~w6272) | (w7092 & w16189) | (~w6272 & w16189);
assign w7094 = ~w7091 & w7093;
assign w7095 = pi149 & pi258;
assign w7096 = pi147 & pi260;
assign w7097 = w7095 & ~w7096;
assign w7098 = ~w7095 & w7096;
assign w7099 = ~w7097 & ~w7098;
assign w7100 = ~w7089 & w16190;
assign w7101 = (w7099 & w7089) | (w7099 & w16191) | (w7089 & w16191);
assign w7102 = ~w7100 & ~w7101;
assign w7103 = w7087 & w7102;
assign w7104 = ~w7087 & ~w7102;
assign w7105 = ~w7103 & ~w7104;
assign w7106 = w6922 & ~w7105;
assign w7107 = ~w6922 & w7105;
assign w7108 = ~w7106 & ~w7107;
assign w7109 = (~w6908 & w7108) | (~w6908 & w16192) | (w7108 & w16192);
assign w7110 = ~w7108 & w16193;
assign w7111 = ~w7109 & ~w7110;
assign w7112 = w6907 & w7111;
assign w7113 = ~w6907 & ~w7111;
assign w7114 = ~w7112 & ~w7113;
assign w7115 = pi325 & w5194;
assign w7116 = ~w6287 & ~w6290;
assign w7117 = w7115 & ~w7116;
assign w7118 = ~w7115 & w7116;
assign w7119 = ~w7117 & ~w7118;
assign w7120 = w7114 & w7119;
assign w7121 = ~w7114 & ~w7119;
assign w7122 = ~w7120 & ~w7121;
assign w7123 = ~w6903 & w7122;
assign w7124 = w6903 & ~w7122;
assign w7125 = ~w7123 & ~w7124;
assign w7126 = w6901 & w7125;
assign w7127 = ~w6901 & ~w7125;
assign w7128 = ~w7126 & ~w7127;
assign w7129 = ~w6888 & w7128;
assign w7130 = w6888 & ~w7128;
assign w7131 = ~w7129 & ~w7130;
assign w7132 = ~w6072 & ~w6319;
assign w7133 = w7131 & ~w7132;
assign w7134 = ~w7131 & w7132;
assign w7135 = ~w7133 & ~w7134;
assign w7136 = w6887 & ~w7135;
assign w7137 = ~w6887 & w7135;
assign w7138 = ~w7136 & ~w7137;
assign w7139 = pi330 & ~w3183;
assign w7140 = ~pi329 & w7139;
assign w7141 = ~w6328 & w7140;
assign w7142 = ~w6325 & w7141;
assign w7143 = w6331 & ~w7140;
assign w7144 = ~w6328 & ~w7139;
assign w7145 = ~w3183 & ~w6329;
assign w7146 = ~w7144 & ~w7145;
assign w7147 = ~w7142 & ~w7146;
assign w7148 = ~w7143 & w7147;
assign w7149 = w7138 & w7148;
assign w7150 = ~w7138 & ~w7148;
assign w7151 = ~w7149 & ~w7150;
assign w7152 = w6334 & ~w6335;
assign w7153 = ~w6334 & w6335;
assign w7154 = w6333 & w6336;
assign w7155 = ~w6333 & ~w6336;
assign w7156 = ~w7154 & ~w7155;
assign w7157 = ~w7153 & ~w7156;
assign w7158 = ~w7152 & ~w7157;
assign w7159 = w7151 & ~w7158;
assign w7160 = ~w7151 & w7158;
assign w7161 = ~w7159 & ~w7160;
assign w7162 = pi333 & ~w2170;
assign w7163 = w7161 & ~w7162;
assign w7164 = ~w7161 & w7162;
assign w7165 = ~w7163 & ~w7164;
assign w7166 = w6881 & w7165;
assign w7167 = ~w6881 & ~w7165;
assign w7168 = ~w7166 & ~w7167;
assign w7169 = ~w6866 & ~w7168;
assign w7170 = w6866 & w7168;
assign w7171 = ~w7169 & ~w7170;
assign w7172 = w6865 & w7171;
assign w7173 = ~w6865 & ~w7171;
assign w7174 = ~w7172 & ~w7173;
assign w7175 = w6864 & w7174;
assign w7176 = ~w6864 & ~w7174;
assign w7177 = ~w7175 & ~w7176;
assign w7178 = ~w6859 & ~w7177;
assign w7179 = w6859 & w7177;
assign w7180 = ~w7178 & ~w7179;
assign w7181 = pi337 & w1101;
assign w7182 = ~w6050 & w6057;
assign w7183 = w6050 & ~w6057;
assign w7184 = ~w6048 & ~w6849;
assign w7185 = (~w7183 & ~w6048) | (~w7183 & w15921) | (~w6048 & w15921);
assign w7186 = ~w7184 & w7185;
assign w7187 = ~w7182 & ~w7186;
assign w7188 = (w7181 & w7186) | (w7181 & w16443) | (w7186 & w16443);
assign w7189 = ~w7186 & w16444;
assign w7190 = ~w7188 & ~w7189;
assign w7191 = w7180 & w7190;
assign w7192 = ~w7180 & ~w7190;
assign w7193 = ~w7191 & ~w7192;
assign w7194 = w6845 & w7193;
assign w7195 = ~w6845 & ~w7193;
assign w7196 = ~w7194 & ~w7195;
assign w7197 = w6839 & ~w7196;
assign w7198 = ~w6839 & w7196;
assign w7199 = ~w7197 & ~w7198;
assign w7200 = ~w6834 & w7199;
assign w7201 = w6834 & ~w7199;
assign w7202 = ~w7200 & ~w7201;
assign w7203 = w6828 & w7202;
assign w7204 = ~w6828 & ~w7202;
assign w7205 = ~w7203 & ~w7204;
assign w7206 = w6824 & w7205;
assign w7207 = ~w6824 & ~w7205;
assign w7208 = ~w7206 & ~w7207;
assign w7209 = w6820 & w7208;
assign w7210 = ~w6820 & ~w7208;
assign w7211 = ~w7209 & ~w7210;
assign w7212 = ~w6380 & ~w6383;
assign w7213 = pi279 & ~w7212;
assign w7214 = ~pi279 & w7212;
assign w7215 = ~w7213 & ~w7214;
assign w7216 = w7211 & ~w7215;
assign w7217 = ~w7211 & w7215;
assign w7218 = ~w7216 & ~w7217;
assign w7219 = ~w6819 & ~w7218;
assign w7220 = w6819 & w7218;
assign w7221 = ~w135 & ~w7219;
assign w7222 = ~w7220 & w7221;
assign w7223 = pi161 & ~w182;
assign w7224 = ~w7222 & w7223;
assign w7225 = ~pi160 & ~w6598;
assign w7226 = ~w7224 & w7225;
assign w7227 = ~pi086 & ~pi161;
assign w7228 = pi128 & pi299;
assign w7229 = pi300 & w464;
assign w7230 = ~w6813 & ~w7229;
assign w7231 = ~pi129 & w6813;
assign w7232 = ~w7230 & ~w7231;
assign w7233 = pi302 & w709;
assign w7234 = pi304 & w855;
assign w7235 = pi306 & w1220;
assign w7236 = pi307 & w1420;
assign w7237 = pi308 & w1693;
assign w7238 = pi309 & w1954;
assign w7239 = ~w6750 & ~w6755;
assign w7240 = ~w7238 & ~w7239;
assign w7241 = w7238 & w7239;
assign w7242 = ~w7240 & ~w7241;
assign w7243 = pi310 & ~w2473;
assign w7244 = pi311 & w2801;
assign w7245 = pi312 & w2925;
assign w7246 = pi314 & w3710;
assign w7247 = pi315 & w4382;
assign w7248 = ~w6703 & ~w6706;
assign w7249 = ~w7247 & ~w7248;
assign w7250 = w7247 & w7248;
assign w7251 = ~w7249 & ~w7250;
assign w7252 = pi316 & w4539;
assign w7253 = pi317 & w5316;
assign w7254 = ~w6682 & ~w6692;
assign w7255 = w7253 & ~w7254;
assign w7256 = ~w7253 & w7254;
assign w7257 = ~w7255 & ~w7256;
assign w7258 = pi318 & w5862;
assign w7259 = pi319 & w6437;
assign w7260 = pi320 & w6652;
assign w7261 = ~w6425 & ~w6636;
assign w7262 = w6647 & w7261;
assign w7263 = ~pi150 & w7262;
assign w7264 = pi150 & ~w7262;
assign w7265 = ~w7263 & ~w7264;
assign w7266 = pi149 & w7265;
assign w7267 = ~pi149 & ~w7265;
assign w7268 = ~w7266 & ~w7267;
assign w7269 = pi321 & w7268;
assign w7270 = ~w6635 & ~w6657;
assign w7271 = ~w6656 & ~w7270;
assign w7272 = ~w7269 & ~w7271;
assign w7273 = w7269 & w7271;
assign w7274 = ~w7272 & ~w7273;
assign w7275 = w7260 & ~w7274;
assign w7276 = ~w7260 & w7274;
assign w7277 = ~w7275 & ~w7276;
assign w7278 = w7259 & ~w7277;
assign w7279 = ~w7259 & w7277;
assign w7280 = ~w7278 & ~w7279;
assign w7281 = ~w6663 & ~w6672;
assign w7282 = w7280 & w7281;
assign w7283 = ~w7280 & ~w7281;
assign w7284 = ~w7282 & ~w7283;
assign w7285 = ~w7258 & ~w7284;
assign w7286 = w7258 & w7284;
assign w7287 = ~w7285 & ~w7286;
assign w7288 = ~w6669 & ~w6680;
assign w7289 = w7287 & ~w7288;
assign w7290 = ~w7287 & w7288;
assign w7291 = ~w7289 & ~w7290;
assign w7292 = w7257 & w7291;
assign w7293 = ~w7257 & ~w7291;
assign w7294 = ~w7292 & ~w7293;
assign w7295 = ~w6697 & ~w7294;
assign w7296 = ~w6699 & w7295;
assign w7297 = w6697 & w7294;
assign w7298 = ~w7296 & ~w7297;
assign w7299 = w7252 & ~w7298;
assign w7300 = w6454 & w6698;
assign w7301 = ~w6631 & ~w7252;
assign w7302 = ~w6697 & w7301;
assign w7303 = ~w7300 & ~w7302;
assign w7304 = w7294 & ~w7303;
assign w7305 = ~w4539 & ~w7294;
assign w7306 = ~w6696 & ~w7305;
assign w7307 = ~w4539 & ~w7306;
assign w7308 = ~w7296 & w7307;
assign w7309 = ~w7304 & ~w7308;
assign w7310 = ~w7299 & w7309;
assign w7311 = ~w7251 & w7310;
assign w7312 = w7251 & ~w7310;
assign w7313 = ~w7311 & ~w7312;
assign w7314 = w7246 & w7313;
assign w7315 = ~w7246 & ~w7313;
assign w7316 = ~w7314 & ~w7315;
assign w7317 = ~w6627 & ~w6709;
assign w7318 = w7316 & ~w7317;
assign w7319 = ~w7316 & w7317;
assign w7320 = ~w7318 & ~w7319;
assign w7321 = pi313 & w3304;
assign w7322 = ~w2925 & ~w6711;
assign w7323 = w6716 & ~w7322;
assign w7324 = ~w6713 & ~w7323;
assign w7325 = w7321 & ~w7324;
assign w7326 = ~w7321 & w7324;
assign w7327 = ~w7325 & ~w7326;
assign w7328 = w7320 & w7327;
assign w7329 = ~w7320 & ~w7327;
assign w7330 = ~w7328 & ~w7329;
assign w7331 = ~w7245 & ~w7330;
assign w7332 = w7245 & w7330;
assign w7333 = ~w7331 & ~w7332;
assign w7334 = ~w6623 & ~w6721;
assign w7335 = ~w7333 & ~w7334;
assign w7336 = w7333 & w7334;
assign w7337 = ~w7335 & ~w7336;
assign w7338 = ~w6723 & ~w6727;
assign w7339 = w7337 & w7338;
assign w7340 = ~w7337 & ~w7338;
assign w7341 = ~w7339 & ~w7340;
assign w7342 = w7244 & w7341;
assign w7343 = ~w7244 & ~w7341;
assign w7344 = ~w7342 & ~w7343;
assign w7345 = ~w6745 & w6748;
assign w7346 = w7344 & w7345;
assign w7347 = ~w7344 & ~w7345;
assign w7348 = ~w7346 & ~w7347;
assign w7349 = w7243 & ~w7348;
assign w7350 = ~w7243 & w7348;
assign w7351 = ~w7349 & ~w7350;
assign w7352 = w7242 & w7351;
assign w7353 = ~w7242 & ~w7351;
assign w7354 = ~w7352 & ~w7353;
assign w7355 = w7237 & ~w7354;
assign w7356 = ~w7237 & w7354;
assign w7357 = ~w7355 & ~w7356;
assign w7358 = ~w6617 & ~w6757;
assign w7359 = w7357 & ~w7358;
assign w7360 = ~w7357 & w7358;
assign w7361 = ~w7359 & ~w7360;
assign w7362 = ~w6760 & ~w6764;
assign w7363 = w7361 & ~w7362;
assign w7364 = ~w7361 & w7362;
assign w7365 = ~w7363 & ~w7364;
assign w7366 = w7236 & ~w7365;
assign w7367 = ~w7236 & w7365;
assign w7368 = ~w7366 & ~w7367;
assign w7369 = w7235 & ~w7368;
assign w7370 = ~w7235 & w7368;
assign w7371 = ~w7369 & ~w7370;
assign w7372 = pi306 & w6770;
assign w7373 = ~w6777 & ~w7372;
assign w7374 = ~w7371 & w7373;
assign w7375 = w7371 & ~w7373;
assign w7376 = ~w7374 & ~w7375;
assign w7377 = pi305 & w1159;
assign w7378 = ~w6787 & ~w6791;
assign w7379 = w7377 & ~w7378;
assign w7380 = ~w7377 & w7378;
assign w7381 = ~w7379 & ~w7380;
assign w7382 = w7376 & w7381;
assign w7383 = ~w7376 & ~w7381;
assign w7384 = ~w7382 & ~w7383;
assign w7385 = w7234 & w7384;
assign w7386 = ~w7234 & ~w7384;
assign w7387 = ~w7385 & ~w7386;
assign w7388 = ~w6610 & ~w6794;
assign w7389 = w7387 & ~w7388;
assign w7390 = ~w7387 & w7388;
assign w7391 = ~w7389 & ~w7390;
assign w7392 = ~w6607 & ~w6798;
assign w7393 = ~w6799 & ~w7392;
assign w7394 = ~w7391 & ~w7393;
assign w7395 = w7391 & w7393;
assign w7396 = ~w7394 & ~w7395;
assign w7397 = pi303 & w698;
assign w7398 = w7396 & w7397;
assign w7399 = ~w7396 & ~w7397;
assign w7400 = ~w7398 & ~w7399;
assign w7401 = w7233 & w7400;
assign w7402 = ~w7233 & ~w7400;
assign w7403 = ~w7401 & ~w7402;
assign w7404 = ~w6604 & ~w6804;
assign w7405 = w7403 & w7404;
assign w7406 = ~w7403 & ~w7404;
assign w7407 = ~w7405 & ~w7406;
assign w7408 = ~w651 & ~w5426;
assign w7409 = ~w6809 & ~w7408;
assign w7410 = w6390 & w6586;
assign w7411 = ~w463 & ~w6809;
assign w7412 = pi130 & ~w7410;
assign w7413 = ~w7411 & w7412;
assign w7414 = ~w7409 & ~w7413;
assign w7415 = pi301 & ~w7414;
assign w7416 = ~w6807 & w7410;
assign w7417 = w653 & w7416;
assign w7418 = ~w7415 & ~w7417;
assign w7419 = w7407 & ~w7418;
assign w7420 = ~w7407 & w7418;
assign w7421 = ~w7419 & ~w7420;
assign w7422 = w7232 & w7421;
assign w7423 = ~w7232 & ~w7421;
assign w7424 = ~w7422 & ~w7423;
assign w7425 = w7228 & w7424;
assign w7426 = ~w7228 & ~w7424;
assign w7427 = ~w7425 & ~w7426;
assign w7428 = ~w6818 & ~w7220;
assign w7429 = w7427 & w7428;
assign w7430 = ~w7427 & ~w7428;
assign w7431 = ~w7429 & ~w7430;
assign w7432 = ~w7213 & ~w7217;
assign w7433 = pi344 & w456;
assign w7434 = pi343 & w466;
assign w7435 = ~w7209 & ~w7434;
assign w7436 = w466 & w7209;
assign w7437 = ~w7435 & ~w7436;
assign w7438 = pi342 & ~w537;
assign w7439 = pi341 & ~w615;
assign w7440 = ~w6826 & ~w7203;
assign w7441 = ~w7439 & w7440;
assign w7442 = w7439 & ~w7440;
assign w7443 = ~w7441 & ~w7442;
assign w7444 = ~w6837 & ~w7197;
assign w7445 = pi338 & w1101;
assign w7446 = w6842 & w7445;
assign w7447 = ~pi337 & w7445;
assign w7448 = ~w6844 & w7445;
assign w7449 = w6843 & ~w7181;
assign w7450 = ~w7448 & ~w7449;
assign w7451 = w7180 & ~w7187;
assign w7452 = ~w7180 & w7187;
assign w7453 = ~w7451 & ~w7452;
assign w7454 = ~w7447 & w7453;
assign w7455 = ~w7450 & w7454;
assign w7456 = ~pi337 & w7448;
assign w7457 = ~w7453 & w7456;
assign w7458 = pi338 & ~w1101;
assign w7459 = w6844 & w7458;
assign w7460 = ~w7446 & ~w7459;
assign w7461 = ~w7457 & w7460;
assign w7462 = ~w7455 & w7461;
assign w7463 = pi339 & ~w955;
assign w7464 = pi337 & w1339;
assign w7465 = (w7180 & w17601) | (w7180 & w17602) | (w17601 & w17602);
assign w7466 = ~w7464 & w17691;
assign w7467 = ~w7465 & ~w7466;
assign w7468 = pi335 & ~w1865;
assign w7469 = ~w7468 & w17692;
assign w7470 = (w7174 & w17603) | (w7174 & w17604) | (w17603 & w17604);
assign w7471 = ~w7469 & ~w7470;
assign w7472 = pi334 & ~w2170;
assign w7473 = ~w7169 & ~w7472;
assign w7474 = ~w7172 & w7473;
assign w7475 = w1865 & ~w7169;
assign w7476 = ~w7170 & w7472;
assign w7477 = ~w7475 & w7476;
assign w7478 = ~w7474 & ~w7477;
assign w7479 = pi333 & ~w2373;
assign w7480 = pi332 & w2698;
assign w7481 = (w7480 & w6869) | (w7480 & w16447) | (w6869 & w16447);
assign w7482 = ~pi331 & w7481;
assign w7483 = ~w7161 & w7482;
assign w7484 = ~pi332 & w6867;
assign w7485 = ~w6872 & ~w7484;
assign w7486 = pi332 & ~w2698;
assign w7487 = (w7486 & ~w6869) | (w7486 & w17605) | (~w6869 & w17605);
assign w7488 = ~w7481 & ~w7487;
assign w7489 = (~w15922 & w16609) | (~w15922 & w16610) | (w16609 & w16610);
assign w7490 = ~w7483 & ~w7489;
assign w7491 = pi331 & ~w3183;
assign w7492 = (~w6329 & ~w7156) | (~w6329 & w15923) | (~w7156 & w15923);
assign w7493 = (~w3183 & w7138) | (~w3183 & w15924) | (w7138 & w15924);
assign w7494 = w7138 & w7492;
assign w7495 = (~w3568 & ~w7138) | (~w3568 & w15925) | (~w7138 & w15925);
assign w7496 = ~w7493 & w7495;
assign w7497 = ~w3183 & w3568;
assign w7498 = (w7497 & w7138) | (w7497 & w16448) | (w7138 & w16448);
assign w7499 = pi330 & ~w3568;
assign w7500 = w7494 & ~w7499;
assign w7501 = ~w7500 & w17693;
assign w7502 = ~w7491 & w7501;
assign w7503 = w7491 & ~w7501;
assign w7504 = ~w7502 & ~w7503;
assign w7505 = w7490 & ~w7504;
assign w7506 = ~w7490 & w7504;
assign w7507 = ~w7505 & ~w7506;
assign w7508 = w7479 & w7507;
assign w7509 = ~w7479 & ~w7507;
assign w7510 = ~w7508 & ~w7509;
assign w7511 = w6875 & ~w7162;
assign w7512 = ~w6875 & w7162;
assign w7513 = w6874 & w7161;
assign w7514 = ~w6874 & ~w7161;
assign w7515 = ~w7513 & ~w7514;
assign w7516 = ~w6873 & ~w7515;
assign w7517 = w6873 & w7515;
assign w7518 = ~w7516 & ~w7517;
assign w7519 = (~w7511 & w7518) | (~w7511 & w15926) | (w7518 & w15926);
assign w7520 = pi328 & ~w4708;
assign w7521 = ~w7129 & ~w7133;
assign w7522 = w7520 & w7521;
assign w7523 = ~w7520 & ~w7521;
assign w7524 = ~w7522 & ~w7523;
assign w7525 = pi326 & w5194;
assign w7526 = pi327 & ~w4854;
assign w7527 = w7525 & ~w7526;
assign w7528 = ~w7525 & w7526;
assign w7529 = ~w7527 & ~w7528;
assign w7530 = ~w6889 & ~w6890;
assign w7531 = w6889 & w6890;
assign w7532 = ~w6895 & w7125;
assign w7533 = w6895 & ~w7125;
assign w7534 = ~w7531 & ~w7532;
assign w7535 = ~w7533 & w7534;
assign w7536 = ~w7530 & ~w7535;
assign w7537 = w7529 & w7536;
assign w7538 = ~w7529 & ~w7536;
assign w7539 = ~w7537 & ~w7538;
assign w7540 = pi325 & w5714;
assign w7541 = pi324 & w6283;
assign w7542 = ~w7111 & ~w7116;
assign w7543 = w7111 & w7116;
assign w7544 = ~w6905 & ~w7542;
assign w7545 = ~w7543 & w7544;
assign w7546 = ~w6906 & ~w7545;
assign w7547 = ~w7541 & ~w7546;
assign w7548 = w7541 & w7546;
assign w7549 = ~w7547 & ~w7548;
assign w7550 = pi323 & ~w7108;
assign w7551 = ~w6919 & ~w7105;
assign w7552 = ~w6921 & w7105;
assign w7553 = ~w7551 & ~w7552;
assign w7554 = ~w7094 & w7096;
assign w7555 = ~w7094 & ~w7096;
assign w7556 = ~w7087 & w7555;
assign w7557 = (~w7089 & ~w7087) | (~w7089 & w15927) | (~w7087 & w15927);
assign w7558 = ~w7556 & w7557;
assign w7559 = pi147 & pi261;
assign w7560 = (~w7077 & ~w7078) | (~w7077 & w15928) | (~w7078 & w15928);
assign w7561 = pi145 & pi263;
assign w7562 = pi144 & pi264;
assign w7563 = (~w7051 & ~w7053) | (~w7051 & w16611) | (~w7053 & w16611);
assign w7564 = pi141 & pi267;
assign w7565 = ~w7030 & ~w7034;
assign w7566 = pi139 & pi269;
assign w7567 = pi138 & pi270;
assign w7568 = ~w7006 & ~w7010;
assign w7569 = pi135 & pi273;
assign w7570 = (~w6982 & ~w6983) | (~w6982 & w16450) | (~w6983 & w16450);
assign w7571 = pi134 & pi274;
assign w7572 = pi133 & pi275;
assign w7573 = pi132 & pi276;
assign w7574 = pi131 & pi277;
assign w7575 = pi130 & pi278;
assign w7576 = pi128 & pi280;
assign w7577 = pi129 & pi279;
assign w7578 = ~w6937 & w6944;
assign w7579 = ~w7577 & ~w7578;
assign w7580 = ~w6135 & ~w7578;
assign w7581 = w7577 & ~w7580;
assign w7582 = ~w7579 & ~w7581;
assign w7583 = w7576 & ~w7582;
assign w7584 = ~w7576 & w7582;
assign w7585 = ~w7583 & ~w7584;
assign w7586 = w7575 & ~w7585;
assign w7587 = ~w7575 & w7585;
assign w7588 = ~w7586 & ~w7587;
assign w7589 = w6953 & ~w6958;
assign w7590 = w7588 & ~w7589;
assign w7591 = ~w7588 & w7589;
assign w7592 = ~w7590 & ~w7591;
assign w7593 = w7574 & ~w7592;
assign w7594 = ~w7574 & w7592;
assign w7595 = ~w7593 & ~w7594;
assign w7596 = ~w6961 & ~w6964;
assign w7597 = w7595 & w7596;
assign w7598 = ~w7595 & ~w7596;
assign w7599 = ~w7597 & ~w7598;
assign w7600 = w7573 & w7599;
assign w7601 = ~w7573 & ~w7599;
assign w7602 = ~w7600 & ~w7601;
assign w7603 = ~w6967 & ~w6972;
assign w7604 = w7602 & w7603;
assign w7605 = ~w7602 & ~w7603;
assign w7606 = ~w7604 & ~w7605;
assign w7607 = w7572 & ~w7606;
assign w7608 = ~w7572 & w7606;
assign w7609 = ~w7607 & ~w7608;
assign w7610 = (~w6976 & ~w6977) | (~w6976 & w16451) | (~w6977 & w16451);
assign w7611 = ~w7609 & ~w7610;
assign w7612 = w7609 & w7610;
assign w7613 = ~w7611 & ~w7612;
assign w7614 = w7571 & w7613;
assign w7615 = ~w7571 & ~w7613;
assign w7616 = ~w7614 & ~w7615;
assign w7617 = w7570 & w7616;
assign w7618 = ~w7570 & ~w7616;
assign w7619 = ~w7617 & ~w7618;
assign w7620 = w7569 & ~w7619;
assign w7621 = ~w7569 & w7619;
assign w7622 = ~w7620 & ~w7621;
assign w7623 = (~w6993 & ~w6988) | (~w6993 & w16452) | (~w6988 & w16452);
assign w7624 = ~w6990 & ~w7623;
assign w7625 = ~w7622 & w7624;
assign w7626 = w7622 & ~w7624;
assign w7627 = ~w7625 & ~w7626;
assign w7628 = ~w6992 & w6999;
assign w7629 = ~w7002 & ~w7628;
assign w7630 = w7627 & ~w7629;
assign w7631 = ~w7627 & w7629;
assign w7632 = ~w7630 & ~w7631;
assign w7633 = pi137 & pi271;
assign w7634 = pi136 & pi272;
assign w7635 = w7633 & ~w7634;
assign w7636 = ~w7633 & w7634;
assign w7637 = ~w7635 & ~w7636;
assign w7638 = w7632 & w7637;
assign w7639 = ~w7632 & ~w7637;
assign w7640 = ~w7638 & ~w7639;
assign w7641 = w7568 & ~w7640;
assign w7642 = ~w7568 & w7640;
assign w7643 = ~w7641 & ~w7642;
assign w7644 = w7567 & ~w7643;
assign w7645 = ~w7567 & w7643;
assign w7646 = ~w7644 & ~w7645;
assign w7647 = ~w7014 & ~w7017;
assign w7648 = ~w7013 & ~w7647;
assign w7649 = w7646 & w7648;
assign w7650 = ~w7646 & ~w7648;
assign w7651 = ~w7649 & ~w7650;
assign w7652 = ~w7566 & ~w7651;
assign w7653 = w7566 & w7651;
assign w7654 = ~w7652 & ~w7653;
assign w7655 = pi140 & pi268;
assign w7656 = ~w7016 & w7023;
assign w7657 = ~w7027 & ~w7656;
assign w7658 = w7655 & ~w7657;
assign w7659 = ~w7655 & w7657;
assign w7660 = ~w7658 & ~w7659;
assign w7661 = w7654 & w7660;
assign w7662 = ~w7654 & ~w7660;
assign w7663 = ~w7661 & ~w7662;
assign w7664 = w7565 & ~w7663;
assign w7665 = ~w7565 & w7663;
assign w7666 = ~w7664 & ~w7665;
assign w7667 = w7564 & ~w7666;
assign w7668 = ~w7564 & w7666;
assign w7669 = ~w7667 & ~w7668;
assign w7670 = (w15916 & w17606) | (w15916 & w17607) | (w17606 & w17607);
assign w7671 = ~w7037 & ~w7670;
assign w7672 = w7669 & w7671;
assign w7673 = ~w7669 & ~w7671;
assign w7674 = ~w7672 & ~w7673;
assign w7675 = w7040 & w7047;
assign w7676 = (w7674 & w7048) | (w7674 & w16453) | (w7048 & w16453);
assign w7677 = ~w7048 & w16454;
assign w7678 = ~w7676 & ~w7677;
assign w7679 = pi142 & pi266;
assign w7680 = pi143 & pi265;
assign w7681 = ~w7679 & w7680;
assign w7682 = w7679 & ~w7680;
assign w7683 = ~w7681 & ~w7682;
assign w7684 = w7678 & w7683;
assign w7685 = ~w7678 & ~w7683;
assign w7686 = ~w7684 & ~w7685;
assign w7687 = w7563 & ~w7686;
assign w7688 = ~w7563 & w7686;
assign w7689 = ~w7687 & ~w7688;
assign w7690 = w7562 & ~w7689;
assign w7691 = ~w7562 & w7689;
assign w7692 = ~w7690 & ~w7691;
assign w7693 = (w7066 & ~w7061) | (w7066 & w15929) | (~w7061 & w15929);
assign w7694 = ~w7063 & ~w7693;
assign w7695 = w7692 & ~w7694;
assign w7696 = ~w7692 & w7694;
assign w7697 = ~w7695 & ~w7696;
assign w7698 = ~w7561 & ~w7697;
assign w7699 = w7561 & w7697;
assign w7700 = ~w7698 & ~w7699;
assign w7701 = pi146 & pi262;
assign w7702 = w7065 & w7072;
assign w7703 = ~w7073 & ~w7702;
assign w7704 = w7701 & ~w7703;
assign w7705 = ~w7701 & w7703;
assign w7706 = ~w7704 & ~w7705;
assign w7707 = w7700 & w7706;
assign w7708 = ~w7700 & ~w7706;
assign w7709 = ~w7707 & ~w7708;
assign w7710 = w7560 & ~w7709;
assign w7711 = ~w7560 & w7709;
assign w7712 = ~w7710 & ~w7711;
assign w7713 = ~w7559 & ~w7712;
assign w7714 = w7559 & w7712;
assign w7715 = ~w7713 & ~w7714;
assign w7716 = (~w7096 & ~w7083) | (~w7096 & w15930) | (~w7083 & w15930);
assign w7717 = ~w7086 & ~w7716;
assign w7718 = w7715 & w7717;
assign w7719 = ~w7715 & ~w7717;
assign w7720 = ~w7718 & ~w7719;
assign w7721 = w7558 & w7720;
assign w7722 = ~w7558 & ~w7720;
assign w7723 = ~w7721 & ~w7722;
assign w7724 = w7095 & ~w7105;
assign w7725 = pi149 & pi259;
assign w7726 = pi148 & pi260;
assign w7727 = pi150 & pi258;
assign w7728 = w7726 & ~w7727;
assign w7729 = ~w7726 & w7727;
assign w7730 = ~w7728 & ~w7729;
assign w7731 = w7725 & ~w7730;
assign w7732 = ~w7725 & w7730;
assign w7733 = ~w7731 & ~w7732;
assign w7734 = w7724 & ~w7733;
assign w7735 = ~w7724 & w7733;
assign w7736 = ~w7734 & ~w7735;
assign w7737 = w7723 & w7736;
assign w7738 = ~w7723 & ~w7736;
assign w7739 = ~w7737 & ~w7738;
assign w7740 = w7553 & ~w7739;
assign w7741 = ~w7553 & w7739;
assign w7742 = ~w7740 & ~w7741;
assign w7743 = pi322 & w7742;
assign w7744 = (~w7550 & ~w7742) | (~w7550 & w15931) | (~w7742 & w15931);
assign w7745 = w7742 & w15932;
assign w7746 = ~w7744 & ~w7745;
assign w7747 = ~w7110 & w7116;
assign w7748 = ~w7109 & ~w7747;
assign w7749 = ~w7746 & w7748;
assign w7750 = w7746 & ~w7748;
assign w7751 = ~w7749 & ~w7750;
assign w7752 = w7549 & ~w7751;
assign w7753 = ~w7549 & w7751;
assign w7754 = ~w7752 & ~w7753;
assign w7755 = w7540 & w7754;
assign w7756 = ~w7540 & ~w7754;
assign w7757 = ~w7755 & ~w7756;
assign w7758 = ~w6892 & w7122;
assign w7759 = ~w7115 & ~w7122;
assign w7760 = ~w7758 & ~w7759;
assign w7761 = w6892 & ~w7122;
assign w7762 = ~w7758 & ~w7761;
assign w7763 = ~w6891 & w7762;
assign w7764 = w6903 & ~w7763;
assign w7765 = w6891 & ~w7762;
assign w7766 = ~w7764 & ~w7765;
assign w7767 = w7760 & ~w7766;
assign w7768 = ~w7760 & w7766;
assign w7769 = ~w7767 & ~w7768;
assign w7770 = w7757 & w7769;
assign w7771 = ~w7757 & ~w7769;
assign w7772 = ~w7770 & ~w7771;
assign w7773 = w7539 & w7772;
assign w7774 = ~w7539 & ~w7772;
assign w7775 = ~w7773 & ~w7774;
assign w7776 = ~w7524 & w7775;
assign w7777 = w7524 & ~w7775;
assign w7778 = ~w7776 & ~w7777;
assign w7779 = pi329 & w3979;
assign w7780 = ~w6885 & ~w7136;
assign w7781 = w7779 & ~w7780;
assign w7782 = ~w7779 & w7780;
assign w7783 = ~w7781 & ~w7782;
assign w7784 = ~w7778 & ~w7783;
assign w7785 = w7778 & w7783;
assign w7786 = ~w7784 & ~w7785;
assign w7787 = ~w7160 & ~w7513;
assign w7788 = ~w7786 & w7787;
assign w7789 = w7786 & ~w7787;
assign w7790 = ~w7788 & ~w7789;
assign w7791 = w7519 & ~w7790;
assign w7792 = ~w7519 & w7790;
assign w7793 = ~w7791 & ~w7792;
assign w7794 = w7510 & w7793;
assign w7795 = ~w7510 & ~w7793;
assign w7796 = ~w7794 & ~w7795;
assign w7797 = w7478 & ~w7796;
assign w7798 = ~w7478 & w7796;
assign w7799 = ~w7797 & ~w7798;
assign w7800 = w7471 & ~w7799;
assign w7801 = ~w7471 & w7799;
assign w7802 = ~w7800 & ~w7801;
assign w7803 = pi336 & w1602;
assign w7804 = ~w7803 & w17694;
assign w7805 = (w7177 & w17608) | (w7177 & w17609) | (w17608 & w17609);
assign w7806 = ~w7804 & ~w7805;
assign w7807 = w7802 & ~w7806;
assign w7808 = ~w7802 & w7806;
assign w7809 = ~w7807 & ~w7808;
assign w7810 = ~w7467 & w7809;
assign w7811 = w7467 & ~w7809;
assign w7812 = ~w7810 & ~w7811;
assign w7813 = w7463 & w7812;
assign w7814 = ~w7463 & ~w7812;
assign w7815 = ~w7813 & ~w7814;
assign w7816 = w7462 & w7815;
assign w7817 = ~w7462 & ~w7815;
assign w7818 = ~w7816 & ~w7817;
assign w7819 = w7444 & ~w7818;
assign w7820 = ~w7444 & w7818;
assign w7821 = ~w7819 & ~w7820;
assign w7822 = pi340 & ~w793;
assign w7823 = ~w6833 & ~w7201;
assign w7824 = ~w7822 & w7823;
assign w7825 = w7822 & ~w7823;
assign w7826 = ~w7824 & ~w7825;
assign w7827 = w7821 & w7826;
assign w7828 = ~w7821 & ~w7826;
assign w7829 = ~w7827 & ~w7828;
assign w7830 = w7443 & w7829;
assign w7831 = ~w7443 & ~w7829;
assign w7832 = ~w7830 & ~w7831;
assign w7833 = ~w6823 & ~w7206;
assign w7834 = ~w7832 & ~w7833;
assign w7835 = w7832 & w7833;
assign w7836 = ~w7834 & ~w7835;
assign w7837 = w7438 & w7836;
assign w7838 = ~w7438 & ~w7836;
assign w7839 = ~w7837 & ~w7838;
assign w7840 = w7437 & w7839;
assign w7841 = ~w7437 & ~w7839;
assign w7842 = ~w7840 & ~w7841;
assign w7843 = w7433 & w7842;
assign w7844 = ~w7433 & ~w7842;
assign w7845 = ~w7843 & ~w7844;
assign w7846 = ~w7432 & ~w7845;
assign w7847 = w7432 & w7845;
assign w7848 = ~w7846 & ~w7847;
assign w7849 = ~w7431 & ~w7848;
assign w7850 = w7431 & w7848;
assign w7851 = ~w135 & ~w7849;
assign w7852 = ~w7850 & w7851;
assign w7853 = ~pi280 & w7852;
assign w7854 = pi280 & ~w7852;
assign w7855 = pi161 & ~w7853;
assign w7856 = ~w7854 & w7855;
assign w7857 = ~pi160 & ~w7227;
assign w7858 = ~w7856 & w7857;
assign w7859 = ~pi087 & ~pi161;
assign w7860 = pi128 & pi298;
assign w7861 = ~pi129 & w7425;
assign w7862 = pi299 & w464;
assign w7863 = ~w7425 & ~w7862;
assign w7864 = ~w7861 & ~w7863;
assign w7865 = pi300 & ~w653;
assign w7866 = pi301 & w709;
assign w7867 = pi302 & w698;
assign w7868 = ~w7401 & ~w7405;
assign w7869 = ~w7867 & w7868;
assign w7870 = w7867 & ~w7868;
assign w7871 = ~w7869 & ~w7870;
assign w7872 = pi303 & w855;
assign w7873 = ~w7395 & ~w7398;
assign w7874 = ~w7872 & w7873;
assign w7875 = w7872 & ~w7873;
assign w7876 = ~w7874 & ~w7875;
assign w7877 = pi304 & w1159;
assign w7878 = ~w7385 & ~w7389;
assign w7879 = ~w7877 & w7878;
assign w7880 = w7877 & ~w7878;
assign w7881 = ~w7879 & ~w7880;
assign w7882 = pi306 & w1420;
assign w7883 = ~w7369 & ~w7375;
assign w7884 = ~w7882 & w7883;
assign w7885 = w7882 & ~w7883;
assign w7886 = ~w7884 & ~w7885;
assign w7887 = pi307 & w1693;
assign w7888 = pi308 & w1954;
assign w7889 = ~w7355 & ~w7359;
assign w7890 = w7888 & ~w7889;
assign w7891 = ~w7888 & w7889;
assign w7892 = ~w7890 & ~w7891;
assign w7893 = pi309 & ~w2473;
assign w7894 = pi311 & w2925;
assign w7895 = ~w7331 & ~w7336;
assign w7896 = pi312 & w3304;
assign w7897 = pi314 & w4382;
assign w7898 = pi315 & w4539;
assign w7899 = pi316 & w5316;
assign w7900 = pi317 & w5862;
assign w7901 = pi318 & w6437;
assign w7902 = pi319 & w6652;
assign w7903 = pi150 & ~pi151;
assign w7904 = ~pi150 & pi151;
assign w7905 = ~w7903 & ~w7904;
assign w7906 = ~w7264 & ~w7266;
assign w7907 = w7905 & w7906;
assign w7908 = ~w7905 & ~w7906;
assign w7909 = ~w7907 & ~w7908;
assign w7910 = pi321 & w7909;
assign w7911 = pi320 & w7268;
assign w7912 = ~w7260 & ~w7273;
assign w7913 = ~w7272 & ~w7912;
assign w7914 = w7911 & ~w7913;
assign w7915 = ~w7911 & w7913;
assign w7916 = ~w7914 & ~w7915;
assign w7917 = w7910 & w7916;
assign w7918 = ~w7910 & ~w7916;
assign w7919 = ~w7917 & ~w7918;
assign w7920 = w7902 & ~w7919;
assign w7921 = ~w7902 & w7919;
assign w7922 = ~w7920 & ~w7921;
assign w7923 = ~w7278 & ~w7282;
assign w7924 = w7922 & w7923;
assign w7925 = ~w7922 & ~w7923;
assign w7926 = ~w7924 & ~w7925;
assign w7927 = ~w7901 & w7926;
assign w7928 = w7901 & ~w7926;
assign w7929 = ~w7927 & ~w7928;
assign w7930 = ~w7286 & ~w7289;
assign w7931 = w7929 & ~w7930;
assign w7932 = ~w7929 & w7930;
assign w7933 = ~w7931 & ~w7932;
assign w7934 = w7900 & w7933;
assign w7935 = ~w7900 & ~w7933;
assign w7936 = ~w7934 & ~w7935;
assign w7937 = ~w7255 & ~w7292;
assign w7938 = w7936 & w7937;
assign w7939 = ~w7936 & ~w7937;
assign w7940 = ~w7938 & ~w7939;
assign w7941 = w4539 & ~w7295;
assign w7942 = w4382 & w7306;
assign w7943 = ~w7941 & ~w7942;
assign w7944 = pi316 & ~w7943;
assign w7945 = ~w7297 & ~w7944;
assign w7946 = ~w7940 & ~w7945;
assign w7947 = w7940 & w7945;
assign w7948 = ~w7946 & ~w7947;
assign w7949 = w7899 & ~w7948;
assign w7950 = ~w7899 & w7948;
assign w7951 = ~w7949 & ~w7950;
assign w7952 = w7898 & ~w7951;
assign w7953 = ~w7898 & w7951;
assign w7954 = ~w7952 & ~w7953;
assign w7955 = ~w7250 & ~w7312;
assign w7956 = w7954 & w7955;
assign w7957 = ~w7954 & ~w7955;
assign w7958 = ~w7956 & ~w7957;
assign w7959 = w7897 & ~w7958;
assign w7960 = ~w7897 & w7958;
assign w7961 = ~w7959 & ~w7960;
assign w7962 = ~w7314 & ~w7318;
assign w7963 = w7961 & w7962;
assign w7964 = ~w7961 & ~w7962;
assign w7965 = ~w7963 & ~w7964;
assign w7966 = pi313 & w3710;
assign w7967 = ~w7965 & w7966;
assign w7968 = w7965 & ~w7966;
assign w7969 = ~w7967 & ~w7968;
assign w7970 = ~w7325 & ~w7328;
assign w7971 = ~w7969 & ~w7970;
assign w7972 = w7969 & w7970;
assign w7973 = ~w7971 & ~w7972;
assign w7974 = ~w7896 & w7973;
assign w7975 = w7896 & ~w7973;
assign w7976 = ~w7974 & ~w7975;
assign w7977 = w7895 & w7976;
assign w7978 = ~w7895 & ~w7976;
assign w7979 = ~w7977 & ~w7978;
assign w7980 = w7894 & w7979;
assign w7981 = ~w7894 & ~w7979;
assign w7982 = ~w7980 & ~w7981;
assign w7983 = ~w7340 & ~w7342;
assign w7984 = w7982 & ~w7983;
assign w7985 = ~w7982 & w7983;
assign w7986 = ~w7984 & ~w7985;
assign w7987 = ~w7347 & ~w7986;
assign w7988 = ~pi310 & ~w7986;
assign w7989 = ~w2473 & ~w7347;
assign w7990 = ~w7346 & w7986;
assign w7991 = ~w7989 & w7990;
assign w7992 = w2801 & ~w7987;
assign w7993 = ~w7988 & w7992;
assign w7994 = ~w7991 & w7993;
assign w7995 = w7347 & w7986;
assign w7996 = ~w7987 & ~w7995;
assign w7997 = ~w2801 & ~w7350;
assign w7998 = ~w7996 & w7997;
assign w7999 = ~w2801 & ~w7986;
assign w8000 = ~w7988 & ~w7999;
assign w8001 = w7346 & w8000;
assign w8002 = w2801 & w7986;
assign w8003 = ~w7989 & ~w8002;
assign w8004 = pi310 & ~w7999;
assign w8005 = ~w8003 & w8004;
assign w8006 = ~w8001 & ~w8005;
assign w8007 = ~w7243 & w8000;
assign w8008 = w8006 & w8007;
assign w8009 = ~w7994 & ~w7998;
assign w8010 = ~w8008 & w8009;
assign w8011 = ~w7893 & w8010;
assign w8012 = w7893 & ~w8010;
assign w8013 = ~w8011 & ~w8012;
assign w8014 = ~w7240 & ~w7352;
assign w8015 = w8013 & w8014;
assign w8016 = ~w8013 & ~w8014;
assign w8017 = ~w8015 & ~w8016;
assign w8018 = ~w7892 & w8017;
assign w8019 = w7892 & ~w8017;
assign w8020 = ~w8018 & ~w8019;
assign w8021 = w7887 & ~w8020;
assign w8022 = ~w7887 & w8020;
assign w8023 = ~w8021 & ~w8022;
assign w8024 = ~w7364 & ~w7367;
assign w8025 = w8023 & w8024;
assign w8026 = ~w8023 & ~w8024;
assign w8027 = ~w8025 & ~w8026;
assign w8028 = w7886 & w8027;
assign w8029 = ~w7886 & ~w8027;
assign w8030 = ~w8028 & ~w8029;
assign w8031 = pi305 & w1220;
assign w8032 = w8030 & w8031;
assign w8033 = ~w8030 & ~w8031;
assign w8034 = ~w8032 & ~w8033;
assign w8035 = ~w7379 & ~w7382;
assign w8036 = w8034 & ~w8035;
assign w8037 = ~w8034 & w8035;
assign w8038 = ~w8036 & ~w8037;
assign w8039 = w7881 & w8038;
assign w8040 = ~w7881 & ~w8038;
assign w8041 = ~w8039 & ~w8040;
assign w8042 = ~w7876 & ~w8041;
assign w8043 = w7876 & w8041;
assign w8044 = ~w8042 & ~w8043;
assign w8045 = w7871 & w8044;
assign w8046 = ~w7871 & ~w8044;
assign w8047 = ~w8045 & ~w8046;
assign w8048 = w7866 & w8047;
assign w8049 = ~w7866 & ~w8047;
assign w8050 = ~w8048 & ~w8049;
assign w8051 = pi130 & w7416;
assign w8052 = w464 & ~w653;
assign w8053 = ~w6806 & w8052;
assign w8054 = ~w8051 & ~w8053;
assign w8055 = pi301 & ~w8054;
assign w8056 = ~w7419 & ~w8055;
assign w8057 = ~w8050 & w8056;
assign w8058 = w8050 & ~w8056;
assign w8059 = ~w8057 & ~w8058;
assign w8060 = w7407 & w8055;
assign w8061 = ~w8056 & ~w8060;
assign w8062 = ~w7230 & ~w7420;
assign w8063 = ~w8061 & w8062;
assign w8064 = ~w7231 & ~w8063;
assign w8065 = w8059 & ~w8064;
assign w8066 = ~w8059 & w8064;
assign w8067 = ~w8065 & ~w8066;
assign w8068 = w7865 & w8067;
assign w8069 = ~w7865 & ~w8067;
assign w8070 = ~w8068 & ~w8069;
assign w8071 = w7864 & w8070;
assign w8072 = ~w7864 & ~w8070;
assign w8073 = ~w8071 & ~w8072;
assign w8074 = w7860 & w8073;
assign w8075 = ~w7860 & ~w8073;
assign w8076 = ~w8074 & ~w8075;
assign w8077 = pi280 & w7848;
assign w8078 = ~w7846 & ~w8077;
assign w8079 = ~pi281 & w8078;
assign w8080 = pi281 & ~w8078;
assign w8081 = ~w8079 & ~w8080;
assign w8082 = pi345 & w456;
assign w8083 = pi344 & w466;
assign w8084 = pi343 & ~w537;
assign w8085 = (~w7436 & ~w7839) | (~w7436 & w17610) | (~w7839 & w17610);
assign w8086 = w8084 & ~w8085;
assign w8087 = ~w8084 & w8085;
assign w8088 = ~w8086 & ~w8087;
assign w8089 = pi340 & ~w955;
assign w8090 = ~w7824 & ~w7827;
assign w8091 = w8089 & w8090;
assign w8092 = ~w8089 & ~w8090;
assign w8093 = ~w8091 & ~w8092;
assign w8094 = pi338 & w1339;
assign w8095 = w7445 & ~w7812;
assign w8096 = ~w6844 & ~w7193;
assign w8097 = ~w1101 & w7812;
assign w8098 = w6843 & ~w8096;
assign w8099 = ~w8097 & w8098;
assign w8100 = ~w8095 & ~w8099;
assign w8101 = w8094 & ~w8100;
assign w8102 = ~w8094 & w8100;
assign w8103 = ~w8101 & ~w8102;
assign w8104 = pi337 & w1602;
assign w8105 = ~w7466 & ~w7811;
assign w8106 = w8104 & w8105;
assign w8107 = ~w8104 & ~w8105;
assign w8108 = ~w8106 & ~w8107;
assign w8109 = pi336 & ~w1865;
assign w8110 = ~w7805 & ~w7808;
assign w8111 = w8109 & ~w8110;
assign w8112 = ~w8109 & w8110;
assign w8113 = ~w8111 & ~w8112;
assign w8114 = pi333 & w2698;
assign w8115 = pi334 & ~w2373;
assign w8116 = (w8115 & w7797) | (w8115 & w16456) | (w7797 & w16456);
assign w8117 = ~w7797 & w16457;
assign w8118 = ~w8116 & ~w8117;
assign w8119 = w8114 & ~w8118;
assign w8120 = ~w8114 & w8118;
assign w8121 = ~w8119 & ~w8120;
assign w8122 = pi335 & ~w2170;
assign w8123 = ~w7479 & ~w7519;
assign w8124 = w7479 & w7519;
assign w8125 = ~w7504 & w7790;
assign w8126 = w7504 & ~w7790;
assign w8127 = ~w8125 & ~w8126;
assign w8128 = w7490 & w8127;
assign w8129 = ~w7490 & ~w8127;
assign w8130 = ~w8128 & ~w8129;
assign w8131 = ~w8124 & ~w8130;
assign w8132 = ~w8123 & ~w8131;
assign w8133 = w8122 & ~w8132;
assign w8134 = ~w8122 & w8132;
assign w8135 = ~w8133 & ~w8134;
assign w8136 = ~w8121 & w8135;
assign w8137 = w8121 & ~w8135;
assign w8138 = ~w8136 & ~w8137;
assign w8139 = pi332 & ~w3183;
assign w8140 = pi332 & w6871;
assign w8141 = ~w7517 & ~w8140;
assign w8142 = w7480 & ~w8141;
assign w8143 = ~w7480 & w8141;
assign w8144 = ~w8127 & ~w8143;
assign w8145 = ~w8142 & ~w8144;
assign w8146 = ~w8139 & w8145;
assign w8147 = w8139 & ~w8145;
assign w8148 = ~w8146 & ~w8147;
assign w8149 = ~w7499 & w7501;
assign w8150 = w7786 & ~w8149;
assign w8151 = ~w7496 & w7499;
assign w8152 = ~w8150 & ~w8151;
assign w8153 = pi330 & w3979;
assign w8154 = w8152 & ~w8153;
assign w8155 = ~w8152 & w8153;
assign w8156 = ~w8154 & ~w8155;
assign w8157 = ~w7522 & ~w7777;
assign w8158 = ~w7755 & ~w7760;
assign w8159 = ~w7756 & ~w8158;
assign w8160 = ~w7745 & ~w7748;
assign w8161 = ~w7744 & ~w8160;
assign w8162 = pi323 & w7742;
assign w8163 = ~w7551 & ~w7739;
assign w8164 = ~w7552 & w7739;
assign w8165 = ~w8163 & ~w8164;
assign w8166 = pi151 & pi258;
assign w8167 = pi150 & pi259;
assign w8168 = (~w8167 & ~w7739) | (~w8167 & w15933) | (~w7739 & w15933);
assign w8169 = w7739 & w15934;
assign w8170 = ~w8168 & ~w8169;
assign w8171 = pi259 & w7724;
assign w8172 = w7558 & w7726;
assign w8173 = ~w7558 & ~w7726;
assign w8174 = ~w8172 & ~w8173;
assign w8175 = ~w7720 & ~w8174;
assign w8176 = ~w7724 & ~w7725;
assign w8177 = w7720 & w8174;
assign w8178 = ~w8175 & ~w8176;
assign w8179 = (~w8171 & ~w8178) | (~w8171 & w16194) | (~w8178 & w16194);
assign w8180 = (~w8172 & ~w7720) | (~w8172 & w15935) | (~w7720 & w15935);
assign w8181 = pi146 & pi263;
assign w8182 = pi143 & pi266;
assign w8183 = ~w7667 & ~w7672;
assign w8184 = pi140 & pi269;
assign w8185 = ~w7653 & ~w7657;
assign w8186 = ~w7652 & ~w8185;
assign w8187 = pi137 & pi272;
assign w8188 = pi136 & pi273;
assign w8189 = pi135 & pi274;
assign w8190 = ~w7621 & ~w7626;
assign w8191 = pi134 & pi275;
assign w8192 = pi133 & pi276;
assign w8193 = pi132 & pi277;
assign w8194 = pi131 & pi278;
assign w8195 = pi130 & pi279;
assign w8196 = w7576 & ~w7579;
assign w8197 = ~w7581 & ~w8196;
assign w8198 = pi128 & pi281;
assign w8199 = pi129 & pi280;
assign w8200 = ~w8198 & ~w8199;
assign w8201 = pi129 & pi281;
assign w8202 = w7576 & w8201;
assign w8203 = ~w8200 & ~w8202;
assign w8204 = w8197 & ~w8203;
assign w8205 = ~w8197 & w8203;
assign w8206 = ~w8204 & ~w8205;
assign w8207 = w8195 & w8206;
assign w8208 = ~w8195 & ~w8206;
assign w8209 = ~w8207 & ~w8208;
assign w8210 = ~w7587 & ~w7590;
assign w8211 = w8209 & w8210;
assign w8212 = ~w8209 & ~w8210;
assign w8213 = ~w8211 & ~w8212;
assign w8214 = w8194 & w8213;
assign w8215 = ~w8194 & ~w8213;
assign w8216 = ~w8214 & ~w8215;
assign w8217 = ~w7593 & ~w7597;
assign w8218 = ~w8216 & w8217;
assign w8219 = w8216 & ~w8217;
assign w8220 = ~w8218 & ~w8219;
assign w8221 = w8193 & w8220;
assign w8222 = ~w8193 & ~w8220;
assign w8223 = ~w8221 & ~w8222;
assign w8224 = ~w7601 & ~w7604;
assign w8225 = w8223 & ~w8224;
assign w8226 = ~w8223 & w8224;
assign w8227 = ~w8225 & ~w8226;
assign w8228 = ~w8192 & w8227;
assign w8229 = w8192 & ~w8227;
assign w8230 = ~w8228 & ~w8229;
assign w8231 = ~w7607 & ~w7612;
assign w8232 = w8230 & ~w8231;
assign w8233 = ~w8230 & w8231;
assign w8234 = ~w8232 & ~w8233;
assign w8235 = ~w8191 & ~w8234;
assign w8236 = w8191 & w8234;
assign w8237 = ~w8235 & ~w8236;
assign w8238 = ~w7615 & ~w7617;
assign w8239 = w8237 & w8238;
assign w8240 = ~w8237 & ~w8238;
assign w8241 = ~w8239 & ~w8240;
assign w8242 = ~w8190 & ~w8241;
assign w8243 = w8190 & w8241;
assign w8244 = ~w8242 & ~w8243;
assign w8245 = w8189 & ~w8244;
assign w8246 = ~w8189 & w8244;
assign w8247 = ~w8245 & ~w8246;
assign w8248 = ~w8188 & w8247;
assign w8249 = w8188 & ~w8247;
assign w8250 = ~w8248 & ~w8249;
assign w8251 = ~w7631 & ~w7634;
assign w8252 = ~w7630 & ~w8251;
assign w8253 = ~w8250 & w8252;
assign w8254 = w8250 & ~w8252;
assign w8255 = ~w8253 & ~w8254;
assign w8256 = ~w8187 & w8255;
assign w8257 = w8187 & ~w8255;
assign w8258 = ~w8256 & ~w8257;
assign w8259 = ~w7633 & w7640;
assign w8260 = ~w7641 & ~w8259;
assign w8261 = w8258 & w8260;
assign w8262 = ~w8258 & ~w8260;
assign w8263 = ~w8261 & ~w8262;
assign w8264 = ~w7644 & ~w7649;
assign w8265 = w8263 & ~w8264;
assign w8266 = ~w8263 & w8264;
assign w8267 = ~w8265 & ~w8266;
assign w8268 = pi139 & pi270;
assign w8269 = pi138 & pi271;
assign w8270 = w8268 & ~w8269;
assign w8271 = ~w8268 & w8269;
assign w8272 = ~w8270 & ~w8271;
assign w8273 = w8267 & w8272;
assign w8274 = ~w8267 & ~w8272;
assign w8275 = ~w8273 & ~w8274;
assign w8276 = w8186 & ~w8275;
assign w8277 = ~w8186 & w8275;
assign w8278 = ~w8276 & ~w8277;
assign w8279 = ~w8184 & ~w8278;
assign w8280 = w8184 & w8278;
assign w8281 = ~w8279 & ~w8280;
assign w8282 = ~w7655 & w7663;
assign w8283 = ~w7664 & ~w8282;
assign w8284 = w8281 & w8283;
assign w8285 = ~w8281 & ~w8283;
assign w8286 = ~w8284 & ~w8285;
assign w8287 = ~w8183 & w8286;
assign w8288 = w8183 & ~w8286;
assign w8289 = ~w8287 & ~w8288;
assign w8290 = pi142 & pi267;
assign w8291 = pi141 & pi268;
assign w8292 = w8290 & ~w8291;
assign w8293 = ~w8290 & w8291;
assign w8294 = ~w8292 & ~w8293;
assign w8295 = w8289 & w8294;
assign w8296 = ~w8289 & ~w8294;
assign w8297 = ~w8295 & ~w8296;
assign w8298 = ~w7679 & ~w7676;
assign w8299 = ~w7677 & ~w8298;
assign w8300 = ~w8297 & w8299;
assign w8301 = w8297 & ~w8299;
assign w8302 = ~w8300 & ~w8301;
assign w8303 = w8182 & w8302;
assign w8304 = ~w8182 & ~w8302;
assign w8305 = ~w8303 & ~w8304;
assign w8306 = ~w7680 & w7686;
assign w8307 = ~w7687 & ~w8306;
assign w8308 = w8305 & ~w8307;
assign w8309 = ~w8305 & w8307;
assign w8310 = ~w8308 & ~w8309;
assign w8311 = (~w7690 & w7694) | (~w7690 & w16612) | (w7694 & w16612);
assign w8312 = w8310 & w8311;
assign w8313 = ~w8310 & ~w8311;
assign w8314 = ~w8312 & ~w8313;
assign w8315 = pi145 & pi264;
assign w8316 = pi144 & pi265;
assign w8317 = w8315 & ~w8316;
assign w8318 = ~w8315 & w8316;
assign w8319 = ~w8317 & ~w8318;
assign w8320 = w8314 & w8319;
assign w8321 = ~w8314 & ~w8319;
assign w8322 = ~w8320 & ~w8321;
assign w8323 = ~w7698 & ~w7703;
assign w8324 = ~w7699 & ~w8323;
assign w8325 = ~w8322 & ~w8324;
assign w8326 = w8322 & w8324;
assign w8327 = ~w8325 & ~w8326;
assign w8328 = w8181 & w8327;
assign w8329 = ~w8181 & ~w8327;
assign w8330 = ~w8328 & ~w8329;
assign w8331 = w7701 & ~w7709;
assign w8332 = ~w7711 & ~w8331;
assign w8333 = w8330 & ~w8332;
assign w8334 = ~w8330 & w8332;
assign w8335 = ~w8333 & ~w8334;
assign w8336 = ~w7714 & ~w7717;
assign w8337 = ~w7713 & ~w8336;
assign w8338 = ~w8335 & ~w8337;
assign w8339 = w8335 & w8337;
assign w8340 = ~w8338 & ~w8339;
assign w8341 = pi149 & pi260;
assign w8342 = pi148 & pi261;
assign w8343 = pi147 & pi262;
assign w8344 = ~w8342 & w8343;
assign w8345 = w8342 & ~w8343;
assign w8346 = ~w8344 & ~w8345;
assign w8347 = w8341 & ~w8346;
assign w8348 = ~w8341 & w8346;
assign w8349 = ~w8347 & ~w8348;
assign w8350 = w8340 & ~w8349;
assign w8351 = ~w8340 & w8349;
assign w8352 = ~w8350 & ~w8351;
assign w8353 = w8180 & ~w8352;
assign w8354 = ~w8180 & w8352;
assign w8355 = ~w8353 & ~w8354;
assign w8356 = w8179 & w8355;
assign w8357 = ~w8179 & ~w8355;
assign w8358 = ~w8356 & ~w8357;
assign w8359 = w8170 & w8358;
assign w8360 = ~w8170 & ~w8358;
assign w8361 = ~w8359 & ~w8360;
assign w8362 = ~w8166 & ~w8361;
assign w8363 = w8166 & w8361;
assign w8364 = ~w8362 & ~w8363;
assign w8365 = w8165 & ~w8364;
assign w8366 = ~w8165 & w8364;
assign w8367 = ~w8365 & ~w8366;
assign w8368 = (w8162 & w8367) | (w8162 & w15936) | (w8367 & w15936);
assign w8369 = ~w8367 & w15937;
assign w8370 = ~w8368 & ~w8369;
assign w8371 = w8161 & ~w8370;
assign w8372 = ~w8161 & w8370;
assign w8373 = ~w8371 & ~w8372;
assign w8374 = pi325 & w6283;
assign w8375 = pi324 & ~w7108;
assign w8376 = ~w7548 & ~w7752;
assign w8377 = ~w8375 & w8376;
assign w8378 = w8375 & ~w8376;
assign w8379 = ~w8377 & ~w8378;
assign w8380 = w8374 & ~w8379;
assign w8381 = ~w8374 & w8379;
assign w8382 = ~w8380 & ~w8381;
assign w8383 = w8373 & w8382;
assign w8384 = ~w8373 & ~w8382;
assign w8385 = ~w8383 & ~w8384;
assign w8386 = w8159 & ~w8385;
assign w8387 = ~w8159 & w8385;
assign w8388 = ~w8386 & ~w8387;
assign w8389 = w7526 & w7536;
assign w8390 = ~w7526 & ~w7536;
assign w8391 = w7525 & w7772;
assign w8392 = (~w8390 & w7772) | (~w8390 & w16195) | (w7772 & w16195);
assign w8393 = ~w8391 & w8392;
assign w8394 = ~w8389 & ~w8393;
assign w8395 = ~w7766 & ~w7772;
assign w8396 = ~w8391 & ~w8395;
assign w8397 = pi327 & w5194;
assign w8398 = pi326 & w5714;
assign w8399 = w8397 & ~w8398;
assign w8400 = ~w8397 & w8398;
assign w8401 = ~w8399 & ~w8400;
assign w8402 = w8396 & ~w8401;
assign w8403 = ~w8396 & w8401;
assign w8404 = ~w8402 & ~w8403;
assign w8405 = w8394 & ~w8404;
assign w8406 = ~w8394 & w8404;
assign w8407 = ~w8405 & ~w8406;
assign w8408 = w8388 & w8407;
assign w8409 = ~w8388 & ~w8407;
assign w8410 = ~w8408 & ~w8409;
assign w8411 = w8157 & w8410;
assign w8412 = ~w8157 & ~w8410;
assign w8413 = ~w8411 & ~w8412;
assign w8414 = pi328 & ~w4854;
assign w8415 = (~w7781 & ~w7778) | (~w7781 & w16196) | (~w7778 & w16196);
assign w8416 = pi329 & ~w4708;
assign w8417 = ~w8415 & w8416;
assign w8418 = w8415 & ~w8416;
assign w8419 = ~w8417 & ~w8418;
assign w8420 = w8414 & ~w8419;
assign w8421 = ~w8414 & w8419;
assign w8422 = ~w8420 & ~w8421;
assign w8423 = w8413 & w8422;
assign w8424 = ~w8413 & ~w8422;
assign w8425 = ~w8423 & ~w8424;
assign w8426 = w8156 & ~w8425;
assign w8427 = ~w8156 & w8425;
assign w8428 = ~w8426 & ~w8427;
assign w8429 = w7491 & ~w7787;
assign w8430 = w8150 & ~w8151;
assign w8431 = w7501 & ~w7786;
assign w8432 = ~w7491 & w7787;
assign w8433 = ~w8431 & ~w8432;
assign w8434 = ~w8430 & w8433;
assign w8435 = ~w8429 & ~w8434;
assign w8436 = pi331 & ~w3568;
assign w8437 = w8435 & ~w8436;
assign w8438 = ~w8435 & w8436;
assign w8439 = ~w8437 & ~w8438;
assign w8440 = w8428 & w8439;
assign w8441 = ~w8428 & ~w8439;
assign w8442 = ~w8440 & ~w8441;
assign w8443 = w8148 & w8442;
assign w8444 = ~w8148 & ~w8442;
assign w8445 = ~w8443 & ~w8444;
assign w8446 = ~w7469 & ~w7800;
assign w8447 = ~w8445 & w8446;
assign w8448 = w8445 & ~w8446;
assign w8449 = ~w8447 & ~w8448;
assign w8450 = w8138 & w8449;
assign w8451 = ~w8138 & ~w8449;
assign w8452 = ~w8450 & ~w8451;
assign w8453 = w8113 & ~w8452;
assign w8454 = ~w8113 & w8452;
assign w8455 = ~w8453 & ~w8454;
assign w8456 = w8108 & ~w8455;
assign w8457 = ~w8108 & w8455;
assign w8458 = ~w8456 & ~w8457;
assign w8459 = ~w8103 & ~w8458;
assign w8460 = w8103 & w8458;
assign w8461 = ~w8459 & ~w8460;
assign w8462 = ~w7463 & ~w7818;
assign w8463 = ~w7820 & ~w8462;
assign w8464 = pi339 & w1101;
assign w8465 = ~w8463 & ~w8464;
assign w8466 = w8463 & w8464;
assign w8467 = ~w8465 & ~w8466;
assign w8468 = ~w8461 & ~w8467;
assign w8469 = w8461 & w8467;
assign w8470 = ~w8468 & ~w8469;
assign w8471 = w8093 & ~w8470;
assign w8472 = ~w8093 & w8470;
assign w8473 = ~w8471 & ~w8472;
assign w8474 = ~w7441 & ~w7830;
assign w8475 = pi341 & ~w793;
assign w8476 = w8474 & w8475;
assign w8477 = ~w8474 & ~w8475;
assign w8478 = ~w8476 & ~w8477;
assign w8479 = w8473 & ~w8478;
assign w8480 = ~w8473 & w8478;
assign w8481 = ~w8479 & ~w8480;
assign w8482 = pi342 & ~w615;
assign w8483 = w537 & ~w7834;
assign w8484 = ~w7835 & w8482;
assign w8485 = ~w8483 & w8484;
assign w8486 = ~w7834 & ~w8482;
assign w8487 = ~w7837 & w8486;
assign w8488 = ~w8485 & ~w8487;
assign w8489 = w8481 & w8488;
assign w8490 = ~w8481 & ~w8488;
assign w8491 = ~w8489 & ~w8490;
assign w8492 = w8088 & w8491;
assign w8493 = ~w8088 & ~w8491;
assign w8494 = ~w8492 & ~w8493;
assign w8495 = w7843 & w8494;
assign w8496 = ~w7843 & ~w8494;
assign w8497 = ~w8495 & ~w8496;
assign w8498 = w8083 & ~w8497;
assign w8499 = ~w8083 & w8497;
assign w8500 = ~w8498 & ~w8499;
assign w8501 = ~w8082 & w8500;
assign w8502 = w8082 & ~w8500;
assign w8503 = ~w8501 & ~w8502;
assign w8504 = w8081 & ~w8503;
assign w8505 = ~w8081 & w8503;
assign w8506 = ~w8504 & ~w8505;
assign w8507 = w8076 & ~w8506;
assign w8508 = ~w8076 & w8506;
assign w8509 = ~w8507 & ~w8508;
assign w8510 = ~pi280 & ~w7848;
assign w8511 = ~w7429 & ~w8077;
assign w8512 = ~w8510 & w8511;
assign w8513 = ~w7430 & ~w8512;
assign w8514 = ~w8509 & w8513;
assign w8515 = w8509 & ~w8513;
assign w8516 = ~w135 & ~w8514;
assign w8517 = ~w8515 & w8516;
assign w8518 = pi161 & ~w189;
assign w8519 = ~w8517 & w8518;
assign w8520 = ~pi160 & ~w7859;
assign w8521 = ~w8519 & w8520;
assign w8522 = ~pi088 & ~pi161;
assign w8523 = pi346 & w456;
assign w8524 = w466 & w8502;
assign w8525 = pi345 & w466;
assign w8526 = ~w8502 & ~w8525;
assign w8527 = ~w8524 & ~w8526;
assign w8528 = pi344 & ~w537;
assign w8529 = ~w466 & ~w8495;
assign w8530 = ~w8496 & ~w8529;
assign w8531 = w8528 & w8530;
assign w8532 = ~w8499 & w8530;
assign w8533 = ~w8528 & ~w8532;
assign w8534 = ~w8531 & ~w8533;
assign w8535 = ~w8086 & ~w8492;
assign w8536 = pi343 & ~w615;
assign w8537 = w8535 & ~w8536;
assign w8538 = ~w8535 & w8536;
assign w8539 = ~w8537 & ~w8538;
assign w8540 = pi342 & ~w793;
assign w8541 = ~w8485 & ~w8489;
assign w8542 = w8540 & ~w8541;
assign w8543 = ~w8540 & w8541;
assign w8544 = ~w8542 & ~w8543;
assign w8545 = pi340 & w1101;
assign w8546 = ~w8092 & ~w8471;
assign w8547 = ~w8545 & ~w8546;
assign w8548 = w8545 & w8546;
assign w8549 = ~w8547 & ~w8548;
assign w8550 = ~w8101 & ~w8460;
assign w8551 = ~w1602 & w8550;
assign w8552 = w1602 & ~w8550;
assign w8553 = pi338 & ~w8551;
assign w8554 = ~w8552 & w8553;
assign w8555 = pi337 & ~w1865;
assign w8556 = ~w8106 & ~w8456;
assign w8557 = w8555 & ~w8556;
assign w8558 = ~w8555 & w8556;
assign w8559 = ~w8557 & ~w8558;
assign w8560 = pi336 & ~w2170;
assign w8561 = ~w8112 & ~w8453;
assign w8562 = ~w8560 & ~w8561;
assign w8563 = w8560 & w8561;
assign w8564 = ~w8562 & ~w8563;
assign w8565 = pi333 & ~w3183;
assign w8566 = ~w8132 & ~w8445;
assign w8567 = w8132 & w8445;
assign w8568 = (~w8114 & ~w8445) | (~w8114 & w16197) | (~w8445 & w16197);
assign w8569 = ~w8566 & ~w8568;
assign w8570 = w8565 & w8569;
assign w8571 = ~w8565 & ~w8569;
assign w8572 = ~w8570 & ~w8571;
assign w8573 = pi331 & w3979;
assign w8574 = (~w8438 & ~w8428) | (~w8438 & w16458) | (~w8428 & w16458);
assign w8575 = ~w8573 & w8574;
assign w8576 = w8573 & ~w8574;
assign w8577 = ~w8575 & ~w8576;
assign w8578 = pi330 & ~w4708;
assign w8579 = ~w8155 & ~w8426;
assign w8580 = ~w8578 & w8579;
assign w8581 = w8578 & ~w8579;
assign w8582 = ~w8580 & ~w8581;
assign w8583 = ~w8417 & ~w8425;
assign w8584 = ~w8418 & ~w8583;
assign w8585 = ~w8396 & w8398;
assign w8586 = w8396 & ~w8398;
assign w8587 = ~w8585 & ~w8586;
assign w8588 = w8388 & w8587;
assign w8589 = ~w8388 & ~w8587;
assign w8590 = ~w8588 & ~w8589;
assign w8591 = w8397 & w8590;
assign w8592 = ~w8397 & ~w8590;
assign w8593 = ~w8394 & ~w8592;
assign w8594 = ~w8591 & ~w8593;
assign w8595 = w8374 & w8385;
assign w8596 = ~w8386 & ~w8595;
assign w8597 = pi324 & w7742;
assign w8598 = pi151 & pi259;
assign w8599 = ~w8164 & w8364;
assign w8600 = ~w8598 & w17695;
assign w8601 = (w8364 & w16198) | (w8364 & w16199) | (w16198 & w16199);
assign w8602 = ~w8600 & ~w8601;
assign w8603 = pi150 & pi260;
assign w8604 = (~w8169 & ~w8358) | (~w8169 & w16200) | (~w8358 & w16200);
assign w8605 = w8603 & ~w8604;
assign w8606 = ~w8603 & w8604;
assign w8607 = ~w8605 & ~w8606;
assign w8608 = w8340 & w8344;
assign w8609 = ~w8342 & ~w8343;
assign w8610 = ~w8340 & w8609;
assign w8611 = ~w8608 & ~w8610;
assign w8612 = ~w8180 & w8611;
assign w8613 = pi148 & pi262;
assign w8614 = w8340 & w8345;
assign w8615 = w8342 & w8343;
assign w8616 = ~w8340 & w8615;
assign w8617 = ~w8614 & ~w8616;
assign w8618 = w8613 & w8617;
assign w8619 = ~w8612 & w8618;
assign w8620 = ~w8613 & ~w8617;
assign w8621 = ~w8180 & ~w8613;
assign w8622 = w8611 & w8621;
assign w8623 = ~w8620 & ~w8622;
assign w8624 = ~w8619 & w8623;
assign w8625 = pi147 & pi263;
assign w8626 = (~w8328 & ~w8330) | (~w8328 & w17611) | (~w8330 & w17611);
assign w8627 = pi145 & pi265;
assign w8628 = pi144 & pi266;
assign w8629 = ~w8304 & ~w8308;
assign w8630 = pi142 & pi268;
assign w8631 = pi141 & pi269;
assign w8632 = pi140 & pi270;
assign w8633 = ~w8280 & ~w8283;
assign w8634 = ~w8279 & ~w8633;
assign w8635 = w8632 & w8634;
assign w8636 = ~w8632 & ~w8634;
assign w8637 = ~w8635 & ~w8636;
assign w8638 = w8268 & w8275;
assign w8639 = ~w8276 & ~w8638;
assign w8640 = pi139 & pi271;
assign w8641 = pi138 & pi272;
assign w8642 = ~w8265 & ~w8269;
assign w8643 = ~w8266 & ~w8642;
assign w8644 = ~w8641 & ~w8643;
assign w8645 = w8641 & w8643;
assign w8646 = ~w8644 & ~w8645;
assign w8647 = pi137 & pi273;
assign w8648 = ~w8257 & ~w8261;
assign w8649 = pi136 & pi274;
assign w8650 = ~w8248 & ~w8254;
assign w8651 = pi135 & pi275;
assign w8652 = pi134 & pi276;
assign w8653 = pi133 & pi277;
assign w8654 = pi132 & pi278;
assign w8655 = ~w8222 & ~w8225;
assign w8656 = ~w8654 & ~w8655;
assign w8657 = w8654 & w8655;
assign w8658 = ~w8656 & ~w8657;
assign w8659 = pi131 & pi279;
assign w8660 = pi130 & pi280;
assign w8661 = pi128 & pi282;
assign w8662 = ~w8202 & ~w8205;
assign w8663 = w8661 & ~w8662;
assign w8664 = ~w8661 & w8662;
assign w8665 = ~w8663 & ~w8664;
assign w8666 = w8201 & w8665;
assign w8667 = ~w8201 & ~w8665;
assign w8668 = ~w8666 & ~w8667;
assign w8669 = w8660 & w8668;
assign w8670 = ~w8660 & ~w8668;
assign w8671 = ~w8669 & ~w8670;
assign w8672 = ~w8207 & ~w8211;
assign w8673 = w8671 & w8672;
assign w8674 = ~w8671 & ~w8672;
assign w8675 = ~w8673 & ~w8674;
assign w8676 = w8659 & ~w8675;
assign w8677 = ~w8659 & w8675;
assign w8678 = ~w8676 & ~w8677;
assign w8679 = ~w8214 & ~w8219;
assign w8680 = w8678 & ~w8679;
assign w8681 = ~w8678 & w8679;
assign w8682 = ~w8680 & ~w8681;
assign w8683 = w8658 & w8682;
assign w8684 = ~w8658 & ~w8682;
assign w8685 = ~w8683 & ~w8684;
assign w8686 = ~w8229 & ~w8232;
assign w8687 = w8685 & ~w8686;
assign w8688 = ~w8685 & w8686;
assign w8689 = ~w8687 & ~w8688;
assign w8690 = w8653 & ~w8689;
assign w8691 = ~w8653 & w8689;
assign w8692 = ~w8690 & ~w8691;
assign w8693 = ~w8236 & ~w8239;
assign w8694 = ~w8692 & ~w8693;
assign w8695 = w8692 & w8693;
assign w8696 = ~w8694 & ~w8695;
assign w8697 = w8652 & w8696;
assign w8698 = ~w8652 & ~w8696;
assign w8699 = ~w8697 & ~w8698;
assign w8700 = w8651 & w8699;
assign w8701 = ~w8651 & ~w8699;
assign w8702 = ~w8700 & ~w8701;
assign w8703 = ~w8242 & ~w8246;
assign w8704 = ~w8702 & w8703;
assign w8705 = w8702 & ~w8703;
assign w8706 = ~w8704 & ~w8705;
assign w8707 = ~w8650 & w8706;
assign w8708 = w8650 & ~w8706;
assign w8709 = ~w8707 & ~w8708;
assign w8710 = w8649 & ~w8709;
assign w8711 = ~w8649 & w8709;
assign w8712 = ~w8710 & ~w8711;
assign w8713 = ~w8648 & ~w8712;
assign w8714 = w8648 & w8712;
assign w8715 = ~w8713 & ~w8714;
assign w8716 = w8647 & ~w8715;
assign w8717 = ~w8647 & w8715;
assign w8718 = ~w8716 & ~w8717;
assign w8719 = w8646 & ~w8718;
assign w8720 = ~w8646 & w8718;
assign w8721 = ~w8719 & ~w8720;
assign w8722 = ~w8640 & ~w8721;
assign w8723 = w8640 & w8721;
assign w8724 = ~w8722 & ~w8723;
assign w8725 = w8639 & ~w8724;
assign w8726 = ~w8639 & w8724;
assign w8727 = ~w8725 & ~w8726;
assign w8728 = ~w8637 & w8727;
assign w8729 = w8637 & ~w8727;
assign w8730 = ~w8728 & ~w8729;
assign w8731 = w8631 & ~w8730;
assign w8732 = ~w8631 & w8730;
assign w8733 = ~w8731 & ~w8732;
assign w8734 = ~w8287 & ~w8291;
assign w8735 = ~w8288 & ~w8734;
assign w8736 = w8733 & w8735;
assign w8737 = ~w8733 & ~w8735;
assign w8738 = ~w8736 & ~w8737;
assign w8739 = ~w8630 & ~w8738;
assign w8740 = w8630 & w8738;
assign w8741 = ~w8739 & ~w8740;
assign w8742 = pi143 & pi267;
assign w8743 = w8290 & w8297;
assign w8744 = ~w8300 & ~w8743;
assign w8745 = w8742 & ~w8744;
assign w8746 = ~w8742 & w8744;
assign w8747 = ~w8745 & ~w8746;
assign w8748 = w8741 & ~w8747;
assign w8749 = ~w8741 & w8747;
assign w8750 = ~w8748 & ~w8749;
assign w8751 = w8629 & ~w8750;
assign w8752 = ~w8629 & w8750;
assign w8753 = ~w8751 & ~w8752;
assign w8754 = w8628 & w8753;
assign w8755 = ~w8628 & ~w8753;
assign w8756 = ~w8754 & ~w8755;
assign w8757 = (w8316 & ~w8311) | (w8316 & w16459) | (~w8311 & w16459);
assign w8758 = ~w8313 & ~w8757;
assign w8759 = w8756 & ~w8758;
assign w8760 = ~w8756 & w8758;
assign w8761 = ~w8759 & ~w8760;
assign w8762 = ~w8627 & ~w8761;
assign w8763 = w8627 & w8761;
assign w8764 = ~w8762 & ~w8763;
assign w8765 = pi146 & pi264;
assign w8766 = w8315 & w8322;
assign w8767 = ~w8325 & ~w8766;
assign w8768 = w8765 & ~w8767;
assign w8769 = ~w8765 & w8767;
assign w8770 = ~w8768 & ~w8769;
assign w8771 = w8764 & ~w8770;
assign w8772 = ~w8764 & w8770;
assign w8773 = ~w8771 & ~w8772;
assign w8774 = w8626 & ~w8773;
assign w8775 = ~w8626 & w8773;
assign w8776 = ~w8774 & ~w8775;
assign w8777 = w8625 & ~w8776;
assign w8778 = ~w8625 & w8776;
assign w8779 = ~w8777 & ~w8778;
assign w8780 = ~w8339 & ~w8343;
assign w8781 = ~w8338 & ~w8780;
assign w8782 = w8779 & w8781;
assign w8783 = ~w8779 & ~w8781;
assign w8784 = ~w8782 & ~w8783;
assign w8785 = w8624 & w8784;
assign w8786 = ~w8624 & ~w8784;
assign w8787 = ~w8785 & ~w8786;
assign w8788 = ~w8179 & w8341;
assign w8789 = w8179 & ~w8341;
assign w8790 = w8611 & w8617;
assign w8791 = w8180 & ~w8790;
assign w8792 = ~w8180 & w8790;
assign w8793 = ~w8791 & ~w8792;
assign w8794 = (~w8788 & ~w8793) | (~w8788 & w15939) | (~w8793 & w15939);
assign w8795 = ~w8787 & ~w8794;
assign w8796 = w8787 & w8794;
assign w8797 = ~w8795 & ~w8796;
assign w8798 = pi149 & pi261;
assign w8799 = w8797 & w8798;
assign w8800 = ~w8797 & ~w8798;
assign w8801 = ~w8799 & ~w8800;
assign w8802 = w8607 & w8801;
assign w8803 = ~w8607 & ~w8801;
assign w8804 = ~w8802 & ~w8803;
assign w8805 = w8602 & w8804;
assign w8806 = ~w8602 & ~w8804;
assign w8807 = ~w8805 & ~w8806;
assign w8808 = pi152 & pi258;
assign w8809 = ~w8362 & w8808;
assign w8810 = w8362 & ~w8808;
assign w8811 = ~w8809 & ~w8810;
assign w8812 = w8807 & w8811;
assign w8813 = ~w8807 & ~w8811;
assign w8814 = ~w8812 & ~w8813;
assign w8815 = pi322 & w8814;
assign w8816 = pi323 & ~w8367;
assign w8817 = ~w8371 & ~w8816;
assign w8818 = (~w7743 & w8370) | (~w7743 & w16201) | (w8370 & w16201);
assign w8819 = w8816 & ~w8818;
assign w8820 = ~w8817 & ~w8819;
assign w8821 = w8815 & w8820;
assign w8822 = ~w8815 & ~w8820;
assign w8823 = ~w8821 & ~w8822;
assign w8824 = w8597 & w8823;
assign w8825 = ~w8597 & ~w8823;
assign w8826 = ~w8824 & ~w8825;
assign w8827 = w8596 & ~w8826;
assign w8828 = ~w8596 & w8826;
assign w8829 = ~w8827 & ~w8828;
assign w8830 = (~w8585 & ~w8388) | (~w8585 & w16202) | (~w8388 & w16202);
assign w8831 = ~w8373 & ~w8378;
assign w8832 = ~w8377 & ~w8831;
assign w8833 = pi326 & w6283;
assign w8834 = pi325 & ~w7108;
assign w8835 = w8833 & ~w8834;
assign w8836 = ~w8833 & w8834;
assign w8837 = ~w8835 & ~w8836;
assign w8838 = w8832 & ~w8837;
assign w8839 = ~w8832 & w8837;
assign w8840 = ~w8838 & ~w8839;
assign w8841 = w8830 & ~w8840;
assign w8842 = ~w8830 & w8840;
assign w8843 = ~w8841 & ~w8842;
assign w8844 = w8829 & w8843;
assign w8845 = ~w8829 & ~w8843;
assign w8846 = ~w8844 & ~w8845;
assign w8847 = ~w8594 & w8846;
assign w8848 = w8594 & ~w8846;
assign w8849 = ~w8847 & ~w8848;
assign w8850 = (w8414 & ~w8410) | (w8414 & w16203) | (~w8410 & w16203);
assign w8851 = ~w8412 & ~w8850;
assign w8852 = pi328 & w5194;
assign w8853 = pi329 & ~w4854;
assign w8854 = pi327 & w5714;
assign w8855 = w8853 & ~w8854;
assign w8856 = ~w8853 & w8854;
assign w8857 = ~w8855 & ~w8856;
assign w8858 = w8852 & ~w8857;
assign w8859 = ~w8852 & w8857;
assign w8860 = ~w8858 & ~w8859;
assign w8861 = w8851 & ~w8860;
assign w8862 = ~w8851 & w8860;
assign w8863 = ~w8861 & ~w8862;
assign w8864 = w8849 & w8863;
assign w8865 = ~w8849 & ~w8863;
assign w8866 = ~w8864 & ~w8865;
assign w8867 = w8584 & w8866;
assign w8868 = ~w8584 & ~w8866;
assign w8869 = ~w8867 & ~w8868;
assign w8870 = w8582 & w8869;
assign w8871 = ~w8582 & ~w8869;
assign w8872 = ~w8870 & ~w8871;
assign w8873 = w8577 & ~w8872;
assign w8874 = ~w8577 & w8872;
assign w8875 = ~w8873 & ~w8874;
assign w8876 = pi332 & ~w3568;
assign w8877 = ~w8147 & ~w8443;
assign w8878 = ~w8876 & w8877;
assign w8879 = w8876 & ~w8877;
assign w8880 = ~w8878 & ~w8879;
assign w8881 = ~w8875 & w8880;
assign w8882 = w8875 & ~w8880;
assign w8883 = ~w8881 & ~w8882;
assign w8884 = ~w8572 & ~w8883;
assign w8885 = w8572 & w8883;
assign w8886 = ~w8884 & ~w8885;
assign w8887 = pi335 & ~w2373;
assign w8888 = ~w8566 & ~w8567;
assign w8889 = ~w8114 & w8117;
assign w8890 = pi334 & w2698;
assign w8891 = ~pi333 & w8890;
assign w8892 = ~pi334 & w8114;
assign w8893 = ~w8891 & ~w8892;
assign w8894 = ~w8116 & w8893;
assign w8895 = ~w8889 & w8894;
assign w8896 = ~w8116 & ~w8890;
assign w8897 = w2698 & ~w8117;
assign w8898 = ~w8896 & ~w8897;
assign w8899 = ~w8116 & w8891;
assign w8900 = ~w8888 & w8899;
assign w8901 = (~w8898 & ~w8888) | (~w8898 & w16204) | (~w8888 & w16204);
assign w8902 = ~w8900 & w8901;
assign w8903 = ~w8887 & w8902;
assign w8904 = w8887 & ~w8902;
assign w8905 = ~w8903 & ~w8904;
assign w8906 = w8886 & w8905;
assign w8907 = ~w8886 & ~w8905;
assign w8908 = ~w8906 & ~w8907;
assign w8909 = ~w8121 & w8888;
assign w8910 = w8121 & ~w8888;
assign w8911 = ~w8909 & ~w8910;
assign w8912 = ~w8446 & ~w8911;
assign w8913 = w8446 & w8911;
assign w8914 = ~w8122 & ~w8913;
assign w8915 = ~w8912 & ~w8914;
assign w8916 = w8908 & w8915;
assign w8917 = ~w8908 & ~w8915;
assign w8918 = ~w8916 & ~w8917;
assign w8919 = w8564 & w8918;
assign w8920 = ~w8564 & ~w8918;
assign w8921 = ~w8919 & ~w8920;
assign w8922 = ~w8559 & w8921;
assign w8923 = w8559 & ~w8921;
assign w8924 = ~w8922 & ~w8923;
assign w8925 = w8554 & ~w8924;
assign w8926 = ~w8554 & w8924;
assign w8927 = ~w8925 & ~w8926;
assign w8928 = pi339 & w1339;
assign w8929 = ~w8466 & ~w8469;
assign w8930 = w8928 & ~w8929;
assign w8931 = ~w8928 & w8929;
assign w8932 = ~w8930 & ~w8931;
assign w8933 = w8927 & w8932;
assign w8934 = ~w8927 & ~w8932;
assign w8935 = ~w8933 & ~w8934;
assign w8936 = w8549 & ~w8935;
assign w8937 = ~w8549 & w8935;
assign w8938 = ~w8936 & ~w8937;
assign w8939 = pi341 & ~w955;
assign w8940 = ~w8476 & ~w8480;
assign w8941 = ~w8939 & w8940;
assign w8942 = w8939 & ~w8940;
assign w8943 = ~w8941 & ~w8942;
assign w8944 = w8938 & w8943;
assign w8945 = ~w8938 & ~w8943;
assign w8946 = ~w8944 & ~w8945;
assign w8947 = w8544 & ~w8946;
assign w8948 = ~w8544 & w8946;
assign w8949 = ~w8947 & ~w8948;
assign w8950 = w8539 & w8949;
assign w8951 = ~w8539 & ~w8949;
assign w8952 = ~w8950 & ~w8951;
assign w8953 = w8534 & w8952;
assign w8954 = ~w8534 & ~w8952;
assign w8955 = ~w8953 & ~w8954;
assign w8956 = w8527 & w8955;
assign w8957 = ~w8527 & ~w8955;
assign w8958 = ~w8956 & ~w8957;
assign w8959 = ~w8523 & ~w8958;
assign w8960 = w8523 & w8958;
assign w8961 = ~w8959 & ~w8960;
assign w8962 = ~w8080 & ~w8504;
assign w8963 = ~w8961 & ~w8962;
assign w8964 = w8961 & w8962;
assign w8965 = ~w8963 & ~w8964;
assign w8966 = pi282 & w8965;
assign w8967 = ~pi282 & ~w8965;
assign w8968 = ~w8966 & ~w8967;
assign w8969 = ~w8508 & ~w8515;
assign w8970 = pi128 & pi297;
assign w8971 = pi298 & w464;
assign w8972 = ~w8074 & ~w8971;
assign w8973 = ~pi129 & w8074;
assign w8974 = ~w8972 & ~w8973;
assign w8975 = pi300 & w709;
assign w8976 = pi301 & w698;
assign w8977 = ~w8048 & ~w8058;
assign w8978 = pi302 & w855;
assign w8979 = pi304 & w1220;
assign w8980 = pi305 & w1420;
assign w8981 = ~w8032 & ~w8036;
assign w8982 = w8980 & ~w8981;
assign w8983 = ~w8980 & w8981;
assign w8984 = ~w8982 & ~w8983;
assign w8985 = pi306 & w1693;
assign w8986 = pi307 & w1954;
assign w8987 = pi308 & ~w2473;
assign w8988 = pi309 & w2801;
assign w8989 = ~w8012 & ~w8015;
assign w8990 = pi310 & w2925;
assign w8991 = pi311 & w3304;
assign w8992 = pi312 & w3710;
assign w8993 = pi314 & w4539;
assign w8994 = ~w7953 & ~w7956;
assign w8995 = pi315 & w5316;
assign w8996 = pi316 & w5862;
assign w8997 = pi317 & w6437;
assign w8998 = pi318 & w6652;
assign w8999 = pi319 & w7268;
assign w9000 = w7268 & w7913;
assign w9001 = ~w7909 & ~w9000;
assign w9002 = pi320 & ~w9001;
assign w9003 = w7268 & w7909;
assign w9004 = pi151 & ~pi152;
assign w9005 = ~pi151 & pi152;
assign w9006 = ~w9004 & ~w9005;
assign w9007 = ~pi151 & w7262;
assign w9008 = ~w7904 & ~w9007;
assign w9009 = w9006 & ~w9008;
assign w9010 = ~pi149 & ~w9009;
assign w9011 = ~w7262 & w9004;
assign w9012 = pi152 & w7903;
assign w9013 = pi149 & ~w9012;
assign w9014 = ~w9011 & w9013;
assign w9015 = ~w9010 & ~w9014;
assign w9016 = pi152 & ~w7262;
assign w9017 = ~pi150 & ~w9016;
assign w9018 = ~w9006 & ~w9007;
assign w9019 = ~w9017 & ~w9018;
assign w9020 = ~pi150 & ~w9006;
assign w9021 = ~w9019 & ~w9020;
assign w9022 = ~w9015 & ~w9021;
assign w9023 = ~w9001 & w9022;
assign w9024 = w7909 & w7913;
assign w9025 = ~w9003 & ~w9024;
assign w9026 = ~w9023 & w9025;
assign w9027 = pi321 & ~w9026;
assign w9028 = w9002 & ~w9027;
assign w9029 = ~pi320 & ~w9022;
assign w9030 = pi320 & w9022;
assign w9031 = ~w9029 & ~w9030;
assign w9032 = w9024 & w9031;
assign w9033 = w9002 & ~w9003;
assign w9034 = w9022 & ~w9033;
assign w9035 = ~w9024 & ~w9034;
assign w9036 = pi321 & ~w9032;
assign w9037 = ~w9035 & w9036;
assign w9038 = ~w9028 & ~w9037;
assign w9039 = w8999 & ~w9038;
assign w9040 = ~w8999 & w9038;
assign w9041 = ~w9039 & ~w9040;
assign w9042 = ~w7921 & ~w7924;
assign w9043 = w9041 & w9042;
assign w9044 = ~w9041 & ~w9042;
assign w9045 = ~w9043 & ~w9044;
assign w9046 = ~w8998 & ~w9045;
assign w9047 = w8998 & w9045;
assign w9048 = ~w9046 & ~w9047;
assign w9049 = ~w7928 & ~w7931;
assign w9050 = w9048 & ~w9049;
assign w9051 = ~w9048 & w9049;
assign w9052 = ~w9050 & ~w9051;
assign w9053 = ~w8997 & ~w9052;
assign w9054 = w8997 & w9052;
assign w9055 = ~w9053 & ~w9054;
assign w9056 = ~w7935 & ~w7938;
assign w9057 = w9055 & ~w9056;
assign w9058 = ~w9055 & w9056;
assign w9059 = ~w9057 & ~w9058;
assign w9060 = w8996 & ~w9059;
assign w9061 = ~w8996 & w9059;
assign w9062 = ~w9060 & ~w9061;
assign w9063 = w7899 & ~w7947;
assign w9064 = ~w7946 & ~w9063;
assign w9065 = ~w9062 & w9064;
assign w9066 = w9062 & ~w9064;
assign w9067 = ~w9065 & ~w9066;
assign w9068 = ~w8995 & ~w9067;
assign w9069 = w8995 & w9067;
assign w9070 = ~w9068 & ~w9069;
assign w9071 = w8994 & w9070;
assign w9072 = ~w8994 & ~w9070;
assign w9073 = ~w9071 & ~w9072;
assign w9074 = w8993 & w9073;
assign w9075 = ~w8993 & ~w9073;
assign w9076 = ~w9074 & ~w9075;
assign w9077 = ~w7960 & ~w7963;
assign w9078 = w9076 & w9077;
assign w9079 = ~w9076 & ~w9077;
assign w9080 = ~w9078 & ~w9079;
assign w9081 = pi313 & w4382;
assign w9082 = ~w7968 & ~w7972;
assign w9083 = w9081 & w9082;
assign w9084 = ~w9081 & ~w9082;
assign w9085 = ~w9083 & ~w9084;
assign w9086 = w9080 & w9085;
assign w9087 = ~w9080 & ~w9085;
assign w9088 = ~w9086 & ~w9087;
assign w9089 = ~w8992 & ~w9088;
assign w9090 = w8992 & w9088;
assign w9091 = ~w9089 & ~w9090;
assign w9092 = ~w7975 & ~w7977;
assign w9093 = ~w9091 & ~w9092;
assign w9094 = w9091 & w9092;
assign w9095 = ~w9093 & ~w9094;
assign w9096 = ~w7980 & ~w7984;
assign w9097 = w9095 & w9096;
assign w9098 = ~w9095 & ~w9096;
assign w9099 = ~w9097 & ~w9098;
assign w9100 = w8991 & w9099;
assign w9101 = ~w8991 & ~w9099;
assign w9102 = ~w9100 & ~w9101;
assign w9103 = w8006 & ~w9102;
assign w9104 = ~w8006 & w9102;
assign w9105 = ~w9103 & ~w9104;
assign w9106 = w8990 & ~w9105;
assign w9107 = ~w8990 & ~w9104;
assign w9108 = ~w9103 & w9107;
assign w9109 = ~w9106 & ~w9108;
assign w9110 = w8989 & w9109;
assign w9111 = ~w8989 & ~w9109;
assign w9112 = ~w9110 & ~w9111;
assign w9113 = w8988 & ~w9112;
assign w9114 = ~w8988 & w9112;
assign w9115 = ~w9113 & ~w9114;
assign w9116 = w8987 & ~w9115;
assign w9117 = ~w8987 & w9115;
assign w9118 = ~w9116 & ~w9117;
assign w9119 = ~w7891 & ~w8019;
assign w9120 = w9118 & w9119;
assign w9121 = ~w9118 & ~w9119;
assign w9122 = ~w9120 & ~w9121;
assign w9123 = ~w8021 & ~w8025;
assign w9124 = w9122 & ~w9123;
assign w9125 = ~w9122 & w9123;
assign w9126 = ~w9124 & ~w9125;
assign w9127 = w8986 & w9126;
assign w9128 = ~w8986 & ~w9126;
assign w9129 = ~w9127 & ~w9128;
assign w9130 = ~w7885 & ~w8028;
assign w9131 = w9129 & ~w9130;
assign w9132 = ~w9129 & w9130;
assign w9133 = ~w9131 & ~w9132;
assign w9134 = w8985 & w9133;
assign w9135 = ~w8985 & ~w9133;
assign w9136 = ~w9134 & ~w9135;
assign w9137 = w8984 & w9136;
assign w9138 = ~w8984 & ~w9136;
assign w9139 = ~w9137 & ~w9138;
assign w9140 = w8979 & w9139;
assign w9141 = ~w8979 & ~w9139;
assign w9142 = ~w9140 & ~w9141;
assign w9143 = ~w7880 & ~w8039;
assign w9144 = w9142 & ~w9143;
assign w9145 = ~w9142 & w9143;
assign w9146 = ~w9144 & ~w9145;
assign w9147 = ~w7875 & ~w8043;
assign w9148 = ~w9146 & w9147;
assign w9149 = w9146 & ~w9147;
assign w9150 = ~w9148 & ~w9149;
assign w9151 = pi303 & w1159;
assign w9152 = w9150 & w9151;
assign w9153 = ~w9150 & ~w9151;
assign w9154 = ~w9152 & ~w9153;
assign w9155 = ~w7870 & ~w8045;
assign w9156 = w9154 & ~w9155;
assign w9157 = ~w9154 & w9155;
assign w9158 = ~w9156 & ~w9157;
assign w9159 = w8978 & ~w9158;
assign w9160 = ~w8978 & w9158;
assign w9161 = ~w9159 & ~w9160;
assign w9162 = w8977 & w9161;
assign w9163 = ~w8977 & ~w9161;
assign w9164 = ~w9162 & ~w9163;
assign w9165 = w8976 & w9164;
assign w9166 = ~w8976 & ~w9164;
assign w9167 = ~w9165 & ~w9166;
assign w9168 = w8975 & w9167;
assign w9169 = ~w8975 & ~w9167;
assign w9170 = ~w9168 & ~w9169;
assign w9171 = ~w8065 & ~w8068;
assign w9172 = w9170 & w9171;
assign w9173 = ~w9170 & ~w9171;
assign w9174 = ~w9172 & ~w9173;
assign w9175 = pi299 & ~w653;
assign w9176 = ~w7861 & ~w8071;
assign w9177 = w9175 & ~w9176;
assign w9178 = ~w9175 & w9176;
assign w9179 = ~w9177 & ~w9178;
assign w9180 = w9174 & ~w9179;
assign w9181 = ~w9174 & w9179;
assign w9182 = ~w9180 & ~w9181;
assign w9183 = w8974 & w9182;
assign w9184 = ~w8974 & ~w9182;
assign w9185 = ~w9183 & ~w9184;
assign w9186 = w8970 & ~w9185;
assign w9187 = ~w8970 & w9185;
assign w9188 = ~w9186 & ~w9187;
assign w9189 = w8969 & ~w9188;
assign w9190 = ~w8969 & w9188;
assign w9191 = ~w9189 & ~w9190;
assign w9192 = ~w8968 & ~w9191;
assign w9193 = w8968 & w9191;
assign w9194 = ~w135 & ~w9192;
assign w9195 = ~w9193 & w9194;
assign w9196 = pi161 & ~w193;
assign w9197 = ~w9195 & w9196;
assign w9198 = ~pi160 & ~w8522;
assign w9199 = ~w9197 & w9198;
assign w9200 = ~pi089 & ~pi161;
assign w9201 = pi283 & w135;
assign w9202 = ~w9190 & ~w9193;
assign w9203 = pi128 & pi296;
assign w9204 = pi129 & ~pi297;
assign w9205 = ~w9186 & ~w9204;
assign w9206 = pi298 & ~w653;
assign w9207 = ~w8973 & ~w9183;
assign w9208 = w9206 & ~w9207;
assign w9209 = ~w9206 & w9207;
assign w9210 = ~w9208 & ~w9209;
assign w9211 = pi299 & w709;
assign w9212 = ~w9177 & ~w9181;
assign w9213 = w9211 & ~w9212;
assign w9214 = ~w9211 & w9212;
assign w9215 = ~w9213 & ~w9214;
assign w9216 = ~w9169 & ~w9172;
assign w9217 = pi300 & w698;
assign w9218 = w9216 & w9217;
assign w9219 = ~w9216 & ~w9217;
assign w9220 = ~w9218 & ~w9219;
assign w9221 = pi301 & w855;
assign w9222 = pi303 & w1220;
assign w9223 = ~w9140 & ~w9144;
assign w9224 = pi304 & w1420;
assign w9225 = ~w9223 & w9224;
assign w9226 = w9223 & ~w9224;
assign w9227 = ~w9225 & ~w9226;
assign w9228 = pi305 & w1693;
assign w9229 = pi307 & ~w2473;
assign w9230 = pi308 & w2801;
assign w9231 = ~w9116 & ~w9120;
assign w9232 = w9230 & ~w9231;
assign w9233 = ~w9230 & w9231;
assign w9234 = ~w9232 & ~w9233;
assign w9235 = pi309 & w2925;
assign w9236 = pi310 & w3304;
assign w9237 = pi311 & w3710;
assign w9238 = ~w9089 & ~w9094;
assign w9239 = pi312 & w4382;
assign w9240 = pi313 & w4539;
assign w9241 = pi314 & w5316;
assign w9242 = pi315 & w5862;
assign w9243 = pi316 & w6437;
assign w9244 = pi317 & w6652;
assign w9245 = pi318 & w7268;
assign w9246 = pi319 & w7909;
assign w9247 = ~pi153 & w9006;
assign w9248 = pi152 & pi153;
assign w9249 = pi151 & pi153;
assign w9250 = ~w9016 & ~w9249;
assign w9251 = pi150 & ~w9250;
assign w9252 = ~w9248 & w9251;
assign w9253 = pi153 & w9005;
assign w9254 = ~pi152 & ~pi153;
assign w9255 = w7262 & w9254;
assign w9256 = ~w9253 & ~w9255;
assign w9257 = ~pi150 & ~w9256;
assign w9258 = ~pi150 & w9254;
assign w9259 = w9007 & w9248;
assign w9260 = ~w9258 & ~w9259;
assign w9261 = ~pi149 & ~w9260;
assign w9262 = pi150 & pi152;
assign w9263 = ~pi153 & ~w9262;
assign w9264 = pi153 & ~w9011;
assign w9265 = pi149 & ~w9263;
assign w9266 = ~w9264 & w9265;
assign w9267 = ~w9247 & ~w9257;
assign w9268 = ~w9266 & w9267;
assign w9269 = ~w9252 & ~w9261;
assign w9270 = w9268 & w9269;
assign w9271 = pi321 & w9270;
assign w9272 = pi320 & w9027;
assign w9273 = ~w9271 & ~w9272;
assign w9274 = w9270 & w9272;
assign w9275 = ~w9273 & ~w9274;
assign w9276 = w9030 & w9275;
assign w9277 = ~w9030 & ~w9275;
assign w9278 = ~w9276 & ~w9277;
assign w9279 = ~w9039 & ~w9043;
assign w9280 = w9278 & ~w9279;
assign w9281 = ~w9278 & w9279;
assign w9282 = ~w9280 & ~w9281;
assign w9283 = w9246 & ~w9282;
assign w9284 = ~w9246 & w9282;
assign w9285 = ~w9283 & ~w9284;
assign w9286 = w9245 & ~w9285;
assign w9287 = ~w9245 & w9285;
assign w9288 = ~w9286 & ~w9287;
assign w9289 = ~w9047 & ~w9050;
assign w9290 = w9288 & ~w9289;
assign w9291 = ~w9288 & w9289;
assign w9292 = ~w9290 & ~w9291;
assign w9293 = w9244 & w9292;
assign w9294 = ~w9244 & ~w9292;
assign w9295 = ~w9293 & ~w9294;
assign w9296 = ~w9053 & ~w9057;
assign w9297 = w9295 & ~w9296;
assign w9298 = ~w9295 & w9296;
assign w9299 = ~w9297 & ~w9298;
assign w9300 = ~w9060 & ~w9066;
assign w9301 = ~w9299 & ~w9300;
assign w9302 = w9299 & w9300;
assign w9303 = ~w9301 & ~w9302;
assign w9304 = ~w9243 & w9303;
assign w9305 = w9243 & ~w9303;
assign w9306 = ~w9304 & ~w9305;
assign w9307 = w9242 & ~w9306;
assign w9308 = ~w9242 & w9306;
assign w9309 = ~w9307 & ~w9308;
assign w9310 = ~w9069 & ~w9071;
assign w9311 = ~w9309 & w9310;
assign w9312 = w9309 & ~w9310;
assign w9313 = ~w9311 & ~w9312;
assign w9314 = w9241 & w9313;
assign w9315 = ~w9241 & ~w9313;
assign w9316 = ~w9314 & ~w9315;
assign w9317 = ~w9074 & ~w9078;
assign w9318 = w9316 & w9317;
assign w9319 = ~w9316 & ~w9317;
assign w9320 = ~w9318 & ~w9319;
assign w9321 = ~w9240 & w9320;
assign w9322 = w9240 & ~w9320;
assign w9323 = ~w9321 & ~w9322;
assign w9324 = ~w9083 & ~w9086;
assign w9325 = w9323 & ~w9324;
assign w9326 = ~w9323 & w9324;
assign w9327 = ~w9325 & ~w9326;
assign w9328 = w9239 & w9327;
assign w9329 = ~w9239 & ~w9327;
assign w9330 = ~w9328 & ~w9329;
assign w9331 = w9238 & ~w9330;
assign w9332 = ~w9238 & w9330;
assign w9333 = ~w9331 & ~w9332;
assign w9334 = ~w9237 & w9333;
assign w9335 = w9237 & ~w9333;
assign w9336 = ~w9334 & ~w9335;
assign w9337 = ~w9098 & ~w9100;
assign w9338 = w9336 & w9337;
assign w9339 = ~w9336 & ~w9337;
assign w9340 = ~w9338 & ~w9339;
assign w9341 = ~w9103 & w9340;
assign w9342 = w9103 & ~w9340;
assign w9343 = ~w9341 & ~w9342;
assign w9344 = ~w9105 & w9236;
assign w9345 = w9343 & w9344;
assign w9346 = w2925 & w3304;
assign w9347 = w9105 & w9346;
assign w9348 = ~w9340 & w9347;
assign w9349 = w9236 & ~w9340;
assign w9350 = ~w9236 & w9340;
assign w9351 = w9107 & ~w9349;
assign w9352 = ~w9350 & w9351;
assign w9353 = ~w3304 & ~w9108;
assign w9354 = ~w9343 & w9353;
assign w9355 = ~w9345 & ~w9348;
assign w9356 = ~w9352 & ~w9354;
assign w9357 = w9355 & w9356;
assign w9358 = ~w9235 & w9357;
assign w9359 = w9235 & ~w9357;
assign w9360 = ~w9358 & ~w9359;
assign w9361 = ~w9110 & ~w9114;
assign w9362 = ~w9360 & ~w9361;
assign w9363 = w9360 & w9361;
assign w9364 = ~w9362 & ~w9363;
assign w9365 = w9234 & ~w9364;
assign w9366 = ~w9234 & w9364;
assign w9367 = ~w9365 & ~w9366;
assign w9368 = w9229 & ~w9367;
assign w9369 = ~w9229 & w9367;
assign w9370 = ~w9368 & ~w9369;
assign w9371 = ~w9124 & ~w9127;
assign w9372 = w9370 & ~w9371;
assign w9373 = ~w9370 & w9371;
assign w9374 = ~w9372 & ~w9373;
assign w9375 = ~w9131 & ~w9374;
assign w9376 = w1693 & ~w9132;
assign w9377 = w9375 & ~w9376;
assign w9378 = w1954 & ~w9377;
assign w9379 = ~w9132 & w9374;
assign w9380 = pi306 & ~w9379;
assign w9381 = ~w9375 & ~w9380;
assign w9382 = w9378 & ~w9381;
assign w9383 = w9132 & ~w9374;
assign w9384 = ~w8985 & ~w9131;
assign w9385 = w9379 & ~w9384;
assign w9386 = ~w9383 & ~w9385;
assign w9387 = ~w1954 & ~w9386;
assign w9388 = pi306 & w1954;
assign w9389 = ~w9374 & w9388;
assign w9390 = w9374 & ~w9388;
assign w9391 = w9384 & ~w9389;
assign w9392 = ~w9390 & w9391;
assign w9393 = ~w9382 & ~w9392;
assign w9394 = ~w9387 & w9393;
assign w9395 = ~w9228 & ~w9394;
assign w9396 = w9228 & w9394;
assign w9397 = ~w9395 & ~w9396;
assign w9398 = ~w8982 & ~w9137;
assign w9399 = w9397 & w9398;
assign w9400 = ~w9397 & ~w9398;
assign w9401 = ~w9399 & ~w9400;
assign w9402 = w9227 & ~w9401;
assign w9403 = ~w9227 & w9401;
assign w9404 = ~w9402 & ~w9403;
assign w9405 = ~w9222 & ~w9404;
assign w9406 = w9222 & w9404;
assign w9407 = ~w9405 & ~w9406;
assign w9408 = ~w9149 & ~w9152;
assign w9409 = w9407 & w9408;
assign w9410 = ~w9407 & ~w9408;
assign w9411 = ~w9409 & ~w9410;
assign w9412 = ~w9157 & ~w9411;
assign w9413 = pi302 & w1159;
assign w9414 = ~w9156 & w9411;
assign w9415 = w9413 & ~w9414;
assign w9416 = ~w9412 & w9415;
assign w9417 = w9157 & w9411;
assign w9418 = ~w9412 & ~w9417;
assign w9419 = ~w1159 & ~w9160;
assign w9420 = ~w9418 & w9419;
assign w9421 = ~w9411 & w9413;
assign w9422 = w9411 & ~w9413;
assign w9423 = ~w9421 & ~w9422;
assign w9424 = ~w8978 & ~w9156;
assign w9425 = ~w9423 & w9424;
assign w9426 = w1213 & ~w9157;
assign w9427 = w9414 & w9426;
assign w9428 = ~w9416 & ~w9427;
assign w9429 = ~w9420 & ~w9425;
assign w9430 = w9428 & w9429;
assign w9431 = ~w9221 & ~w9430;
assign w9432 = w9221 & w9430;
assign w9433 = ~w9431 & ~w9432;
assign w9434 = ~w9163 & ~w9165;
assign w9435 = ~w9433 & w9434;
assign w9436 = w9433 & ~w9434;
assign w9437 = ~w9435 & ~w9436;
assign w9438 = ~w9220 & ~w9437;
assign w9439 = w9220 & w9437;
assign w9440 = ~w9438 & ~w9439;
assign w9441 = w9215 & w9440;
assign w9442 = ~w9215 & ~w9440;
assign w9443 = ~w9441 & ~w9442;
assign w9444 = w9210 & w9443;
assign w9445 = ~w9210 & ~w9443;
assign w9446 = ~w9444 & ~w9445;
assign w9447 = pi129 & ~w9446;
assign w9448 = ~pi129 & w9446;
assign w9449 = ~w9447 & ~w9448;
assign w9450 = w9205 & w9449;
assign w9451 = ~w9205 & ~w9449;
assign w9452 = ~w9450 & ~w9451;
assign w9453 = w9203 & w9452;
assign w9454 = ~w9203 & ~w9452;
assign w9455 = ~w9453 & ~w9454;
assign w9456 = pi347 & w456;
assign w9457 = pi345 & ~w537;
assign w9458 = ~w8524 & ~w8956;
assign w9459 = ~w9457 & w9458;
assign w9460 = w9457 & ~w9458;
assign w9461 = ~w9459 & ~w9460;
assign w9462 = pi344 & ~w615;
assign w9463 = ~w8531 & ~w8953;
assign w9464 = w9462 & ~w9463;
assign w9465 = ~w9462 & w9463;
assign w9466 = ~w9464 & ~w9465;
assign w9467 = pi343 & ~w793;
assign w9468 = ~w8538 & ~w8950;
assign w9469 = ~w9467 & w9468;
assign w9470 = w9467 & ~w9468;
assign w9471 = ~w9469 & ~w9470;
assign w9472 = pi342 & ~w955;
assign w9473 = ~w8542 & ~w8947;
assign w9474 = w9472 & ~w9473;
assign w9475 = ~w9472 & w9473;
assign w9476 = ~w9474 & ~w9475;
assign w9477 = pi340 & w1339;
assign w9478 = ~w8547 & ~w8936;
assign w9479 = w9477 & w9478;
assign w9480 = ~w9477 & ~w9478;
assign w9481 = ~w9479 & ~w9480;
assign w9482 = pi339 & w1602;
assign w9483 = ~w8930 & ~w8933;
assign w9484 = w9482 & ~w9483;
assign w9485 = ~w9482 & w9483;
assign w9486 = ~w9484 & ~w9485;
assign w9487 = pi337 & ~w2170;
assign w9488 = ~w8557 & ~w8921;
assign w9489 = ~w8558 & ~w9488;
assign w9490 = ~w9487 & ~w9489;
assign w9491 = w9487 & w9489;
assign w9492 = ~w9490 & ~w9491;
assign w9493 = pi336 & ~w2373;
assign w9494 = (~w8563 & ~w8918) | (~w8563 & w16205) | (~w8918 & w16205);
assign w9495 = ~w9493 & w9494;
assign w9496 = w9493 & ~w9494;
assign w9497 = ~w9495 & ~w9496;
assign w9498 = w8887 & ~w8908;
assign w9499 = ~w8916 & ~w9498;
assign w9500 = pi335 & w2698;
assign w9501 = w9499 & ~w9500;
assign w9502 = ~w9499 & w9500;
assign w9503 = ~w9501 & ~w9502;
assign w9504 = pi334 & ~w3183;
assign w9505 = ~w8886 & ~w8890;
assign w9506 = ~w8116 & w8911;
assign w9507 = ~w8117 & ~w9506;
assign w9508 = (~w9507 & ~w8886) | (~w9507 & w16460) | (~w8886 & w16460);
assign w9509 = ~w9505 & ~w9508;
assign w9510 = w9504 & w9509;
assign w9511 = ~w9504 & ~w9509;
assign w9512 = ~w9510 & ~w9511;
assign w9513 = pi333 & ~w3568;
assign w9514 = ~w8570 & ~w8885;
assign w9515 = ~w9513 & w9514;
assign w9516 = w9513 & ~w9514;
assign w9517 = ~w9515 & ~w9516;
assign w9518 = w8875 & w8877;
assign w9519 = ~w3568 & w3979;
assign w9520 = ~w8875 & ~w8877;
assign w9521 = ~w9519 & ~w9520;
assign w9522 = pi332 & w3979;
assign w9523 = ~w9518 & w9522;
assign w9524 = ~w9521 & w9523;
assign w9525 = w8876 & ~w9518;
assign w9526 = ~w9520 & ~w9522;
assign w9527 = ~w9525 & w9526;
assign w9528 = ~w9524 & ~w9527;
assign w9529 = pi329 & w5194;
assign w9530 = w8853 & ~w8866;
assign w9531 = ~w8867 & ~w9530;
assign w9532 = w8849 & w8854;
assign w9533 = ~w8847 & ~w9532;
assign w9534 = ~w8851 & w8852;
assign w9535 = w8851 & ~w8852;
assign w9536 = ~w8849 & ~w8854;
assign w9537 = (~w9535 & ~w8849) | (~w9535 & w16206) | (~w8849 & w16206);
assign w9538 = ~w9536 & w9537;
assign w9539 = ~w9534 & ~w9538;
assign w9540 = ~w9533 & w9539;
assign w9541 = w9533 & ~w9539;
assign w9542 = ~w9540 & ~w9541;
assign w9543 = pi324 & ~w8367;
assign w9544 = pi323 & w8814;
assign w9545 = ~w8163 & ~w8364;
assign w9546 = pi258 & w8361;
assign w9547 = ~pi259 & ~w9546;
assign w9548 = pi151 & ~w9547;
assign w9549 = w458 & w8361;
assign w9550 = w9548 & ~w9549;
assign w9551 = w8804 & ~w9550;
assign w9552 = ~w8804 & w9550;
assign w9553 = ~w9551 & ~w9552;
assign w9554 = ~w8808 & w9553;
assign w9555 = w8808 & ~w9553;
assign w9556 = ~w9554 & ~w9555;
assign w9557 = ~w9545 & w9556;
assign w9558 = ~w8599 & ~w9557;
assign w9559 = pi151 & pi260;
assign w9560 = ~w9559 & w17696;
assign w9561 = pi260 & ~w9547;
assign w9562 = (w9561 & w8804) | (w9561 & w16207) | (w8804 & w16207);
assign w9563 = ~w9560 & ~w9562;
assign w9564 = (~w8605 & ~w8801) | (~w8605 & w15941) | (~w8801 & w15941);
assign w9565 = ~w8613 & w8623;
assign w9566 = ~w8786 & ~w9565;
assign w9567 = (~w8777 & ~w8779) | (~w8777 & w17612) | (~w8779 & w17612);
assign w9568 = pi146 & pi265;
assign w9569 = ~w8755 & ~w8758;
assign w9570 = ~w8754 & ~w9569;
assign w9571 = w8742 & w8750;
assign w9572 = ~w8751 & ~w9571;
assign w9573 = pi143 & pi268;
assign w9574 = pi140 & pi271;
assign w9575 = w8639 & ~w8723;
assign w9576 = ~w8722 & ~w9575;
assign w9577 = ~w8645 & w8718;
assign w9578 = ~w8644 & ~w9577;
assign w9579 = pi137 & pi274;
assign w9580 = pi136 & pi275;
assign w9581 = pi135 & pi276;
assign w9582 = pi134 & pi277;
assign w9583 = pi133 & pi278;
assign w9584 = ~w8688 & ~w8691;
assign w9585 = pi132 & pi279;
assign w9586 = pi131 & pi280;
assign w9587 = ~w8670 & ~w8673;
assign w9588 = pi129 & pi282;
assign w9589 = pi128 & pi283;
assign w9590 = ~w9588 & ~w9589;
assign w9591 = pi129 & pi283;
assign w9592 = w8661 & w9591;
assign w9593 = ~w9590 & ~w9592;
assign w9594 = ~pi281 & w8663;
assign w9595 = pi130 & pi281;
assign w9596 = pi129 & ~w8664;
assign w9597 = w9595 & ~w9596;
assign w9598 = ~w9594 & ~w9597;
assign w9599 = ~w9593 & ~w9598;
assign w9600 = ~w8201 & ~w8663;
assign w9601 = w9593 & ~w9595;
assign w9602 = w9600 & w9601;
assign w9603 = ~w8664 & w9593;
assign w9604 = w646 & ~w9594;
assign w9605 = w9603 & w9604;
assign w9606 = ~w8664 & ~w9600;
assign w9607 = ~w9593 & ~w9606;
assign w9608 = ~pi130 & ~w9603;
assign w9609 = ~w9607 & w9608;
assign w9610 = ~w9602 & ~w9605;
assign w9611 = ~w9599 & w9610;
assign w9612 = ~w9609 & w9611;
assign w9613 = w9587 & ~w9612;
assign w9614 = ~w9587 & w9612;
assign w9615 = ~w9613 & ~w9614;
assign w9616 = w9586 & w9615;
assign w9617 = ~w9586 & ~w9615;
assign w9618 = ~w9616 & ~w9617;
assign w9619 = ~w8676 & ~w8680;
assign w9620 = w9618 & w9619;
assign w9621 = ~w9618 & ~w9619;
assign w9622 = ~w9620 & ~w9621;
assign w9623 = w9585 & ~w9622;
assign w9624 = ~w9585 & w9622;
assign w9625 = ~w9623 & ~w9624;
assign w9626 = ~w8657 & ~w8683;
assign w9627 = ~w9625 & w9626;
assign w9628 = w9625 & ~w9626;
assign w9629 = ~w9627 & ~w9628;
assign w9630 = ~w9584 & ~w9629;
assign w9631 = w9584 & w9629;
assign w9632 = ~w9630 & ~w9631;
assign w9633 = w9583 & w9632;
assign w9634 = ~w9583 & ~w9632;
assign w9635 = ~w9633 & ~w9634;
assign w9636 = ~w9582 & ~w9635;
assign w9637 = w9582 & w9635;
assign w9638 = ~w9636 & ~w9637;
assign w9639 = ~w8694 & ~w8697;
assign w9640 = ~w9638 & w9639;
assign w9641 = w9638 & ~w9639;
assign w9642 = ~w9640 & ~w9641;
assign w9643 = ~w8701 & ~w8705;
assign w9644 = w9642 & w9643;
assign w9645 = ~w9642 & ~w9643;
assign w9646 = ~w9644 & ~w9645;
assign w9647 = w9581 & w9646;
assign w9648 = ~w9581 & ~w9646;
assign w9649 = ~w9647 & ~w9648;
assign w9650 = ~w9580 & ~w9649;
assign w9651 = w9580 & w9649;
assign w9652 = ~w9650 & ~w9651;
assign w9653 = w8649 & ~w8707;
assign w9654 = ~w8708 & ~w9653;
assign w9655 = w9652 & ~w9654;
assign w9656 = ~w9652 & w9654;
assign w9657 = ~w9655 & ~w9656;
assign w9658 = w9579 & w9657;
assign w9659 = ~w9579 & ~w9657;
assign w9660 = ~w9658 & ~w9659;
assign w9661 = w8647 & ~w8714;
assign w9662 = ~w8713 & ~w9661;
assign w9663 = w9660 & w9662;
assign w9664 = ~w9660 & ~w9662;
assign w9665 = ~w9663 & ~w9664;
assign w9666 = ~w9578 & w9665;
assign w9667 = w9578 & ~w9665;
assign w9668 = ~w9666 & ~w9667;
assign w9669 = pi139 & pi272;
assign w9670 = pi138 & pi273;
assign w9671 = w9669 & ~w9670;
assign w9672 = ~w9669 & w9670;
assign w9673 = ~w9671 & ~w9672;
assign w9674 = w9668 & w9673;
assign w9675 = ~w9668 & ~w9673;
assign w9676 = ~w9674 & ~w9675;
assign w9677 = ~w9576 & w9676;
assign w9678 = w9576 & ~w9676;
assign w9679 = ~w9677 & ~w9678;
assign w9680 = ~w9574 & ~w9679;
assign w9681 = w9574 & w9679;
assign w9682 = ~w9680 & ~w9681;
assign w9683 = ~w8636 & ~w8729;
assign w9684 = ~w9682 & w9683;
assign w9685 = w9682 & ~w9683;
assign w9686 = ~w9684 & ~w9685;
assign w9687 = ~w8731 & ~w8735;
assign w9688 = ~w8732 & ~w9687;
assign w9689 = ~w9686 & w9688;
assign w9690 = w9686 & ~w9688;
assign w9691 = ~w9689 & ~w9690;
assign w9692 = pi142 & pi269;
assign w9693 = pi141 & pi270;
assign w9694 = w9692 & ~w9693;
assign w9695 = ~w9692 & w9693;
assign w9696 = ~w9694 & ~w9695;
assign w9697 = w9691 & w9696;
assign w9698 = ~w9691 & ~w9696;
assign w9699 = ~w9697 & ~w9698;
assign w9700 = ~w8740 & w8744;
assign w9701 = ~w8739 & ~w9700;
assign w9702 = ~w9699 & w9701;
assign w9703 = w9699 & ~w9701;
assign w9704 = ~w9702 & ~w9703;
assign w9705 = ~w9573 & ~w9704;
assign w9706 = w9573 & w9704;
assign w9707 = ~w9705 & ~w9706;
assign w9708 = w9572 & ~w9707;
assign w9709 = ~w9572 & w9707;
assign w9710 = ~w9708 & ~w9709;
assign w9711 = w9570 & ~w9710;
assign w9712 = ~w9570 & w9710;
assign w9713 = ~w9711 & ~w9712;
assign w9714 = pi145 & pi266;
assign w9715 = pi144 & pi267;
assign w9716 = w9714 & ~w9715;
assign w9717 = ~w9714 & w9715;
assign w9718 = ~w9716 & ~w9717;
assign w9719 = w9713 & w9718;
assign w9720 = ~w9713 & ~w9718;
assign w9721 = ~w9719 & ~w9720;
assign w9722 = ~w8762 & ~w8767;
assign w9723 = ~w8763 & ~w9722;
assign w9724 = w9721 & ~w9723;
assign w9725 = ~w9721 & w9723;
assign w9726 = ~w9724 & ~w9725;
assign w9727 = w9568 & ~w9726;
assign w9728 = ~w9568 & w9726;
assign w9729 = ~w9727 & ~w9728;
assign w9730 = ~w8765 & w8773;
assign w9731 = ~w8774 & ~w9730;
assign w9732 = w9729 & w9731;
assign w9733 = ~w9729 & ~w9731;
assign w9734 = ~w9732 & ~w9733;
assign w9735 = w9567 & ~w9734;
assign w9736 = ~w9567 & w9734;
assign w9737 = ~w9735 & ~w9736;
assign w9738 = pi148 & pi263;
assign w9739 = pi147 & pi264;
assign w9740 = w9738 & ~w9739;
assign w9741 = ~w9738 & w9739;
assign w9742 = ~w9740 & ~w9741;
assign w9743 = w9737 & w9742;
assign w9744 = ~w9737 & ~w9742;
assign w9745 = ~w9743 & ~w9744;
assign w9746 = w9566 & ~w9745;
assign w9747 = ~w9566 & w9745;
assign w9748 = ~w9746 & ~w9747;
assign w9749 = (~pi261 & w8787) | (~pi261 & w15942) | (w8787 & w15942);
assign w9750 = pi149 & pi262;
assign w9751 = (w9750 & ~w8787) | (w9750 & w15943) | (~w8787 & w15943);
assign w9752 = ~w9749 & w9751;
assign w9753 = w8787 & w15944;
assign w9754 = pi149 & ~w925;
assign w9755 = (~w9754 & w8787) | (~w9754 & w15945) | (w8787 & w15945);
assign w9756 = ~w9753 & ~w9755;
assign w9757 = ~w9752 & w9756;
assign w9758 = w9748 & w9757;
assign w9759 = ~w9748 & ~w9757;
assign w9760 = ~w9758 & ~w9759;
assign w9761 = w9564 & ~w9760;
assign w9762 = ~w9564 & w9760;
assign w9763 = ~w9761 & ~w9762;
assign w9764 = pi150 & pi261;
assign w9765 = ~w9763 & w9764;
assign w9766 = w9763 & ~w9764;
assign w9767 = ~w9765 & ~w9766;
assign w9768 = w9563 & ~w9767;
assign w9769 = ~w9563 & w9767;
assign w9770 = ~w9768 & ~w9769;
assign w9771 = pi153 & pi258;
assign w9772 = pi152 & pi259;
assign w9773 = w9771 & ~w9772;
assign w9774 = ~w9771 & w9772;
assign w9775 = ~w9773 & ~w9774;
assign w9776 = (w9775 & ~w9553) | (w9775 & w16208) | (~w9553 & w16208);
assign w9777 = w9553 & w16209;
assign w9778 = ~w9776 & ~w9777;
assign w9779 = w9770 & w9778;
assign w9780 = ~w9770 & ~w9778;
assign w9781 = ~w9779 & ~w9780;
assign w9782 = w9558 & ~w9781;
assign w9783 = ~w9558 & w9781;
assign w9784 = ~w9782 & ~w9783;
assign w9785 = ~w8819 & ~w8821;
assign w9786 = ~w9784 & w16210;
assign w9787 = (w9785 & w9784) | (w9785 & w16211) | (w9784 & w16211);
assign w9788 = ~w9786 & ~w9787;
assign w9789 = w9544 & w9788;
assign w9790 = ~w9544 & ~w9788;
assign w9791 = ~w9789 & ~w9790;
assign w9792 = w9543 & w9791;
assign w9793 = ~w9543 & ~w9791;
assign w9794 = ~w9792 & ~w9793;
assign w9795 = w8826 & w8832;
assign w9796 = ~w8826 & ~w8832;
assign w9797 = ~w9795 & ~w9796;
assign w9798 = w8834 & w9797;
assign w9799 = ~w8834 & ~w9797;
assign w9800 = (~w8596 & w9797) | (~w8596 & w16212) | (w9797 & w16212);
assign w9801 = ~w9798 & ~w9800;
assign w9802 = ~w8824 & ~w9795;
assign w9803 = pi326 & ~w7108;
assign w9804 = pi325 & w7742;
assign w9805 = ~w9803 & w9804;
assign w9806 = w9803 & ~w9804;
assign w9807 = ~w9805 & ~w9806;
assign w9808 = w9802 & ~w9807;
assign w9809 = ~w9802 & w9807;
assign w9810 = ~w9808 & ~w9809;
assign w9811 = w9801 & ~w9810;
assign w9812 = ~w9801 & w9810;
assign w9813 = ~w9811 & ~w9812;
assign w9814 = w9794 & w9813;
assign w9815 = ~w9794 & ~w9813;
assign w9816 = ~w9814 & ~w9815;
assign w9817 = ~w8830 & w8833;
assign w9818 = w8830 & ~w8833;
assign w9819 = ~w9798 & ~w9799;
assign w9820 = ~w8596 & w9819;
assign w9821 = (~w9818 & w9819) | (~w9818 & w16213) | (w9819 & w16213);
assign w9822 = ~w9820 & w9821;
assign w9823 = ~w9817 & ~w9822;
assign w9824 = pi327 & w6283;
assign w9825 = pi328 & w5714;
assign w9826 = ~w9824 & w9825;
assign w9827 = w9824 & ~w9825;
assign w9828 = ~w9826 & ~w9827;
assign w9829 = ~w9822 & w16461;
assign w9830 = (w9828 & w9822) | (w9828 & w16462) | (w9822 & w16462);
assign w9831 = ~w9829 & ~w9830;
assign w9832 = w9816 & ~w9831;
assign w9833 = ~w9816 & w9831;
assign w9834 = ~w9832 & ~w9833;
assign w9835 = w9542 & w9834;
assign w9836 = ~w9542 & ~w9834;
assign w9837 = ~w9835 & ~w9836;
assign w9838 = w9531 & ~w9837;
assign w9839 = ~w9531 & w9837;
assign w9840 = ~w9838 & ~w9839;
assign w9841 = ~w9529 & w9840;
assign w9842 = w9529 & ~w9840;
assign w9843 = ~w9841 & ~w9842;
assign w9844 = pi330 & ~w4854;
assign w9845 = ~w8581 & ~w8870;
assign w9846 = ~w9844 & w9845;
assign w9847 = w9844 & ~w9845;
assign w9848 = ~w9846 & ~w9847;
assign w9849 = pi331 & ~w4708;
assign w9850 = (w8872 & w16463) | (w8872 & w16464) | (w16463 & w16464);
assign w9851 = ~w9849 & w17697;
assign w9852 = ~w9850 & ~w9851;
assign w9853 = w9848 & ~w9852;
assign w9854 = ~w9848 & w9852;
assign w9855 = ~w9853 & ~w9854;
assign w9856 = w9843 & w9855;
assign w9857 = ~w9843 & ~w9855;
assign w9858 = ~w9856 & ~w9857;
assign w9859 = w9528 & w9858;
assign w9860 = ~w9528 & ~w9858;
assign w9861 = ~w9859 & ~w9860;
assign w9862 = w9517 & ~w9861;
assign w9863 = ~w9517 & w9861;
assign w9864 = ~w9862 & ~w9863;
assign w9865 = ~w9512 & w9864;
assign w9866 = w9512 & ~w9864;
assign w9867 = ~w9865 & ~w9866;
assign w9868 = w9503 & ~w9867;
assign w9869 = ~w9503 & w9867;
assign w9870 = ~w9868 & ~w9869;
assign w9871 = w9497 & w9870;
assign w9872 = ~w9497 & ~w9870;
assign w9873 = ~w9871 & ~w9872;
assign w9874 = w9492 & ~w9873;
assign w9875 = ~w9492 & w9873;
assign w9876 = ~w9874 & ~w9875;
assign w9877 = pi338 & ~w1865;
assign w9878 = ~w8552 & w8924;
assign w9879 = ~w8551 & w9877;
assign w9880 = ~w9878 & w9879;
assign w9881 = ~w8552 & ~w9877;
assign w9882 = ~w8925 & w9881;
assign w9883 = ~w9880 & ~w9882;
assign w9884 = w9876 & w9883;
assign w9885 = ~w9876 & ~w9883;
assign w9886 = ~w9884 & ~w9885;
assign w9887 = ~w9486 & ~w9886;
assign w9888 = w9486 & w9886;
assign w9889 = ~w9887 & ~w9888;
assign w9890 = w9481 & w9889;
assign w9891 = ~w9481 & ~w9889;
assign w9892 = ~w9890 & ~w9891;
assign w9893 = ~w8941 & ~w8944;
assign w9894 = pi341 & w1101;
assign w9895 = w9893 & w9894;
assign w9896 = ~w9893 & ~w9894;
assign w9897 = ~w9895 & ~w9896;
assign w9898 = w9892 & w9897;
assign w9899 = ~w9892 & ~w9897;
assign w9900 = ~w9898 & ~w9899;
assign w9901 = ~w9476 & w9900;
assign w9902 = w9476 & ~w9900;
assign w9903 = ~w9901 & ~w9902;
assign w9904 = ~w9471 & w9903;
assign w9905 = w9471 & ~w9903;
assign w9906 = ~w9904 & ~w9905;
assign w9907 = w9466 & w9906;
assign w9908 = ~w9466 & ~w9906;
assign w9909 = ~w9907 & ~w9908;
assign w9910 = w9461 & w9909;
assign w9911 = ~w9461 & ~w9909;
assign w9912 = ~w9910 & ~w9911;
assign w9913 = w466 & w9912;
assign w9914 = ~w466 & ~w9912;
assign w9915 = ~w9913 & ~w9914;
assign w9916 = ~pi346 & w466;
assign w9917 = ~w8960 & ~w9916;
assign w9918 = ~w9915 & w9917;
assign w9919 = w9915 & ~w9917;
assign w9920 = ~w9918 & ~w9919;
assign w9921 = w9456 & w9920;
assign w9922 = ~w9456 & ~w9920;
assign w9923 = ~w9921 & ~w9922;
assign w9924 = ~w8963 & ~w8966;
assign w9925 = ~w9923 & ~w9924;
assign w9926 = w9923 & w9924;
assign w9927 = ~w9925 & ~w9926;
assign w9928 = pi283 & w9927;
assign w9929 = ~pi283 & ~w9927;
assign w9930 = ~w9928 & ~w9929;
assign w9931 = ~w9455 & w9930;
assign w9932 = w9455 & ~w9930;
assign w9933 = ~w9931 & ~w9932;
assign w9934 = w9202 & ~w9933;
assign w9935 = ~w9202 & ~w9932;
assign w9936 = ~w9931 & w9935;
assign w9937 = ~w135 & ~w9934;
assign w9938 = ~w9936 & w9937;
assign w9939 = pi161 & ~w9201;
assign w9940 = ~w9938 & w9939;
assign w9941 = ~pi160 & ~w9200;
assign w9942 = ~w9940 & w9941;
assign w9943 = ~pi090 & ~pi161;
assign w9944 = pi284 & w135;
assign w9945 = pi128 & pi295;
assign w9946 = pi296 & w464;
assign w9947 = ~w9453 & ~w9946;
assign w9948 = ~pi129 & w9453;
assign w9949 = ~w9947 & ~w9948;
assign w9950 = pi298 & w709;
assign w9951 = pi299 & w698;
assign w9952 = pi300 & w855;
assign w9953 = pi302 & w1220;
assign w9954 = pi303 & w1420;
assign w9955 = ~w9405 & ~w9409;
assign w9956 = pi304 & w1693;
assign w9957 = pi305 & w1954;
assign w9958 = pi306 & ~w2473;
assign w9959 = pi307 & w2801;
assign w9960 = pi308 & w2925;
assign w9961 = pi309 & w3304;
assign w9962 = pi310 & w3710;
assign w9963 = pi311 & w4382;
assign w9964 = pi312 & w4539;
assign w9965 = pi313 & w5316;
assign w9966 = pi314 & w5862;
assign w9967 = pi315 & w6437;
assign w9968 = ~w9307 & ~w9312;
assign w9969 = ~w9967 & w9968;
assign w9970 = w9967 & ~w9968;
assign w9971 = ~w9969 & ~w9970;
assign w9972 = pi317 & w7268;
assign w9973 = ~w9294 & ~w9297;
assign w9974 = w9972 & w9973;
assign w9975 = ~w9972 & ~w9973;
assign w9976 = ~w9974 & ~w9975;
assign w9977 = pi318 & w7909;
assign w9978 = pi319 & w9022;
assign w9979 = ~w9027 & ~w9270;
assign w9980 = ~pi151 & ~pi153;
assign w9981 = pi152 & ~w9980;
assign w9982 = ~w7262 & w9249;
assign w9983 = ~w9262 & ~w9982;
assign w9984 = pi149 & ~w9983;
assign w9985 = ~w9251 & ~w9981;
assign w9986 = ~w9984 & w9985;
assign w9987 = ~pi154 & w9986;
assign w9988 = pi154 & ~w9986;
assign w9989 = ~w9987 & ~w9988;
assign w9990 = pi153 & w9989;
assign w9991 = ~pi153 & ~w9989;
assign w9992 = ~w9990 & ~w9991;
assign w9993 = ~w9270 & w9992;
assign w9994 = ~w9022 & ~w9270;
assign w9995 = pi320 & ~w9994;
assign w9996 = ~w9022 & ~w9992;
assign w9997 = ~w9272 & w9996;
assign w9998 = w9271 & ~w9997;
assign w9999 = ~w9993 & w9995;
assign w10000 = ~w9979 & w9999;
assign w10001 = ~w9998 & w10000;
assign w10002 = w9022 & ~w9027;
assign w10003 = w9995 & ~w10002;
assign w10004 = ~w9274 & w10003;
assign w10005 = pi321 & w9992;
assign w10006 = ~w10004 & w10005;
assign w10007 = ~w10001 & ~w10006;
assign w10008 = w9978 & ~w10007;
assign w10009 = w9280 & w10008;
assign w10010 = w9281 & w10007;
assign w10011 = w9978 & w10010;
assign w10012 = ~w9978 & w10007;
assign w10013 = ~w9246 & ~w10008;
assign w10014 = ~w10012 & w10013;
assign w10015 = ~w9280 & w10014;
assign w10016 = w7909 & w9022;
assign w10017 = ~w10007 & w10016;
assign w10018 = w9282 & w10017;
assign w10019 = ~w9281 & ~w10007;
assign w10020 = ~w9022 & ~w10010;
assign w10021 = ~w10019 & w10020;
assign w10022 = ~w9284 & w10021;
assign w10023 = ~w10011 & ~w10015;
assign w10024 = ~w10018 & w10023;
assign w10025 = ~w10022 & w10024;
assign w10026 = ~w10009 & w10025;
assign w10027 = w9977 & ~w10026;
assign w10028 = ~w9977 & w10026;
assign w10029 = ~w10027 & ~w10028;
assign w10030 = ~w9286 & ~w9290;
assign w10031 = w10029 & ~w10030;
assign w10032 = ~w10029 & w10030;
assign w10033 = ~w10031 & ~w10032;
assign w10034 = w9976 & w10033;
assign w10035 = ~w9976 & ~w10033;
assign w10036 = ~w10034 & ~w10035;
assign w10037 = w9302 & ~w10036;
assign w10038 = pi316 & w6652;
assign w10039 = w10037 & w10038;
assign w10040 = ~w10036 & ~w10038;
assign w10041 = w10036 & w10038;
assign w10042 = ~w9243 & ~w10040;
assign w10043 = ~w10041 & w10042;
assign w10044 = ~w9302 & w10036;
assign w10045 = w6437 & w6652;
assign w10046 = w10044 & w10045;
assign w10047 = ~w9301 & ~w10043;
assign w10048 = ~w10046 & w10047;
assign w10049 = ~pi316 & ~w10036;
assign w10050 = ~w10041 & ~w10049;
assign w10051 = w9301 & w10050;
assign w10052 = ~w10048 & ~w10051;
assign w10053 = ~w6652 & ~w10037;
assign w10054 = ~w10044 & w10053;
assign w10055 = ~w9304 & w10054;
assign w10056 = ~w10039 & ~w10052;
assign w10057 = ~w10055 & w10056;
assign w10058 = ~w9971 & w10057;
assign w10059 = w9971 & ~w10057;
assign w10060 = ~w10058 & ~w10059;
assign w10061 = w9966 & w10060;
assign w10062 = ~w9966 & ~w10060;
assign w10063 = ~w10061 & ~w10062;
assign w10064 = ~w9315 & ~w9318;
assign w10065 = w10063 & w10064;
assign w10066 = ~w10063 & ~w10064;
assign w10067 = ~w10065 & ~w10066;
assign w10068 = ~w9322 & ~w9325;
assign w10069 = ~w10067 & w10068;
assign w10070 = w10067 & ~w10068;
assign w10071 = ~w10069 & ~w10070;
assign w10072 = w9965 & w10071;
assign w10073 = ~w9965 & ~w10071;
assign w10074 = ~w10072 & ~w10073;
assign w10075 = ~w9964 & ~w10074;
assign w10076 = w9964 & w10074;
assign w10077 = ~w10075 & ~w10076;
assign w10078 = ~w9329 & ~w9332;
assign w10079 = ~w10077 & w10078;
assign w10080 = w10077 & ~w10078;
assign w10081 = ~w10079 & ~w10080;
assign w10082 = ~w9334 & ~w9338;
assign w10083 = w10081 & ~w10082;
assign w10084 = ~w10081 & w10082;
assign w10085 = ~w10083 & ~w10084;
assign w10086 = w9963 & w10085;
assign w10087 = ~w9963 & ~w10085;
assign w10088 = ~w10086 & ~w10087;
assign w10089 = ~w9349 & ~w9357;
assign w10090 = ~w9350 & ~w10089;
assign w10091 = w10088 & w10090;
assign w10092 = ~w10088 & ~w10090;
assign w10093 = ~w10091 & ~w10092;
assign w10094 = w9962 & ~w10093;
assign w10095 = ~w9962 & w10093;
assign w10096 = ~w10094 & ~w10095;
assign w10097 = w9961 & ~w10096;
assign w10098 = ~w9961 & w10096;
assign w10099 = ~w10097 & ~w10098;
assign w10100 = ~w9359 & ~w9363;
assign w10101 = w10099 & ~w10100;
assign w10102 = ~w10099 & w10100;
assign w10103 = ~w10101 & ~w10102;
assign w10104 = ~w9960 & ~w10103;
assign w10105 = w9960 & w10103;
assign w10106 = ~w10104 & ~w10105;
assign w10107 = ~w9233 & ~w9365;
assign w10108 = w10106 & w10107;
assign w10109 = ~w10106 & ~w10107;
assign w10110 = ~w10108 & ~w10109;
assign w10111 = ~w9368 & ~w9372;
assign w10112 = w10110 & ~w10111;
assign w10113 = ~w10110 & w10111;
assign w10114 = ~w10112 & ~w10113;
assign w10115 = w9959 & w10114;
assign w10116 = ~w9959 & ~w10114;
assign w10117 = ~w10115 & ~w10116;
assign w10118 = pi306 & w9378;
assign w10119 = ~w9385 & ~w10118;
assign w10120 = ~w10117 & w10119;
assign w10121 = w10117 & ~w10119;
assign w10122 = ~w10120 & ~w10121;
assign w10123 = w9958 & w10122;
assign w10124 = ~w9958 & ~w10122;
assign w10125 = ~w10123 & ~w10124;
assign w10126 = w9957 & w10125;
assign w10127 = ~w9957 & ~w10125;
assign w10128 = ~w10126 & ~w10127;
assign w10129 = ~w9395 & ~w9399;
assign w10130 = ~w10128 & w10129;
assign w10131 = w10128 & ~w10129;
assign w10132 = ~w10130 & ~w10131;
assign w10133 = ~w9956 & w10132;
assign w10134 = w9956 & ~w10132;
assign w10135 = ~w10133 & ~w10134;
assign w10136 = ~w9225 & ~w9402;
assign w10137 = ~w10135 & w10136;
assign w10138 = w10135 & ~w10136;
assign w10139 = ~w10137 & ~w10138;
assign w10140 = w9955 & w10139;
assign w10141 = ~w9955 & ~w10139;
assign w10142 = ~w10140 & ~w10141;
assign w10143 = w9954 & w10142;
assign w10144 = ~w9954 & ~w10142;
assign w10145 = ~w10143 & ~w10144;
assign w10146 = w9953 & w10145;
assign w10147 = ~w9953 & ~w10145;
assign w10148 = ~w10146 & ~w10147;
assign w10149 = ~w9422 & ~w9430;
assign w10150 = ~w9415 & ~w10149;
assign w10151 = ~w10148 & w10150;
assign w10152 = w10148 & ~w10150;
assign w10153 = ~w10151 & ~w10152;
assign w10154 = pi301 & w1159;
assign w10155 = ~w9432 & w9434;
assign w10156 = ~w9431 & ~w10155;
assign w10157 = ~w10154 & ~w10156;
assign w10158 = w10154 & w10156;
assign w10159 = ~w10157 & ~w10158;
assign w10160 = w10153 & w10159;
assign w10161 = ~w10153 & ~w10159;
assign w10162 = ~w10160 & ~w10161;
assign w10163 = w9952 & w10162;
assign w10164 = ~w9952 & ~w10162;
assign w10165 = ~w10163 & ~w10164;
assign w10166 = ~w9218 & ~w9439;
assign w10167 = w10165 & ~w10166;
assign w10168 = ~w10165 & w10166;
assign w10169 = ~w10167 & ~w10168;
assign w10170 = ~w9213 & ~w9441;
assign w10171 = w10169 & ~w10170;
assign w10172 = ~w10169 & w10170;
assign w10173 = ~w10171 & ~w10172;
assign w10174 = w9951 & w10173;
assign w10175 = ~w9951 & ~w10173;
assign w10176 = ~w10174 & ~w10175;
assign w10177 = w9950 & w10176;
assign w10178 = ~w9950 & ~w10176;
assign w10179 = ~w10177 & ~w10178;
assign w10180 = ~w9208 & ~w9444;
assign w10181 = ~w10179 & w10180;
assign w10182 = w10179 & ~w10180;
assign w10183 = ~w10181 & ~w10182;
assign w10184 = w705 & ~w9446;
assign w10185 = ~w5426 & ~w10184;
assign w10186 = ~w9449 & ~w10185;
assign w10187 = w8970 & w9185;
assign w10188 = pi128 & w9448;
assign w10189 = pi130 & ~w10187;
assign w10190 = ~w9447 & w10189;
assign w10191 = ~w10188 & w10190;
assign w10192 = ~w10186 & ~w10191;
assign w10193 = pi297 & ~w10192;
assign w10194 = ~w9447 & w10187;
assign w10195 = w653 & w10194;
assign w10196 = ~w10193 & ~w10195;
assign w10197 = w10183 & ~w10196;
assign w10198 = ~w10183 & w10196;
assign w10199 = ~w10197 & ~w10198;
assign w10200 = w9949 & ~w10199;
assign w10201 = ~w9949 & w10199;
assign w10202 = ~w10200 & ~w10201;
assign w10203 = w9945 & ~w10202;
assign w10204 = ~w9945 & w10202;
assign w10205 = ~w10203 & ~w10204;
assign w10206 = ~w9931 & ~w9935;
assign w10207 = w10205 & w10206;
assign w10208 = ~w10205 & ~w10206;
assign w10209 = ~w10207 & ~w10208;
assign w10210 = ~w9925 & ~w9928;
assign w10211 = pi284 & ~w10210;
assign w10212 = ~pi284 & w10210;
assign w10213 = ~w10211 & ~w10212;
assign w10214 = pi348 & w456;
assign w10215 = pi347 & w466;
assign w10216 = ~w9921 & ~w10215;
assign w10217 = w466 & w9921;
assign w10218 = ~w10216 & ~w10217;
assign w10219 = w456 & w8958;
assign w10220 = ~w9913 & ~w10219;
assign w10221 = ~w9914 & ~w10220;
assign w10222 = w537 & ~w10221;
assign w10223 = pi346 & ~w10222;
assign w10224 = ~w537 & w10221;
assign w10225 = ~w9460 & ~w9910;
assign w10226 = pi345 & ~w615;
assign w10227 = ~w10225 & w10226;
assign w10228 = w10225 & ~w10226;
assign w10229 = ~w10227 & ~w10228;
assign w10230 = pi342 & w1101;
assign w10231 = ~w9475 & ~w9902;
assign w10232 = ~w10230 & ~w10231;
assign w10233 = w10230 & w10231;
assign w10234 = ~w10232 & ~w10233;
assign w10235 = pi341 & w1339;
assign w10236 = ~w9895 & ~w9898;
assign w10237 = w10235 & ~w10236;
assign w10238 = ~w10235 & w10236;
assign w10239 = ~w10237 & ~w10238;
assign w10240 = ~w9479 & ~w9890;
assign w10241 = pi340 & w1602;
assign w10242 = ~w10240 & w10241;
assign w10243 = w10240 & ~w10241;
assign w10244 = ~w10242 & ~w10243;
assign w10245 = ~w9484 & ~w9888;
assign w10246 = pi339 & ~w1865;
assign w10247 = w10245 & ~w10246;
assign w10248 = ~w10245 & w10246;
assign w10249 = ~w10247 & ~w10248;
assign w10250 = pi337 & ~w2373;
assign w10251 = ~w9491 & ~w9874;
assign w10252 = pi336 & w2698;
assign w10253 = ~w9867 & w16465;
assign w10254 = ~w9495 & ~w9503;
assign w10255 = w9867 & w10254;
assign w10256 = ~w9496 & ~w10255;
assign w10257 = (w10252 & ~w10256) | (w10252 & w16466) | (~w10256 & w16466);
assign w10258 = w10256 & w16467;
assign w10259 = ~w10257 & ~w10258;
assign w10260 = pi335 & ~w3183;
assign w10261 = pi334 & ~w3568;
assign w10262 = (~w9510 & w9864) | (~w9510 & w16468) | (w9864 & w16468);
assign w10263 = w10261 & ~w10262;
assign w10264 = ~w10261 & w10262;
assign w10265 = ~w10263 & ~w10264;
assign w10266 = w10260 & ~w10265;
assign w10267 = ~w10260 & w10265;
assign w10268 = ~w10266 & ~w10267;
assign w10269 = w10259 & w10268;
assign w10270 = ~w10259 & ~w10268;
assign w10271 = ~w10269 & ~w10270;
assign w10272 = ~w9501 & ~w9868;
assign w10273 = (~w9515 & w9861) | (~w9515 & w16469) | (w9861 & w16469);
assign w10274 = pi329 & w5714;
assign w10275 = (~w9838 & ~w9840) | (~w9838 & w16470) | (~w9840 & w16470);
assign w10276 = ~w10274 & ~w10275;
assign w10277 = w10274 & w10275;
assign w10278 = ~w10276 & ~w10277;
assign w10279 = pi328 & w6283;
assign w10280 = w9539 & ~w9825;
assign w10281 = ~w9539 & w9825;
assign w10282 = ~w9816 & ~w9823;
assign w10283 = w9816 & w9823;
assign w10284 = ~w10282 & ~w10283;
assign w10285 = (w9824 & w9532) | (w9824 & w16471) | (w9532 & w16471);
assign w10286 = ~w9532 & w16472;
assign w10287 = ~w10285 & ~w10286;
assign w10288 = w10284 & ~w10287;
assign w10289 = ~w10284 & w10287;
assign w10290 = ~w10281 & ~w10288;
assign w10291 = ~w10289 & w10290;
assign w10292 = ~w10280 & ~w10291;
assign w10293 = w10279 & w10292;
assign w10294 = ~w10279 & ~w10292;
assign w10295 = ~w10293 & ~w10294;
assign w10296 = pi322 & pi323;
assign w10297 = ~w9553 & w16215;
assign w10298 = (~w9772 & w9553) | (~w9772 & w16216) | (w9553 & w16216);
assign w10299 = ~w10297 & ~w10298;
assign w10300 = w9770 & w10299;
assign w10301 = ~w9770 & ~w10299;
assign w10302 = ~w10300 & ~w10301;
assign w10303 = w9771 & w10302;
assign w10304 = pi154 & pi258;
assign w10305 = (w10304 & ~w10302) | (w10304 & w16217) | (~w10302 & w16217);
assign w10306 = pi153 & w10305;
assign w10307 = w10302 & w16218;
assign w10308 = ~pi153 & ~w10304;
assign w10309 = pi259 & ~w10308;
assign w10310 = (w10309 & ~w10302) | (w10309 & w16473) | (~w10302 & w16473);
assign w10311 = ~w10306 & w10310;
assign w10312 = ~w10305 & ~w10307;
assign w10313 = w5690 & ~w10312;
assign w10314 = ~w10311 & ~w10313;
assign w10315 = pi151 & pi261;
assign w10316 = pi150 & pi262;
assign w10317 = ~w9762 & ~w9764;
assign w10318 = (~w10316 & w10317) | (~w10316 & w16219) | (w10317 & w16219);
assign w10319 = ~w10317 & w16220;
assign w10320 = ~w10318 & ~w10319;
assign w10321 = pi149 & pi263;
assign w10322 = (~w8795 & ~w8797) | (~w8795 & w15946) | (~w8797 & w15946);
assign w10323 = (~w9750 & w10322) | (~w9750 & w16221) | (w10322 & w16221);
assign w10324 = ~w10323 & w15947;
assign w10325 = (~w10321 & w10323) | (~w10321 & w15948) | (w10323 & w15948);
assign w10326 = ~w10324 & ~w10325;
assign w10327 = w9738 & w9745;
assign w10328 = ~w9746 & ~w10327;
assign w10329 = pi148 & pi264;
assign w10330 = pi147 & pi265;
assign w10331 = pi146 & pi266;
assign w10332 = ~w9728 & w9731;
assign w10333 = (w10331 & w10332) | (w10331 & w15949) | (w10332 & w15949);
assign w10334 = ~w10332 & w15950;
assign w10335 = ~w10333 & ~w10334;
assign w10336 = pi144 & pi268;
assign w10337 = pi143 & pi269;
assign w10338 = w9572 & ~w9706;
assign w10339 = ~w10338 & w15951;
assign w10340 = (~w10337 & w10338) | (~w10337 & w15952) | (w10338 & w15952);
assign w10341 = ~w10339 & ~w10340;
assign w10342 = pi142 & pi270;
assign w10343 = pi141 & pi271;
assign w10344 = pi140 & pi272;
assign w10345 = ~w9681 & ~w9683;
assign w10346 = ~w10345 & w15953;
assign w10347 = (~w10344 & w10345) | (~w10344 & w15954) | (w10345 & w15954);
assign w10348 = ~w10346 & ~w10347;
assign w10349 = pi139 & pi273;
assign w10350 = w9669 & w9676;
assign w10351 = ~w9678 & ~w10350;
assign w10352 = pi138 & pi274;
assign w10353 = pi137 & pi275;
assign w10354 = pi136 & pi276;
assign w10355 = pi135 & pi277;
assign w10356 = (~w9637 & ~w9638) | (~w9637 & w15955) | (~w9638 & w15955);
assign w10357 = pi134 & pi278;
assign w10358 = (pi133 & w9584) | (pi133 & w16222) | (w9584 & w16222);
assign w10359 = pi133 & pi279;
assign w10360 = pi132 & pi280;
assign w10361 = pi131 & pi281;
assign w10362 = pi130 & pi282;
assign w10363 = pi128 & pi284;
assign w10364 = ~w9600 & w9603;
assign w10365 = ~w9592 & ~w10364;
assign w10366 = w10363 & ~w10365;
assign w10367 = ~w10363 & w10365;
assign w10368 = ~w10366 & ~w10367;
assign w10369 = w9591 & ~w10368;
assign w10370 = ~w9591 & w10368;
assign w10371 = ~w10369 & ~w10370;
assign w10372 = ~w9607 & ~w10364;
assign w10373 = (~w10372 & w8673) | (~w10372 & w16223) | (w8673 & w16223);
assign w10374 = (~w9595 & w8673) | (~w9595 & w16474) | (w8673 & w16474);
assign w10375 = ~w10373 & ~w10374;
assign w10376 = ~w10371 & w10375;
assign w10377 = w10371 & ~w10375;
assign w10378 = ~w10376 & ~w10377;
assign w10379 = w10362 & w10378;
assign w10380 = ~w10362 & ~w10378;
assign w10381 = ~w10379 & ~w10380;
assign w10382 = w10361 & w10381;
assign w10383 = ~w10361 & ~w10381;
assign w10384 = ~w10382 & ~w10383;
assign w10385 = ~w9617 & ~w9620;
assign w10386 = w10384 & ~w10385;
assign w10387 = ~w10384 & w10385;
assign w10388 = ~w10386 & ~w10387;
assign w10389 = w10360 & ~w10388;
assign w10390 = ~w10360 & w10388;
assign w10391 = ~w10389 & ~w10390;
assign w10392 = (~w9623 & w9626) | (~w9623 & w16224) | (w9626 & w16224);
assign w10393 = w10391 & ~w10392;
assign w10394 = ~w10391 & w10392;
assign w10395 = ~w10393 & ~w10394;
assign w10396 = w10359 & w10395;
assign w10397 = ~w10359 & ~w10395;
assign w10398 = ~w10396 & ~w10397;
assign w10399 = w10358 & w10398;
assign w10400 = ~w10358 & ~w10398;
assign w10401 = ~w10399 & ~w10400;
assign w10402 = w10357 & ~w10401;
assign w10403 = ~pi134 & ~w10358;
assign w10404 = ~pi278 & ~w9631;
assign w10405 = ~w10403 & ~w10404;
assign w10406 = w10398 & ~w10405;
assign w10407 = pi133 & w10357;
assign w10408 = ~w10398 & ~w10407;
assign w10409 = w10405 & w10408;
assign w10410 = ~w10402 & w16225;
assign w10411 = ~w10356 & ~w10410;
assign w10412 = w10356 & w10410;
assign w10413 = ~w10411 & ~w10412;
assign w10414 = w10355 & w10413;
assign w10415 = ~w10355 & ~w10413;
assign w10416 = ~w10414 & ~w10415;
assign w10417 = (~w9644 & ~w9646) | (~w9644 & w15957) | (~w9646 & w15957);
assign w10418 = w10416 & ~w10417;
assign w10419 = ~w10416 & w10417;
assign w10420 = ~w10418 & ~w10419;
assign w10421 = ~w9650 & ~w9654;
assign w10422 = ~w10421 & w15958;
assign w10423 = (w10420 & w10421) | (w10420 & w15959) | (w10421 & w15959);
assign w10424 = ~w10422 & ~w10423;
assign w10425 = w10354 & ~w10424;
assign w10426 = ~w10354 & w10424;
assign w10427 = ~w10425 & ~w10426;
assign w10428 = ~w9658 & w9662;
assign w10429 = ~w9659 & ~w10428;
assign w10430 = ~w10427 & w10429;
assign w10431 = w10427 & ~w10429;
assign w10432 = ~w10430 & ~w10431;
assign w10433 = w10353 & w10432;
assign w10434 = ~w10353 & ~w10432;
assign w10435 = ~w10433 & ~w10434;
assign w10436 = w10352 & w10435;
assign w10437 = ~w10352 & ~w10435;
assign w10438 = ~w10436 & ~w10437;
assign w10439 = (w9670 & w9578) | (w9670 & w16475) | (w9578 & w16475);
assign w10440 = ~w9667 & ~w10439;
assign w10441 = w10438 & ~w10440;
assign w10442 = ~w10438 & w10440;
assign w10443 = ~w10441 & ~w10442;
assign w10444 = ~w10351 & w10443;
assign w10445 = w10351 & ~w10443;
assign w10446 = ~w10444 & ~w10445;
assign w10447 = w10349 & w10446;
assign w10448 = ~w10349 & ~w10446;
assign w10449 = ~w10447 & ~w10448;
assign w10450 = w10348 & ~w10449;
assign w10451 = ~w10348 & w10449;
assign w10452 = ~w10450 & ~w10451;
assign w10453 = w10343 & ~w10452;
assign w10454 = ~w10343 & w10452;
assign w10455 = ~w10453 & ~w10454;
assign w10456 = ~w9690 & w9693;
assign w10457 = ~w9689 & ~w10456;
assign w10458 = w10455 & ~w10457;
assign w10459 = ~w10455 & w10457;
assign w10460 = ~w10458 & ~w10459;
assign w10461 = w9692 & w9699;
assign w10462 = ~w9702 & ~w10461;
assign w10463 = w10460 & ~w10462;
assign w10464 = ~w10460 & w10462;
assign w10465 = ~w10463 & ~w10464;
assign w10466 = w10342 & w10465;
assign w10467 = ~w10342 & ~w10465;
assign w10468 = ~w10466 & ~w10467;
assign w10469 = w10341 & w10468;
assign w10470 = ~w10341 & ~w10468;
assign w10471 = ~w10469 & ~w10470;
assign w10472 = w10336 & w10471;
assign w10473 = ~w10336 & ~w10471;
assign w10474 = ~w10472 & ~w10473;
assign w10475 = ~w9711 & w9715;
assign w10476 = ~w9712 & ~w10475;
assign w10477 = w10474 & w10476;
assign w10478 = ~w10474 & ~w10476;
assign w10479 = ~w10477 & ~w10478;
assign w10480 = ~w9714 & w9721;
assign w10481 = ~w9725 & ~w10480;
assign w10482 = w10479 & ~w10481;
assign w10483 = ~w10479 & w10481;
assign w10484 = ~w10482 & ~w10483;
assign w10485 = pi145 & pi267;
assign w10486 = ~w10484 & w10485;
assign w10487 = w10484 & ~w10485;
assign w10488 = ~w10486 & ~w10487;
assign w10489 = w10335 & ~w10488;
assign w10490 = ~w10335 & w10488;
assign w10491 = ~w10489 & ~w10490;
assign w10492 = w10330 & w10491;
assign w10493 = ~w10330 & ~w10491;
assign w10494 = ~w10492 & ~w10493;
assign w10495 = (~w9739 & w9567) | (~w9739 & w16476) | (w9567 & w16476);
assign w10496 = ~w9735 & ~w10495;
assign w10497 = w10494 & w10496;
assign w10498 = ~w10494 & ~w10496;
assign w10499 = ~w10497 & ~w10498;
assign w10500 = w10329 & w10499;
assign w10501 = ~w10329 & ~w10499;
assign w10502 = ~w10500 & ~w10501;
assign w10503 = w10328 & ~w10502;
assign w10504 = ~w10328 & w10502;
assign w10505 = ~w10503 & ~w10504;
assign w10506 = w10326 & ~w10505;
assign w10507 = ~w10326 & w10505;
assign w10508 = ~w10506 & ~w10507;
assign w10509 = w10320 & ~w10508;
assign w10510 = ~w10320 & w10508;
assign w10511 = ~w10509 & ~w10510;
assign w10512 = ~w10315 & ~w10511;
assign w10513 = w10315 & w10511;
assign w10514 = ~w10512 & ~w10513;
assign w10515 = pi151 & w9562;
assign w10516 = ~w9768 & ~w10515;
assign w10517 = w10514 & ~w10516;
assign w10518 = ~w10514 & w10516;
assign w10519 = ~w10517 & ~w10518;
assign w10520 = (~w10297 & ~w9770) | (~w10297 & w16226) | (~w9770 & w16226);
assign w10521 = pi152 & pi260;
assign w10522 = ~w10520 & w10521;
assign w10523 = w10520 & ~w10521;
assign w10524 = ~w10522 & ~w10523;
assign w10525 = w10519 & w10524;
assign w10526 = ~w10519 & ~w10524;
assign w10527 = ~w10525 & ~w10526;
assign w10528 = w10314 & w10527;
assign w10529 = ~w10314 & ~w10527;
assign w10530 = ~w10528 & ~w10529;
assign w10531 = ~w9771 & ~w10302;
assign w10532 = ~w10303 & ~w10531;
assign w10533 = ~w8599 & ~w9556;
assign w10534 = w10532 & w10533;
assign w10535 = w9556 & ~w9784;
assign w10536 = w8599 & ~w9556;
assign w10537 = ~w10532 & w10536;
assign w10538 = ~w10535 & ~w10537;
assign w10539 = ~w10530 & w10538;
assign w10540 = (w10296 & ~w10530) | (w10296 & w15960) | (~w10530 & w15960);
assign w10541 = ~w10539 & w10540;
assign w10542 = pi323 & ~w9784;
assign w10543 = w9557 & ~w10532;
assign w10544 = ~w10534 & ~w10543;
assign w10545 = w10530 & w10544;
assign w10546 = (pi322 & w10530) | (pi322 & w15961) | (w10530 & w15961);
assign w10547 = ~w10545 & w10546;
assign w10548 = ~w10542 & ~w10547;
assign w10549 = ~w9786 & ~w9789;
assign w10550 = (~w10549 & w10548) | (~w10549 & w16227) | (w10548 & w16227);
assign w10551 = ~w10541 & w10549;
assign w10552 = ~w10548 & w10551;
assign w10553 = ~w10550 & ~w10552;
assign w10554 = pi325 & ~w8367;
assign w10555 = pi324 & w8814;
assign w10556 = w9794 & ~w9802;
assign w10557 = ~w10555 & w17698;
assign w10558 = (w9794 & w16228) | (w9794 & w16229) | (w16228 & w16229);
assign w10559 = ~w10557 & ~w10558;
assign w10560 = w10554 & ~w10559;
assign w10561 = ~w10554 & w10559;
assign w10562 = ~w10560 & ~w10561;
assign w10563 = w10553 & w10562;
assign w10564 = ~w10553 & ~w10562;
assign w10565 = ~w10563 & ~w10564;
assign w10566 = ~w9794 & w9802;
assign w10567 = ~w10556 & ~w10566;
assign w10568 = w9804 & w10567;
assign w10569 = ~w9804 & ~w10567;
assign w10570 = ~w9801 & ~w10569;
assign w10571 = ~w10568 & ~w10570;
assign w10572 = w10565 & ~w10571;
assign w10573 = ~w10565 & w10571;
assign w10574 = ~w10572 & ~w10573;
assign w10575 = pi326 & w7742;
assign w10576 = w9803 & w9816;
assign w10577 = ~w10282 & ~w10576;
assign w10578 = w10575 & ~w10577;
assign w10579 = ~w10575 & w10577;
assign w10580 = ~w10578 & ~w10579;
assign w10581 = pi327 & ~w7108;
assign w10582 = (w10284 & w16477) | (w10284 & w16478) | (w16477 & w16478);
assign w10583 = ~w10581 & w17699;
assign w10584 = ~w10582 & ~w10583;
assign w10585 = w10580 & ~w10584;
assign w10586 = ~w10580 & w10584;
assign w10587 = ~w10585 & ~w10586;
assign w10588 = w10574 & w10587;
assign w10589 = ~w10574 & ~w10587;
assign w10590 = ~w10588 & ~w10589;
assign w10591 = w10295 & ~w10590;
assign w10592 = ~w10295 & w10590;
assign w10593 = ~w10591 & ~w10592;
assign w10594 = w10278 & w10593;
assign w10595 = ~w10278 & ~w10593;
assign w10596 = ~w10594 & ~w10595;
assign w10597 = (~w9847 & w9843) | (~w9847 & w15964) | (w9843 & w15964);
assign w10598 = pi330 & w5194;
assign w10599 = w10597 & ~w10598;
assign w10600 = ~w9843 & w16230;
assign w10601 = w5194 & ~w10597;
assign w10602 = ~w10600 & w10601;
assign w10603 = ~w10599 & ~w10602;
assign w10604 = w10596 & w10603;
assign w10605 = ~w10596 & ~w10603;
assign w10606 = ~w10604 & ~w10605;
assign w10607 = ~w10273 & w10606;
assign w10608 = w10273 & ~w10606;
assign w10609 = ~w10607 & ~w10608;
assign w10610 = pi331 & ~w4854;
assign w10611 = pi332 & ~w4708;
assign w10612 = (~w9524 & ~w9858) | (~w9524 & w16231) | (~w9858 & w16231);
assign w10613 = w10611 & ~w10612;
assign w10614 = ~w10611 & w10612;
assign w10615 = ~w10613 & ~w10614;
assign w10616 = w10610 & w10615;
assign w10617 = ~w10610 & ~w10615;
assign w10618 = ~w10616 & ~w10617;
assign w10619 = w10609 & w10618;
assign w10620 = ~w10609 & ~w10618;
assign w10621 = ~w10619 & ~w10620;
assign w10622 = pi333 & w3979;
assign w10623 = ~w9850 & w9858;
assign w10624 = ~w9851 & ~w10623;
assign w10625 = ~w10622 & w10624;
assign w10626 = w10622 & ~w10624;
assign w10627 = ~w10625 & ~w10626;
assign w10628 = w10621 & w10627;
assign w10629 = ~w10621 & ~w10627;
assign w10630 = ~w10628 & ~w10629;
assign w10631 = w10272 & ~w10630;
assign w10632 = ~w10272 & w10630;
assign w10633 = ~w10631 & ~w10632;
assign w10634 = w10271 & w10633;
assign w10635 = ~w10271 & ~w10633;
assign w10636 = ~w10634 & ~w10635;
assign w10637 = w10251 & ~w10636;
assign w10638 = ~w10251 & w10636;
assign w10639 = ~w10637 & ~w10638;
assign w10640 = ~w10250 & ~w10639;
assign w10641 = w10250 & w10639;
assign w10642 = ~w10640 & ~w10641;
assign w10643 = ~w2170 & w9880;
assign w10644 = pi338 & ~w2170;
assign w10645 = ~w9880 & ~w10644;
assign w10646 = ~w10643 & ~w10645;
assign w10647 = w9884 & ~w10646;
assign w10648 = ~w9884 & w10646;
assign w10649 = ~w10647 & ~w10648;
assign w10650 = w10642 & w10649;
assign w10651 = ~w10642 & ~w10649;
assign w10652 = ~w10650 & ~w10651;
assign w10653 = w10249 & ~w10652;
assign w10654 = ~w10249 & w10652;
assign w10655 = ~w10653 & ~w10654;
assign w10656 = ~w10244 & ~w10655;
assign w10657 = w10244 & w10655;
assign w10658 = ~w10656 & ~w10657;
assign w10659 = w10239 & w10658;
assign w10660 = ~w10239 & ~w10658;
assign w10661 = ~w10659 & ~w10660;
assign w10662 = ~w10234 & ~w10661;
assign w10663 = w10234 & w10661;
assign w10664 = ~w10662 & ~w10663;
assign w10665 = pi343 & ~w955;
assign w10666 = ~w9470 & ~w9905;
assign w10667 = w10665 & ~w10666;
assign w10668 = ~w10665 & w10666;
assign w10669 = ~w10667 & ~w10668;
assign w10670 = w10664 & w10669;
assign w10671 = ~w10664 & ~w10669;
assign w10672 = ~w10670 & ~w10671;
assign w10673 = pi344 & ~w793;
assign w10674 = (~w9464 & ~w9466) | (~w9464 & w15965) | (~w9466 & w15965);
assign w10675 = w10673 & ~w10674;
assign w10676 = ~w10673 & w10674;
assign w10677 = ~w10675 & ~w10676;
assign w10678 = w10672 & w10677;
assign w10679 = ~w10672 & ~w10677;
assign w10680 = ~w10678 & ~w10679;
assign w10681 = w10229 & w10680;
assign w10682 = ~w10229 & ~w10680;
assign w10683 = ~w10681 & ~w10682;
assign w10684 = (w10683 & ~w10223) | (w10683 & w15966) | (~w10223 & w15966);
assign w10685 = w10223 & w10978;
assign w10686 = ~w10684 & ~w10685;
assign w10687 = w10218 & ~w10686;
assign w10688 = ~w10218 & w10686;
assign w10689 = ~w10687 & ~w10688;
assign w10690 = w10214 & w10689;
assign w10691 = ~w10214 & ~w10689;
assign w10692 = ~w10690 & ~w10691;
assign w10693 = w10213 & ~w10692;
assign w10694 = ~w10213 & w10692;
assign w10695 = ~w10693 & ~w10694;
assign w10696 = w10209 & ~w10695;
assign w10697 = ~w10209 & w10695;
assign w10698 = ~w10696 & ~w10697;
assign w10699 = ~w135 & ~w10698;
assign w10700 = pi161 & ~w9944;
assign w10701 = ~w10699 & w10700;
assign w10702 = ~pi160 & ~w9943;
assign w10703 = ~w10701 & w10702;
assign w10704 = ~pi091 & ~pi161;
assign w10705 = pi128 & pi294;
assign w10706 = ~pi129 & w10203;
assign w10707 = pi295 & w464;
assign w10708 = ~w10203 & ~w10707;
assign w10709 = ~w10706 & ~w10708;
assign w10710 = pi296 & ~w653;
assign w10711 = pi297 & w709;
assign w10712 = pi298 & w698;
assign w10713 = (~w10177 & ~w10179) | (~w10177 & w15967) | (~w10179 & w15967);
assign w10714 = pi300 & w1159;
assign w10715 = ~w10163 & ~w10167;
assign w10716 = pi301 & w1220;
assign w10717 = pi302 & w1420;
assign w10718 = pi303 & w1693;
assign w10719 = w10140 & ~w10718;
assign w10720 = w9955 & w16232;
assign w10721 = (w1420 & w9955) | (w1420 & w16233) | (w9955 & w16233);
assign w10722 = ~w1693 & ~w10721;
assign w10723 = w1693 & w10721;
assign w10724 = pi303 & ~w10720;
assign w10725 = ~w10722 & w10724;
assign w10726 = (~w10719 & ~w10725) | (~w10719 & w16479) | (~w10725 & w16479);
assign w10727 = pi304 & w1954;
assign w10728 = ~w10134 & ~w10138;
assign w10729 = w10727 & ~w10728;
assign w10730 = ~w10727 & w10728;
assign w10731 = ~w10729 & ~w10730;
assign w10732 = pi307 & w2925;
assign w10733 = pi309 & w3710;
assign w10734 = pi311 & w4539;
assign w10735 = ~w10075 & ~w10080;
assign w10736 = pi312 & w5316;
assign w10737 = w10735 & w10736;
assign w10738 = ~w10735 & ~w10736;
assign w10739 = ~w10737 & ~w10738;
assign w10740 = pi314 & w6437;
assign w10741 = pi315 & w6652;
assign w10742 = pi316 & w7268;
assign w10743 = pi317 & w7909;
assign w10744 = pi318 & w9022;
assign w10745 = ~w10027 & ~w10031;
assign w10746 = pi319 & w9270;
assign w10747 = ~pi155 & w9986;
assign w10748 = pi155 & ~w9986;
assign w10749 = ~w10747 & ~w10748;
assign w10750 = ~w9987 & ~w9990;
assign w10751 = w10749 & w10750;
assign w10752 = ~w10749 & ~w10750;
assign w10753 = ~w10751 & ~w10752;
assign w10754 = pi321 & w10753;
assign w10755 = ~w9274 & ~w9276;
assign w10756 = w9270 & ~w10755;
assign w10757 = ~w9993 & ~w10756;
assign w10758 = w9992 & ~w10755;
assign w10759 = pi320 & ~w10758;
assign w10760 = ~w10757 & w10759;
assign w10761 = w10754 & ~w10760;
assign w10762 = ~w9992 & ~w10754;
assign w10763 = w10756 & ~w10762;
assign w10764 = ~w9271 & w9992;
assign w10765 = ~w10754 & w10764;
assign w10766 = ~w9276 & w10765;
assign w10767 = ~w10756 & ~w10766;
assign w10768 = pi320 & ~w10763;
assign w10769 = ~w10767 & w10768;
assign w10770 = ~w10761 & ~w10769;
assign w10771 = ~w10008 & ~w10025;
assign w10772 = ~w10012 & ~w10771;
assign w10773 = ~w10770 & w10772;
assign w10774 = w10770 & ~w10772;
assign w10775 = ~w10773 & ~w10774;
assign w10776 = w10746 & ~w10775;
assign w10777 = ~w10746 & w10775;
assign w10778 = ~w10776 & ~w10777;
assign w10779 = ~w10745 & ~w10778;
assign w10780 = w10745 & w10778;
assign w10781 = ~w10779 & ~w10780;
assign w10782 = w10744 & ~w10781;
assign w10783 = ~w10744 & w10781;
assign w10784 = ~w10782 & ~w10783;
assign w10785 = w10743 & ~w10784;
assign w10786 = ~w10743 & w10784;
assign w10787 = ~w10785 & ~w10786;
assign w10788 = ~w9974 & ~w10034;
assign w10789 = w10787 & ~w10788;
assign w10790 = ~w10787 & w10788;
assign w10791 = ~w10789 & ~w10790;
assign w10792 = ~w10041 & ~w10057;
assign w10793 = ~w10040 & ~w10792;
assign w10794 = w10791 & w10793;
assign w10795 = ~w10791 & ~w10793;
assign w10796 = ~w10794 & ~w10795;
assign w10797 = w10742 & w10796;
assign w10798 = ~w10742 & ~w10796;
assign w10799 = ~w10797 & ~w10798;
assign w10800 = w10741 & w10799;
assign w10801 = ~w10741 & ~w10799;
assign w10802 = ~w10800 & ~w10801;
assign w10803 = ~w9970 & ~w10059;
assign w10804 = w10802 & w10803;
assign w10805 = ~w10802 & ~w10803;
assign w10806 = ~w10804 & ~w10805;
assign w10807 = w10740 & ~w10806;
assign w10808 = ~w10740 & w10806;
assign w10809 = ~w10807 & ~w10808;
assign w10810 = ~w10061 & ~w10065;
assign w10811 = ~w10809 & w10810;
assign w10812 = w10809 & ~w10810;
assign w10813 = ~w10811 & ~w10812;
assign w10814 = pi313 & w5862;
assign w10815 = ~w10813 & ~w10814;
assign w10816 = w10813 & w10814;
assign w10817 = ~w10815 & ~w10816;
assign w10818 = ~w10070 & ~w10072;
assign w10819 = ~w10817 & w10818;
assign w10820 = w10817 & ~w10818;
assign w10821 = ~w10819 & ~w10820;
assign w10822 = ~w10739 & w10821;
assign w10823 = w10739 & ~w10821;
assign w10824 = ~w10822 & ~w10823;
assign w10825 = w10734 & ~w10824;
assign w10826 = ~w10734 & w10824;
assign w10827 = ~w10825 & ~w10826;
assign w10828 = ~w10084 & ~w10086;
assign w10829 = w10827 & w10828;
assign w10830 = ~w10827 & ~w10828;
assign w10831 = ~w10829 & ~w10830;
assign w10832 = ~w10092 & ~w10831;
assign w10833 = ~w10095 & w10832;
assign w10834 = w3710 & ~w10092;
assign w10835 = ~w10091 & w10831;
assign w10836 = ~w10834 & w10835;
assign w10837 = ~w10833 & ~w10836;
assign w10838 = pi310 & w4382;
assign w10839 = ~w10837 & w10838;
assign w10840 = ~w4382 & ~w10095;
assign w10841 = w10837 & w10840;
assign w10842 = ~w9962 & ~w10838;
assign w10843 = ~w10831 & w10842;
assign w10844 = ~w10091 & w10843;
assign w10845 = ~w10839 & ~w10844;
assign w10846 = ~w10841 & w10845;
assign w10847 = w10733 & ~w10846;
assign w10848 = ~w10733 & w10846;
assign w10849 = ~w10847 & ~w10848;
assign w10850 = ~w10097 & ~w10101;
assign w10851 = ~w10849 & w10850;
assign w10852 = w10849 & ~w10850;
assign w10853 = ~w10851 & ~w10852;
assign w10854 = (~w10105 & ~w10106) | (~w10105 & w16234) | (~w10106 & w16234);
assign w10855 = pi308 & w3304;
assign w10856 = w10854 & ~w10855;
assign w10857 = ~w10854 & w10855;
assign w10858 = ~w10856 & ~w10857;
assign w10859 = w10853 & w10858;
assign w10860 = ~w10853 & ~w10858;
assign w10861 = ~w10859 & ~w10860;
assign w10862 = w10732 & w10861;
assign w10863 = ~w10732 & ~w10861;
assign w10864 = ~w10862 & ~w10863;
assign w10865 = (~w10112 & ~w10114) | (~w10112 & w16480) | (~w10114 & w16480);
assign w10866 = w10864 & ~w10865;
assign w10867 = ~w10864 & w10865;
assign w10868 = ~w10866 & ~w10867;
assign w10869 = ~w10120 & w10868;
assign w10870 = ~w9958 & ~w10121;
assign w10871 = w10869 & ~w10870;
assign w10872 = w10120 & ~w10868;
assign w10873 = ~w10871 & ~w10872;
assign w10874 = ~w2801 & ~w10873;
assign w10875 = w10122 & w16481;
assign w10876 = ~w10121 & ~w10868;
assign w10877 = pi306 & ~w10869;
assign w10878 = ~w10876 & w10877;
assign w10879 = (w2801 & w10878) | (w2801 & w16482) | (w10878 & w16482);
assign w10880 = pi306 & w2801;
assign w10881 = w10868 & ~w10880;
assign w10882 = ~w10868 & w10880;
assign w10883 = w10870 & ~w10881;
assign w10884 = ~w10882 & w10883;
assign w10885 = ~w10879 & ~w10884;
assign w10886 = ~w10874 & w10885;
assign w10887 = pi305 & ~w2473;
assign w10888 = w10886 & w10887;
assign w10889 = ~w10886 & ~w10887;
assign w10890 = ~w10888 & ~w10889;
assign w10891 = ~w10127 & ~w10131;
assign w10892 = ~w10890 & w10891;
assign w10893 = w10890 & ~w10891;
assign w10894 = ~w10892 & ~w10893;
assign w10895 = ~w10731 & w10894;
assign w10896 = w10731 & ~w10894;
assign w10897 = ~w10895 & ~w10896;
assign w10898 = w10726 & w10897;
assign w10899 = ~w10726 & ~w10897;
assign w10900 = ~w10898 & ~w10899;
assign w10901 = w10717 & ~w10900;
assign w10902 = ~w10717 & w10900;
assign w10903 = ~w10901 & ~w10902;
assign w10904 = (~w10146 & w10150) | (~w10146 & w16483) | (w10150 & w16483);
assign w10905 = ~w10903 & w10904;
assign w10906 = w10903 & ~w10904;
assign w10907 = ~w10905 & ~w10906;
assign w10908 = ~w10716 & ~w10907;
assign w10909 = w10716 & w10907;
assign w10910 = ~w10908 & ~w10909;
assign w10911 = ~w10158 & ~w10160;
assign w10912 = w10910 & ~w10911;
assign w10913 = ~w10910 & w10911;
assign w10914 = ~w10912 & ~w10913;
assign w10915 = (w10914 & w10167) | (w10914 & w16484) | (w10167 & w16484);
assign w10916 = ~w10167 & w16485;
assign w10917 = ~w10915 & ~w10916;
assign w10918 = w10714 & w10917;
assign w10919 = ~w10714 & ~w10917;
assign w10920 = ~w10918 & ~w10919;
assign w10921 = pi299 & w855;
assign w10922 = (~w10171 & ~w10173) | (~w10171 & w15968) | (~w10173 & w15968);
assign w10923 = w10921 & ~w10922;
assign w10924 = ~w10921 & w10922;
assign w10925 = ~w10923 & ~w10924;
assign w10926 = w10920 & w10925;
assign w10927 = ~w10920 & ~w10925;
assign w10928 = ~w10926 & ~w10927;
assign w10929 = ~w10713 & w10928;
assign w10930 = w10713 & ~w10928;
assign w10931 = ~w10929 & ~w10930;
assign w10932 = w10712 & w10931;
assign w10933 = ~w10712 & ~w10931;
assign w10934 = ~w10932 & ~w10933;
assign w10935 = w10711 & w10934;
assign w10936 = ~w10711 & ~w10934;
assign w10937 = ~w10935 & ~w10936;
assign w10938 = w651 & w9446;
assign w10939 = ~w10188 & ~w10194;
assign w10940 = pi130 & ~w10939;
assign w10941 = ~w10938 & ~w10940;
assign w10942 = pi297 & ~w10941;
assign w10943 = ~w10197 & ~w10942;
assign w10944 = ~w10937 & w10943;
assign w10945 = w10937 & ~w10943;
assign w10946 = ~w10944 & ~w10945;
assign w10947 = w10183 & w10942;
assign w10948 = ~w10943 & ~w10947;
assign w10949 = ~w9947 & ~w10198;
assign w10950 = ~w10948 & w10949;
assign w10951 = ~w9948 & ~w10950;
assign w10952 = w10946 & ~w10951;
assign w10953 = ~w10946 & w10951;
assign w10954 = ~w10952 & ~w10953;
assign w10955 = w10710 & w10954;
assign w10956 = ~w10710 & ~w10954;
assign w10957 = ~w10955 & ~w10956;
assign w10958 = w10709 & w10957;
assign w10959 = ~w10709 & ~w10957;
assign w10960 = ~w10958 & ~w10959;
assign w10961 = w10705 & w10960;
assign w10962 = ~w10705 & ~w10960;
assign w10963 = ~w10961 & ~w10962;
assign w10964 = ~w10211 & ~w10693;
assign w10965 = ~pi285 & w10964;
assign w10966 = pi285 & ~w10964;
assign w10967 = ~w10965 & ~w10966;
assign w10968 = pi349 & w456;
assign w10969 = pi348 & w466;
assign w10970 = ~w10690 & ~w10969;
assign w10971 = w466 & w10690;
assign w10972 = ~w10970 & ~w10971;
assign w10973 = pi347 & ~w537;
assign w10974 = (w10973 & w10687) | (w10973 & w16235) | (w10687 & w16235);
assign w10975 = ~w10687 & w16236;
assign w10976 = ~w10974 & ~w10975;
assign w10977 = pi346 & ~w615;
assign w10978 = ~w10224 & ~w10683;
assign w10979 = w10223 & ~w10978;
assign w10980 = ~w10977 & ~w10979;
assign w10981 = ~w615 & w10979;
assign w10982 = ~w10980 & ~w10981;
assign w10983 = pi345 & ~w793;
assign w10984 = pi344 & ~w955;
assign w10985 = (~w10672 & w16613) | (~w10672 & w16614) | (w16613 & w16614);
assign w10986 = (w10672 & w16615) | (w10672 & w16616) | (w16615 & w16616);
assign w10987 = ~w10985 & ~w10986;
assign w10988 = pi343 & w1101;
assign w10989 = ~w10988 & w17700;
assign w10990 = (w10664 & w16237) | (w10664 & w16238) | (w16237 & w16238);
assign w10991 = ~w10989 & ~w10990;
assign w10992 = pi342 & w1339;
assign w10993 = (~w10233 & ~w10661) | (~w10233 & w15971) | (~w10661 & w15971);
assign w10994 = (w10661 & w16239) | (w10661 & w16240) | (w16239 & w16240);
assign w10995 = ~w10992 & w10993;
assign w10996 = ~w10994 & ~w10995;
assign w10997 = pi341 & w1602;
assign w10998 = ~w10997 & w17701;
assign w10999 = (w10658 & w16241) | (w10658 & w16242) | (w16241 & w16242);
assign w11000 = ~w10998 & ~w10999;
assign w11001 = pi340 & ~w1865;
assign w11002 = (~w10242 & ~w10655) | (~w10242 & w15973) | (~w10655 & w15973);
assign w11003 = ~w11001 & w11002;
assign w11004 = (w10655 & w16243) | (w10655 & w16244) | (w16243 & w16244);
assign w11005 = ~w11003 & ~w11004;
assign w11006 = pi337 & w2698;
assign w11007 = ~w10638 & ~w10641;
assign w11008 = ~w11006 & w11007;
assign w11009 = w11006 & ~w11007;
assign w11010 = ~w11008 & ~w11009;
assign w11011 = pi335 & ~w3568;
assign w11012 = w10260 & w10272;
assign w11013 = ~w10260 & ~w10272;
assign w11014 = ~w10262 & w10630;
assign w11015 = w10262 & ~w10630;
assign w11016 = ~w11014 & ~w11015;
assign w11017 = ~w10261 & ~w11016;
assign w11018 = (~w11013 & ~w11016) | (~w11013 & w16245) | (~w11016 & w16245);
assign w11019 = ~w11017 & w11018;
assign w11020 = ~w11012 & ~w11019;
assign w11021 = ~w11011 & w11020;
assign w11022 = w11011 & ~w11020;
assign w11023 = ~w11021 & ~w11022;
assign w11024 = pi334 & w3979;
assign w11025 = (~w11014 & ~w11016) | (~w11014 & w16246) | (~w11016 & w16246);
assign w11026 = ~w11024 & w11025;
assign w11027 = w3979 & ~w11025;
assign w11028 = ~w11026 & ~w11027;
assign w11029 = pi333 & ~w4708;
assign w11030 = w10273 & w10622;
assign w11031 = ~w10273 & ~w10622;
assign w11032 = ~w10606 & ~w10624;
assign w11033 = w10606 & w10624;
assign w11034 = ~w11032 & ~w11033;
assign w11035 = ~w10618 & w11034;
assign w11036 = w10618 & ~w11034;
assign w11037 = ~w11035 & ~w11036;
assign w11038 = ~w11031 & ~w11037;
assign w11039 = ~w11030 & ~w11038;
assign w11040 = w11029 & ~w11039;
assign w11041 = ~w11029 & w11039;
assign w11042 = ~w11040 & ~w11041;
assign w11043 = pi330 & w5714;
assign w11044 = w10596 & ~w10597;
assign w11045 = ~w11043 & w11044;
assign w11046 = w5194 & ~w5714;
assign w11047 = ~w10596 & w10597;
assign w11048 = (w5194 & w10596) | (w5194 & w10601) | (w10596 & w10601);
assign w11049 = ~w11044 & ~w11048;
assign w11050 = ~w11046 & ~w11049;
assign w11051 = w10598 & ~w11047;
assign w11052 = ~w11043 & ~w11051;
assign w11053 = ~w11050 & ~w11052;
assign w11054 = ~w11045 & ~w11053;
assign w11055 = ~w10293 & ~w10591;
assign w11056 = pi327 & w7742;
assign w11057 = (~w10582 & ~w10590) | (~w10582 & w16247) | (~w10590 & w16247);
assign w11058 = w11056 & ~w11057;
assign w11059 = ~w11056 & w11057;
assign w11060 = ~w11058 & ~w11059;
assign w11061 = w10554 & ~w10565;
assign w11062 = ~w10572 & ~w11061;
assign w11063 = ~w9782 & ~w10533;
assign w11064 = ~w10537 & w11063;
assign w11065 = w10530 & w11064;
assign w11066 = ~w10530 & ~w11064;
assign w11067 = ~w11065 & ~w11066;
assign w11068 = ~w10532 & ~w11067;
assign w11069 = w10532 & w11067;
assign w11070 = ~w11068 & ~w11069;
assign w11071 = pi323 & ~w11070;
assign w11072 = ~pi322 & ~w11071;
assign w11073 = ~w10530 & ~w10532;
assign w11074 = pi152 & pi261;
assign w11075 = (~w10513 & ~w10514) | (~w10513 & w15974) | (~w10514 & w15974);
assign w11076 = pi149 & pi264;
assign w11077 = pi148 & pi265;
assign w11078 = w10328 & ~w10500;
assign w11079 = ~w11078 & w15975;
assign w11080 = (~w11077 & w11078) | (~w11077 & w15976) | (w11078 & w15976);
assign w11081 = ~w11079 & ~w11080;
assign w11082 = pi147 & pi266;
assign w11083 = (~w10492 & ~w10494) | (~w10492 & w16486) | (~w10494 & w16486);
assign w11084 = pi146 & pi267;
assign w11085 = pi145 & pi268;
assign w11086 = (~w10485 & w10479) | (~w10485 & w15977) | (w10479 & w15977);
assign w11087 = (~w11085 & w11086) | (~w11085 & w16487) | (w11086 & w16487);
assign w11088 = ~w11086 & w16488;
assign w11089 = ~w11087 & ~w11088;
assign w11090 = pi144 & pi269;
assign w11091 = ~w10473 & ~w10477;
assign w11092 = pi143 & pi270;
assign w11093 = ~w10463 & ~w10466;
assign w11094 = ~w10453 & ~w10458;
assign w11095 = pi140 & pi273;
assign w11096 = pi139 & pi274;
assign w11097 = pi138 & pi275;
assign w11098 = pi137 & pi276;
assign w11099 = pi136 & pi277;
assign w11100 = pi135 & pi278;
assign w11101 = pi134 & pi279;
assign w11102 = pi133 & pi280;
assign w11103 = pi132 & pi281;
assign w11104 = ~w10383 & ~w10386;
assign w11105 = pi129 & pi284;
assign w11106 = pi128 & pi285;
assign w11107 = ~w11105 & ~w11106;
assign w11108 = w11105 & w11106;
assign w11109 = ~w11107 & ~w11108;
assign w11110 = ~w9591 & ~w10366;
assign w11111 = pi130 & pi283;
assign w11112 = w11110 & ~w11111;
assign w11113 = ~pi283 & w10366;
assign w11114 = pi129 & ~w10367;
assign w11115 = ~w11113 & w11114;
assign w11116 = pi130 & w11115;
assign w11117 = ~w11112 & ~w11116;
assign w11118 = w11109 & ~w11117;
assign w11119 = ~w10367 & w11109;
assign w11120 = ~w10367 & ~w11110;
assign w11121 = ~w11109 & ~w11120;
assign w11122 = ~pi130 & ~w11119;
assign w11123 = ~w11121 & w11122;
assign w11124 = ~w11111 & ~w11113;
assign w11125 = ~w11109 & ~w11115;
assign w11126 = ~w11124 & w11125;
assign w11127 = ~w11123 & ~w11126;
assign w11128 = ~w11118 & w11127;
assign w11129 = ~w10376 & ~w11128;
assign w11130 = w10362 & ~w10377;
assign w11131 = w11129 & ~w11130;
assign w11132 = pi130 & ~w10377;
assign w11133 = w11128 & w11132;
assign w11134 = ~w11131 & ~w11133;
assign w11135 = ~pi131 & w11134;
assign w11136 = w10376 & w11128;
assign w11137 = ~pi282 & ~w11129;
assign w11138 = ~w11136 & w11137;
assign w11139 = ~w11135 & ~w11138;
assign w11140 = pi131 & pi282;
assign w11141 = ~w11134 & w11140;
assign w11142 = w11139 & ~w11141;
assign w11143 = ~w11104 & w11142;
assign w11144 = w11104 & ~w11142;
assign w11145 = ~w11143 & ~w11144;
assign w11146 = w11103 & ~w11145;
assign w11147 = ~w11103 & w11145;
assign w11148 = ~w11146 & ~w11147;
assign w11149 = ~w10389 & ~w10393;
assign w11150 = w11148 & ~w11149;
assign w11151 = ~w11148 & w11149;
assign w11152 = ~w11150 & ~w11151;
assign w11153 = w11102 & w11152;
assign w11154 = ~w11102 & ~w11152;
assign w11155 = ~w11153 & ~w11154;
assign w11156 = w10399 & ~w10404;
assign w11157 = ~w10396 & ~w11156;
assign w11158 = w11155 & ~w11157;
assign w11159 = ~w11155 & w11157;
assign w11160 = ~w11158 & ~w11159;
assign w11161 = ~w11101 & ~w11160;
assign w11162 = w11101 & w11160;
assign w11163 = ~w11161 & ~w11162;
assign w11164 = w10357 & w10401;
assign w11165 = (~w11164 & w10356) | (~w11164 & w16489) | (w10356 & w16489);
assign w11166 = ~w11163 & ~w11165;
assign w11167 = w11163 & w11165;
assign w11168 = ~w11166 & ~w11167;
assign w11169 = ~w10418 & w16248;
assign w11170 = (~w11168 & w10418) | (~w11168 & w16249) | (w10418 & w16249);
assign w11171 = ~w11169 & ~w11170;
assign w11172 = w11100 & w11171;
assign w11173 = ~w11100 & ~w11171;
assign w11174 = ~w11172 & ~w11173;
assign w11175 = w10354 & ~w10422;
assign w11176 = ~w10423 & ~w11175;
assign w11177 = w11174 & ~w11176;
assign w11178 = ~w11174 & w11176;
assign w11179 = ~w11177 & ~w11178;
assign w11180 = w11099 & ~w11179;
assign w11181 = ~w11099 & w11179;
assign w11182 = ~w11180 & ~w11181;
assign w11183 = ~w11098 & w11182;
assign w11184 = w11098 & ~w11182;
assign w11185 = ~w11183 & ~w11184;
assign w11186 = (~w10430 & ~w10432) | (~w10430 & w16250) | (~w10432 & w16250);
assign w11187 = w11185 & ~w11186;
assign w11188 = ~w11185 & w11186;
assign w11189 = ~w11187 & ~w11188;
assign w11190 = ~w10437 & ~w10440;
assign w11191 = ~w10436 & ~w11190;
assign w11192 = w11189 & ~w11191;
assign w11193 = ~w11189 & w11191;
assign w11194 = ~w11192 & ~w11193;
assign w11195 = w11097 & w11194;
assign w11196 = ~w11097 & ~w11194;
assign w11197 = ~w11195 & ~w11196;
assign w11198 = w11096 & w11197;
assign w11199 = ~w11096 & ~w11197;
assign w11200 = ~w11198 & ~w11199;
assign w11201 = ~w10444 & ~w10447;
assign w11202 = w11200 & ~w11201;
assign w11203 = ~w11200 & w11201;
assign w11204 = ~w11202 & ~w11203;
assign w11205 = ~w11095 & ~w11204;
assign w11206 = w11095 & w11204;
assign w11207 = ~w11205 & ~w11206;
assign w11208 = ~w10347 & ~w10450;
assign w11209 = ~w11207 & w11208;
assign w11210 = w11207 & ~w11208;
assign w11211 = ~w11209 & ~w11210;
assign w11212 = w11094 & w11211;
assign w11213 = ~w11094 & ~w11211;
assign w11214 = ~w11212 & ~w11213;
assign w11215 = pi142 & pi271;
assign w11216 = pi141 & pi272;
assign w11217 = w11215 & ~w11216;
assign w11218 = ~w11215 & w11216;
assign w11219 = ~w11217 & ~w11218;
assign w11220 = w11214 & w11219;
assign w11221 = ~w11214 & ~w11219;
assign w11222 = ~w11220 & ~w11221;
assign w11223 = ~w11093 & ~w11222;
assign w11224 = w11093 & w11222;
assign w11225 = ~w11223 & ~w11224;
assign w11226 = w11092 & w11225;
assign w11227 = ~w11092 & ~w11225;
assign w11228 = ~w11226 & ~w11227;
assign w11229 = ~w10339 & ~w10469;
assign w11230 = ~w11228 & w11229;
assign w11231 = w11228 & ~w11229;
assign w11232 = ~w11230 & ~w11231;
assign w11233 = ~w11091 & ~w11232;
assign w11234 = w11091 & w11232;
assign w11235 = ~w11233 & ~w11234;
assign w11236 = w11090 & w11235;
assign w11237 = ~w11090 & ~w11235;
assign w11238 = ~w11236 & ~w11237;
assign w11239 = ~w11089 & ~w11238;
assign w11240 = w11089 & w11238;
assign w11241 = ~w11239 & ~w11240;
assign w11242 = w11084 & w11241;
assign w11243 = ~w11084 & ~w11241;
assign w11244 = ~w11242 & ~w11243;
assign w11245 = (~w10333 & ~w10335) | (~w10333 & w16490) | (~w10335 & w16490);
assign w11246 = ~w11244 & w11245;
assign w11247 = w11244 & ~w11245;
assign w11248 = ~w11246 & ~w11247;
assign w11249 = w11083 & ~w11248;
assign w11250 = ~w11083 & w11248;
assign w11251 = ~w11249 & ~w11250;
assign w11252 = ~w11082 & w11251;
assign w11253 = w11082 & ~w11251;
assign w11254 = ~w11252 & ~w11253;
assign w11255 = w11081 & ~w11254;
assign w11256 = ~w11081 & w11254;
assign w11257 = ~w11255 & ~w11256;
assign w11258 = ~w11076 & ~w11257;
assign w11259 = w11076 & w11257;
assign w11260 = ~w11258 & ~w11259;
assign w11261 = ~w10325 & ~w10506;
assign w11262 = w11260 & ~w11261;
assign w11263 = ~w11260 & w11261;
assign w11264 = ~w11262 & ~w11263;
assign w11265 = (~w10319 & ~w10320) | (~w10319 & w15978) | (~w10320 & w15978);
assign w11266 = pi151 & pi262;
assign w11267 = pi150 & pi263;
assign w11268 = w11266 & ~w11267;
assign w11269 = ~w11266 & w11267;
assign w11270 = ~w11268 & ~w11269;
assign w11271 = (w15978 & w16251) | (w15978 & w16252) | (w16251 & w16252);
assign w11272 = (~w15978 & w16253) | (~w15978 & w16254) | (w16253 & w16254);
assign w11273 = ~w11271 & ~w11272;
assign w11274 = w11264 & w11273;
assign w11275 = ~w11264 & ~w11273;
assign w11276 = ~w11274 & ~w11275;
assign w11277 = w11075 & w11276;
assign w11278 = ~w11075 & ~w11276;
assign w11279 = ~w11277 & ~w11278;
assign w11280 = ~w11074 & w11279;
assign w11281 = w11074 & ~w11279;
assign w11282 = ~w11280 & ~w11281;
assign w11283 = ~w10522 & ~w10525;
assign w11284 = w11282 & w11283;
assign w11285 = ~w11282 & ~w11283;
assign w11286 = ~w11284 & ~w11285;
assign w11287 = (w10303 & w10527) | (w10303 & w16491) | (w10527 & w16491);
assign w11288 = pi153 & pi259;
assign w11289 = w10527 & w11288;
assign w11290 = ~w11287 & ~w11289;
assign w11291 = w11286 & w11290;
assign w11292 = ~w11286 & ~w11290;
assign w11293 = ~w11291 & ~w11292;
assign w11294 = w10304 & w10530;
assign w11295 = pi154 & pi259;
assign w11296 = pi153 & pi260;
assign w11297 = pi155 & pi258;
assign w11298 = w11296 & ~w11297;
assign w11299 = ~w11296 & w11297;
assign w11300 = ~w11298 & ~w11299;
assign w11301 = w11295 & ~w11300;
assign w11302 = ~w11295 & w11300;
assign w11303 = ~w11301 & ~w11302;
assign w11304 = w10530 & w16492;
assign w11305 = (w11303 & ~w10530) | (w11303 & w16493) | (~w10530 & w16493);
assign w11306 = ~w11304 & ~w11305;
assign w11307 = w11293 & w11306;
assign w11308 = ~w11293 & ~w11306;
assign w11309 = ~w11307 & ~w11308;
assign w11310 = ~w11064 & w11309;
assign w11311 = w11309 & w15979;
assign w11312 = w10530 & w10543;
assign w11313 = ~w11069 & ~w11312;
assign w11314 = ~w11309 & ~w11313;
assign w11315 = ~w11311 & ~w11314;
assign w11316 = w10296 & ~w11315;
assign w11317 = w11065 & w11309;
assign w11318 = ~w11065 & ~w11309;
assign w11319 = ~w11317 & ~w11318;
assign w11320 = ~w11068 & ~w11073;
assign w11321 = ~w11319 & w11320;
assign w11322 = ~w10530 & w11064;
assign w11323 = ~w10543 & ~w11322;
assign w11324 = (~w11071 & w11309) | (~w11071 & w16255) | (w11309 & w16255);
assign w11325 = ~w11311 & w11324;
assign w11326 = ~w11321 & w11325;
assign w11327 = (~w11072 & w11315) | (~w11072 & w16256) | (w11315 & w16256);
assign w11328 = ~w11326 & w11327;
assign w11329 = pi324 & ~w9784;
assign w11330 = ~w10552 & ~w10558;
assign w11331 = (~w10557 & ~w11330) | (~w10557 & w16257) | (~w11330 & w16257);
assign w11332 = w11329 & w11331;
assign w11333 = ~w11329 & ~w11331;
assign w11334 = ~w11332 & ~w11333;
assign w11335 = pi325 & w8814;
assign w11336 = ~w10548 & ~w10551;
assign w11337 = w11335 & ~w11336;
assign w11338 = ~w11335 & w11336;
assign w11339 = ~w11337 & ~w11338;
assign w11340 = w11334 & ~w11339;
assign w11341 = ~w11334 & w11339;
assign w11342 = ~w11340 & ~w11341;
assign w11343 = w11328 & w11342;
assign w11344 = ~w11328 & ~w11342;
assign w11345 = ~w11343 & ~w11344;
assign w11346 = ~w11062 & w11345;
assign w11347 = w11062 & ~w11345;
assign w11348 = ~w11346 & ~w11347;
assign w11349 = pi326 & ~w8367;
assign w11350 = (~w10578 & ~w10574) | (~w10578 & w16494) | (~w10574 & w16494);
assign w11351 = ~w11349 & w11350;
assign w11352 = w11349 & ~w11350;
assign w11353 = ~w11351 & ~w11352;
assign w11354 = w11348 & w11353;
assign w11355 = ~w11348 & ~w11353;
assign w11356 = ~w11354 & ~w11355;
assign w11357 = w11060 & w11356;
assign w11358 = ~w11060 & ~w11356;
assign w11359 = ~w11357 & ~w11358;
assign w11360 = w11055 & ~w11359;
assign w11361 = ~w11055 & w11359;
assign w11362 = ~w11360 & ~w11361;
assign w11363 = pi328 & ~w7108;
assign w11364 = pi329 & w6283;
assign w11365 = ~w10594 & w16258;
assign w11366 = (w11364 & w10594) | (w11364 & w16259) | (w10594 & w16259);
assign w11367 = ~w11365 & ~w11366;
assign w11368 = w11363 & ~w11367;
assign w11369 = ~w11363 & w11367;
assign w11370 = ~w11368 & ~w11369;
assign w11371 = w11362 & w11370;
assign w11372 = ~w11362 & ~w11370;
assign w11373 = ~w11371 & ~w11372;
assign w11374 = ~w11054 & ~w11373;
assign w11375 = w11054 & w11373;
assign w11376 = ~w11374 & ~w11375;
assign w11377 = pi331 & w5194;
assign w11378 = ~w10610 & ~w11033;
assign w11379 = ~w11032 & ~w11378;
assign w11380 = w11377 & w11379;
assign w11381 = ~w11377 & ~w11379;
assign w11382 = ~w11380 & ~w11381;
assign w11383 = ~w11376 & ~w11382;
assign w11384 = w11376 & w11382;
assign w11385 = ~w11383 & ~w11384;
assign w11386 = pi332 & ~w4854;
assign w11387 = ~pi331 & w11386;
assign w11388 = ~w10613 & w11387;
assign w11389 = ~w11034 & w11388;
assign w11390 = ~w4854 & ~w10614;
assign w11391 = ~w10613 & ~w11386;
assign w11392 = ~w11390 & ~w11391;
assign w11393 = w10615 & ~w11388;
assign w11394 = w11034 & w11393;
assign w11395 = ~w11389 & ~w11392;
assign w11396 = ~w11394 & w11395;
assign w11397 = w11385 & w11396;
assign w11398 = ~w11385 & ~w11396;
assign w11399 = ~w11397 & ~w11398;
assign w11400 = w11042 & ~w11399;
assign w11401 = ~w11042 & w11399;
assign w11402 = ~w11400 & ~w11401;
assign w11403 = w11028 & ~w11402;
assign w11404 = ~w11028 & w11402;
assign w11405 = ~w11403 & ~w11404;
assign w11406 = w11023 & ~w11405;
assign w11407 = ~w11023 & w11405;
assign w11408 = ~w11406 & ~w11407;
assign w11409 = pi336 & ~w3183;
assign w11410 = ~w10258 & ~w10636;
assign w11411 = ~w10257 & ~w11410;
assign w11412 = w11409 & ~w11411;
assign w11413 = ~w11409 & w11411;
assign w11414 = ~w11412 & ~w11413;
assign w11415 = w11408 & w11414;
assign w11416 = ~w11408 & ~w11414;
assign w11417 = ~w11415 & ~w11416;
assign w11418 = w11010 & w11417;
assign w11419 = ~w11010 & ~w11417;
assign w11420 = ~w11418 & ~w11419;
assign w11421 = (~w10248 & w10652) | (~w10248 & w15980) | (w10652 & w15980);
assign w11422 = pi338 & ~w2373;
assign w11423 = ~w10644 & w17702;
assign w11424 = ~w11422 & ~w11423;
assign w11425 = (w9876 & w16495) | (w9876 & w16496) | (w16495 & w16496);
assign w11426 = w11422 & ~w11425;
assign w11427 = pi337 & w11426;
assign w11428 = ~w11424 & ~w11427;
assign w11429 = w10639 & ~w11428;
assign w11430 = ~w11422 & ~w11425;
assign w11431 = ~w2373 & ~w11423;
assign w11432 = ~w11430 & ~w11431;
assign w11433 = ~pi337 & w11426;
assign w11434 = (~w11432 & w10639) | (~w11432 & w16261) | (w10639 & w16261);
assign w11435 = ~w11429 & w11434;
assign w11436 = pi339 & ~w2170;
assign w11437 = w11435 & ~w11436;
assign w11438 = ~w11435 & w11436;
assign w11439 = ~w11437 & ~w11438;
assign w11440 = w11421 & ~w11439;
assign w11441 = ~w11421 & w11439;
assign w11442 = ~w11440 & ~w11441;
assign w11443 = w11420 & w11442;
assign w11444 = ~w11420 & ~w11442;
assign w11445 = ~w11443 & ~w11444;
assign w11446 = w11005 & w11445;
assign w11447 = ~w11005 & ~w11445;
assign w11448 = ~w11446 & ~w11447;
assign w11449 = w11000 & w11448;
assign w11450 = ~w11000 & ~w11448;
assign w11451 = ~w11449 & ~w11450;
assign w11452 = w10996 & w11451;
assign w11453 = ~w10996 & ~w11451;
assign w11454 = ~w11452 & ~w11453;
assign w11455 = w10991 & w11454;
assign w11456 = ~w10991 & ~w11454;
assign w11457 = ~w11455 & ~w11456;
assign w11458 = w10987 & w11457;
assign w11459 = ~w10987 & ~w11457;
assign w11460 = ~w11458 & ~w11459;
assign w11461 = ~w10227 & ~w10681;
assign w11462 = w11460 & ~w11461;
assign w11463 = ~w11460 & w11461;
assign w11464 = ~w11462 & ~w11463;
assign w11465 = w10983 & w11464;
assign w11466 = ~w10983 & ~w11464;
assign w11467 = ~w11465 & ~w11466;
assign w11468 = w10982 & w11467;
assign w11469 = ~w10982 & ~w11467;
assign w11470 = ~w11468 & ~w11469;
assign w11471 = w10976 & w11470;
assign w11472 = ~w10976 & ~w11470;
assign w11473 = ~w11471 & ~w11472;
assign w11474 = w10972 & w11473;
assign w11475 = ~w10972 & ~w11473;
assign w11476 = ~w11474 & ~w11475;
assign w11477 = ~w10968 & ~w11476;
assign w11478 = w10968 & w11476;
assign w11479 = ~w11477 & ~w11478;
assign w11480 = w10967 & w11479;
assign w11481 = ~w10967 & ~w11479;
assign w11482 = ~w11480 & ~w11481;
assign w11483 = w10963 & w11482;
assign w11484 = ~w10963 & ~w11482;
assign w11485 = ~w11483 & ~w11484;
assign w11486 = ~w10207 & ~w10696;
assign w11487 = ~w11485 & ~w11486;
assign w11488 = w11485 & w11486;
assign w11489 = ~w135 & ~w11487;
assign w11490 = ~w11488 & w11489;
assign w11491 = pi161 & ~w203;
assign w11492 = ~w11490 & w11491;
assign w11493 = ~pi160 & ~w10704;
assign w11494 = ~w11492 & w11493;
assign w11495 = ~pi092 & ~pi161;
assign w11496 = ~w11484 & ~w11488;
assign w11497 = pi128 & pi293;
assign w11498 = pi294 & w464;
assign w11499 = (~w11498 & ~w10960) | (~w11498 & w16262) | (~w10960 & w16262);
assign w11500 = w10960 & w16263;
assign w11501 = ~w11499 & ~w11500;
assign w11502 = pi295 & ~w653;
assign w11503 = (~w10706 & ~w10957) | (~w10706 & w16264) | (~w10957 & w16264);
assign w11504 = ~w11502 & w11503;
assign w11505 = w11502 & ~w11503;
assign w11506 = ~w11504 & ~w11505;
assign w11507 = pi297 & w698;
assign w11508 = (~w10935 & ~w10937) | (~w10935 & w16265) | (~w10937 & w16265);
assign w11509 = (~w10929 & ~w10931) | (~w10929 & w16266) | (~w10931 & w16266);
assign w11510 = pi299 & w1159;
assign w11511 = pi301 & w1420;
assign w11512 = pi302 & w1693;
assign w11513 = pi303 & w1954;
assign w11514 = ~w10718 & ~w10897;
assign w11515 = w10718 & w10897;
assign w11516 = ~w10140 & ~w10143;
assign w11517 = ~w11515 & w11516;
assign w11518 = ~w11514 & ~w11517;
assign w11519 = w11513 & w11518;
assign w11520 = ~w11513 & ~w11518;
assign w11521 = ~w11519 & ~w11520;
assign w11522 = pi304 & ~w2473;
assign w11523 = pi305 & w2801;
assign w11524 = pi306 & w2925;
assign w11525 = pi307 & w3304;
assign w11526 = pi308 & w3710;
assign w11527 = pi309 & w4382;
assign w11528 = ~w10847 & ~w10852;
assign w11529 = pi310 & w4539;
assign w11530 = pi311 & w5316;
assign w11531 = pi312 & w5862;
assign w11532 = pi313 & w6437;
assign w11533 = pi314 & w6652;
assign w11534 = ~w10801 & ~w10804;
assign w11535 = pi315 & w7268;
assign w11536 = pi316 & w7909;
assign w11537 = pi317 & w9022;
assign w11538 = ~w10780 & ~w10783;
assign w11539 = pi319 & w9992;
assign w11540 = ~pi155 & ~pi156;
assign w11541 = pi155 & pi156;
assign w11542 = ~w11540 & ~w11541;
assign w11543 = pi154 & w11542;
assign w11544 = ~w10747 & w11543;
assign w11545 = pi156 & w11543;
assign w11546 = ~pi156 & w10748;
assign w11547 = pi153 & ~w11545;
assign w11548 = ~w11546 & w11547;
assign w11549 = w9986 & w11540;
assign w11550 = ~pi154 & w11541;
assign w11551 = ~pi153 & ~w11550;
assign w11552 = ~w11549 & w11551;
assign w11553 = ~w11548 & ~w11552;
assign w11554 = ~pi154 & ~w11542;
assign w11555 = ~w10748 & w11554;
assign w11556 = ~w11544 & ~w11555;
assign w11557 = ~w11553 & w11556;
assign w11558 = pi321 & w11557;
assign w11559 = w9992 & ~w10766;
assign w11560 = ~w10763 & ~w11559;
assign w11561 = ~w10753 & w11560;
assign w11562 = pi320 & ~w11560;
assign w11563 = w10753 & w11562;
assign w11564 = pi320 & ~w11561;
assign w11565 = ~w11563 & w11564;
assign w11566 = ~w11558 & w11565;
assign w11567 = w11558 & ~w11565;
assign w11568 = ~w11566 & ~w11567;
assign w11569 = ~w11539 & w11568;
assign w11570 = w11539 & ~w11568;
assign w11571 = ~w11569 & ~w11570;
assign w11572 = pi319 & ~w10774;
assign w11573 = ~w11571 & w11572;
assign w11574 = ~w10774 & ~w10777;
assign w11575 = ~w11570 & ~w11574;
assign w11576 = ~w11569 & w11575;
assign w11577 = ~pi318 & ~w11573;
assign w11578 = ~w11576 & w11577;
assign w11579 = w10773 & ~w11571;
assign w11580 = ~w10773 & w11571;
assign w11581 = ~w9270 & ~w11579;
assign w11582 = ~w11580 & w11581;
assign w11583 = ~w11578 & ~w11582;
assign w11584 = w11571 & ~w11572;
assign w11585 = ~w11573 & ~w11584;
assign w11586 = pi318 & w9270;
assign w11587 = ~w11585 & w11586;
assign w11588 = w11583 & ~w11587;
assign w11589 = w11538 & ~w11588;
assign w11590 = ~w11538 & w11588;
assign w11591 = ~w11589 & ~w11590;
assign w11592 = ~w11537 & w11591;
assign w11593 = w11537 & ~w11591;
assign w11594 = ~w11592 & ~w11593;
assign w11595 = ~w10785 & ~w10789;
assign w11596 = w11594 & w11595;
assign w11597 = ~w11594 & ~w11595;
assign w11598 = ~w11596 & ~w11597;
assign w11599 = w11536 & ~w11598;
assign w11600 = ~w11536 & w11598;
assign w11601 = ~w11599 & ~w11600;
assign w11602 = ~w10794 & ~w10797;
assign w11603 = ~w11601 & w11602;
assign w11604 = w11601 & ~w11602;
assign w11605 = ~w11603 & ~w11604;
assign w11606 = ~w11535 & ~w11605;
assign w11607 = w11535 & w11605;
assign w11608 = ~w11606 & ~w11607;
assign w11609 = w11534 & w11608;
assign w11610 = ~w11534 & ~w11608;
assign w11611 = ~w11609 & ~w11610;
assign w11612 = w11533 & w11611;
assign w11613 = ~w11533 & ~w11611;
assign w11614 = ~w11612 & ~w11613;
assign w11615 = ~w10807 & ~w10812;
assign w11616 = w11614 & ~w11615;
assign w11617 = ~w11614 & w11615;
assign w11618 = ~w11616 & ~w11617;
assign w11619 = ~w11532 & ~w11618;
assign w11620 = w11532 & w11618;
assign w11621 = ~w11619 & ~w11620;
assign w11622 = ~w10816 & ~w10820;
assign w11623 = w11621 & ~w11622;
assign w11624 = ~w11621 & w11622;
assign w11625 = ~w11623 & ~w11624;
assign w11626 = ~w11531 & ~w11625;
assign w11627 = w11531 & w11625;
assign w11628 = ~w11626 & ~w11627;
assign w11629 = ~w10738 & ~w10823;
assign w11630 = w11628 & ~w11629;
assign w11631 = ~w11628 & w11629;
assign w11632 = ~w11630 & ~w11631;
assign w11633 = ~w10826 & ~w10829;
assign w11634 = w11632 & ~w11633;
assign w11635 = ~w11632 & w11633;
assign w11636 = ~w11634 & ~w11635;
assign w11637 = w11530 & w11636;
assign w11638 = ~w11530 & ~w11636;
assign w11639 = ~w11637 & ~w11638;
assign w11640 = ~w10833 & ~w10838;
assign w11641 = ~w10836 & ~w11640;
assign w11642 = w11639 & w11641;
assign w11643 = ~w11639 & ~w11641;
assign w11644 = ~w11642 & ~w11643;
assign w11645 = w11529 & ~w11644;
assign w11646 = ~w11529 & w11644;
assign w11647 = ~w11645 & ~w11646;
assign w11648 = ~w11528 & ~w11647;
assign w11649 = w11528 & w11647;
assign w11650 = ~w11648 & ~w11649;
assign w11651 = w11527 & ~w11650;
assign w11652 = ~w11527 & w11650;
assign w11653 = ~w11651 & ~w11652;
assign w11654 = ~w11526 & w11653;
assign w11655 = w11526 & ~w11653;
assign w11656 = ~w11654 & ~w11655;
assign w11657 = ~w10857 & ~w10859;
assign w11658 = w11656 & ~w11657;
assign w11659 = ~w11656 & w11657;
assign w11660 = ~w11658 & ~w11659;
assign w11661 = ~w10862 & ~w10866;
assign w11662 = w11660 & ~w11661;
assign w11663 = ~w11660 & w11661;
assign w11664 = ~w11662 & ~w11663;
assign w11665 = w11525 & w11664;
assign w11666 = ~w11525 & ~w11664;
assign w11667 = ~w11665 & ~w11666;
assign w11668 = w10880 & ~w10885;
assign w11669 = ~w10871 & ~w11668;
assign w11670 = ~w11667 & w11669;
assign w11671 = w11667 & ~w11669;
assign w11672 = ~w11670 & ~w11671;
assign w11673 = w11524 & w11672;
assign w11674 = ~w11524 & ~w11672;
assign w11675 = ~w11673 & ~w11674;
assign w11676 = ~w11523 & ~w11675;
assign w11677 = w11523 & w11675;
assign w11678 = ~w11676 & ~w11677;
assign w11679 = ~w10889 & ~w10893;
assign w11680 = w11678 & w11679;
assign w11681 = ~w11678 & ~w11679;
assign w11682 = ~w11680 & ~w11681;
assign w11683 = ~w11522 & ~w11682;
assign w11684 = w11522 & w11682;
assign w11685 = ~w11683 & ~w11684;
assign w11686 = ~w10729 & ~w10896;
assign w11687 = ~w11685 & w11686;
assign w11688 = w11685 & ~w11686;
assign w11689 = ~w11687 & ~w11688;
assign w11690 = ~w11521 & ~w11689;
assign w11691 = w11521 & w11689;
assign w11692 = ~w11690 & ~w11691;
assign w11693 = ~w10901 & ~w10906;
assign w11694 = w11692 & ~w11693;
assign w11695 = ~w11692 & w11693;
assign w11696 = ~w11694 & ~w11695;
assign w11697 = w11512 & ~w11696;
assign w11698 = ~w11512 & w11696;
assign w11699 = ~w11697 & ~w11698;
assign w11700 = w11511 & ~w11699;
assign w11701 = ~w11511 & w11699;
assign w11702 = ~w11700 & ~w11701;
assign w11703 = ~w10909 & ~w10912;
assign w11704 = ~w11702 & w11703;
assign w11705 = w11702 & ~w11703;
assign w11706 = ~w11704 & ~w11705;
assign w11707 = pi300 & w1220;
assign w11708 = ~w10715 & w16267;
assign w11709 = ~w1220 & w10714;
assign w11710 = (w11709 & ~w10715) | (w11709 & w16268) | (~w10715 & w16268);
assign w11711 = (w1159 & ~w10715) | (w1159 & w16269) | (~w10715 & w16269);
assign w11712 = (w11707 & w10715) | (w11707 & w16270) | (w10715 & w16270);
assign w11713 = ~w11711 & w11712;
assign w11714 = ~w11708 & ~w11710;
assign w11715 = ~w11713 & w11714;
assign w11716 = w11706 & w11715;
assign w11717 = ~w11706 & ~w11715;
assign w11718 = ~w11716 & ~w11717;
assign w11719 = (~w10923 & ~w10925) | (~w10923 & w16271) | (~w10925 & w16271);
assign w11720 = w11718 & w11719;
assign w11721 = ~w11718 & ~w11719;
assign w11722 = ~w11720 & ~w11721;
assign w11723 = w11510 & ~w11722;
assign w11724 = ~w11510 & w11722;
assign w11725 = ~w11723 & ~w11724;
assign w11726 = ~w11509 & ~w11725;
assign w11727 = w11509 & w11725;
assign w11728 = ~w11726 & ~w11727;
assign w11729 = pi298 & w855;
assign w11730 = ~w11728 & w11729;
assign w11731 = w11728 & ~w11729;
assign w11732 = ~w11730 & ~w11731;
assign w11733 = ~w11508 & ~w11732;
assign w11734 = w11508 & w11732;
assign w11735 = ~w11733 & ~w11734;
assign w11736 = w11507 & w11735;
assign w11737 = ~w11507 & ~w11735;
assign w11738 = ~w11736 & ~w11737;
assign w11739 = pi296 & w709;
assign w11740 = (~w10952 & ~w10954) | (~w10952 & w16272) | (~w10954 & w16272);
assign w11741 = w11739 & ~w11740;
assign w11742 = ~w11739 & w11740;
assign w11743 = ~w11741 & ~w11742;
assign w11744 = w11738 & w11743;
assign w11745 = ~w11738 & ~w11743;
assign w11746 = ~w11744 & ~w11745;
assign w11747 = ~w11506 & w11746;
assign w11748 = w11506 & ~w11746;
assign w11749 = ~w11747 & ~w11748;
assign w11750 = w11501 & ~w11749;
assign w11751 = ~w11501 & w11749;
assign w11752 = ~w11750 & ~w11751;
assign w11753 = w11497 & w11752;
assign w11754 = ~w11497 & ~w11752;
assign w11755 = ~w11753 & ~w11754;
assign w11756 = w11496 & w11755;
assign w11757 = ~w11496 & ~w11755;
assign w11758 = ~w11756 & ~w11757;
assign w11759 = pi350 & w456;
assign w11760 = pi348 & ~w537;
assign w11761 = (~w10971 & ~w11473) | (~w10971 & w16273) | (~w11473 & w16273);
assign w11762 = w11760 & ~w11761;
assign w11763 = ~w11760 & w11761;
assign w11764 = ~w11762 & ~w11763;
assign w11765 = pi345 & ~w955;
assign w11766 = ~pi346 & w10983;
assign w11767 = (w10983 & ~w10979) | (w10983 & w16274) | (~w10979 & w16274);
assign w11768 = pi346 & ~w793;
assign w11769 = (~w11768 & w10979) | (~w11768 & w16275) | (w10979 & w16275);
assign w11770 = ~w11767 & ~w11769;
assign w11771 = w11464 & ~w11766;
assign w11772 = ~w11770 & w11771;
assign w11773 = w10979 & w16276;
assign w11774 = ~w10979 & w16277;
assign w11775 = ~pi345 & w11768;
assign w11776 = (w11775 & ~w10979) | (w11775 & w16278) | (~w10979 & w16278);
assign w11777 = ~w11464 & w11776;
assign w11778 = ~w11773 & ~w11774;
assign w11779 = ~w11777 & w11778;
assign w11780 = ~w11772 & w11779;
assign w11781 = ~w11765 & w11780;
assign w11782 = w11765 & ~w11780;
assign w11783 = ~w11781 & ~w11782;
assign w11784 = pi347 & ~w615;
assign w11785 = ~w1339 & ~w11451;
assign w11786 = w1339 & w11451;
assign w11787 = w10993 & ~w11786;
assign w11788 = pi342 & w1602;
assign w11789 = ~w11785 & w11788;
assign w11790 = ~w11787 & w11789;
assign w11791 = ~w10994 & ~w11788;
assign w11792 = ~w11452 & w11791;
assign w11793 = ~w11790 & ~w11792;
assign w11794 = ~w11003 & w11445;
assign w11795 = pi340 & ~w2170;
assign w11796 = w11794 & ~w11795;
assign w11797 = w1865 & w11002;
assign w11798 = w11445 & ~w11797;
assign w11799 = ~w11004 & ~w11798;
assign w11800 = ~w2170 & ~w11799;
assign w11801 = ~w11004 & ~w11795;
assign w11802 = pi340 & ~w11801;
assign w11803 = ~w11800 & w11802;
assign w11804 = ~w11796 & ~w11803;
assign w11805 = ~w11421 & w11436;
assign w11806 = w11421 & ~w11436;
assign w11807 = w11420 & ~w11435;
assign w11808 = ~w11420 & w11435;
assign w11809 = (~w11806 & ~w11420) | (~w11806 & w16279) | (~w11420 & w16279);
assign w11810 = ~w11808 & w11809;
assign w11811 = ~w11805 & ~w11810;
assign w11812 = ~w11804 & w11811;
assign w11813 = w11804 & ~w11811;
assign w11814 = ~w11812 & ~w11813;
assign w11815 = pi341 & ~w1865;
assign w11816 = ~w10999 & ~w11449;
assign w11817 = ~w11815 & w11816;
assign w11818 = w11815 & ~w11816;
assign w11819 = ~w11817 & ~w11818;
assign w11820 = pi339 & ~w2373;
assign w11821 = ~w10642 & ~w11425;
assign w11822 = w11431 & ~w11821;
assign w11823 = ~w2698 & w11822;
assign w11824 = pi338 & w2698;
assign w11825 = ~w11822 & w11824;
assign w11826 = ~w11823 & ~w11825;
assign w11827 = w11420 & w16280;
assign w11828 = (w11826 & ~w11420) | (w11826 & w16281) | (~w11420 & w16281);
assign w11829 = ~w11827 & ~w11828;
assign w11830 = ~w11408 & w11411;
assign w11831 = ~w11408 & w16282;
assign w11832 = w3183 & ~w3568;
assign w11833 = w11411 & w11832;
assign w11834 = ~w3568 & ~w11412;
assign w11835 = ~w11408 & w11834;
assign w11836 = ~w7497 & ~w11833;
assign w11837 = ~w11835 & w11836;
assign w11838 = pi336 & ~w11831;
assign w11839 = ~w11837 & w11838;
assign w11840 = pi337 & ~w3183;
assign w11841 = ~w11839 & w11840;
assign w11842 = w11408 & ~w11411;
assign w11843 = pi336 & ~w3568;
assign w11844 = w11842 & ~w11843;
assign w11845 = ~w11839 & ~w11844;
assign w11846 = ~w11840 & ~w11845;
assign w11847 = ~w11841 & ~w11846;
assign w11848 = w11829 & w11847;
assign w11849 = ~w11829 & ~w11847;
assign w11850 = ~w11848 & ~w11849;
assign w11851 = pi335 & w3979;
assign w11852 = ~w11022 & ~w11406;
assign w11853 = ~w11851 & w11852;
assign w11854 = w11851 & ~w11852;
assign w11855 = ~w11853 & ~w11854;
assign w11856 = pi333 & ~w4854;
assign w11857 = pi332 & w5194;
assign w11858 = ~w10614 & w11037;
assign w11859 = ~w10613 & ~w11858;
assign w11860 = ~w11386 & w11859;
assign w11861 = w11386 & ~w11859;
assign w11862 = (~w11860 & w11385) | (~w11860 & w16283) | (w11385 & w16283);
assign w11863 = w11857 & w11862;
assign w11864 = ~w11857 & ~w11862;
assign w11865 = ~w11863 & ~w11864;
assign w11866 = ~w11380 & ~w11384;
assign w11867 = ~w11865 & w11866;
assign w11868 = w11865 & ~w11866;
assign w11869 = ~w11867 & ~w11868;
assign w11870 = pi328 & w7742;
assign w11871 = ~w11361 & ~w11363;
assign w11872 = ~w11360 & ~w11871;
assign w11873 = w11335 & ~w11345;
assign w11874 = ~w11346 & ~w11873;
assign w11875 = ~w11068 & w11319;
assign w11876 = ~w11066 & ~w11309;
assign w11877 = ~w10532 & ~w11310;
assign w11878 = ~w11876 & w11877;
assign w11879 = ~w11875 & ~w11878;
assign w11880 = pi323 & w11879;
assign w11881 = ~w10530 & ~w11311;
assign w11882 = w10532 & ~w10533;
assign w11883 = ~w11309 & w11882;
assign w11884 = ~w11881 & ~w11883;
assign w11885 = pi153 & pi261;
assign w11886 = (w11296 & ~w11286) | (w11296 & w15981) | (~w11286 & w15981);
assign w11887 = ~w11292 & ~w11886;
assign w11888 = w11885 & ~w11887;
assign w11889 = ~w11885 & w11887;
assign w11890 = ~w11888 & ~w11889;
assign w11891 = pi152 & pi262;
assign w11892 = (~w11280 & ~w11282) | (~w11280 & w16284) | (~w11282 & w16284);
assign w11893 = ~w11891 & ~w11892;
assign w11894 = w11891 & w11892;
assign w11895 = ~w11893 & ~w11894;
assign w11896 = pi150 & pi264;
assign w11897 = (~w11258 & ~w11260) | (~w11258 & w16285) | (~w11260 & w16285);
assign w11898 = pi147 & pi267;
assign w11899 = pi146 & pi268;
assign w11900 = (w11245 & ~w11241) | (w11245 & w15982) | (~w11241 & w15982);
assign w11901 = ~w11900 & w17613;
assign w11902 = (~w11899 & w11900) | (~w11899 & w17614) | (w11900 & w17614);
assign w11903 = ~w11901 & ~w11902;
assign w11904 = pi145 & pi269;
assign w11905 = pi144 & pi270;
assign w11906 = pi143 & pi271;
assign w11907 = (w11229 & ~w11225) | (w11229 & w15983) | (~w11225 & w15983);
assign w11908 = ~w11227 & ~w11907;
assign w11909 = w11906 & w11908;
assign w11910 = ~w11906 & ~w11908;
assign w11911 = ~w11909 & ~w11910;
assign w11912 = pi142 & pi272;
assign w11913 = pi141 & pi273;
assign w11914 = pi139 & pi275;
assign w11915 = (~w11198 & ~w11200) | (~w11198 & w16286) | (~w11200 & w16286);
assign w11916 = pi138 & pi276;
assign w11917 = pi137 & pi277;
assign w11918 = (~w11184 & ~w11185) | (~w11184 & w16287) | (~w11185 & w16287);
assign w11919 = ~w11917 & w11918;
assign w11920 = w11917 & ~w11918;
assign w11921 = ~w11919 & ~w11920;
assign w11922 = pi135 & pi279;
assign w11923 = pi134 & pi280;
assign w11924 = ~w11161 & ~w11167;
assign w11925 = pi133 & pi281;
assign w11926 = pi132 & pi282;
assign w11927 = pi131 & pi283;
assign w11928 = w11139 & ~w11143;
assign w11929 = ~w11927 & ~w11928;
assign w11930 = w11927 & w11928;
assign w11931 = ~w11929 & ~w11930;
assign w11932 = pi130 & pi284;
assign w11933 = w11109 & w11120;
assign w11934 = ~w11121 & ~w11933;
assign w11935 = ~w11111 & ~w11934;
assign w11936 = w11111 & w11934;
assign w11937 = ~w10376 & ~w11936;
assign w11938 = ~w11130 & w11937;
assign w11939 = ~w11935 & ~w11938;
assign w11940 = ~w11932 & ~w11939;
assign w11941 = w11932 & w11939;
assign w11942 = ~w11940 & ~w11941;
assign w11943 = pi129 & pi285;
assign w11944 = pi128 & pi286;
assign w11945 = ~w11108 & ~w11933;
assign w11946 = w11944 & ~w11945;
assign w11947 = ~w11944 & w11945;
assign w11948 = ~w11946 & ~w11947;
assign w11949 = w11943 & ~w11948;
assign w11950 = ~w11943 & w11948;
assign w11951 = ~w11949 & ~w11950;
assign w11952 = w11942 & ~w11951;
assign w11953 = ~w11942 & w11951;
assign w11954 = ~w11952 & ~w11953;
assign w11955 = w11931 & w11954;
assign w11956 = ~w11931 & ~w11954;
assign w11957 = ~w11955 & ~w11956;
assign w11958 = w11926 & w11957;
assign w11959 = ~w11926 & ~w11957;
assign w11960 = ~w11958 & ~w11959;
assign w11961 = ~w11146 & ~w11150;
assign w11962 = w11960 & ~w11961;
assign w11963 = ~w11960 & w11961;
assign w11964 = ~w11962 & ~w11963;
assign w11965 = ~w11153 & ~w11158;
assign w11966 = w11964 & ~w11965;
assign w11967 = ~w11964 & w11965;
assign w11968 = ~w11966 & ~w11967;
assign w11969 = w11925 & w11968;
assign w11970 = ~w11925 & ~w11968;
assign w11971 = ~w11969 & ~w11970;
assign w11972 = w11924 & w11971;
assign w11973 = ~w11924 & ~w11971;
assign w11974 = ~w11972 & ~w11973;
assign w11975 = w11923 & ~w11974;
assign w11976 = ~w11923 & w11974;
assign w11977 = ~w11975 & ~w11976;
assign w11978 = w11922 & ~w11977;
assign w11979 = ~w11922 & w11977;
assign w11980 = ~w11978 & ~w11979;
assign w11981 = ~w11170 & ~w11172;
assign w11982 = w11980 & ~w11981;
assign w11983 = ~w11980 & w11981;
assign w11984 = ~w11982 & ~w11983;
assign w11985 = pi136 & pi278;
assign w11986 = ~w11984 & ~w11985;
assign w11987 = w11984 & w11985;
assign w11988 = ~w11986 & ~w11987;
assign w11989 = ~w11178 & ~w11181;
assign w11990 = w11988 & ~w11989;
assign w11991 = ~w11988 & w11989;
assign w11992 = ~w11990 & ~w11991;
assign w11993 = w11921 & ~w11992;
assign w11994 = ~w11921 & w11992;
assign w11995 = ~w11993 & ~w11994;
assign w11996 = w11916 & w11995;
assign w11997 = ~w11916 & ~w11995;
assign w11998 = ~w11996 & ~w11997;
assign w11999 = (~w11192 & ~w11194) | (~w11192 & w16288) | (~w11194 & w16288);
assign w12000 = ~w11998 & w11999;
assign w12001 = w11998 & ~w11999;
assign w12002 = ~w12000 & ~w12001;
assign w12003 = ~w11915 & w12002;
assign w12004 = w11915 & ~w12002;
assign w12005 = ~w12003 & ~w12004;
assign w12006 = w11914 & w12005;
assign w12007 = ~w11914 & ~w12005;
assign w12008 = ~w12006 & ~w12007;
assign w12009 = pi140 & pi274;
assign w12010 = (~w11208 & ~w11204) | (~w11208 & w15984) | (~w11204 & w15984);
assign w12011 = ~w11205 & ~w12010;
assign w12012 = ~w12009 & ~w12011;
assign w12013 = w12009 & w12011;
assign w12014 = ~w12012 & ~w12013;
assign w12015 = ~w12008 & w12014;
assign w12016 = w12008 & ~w12014;
assign w12017 = ~w12015 & ~w12016;
assign w12018 = w11913 & ~w12017;
assign w12019 = ~w11913 & w12017;
assign w12020 = ~w12018 & ~w12019;
assign w12021 = (w11216 & ~w11211) | (w11216 & w16497) | (~w11211 & w16497);
assign w12022 = ~w11213 & ~w12021;
assign w12023 = w12020 & ~w12022;
assign w12024 = ~w12020 & w12022;
assign w12025 = ~w12023 & ~w12024;
assign w12026 = w11215 & w11222;
assign w12027 = ~w11223 & ~w12026;
assign w12028 = w12025 & ~w12027;
assign w12029 = ~w12025 & w12027;
assign w12030 = ~w12028 & ~w12029;
assign w12031 = w11912 & w12030;
assign w12032 = ~w11912 & ~w12030;
assign w12033 = ~w12031 & ~w12032;
assign w12034 = w11911 & w12033;
assign w12035 = ~w11911 & ~w12033;
assign w12036 = ~w12034 & ~w12035;
assign w12037 = ~w11905 & ~w12036;
assign w12038 = w11905 & w12036;
assign w12039 = ~w12037 & ~w12038;
assign w12040 = (~w11234 & ~w11235) | (~w11234 & w16289) | (~w11235 & w16289);
assign w12041 = w12039 & ~w12040;
assign w12042 = ~w12039 & w12040;
assign w12043 = ~w12041 & ~w12042;
assign w12044 = (~w11088 & ~w11238) | (~w11088 & w16290) | (~w11238 & w16290);
assign w12045 = ~w12043 & w12044;
assign w12046 = w12043 & ~w12044;
assign w12047 = ~w12045 & ~w12046;
assign w12048 = w11904 & w12047;
assign w12049 = ~w11904 & ~w12047;
assign w12050 = ~w12048 & ~w12049;
assign w12051 = w11903 & w12050;
assign w12052 = ~w11903 & ~w12050;
assign w12053 = ~w12051 & ~w12052;
assign w12054 = ~w11898 & ~w12053;
assign w12055 = w11898 & w12053;
assign w12056 = ~w12054 & ~w12055;
assign w12057 = (~w11249 & ~w11251) | (~w11249 & w16291) | (~w11251 & w16291);
assign w12058 = w12056 & w12057;
assign w12059 = ~w12056 & ~w12057;
assign w12060 = ~w12058 & ~w12059;
assign w12061 = (~w11079 & ~w11081) | (~w11079 & w17615) | (~w11081 & w17615);
assign w12062 = ~w12060 & w12061;
assign w12063 = w12060 & ~w12061;
assign w12064 = ~w12062 & ~w12063;
assign w12065 = pi148 & pi266;
assign w12066 = pi149 & pi265;
assign w12067 = ~w12065 & w12066;
assign w12068 = w12065 & ~w12066;
assign w12069 = ~w12067 & ~w12068;
assign w12070 = w12064 & w12069;
assign w12071 = ~w12064 & ~w12069;
assign w12072 = ~w12070 & ~w12071;
assign w12073 = ~w11897 & ~w12072;
assign w12074 = w11897 & w12072;
assign w12075 = ~w12073 & ~w12074;
assign w12076 = w11896 & ~w12075;
assign w12077 = ~w11896 & w12075;
assign w12078 = ~w12076 & ~w12077;
assign w12079 = w11264 & w11265;
assign w12080 = ~w11264 & ~w11265;
assign w12081 = ~w11267 & ~w12080;
assign w12082 = ~w12079 & ~w12081;
assign w12083 = w12078 & w12082;
assign w12084 = ~w12078 & ~w12082;
assign w12085 = ~w12083 & ~w12084;
assign w12086 = ~w11266 & ~w11276;
assign w12087 = ~w11277 & ~w12086;
assign w12088 = ~w12085 & ~w12087;
assign w12089 = w12085 & w12087;
assign w12090 = ~w12088 & ~w12089;
assign w12091 = pi151 & pi263;
assign w12092 = ~w12090 & w12091;
assign w12093 = w12090 & ~w12091;
assign w12094 = ~w12092 & ~w12093;
assign w12095 = ~w11895 & w12094;
assign w12096 = w11895 & ~w12094;
assign w12097 = ~w12095 & ~w12096;
assign w12098 = w11890 & w12097;
assign w12099 = ~w11890 & ~w12097;
assign w12100 = ~w12098 & ~w12099;
assign w12101 = ~w11293 & ~w11296;
assign w12102 = w11293 & w11296;
assign w12103 = ~w12101 & ~w12102;
assign w12104 = (w11294 & w12103) | (w11294 & w15985) | (w12103 & w15985);
assign w12105 = w11295 & w12103;
assign w12106 = ~w12104 & ~w12105;
assign w12107 = w12100 & ~w12106;
assign w12108 = ~w12100 & w12106;
assign w12109 = ~w12107 & ~w12108;
assign w12110 = pi155 & pi259;
assign w12111 = (~w12110 & ~w11309) | (~w12110 & w15986) | (~w11309 & w15986);
assign w12112 = w11309 & w15987;
assign w12113 = ~w12111 & ~w12112;
assign w12114 = pi154 & pi260;
assign w12115 = pi156 & pi258;
assign w12116 = ~w12114 & w12115;
assign w12117 = w12114 & ~w12115;
assign w12118 = ~w12116 & ~w12117;
assign w12119 = w12113 & ~w12118;
assign w12120 = ~w12113 & w12118;
assign w12121 = ~w12119 & ~w12120;
assign w12122 = w12109 & w12121;
assign w12123 = ~w12109 & ~w12121;
assign w12124 = ~w12122 & ~w12123;
assign w12125 = w11884 & w12124;
assign w12126 = ~w11884 & ~w12124;
assign w12127 = ~w12125 & ~w12126;
assign w12128 = ~w11309 & ~w12127;
assign w12129 = w11309 & w12127;
assign w12130 = ~w12128 & ~w12129;
assign w12131 = (~w11880 & ~w12130) | (~w11880 & w15988) | (~w12130 & w15988);
assign w12132 = w12130 & w15989;
assign w12133 = ~w12131 & ~w12132;
assign w12134 = pi324 & ~w11070;
assign w12135 = w11328 & w11336;
assign w12136 = (~w11336 & w11326) | (~w11336 & w16292) | (w11326 & w16292);
assign w12137 = (w11326 & w16293) | (w11326 & w16294) | (w16293 & w16294);
assign w12138 = ~w12136 & w12137;
assign w12139 = ~w11332 & ~w12138;
assign w12140 = ~w12134 & w12139;
assign w12141 = w12134 & ~w12139;
assign w12142 = ~w12140 & ~w12141;
assign w12143 = pi325 & ~w9784;
assign w12144 = ~w11316 & ~w12135;
assign w12145 = ~w12143 & w12144;
assign w12146 = w12143 & ~w12144;
assign w12147 = ~w12145 & ~w12146;
assign w12148 = w12142 & ~w12147;
assign w12149 = ~w12142 & w12147;
assign w12150 = ~w12148 & ~w12149;
assign w12151 = w12133 & w12150;
assign w12152 = ~w12133 & ~w12150;
assign w12153 = ~w12151 & ~w12152;
assign w12154 = w11874 & w12153;
assign w12155 = ~w11874 & ~w12153;
assign w12156 = ~w12154 & ~w12155;
assign w12157 = pi327 & ~w8367;
assign w12158 = (w15991 & ~w11356) | (w15991 & w16295) | (~w11356 & w16295);
assign w12159 = (w11356 & w16296) | (w11356 & w16297) | (w16296 & w16297);
assign w12160 = ~w12158 & ~w12159;
assign w12161 = pi326 & w8814;
assign w12162 = ~w11352 & ~w11354;
assign w12163 = w12161 & ~w12162;
assign w12164 = ~w12161 & w12162;
assign w12165 = ~w12163 & ~w12164;
assign w12166 = w12160 & ~w12165;
assign w12167 = ~w12160 & w12165;
assign w12168 = ~w12166 & ~w12167;
assign w12169 = w12156 & w12168;
assign w12170 = ~w12156 & ~w12168;
assign w12171 = ~w12169 & ~w12170;
assign w12172 = ~w11872 & w12171;
assign w12173 = w11872 & ~w12171;
assign w12174 = ~w12172 & ~w12173;
assign w12175 = ~w11870 & w12174;
assign w12176 = w11870 & ~w12174;
assign w12177 = ~w12175 & ~w12176;
assign w12178 = pi329 & ~w7108;
assign w12179 = ~w11366 & ~w11373;
assign w12180 = ~w11365 & ~w12179;
assign w12181 = ~w12178 & ~w12180;
assign w12182 = w12178 & w12180;
assign w12183 = ~w12181 & ~w12182;
assign w12184 = w12177 & ~w12183;
assign w12185 = ~w12177 & w12183;
assign w12186 = ~w12184 & ~w12185;
assign w12187 = pi331 & w5714;
assign w12188 = pi330 & w6283;
assign w12189 = w11043 & ~w11049;
assign w12190 = ~w11374 & ~w12189;
assign w12191 = w12188 & ~w12190;
assign w12192 = ~w12188 & w12190;
assign w12193 = ~w12191 & ~w12192;
assign w12194 = w12187 & ~w12193;
assign w12195 = ~w12187 & w12193;
assign w12196 = ~w12194 & ~w12195;
assign w12197 = w12186 & ~w12196;
assign w12198 = ~w12186 & w12196;
assign w12199 = ~w12197 & ~w12198;
assign w12200 = w11869 & w12199;
assign w12201 = ~w11869 & ~w12199;
assign w12202 = ~w12200 & ~w12201;
assign w12203 = w11856 & w12202;
assign w12204 = ~w11856 & ~w12202;
assign w12205 = ~w12203 & ~w12204;
assign w12206 = (~w4708 & w11025) | (~w4708 & w12209) | (w11025 & w12209);
assign w12207 = ~w11402 & w12206;
assign w12208 = ~w11025 & w15993;
assign w12209 = ~w3979 & ~w4708;
assign w12210 = w11025 & w12209;
assign w12211 = ~w12208 & ~w12210;
assign w12212 = (pi334 & w12207) | (pi334 & w15994) | (w12207 & w15994);
assign w12213 = pi334 & ~w4708;
assign w12214 = ~w11026 & w11402;
assign w12215 = ~w12213 & w12214;
assign w12216 = ~w12212 & ~w12215;
assign w12217 = ~w11040 & ~w11400;
assign w12218 = ~w12216 & w12217;
assign w12219 = w12216 & ~w12217;
assign w12220 = ~w12218 & ~w12219;
assign w12221 = w12205 & w12220;
assign w12222 = ~w12205 & ~w12220;
assign w12223 = ~w12221 & ~w12222;
assign w12224 = w11855 & ~w12223;
assign w12225 = ~w11855 & w12223;
assign w12226 = ~w12224 & ~w12225;
assign w12227 = (~w11009 & ~w11417) | (~w11009 & w16298) | (~w11417 & w16298);
assign w12228 = ~w12226 & w12227;
assign w12229 = w12226 & ~w12227;
assign w12230 = ~w12228 & ~w12229;
assign w12231 = w11850 & w12230;
assign w12232 = ~w11850 & ~w12230;
assign w12233 = ~w12231 & ~w12232;
assign w12234 = w11820 & ~w12233;
assign w12235 = ~w11820 & w12233;
assign w12236 = ~w12234 & ~w12235;
assign w12237 = w11819 & ~w12236;
assign w12238 = ~w11819 & w12236;
assign w12239 = ~w12237 & ~w12238;
assign w12240 = w11814 & w12239;
assign w12241 = ~w11814 & ~w12239;
assign w12242 = ~w12240 & ~w12241;
assign w12243 = w11793 & w12242;
assign w12244 = ~w11793 & ~w12242;
assign w12245 = ~w12243 & ~w12244;
assign w12246 = pi344 & w1101;
assign w12247 = (w15995 & ~w11457) | (w15995 & w16617) | (~w11457 & w16617);
assign w12248 = (w11457 & w16618) | (w11457 & w16619) | (w16618 & w16619);
assign w12249 = ~w12247 & ~w12248;
assign w12250 = ~w10990 & ~w11455;
assign w12251 = pi343 & w1339;
assign w12252 = w12250 & ~w12251;
assign w12253 = ~w12250 & w12251;
assign w12254 = ~w12252 & ~w12253;
assign w12255 = w12249 & ~w12254;
assign w12256 = ~w12249 & w12254;
assign w12257 = ~w12255 & ~w12256;
assign w12258 = w12245 & w12257;
assign w12259 = ~w12245 & ~w12257;
assign w12260 = ~w12258 & ~w12259;
assign w12261 = ~w11784 & w12260;
assign w12262 = w11784 & ~w12260;
assign w12263 = ~w12261 & ~w12262;
assign w12264 = w11783 & w12263;
assign w12265 = ~w11783 & ~w12263;
assign w12266 = ~w12264 & ~w12265;
assign w12267 = (~w10974 & ~w11470) | (~w10974 & w16299) | (~w11470 & w16299);
assign w12268 = ~w11462 & ~w11465;
assign w12269 = (w12268 & w11471) | (w12268 & w15997) | (w11471 & w15997);
assign w12270 = ~w11471 & w15998;
assign w12271 = ~w12269 & ~w12270;
assign w12272 = w12266 & w12271;
assign w12273 = ~w12266 & ~w12271;
assign w12274 = ~w12272 & ~w12273;
assign w12275 = w11764 & ~w12274;
assign w12276 = ~w11764 & w12274;
assign w12277 = ~w12275 & ~w12276;
assign w12278 = pi349 & w466;
assign w12279 = (~w12278 & ~w11476) | (~w12278 & w16300) | (~w11476 & w16300);
assign w12280 = w11476 & w16301;
assign w12281 = ~w12279 & ~w12280;
assign w12282 = w12277 & w12281;
assign w12283 = ~w12277 & ~w12281;
assign w12284 = ~w12282 & ~w12283;
assign w12285 = w11759 & w12284;
assign w12286 = ~w11759 & ~w12284;
assign w12287 = ~w12285 & ~w12286;
assign w12288 = pi286 & ~w12287;
assign w12289 = ~pi286 & w12287;
assign w12290 = ~w12288 & ~w12289;
assign w12291 = ~w10965 & ~w11480;
assign w12292 = w12290 & w12291;
assign w12293 = ~w12290 & ~w12291;
assign w12294 = ~w12292 & ~w12293;
assign w12295 = ~w11758 & ~w12294;
assign w12296 = w11758 & w12294;
assign w12297 = ~w135 & ~w12295;
assign w12298 = ~w12296 & w12297;
assign w12299 = pi161 & ~w207;
assign w12300 = ~w12298 & w12299;
assign w12301 = ~pi160 & ~w11495;
assign w12302 = ~w12300 & w12301;
assign w12303 = ~pi093 & ~pi161;
assign w12304 = pi128 & pi292;
assign w12305 = w11497 & ~w11752;
assign w12306 = pi129 & ~pi293;
assign w12307 = ~w12305 & ~w12306;
assign w12308 = pi294 & ~w653;
assign w12309 = (~w11500 & w11749) | (~w11500 & w15999) | (w11749 & w15999);
assign w12310 = w12308 & ~w12309;
assign w12311 = ~w12308 & w12309;
assign w12312 = ~w12310 & ~w12311;
assign w12313 = pi296 & w698;
assign w12314 = w855 & w11728;
assign w12315 = pi299 & w1220;
assign w12316 = (w11510 & ~w11719) | (w11510 & w16000) | (~w11719 & w16000);
assign w12317 = ~w11721 & ~w12316;
assign w12318 = w12315 & ~w12317;
assign w12319 = ~w12315 & w12317;
assign w12320 = ~w12318 & ~w12319;
assign w12321 = pi300 & w1420;
assign w12322 = w11706 & w11707;
assign w12323 = ~w10915 & ~w10918;
assign w12324 = ~w12322 & w12323;
assign w12325 = ~w11706 & ~w11707;
assign w12326 = ~w12324 & ~w12325;
assign w12327 = ~w12321 & ~w12326;
assign w12328 = w12321 & w12326;
assign w12329 = ~w12327 & ~w12328;
assign w12330 = pi301 & w1693;
assign w12331 = pi303 & ~w2473;
assign w12332 = pi305 & w2925;
assign w12333 = pi307 & w3710;
assign w12334 = pi309 & w4539;
assign w12335 = pi311 & w5862;
assign w12336 = ~w11635 & ~w11637;
assign w12337 = ~w11626 & ~w11630;
assign w12338 = pi312 & w6437;
assign w12339 = w12337 & w12338;
assign w12340 = ~w12337 & ~w12338;
assign w12341 = ~w12339 & ~w12340;
assign w12342 = pi314 & w7268;
assign w12343 = pi315 & w7909;
assign w12344 = ~w11607 & ~w11609;
assign w12345 = ~w12343 & w12344;
assign w12346 = w12343 & ~w12344;
assign w12347 = ~w12345 & ~w12346;
assign w12348 = pi316 & w9022;
assign w12349 = pi317 & w9270;
assign w12350 = pi318 & w9992;
assign w12351 = pi319 & w10753;
assign w12352 = pi156 & ~pi157;
assign w12353 = ~pi156 & pi157;
assign w12354 = ~w12352 & ~w12353;
assign w12355 = ~w11540 & ~w11557;
assign w12356 = ~w11541 & ~w12355;
assign w12357 = w12354 & w12356;
assign w12358 = ~w12354 & ~w12356;
assign w12359 = ~w12357 & ~w12358;
assign w12360 = pi321 & w12359;
assign w12361 = w11558 & ~w11560;
assign w12362 = ~w10753 & w11557;
assign w12363 = ~w11563 & ~w12362;
assign w12364 = pi320 & w12359;
assign w12365 = ~w12361 & w12364;
assign w12366 = ~w12363 & w12365;
assign w12367 = w12360 & ~w12366;
assign w12368 = w11563 & ~w12360;
assign w12369 = ~w11557 & ~w12368;
assign w12370 = ~w10753 & ~w12359;
assign w12371 = ~w11562 & w12370;
assign w12372 = w11558 & ~w12371;
assign w12373 = pi320 & ~w12372;
assign w12374 = ~w12369 & w12373;
assign w12375 = ~w12367 & ~w12374;
assign w12376 = w12351 & ~w12375;
assign w12377 = ~w12351 & w12375;
assign w12378 = ~w12376 & ~w12377;
assign w12379 = ~w11569 & ~w11575;
assign w12380 = ~w12378 & ~w12379;
assign w12381 = w12378 & w12379;
assign w12382 = ~w12380 & ~w12381;
assign w12383 = w12350 & w12382;
assign w12384 = ~w12350 & ~w12382;
assign w12385 = ~w12383 & ~w12384;
assign w12386 = w11583 & ~w11590;
assign w12387 = w12385 & ~w12386;
assign w12388 = ~w12385 & w12386;
assign w12389 = ~w12387 & ~w12388;
assign w12390 = w12349 & ~w12389;
assign w12391 = ~w12349 & w12389;
assign w12392 = ~w12390 & ~w12391;
assign w12393 = ~w11592 & ~w11596;
assign w12394 = w12392 & w12393;
assign w12395 = ~w12392 & ~w12393;
assign w12396 = ~w12394 & ~w12395;
assign w12397 = ~w11599 & ~w11604;
assign w12398 = w12396 & ~w12397;
assign w12399 = ~w12396 & w12397;
assign w12400 = ~w12398 & ~w12399;
assign w12401 = w12348 & w12400;
assign w12402 = ~w12348 & ~w12400;
assign w12403 = ~w12401 & ~w12402;
assign w12404 = w12347 & w12403;
assign w12405 = ~w12347 & ~w12403;
assign w12406 = ~w12404 & ~w12405;
assign w12407 = w12342 & w12406;
assign w12408 = ~w12342 & ~w12406;
assign w12409 = ~w12407 & ~w12408;
assign w12410 = ~w11612 & ~w11616;
assign w12411 = w12409 & w12410;
assign w12412 = ~w12409 & ~w12410;
assign w12413 = ~w12411 & ~w12412;
assign w12414 = pi313 & w6652;
assign w12415 = ~w12413 & w12414;
assign w12416 = w12413 & ~w12414;
assign w12417 = ~w12415 & ~w12416;
assign w12418 = ~w11620 & ~w11623;
assign w12419 = w12417 & ~w12418;
assign w12420 = ~w12417 & w12418;
assign w12421 = ~w12419 & ~w12420;
assign w12422 = w12341 & w12421;
assign w12423 = ~w12341 & ~w12421;
assign w12424 = ~w12422 & ~w12423;
assign w12425 = w12336 & ~w12424;
assign w12426 = ~w12336 & w12424;
assign w12427 = ~w12425 & ~w12426;
assign w12428 = w12335 & ~w12427;
assign w12429 = ~w12335 & w12427;
assign w12430 = ~w12428 & ~w12429;
assign w12431 = w5316 & ~w12430;
assign w12432 = w4539 & w12431;
assign w12433 = ~w11641 & w12432;
assign w12434 = pi310 & w5316;
assign w12435 = w12430 & ~w12434;
assign w12436 = ~w12430 & w12434;
assign w12437 = ~w12435 & ~w12436;
assign w12438 = w11642 & ~w12437;
assign w12439 = ~w5316 & w11529;
assign w12440 = w12430 & w12439;
assign w12441 = ~w12433 & ~w12440;
assign w12442 = ~w12438 & w12441;
assign w12443 = ~w11643 & ~w12442;
assign w12444 = w11641 & w12432;
assign w12445 = ~w11641 & ~w12431;
assign w12446 = ~w12435 & w12445;
assign w12447 = ~w12444 & ~w12446;
assign w12448 = ~w11639 & ~w12447;
assign w12449 = ~w11529 & ~w11642;
assign w12450 = w12437 & w12449;
assign w12451 = ~w12448 & ~w12450;
assign w12452 = ~w12443 & w12451;
assign w12453 = w12334 & ~w12452;
assign w12454 = ~w12334 & w12452;
assign w12455 = ~w12453 & ~w12454;
assign w12456 = ~w11655 & ~w11658;
assign w12457 = pi308 & w4382;
assign w12458 = ~w11649 & ~w11652;
assign w12459 = ~w12457 & ~w12458;
assign w12460 = ~w4382 & ~w11648;
assign w12461 = ~w11527 & ~w12460;
assign w12462 = pi308 & ~w11649;
assign w12463 = ~w12461 & w12462;
assign w12464 = ~w12459 & ~w12463;
assign w12465 = w12456 & ~w12464;
assign w12466 = ~w12456 & w12464;
assign w12467 = ~w12465 & ~w12466;
assign w12468 = w12455 & w12467;
assign w12469 = ~w12455 & ~w12467;
assign w12470 = ~w12468 & ~w12469;
assign w12471 = w12333 & w12470;
assign w12472 = ~w12333 & ~w12470;
assign w12473 = ~w12471 & ~w12472;
assign w12474 = ~w11662 & ~w11665;
assign w12475 = ~w12473 & w12474;
assign w12476 = w12473 & ~w12474;
assign w12477 = ~w12475 & ~w12476;
assign w12478 = pi306 & w3304;
assign w12479 = ~w12477 & ~w12478;
assign w12480 = w12477 & w12478;
assign w12481 = ~w12479 & ~w12480;
assign w12482 = ~w11669 & w12481;
assign w12483 = w9346 & ~w12477;
assign w12484 = w11669 & w12483;
assign w12485 = ~w3304 & w11524;
assign w12486 = w12477 & w12485;
assign w12487 = ~w12484 & ~w12486;
assign w12488 = ~w12482 & w12487;
assign w12489 = w11667 & ~w12488;
assign w12490 = ~w11667 & w12483;
assign w12491 = ~w12486 & ~w12490;
assign w12492 = ~w11669 & ~w12491;
assign w12493 = ~w11671 & ~w12481;
assign w12494 = ~w11673 & w12493;
assign w12495 = ~w12492 & ~w12494;
assign w12496 = ~w12489 & w12495;
assign w12497 = ~w12332 & ~w12496;
assign w12498 = w12332 & w12496;
assign w12499 = ~w12497 & ~w12498;
assign w12500 = ~w11677 & ~w11680;
assign w12501 = w12499 & w12500;
assign w12502 = ~w12499 & ~w12500;
assign w12503 = ~w12501 & ~w12502;
assign w12504 = pi304 & w2801;
assign w12505 = ~w11684 & w11686;
assign w12506 = ~w11683 & ~w12505;
assign w12507 = ~w12504 & ~w12506;
assign w12508 = w12504 & w12506;
assign w12509 = ~w12507 & ~w12508;
assign w12510 = w12503 & ~w12509;
assign w12511 = ~w12503 & w12509;
assign w12512 = ~w12510 & ~w12511;
assign w12513 = w12331 & w12512;
assign w12514 = ~w12331 & ~w12512;
assign w12515 = ~w12513 & ~w12514;
assign w12516 = ~w11519 & ~w11691;
assign w12517 = w12515 & ~w12516;
assign w12518 = ~w12515 & w12516;
assign w12519 = ~w12517 & ~w12518;
assign w12520 = ~w11695 & w12519;
assign w12521 = w11695 & ~w12519;
assign w12522 = ~w12520 & ~w12521;
assign w12523 = ~w1954 & ~w11698;
assign w12524 = ~w12522 & w12523;
assign w12525 = pi302 & w1954;
assign w12526 = ~w12519 & w12525;
assign w12527 = w12519 & ~w12525;
assign w12528 = ~w11512 & ~w11694;
assign w12529 = ~w12526 & w12528;
assign w12530 = ~w12527 & w12529;
assign w12531 = ~w11694 & ~w12519;
assign w12532 = w1693 & ~w11695;
assign w12533 = w12531 & ~w12532;
assign w12534 = pi302 & ~w12520;
assign w12535 = ~w12531 & ~w12534;
assign w12536 = w1954 & ~w12533;
assign w12537 = ~w12535 & w12536;
assign w12538 = ~w12524 & ~w12530;
assign w12539 = ~w12537 & w12538;
assign w12540 = ~w12330 & ~w12539;
assign w12541 = w12330 & w12539;
assign w12542 = ~w12540 & ~w12541;
assign w12543 = ~w11700 & ~w11705;
assign w12544 = w12542 & w12543;
assign w12545 = ~w12542 & ~w12543;
assign w12546 = ~w12544 & ~w12545;
assign w12547 = w12329 & ~w12546;
assign w12548 = ~w12329 & w12546;
assign w12549 = ~w12547 & ~w12548;
assign w12550 = ~w12320 & w12549;
assign w12551 = w12320 & ~w12549;
assign w12552 = ~w12550 & ~w12551;
assign w12553 = (pi298 & w12552) | (pi298 & w16498) | (w12552 & w16498);
assign w12554 = ~w12314 & ~w12553;
assign w12555 = pi298 & w11727;
assign w12556 = w12552 & ~w12555;
assign w12557 = w1159 & ~w12556;
assign w12558 = ~w12554 & w12557;
assign w12559 = ~w11726 & ~w11729;
assign w12560 = ~w11727 & ~w12559;
assign w12561 = ~w11727 & ~w12552;
assign w12562 = (~w1159 & w12560) | (~w1159 & w16001) | (w12560 & w16001);
assign w12563 = ~w12561 & w12562;
assign w12564 = pi298 & w1159;
assign w12565 = ~w12552 & w12564;
assign w12566 = w12552 & ~w12564;
assign w12567 = w12559 & ~w12565;
assign w12568 = ~w12566 & w12567;
assign w12569 = ~w12563 & ~w12568;
assign w12570 = ~w12558 & w12569;
assign w12571 = (w855 & w11733) | (w855 & w15823) | (w11733 & w15823);
assign w12572 = w698 & ~w855;
assign w12573 = ~w12570 & ~w12572;
assign w12574 = pi297 & ~w11734;
assign w12575 = (w12574 & ~w12570) | (w12574 & w12580) | (~w12570 & w12580);
assign w12576 = ~w12573 & w12575;
assign w12577 = pi297 & w855;
assign w12578 = ~w11733 & ~w12577;
assign w12579 = ~w12570 & ~w12578;
assign w12580 = w12571 & w12574;
assign w12581 = w12579 & ~w12580;
assign w12582 = ~w11736 & w12578;
assign w12583 = w12570 & w12582;
assign w12584 = ~w12581 & ~w12583;
assign w12585 = ~w12576 & w12584;
assign w12586 = (~w11741 & ~w11743) | (~w11741 & w16002) | (~w11743 & w16002);
assign w12587 = ~w12585 & w12586;
assign w12588 = w12585 & ~w12586;
assign w12589 = ~w12587 & ~w12588;
assign w12590 = w12313 & ~w12589;
assign w12591 = ~w12313 & w12589;
assign w12592 = ~w12590 & ~w12591;
assign w12593 = pi295 & w709;
assign w12594 = ~w11504 & ~w11748;
assign w12595 = (w12593 & w11748) | (w12593 & w16003) | (w11748 & w16003);
assign w12596 = ~w11748 & w16004;
assign w12597 = ~w12595 & ~w12596;
assign w12598 = w12592 & w12597;
assign w12599 = ~w12592 & ~w12597;
assign w12600 = ~w12598 & ~w12599;
assign w12601 = w12312 & w12600;
assign w12602 = ~w12312 & ~w12600;
assign w12603 = ~w12601 & ~w12602;
assign w12604 = pi129 & ~w12603;
assign w12605 = ~pi129 & w12603;
assign w12606 = ~w12604 & ~w12605;
assign w12607 = w12307 & w12606;
assign w12608 = ~w12307 & ~w12606;
assign w12609 = ~w12607 & ~w12608;
assign w12610 = w12304 & w12609;
assign w12611 = ~w12304 & ~w12609;
assign w12612 = ~w12610 & ~w12611;
assign w12613 = pi351 & w456;
assign w12614 = pi349 & ~w537;
assign w12615 = (~w12280 & ~w12277) | (~w12280 & w16005) | (~w12277 & w16005);
assign w12616 = ~w12614 & w12615;
assign w12617 = w12614 & ~w12615;
assign w12618 = ~w12616 & ~w12617;
assign w12619 = pi348 & ~w615;
assign w12620 = (w12619 & w12275) | (w12619 & w16006) | (w12275 & w16006);
assign w12621 = ~w12275 & w16007;
assign w12622 = ~w12620 & ~w12621;
assign w12623 = pi346 & ~w955;
assign w12624 = ~w12260 & ~w12268;
assign w12625 = (~w11765 & w12260) | (~w11765 & w16302) | (w12260 & w16302);
assign w12626 = w12260 & w12268;
assign w12627 = (~w10981 & ~w11467) | (~w10981 & w16008) | (~w11467 & w16008);
assign w12628 = ~w11768 & w12627;
assign w12629 = ~w12626 & ~w12628;
assign w12630 = w12625 & w12629;
assign w12631 = w12629 & w16303;
assign w12632 = w11768 & ~w12627;
assign w12633 = ~w12623 & ~w12632;
assign w12634 = ~w955 & ~w12628;
assign w12635 = ~w12633 & ~w12634;
assign w12636 = ~w12624 & ~w12626;
assign w12637 = ~pi345 & w12636;
assign w12638 = pi345 & ~w12636;
assign w12639 = w12623 & ~w12632;
assign w12640 = ~w12637 & w12639;
assign w12641 = ~w12638 & w12640;
assign w12642 = ~w12631 & ~w12635;
assign w12643 = ~w12641 & w12642;
assign w12644 = ~w12625 & ~w12626;
assign w12645 = pi341 & ~w2170;
assign w12646 = pi339 & w2698;
assign w12647 = ~w11810 & w16009;
assign w12648 = (w11820 & w11810) | (w11820 & w16010) | (w11810 & w16010);
assign w12649 = ~w12647 & ~w12648;
assign w12650 = w12233 & w12649;
assign w12651 = ~w12647 & ~w12650;
assign w12652 = w12646 & w12651;
assign w12653 = ~w12646 & ~w12651;
assign w12654 = ~w12652 & ~w12653;
assign w12655 = pi338 & ~w3183;
assign w12656 = ~w11807 & ~w11822;
assign w12657 = ~w11824 & w12656;
assign w12658 = w11824 & ~w12656;
assign w12659 = w11847 & w12230;
assign w12660 = ~w11847 & ~w12230;
assign w12661 = ~w12658 & ~w12659;
assign w12662 = ~w12660 & w12661;
assign w12663 = ~w12657 & ~w12662;
assign w12664 = ~w12655 & w12663;
assign w12665 = w12655 & ~w12663;
assign w12666 = ~w12664 & ~w12665;
assign w12667 = w12654 & ~w12666;
assign w12668 = ~w12654 & w12666;
assign w12669 = ~w12667 & ~w12668;
assign w12670 = pi340 & ~w2373;
assign w12671 = ~w11794 & w11801;
assign w12672 = w12233 & w16011;
assign w12673 = ~w12649 & ~w12671;
assign w12674 = w11795 & ~w11799;
assign w12675 = (~w12674 & w12233) | (~w12674 & w16012) | (w12233 & w16012);
assign w12676 = ~w12672 & w12675;
assign w12677 = ~w12670 & w12676;
assign w12678 = w12670 & ~w12676;
assign w12679 = ~w12677 & ~w12678;
assign w12680 = pi335 & ~w4708;
assign w12681 = ~w11854 & ~w12224;
assign w12682 = pi331 & w6283;
assign w12683 = ~w12186 & ~w12193;
assign w12684 = w12186 & w12193;
assign w12685 = ~w12683 & ~w12684;
assign w12686 = w12187 & w12685;
assign w12687 = w11866 & ~w12686;
assign w12688 = ~w12187 & ~w12685;
assign w12689 = ~w12687 & ~w12688;
assign w12690 = ~w12682 & ~w12689;
assign w12691 = w12682 & w12689;
assign w12692 = ~w12690 & ~w12691;
assign w12693 = ~w12182 & ~w12185;
assign w12694 = pi327 & w8814;
assign w12695 = ~w12133 & ~w12144;
assign w12696 = (w12144 & ~w12130) | (w12144 & w16304) | (~w12130 & w16304);
assign w12697 = ~w12131 & w12696;
assign w12698 = ~w12141 & ~w12695;
assign w12699 = ~w12697 & w12698;
assign w12700 = ~w12140 & ~w12699;
assign w12701 = w11309 & ~w11881;
assign w12702 = w12124 & ~w12701;
assign w12703 = ~w12124 & ~w12128;
assign w12704 = ~w12702 & ~w12703;
assign w12705 = pi157 & pi258;
assign w12706 = pi155 & pi260;
assign w12707 = ~w12108 & w12114;
assign w12708 = ~w12107 & w12707;
assign w12709 = (~w12111 & w12109) | (~w12111 & w16013) | (w12109 & w16013);
assign w12710 = ~w12708 & w12709;
assign w12711 = ~w12710 & w16499;
assign w12712 = (w12706 & w12710) | (w12706 & w16500) | (w12710 & w16500);
assign w12713 = ~w12711 & ~w12712;
assign w12714 = pi154 & pi261;
assign w12715 = pi151 & pi264;
assign w12716 = (~w12091 & ~w12085) | (~w12091 & w16501) | (~w12085 & w16501);
assign w12717 = ~w12088 & ~w12716;
assign w12718 = w12715 & w12717;
assign w12719 = ~w12715 & ~w12717;
assign w12720 = ~w12718 & ~w12719;
assign w12721 = pi150 & pi265;
assign w12722 = pi148 & pi267;
assign w12723 = pi147 & pi268;
assign w12724 = pi146 & pi269;
assign w12725 = pi145 & pi270;
assign w12726 = pi144 & pi271;
assign w12727 = ~w12041 & w16014;
assign w12728 = (w12726 & w12041) | (w12726 & w16015) | (w12041 & w16015);
assign w12729 = ~w12727 & ~w12728;
assign w12730 = pi143 & pi272;
assign w12731 = pi142 & pi273;
assign w12732 = pi141 & pi274;
assign w12733 = pi140 & pi275;
assign w12734 = pi139 & pi276;
assign w12735 = pi138 & pi277;
assign w12736 = pi137 & pi278;
assign w12737 = pi136 & pi279;
assign w12738 = pi135 & pi280;
assign w12739 = ~w11978 & ~w11982;
assign w12740 = pi133 & pi282;
assign w12741 = pi132 & pi283;
assign w12742 = (~w11958 & ~w11960) | (~w11958 & w16016) | (~w11960 & w16016);
assign w12743 = w12741 & ~w12742;
assign w12744 = ~w12741 & w12742;
assign w12745 = ~w12743 & ~w12744;
assign w12746 = pi131 & pi284;
assign w12747 = ~w11930 & ~w11955;
assign w12748 = ~w12746 & w12747;
assign w12749 = w12746 & ~w12747;
assign w12750 = ~w12748 & ~w12749;
assign w12751 = ~w11941 & ~w11952;
assign w12752 = pi129 & pi286;
assign w12753 = pi128 & pi287;
assign w12754 = w12752 & ~w12753;
assign w12755 = ~w12752 & w12753;
assign w12756 = ~w12754 & ~w12755;
assign w12757 = ~w11943 & ~w11946;
assign w12758 = pi130 & pi285;
assign w12759 = w12757 & ~w12758;
assign w12760 = ~pi285 & w11946;
assign w12761 = w646 & ~w11947;
assign w12762 = ~w12760 & w12761;
assign w12763 = ~w12756 & ~w12759;
assign w12764 = ~w12762 & w12763;
assign w12765 = w12758 & ~w12761;
assign w12766 = w12756 & ~w12760;
assign w12767 = ~w12765 & w12766;
assign w12768 = ~w12764 & ~w12767;
assign w12769 = ~w11947 & ~w12757;
assign w12770 = w12756 & ~w12769;
assign w12771 = ~w12756 & w12769;
assign w12772 = ~w12770 & ~w12771;
assign w12773 = ~pi130 & ~w11950;
assign w12774 = w12772 & w12773;
assign w12775 = ~w12768 & ~w12774;
assign w12776 = ~w12751 & w12775;
assign w12777 = w12751 & ~w12775;
assign w12778 = ~w12776 & ~w12777;
assign w12779 = w12750 & ~w12778;
assign w12780 = ~w12750 & w12778;
assign w12781 = ~w12779 & ~w12780;
assign w12782 = w12745 & w12781;
assign w12783 = ~w12745 & ~w12781;
assign w12784 = ~w12782 & ~w12783;
assign w12785 = w12740 & w12784;
assign w12786 = ~w12740 & ~w12784;
assign w12787 = ~w12785 & ~w12786;
assign w12788 = ~w11966 & ~w11969;
assign w12789 = w12787 & ~w12788;
assign w12790 = ~w12787 & w12788;
assign w12791 = ~w12789 & ~w12790;
assign w12792 = ~w11973 & w12791;
assign w12793 = pi134 & pi281;
assign w12794 = ~w11972 & ~w12791;
assign w12795 = pi280 & ~w11973;
assign w12796 = w12794 & ~w12795;
assign w12797 = w12793 & ~w12796;
assign w12798 = ~w12792 & w12797;
assign w12799 = w12794 & w12795;
assign w12800 = pi281 & ~w12799;
assign w12801 = ~w11923 & ~w11972;
assign w12802 = w12792 & ~w12801;
assign w12803 = w11973 & ~w12791;
assign w12804 = ~pi281 & ~w12803;
assign w12805 = ~w12802 & w12804;
assign w12806 = ~w12800 & ~w12805;
assign w12807 = w12791 & ~w12793;
assign w12808 = ~w12791 & w12793;
assign w12809 = w12801 & ~w12807;
assign w12810 = ~w12808 & w12809;
assign w12811 = ~w12798 & ~w12810;
assign w12812 = ~w12806 & w12811;
assign w12813 = w12739 & ~w12812;
assign w12814 = ~w12739 & w12812;
assign w12815 = ~w12813 & ~w12814;
assign w12816 = ~w12738 & w12815;
assign w12817 = w12738 & ~w12815;
assign w12818 = ~w12816 & ~w12817;
assign w12819 = ~w12737 & w12818;
assign w12820 = w12737 & ~w12818;
assign w12821 = ~w12819 & ~w12820;
assign w12822 = ~w11986 & ~w11990;
assign w12823 = ~w12821 & ~w12822;
assign w12824 = w12821 & w12822;
assign w12825 = ~w12823 & ~w12824;
assign w12826 = ~w12736 & ~w12825;
assign w12827 = w12736 & w12825;
assign w12828 = ~w12826 & ~w12827;
assign w12829 = ~w11920 & ~w11993;
assign w12830 = w12828 & ~w12829;
assign w12831 = ~w12828 & w12829;
assign w12832 = ~w12830 & ~w12831;
assign w12833 = ~w11996 & w11999;
assign w12834 = ~w11997 & ~w12833;
assign w12835 = w12832 & w12834;
assign w12836 = ~w12832 & ~w12834;
assign w12837 = ~w12835 & ~w12836;
assign w12838 = w12735 & w12837;
assign w12839 = ~w12735 & ~w12837;
assign w12840 = ~w12838 & ~w12839;
assign w12841 = w12734 & w12840;
assign w12842 = ~w12734 & ~w12840;
assign w12843 = ~w12841 & ~w12842;
assign w12844 = (~w12003 & ~w12005) | (~w12003 & w16017) | (~w12005 & w16017);
assign w12845 = w12843 & ~w12844;
assign w12846 = ~w12843 & w12844;
assign w12847 = ~w12845 & ~w12846;
assign w12848 = w12733 & w12847;
assign w12849 = ~w12733 & ~w12847;
assign w12850 = ~w12848 & ~w12849;
assign w12851 = ~w12012 & ~w12015;
assign w12852 = w12850 & w12851;
assign w12853 = ~w12850 & ~w12851;
assign w12854 = ~w12852 & ~w12853;
assign w12855 = (~w12018 & ~w12020) | (~w12018 & w16018) | (~w12020 & w16018);
assign w12856 = w12854 & ~w12855;
assign w12857 = ~w12854 & w12855;
assign w12858 = ~w12856 & ~w12857;
assign w12859 = w12732 & w12858;
assign w12860 = ~w12732 & ~w12858;
assign w12861 = ~w12859 & ~w12860;
assign w12862 = w12731 & w12861;
assign w12863 = ~w12731 & ~w12861;
assign w12864 = ~w12862 & ~w12863;
assign w12865 = ~w12028 & ~w12031;
assign w12866 = ~w12864 & w12865;
assign w12867 = w12864 & ~w12865;
assign w12868 = ~w12866 & ~w12867;
assign w12869 = w12730 & w12868;
assign w12870 = ~w12730 & ~w12868;
assign w12871 = ~w12869 & ~w12870;
assign w12872 = ~w11909 & ~w12034;
assign w12873 = w12871 & ~w12872;
assign w12874 = ~w12871 & w12872;
assign w12875 = ~w12873 & ~w12874;
assign w12876 = w12729 & w12875;
assign w12877 = ~w12729 & ~w12875;
assign w12878 = ~w12876 & ~w12877;
assign w12879 = ~w12725 & ~w12878;
assign w12880 = w12725 & w12878;
assign w12881 = ~w12879 & ~w12880;
assign w12882 = ~w12046 & ~w12048;
assign w12883 = ~w12881 & w12882;
assign w12884 = w12881 & ~w12882;
assign w12885 = ~w12883 & ~w12884;
assign w12886 = w12724 & w12885;
assign w12887 = ~w12724 & ~w12885;
assign w12888 = ~w12886 & ~w12887;
assign w12889 = ~w11901 & ~w12051;
assign w12890 = w12888 & ~w12889;
assign w12891 = ~w12888 & w12889;
assign w12892 = ~w12890 & ~w12891;
assign w12893 = ~w12055 & ~w12058;
assign w12894 = ~w12892 & w12893;
assign w12895 = w12892 & ~w12893;
assign w12896 = ~w12894 & ~w12895;
assign w12897 = w12723 & w12896;
assign w12898 = ~w12723 & ~w12896;
assign w12899 = ~w12897 & ~w12898;
assign w12900 = ~w12722 & ~w12899;
assign w12901 = w12722 & w12899;
assign w12902 = ~w12900 & ~w12901;
assign w12903 = ~w12063 & ~w12065;
assign w12904 = ~w12062 & ~w12903;
assign w12905 = ~w12902 & w12904;
assign w12906 = w12902 & ~w12904;
assign w12907 = ~w12905 & ~w12906;
assign w12908 = pi149 & pi266;
assign w12909 = ~w12066 & w12072;
assign w12910 = ~w12073 & ~w12909;
assign w12911 = w12908 & w12910;
assign w12912 = ~w12908 & ~w12910;
assign w12913 = ~w12911 & ~w12912;
assign w12914 = w12907 & ~w12913;
assign w12915 = ~w12907 & w12913;
assign w12916 = ~w12914 & ~w12915;
assign w12917 = ~w12076 & ~w12083;
assign w12918 = w12916 & ~w12917;
assign w12919 = ~w12916 & w12917;
assign w12920 = ~w12918 & ~w12919;
assign w12921 = w12721 & w12920;
assign w12922 = ~w12721 & ~w12920;
assign w12923 = ~w12921 & ~w12922;
assign w12924 = w12720 & w12923;
assign w12925 = ~w12720 & ~w12923;
assign w12926 = ~w12924 & ~w12925;
assign w12927 = pi152 & pi263;
assign w12928 = (w12927 & w16019) | (w12927 & w12096) | (w16019 & w12096);
assign w12929 = (w16020 & w12094) | (w16020 & w16502) | (w12094 & w16502);
assign w12930 = ~w12928 & ~w12929;
assign w12931 = ~w12926 & ~w12930;
assign w12932 = w12926 & w12930;
assign w12933 = ~w12931 & ~w12932;
assign w12934 = pi153 & pi262;
assign w12935 = (w12934 & w12098) | (w12934 & w16021) | (w12098 & w16021);
assign w12936 = ~w12098 & w16022;
assign w12937 = ~w12935 & ~w12936;
assign w12938 = ~w12933 & w12937;
assign w12939 = w12933 & ~w12937;
assign w12940 = ~w12938 & ~w12939;
assign w12941 = w12714 & ~w12940;
assign w12942 = ~w12714 & w12940;
assign w12943 = ~w12941 & ~w12942;
assign w12944 = ~w12107 & ~w12707;
assign w12945 = ~w12943 & w12944;
assign w12946 = w12943 & ~w12944;
assign w12947 = ~w12945 & ~w12946;
assign w12948 = w12713 & ~w12947;
assign w12949 = ~w12713 & w12947;
assign w12950 = ~w12948 & ~w12949;
assign w12951 = w12115 & ~w12124;
assign w12952 = pi259 & w12951;
assign w12953 = pi156 & pi259;
assign w12954 = ~w12951 & ~w12953;
assign w12955 = ~w12952 & ~w12954;
assign w12956 = ~w12950 & w12955;
assign w12957 = w12950 & ~w12955;
assign w12958 = ~w12956 & ~w12957;
assign w12959 = ~w12705 & ~w12958;
assign w12960 = w12705 & w12958;
assign w12961 = ~w12959 & ~w12960;
assign w12962 = w12704 & w12961;
assign w12963 = ~w12704 & ~w12961;
assign w12964 = ~w12962 & ~w12963;
assign w12965 = pi322 & w12964;
assign w12966 = pi324 & w11879;
assign w12967 = pi323 & w12130;
assign w12968 = ~w12131 & ~w12696;
assign w12969 = w12967 & w12968;
assign w12970 = ~w12967 & ~w12968;
assign w12971 = ~w12969 & ~w12970;
assign w12972 = ~w12966 & w12971;
assign w12973 = w12966 & ~w12971;
assign w12974 = ~w12972 & ~w12973;
assign w12975 = w12964 & w16023;
assign w12976 = (~w12974 & ~w12964) | (~w12974 & w16024) | (~w12964 & w16024);
assign w12977 = ~w12975 & ~w12976;
assign w12978 = ~w12700 & w12977;
assign w12979 = w12700 & ~w12977;
assign w12980 = ~w12978 & ~w12979;
assign w12981 = w12143 & w12153;
assign w12982 = ~w12155 & ~w12981;
assign w12983 = pi325 & ~w11070;
assign w12984 = w12982 & ~w12983;
assign w12985 = ~w12982 & w12983;
assign w12986 = ~w12984 & ~w12985;
assign w12987 = pi326 & ~w9784;
assign w12988 = ~w12987 & w17703;
assign w12989 = (w12156 & w16503) | (w12156 & w16504) | (w16503 & w16504);
assign w12990 = ~w12988 & ~w12989;
assign w12991 = w12986 & ~w12990;
assign w12992 = ~w12986 & w12990;
assign w12993 = ~w12991 & ~w12992;
assign w12994 = w12980 & w12993;
assign w12995 = ~w12980 & ~w12993;
assign w12996 = ~w12994 & ~w12995;
assign w12997 = ~w12694 & w12996;
assign w12998 = w12694 & ~w12996;
assign w12999 = ~w12997 & ~w12998;
assign w13000 = pi328 & ~w8367;
assign w13001 = w13000 & w17704;
assign w13002 = (w12174 & w16505) | (w12174 & w16506) | (w16505 & w16506);
assign w13003 = ~w13001 & ~w13002;
assign w13004 = pi329 & w7742;
assign w13005 = ~w12159 & ~w12171;
assign w13006 = ~w12158 & ~w13005;
assign w13007 = w13004 & ~w13006;
assign w13008 = ~w13004 & w13006;
assign w13009 = ~w13007 & ~w13008;
assign w13010 = w13003 & ~w13009;
assign w13011 = ~w13003 & w13009;
assign w13012 = ~w13010 & ~w13011;
assign w13013 = w12999 & w13012;
assign w13014 = ~w12999 & ~w13012;
assign w13015 = ~w13013 & ~w13014;
assign w13016 = ~w12693 & ~w13015;
assign w13017 = w12693 & w13015;
assign w13018 = ~w13016 & ~w13017;
assign w13019 = pi330 & ~w7108;
assign w13020 = ~w12191 & ~w12684;
assign w13021 = w13019 & ~w13020;
assign w13022 = ~w13019 & w13020;
assign w13023 = ~w13021 & ~w13022;
assign w13024 = w13018 & ~w13023;
assign w13025 = ~w13018 & w13023;
assign w13026 = ~w13024 & ~w13025;
assign w13027 = w12692 & w13026;
assign w13028 = ~w12692 & ~w13026;
assign w13029 = ~w13027 & ~w13028;
assign w13030 = w12205 & w12217;
assign w13031 = ~w12204 & ~w13030;
assign w13032 = w13029 & w13031;
assign w13033 = ~w13029 & ~w13031;
assign w13034 = ~w13032 & ~w13033;
assign w13035 = ~w11027 & ~w12214;
assign w13036 = ~w12213 & w13035;
assign w13037 = w12213 & ~w13035;
assign w13038 = ~w12205 & ~w12217;
assign w13039 = (~w13037 & ~w12205) | (~w13037 & w16025) | (~w12205 & w16025);
assign w13040 = ~w13038 & w13039;
assign w13041 = ~w13036 & ~w13040;
assign w13042 = pi334 & ~w4854;
assign w13043 = (~w11863 & w12202) | (~w11863 & w16026) | (w12202 & w16026);
assign w13044 = pi333 & w5194;
assign w13045 = pi332 & w5714;
assign w13046 = w13044 & ~w13045;
assign w13047 = ~w13044 & w13045;
assign w13048 = ~w13046 & ~w13047;
assign w13049 = w13043 & w13048;
assign w13050 = ~w13043 & ~w13048;
assign w13051 = ~w13049 & ~w13050;
assign w13052 = ~w13042 & w13051;
assign w13053 = w13042 & ~w13051;
assign w13054 = ~w13052 & ~w13053;
assign w13055 = w13041 & ~w13054;
assign w13056 = ~w13041 & w13054;
assign w13057 = ~w13055 & ~w13056;
assign w13058 = w13034 & w13057;
assign w13059 = ~w13034 & ~w13057;
assign w13060 = ~w13058 & ~w13059;
assign w13061 = ~w12681 & w13060;
assign w13062 = w12681 & ~w13060;
assign w13063 = ~w13061 & ~w13062;
assign w13064 = w12680 & w13063;
assign w13065 = ~w12680 & ~w13063;
assign w13066 = ~w13064 & ~w13065;
assign w13067 = pi336 & w3979;
assign w13068 = ~w11845 & w12226;
assign w13069 = w3183 & ~w11842;
assign w13070 = ~w11830 & w11843;
assign w13071 = ~w13069 & w13070;
assign w13072 = ~w13068 & ~w13071;
assign w13073 = w13067 & ~w13072;
assign w13074 = ~w13067 & w13072;
assign w13075 = ~w13073 & ~w13074;
assign w13076 = pi337 & ~w3568;
assign w13077 = w11840 & ~w12227;
assign w13078 = ~w11840 & w12227;
assign w13079 = w11845 & ~w12226;
assign w13080 = (~w13078 & ~w12226) | (~w13078 & w16027) | (~w12226 & w16027);
assign w13081 = ~w13079 & w13080;
assign w13082 = ~w13077 & ~w13081;
assign w13083 = w13076 & ~w13082;
assign w13084 = ~w13076 & w13082;
assign w13085 = ~w13083 & ~w13084;
assign w13086 = w13075 & ~w13085;
assign w13087 = ~w13075 & w13085;
assign w13088 = ~w13086 & ~w13087;
assign w13089 = w13066 & w13088;
assign w13090 = ~w13066 & ~w13088;
assign w13091 = ~w13089 & ~w13090;
assign w13092 = w12679 & ~w13091;
assign w13093 = ~w12679 & w13091;
assign w13094 = ~w13092 & ~w13093;
assign w13095 = w12669 & w13094;
assign w13096 = ~w12669 & ~w13094;
assign w13097 = ~w13095 & ~w13096;
assign w13098 = w12645 & w13097;
assign w13099 = ~w12645 & ~w13097;
assign w13100 = ~w13098 & ~w13099;
assign w13101 = ~w11817 & ~w12242;
assign w13102 = ~w11818 & ~w13101;
assign w13103 = w13100 & ~w13102;
assign w13104 = ~w13100 & w13102;
assign w13105 = ~w13103 & ~w13104;
assign w13106 = ~w12245 & ~w12253;
assign w13107 = ~w12252 & ~w13106;
assign w13108 = pi343 & w1602;
assign w13109 = pi342 & ~w1865;
assign w13110 = ~w11792 & w12242;
assign w13111 = w12242 & w16028;
assign w13112 = w1865 & w11790;
assign w13113 = ~w11790 & w13109;
assign w13114 = ~w13112 & ~w13113;
assign w13115 = (~w13114 & ~w12242) | (~w13114 & w16029) | (~w12242 & w16029);
assign w13116 = ~w13111 & ~w13115;
assign w13117 = w13108 & ~w13116;
assign w13118 = ~w13108 & w13116;
assign w13119 = ~w13117 & ~w13118;
assign w13120 = w13107 & ~w13119;
assign w13121 = ~w13107 & w13119;
assign w13122 = ~w13120 & ~w13121;
assign w13123 = w13105 & w13122;
assign w13124 = ~w13105 & ~w13122;
assign w13125 = ~w13123 & ~w13124;
assign w13126 = w12644 & ~w13125;
assign w13127 = ~w12644 & w13125;
assign w13128 = ~w13126 & ~w13127;
assign w13129 = ~w12643 & ~w13128;
assign w13130 = w12643 & w13128;
assign w13131 = ~w13129 & ~w13130;
assign w13132 = w11784 & ~w12267;
assign w13133 = ~w11471 & w16030;
assign w13134 = w11783 & w12636;
assign w13135 = ~w11783 & ~w12636;
assign w13136 = ~w13133 & ~w13134;
assign w13137 = (~w13132 & ~w13136) | (~w13132 & w16031) | (~w13136 & w16031);
assign w13138 = pi347 & ~w793;
assign w13139 = (~w12247 & w12260) | (~w12247 & w16307) | (w12260 & w16307);
assign w13140 = pi345 & w1101;
assign w13141 = pi344 & w1339;
assign w13142 = w13140 & ~w13141;
assign w13143 = ~w13140 & w13141;
assign w13144 = ~w13142 & ~w13143;
assign w13145 = ~w13139 & w13144;
assign w13146 = w13139 & ~w13144;
assign w13147 = ~w13145 & ~w13146;
assign w13148 = w13138 & ~w13147;
assign w13149 = ~w13138 & w13147;
assign w13150 = ~w13148 & ~w13149;
assign w13151 = w13137 & ~w13150;
assign w13152 = ~w13137 & w13150;
assign w13153 = ~w13151 & ~w13152;
assign w13154 = w13131 & w13153;
assign w13155 = ~w13131 & ~w13153;
assign w13156 = ~w13154 & ~w13155;
assign w13157 = w12622 & w13156;
assign w13158 = ~w12622 & ~w13156;
assign w13159 = ~w13157 & ~w13158;
assign w13160 = w12618 & w13159;
assign w13161 = ~w12618 & ~w13159;
assign w13162 = ~w13160 & ~w13161;
assign w13163 = w456 & w12284;
assign w13164 = ~w466 & ~w13163;
assign w13165 = w971 & w12284;
assign w13166 = pi350 & ~w13165;
assign w13167 = ~w13164 & w13166;
assign w13168 = w13162 & w13167;
assign w13169 = ~w13162 & ~w13167;
assign w13170 = ~w13168 & ~w13169;
assign w13171 = w12613 & w13170;
assign w13172 = ~w12613 & ~w13170;
assign w13173 = ~w13171 & ~w13172;
assign w13174 = ~w12288 & ~w12292;
assign w13175 = ~pi287 & w13174;
assign w13176 = pi287 & ~w13174;
assign w13177 = ~w13175 & ~w13176;
assign w13178 = w13173 & ~w13177;
assign w13179 = ~w13173 & w13177;
assign w13180 = ~w13178 & ~w13179;
assign w13181 = ~w11757 & ~w12296;
assign w13182 = ~w13180 & w13181;
assign w13183 = w13180 & ~w13181;
assign w13184 = ~w13182 & ~w13183;
assign w13185 = w12612 & ~w13184;
assign w13186 = ~w12612 & w13184;
assign w13187 = ~w135 & ~w13185;
assign w13188 = ~w13186 & w13187;
assign w13189 = pi161 & ~w211;
assign w13190 = ~w13188 & w13189;
assign w13191 = ~pi160 & ~w12303;
assign w13192 = ~w13190 & w13191;
assign w13193 = ~pi094 & ~pi161;
assign w13194 = pi288 & w135;
assign w13195 = ~w13176 & ~w13179;
assign w13196 = pi288 & ~w13195;
assign w13197 = ~pi288 & w13195;
assign w13198 = ~w13196 & ~w13197;
assign w13199 = pi352 & w456;
assign w13200 = pi351 & w466;
assign w13201 = (~w13200 & ~w13170) | (~w13200 & w16308) | (~w13170 & w16308);
assign w13202 = w13170 & w16309;
assign w13203 = ~w13201 & ~w13202;
assign w13204 = (~w13165 & ~w13162) | (~w13165 & w16310) | (~w13162 & w16310);
assign w13205 = ~w537 & ~w13204;
assign w13206 = w537 & w13204;
assign w13207 = pi350 & ~w13206;
assign w13208 = ~w13205 & w13207;
assign w13209 = w13203 & ~w13208;
assign w13210 = ~w13203 & w13208;
assign w13211 = ~w13209 & ~w13210;
assign w13212 = (~w12617 & ~w13159) | (~w12617 & w16311) | (~w13159 & w16311);
assign w13213 = w13137 & ~w13138;
assign w13214 = ~w13137 & w13138;
assign w13215 = w13131 & w13147;
assign w13216 = ~w13131 & ~w13147;
assign w13217 = ~w13214 & ~w13215;
assign w13218 = ~w13216 & w13217;
assign w13219 = ~w13213 & ~w13218;
assign w13220 = w13212 & ~w13219;
assign w13221 = ~w13212 & w13219;
assign w13222 = ~w13220 & ~w13221;
assign w13223 = pi347 & ~w955;
assign w13224 = pi348 & ~w793;
assign w13225 = (~w12620 & ~w13156) | (~w12620 & w16312) | (~w13156 & w16312);
assign w13226 = ~w13224 & w13225;
assign w13227 = w13224 & ~w13225;
assign w13228 = ~w13226 & ~w13227;
assign w13229 = ~w13223 & w13228;
assign w13230 = w13223 & ~w13228;
assign w13231 = ~w13229 & ~w13230;
assign w13232 = w13222 & ~w13231;
assign w13233 = ~w13222 & w13231;
assign w13234 = ~w13232 & ~w13233;
assign w13235 = pi349 & ~w615;
assign w13236 = w13125 & ~w13139;
assign w13237 = ~w13125 & w13139;
assign w13238 = ~w1339 & ~w13237;
assign w13239 = ~w13236 & ~w13238;
assign w13240 = ~w1602 & ~w13239;
assign w13241 = w1602 & w13239;
assign w13242 = pi344 & ~w13240;
assign w13243 = ~w13241 & w13242;
assign w13244 = pi341 & ~w2373;
assign w13245 = pi339 & ~w3183;
assign w13246 = (w12663 & ~w13091) | (w12663 & w16313) | (~w13091 & w16313);
assign w13247 = ~w3183 & ~w13091;
assign w13248 = ~w13246 & ~w13247;
assign w13249 = ~w3568 & ~w13248;
assign w13250 = w3568 & w13248;
assign w13251 = pi338 & ~w13249;
assign w13252 = ~w13250 & w13251;
assign w13253 = ~w13061 & ~w13064;
assign w13254 = pi332 & w6283;
assign w13255 = ~w13029 & w13043;
assign w13256 = w13029 & ~w13043;
assign w13257 = ~w13255 & ~w13256;
assign w13258 = ~w13045 & w13257;
assign w13259 = ~w13255 & ~w13258;
assign w13260 = ~w13254 & ~w13259;
assign w13261 = ~w5714 & ~w13256;
assign w13262 = w13254 & ~w13255;
assign w13263 = ~w13261 & w13262;
assign w13264 = ~w13260 & ~w13263;
assign w13265 = pi333 & w5714;
assign w13266 = ~w13031 & ~w13044;
assign w13267 = w13031 & w13044;
assign w13268 = w13045 & ~w13257;
assign w13269 = (~w13267 & ~w13257) | (~w13267 & w16314) | (~w13257 & w16314);
assign w13270 = ~w13268 & w13269;
assign w13271 = ~w13266 & ~w13270;
assign w13272 = ~w13265 & ~w13271;
assign w13273 = w13265 & w13271;
assign w13274 = ~w13272 & ~w13273;
assign w13275 = ~w13264 & w13274;
assign w13276 = w13264 & ~w13274;
assign w13277 = ~w13275 & ~w13276;
assign w13278 = pi334 & w5194;
assign w13279 = w13041 & w13042;
assign w13280 = ~w13041 & ~w13042;
assign w13281 = ~w13034 & ~w13051;
assign w13282 = (~w13280 & ~w13034) | (~w13280 & w16315) | (~w13034 & w16315);
assign w13283 = ~w13281 & w13282;
assign w13284 = ~w13279 & ~w13283;
assign w13285 = ~w13278 & w13284;
assign w13286 = w13278 & ~w13284;
assign w13287 = ~w13285 & ~w13286;
assign w13288 = pi331 & ~w7108;
assign w13289 = ~w12691 & ~w13027;
assign w13290 = w13288 & ~w13289;
assign w13291 = ~w13288 & w13289;
assign w13292 = ~w13290 & ~w13291;
assign w13293 = pi330 & w7742;
assign w13294 = ~w13021 & ~w13025;
assign w13295 = w13293 & ~w13294;
assign w13296 = ~w13293 & w13294;
assign w13297 = ~w13295 & ~w13296;
assign w13298 = pi329 & ~w8367;
assign w13299 = w12999 & w13006;
assign w13300 = ~w12998 & ~w13299;
assign w13301 = pi324 & w12130;
assign w13302 = w12966 & w12977;
assign w13303 = ~w12979 & ~w13302;
assign w13304 = w13301 & ~w13303;
assign w13305 = ~w13301 & w13303;
assign w13306 = ~w13304 & ~w13305;
assign w13307 = pi156 & pi260;
assign w13308 = ~w12952 & ~w12956;
assign w13309 = ~w13307 & w13308;
assign w13310 = w13307 & ~w13308;
assign w13311 = ~w13309 & ~w13310;
assign w13312 = pi155 & pi261;
assign w13313 = ~w12711 & ~w12948;
assign w13314 = ~w13312 & ~w13313;
assign w13315 = w13312 & w13313;
assign w13316 = ~w13314 & ~w13315;
assign w13317 = pi154 & pi262;
assign w13318 = pi153 & pi263;
assign w13319 = ~w12936 & ~w12938;
assign w13320 = ~w13318 & ~w13319;
assign w13321 = w13318 & w13319;
assign w13322 = ~w13320 & ~w13321;
assign w13323 = pi150 & pi266;
assign w13324 = ~w12918 & ~w12921;
assign w13325 = w13323 & ~w13324;
assign w13326 = ~w13323 & w13324;
assign w13327 = ~w13325 & ~w13326;
assign w13328 = pi149 & pi267;
assign w13329 = pi148 & pi268;
assign w13330 = pi147 & pi269;
assign w13331 = pi146 & pi270;
assign w13332 = pi145 & pi271;
assign w13333 = ~w12880 & ~w12884;
assign w13334 = ~w13332 & w13333;
assign w13335 = w13332 & ~w13333;
assign w13336 = ~w13334 & ~w13335;
assign w13337 = pi144 & pi272;
assign w13338 = ~w12728 & ~w12876;
assign w13339 = w13337 & ~w13338;
assign w13340 = ~w13337 & w13338;
assign w13341 = ~w13339 & ~w13340;
assign w13342 = pi143 & pi273;
assign w13343 = pi142 & pi274;
assign w13344 = pi141 & pi275;
assign w13345 = ~w12856 & ~w12859;
assign w13346 = ~w13344 & w13345;
assign w13347 = w13344 & ~w13345;
assign w13348 = ~w13346 & ~w13347;
assign w13349 = pi140 & pi276;
assign w13350 = pi139 & pi277;
assign w13351 = pi138 & pi278;
assign w13352 = ~w12835 & ~w12838;
assign w13353 = ~w13351 & w13352;
assign w13354 = w13351 & ~w13352;
assign w13355 = ~w13353 & ~w13354;
assign w13356 = pi137 & pi279;
assign w13357 = ~w12827 & ~w12830;
assign w13358 = ~w13356 & w13357;
assign w13359 = w13356 & ~w13357;
assign w13360 = ~w13358 & ~w13359;
assign w13361 = pi136 & pi280;
assign w13362 = pi135 & pi281;
assign w13363 = ~w12813 & ~w12816;
assign w13364 = w13362 & w13363;
assign w13365 = ~w13362 & ~w13363;
assign w13366 = ~w13364 & ~w13365;
assign w13367 = pi134 & pi282;
assign w13368 = pi133 & pi283;
assign w13369 = pi132 & pi284;
assign w13370 = pi131 & pi285;
assign w13371 = ~w12749 & ~w12779;
assign w13372 = pi130 & pi286;
assign w13373 = pi128 & pi288;
assign w13374 = pi129 & pi287;
assign w13375 = ~w12771 & ~w13374;
assign w13376 = ~w11944 & ~w12771;
assign w13377 = w13374 & ~w13376;
assign w13378 = ~w13375 & ~w13377;
assign w13379 = w13373 & w13378;
assign w13380 = ~w13373 & ~w13378;
assign w13381 = ~w13379 & ~w13380;
assign w13382 = w13372 & w13381;
assign w13383 = ~w13372 & ~w13381;
assign w13384 = ~w13382 & ~w13383;
assign w13385 = w12758 & w12772;
assign w13386 = w12751 & ~w13385;
assign w13387 = ~w12758 & ~w12772;
assign w13388 = ~w13386 & ~w13387;
assign w13389 = ~w13384 & w13388;
assign w13390 = w13384 & ~w13388;
assign w13391 = ~w13389 & ~w13390;
assign w13392 = ~w13371 & ~w13391;
assign w13393 = w13371 & w13391;
assign w13394 = ~w13392 & ~w13393;
assign w13395 = w13370 & w13394;
assign w13396 = ~w13370 & ~w13394;
assign w13397 = ~w13395 & ~w13396;
assign w13398 = w13369 & w13397;
assign w13399 = ~w13369 & ~w13397;
assign w13400 = ~w13398 & ~w13399;
assign w13401 = ~w12743 & ~w12782;
assign w13402 = w13400 & ~w13401;
assign w13403 = ~w13400 & w13401;
assign w13404 = ~w13402 & ~w13403;
assign w13405 = w13368 & w13404;
assign w13406 = ~w13368 & ~w13404;
assign w13407 = ~w13405 & ~w13406;
assign w13408 = ~w12785 & ~w12789;
assign w13409 = w13407 & ~w13408;
assign w13410 = ~w13407 & w13408;
assign w13411 = ~w13409 & ~w13410;
assign w13412 = w13367 & w13411;
assign w13413 = ~w13367 & ~w13411;
assign w13414 = ~w13412 & ~w13413;
assign w13415 = ~w12797 & ~w12802;
assign w13416 = w13414 & ~w13415;
assign w13417 = ~w13414 & w13415;
assign w13418 = ~w13416 & ~w13417;
assign w13419 = w13366 & w13418;
assign w13420 = ~w13366 & ~w13418;
assign w13421 = ~w13419 & ~w13420;
assign w13422 = ~w12820 & ~w12824;
assign w13423 = ~w13421 & w13422;
assign w13424 = w13421 & ~w13422;
assign w13425 = ~w13423 & ~w13424;
assign w13426 = w13361 & w13425;
assign w13427 = ~w13361 & ~w13425;
assign w13428 = ~w13426 & ~w13427;
assign w13429 = w13360 & w13428;
assign w13430 = ~w13360 & ~w13428;
assign w13431 = ~w13429 & ~w13430;
assign w13432 = ~w13355 & ~w13431;
assign w13433 = w13355 & w13431;
assign w13434 = ~w13432 & ~w13433;
assign w13435 = ~w12841 & ~w12845;
assign w13436 = w13434 & ~w13435;
assign w13437 = ~w13434 & w13435;
assign w13438 = ~w13436 & ~w13437;
assign w13439 = w13350 & ~w13438;
assign w13440 = ~w13350 & w13438;
assign w13441 = ~w13439 & ~w13440;
assign w13442 = w13349 & ~w13441;
assign w13443 = ~w13349 & w13441;
assign w13444 = ~w13442 & ~w13443;
assign w13445 = ~w12848 & ~w12852;
assign w13446 = w13444 & ~w13445;
assign w13447 = ~w13444 & w13445;
assign w13448 = ~w13446 & ~w13447;
assign w13449 = ~w13348 & w13448;
assign w13450 = w13348 & ~w13448;
assign w13451 = ~w13449 & ~w13450;
assign w13452 = ~w12862 & ~w12867;
assign w13453 = ~w13451 & ~w13452;
assign w13454 = w13451 & w13452;
assign w13455 = ~w13453 & ~w13454;
assign w13456 = w13343 & w13455;
assign w13457 = ~w13343 & ~w13455;
assign w13458 = ~w13456 & ~w13457;
assign w13459 = w13342 & w13458;
assign w13460 = ~w13342 & ~w13458;
assign w13461 = ~w13459 & ~w13460;
assign w13462 = ~w12869 & ~w12873;
assign w13463 = w13461 & ~w13462;
assign w13464 = ~w13461 & w13462;
assign w13465 = ~w13463 & ~w13464;
assign w13466 = w13341 & w13465;
assign w13467 = ~w13341 & ~w13465;
assign w13468 = ~w13466 & ~w13467;
assign w13469 = w13336 & ~w13468;
assign w13470 = ~w13336 & w13468;
assign w13471 = ~w13469 & ~w13470;
assign w13472 = w13331 & ~w13471;
assign w13473 = ~w13331 & w13471;
assign w13474 = ~w13472 & ~w13473;
assign w13475 = ~w12886 & ~w12890;
assign w13476 = w13474 & ~w13475;
assign w13477 = ~w13474 & w13475;
assign w13478 = ~w13476 & ~w13477;
assign w13479 = ~w13330 & ~w13478;
assign w13480 = w13330 & w13478;
assign w13481 = ~w13479 & ~w13480;
assign w13482 = ~w12895 & ~w12897;
assign w13483 = w13481 & ~w13482;
assign w13484 = ~w13481 & w13482;
assign w13485 = ~w13483 & ~w13484;
assign w13486 = ~w12900 & ~w12906;
assign w13487 = ~w13485 & ~w13486;
assign w13488 = w13485 & w13486;
assign w13489 = ~w13487 & ~w13488;
assign w13490 = w13329 & ~w13489;
assign w13491 = ~w13329 & w13489;
assign w13492 = ~w13490 & ~w13491;
assign w13493 = ~w12911 & ~w12915;
assign w13494 = ~w13492 & ~w13493;
assign w13495 = w13492 & w13493;
assign w13496 = ~w13494 & ~w13495;
assign w13497 = w13328 & w13496;
assign w13498 = ~w13328 & ~w13496;
assign w13499 = ~w13497 & ~w13498;
assign w13500 = w13327 & w13499;
assign w13501 = ~w13327 & ~w13499;
assign w13502 = ~w13500 & ~w13501;
assign w13503 = ~w12718 & ~w12924;
assign w13504 = w13502 & ~w13503;
assign w13505 = ~w13502 & w13503;
assign w13506 = ~w13504 & ~w13505;
assign w13507 = pi151 & pi265;
assign w13508 = pi152 & pi264;
assign w13509 = w13508 & w17705;
assign w13510 = ~w12928 & w17706;
assign w13511 = ~w13509 & ~w13510;
assign w13512 = ~w13507 & ~w13511;
assign w13513 = w13507 & w13511;
assign w13514 = ~w13512 & ~w13513;
assign w13515 = w13506 & w13514;
assign w13516 = ~w13506 & ~w13514;
assign w13517 = ~w13515 & ~w13516;
assign w13518 = w13322 & ~w13517;
assign w13519 = ~w13322 & w13517;
assign w13520 = ~w13518 & ~w13519;
assign w13521 = ~w12941 & ~w12946;
assign w13522 = ~w13520 & ~w13521;
assign w13523 = w13520 & w13521;
assign w13524 = ~w13522 & ~w13523;
assign w13525 = w13317 & w13524;
assign w13526 = ~w13317 & ~w13524;
assign w13527 = ~w13525 & ~w13526;
assign w13528 = w13316 & w13527;
assign w13529 = ~w13316 & ~w13527;
assign w13530 = ~w13528 & ~w13529;
assign w13531 = w13311 & w13530;
assign w13532 = ~w13311 & ~w13530;
assign w13533 = ~w13531 & ~w13532;
assign w13534 = pi158 & pi258;
assign w13535 = pi157 & pi259;
assign w13536 = w13534 & ~w13535;
assign w13537 = ~w13534 & w13535;
assign w13538 = ~w13536 & ~w13537;
assign w13539 = w13533 & w13538;
assign w13540 = ~w13533 & ~w13538;
assign w13541 = ~w13539 & ~w13540;
assign w13542 = ~w12702 & w12959;
assign w13543 = ~w12703 & w12961;
assign w13544 = ~w12702 & ~w13543;
assign w13545 = ~w12959 & ~w13544;
assign w13546 = ~w13542 & ~w13545;
assign w13547 = w13541 & ~w13546;
assign w13548 = ~w13541 & w13546;
assign w13549 = ~w13547 & ~w13548;
assign w13550 = pi322 & w13549;
assign w13551 = w12965 & ~w12970;
assign w13552 = pi323 & w12964;
assign w13553 = ~w12969 & ~w13552;
assign w13554 = ~w13551 & ~w13553;
assign w13555 = (w13554 & ~w13549) | (w13554 & w16033) | (~w13549 & w16033);
assign w13556 = w13549 & w16034;
assign w13557 = ~w13555 & ~w13556;
assign w13558 = w13306 & w13557;
assign w13559 = ~w13306 & ~w13557;
assign w13560 = ~w13558 & ~w13559;
assign w13561 = pi325 & w11879;
assign w13562 = w12980 & ~w12984;
assign w13563 = ~w12985 & ~w13562;
assign w13564 = w13561 & ~w13563;
assign w13565 = ~w13561 & w13563;
assign w13566 = ~w13564 & ~w13565;
assign w13567 = ~w13560 & w13566;
assign w13568 = w13560 & ~w13566;
assign w13569 = ~w13567 & ~w13568;
assign w13570 = pi326 & ~w11070;
assign w13571 = ~w12989 & ~w12996;
assign w13572 = ~w12988 & ~w13571;
assign w13573 = ~w13570 & w13572;
assign w13574 = w13570 & ~w13572;
assign w13575 = ~w13573 & ~w13574;
assign w13576 = w13569 & w13575;
assign w13577 = ~w13569 & ~w13575;
assign w13578 = ~w13576 & ~w13577;
assign w13579 = ~w13300 & ~w13578;
assign w13580 = w13300 & w13578;
assign w13581 = ~w13579 & ~w13580;
assign w13582 = w13298 & ~w13581;
assign w13583 = ~w13298 & w13581;
assign w13584 = ~w13582 & ~w13583;
assign w13585 = pi328 & w8814;
assign w13586 = pi327 & ~w9784;
assign w13587 = ~w13004 & ~w13015;
assign w13588 = ~w13017 & ~w13587;
assign w13589 = ~w12999 & ~w13006;
assign w13590 = (~w13002 & ~w12999) | (~w13002 & w16035) | (~w12999 & w16035);
assign w13591 = ~w13589 & w13590;
assign w13592 = ~w13001 & ~w13591;
assign w13593 = ~w13588 & w13592;
assign w13594 = w13588 & ~w13592;
assign w13595 = ~w13593 & ~w13594;
assign w13596 = w13586 & ~w13595;
assign w13597 = ~w13586 & w13595;
assign w13598 = ~w13596 & ~w13597;
assign w13599 = w13585 & ~w13598;
assign w13600 = ~w13585 & w13598;
assign w13601 = ~w13599 & ~w13600;
assign w13602 = w13584 & w13601;
assign w13603 = ~w13584 & ~w13601;
assign w13604 = ~w13602 & ~w13603;
assign w13605 = w13297 & ~w13604;
assign w13606 = ~w13297 & w13604;
assign w13607 = ~w13605 & ~w13606;
assign w13608 = w13292 & w13607;
assign w13609 = ~w13292 & ~w13607;
assign w13610 = ~w13608 & ~w13609;
assign w13611 = w13287 & ~w13610;
assign w13612 = ~w13287 & w13610;
assign w13613 = ~w13611 & ~w13612;
assign w13614 = w13277 & w13613;
assign w13615 = ~w13277 & ~w13613;
assign w13616 = ~w13614 & ~w13615;
assign w13617 = ~w13253 & w13616;
assign w13618 = w13253 & ~w13616;
assign w13619 = ~w13617 & ~w13618;
assign w13620 = (~w13084 & w13091) | (~w13084 & w16036) | (w13091 & w16036);
assign w13621 = pi336 & ~w4708;
assign w13622 = ~pi335 & w13621;
assign w13623 = ~w13073 & w13622;
assign w13624 = ~w13063 & w13623;
assign w13625 = ~w13073 & ~w13621;
assign w13626 = ~w4708 & ~w13074;
assign w13627 = ~w13625 & ~w13626;
assign w13628 = w13075 & ~w13623;
assign w13629 = w13063 & w13628;
assign w13630 = ~w13624 & ~w13627;
assign w13631 = ~w13629 & w13630;
assign w13632 = pi337 & w3979;
assign w13633 = pi335 & ~w4854;
assign w13634 = w13632 & ~w13633;
assign w13635 = ~w13632 & w13633;
assign w13636 = ~w13634 & ~w13635;
assign w13637 = w13631 & ~w13636;
assign w13638 = ~w13631 & w13636;
assign w13639 = ~w13637 & ~w13638;
assign w13640 = w13620 & ~w13639;
assign w13641 = ~w13620 & w13639;
assign w13642 = ~w13640 & ~w13641;
assign w13643 = w13619 & w13642;
assign w13644 = ~w13619 & ~w13642;
assign w13645 = ~w13643 & ~w13644;
assign w13646 = w13252 & w13645;
assign w13647 = ~w13252 & ~w13645;
assign w13648 = ~w13646 & ~w13647;
assign w13649 = ~w13245 & ~w13648;
assign w13650 = w13245 & w13648;
assign w13651 = ~w13649 & ~w13650;
assign w13652 = pi340 & w2698;
assign w13653 = (~w12677 & ~w13097) | (~w12677 & w16037) | (~w13097 & w16037);
assign w13654 = ~w13652 & ~w13653;
assign w13655 = w13652 & w13653;
assign w13656 = ~w13654 & ~w13655;
assign w13657 = w12666 & w13091;
assign w13658 = ~w12666 & ~w13091;
assign w13659 = ~w12653 & ~w13657;
assign w13660 = ~w13658 & w13659;
assign w13661 = ~w12652 & ~w13660;
assign w13662 = w13656 & ~w13661;
assign w13663 = ~w13656 & w13661;
assign w13664 = ~w13662 & ~w13663;
assign w13665 = w13651 & ~w13664;
assign w13666 = ~w13651 & w13664;
assign w13667 = ~w13665 & ~w13666;
assign w13668 = ~w13244 & w13667;
assign w13669 = w13244 & ~w13667;
assign w13670 = ~w13668 & ~w13669;
assign w13671 = ~w13098 & ~w13103;
assign w13672 = ~w13670 & w13671;
assign w13673 = w13670 & ~w13671;
assign w13674 = ~w13672 & ~w13673;
assign w13675 = pi343 & ~w1865;
assign w13676 = ~w13107 & ~w13108;
assign w13677 = w13107 & w13108;
assign w13678 = ~w13105 & w13116;
assign w13679 = w13105 & ~w13116;
assign w13680 = ~w13678 & ~w13679;
assign w13681 = (~w13676 & w13680) | (~w13676 & w16038) | (w13680 & w16038);
assign w13682 = ~w13675 & ~w13681;
assign w13683 = w13675 & w13681;
assign w13684 = ~w13682 & ~w13683;
assign w13685 = ~w11790 & ~w13110;
assign w13686 = w13109 & ~w13685;
assign w13687 = ~w13109 & w13685;
assign w13688 = w13105 & ~w13687;
assign w13689 = pi342 & ~w2170;
assign w13690 = ~w13686 & ~w13689;
assign w13691 = ~w13688 & w13690;
assign w13692 = pi341 & w13102;
assign w13693 = ~w13097 & w13692;
assign w13694 = w13097 & ~w13692;
assign w13695 = ~w13686 & ~w13693;
assign w13696 = ~w13694 & w13695;
assign w13697 = ~w2170 & ~w13687;
assign w13698 = ~w13696 & w13697;
assign w13699 = ~w13691 & ~w13698;
assign w13700 = w13684 & ~w13699;
assign w13701 = ~w13684 & w13699;
assign w13702 = ~w13700 & ~w13701;
assign w13703 = ~w13674 & w13702;
assign w13704 = w13674 & ~w13702;
assign w13705 = ~w13703 & ~w13704;
assign w13706 = w13243 & w13705;
assign w13707 = ~w13243 & ~w13705;
assign w13708 = ~w13706 & ~w13707;
assign w13709 = pi346 & w1101;
assign w13710 = w12634 & w12638;
assign w13711 = ~w12630 & ~w12632;
assign w13712 = ~w13710 & w13711;
assign w13713 = ~w12623 & w13712;
assign w13714 = w12623 & ~w13712;
assign w13715 = w13128 & w13147;
assign w13716 = ~w13128 & ~w13147;
assign w13717 = ~w13715 & ~w13716;
assign w13718 = (~w13713 & w13717) | (~w13713 & w16039) | (w13717 & w16039);
assign w13719 = ~w13709 & ~w13718;
assign w13720 = w13709 & w13718;
assign w13721 = ~w13719 & ~w13720;
assign w13722 = pi345 & w1339;
assign w13723 = w12644 & w13140;
assign w13724 = ~w12644 & ~w13140;
assign w13725 = ~w13236 & ~w13237;
assign w13726 = ~w13141 & ~w13725;
assign w13727 = (~w13724 & ~w13725) | (~w13724 & w16040) | (~w13725 & w16040);
assign w13728 = ~w13726 & w13727;
assign w13729 = ~w13723 & ~w13728;
assign w13730 = w13722 & ~w13729;
assign w13731 = ~w13722 & w13729;
assign w13732 = ~w13730 & ~w13731;
assign w13733 = w13721 & ~w13732;
assign w13734 = ~w13721 & w13732;
assign w13735 = ~w13733 & ~w13734;
assign w13736 = w13708 & w13735;
assign w13737 = ~w13708 & ~w13735;
assign w13738 = ~w13736 & ~w13737;
assign w13739 = ~w13235 & w13738;
assign w13740 = w13235 & ~w13738;
assign w13741 = ~w13739 & ~w13740;
assign w13742 = w13234 & w13741;
assign w13743 = ~w13234 & ~w13741;
assign w13744 = ~w13742 & ~w13743;
assign w13745 = w13211 & w13744;
assign w13746 = ~w13211 & ~w13744;
assign w13747 = ~w13745 & ~w13746;
assign w13748 = w13199 & ~w13747;
assign w13749 = ~w13199 & w13747;
assign w13750 = ~w13748 & ~w13749;
assign w13751 = w13198 & ~w13750;
assign w13752 = ~w13198 & w13750;
assign w13753 = ~w13751 & ~w13752;
assign w13754 = (~w13183 & ~w13184) | (~w13183 & w16317) | (~w13184 & w16317);
assign w13755 = pi128 & pi291;
assign w13756 = pi294 & w709;
assign w13757 = ~w12310 & ~w12601;
assign w13758 = ~w13756 & w13757;
assign w13759 = w13756 & ~w13757;
assign w13760 = ~w13758 & ~w13759;
assign w13761 = pi297 & w1159;
assign w13762 = pi298 & w1220;
assign w13763 = ~w12560 & ~w12565;
assign w13764 = ~w12566 & ~w13763;
assign w13765 = ~w13762 & ~w13764;
assign w13766 = w13762 & w13764;
assign w13767 = ~w13765 & ~w13766;
assign w13768 = pi300 & w1693;
assign w13769 = pi302 & ~w2473;
assign w13770 = ~w12524 & ~w12525;
assign w13771 = ~w12533 & ~w13770;
assign w13772 = ~w13769 & ~w13771;
assign w13773 = w13769 & w13771;
assign w13774 = ~w13772 & ~w13773;
assign w13775 = pi303 & w2801;
assign w13776 = ~w12513 & ~w12517;
assign w13777 = w13775 & ~w13776;
assign w13778 = ~w13775 & w13776;
assign w13779 = ~w13777 & ~w13778;
assign w13780 = pi304 & w2925;
assign w13781 = pi306 & w3710;
assign w13782 = ~w12479 & ~w12496;
assign w13783 = ~w12480 & ~w13782;
assign w13784 = ~w13781 & w13783;
assign w13785 = w13781 & ~w13783;
assign w13786 = ~w13784 & ~w13785;
assign w13787 = pi307 & w4382;
assign w13788 = ~w12471 & ~w12476;
assign w13789 = w13787 & ~w13788;
assign w13790 = ~w13787 & w13788;
assign w13791 = ~w13789 & ~w13790;
assign w13792 = pi308 & w4539;
assign w13793 = ~w12436 & ~w12451;
assign w13794 = ~w12435 & ~w13793;
assign w13795 = pi312 & w6652;
assign w13796 = pi313 & w7268;
assign w13797 = pi315 & w9022;
assign w13798 = pi316 & w9270;
assign w13799 = pi317 & w9992;
assign w13800 = pi318 & w10753;
assign w13801 = ~w12384 & ~w12387;
assign w13802 = pi319 & w11557;
assign w13803 = ~w12376 & ~w12381;
assign w13804 = w13802 & ~w13803;
assign w13805 = ~w13802 & w13803;
assign w13806 = ~w13804 & ~w13805;
assign w13807 = w12352 & ~w12356;
assign w13808 = w12353 & ~w12355;
assign w13809 = ~w13807 & ~w13808;
assign w13810 = pi158 & w13809;
assign w13811 = ~pi158 & ~w13809;
assign w13812 = ~w13810 & ~w13811;
assign w13813 = pi321 & ~w13812;
assign w13814 = ~w12364 & ~w13813;
assign w13815 = w12364 & w13813;
assign w13816 = ~w13814 & ~w13815;
assign w13817 = ~w12366 & ~w12372;
assign w13818 = w479 & ~w13817;
assign w13819 = ~w13816 & w13818;
assign w13820 = w13816 & ~w13818;
assign w13821 = ~w13819 & ~w13820;
assign w13822 = w13806 & ~w13821;
assign w13823 = ~w13806 & w13821;
assign w13824 = ~w13822 & ~w13823;
assign w13825 = ~w13801 & ~w13824;
assign w13826 = w13801 & w13824;
assign w13827 = ~w13825 & ~w13826;
assign w13828 = w13800 & ~w13827;
assign w13829 = ~w13800 & w13827;
assign w13830 = ~w13828 & ~w13829;
assign w13831 = w13799 & ~w13830;
assign w13832 = ~w13799 & w13830;
assign w13833 = ~w13831 & ~w13832;
assign w13834 = ~w12390 & ~w12394;
assign w13835 = w13833 & ~w13834;
assign w13836 = ~w13833 & w13834;
assign w13837 = ~w13835 & ~w13836;
assign w13838 = ~w12398 & ~w12401;
assign w13839 = ~w13837 & w13838;
assign w13840 = w13837 & ~w13838;
assign w13841 = ~w13839 & ~w13840;
assign w13842 = w13798 & w13841;
assign w13843 = ~w13798 & ~w13841;
assign w13844 = ~w13842 & ~w13843;
assign w13845 = w13797 & w13844;
assign w13846 = ~w13797 & ~w13844;
assign w13847 = ~w13845 & ~w13846;
assign w13848 = ~w12346 & ~w12404;
assign w13849 = ~w13847 & w13848;
assign w13850 = w13847 & ~w13848;
assign w13851 = ~w13849 & ~w13850;
assign w13852 = pi314 & w7909;
assign w13853 = ~w12408 & ~w12411;
assign w13854 = w13852 & w13853;
assign w13855 = ~w13852 & ~w13853;
assign w13856 = ~w13854 & ~w13855;
assign w13857 = ~w13851 & ~w13856;
assign w13858 = w13851 & w13856;
assign w13859 = ~w13857 & ~w13858;
assign w13860 = ~w12415 & ~w12419;
assign w13861 = ~w13859 & w13860;
assign w13862 = w13859 & ~w13860;
assign w13863 = ~w13861 & ~w13862;
assign w13864 = w13796 & w13863;
assign w13865 = ~w13796 & ~w13863;
assign w13866 = ~w13864 & ~w13865;
assign w13867 = ~w13795 & ~w13866;
assign w13868 = w13795 & w13866;
assign w13869 = ~w13867 & ~w13868;
assign w13870 = ~w12339 & ~w12422;
assign w13871 = w13869 & w13870;
assign w13872 = ~w13869 & ~w13870;
assign w13873 = ~w13871 & ~w13872;
assign w13874 = ~w12426 & w13873;
assign w13875 = w5862 & ~w12425;
assign w13876 = w13874 & ~w13875;
assign w13877 = w6437 & ~w13876;
assign w13878 = ~w12425 & ~w13873;
assign w13879 = pi311 & ~w13878;
assign w13880 = ~w13874 & ~w13879;
assign w13881 = w13877 & ~w13880;
assign w13882 = pi311 & w6437;
assign w13883 = ~w12335 & ~w13882;
assign w13884 = w13873 & w13883;
assign w13885 = ~w5862 & w13882;
assign w13886 = ~w13873 & w13885;
assign w13887 = ~w13884 & ~w13886;
assign w13888 = ~w12426 & ~w13887;
assign w13889 = w12425 & w13873;
assign w13890 = ~w13878 & ~w13889;
assign w13891 = ~w6437 & ~w12429;
assign w13892 = ~w13890 & w13891;
assign w13893 = ~w13881 & ~w13888;
assign w13894 = ~w13892 & w13893;
assign w13895 = ~w13794 & ~w13894;
assign w13896 = w13794 & w13894;
assign w13897 = ~w13895 & ~w13896;
assign w13898 = pi310 & w5862;
assign w13899 = w13897 & w13898;
assign w13900 = ~w13897 & ~w13898;
assign w13901 = ~w13899 & ~w13900;
assign w13902 = w12452 & ~w12458;
assign w13903 = w13901 & ~w13902;
assign w13904 = ~w12452 & w12458;
assign w13905 = ~w12334 & ~w13904;
assign w13906 = w13903 & ~w13905;
assign w13907 = ~w13901 & w13902;
assign w13908 = ~w13906 & ~w13907;
assign w13909 = ~w5316 & ~w13908;
assign w13910 = pi309 & w5316;
assign w13911 = ~w13901 & ~w13904;
assign w13912 = w4539 & ~w13902;
assign w13913 = w13911 & ~w13912;
assign w13914 = w13910 & ~w13913;
assign w13915 = ~w13903 & w13914;
assign w13916 = ~w13901 & w13910;
assign w13917 = w13901 & ~w13910;
assign w13918 = w13905 & ~w13916;
assign w13919 = ~w13917 & w13918;
assign w13920 = w5316 & w13912;
assign w13921 = w13911 & w13920;
assign w13922 = ~w13919 & ~w13921;
assign w13923 = ~w13909 & w13922;
assign w13924 = ~w13915 & w13923;
assign w13925 = w13792 & w13924;
assign w13926 = ~w13792 & ~w13924;
assign w13927 = ~w13925 & ~w13926;
assign w13928 = ~w12456 & w12457;
assign w13929 = w12456 & ~w12457;
assign w13930 = w12455 & w12458;
assign w13931 = ~w12455 & ~w12458;
assign w13932 = ~w13930 & ~w13931;
assign w13933 = ~w13929 & w13932;
assign w13934 = ~w13928 & ~w13933;
assign w13935 = ~w13927 & w13934;
assign w13936 = w13927 & ~w13934;
assign w13937 = ~w13935 & ~w13936;
assign w13938 = w13791 & w13937;
assign w13939 = ~w13791 & ~w13937;
assign w13940 = ~w13938 & ~w13939;
assign w13941 = w13786 & w13940;
assign w13942 = ~w13786 & ~w13940;
assign w13943 = ~w13941 & ~w13942;
assign w13944 = ~w12497 & ~w12501;
assign w13945 = w13943 & w13944;
assign w13946 = ~w13943 & ~w13944;
assign w13947 = ~w13945 & ~w13946;
assign w13948 = pi305 & w3304;
assign w13949 = w13947 & w13948;
assign w13950 = ~w13947 & ~w13948;
assign w13951 = ~w13949 & ~w13950;
assign w13952 = ~w13780 & ~w13951;
assign w13953 = w13780 & w13951;
assign w13954 = ~w13952 & ~w13953;
assign w13955 = ~w12508 & ~w12511;
assign w13956 = w13954 & ~w13955;
assign w13957 = ~w13954 & w13955;
assign w13958 = ~w13956 & ~w13957;
assign w13959 = w13779 & ~w13958;
assign w13960 = ~w13779 & w13958;
assign w13961 = ~w13959 & ~w13960;
assign w13962 = w13774 & ~w13961;
assign w13963 = ~w13774 & w13961;
assign w13964 = ~w13962 & ~w13963;
assign w13965 = pi301 & w1954;
assign w13966 = ~w12540 & ~w12544;
assign w13967 = w13965 & w13966;
assign w13968 = ~w13965 & ~w13966;
assign w13969 = ~w13967 & ~w13968;
assign w13970 = ~w13964 & ~w13969;
assign w13971 = w13964 & w13969;
assign w13972 = ~w13970 & ~w13971;
assign w13973 = w13768 & w13972;
assign w13974 = ~w13768 & ~w13972;
assign w13975 = ~w13973 & ~w13974;
assign w13976 = ~w12328 & ~w12547;
assign w13977 = ~w13975 & ~w13976;
assign w13978 = w13975 & w13976;
assign w13979 = ~w13977 & ~w13978;
assign w13980 = pi299 & w1420;
assign w13981 = ~w12319 & ~w12551;
assign w13982 = w13980 & w13981;
assign w13983 = ~w13980 & ~w13981;
assign w13984 = ~w13982 & ~w13983;
assign w13985 = ~w13979 & w13984;
assign w13986 = w13979 & ~w13984;
assign w13987 = ~w13985 & ~w13986;
assign w13988 = w13767 & w13987;
assign w13989 = ~w13767 & ~w13987;
assign w13990 = ~w13988 & ~w13989;
assign w13991 = w13761 & w13990;
assign w13992 = ~w13761 & ~w13990;
assign w13993 = ~w13991 & ~w13992;
assign w13994 = ~w12576 & ~w12579;
assign w13995 = w13993 & ~w13994;
assign w13996 = ~w13993 & w13994;
assign w13997 = ~w13995 & ~w13996;
assign w13998 = pi296 & w855;
assign w13999 = (~w12587 & ~w12589) | (~w12587 & w16041) | (~w12589 & w16041);
assign w14000 = w13998 & w13999;
assign w14001 = ~w13998 & ~w13999;
assign w14002 = ~w14000 & ~w14001;
assign w14003 = w13997 & w14002;
assign w14004 = ~w13997 & ~w14002;
assign w14005 = ~w14003 & ~w14004;
assign w14006 = w12592 & ~w12594;
assign w14007 = w14005 & ~w14006;
assign w14008 = ~w14005 & w14006;
assign w14009 = ~w12592 & w12594;
assign w14010 = ~w12593 & ~w14009;
assign w14011 = ~w14005 & w14010;
assign w14012 = ~w14008 & ~w14011;
assign w14013 = (~w698 & ~w14005) | (~w698 & w16318) | (~w14005 & w16318);
assign w14014 = w14012 & w14013;
assign w14015 = pi295 & w698;
assign w14016 = ~w14005 & ~w14015;
assign w14017 = (w14010 & ~w14005) | (w14010 & w16319) | (~w14005 & w16319);
assign w14018 = ~w14016 & w14017;
assign w14019 = ~w14014 & ~w14018;
assign w14020 = w14005 & w14009;
assign w14021 = ~w14008 & ~w14020;
assign w14022 = w14015 & ~w14021;
assign w14023 = w698 & w709;
assign w14024 = ~w14009 & w14023;
assign w14025 = w14007 & w14024;
assign w14026 = ~w14022 & ~w14025;
assign w14027 = w14019 & w14026;
assign w14028 = w13760 & w14027;
assign w14029 = ~w13760 & ~w14027;
assign w14030 = ~w14028 & ~w14029;
assign w14031 = pi130 & w11753;
assign w14032 = (~pi130 & w12603) | (~pi130 & w16042) | (w12603 & w16042);
assign w14033 = ~pi128 & ~w646;
assign w14034 = ~w12606 & ~w14033;
assign w14035 = ~w14031 & ~w14032;
assign w14036 = ~w14034 & w14035;
assign w14037 = pi293 & w651;
assign w14038 = ~w652 & ~w14037;
assign w14039 = w11753 & w14038;
assign w14040 = ~w12604 & w14039;
assign w14041 = ~w14040 & w17707;
assign w14042 = ~w14030 & ~w14041;
assign w14043 = w14030 & w14041;
assign w14044 = ~w14042 & ~w14043;
assign w14045 = pi292 & w464;
assign w14046 = ~w12610 & ~w14045;
assign w14047 = ~pi129 & w12610;
assign w14048 = ~w14046 & ~w14047;
assign w14049 = ~w14044 & w14048;
assign w14050 = w14044 & ~w14048;
assign w14051 = ~w14049 & ~w14050;
assign w14052 = w13755 & ~w14051;
assign w14053 = ~w13755 & w14051;
assign w14054 = ~w14052 & ~w14053;
assign w14055 = ~w13754 & ~w14054;
assign w14056 = w13754 & w14054;
assign w14057 = ~w14055 & ~w14056;
assign w14058 = ~w13753 & ~w14057;
assign w14059 = w13753 & ~w14056;
assign w14060 = ~w14055 & w14059;
assign w14061 = ~w135 & ~w14058;
assign w14062 = ~w14060 & w14061;
assign w14063 = pi161 & ~w13194;
assign w14064 = ~w14062 & w14063;
assign w14065 = ~pi160 & ~w13193;
assign w14066 = ~w14064 & w14065;
assign w14067 = w8052 & w12603;
assign w14068 = ~w14031 & ~w14067;
assign w14069 = pi293 & ~w12604;
assign w14070 = ~w14068 & w14069;
assign w14071 = ~w653 & ~w14070;
assign w14072 = pi292 & ~w14071;
assign w14073 = ~pi292 & ~w14070;
assign w14074 = ~w14072 & ~w14073;
assign w14075 = pi291 & w464;
assign w14076 = w14042 & ~w14075;
assign w14077 = ~w14042 & w14075;
assign w14078 = ~w14076 & ~w14077;
assign w14079 = pi128 & pi290;
assign w14080 = w14078 & ~w14079;
assign w14081 = ~w14078 & w14079;
assign w14082 = ~w14080 & ~w14081;
assign w14083 = w14074 & w14082;
assign w14084 = ~w14074 & ~w14082;
assign w14085 = ~w14083 & ~w14084;
assign w14086 = pi353 & w456;
assign w14087 = (w13207 & w13744) | (w13207 & w16320) | (w13744 & w16320);
assign w14088 = w14086 & ~w14087;
assign w14089 = ~w14086 & w14087;
assign w14090 = ~w14088 & ~w14089;
assign w14091 = pi294 & w698;
assign w14092 = pi293 & w709;
assign w14093 = ~w14091 & w14092;
assign w14094 = w14091 & ~w14092;
assign w14095 = ~w14093 & ~w14094;
assign w14096 = ~w14095 & w17708;
assign w14097 = (w14044 & w16507) | (w14044 & w16508) | (w16507 & w16508);
assign w14098 = ~w14096 & ~w14097;
assign w14099 = w14090 & w14098;
assign w14100 = ~w14090 & ~w14098;
assign w14101 = ~w14099 & ~w14100;
assign w14102 = w13619 & w13633;
assign w14103 = ~w13619 & ~w13633;
assign w14104 = ~w14102 & ~w14103;
assign w14105 = ~w13066 & ~w13073;
assign w14106 = ~w13074 & ~w14105;
assign w14107 = w13621 & w14106;
assign w14108 = ~w14104 & ~w14107;
assign w14109 = ~w13621 & ~w14106;
assign w14110 = ~w14108 & ~w14109;
assign w14111 = pi339 & ~w3568;
assign w14112 = pi348 & ~w955;
assign w14113 = w14111 & ~w14112;
assign w14114 = ~w14111 & w14112;
assign w14115 = ~w14113 & ~w14114;
assign w14116 = pi347 & w1101;
assign w14117 = w14115 & ~w14116;
assign w14118 = ~w14115 & w14116;
assign w14119 = ~w14117 & ~w14118;
assign w14120 = w14110 & ~w14119;
assign w14121 = ~w14110 & w14119;
assign w14122 = ~w14120 & ~w14121;
assign w14123 = w13219 & ~w13738;
assign w14124 = ~w13219 & w13738;
assign w14125 = (w13223 & ~w13738) | (w13223 & w16044) | (~w13738 & w16044);
assign w14126 = ~w14123 & ~w14125;
assign w14127 = ~w13655 & ~w13667;
assign w14128 = ~w13654 & ~w14127;
assign w14129 = pi323 & w13549;
assign w14130 = w13569 & w13570;
assign w14131 = pi326 & w11879;
assign w14132 = w14130 & ~w14131;
assign w14133 = ~w14130 & w14131;
assign w14134 = ~w14132 & ~w14133;
assign w14135 = w14129 & ~w14134;
assign w14136 = ~w14129 & w14134;
assign w14137 = ~w14135 & ~w14136;
assign w14138 = w14128 & ~w14137;
assign w14139 = ~w14128 & w14137;
assign w14140 = ~w14138 & ~w14139;
assign w14141 = w13550 & ~w13553;
assign w14142 = ~w13551 & ~w14141;
assign w14143 = w13264 & w13610;
assign w14144 = ~w13263 & ~w14143;
assign w14145 = w13541 & w13543;
assign w14146 = w12960 & w13541;
assign w14147 = ~w12960 & ~w13541;
assign w14148 = ~w14146 & ~w14147;
assign w14149 = ~w12702 & ~w12961;
assign w14150 = ~w14148 & w14149;
assign w14151 = ~w14145 & ~w14150;
assign w14152 = w13534 & w14148;
assign w14153 = ~w13412 & ~w13416;
assign w14154 = pi142 & pi275;
assign w14155 = pi141 & pi276;
assign w14156 = w14154 & ~w14155;
assign w14157 = ~w14154 & w14155;
assign w14158 = ~w14156 & ~w14157;
assign w14159 = w14153 & ~w14158;
assign w14160 = ~w14153 & w14158;
assign w14161 = ~w14159 & ~w14160;
assign w14162 = pi150 & pi267;
assign w14163 = pi144 & pi273;
assign w14164 = ~w13487 & ~w13491;
assign w14165 = w14163 & ~w14164;
assign w14166 = ~w14163 & w14164;
assign w14167 = ~w14165 & ~w14166;
assign w14168 = pi146 & pi271;
assign w14169 = w14167 & ~w14168;
assign w14170 = ~w14167 & w14168;
assign w14171 = ~w14169 & ~w14170;
assign w14172 = w14162 & ~w14171;
assign w14173 = ~w14162 & w14171;
assign w14174 = ~w14172 & ~w14173;
assign w14175 = ~w13398 & ~w13402;
assign w14176 = pi131 & pi286;
assign w14177 = w14175 & ~w14176;
assign w14178 = ~w14175 & w14176;
assign w14179 = ~w14177 & ~w14178;
assign w14180 = ~w13377 & ~w13379;
assign w14181 = ~w13383 & ~w13390;
assign w14182 = w14180 & ~w14181;
assign w14183 = ~w14180 & w14181;
assign w14184 = ~w14182 & ~w14183;
assign w14185 = pi152 & pi265;
assign w14186 = w14184 & ~w14185;
assign w14187 = ~w14184 & w14185;
assign w14188 = ~w14186 & ~w14187;
assign w14189 = w14179 & w14188;
assign w14190 = ~w14179 & ~w14188;
assign w14191 = ~w14189 & ~w14190;
assign w14192 = ~w13453 & ~w13456;
assign w14193 = ~w13392 & ~w13395;
assign w14194 = w14192 & ~w14193;
assign w14195 = ~w14192 & w14193;
assign w14196 = ~w14194 & ~w14195;
assign w14197 = pi148 & pi269;
assign w14198 = pi135 & pi282;
assign w14199 = w14197 & ~w14198;
assign w14200 = ~w14197 & w14198;
assign w14201 = ~w14199 & ~w14200;
assign w14202 = ~w13364 & ~w13419;
assign w14203 = w14201 & ~w14202;
assign w14204 = ~w14201 & w14202;
assign w14205 = ~w14203 & ~w14204;
assign w14206 = w14196 & ~w14205;
assign w14207 = ~w14196 & w14205;
assign w14208 = ~w14206 & ~w14207;
assign w14209 = w14191 & ~w14208;
assign w14210 = ~w14191 & w14208;
assign w14211 = ~w14209 & ~w14210;
assign w14212 = ~w13522 & ~w13525;
assign w14213 = ~w13442 & ~w13446;
assign w14214 = pi139 & pi278;
assign w14215 = w14213 & ~w14214;
assign w14216 = ~w14213 & w14214;
assign w14217 = ~w14215 & ~w14216;
assign w14218 = pi133 & pi284;
assign w14219 = pi137 & pi280;
assign w14220 = pi157 & pi260;
assign w14221 = w14219 & ~w14220;
assign w14222 = ~w14219 & w14220;
assign w14223 = ~w14221 & ~w14222;
assign w14224 = w14218 & ~w14223;
assign w14225 = ~w14218 & w14223;
assign w14226 = ~w14224 & ~w14225;
assign w14227 = w14217 & ~w14226;
assign w14228 = ~w14217 & w14226;
assign w14229 = ~w14227 & ~w14228;
assign w14230 = w14212 & ~w14229;
assign w14231 = ~w14212 & w14229;
assign w14232 = ~w14230 & ~w14231;
assign w14233 = w14211 & w14232;
assign w14234 = ~w14211 & ~w14232;
assign w14235 = ~w14233 & ~w14234;
assign w14236 = ~w13504 & ~w13507;
assign w14237 = ~w13505 & ~w14236;
assign w14238 = pi156 & pi261;
assign w14239 = pi159 & pi258;
assign w14240 = w14238 & ~w14239;
assign w14241 = ~w14238 & w14239;
assign w14242 = ~w14240 & ~w14241;
assign w14243 = w14237 & ~w14242;
assign w14244 = ~w14237 & w14242;
assign w14245 = ~w14243 & ~w14244;
assign w14246 = w14235 & ~w14245;
assign w14247 = ~w14235 & w14245;
assign w14248 = ~w14246 & ~w14247;
assign w14249 = w14174 & w14248;
assign w14250 = ~w14174 & ~w14248;
assign w14251 = ~w14249 & ~w14250;
assign w14252 = ~w13494 & ~w13497;
assign w14253 = ~w13334 & ~w13469;
assign w14254 = w14252 & ~w14253;
assign w14255 = ~w14252 & w14253;
assign w14256 = ~w14254 & ~w14255;
assign w14257 = w14251 & ~w14256;
assign w14258 = ~w14251 & w14256;
assign w14259 = ~w14257 & ~w14258;
assign w14260 = w14161 & w14259;
assign w14261 = ~w14161 & ~w14259;
assign w14262 = ~w14260 & ~w14261;
assign w14263 = ~w13310 & ~w13531;
assign w14264 = ~w13320 & ~w13518;
assign w14265 = w14263 & ~w14264;
assign w14266 = ~w14263 & w14264;
assign w14267 = ~w14265 & ~w14266;
assign w14268 = ~w13480 & ~w13483;
assign w14269 = pi145 & pi272;
assign w14270 = w14268 & ~w14269;
assign w14271 = ~w14268 & w14269;
assign w14272 = ~w14270 & ~w14271;
assign w14273 = pi130 & pi287;
assign w14274 = ~w13359 & ~w13429;
assign w14275 = w14273 & ~w14274;
assign w14276 = ~w14273 & w14274;
assign w14277 = ~w14275 & ~w14276;
assign w14278 = w14272 & ~w14277;
assign w14279 = ~w14272 & w14277;
assign w14280 = ~w14278 & ~w14279;
assign w14281 = w14267 & ~w14280;
assign w14282 = ~w14267 & w14280;
assign w14283 = ~w14281 & ~w14282;
assign w14284 = w14262 & ~w14283;
assign w14285 = ~w14262 & w14283;
assign w14286 = ~w14284 & ~w14285;
assign w14287 = w14152 & ~w14286;
assign w14288 = ~w14152 & w14286;
assign w14289 = ~w14287 & ~w14288;
assign w14290 = ~pi259 & ~w13533;
assign w14291 = w12960 & ~w14290;
assign w14292 = w13533 & w13535;
assign w14293 = ~w14291 & ~w14292;
assign w14294 = pi154 & pi263;
assign w14295 = ~w13472 & ~w13476;
assign w14296 = ~w13459 & ~w13463;
assign w14297 = w14295 & ~w14296;
assign w14298 = ~w14295 & w14296;
assign w14299 = ~w14297 & ~w14298;
assign w14300 = w14294 & ~w14299;
assign w14301 = ~w14294 & w14299;
assign w14302 = ~w14300 & ~w14301;
assign w14303 = w14293 & w14302;
assign w14304 = ~w14293 & ~w14302;
assign w14305 = ~w14303 & ~w14304;
assign w14306 = ~w13315 & ~w13528;
assign w14307 = pi155 & pi262;
assign w14308 = w14306 & ~w14307;
assign w14309 = ~w14306 & w14307;
assign w14310 = ~w14308 & ~w14309;
assign w14311 = pi151 & pi266;
assign w14312 = pi158 & pi259;
assign w14313 = ~w13405 & ~w13409;
assign w14314 = w14312 & ~w14313;
assign w14315 = ~w14312 & w14313;
assign w14316 = ~w14314 & ~w14315;
assign w14317 = w14311 & w14316;
assign w14318 = ~w14311 & ~w14316;
assign w14319 = ~w14317 & ~w14318;
assign w14320 = ~w13325 & ~w13500;
assign w14321 = pi138 & pi279;
assign w14322 = w14320 & ~w14321;
assign w14323 = ~w14320 & w14321;
assign w14324 = ~w14322 & ~w14323;
assign w14325 = pi129 & pi288;
assign w14326 = pi140 & pi277;
assign w14327 = pi134 & pi283;
assign w14328 = w14326 & ~w14327;
assign w14329 = ~w14326 & w14327;
assign w14330 = ~w14328 & ~w14329;
assign w14331 = w14325 & ~w14330;
assign w14332 = ~w14325 & w14330;
assign w14333 = ~w14331 & ~w14332;
assign w14334 = ~w13339 & ~w13466;
assign w14335 = ~w13346 & ~w13450;
assign w14336 = pi149 & pi268;
assign w14337 = w14335 & ~w14336;
assign w14338 = ~w14335 & w14336;
assign w14339 = ~w14337 & ~w14338;
assign w14340 = pi128 & pi289;
assign w14341 = ~w13354 & ~w13433;
assign w14342 = w14340 & ~w14341;
assign w14343 = ~w14340 & w14341;
assign w14344 = ~w14342 & ~w14343;
assign w14345 = pi132 & pi285;
assign w14346 = w14344 & ~w14345;
assign w14347 = ~w14344 & w14345;
assign w14348 = ~w14346 & ~w14347;
assign w14349 = w14339 & ~w14348;
assign w14350 = ~w14339 & w14348;
assign w14351 = ~w14349 & ~w14350;
assign w14352 = w14334 & ~w14351;
assign w14353 = ~w14334 & w14351;
assign w14354 = ~w14352 & ~w14353;
assign w14355 = w14333 & w14354;
assign w14356 = ~w14333 & ~w14354;
assign w14357 = ~w14355 & ~w14356;
assign w14358 = pi136 & pi281;
assign w14359 = pi147 & pi270;
assign w14360 = w14358 & ~w14359;
assign w14361 = ~w14358 & w14359;
assign w14362 = ~w14360 & ~w14361;
assign w14363 = w14357 & ~w14362;
assign w14364 = ~w14357 & w14362;
assign w14365 = ~w14363 & ~w14364;
assign w14366 = w14324 & w14365;
assign w14367 = ~w14324 & ~w14365;
assign w14368 = ~w14366 & ~w14367;
assign w14369 = ~w13509 & ~w14368;
assign w14370 = ~w13507 & w14369;
assign w14371 = ~w13510 & w14368;
assign w14372 = w13507 & w14371;
assign w14373 = ~w14370 & ~w14372;
assign w14374 = ~w13506 & ~w14373;
assign w14375 = ~w13513 & w14371;
assign w14376 = ~w14369 & ~w14375;
assign w14377 = w13506 & ~w14370;
assign w14378 = w13511 & ~w14377;
assign w14379 = ~w14376 & ~w14378;
assign w14380 = ~w14374 & ~w14379;
assign w14381 = pi143 & pi274;
assign w14382 = ~w13424 & ~w13426;
assign w14383 = ~w13437 & ~w13440;
assign w14384 = w14382 & ~w14383;
assign w14385 = ~w14382 & w14383;
assign w14386 = ~w14384 & ~w14385;
assign w14387 = pi153 & pi264;
assign w14388 = w14386 & w14387;
assign w14389 = ~w14386 & ~w14387;
assign w14390 = ~w14388 & ~w14389;
assign w14391 = w14381 & ~w14390;
assign w14392 = ~w14381 & w14390;
assign w14393 = ~w14391 & ~w14392;
assign w14394 = w14380 & ~w14393;
assign w14395 = ~w14380 & w14393;
assign w14396 = ~w14394 & ~w14395;
assign w14397 = w14319 & ~w14396;
assign w14398 = ~w14319 & w14396;
assign w14399 = ~w14397 & ~w14398;
assign w14400 = w14310 & ~w14399;
assign w14401 = ~w14310 & w14399;
assign w14402 = ~w14400 & ~w14401;
assign w14403 = w14305 & ~w14402;
assign w14404 = ~w14305 & w14402;
assign w14405 = ~w14403 & ~w14404;
assign w14406 = w14289 & w14405;
assign w14407 = ~w14289 & ~w14405;
assign w14408 = ~w14406 & ~w14407;
assign w14409 = ~w14151 & ~w14408;
assign w14410 = w14151 & w14408;
assign w14411 = pi322 & ~w14409;
assign w14412 = ~w14410 & w14411;
assign w14413 = w14144 & ~w14412;
assign w14414 = ~w14144 & w14412;
assign w14415 = ~w14413 & ~w14414;
assign w14416 = w14142 & ~w14415;
assign w14417 = ~w14142 & w14415;
assign w14418 = ~w14416 & ~w14417;
assign w14419 = ~w13617 & ~w14102;
assign w14420 = pi328 & ~w9784;
assign w14421 = pi338 & w3979;
assign w14422 = w13572 & w13578;
assign w14423 = w14421 & ~w14422;
assign w14424 = ~w14421 & w14422;
assign w14425 = ~w14423 & ~w14424;
assign w14426 = w14420 & ~w14425;
assign w14427 = ~w14420 & w14425;
assign w14428 = ~w14426 & ~w14427;
assign w14429 = w14419 & ~w14428;
assign w14430 = ~w14419 & w14428;
assign w14431 = ~w14429 & ~w14430;
assign w14432 = w14418 & w14431;
assign w14433 = ~w14418 & ~w14431;
assign w14434 = ~w14432 & ~w14433;
assign w14435 = pi331 & w7742;
assign w14436 = pi324 & w12964;
assign w14437 = pi329 & w8814;
assign w14438 = pi334 & w5714;
assign w14439 = w14437 & ~w14438;
assign w14440 = ~w14437 & w14438;
assign w14441 = ~w14439 & ~w14440;
assign w14442 = w14436 & ~w14441;
assign w14443 = ~w14436 & w14441;
assign w14444 = ~w14442 & ~w14443;
assign w14445 = w14435 & ~w14444;
assign w14446 = ~w14435 & w14444;
assign w14447 = ~w14445 & ~w14446;
assign w14448 = w14434 & ~w14447;
assign w14449 = ~w14434 & w14447;
assign w14450 = ~w14448 & ~w14449;
assign w14451 = w14140 & ~w14450;
assign w14452 = ~w14140 & w14450;
assign w14453 = ~w14451 & ~w14452;
assign w14454 = w14126 & w14453;
assign w14455 = ~w14126 & ~w14453;
assign w14456 = ~w14454 & ~w14455;
assign w14457 = pi330 & ~w8367;
assign w14458 = ~w13650 & w13661;
assign w14459 = ~w13649 & ~w14458;
assign w14460 = w14457 & ~w14459;
assign w14461 = ~w14457 & w14459;
assign w14462 = ~w14460 & ~w14461;
assign w14463 = pi346 & w1339;
assign w14464 = (~w13683 & w13705) | (~w13683 & w16322) | (w13705 & w16322);
assign w14465 = w14463 & ~w14464;
assign w14466 = ~w14463 & w14464;
assign w14467 = ~w14465 & ~w14466;
assign w14468 = w14462 & w14467;
assign w14469 = ~w14462 & ~w14467;
assign w14470 = ~w14468 & ~w14469;
assign w14471 = pi344 & w13241;
assign w14472 = (~w14471 & ~w13705) | (~w14471 & w16323) | (~w13705 & w16323);
assign w14473 = w13581 & w13586;
assign w14474 = ~w13581 & ~w13586;
assign w14475 = ~w14473 & ~w14474;
assign w14476 = w13593 & ~w14475;
assign w14477 = ~w13585 & w14476;
assign w14478 = w13298 & w13594;
assign w14479 = w14475 & w14478;
assign w14480 = w13585 & ~w14476;
assign w14481 = ~w13593 & w14475;
assign w14482 = ~w13298 & ~w13594;
assign w14483 = ~w14481 & w14482;
assign w14484 = ~w14480 & w14483;
assign w14485 = ~w14478 & ~w14481;
assign w14486 = w13585 & ~w14482;
assign w14487 = ~w14485 & w14486;
assign w14488 = ~w14477 & ~w14479;
assign w14489 = ~w14484 & w14488;
assign w14490 = ~w14487 & w14489;
assign w14491 = w14472 & ~w14490;
assign w14492 = ~w14472 & w14490;
assign w14493 = ~w14491 & ~w14492;
assign w14494 = ~w13305 & ~w13558;
assign w14495 = pi335 & w5194;
assign w14496 = w14494 & ~w14495;
assign w14497 = ~w14494 & w14495;
assign w14498 = ~w14496 & ~w14497;
assign w14499 = pi325 & w12130;
assign w14500 = pi336 & ~w4854;
assign w14501 = w14499 & ~w14500;
assign w14502 = ~w14499 & w14500;
assign w14503 = ~w14501 & ~w14502;
assign w14504 = pi343 & ~w2170;
assign w14505 = w14503 & ~w14504;
assign w14506 = ~w14503 & w14504;
assign w14507 = ~w14505 & ~w14506;
assign w14508 = w14498 & ~w14507;
assign w14509 = ~w14498 & w14507;
assign w14510 = ~w14508 & ~w14509;
assign w14511 = w14493 & ~w14510;
assign w14512 = ~w14493 & w14510;
assign w14513 = ~w14511 & ~w14512;
assign w14514 = w14470 & w14513;
assign w14515 = ~w14470 & ~w14513;
assign w14516 = ~w14514 & ~w14515;
assign w14517 = w14456 & ~w14516;
assign w14518 = ~w14456 & w14516;
assign w14519 = ~w14517 & ~w14518;
assign w14520 = w14122 & ~w14519;
assign w14521 = ~w14122 & w14519;
assign w14522 = ~w14520 & ~w14521;
assign w14523 = w13748 & ~w14522;
assign w14524 = ~w13748 & w14522;
assign w14525 = ~w14523 & ~w14524;
assign w14526 = w14101 & w14525;
assign w14527 = ~w14101 & ~w14525;
assign w14528 = ~w14526 & ~w14527;
assign w14529 = pi349 & ~w793;
assign w14530 = w13208 & w13744;
assign w14531 = ~w13208 & ~w13744;
assign w14532 = ~w14530 & ~w14531;
assign w14533 = w14529 & w17709;
assign w14534 = w13202 & ~w14529;
assign w14535 = ~w13201 & ~w14529;
assign w14536 = pi350 & ~w615;
assign w14537 = ~pi289 & w14536;
assign w14538 = pi289 & ~w14536;
assign w14539 = ~w14537 & ~w14538;
assign w14540 = w14539 & w17710;
assign w14541 = ~w14533 & w14540;
assign w14542 = (w14532 & w16324) | (w14532 & w16325) | (w16324 & w16325);
assign w14543 = w14529 & ~w14539;
assign w14544 = w14543 & w17709;
assign w14545 = ~w14542 & ~w14544;
assign w14546 = ~w14541 & w14545;
assign w14547 = ~w14123 & ~w14124;
assign w14548 = ~w13231 & w14547;
assign w14549 = w13231 & ~w14547;
assign w14550 = ~w14548 & ~w14549;
assign w14551 = (~w13227 & w14550) | (~w13227 & w16326) | (w14550 & w16326);
assign w14552 = pi337 & ~w4708;
assign w14553 = (~w13691 & w13674) | (~w13691 & w16327) | (w13674 & w16327);
assign w14554 = pi342 & ~w2373;
assign w14555 = w14553 & ~w14554;
assign w14556 = ~w14553 & w14554;
assign w14557 = ~w14555 & ~w14556;
assign w14558 = pi340 & ~w3183;
assign w14559 = w14557 & ~w14558;
assign w14560 = ~w14557 & w14558;
assign w14561 = ~w14559 & ~w14560;
assign w14562 = w14552 & w14561;
assign w14563 = ~w14552 & ~w14561;
assign w14564 = ~w14562 & ~w14563;
assign w14565 = ~w13290 & ~w13608;
assign w14566 = ~w13295 & ~w13605;
assign w14567 = w14565 & ~w14566;
assign w14568 = ~w14565 & w14566;
assign w14569 = ~w14567 & ~w14568;
assign w14570 = ~w13564 & ~w13567;
assign w14571 = pi341 & w2698;
assign w14572 = pi344 & ~w1865;
assign w14573 = w14571 & ~w14572;
assign w14574 = ~w14571 & w14572;
assign w14575 = ~w14573 & ~w14574;
assign w14576 = ~w13579 & ~w14473;
assign w14577 = pi333 & w6283;
assign w14578 = w14576 & ~w14577;
assign w14579 = ~w14576 & w14577;
assign w14580 = ~w14578 & ~w14579;
assign w14581 = pi327 & ~w11070;
assign w14582 = w14580 & ~w14581;
assign w14583 = ~w14580 & w14581;
assign w14584 = ~w14582 & ~w14583;
assign w14585 = w14575 & w14584;
assign w14586 = ~w14575 & ~w14584;
assign w14587 = ~w14585 & ~w14586;
assign w14588 = w14570 & ~w14587;
assign w14589 = ~w14570 & w14587;
assign w14590 = ~w14588 & ~w14589;
assign w14591 = w14569 & ~w14590;
assign w14592 = ~w14569 & w14590;
assign w14593 = ~w14591 & ~w14592;
assign w14594 = w14564 & w14593;
assign w14595 = ~w14564 & ~w14593;
assign w14596 = ~w14594 & ~w14595;
assign w14597 = w13631 & w14104;
assign w14598 = ~w13631 & ~w14104;
assign w14599 = ~w14597 & ~w14598;
assign w14600 = w13632 & ~w14599;
assign w14601 = ~w13620 & ~w14600;
assign w14602 = ~w13632 & w14599;
assign w14603 = ~w14601 & ~w14602;
assign w14604 = (~w13730 & ~w13708) | (~w13730 & w16328) | (~w13708 & w16328);
assign w14605 = pi332 & ~w7108;
assign w14606 = ~w13264 & ~w13610;
assign w14607 = ~w13272 & ~w14143;
assign w14608 = ~w14606 & w14607;
assign w14609 = ~w13273 & ~w14608;
assign w14610 = w14605 & ~w14609;
assign w14611 = ~w14605 & w14609;
assign w14612 = ~w14610 & ~w14611;
assign w14613 = pi338 & w13249;
assign w14614 = ~w13646 & ~w14613;
assign w14615 = ~w13285 & ~w13616;
assign w14616 = ~w13286 & ~w14615;
assign w14617 = w14614 & ~w14616;
assign w14618 = ~w14614 & w14616;
assign w14619 = ~w14617 & ~w14618;
assign w14620 = w14612 & w14619;
assign w14621 = ~w14612 & ~w14619;
assign w14622 = ~w14620 & ~w14621;
assign w14623 = w14604 & ~w14622;
assign w14624 = ~w14604 & w14622;
assign w14625 = ~w14623 & ~w14624;
assign w14626 = w14603 & ~w14625;
assign w14627 = ~w14603 & w14625;
assign w14628 = ~w14626 & ~w14627;
assign w14629 = w14596 & ~w14628;
assign w14630 = ~w14596 & w14628;
assign w14631 = ~w14629 & ~w14630;
assign w14632 = w14551 & w14631;
assign w14633 = ~w14551 & ~w14631;
assign w14634 = ~w14632 & ~w14633;
assign w14635 = pi345 & w1602;
assign w14636 = ~w13669 & ~w13673;
assign w14637 = ~w14635 & w14636;
assign w14638 = w14635 & ~w14636;
assign w14639 = ~w14637 & ~w14638;
assign w14640 = ~w13719 & w13738;
assign w14641 = ~w13720 & ~w14640;
assign w14642 = w14639 & w14641;
assign w14643 = ~w14639 & ~w14641;
assign w14644 = ~w14642 & ~w14643;
assign w14645 = ~w13212 & w13235;
assign w14646 = w13212 & ~w13235;
assign w14647 = (~w14646 & w14550) | (~w14646 & w16329) | (w14550 & w16329);
assign w14648 = w14644 & ~w14647;
assign w14649 = ~w14644 & w14647;
assign w14650 = ~w14648 & ~w14649;
assign w14651 = w14634 & ~w14650;
assign w14652 = ~w14634 & w14650;
assign w14653 = ~w14651 & ~w14652;
assign w14654 = w14546 & ~w14653;
assign w14655 = ~w14546 & w14653;
assign w14656 = ~w14654 & ~w14655;
assign w14657 = w14528 & w14656;
assign w14658 = ~w14528 & ~w14656;
assign w14659 = ~w14657 & ~w14658;
assign w14660 = (~w14055 & ~w13753) | (~w14055 & w16047) | (~w13753 & w16047);
assign w14661 = (~w13196 & w13750) | (~w13196 & w16048) | (w13750 & w16048);
assign w14662 = ~w13974 & ~w13978;
assign w14663 = w13982 & ~w14662;
assign w14664 = ~w13982 & w14662;
assign w14665 = ~w14663 & ~w14664;
assign w14666 = ~w13991 & ~w13995;
assign w14667 = ~w13985 & w14666;
assign w14668 = w13985 & ~w14666;
assign w14669 = ~w14667 & ~w14668;
assign w14670 = ~w13867 & ~w13871;
assign w14671 = w14669 & ~w14670;
assign w14672 = ~w14669 & w14670;
assign w14673 = ~w14671 & ~w14672;
assign w14674 = w14665 & ~w14673;
assign w14675 = ~w14665 & w14673;
assign w14676 = ~w14674 & ~w14675;
assign w14677 = ~w14000 & ~w14003;
assign w14678 = (w14027 & w16509) | (w14027 & w16510) | (w16509 & w16510);
assign w14679 = ~w14677 & w17711;
assign w14680 = ~w14678 & ~w14679;
assign w14681 = pi300 & w1954;
assign w14682 = pi352 & w466;
assign w14683 = w14681 & ~w14682;
assign w14684 = ~w14681 & w14682;
assign w14685 = ~w14683 & ~w14684;
assign w14686 = ~w13945 & ~w13949;
assign w14687 = pi315 & w9270;
assign w14688 = w14686 & ~w14687;
assign w14689 = ~w14686 & w14687;
assign w14690 = ~w14688 & ~w14689;
assign w14691 = pi303 & w2925;
assign w14692 = pi305 & w3710;
assign w14693 = pi316 & w9992;
assign w14694 = ~w13925 & ~w13936;
assign w14695 = w14693 & ~w14694;
assign w14696 = ~w14693 & w14694;
assign w14697 = ~w14695 & ~w14696;
assign w14698 = ~w13862 & ~w13864;
assign w14699 = pi313 & w7909;
assign w14700 = w14698 & ~w14699;
assign w14701 = ~w14698 & w14699;
assign w14702 = ~w14700 & ~w14701;
assign w14703 = pi312 & w7268;
assign w14704 = w14702 & ~w14703;
assign w14705 = ~w14702 & w14703;
assign w14706 = ~w14704 & ~w14705;
assign w14707 = w14697 & ~w14706;
assign w14708 = ~w14697 & w14706;
assign w14709 = ~w14707 & ~w14708;
assign w14710 = w14692 & ~w14709;
assign w14711 = ~w14692 & w14709;
assign w14712 = ~w14710 & ~w14711;
assign w14713 = pi304 & w3304;
assign w14714 = pi295 & w855;
assign w14715 = ~w13840 & ~w13842;
assign w14716 = pi296 & w1159;
assign w14717 = w14715 & ~w14716;
assign w14718 = ~w14715 & w14716;
assign w14719 = ~w14717 & ~w14718;
assign w14720 = w14714 & w14719;
assign w14721 = ~w14714 & ~w14719;
assign w14722 = ~w14720 & ~w14721;
assign w14723 = w14713 & ~w14722;
assign w14724 = ~w14713 & w14722;
assign w14725 = ~w14723 & ~w14724;
assign w14726 = ~w13967 & ~w13971;
assign w14727 = pi306 & w4382;
assign w14728 = w12426 & ~w13873;
assign w14729 = ~w13877 & ~w13878;
assign w14730 = ~w13883 & ~w14729;
assign w14731 = ~w14728 & ~w14730;
assign w14732 = w14727 & ~w14731;
assign w14733 = ~w14727 & w14731;
assign w14734 = ~w14732 & ~w14733;
assign w14735 = w14726 & ~w14734;
assign w14736 = ~w14726 & w14734;
assign w14737 = ~w14735 & ~w14736;
assign w14738 = w14725 & w14737;
assign w14739 = ~w14725 & ~w14737;
assign w14740 = ~w14738 & ~w14739;
assign w14741 = ~w13789 & ~w13938;
assign w14742 = pi309 & w5862;
assign w14743 = pi299 & w1693;
assign w14744 = ~w13835 & w14743;
assign w14745 = w13835 & ~w14743;
assign w14746 = ~w14744 & ~w14745;
assign w14747 = pi308 & w5316;
assign w14748 = w14746 & ~w14747;
assign w14749 = ~w14746 & w14747;
assign w14750 = ~w14748 & ~w14749;
assign w14751 = w14742 & ~w14750;
assign w14752 = ~w14742 & w14750;
assign w14753 = ~w14751 & ~w14752;
assign w14754 = w14741 & ~w14753;
assign w14755 = ~w14741 & w14753;
assign w14756 = ~w14754 & ~w14755;
assign w14757 = w14740 & ~w14756;
assign w14758 = ~w14740 & w14756;
assign w14759 = ~w14757 & ~w14758;
assign w14760 = w14712 & w14759;
assign w14761 = ~w14712 & ~w14759;
assign w14762 = ~w14760 & ~w14761;
assign w14763 = w14691 & ~w14762;
assign w14764 = ~w14691 & w14762;
assign w14765 = ~w14763 & ~w14764;
assign w14766 = w14690 & w14765;
assign w14767 = ~w14690 & ~w14765;
assign w14768 = ~w14766 & ~w14767;
assign w14769 = ~w13953 & ~w13956;
assign w14770 = pi311 & w6652;
assign w14771 = ~w13804 & ~w13822;
assign w14772 = ~w14770 & w14771;
assign w14773 = w14770 & ~w14771;
assign w14774 = ~w14772 & ~w14773;
assign w14775 = w14769 & ~w14774;
assign w14776 = ~w14769 & w14774;
assign w14777 = ~w14775 & ~w14776;
assign w14778 = w14768 & ~w14777;
assign w14779 = ~w14768 & w14777;
assign w14780 = ~w14778 & ~w14779;
assign w14781 = w14685 & w14780;
assign w14782 = ~w14685 & ~w14780;
assign w14783 = ~w14781 & ~w14782;
assign w14784 = ~w13896 & ~w13899;
assign w14785 = pi319 & w12359;
assign w14786 = pi317 & w10753;
assign w14787 = pi320 & ~w13812;
assign w14788 = ~w13854 & ~w13858;
assign w14789 = w14787 & ~w14788;
assign w14790 = ~w14787 & w14788;
assign w14791 = ~w14789 & ~w14790;
assign w14792 = w13831 & w14791;
assign w14793 = ~w13831 & ~w14791;
assign w14794 = ~w14792 & ~w14793;
assign w14795 = w14786 & ~w14794;
assign w14796 = ~w14786 & w14794;
assign w14797 = ~w14795 & ~w14796;
assign w14798 = w14785 & ~w14797;
assign w14799 = ~w14785 & w14797;
assign w14800 = ~w14798 & ~w14799;
assign w14801 = w14784 & ~w14800;
assign w14802 = ~w14784 & w14800;
assign w14803 = ~w14801 & ~w14802;
assign w14804 = w14783 & ~w14803;
assign w14805 = ~w14783 & w14803;
assign w14806 = ~w14804 & ~w14805;
assign w14807 = pi298 & w1420;
assign w14808 = ~w13906 & ~w13914;
assign w14809 = pi318 & w11557;
assign w14810 = w14808 & ~w14809;
assign w14811 = ~w14808 & w14809;
assign w14812 = ~w14810 & ~w14811;
assign w14813 = w14807 & ~w14812;
assign w14814 = ~w14807 & w14812;
assign w14815 = ~w14813 & ~w14814;
assign w14816 = pi301 & ~w2473;
assign w14817 = pi310 & w6437;
assign w14818 = ~w13815 & ~w13818;
assign w14819 = ~w13814 & ~w14818;
assign w14820 = w14817 & ~w14819;
assign w14821 = ~w14817 & w14819;
assign w14822 = ~w14820 & ~w14821;
assign w14823 = w14816 & ~w14822;
assign w14824 = ~w14816 & w14822;
assign w14825 = ~w14823 & ~w14824;
assign w14826 = w14815 & w14825;
assign w14827 = ~w14815 & ~w14825;
assign w14828 = ~w14826 & ~w14827;
assign w14829 = ~w13766 & ~w13988;
assign w14830 = ~w13773 & ~w13962;
assign w14831 = w14829 & ~w14830;
assign w14832 = ~w14829 & w14830;
assign w14833 = ~w14831 & ~w14832;
assign w14834 = ~w13785 & ~w13941;
assign w14835 = ~pi157 & pi158;
assign w14836 = ~pi159 & w14835;
assign w14837 = ~pi156 & w14836;
assign w14838 = pi157 & ~pi158;
assign w14839 = ~pi159 & w14838;
assign w14840 = pi158 & pi159;
assign w14841 = ~w12356 & w14840;
assign w14842 = ~w14839 & ~w14841;
assign w14843 = pi156 & ~w14842;
assign w14844 = ~pi156 & ~pi158;
assign w14845 = pi159 & w14844;
assign w14846 = ~w14836 & ~w14845;
assign w14847 = w12356 & ~w14846;
assign w14848 = ~w12356 & w14839;
assign w14849 = pi159 & ~w14835;
assign w14850 = ~w14838 & w14849;
assign w14851 = ~w14837 & ~w14850;
assign w14852 = ~w14847 & w14851;
assign w14853 = ~w14848 & w14852;
assign w14854 = ~w14843 & w14853;
assign w14855 = pi321 & ~w14854;
assign w14856 = pi302 & w2801;
assign w14857 = w14855 & ~w14856;
assign w14858 = ~w14855 & w14856;
assign w14859 = ~w14857 & ~w14858;
assign w14860 = pi314 & w9022;
assign w14861 = ~w13845 & ~w13850;
assign w14862 = w14860 & ~w14861;
assign w14863 = ~w14860 & w14861;
assign w14864 = ~w14862 & ~w14863;
assign w14865 = w14859 & ~w14864;
assign w14866 = ~w14859 & w14864;
assign w14867 = ~w14865 & ~w14866;
assign w14868 = w14834 & ~w14867;
assign w14869 = ~w14834 & w14867;
assign w14870 = ~w14868 & ~w14869;
assign w14871 = w14833 & ~w14870;
assign w14872 = ~w14833 & w14870;
assign w14873 = ~w14871 & ~w14872;
assign w14874 = w14828 & ~w14873;
assign w14875 = ~w14828 & w14873;
assign w14876 = ~w14874 & ~w14875;
assign w14877 = w14806 & w14876;
assign w14878 = ~w14806 & ~w14876;
assign w14879 = ~w14877 & ~w14878;
assign w14880 = pi297 & w1220;
assign w14881 = ~w13825 & ~w13829;
assign w14882 = w14880 & ~w14881;
assign w14883 = ~w14880 & w14881;
assign w14884 = ~w14882 & ~w14883;
assign w14885 = ~w13778 & ~w13959;
assign w14886 = w14884 & ~w14885;
assign w14887 = ~w14884 & w14885;
assign w14888 = ~w14886 & ~w14887;
assign w14889 = w14879 & ~w14888;
assign w14890 = ~w14879 & w14888;
assign w14891 = ~w14889 & ~w14890;
assign w14892 = pi351 & ~w537;
assign w14893 = pi307 & w4539;
assign w14894 = w14892 & ~w14893;
assign w14895 = ~w14892 & w14893;
assign w14896 = ~w14894 & ~w14895;
assign w14897 = w14019 & w16050;
assign w14898 = (w14896 & ~w14019) | (w14896 & w16051) | (~w14019 & w16051);
assign w14899 = ~w14897 & ~w14898;
assign w14900 = w14891 & w14899;
assign w14901 = ~w14891 & ~w14899;
assign w14902 = ~w14900 & ~w14901;
assign w14903 = w14680 & ~w14902;
assign w14904 = ~w14680 & w14902;
assign w14905 = ~w14903 & ~w14904;
assign w14906 = w14676 & ~w14905;
assign w14907 = ~w14676 & w14905;
assign w14908 = ~w14906 & ~w14907;
assign w14909 = w14052 & ~w14908;
assign w14910 = ~w14052 & w14908;
assign w14911 = ~w14909 & ~w14910;
assign w14912 = w14661 & ~w14911;
assign w14913 = ~w14661 & w14911;
assign w14914 = ~w14912 & ~w14913;
assign w14915 = w14660 & ~w14914;
assign w14916 = ~w14660 & w14914;
assign w14917 = ~w14915 & ~w14916;
assign w14918 = w14659 & w14917;
assign w14919 = ~w14659 & ~w14917;
assign w14920 = ~w14918 & ~w14919;
assign w14921 = ~w135 & ~w14085;
assign w14922 = ~pi289 & w135;
assign w14923 = ~w135 & w14085;
assign w14924 = w14920 & w14923;
assign w14925 = w136 & ~w14922;
assign w14926 = (w14925 & w14920) | (w14925 & w16052) | (w14920 & w16052);
assign w14927 = ~w14924 & w14926;
assign w14928 = pi095 & ~pi160;
assign w14929 = ~pi161 & w14928;
assign w14930 = ~w14927 & ~w14929;
assign w14931 = ~pi063 & ~pi161;
assign w14932 = pi319 & ~w785;
assign w14933 = ~pi319 & w785;
assign w14934 = ~w14932 & ~w14933;
assign w14935 = pi320 & ~w777;
assign w14936 = pi321 & w456;
assign w14937 = ~pi320 & w777;
assign w14938 = ~w14935 & ~w14937;
assign w14939 = w14936 & w14938;
assign w14940 = ~w14935 & ~w14939;
assign w14941 = w14934 & ~w14940;
assign w14942 = ~w14932 & ~w14941;
assign w14943 = ~w596 & w14942;
assign w14944 = w596 & ~w14942;
assign w14945 = ~pi318 & ~w14944;
assign w14946 = ~w14943 & ~w14945;
assign w14947 = ~w773 & ~w14946;
assign w14948 = w773 & w14946;
assign w14949 = ~pi317 & ~w14948;
assign w14950 = ~w14947 & ~w14949;
assign w14951 = ~w1088 & ~w14950;
assign w14952 = w1088 & w14950;
assign w14953 = ~pi316 & ~w14952;
assign w14954 = ~w14951 & ~w14953;
assign w14955 = ~w1082 & ~w14954;
assign w14956 = w1082 & w14954;
assign w14957 = ~pi315 & ~w14956;
assign w14958 = ~w14955 & ~w14957;
assign w14959 = ~w1507 & ~w14958;
assign w14960 = w1507 & w14958;
assign w14961 = ~pi314 & ~w14960;
assign w14962 = ~w14959 & ~w14961;
assign w14963 = ~w1589 & ~w14962;
assign w14964 = w1589 & w14962;
assign w14965 = ~pi313 & ~w14964;
assign w14966 = ~w14963 & ~w14965;
assign w14967 = ~w1859 & ~w14966;
assign w14968 = w1859 & w14966;
assign w14969 = ~pi312 & ~w14968;
assign w14970 = ~w14967 & ~w14969;
assign w14971 = ~w2164 & ~w14970;
assign w14972 = w2164 & w14970;
assign w14973 = ~pi311 & ~w14972;
assign w14974 = ~w14971 & ~w14973;
assign w14975 = ~w2367 & ~w14974;
assign w14976 = w2367 & w14974;
assign w14977 = ~pi310 & ~w14976;
assign w14978 = ~w14975 & ~w14977;
assign w14979 = ~w3177 & ~w14978;
assign w14980 = w3177 & w14978;
assign w14981 = ~pi309 & ~w14980;
assign w14982 = ~w14979 & ~w14981;
assign w14983 = ~w3170 & ~w14982;
assign w14984 = w3170 & w14982;
assign w14985 = ~pi308 & ~w14984;
assign w14986 = ~w14983 & ~w14985;
assign w14987 = ~w3561 & ~w14986;
assign w14988 = w3561 & w14986;
assign w14989 = ~pi307 & ~w14988;
assign w14990 = ~w14987 & ~w14989;
assign w14991 = ~w3975 & ~w14990;
assign w14992 = w3975 & w14990;
assign w14993 = ~pi306 & ~w14992;
assign w14994 = ~w14991 & ~w14993;
assign w14995 = ~w4241 & ~w14994;
assign w14996 = w4241 & w14994;
assign w14997 = ~pi305 & ~w14996;
assign w14998 = ~w14995 & ~w14997;
assign w14999 = ~w5035 & ~w14998;
assign w15000 = w5035 & w14998;
assign w15001 = ~pi304 & ~w15000;
assign w15002 = ~w14999 & ~w15001;
assign w15003 = ~w5705 & ~w15002;
assign w15004 = w5705 & w15002;
assign w15005 = ~pi303 & ~w15004;
assign w15006 = ~w15003 & ~w15005;
assign w15007 = ~w6090 & ~w15006;
assign w15008 = w6090 & w15006;
assign w15009 = ~pi302 & ~w15008;
assign w15010 = ~w15007 & ~w15009;
assign w15011 = ~w6917 & ~w15010;
assign w15012 = w6917 & w15010;
assign w15013 = ~pi301 & ~w15012;
assign w15014 = ~w15011 & ~w15013;
assign w15015 = ~w7105 & ~w15014;
assign w15016 = w7105 & w15014;
assign w15017 = ~pi300 & ~w15016;
assign w15018 = ~w15015 & ~w15017;
assign w15019 = w7739 & ~w15018;
assign w15020 = ~w7739 & w15018;
assign w15021 = ~pi299 & ~w15020;
assign w15022 = ~w15019 & ~w15021;
assign w15023 = ~w8364 & ~w15022;
assign w15024 = w8364 & w15022;
assign w15025 = ~pi298 & ~w15024;
assign w15026 = ~w15023 & ~w15025;
assign w15027 = ~w9556 & ~w15026;
assign w15028 = w9556 & w15026;
assign w15029 = ~pi297 & ~w15028;
assign w15030 = ~w15027 & ~w15029;
assign w15031 = ~w10532 & ~w15030;
assign w15032 = w10532 & w15030;
assign w15033 = ~pi296 & ~w15032;
assign w15034 = ~w15031 & ~w15033;
assign w15035 = w10530 & ~w15034;
assign w15036 = ~w10530 & w15034;
assign w15037 = ~pi295 & ~w15036;
assign w15038 = ~w15035 & ~w15037;
assign w15039 = w11309 & ~w15038;
assign w15040 = ~w11309 & w15038;
assign w15041 = ~pi294 & ~w15040;
assign w15042 = ~w15039 & ~w15041;
assign w15043 = ~w12124 & ~w15042;
assign w15044 = w12124 & w15042;
assign w15045 = ~pi293 & ~w15044;
assign w15046 = ~w15043 & ~w15045;
assign w15047 = ~w12961 & ~w15046;
assign w15048 = w12961 & w15046;
assign w15049 = ~pi292 & ~w15048;
assign w15050 = ~w15047 & ~w15049;
assign w15051 = w14148 & ~w15050;
assign w15052 = ~w14148 & w15050;
assign w15053 = ~pi291 & ~w15052;
assign w15054 = ~w15051 & ~w15053;
assign w15055 = ~w14408 & ~w15054;
assign w15056 = w14408 & w15054;
assign w15057 = ~w15055 & ~w15056;
assign w15058 = ~w135 & ~w15057;
assign w15059 = pi290 & ~w15058;
assign w15060 = ~pi290 & w15058;
assign w15061 = pi161 & ~w15059;
assign w15062 = ~w15060 & w15061;
assign w15063 = ~pi160 & ~w14931;
assign w15064 = ~w15062 & w15063;
assign w15065 = ~pi062 & ~pi161;
assign w15066 = ~w135 & ~w15051;
assign w15067 = w15053 & w15066;
assign w15068 = ~w15052 & w15066;
assign w15069 = pi291 & ~w15068;
assign w15070 = pi161 & ~w15067;
assign w15071 = ~w15069 & w15070;
assign w15072 = ~pi160 & ~w15065;
assign w15073 = ~w15071 & w15072;
assign w15074 = ~pi061 & ~pi161;
assign w15075 = ~w135 & ~w15047;
assign w15076 = w15049 & w15075;
assign w15077 = ~w15048 & w15075;
assign w15078 = pi292 & ~w15077;
assign w15079 = pi161 & ~w15076;
assign w15080 = ~w15078 & w15079;
assign w15081 = ~pi160 & ~w15074;
assign w15082 = ~w15080 & w15081;
assign w15083 = ~pi060 & ~pi161;
assign w15084 = ~w135 & ~w15043;
assign w15085 = w15045 & w15084;
assign w15086 = ~w15044 & w15084;
assign w15087 = pi293 & ~w15086;
assign w15088 = pi161 & ~w15085;
assign w15089 = ~w15087 & w15088;
assign w15090 = ~pi160 & ~w15083;
assign w15091 = ~w15089 & w15090;
assign w15092 = ~pi059 & ~pi161;
assign w15093 = ~w135 & ~w15039;
assign w15094 = w15041 & w15093;
assign w15095 = ~w15040 & w15093;
assign w15096 = pi294 & ~w15095;
assign w15097 = pi161 & ~w15094;
assign w15098 = ~w15096 & w15097;
assign w15099 = ~pi160 & ~w15092;
assign w15100 = ~w15098 & w15099;
assign w15101 = ~pi058 & ~pi161;
assign w15102 = ~w135 & ~w15035;
assign w15103 = w15037 & w15102;
assign w15104 = ~w15036 & w15102;
assign w15105 = pi295 & ~w15104;
assign w15106 = pi161 & ~w15103;
assign w15107 = ~w15105 & w15106;
assign w15108 = ~pi160 & ~w15101;
assign w15109 = ~w15107 & w15108;
assign w15110 = ~pi057 & ~pi161;
assign w15111 = ~w135 & ~w15031;
assign w15112 = w15033 & w15111;
assign w15113 = ~w15032 & w15111;
assign w15114 = pi296 & ~w15113;
assign w15115 = pi161 & ~w15112;
assign w15116 = ~w15114 & w15115;
assign w15117 = ~pi160 & ~w15110;
assign w15118 = ~w15116 & w15117;
assign w15119 = ~pi056 & ~pi161;
assign w15120 = ~w135 & ~w15027;
assign w15121 = w15029 & w15120;
assign w15122 = ~w15028 & w15120;
assign w15123 = pi297 & ~w15122;
assign w15124 = pi161 & ~w15121;
assign w15125 = ~w15123 & w15124;
assign w15126 = ~pi160 & ~w15119;
assign w15127 = ~w15125 & w15126;
assign w15128 = ~pi055 & ~pi161;
assign w15129 = ~w135 & ~w15023;
assign w15130 = w15025 & w15129;
assign w15131 = ~w15024 & w15129;
assign w15132 = pi298 & ~w15131;
assign w15133 = pi161 & ~w15130;
assign w15134 = ~w15132 & w15133;
assign w15135 = ~pi160 & ~w15128;
assign w15136 = ~w15134 & w15135;
assign w15137 = ~pi054 & ~pi161;
assign w15138 = ~w135 & ~w15019;
assign w15139 = w15021 & w15138;
assign w15140 = ~w15020 & w15138;
assign w15141 = pi299 & ~w15140;
assign w15142 = pi161 & ~w15139;
assign w15143 = ~w15141 & w15142;
assign w15144 = ~pi160 & ~w15137;
assign w15145 = ~w15143 & w15144;
assign w15146 = ~pi053 & ~pi161;
assign w15147 = ~w135 & ~w15015;
assign w15148 = w15017 & w15147;
assign w15149 = ~w15016 & w15147;
assign w15150 = pi300 & ~w15149;
assign w15151 = pi161 & ~w15148;
assign w15152 = ~w15150 & w15151;
assign w15153 = ~pi160 & ~w15146;
assign w15154 = ~w15152 & w15153;
assign w15155 = ~pi052 & ~pi161;
assign w15156 = ~w135 & ~w15011;
assign w15157 = w15013 & w15156;
assign w15158 = ~w15012 & w15156;
assign w15159 = pi301 & ~w15158;
assign w15160 = pi161 & ~w15157;
assign w15161 = ~w15159 & w15160;
assign w15162 = ~pi160 & ~w15155;
assign w15163 = ~w15161 & w15162;
assign w15164 = ~pi051 & ~pi161;
assign w15165 = ~w135 & ~w15007;
assign w15166 = w15009 & w15165;
assign w15167 = ~w15008 & w15165;
assign w15168 = pi302 & ~w15167;
assign w15169 = pi161 & ~w15166;
assign w15170 = ~w15168 & w15169;
assign w15171 = ~pi160 & ~w15164;
assign w15172 = ~w15170 & w15171;
assign w15173 = ~pi050 & ~pi161;
assign w15174 = ~w135 & ~w15003;
assign w15175 = w15005 & w15174;
assign w15176 = ~w15004 & w15174;
assign w15177 = pi303 & ~w15176;
assign w15178 = pi161 & ~w15175;
assign w15179 = ~w15177 & w15178;
assign w15180 = ~pi160 & ~w15173;
assign w15181 = ~w15179 & w15180;
assign w15182 = ~pi049 & ~pi161;
assign w15183 = ~w135 & ~w14999;
assign w15184 = ~w15000 & w15183;
assign w15185 = pi304 & ~w15184;
assign w15186 = ~pi304 & w15184;
assign w15187 = pi161 & ~w15185;
assign w15188 = ~w15186 & w15187;
assign w15189 = ~pi160 & ~w15182;
assign w15190 = ~w15188 & w15189;
assign w15191 = ~pi048 & ~pi161;
assign w15192 = ~w135 & ~w14995;
assign w15193 = w14997 & w15192;
assign w15194 = ~w14996 & w15192;
assign w15195 = pi305 & ~w15194;
assign w15196 = pi161 & ~w15193;
assign w15197 = ~w15195 & w15196;
assign w15198 = ~pi160 & ~w15191;
assign w15199 = ~w15197 & w15198;
assign w15200 = ~pi047 & ~pi161;
assign w15201 = ~w135 & ~w14991;
assign w15202 = ~w14992 & w15201;
assign w15203 = ~pi306 & w15202;
assign w15204 = pi306 & ~w15202;
assign w15205 = pi161 & ~w15203;
assign w15206 = ~w15204 & w15205;
assign w15207 = ~pi160 & ~w15200;
assign w15208 = ~w15206 & w15207;
assign w15209 = ~pi046 & ~pi161;
assign w15210 = ~w135 & ~w14987;
assign w15211 = ~w14988 & w15210;
assign w15212 = ~pi307 & w15211;
assign w15213 = pi307 & ~w15211;
assign w15214 = pi161 & ~w15212;
assign w15215 = ~w15213 & w15214;
assign w15216 = ~pi160 & ~w15209;
assign w15217 = ~w15215 & w15216;
assign w15218 = ~pi045 & ~pi161;
assign w15219 = ~w135 & ~w14983;
assign w15220 = w14985 & w15219;
assign w15221 = ~w14984 & w15219;
assign w15222 = pi308 & ~w15221;
assign w15223 = pi161 & ~w15220;
assign w15224 = ~w15222 & w15223;
assign w15225 = ~pi160 & ~w15218;
assign w15226 = ~w15224 & w15225;
assign w15227 = ~pi044 & ~pi161;
assign w15228 = ~w135 & ~w14979;
assign w15229 = ~w14980 & w15228;
assign w15230 = ~pi309 & w15229;
assign w15231 = pi309 & ~w15229;
assign w15232 = pi161 & ~w15230;
assign w15233 = ~w15231 & w15232;
assign w15234 = ~pi160 & ~w15227;
assign w15235 = ~w15233 & w15234;
assign w15236 = ~pi043 & ~pi161;
assign w15237 = ~w135 & ~w14975;
assign w15238 = ~w14976 & w15237;
assign w15239 = ~pi310 & w15238;
assign w15240 = pi310 & ~w15238;
assign w15241 = pi161 & ~w15239;
assign w15242 = ~w15240 & w15241;
assign w15243 = ~pi160 & ~w15236;
assign w15244 = ~w15242 & w15243;
assign w15245 = ~pi042 & ~pi161;
assign w15246 = ~w135 & ~w14971;
assign w15247 = ~w14972 & w15246;
assign w15248 = ~pi311 & w15247;
assign w15249 = pi311 & ~w15247;
assign w15250 = pi161 & ~w15248;
assign w15251 = ~w15249 & w15250;
assign w15252 = ~pi160 & ~w15245;
assign w15253 = ~w15251 & w15252;
assign w15254 = ~pi041 & ~pi161;
assign w15255 = ~w135 & ~w14967;
assign w15256 = ~w14968 & w15255;
assign w15257 = ~pi312 & w15256;
assign w15258 = pi312 & ~w15256;
assign w15259 = pi161 & ~w15257;
assign w15260 = ~w15258 & w15259;
assign w15261 = ~pi160 & ~w15254;
assign w15262 = ~w15260 & w15261;
assign w15263 = ~pi040 & ~pi161;
assign w15264 = ~w135 & ~w14963;
assign w15265 = w14965 & w15264;
assign w15266 = ~w14964 & w15264;
assign w15267 = pi313 & ~w15266;
assign w15268 = pi161 & ~w15265;
assign w15269 = ~w15267 & w15268;
assign w15270 = ~pi160 & ~w15263;
assign w15271 = ~w15269 & w15270;
assign w15272 = ~pi039 & ~pi161;
assign w15273 = ~w135 & ~w14959;
assign w15274 = w14961 & w15273;
assign w15275 = ~w14960 & w15273;
assign w15276 = pi314 & ~w15275;
assign w15277 = pi161 & ~w15274;
assign w15278 = ~w15276 & w15277;
assign w15279 = ~pi160 & ~w15272;
assign w15280 = ~w15278 & w15279;
assign w15281 = ~pi038 & ~pi161;
assign w15282 = ~w135 & ~w14955;
assign w15283 = w14957 & w15282;
assign w15284 = ~w14956 & w15282;
assign w15285 = pi315 & ~w15284;
assign w15286 = pi161 & ~w15283;
assign w15287 = ~w15285 & w15286;
assign w15288 = ~pi160 & ~w15281;
assign w15289 = ~w15287 & w15288;
assign w15290 = ~pi037 & ~pi161;
assign w15291 = ~w135 & ~w14951;
assign w15292 = ~w14952 & w15291;
assign w15293 = ~pi316 & w15292;
assign w15294 = pi316 & ~w15292;
assign w15295 = pi161 & ~w15293;
assign w15296 = ~w15294 & w15295;
assign w15297 = ~pi160 & ~w15290;
assign w15298 = ~w15296 & w15297;
assign w15299 = ~pi036 & ~pi161;
assign w15300 = ~w135 & ~w14947;
assign w15301 = w14949 & w15300;
assign w15302 = ~w14948 & w15300;
assign w15303 = pi317 & ~w15302;
assign w15304 = pi161 & ~w15301;
assign w15305 = ~w15303 & w15304;
assign w15306 = ~pi160 & ~w15299;
assign w15307 = ~w15305 & w15306;
assign w15308 = ~pi035 & ~pi161;
assign w15309 = ~w135 & ~w14943;
assign w15310 = w14945 & w15309;
assign w15311 = ~w14944 & w15309;
assign w15312 = pi318 & ~w15311;
assign w15313 = pi161 & ~w15310;
assign w15314 = ~w15312 & w15313;
assign w15315 = ~pi160 & ~w15308;
assign w15316 = ~w15314 & w15315;
assign w15317 = ~pi034 & ~pi161;
assign w15318 = ~w14934 & w14940;
assign w15319 = ~w14941 & ~w15318;
assign w15320 = ~w135 & w15319;
assign w15321 = pi161 & ~w382;
assign w15322 = ~w15320 & w15321;
assign w15323 = ~pi160 & ~w15317;
assign w15324 = ~w15322 & w15323;
assign w15325 = ~pi033 & ~pi161;
assign w15326 = ~w14936 & ~w14938;
assign w15327 = ~w14939 & ~w15326;
assign w15328 = ~w135 & w15327;
assign w15329 = pi161 & ~w348;
assign w15330 = ~w15328 & w15329;
assign w15331 = ~pi160 & ~w15325;
assign w15332 = ~w15330 & w15331;
assign w15333 = ~pi032 & ~pi161;
assign w15334 = pi258 & w448;
assign w15335 = ~pi321 & w15334;
assign w15336 = pi321 & ~w15334;
assign w15337 = pi161 & ~w15335;
assign w15338 = ~w15336 & w15337;
assign w15339 = ~pi160 & ~w15333;
assign w15340 = ~w15338 & w15339;
assign w15341 = ~pi000 & ~pi161;
assign w15342 = ~pi322 & ~w448;
assign w15343 = pi322 & w448;
assign w15344 = ~w15342 & ~w15343;
assign w15345 = pi161 & ~w15344;
assign w15346 = ~pi160 & ~w15341;
assign w15347 = ~w15345 & w15346;
assign w15348 = ~pi001 & ~pi161;
assign w15349 = ~pi129 & ~pi323;
assign w15350 = pi129 & pi323;
assign w15351 = ~w15349 & ~w15350;
assign w15352 = ~w444 & ~w15351;
assign w15353 = w444 & w15351;
assign w15354 = ~w15352 & ~w15353;
assign w15355 = ~w135 & w15354;
assign w15356 = pi161 & ~w245;
assign w15357 = ~w15355 & w15356;
assign w15358 = ~pi160 & ~w15348;
assign w15359 = ~w15357 & w15358;
assign w15360 = ~pi002 & ~pi161;
assign w15361 = pi130 & pi324;
assign w15362 = ~pi130 & ~pi324;
assign w15363 = ~w15361 & ~w15362;
assign w15364 = ~w15350 & ~w15353;
assign w15365 = ~w15363 & w15364;
assign w15366 = w15363 & ~w15364;
assign w15367 = ~w15365 & ~w15366;
assign w15368 = ~w135 & w15367;
assign w15369 = pi161 & ~w279;
assign w15370 = ~w15368 & w15369;
assign w15371 = ~pi160 & ~w15360;
assign w15372 = ~w15370 & w15371;
assign w15373 = ~pi003 & ~pi161;
assign w15374 = ~w15361 & ~w15366;
assign w15375 = ~pi325 & w15374;
assign w15376 = pi325 & ~w15374;
assign w15377 = ~w15375 & ~w15376;
assign w15378 = pi131 & w15377;
assign w15379 = ~pi131 & ~w15377;
assign w15380 = ~w15378 & ~w15379;
assign w15381 = ~w135 & w15380;
assign w15382 = pi161 & ~w313;
assign w15383 = ~w15381 & w15382;
assign w15384 = ~pi160 & ~w15373;
assign w15385 = ~w15383 & w15384;
assign w15386 = ~pi004 & ~pi161;
assign w15387 = pi132 & pi326;
assign w15388 = ~pi132 & ~pi326;
assign w15389 = ~w15387 & ~w15388;
assign w15390 = ~w15376 & ~w15378;
assign w15391 = ~w135 & ~w15390;
assign w15392 = pi132 & w135;
assign w15393 = ~w15391 & ~w15392;
assign w15394 = w15389 & w15393;
assign w15395 = ~w15389 & ~w15393;
assign w15396 = pi161 & ~w15394;
assign w15397 = ~w15395 & w15396;
assign w15398 = ~pi160 & ~w15386;
assign w15399 = ~w15397 & w15398;
assign w15400 = ~pi005 & ~pi161;
assign w15401 = ~w15388 & ~w15390;
assign w15402 = ~w15387 & ~w15401;
assign w15403 = ~pi327 & w15402;
assign w15404 = pi327 & ~w15402;
assign w15405 = ~w15403 & ~w15404;
assign w15406 = ~pi133 & ~w15405;
assign w15407 = pi133 & w15405;
assign w15408 = ~w15406 & ~w15407;
assign w15409 = ~w135 & w15408;
assign w15410 = pi161 & ~w327;
assign w15411 = ~w15409 & w15410;
assign w15412 = ~pi160 & ~w15400;
assign w15413 = ~w15411 & w15412;
assign w15414 = ~pi006 & ~pi161;
assign w15415 = ~w15404 & ~w15407;
assign w15416 = ~pi328 & w15415;
assign w15417 = pi328 & ~w15415;
assign w15418 = ~w15416 & ~w15417;
assign w15419 = w135 & ~w15415;
assign w15420 = pi134 & ~w135;
assign w15421 = ~w15419 & ~w15420;
assign w15422 = ~w15418 & ~w15421;
assign w15423 = w15418 & w15421;
assign w15424 = pi161 & ~w15422;
assign w15425 = ~w15423 & w15424;
assign w15426 = ~pi160 & ~w15414;
assign w15427 = ~w15425 & w15426;
assign w15428 = ~pi007 & ~pi161;
assign w15429 = pi134 & ~w15416;
assign w15430 = ~w15417 & ~w15429;
assign w15431 = ~pi329 & w15430;
assign w15432 = pi329 & ~w15430;
assign w15433 = ~w15431 & ~w15432;
assign w15434 = ~pi135 & ~w15433;
assign w15435 = pi135 & w15433;
assign w15436 = ~w135 & ~w15434;
assign w15437 = ~w15435 & w15436;
assign w15438 = pi161 & ~w334;
assign w15439 = ~w15437 & w15438;
assign w15440 = ~pi160 & ~w15428;
assign w15441 = ~w15439 & w15440;
assign w15442 = ~pi008 & ~pi161;
assign w15443 = ~w15432 & ~w15435;
assign w15444 = pi330 & ~w15443;
assign w15445 = ~pi330 & w15443;
assign w15446 = ~w15444 & ~w15445;
assign w15447 = ~pi136 & ~w15446;
assign w15448 = pi136 & ~w15445;
assign w15449 = ~w15444 & w15448;
assign w15450 = ~w135 & ~w15447;
assign w15451 = ~w15449 & w15450;
assign w15452 = pi161 & ~w338;
assign w15453 = ~w15451 & w15452;
assign w15454 = ~pi160 & ~w15442;
assign w15455 = ~w15453 & w15454;
assign w15456 = ~pi009 & ~pi161;
assign w15457 = ~w15444 & ~w15448;
assign w15458 = ~pi331 & w15457;
assign w15459 = pi331 & ~w15457;
assign w15460 = ~w15458 & ~w15459;
assign w15461 = w135 & ~w15457;
assign w15462 = pi137 & ~w135;
assign w15463 = ~w15461 & ~w15462;
assign w15464 = ~w15460 & ~w15463;
assign w15465 = w15460 & w15463;
assign w15466 = pi161 & ~w15464;
assign w15467 = ~w15465 & w15466;
assign w15468 = ~pi160 & ~w15456;
assign w15469 = ~w15467 & w15468;
assign w15470 = ~pi010 & ~pi161;
assign w15471 = pi137 & ~w15458;
assign w15472 = ~w15459 & ~w15471;
assign w15473 = ~pi332 & w15472;
assign w15474 = pi332 & ~w15472;
assign w15475 = ~w15473 & ~w15474;
assign w15476 = w135 & ~w15472;
assign w15477 = pi138 & ~w135;
assign w15478 = ~w15476 & ~w15477;
assign w15479 = ~w15475 & ~w15478;
assign w15480 = w15475 & w15478;
assign w15481 = pi161 & ~w15479;
assign w15482 = ~w15480 & w15481;
assign w15483 = ~pi160 & ~w15470;
assign w15484 = ~w15482 & w15483;
assign w15485 = ~pi011 & ~pi161;
assign w15486 = pi138 & ~w15473;
assign w15487 = ~w15474 & ~w15486;
assign w15488 = ~pi333 & w15487;
assign w15489 = pi333 & ~w15487;
assign w15490 = ~w15488 & ~w15489;
assign w15491 = w135 & ~w15487;
assign w15492 = pi139 & ~w135;
assign w15493 = ~w15491 & ~w15492;
assign w15494 = ~w15490 & ~w15493;
assign w15495 = w15490 & w15493;
assign w15496 = pi161 & ~w15494;
assign w15497 = ~w15495 & w15496;
assign w15498 = ~pi160 & ~w15485;
assign w15499 = ~w15497 & w15498;
assign w15500 = ~pi012 & ~pi161;
assign w15501 = pi139 & ~w15488;
assign w15502 = ~w15489 & ~w15501;
assign w15503 = ~pi334 & w15502;
assign w15504 = pi334 & ~w15502;
assign w15505 = ~w15503 & ~w15504;
assign w15506 = w135 & ~w15502;
assign w15507 = pi140 & ~w135;
assign w15508 = ~w15506 & ~w15507;
assign w15509 = ~w15505 & ~w15508;
assign w15510 = w15505 & w15508;
assign w15511 = pi161 & ~w15509;
assign w15512 = ~w15510 & w15511;
assign w15513 = ~pi160 & ~w15500;
assign w15514 = ~w15512 & w15513;
assign w15515 = ~pi013 & ~pi161;
assign w15516 = pi140 & ~w15503;
assign w15517 = ~w15504 & ~w15516;
assign w15518 = ~pi335 & w15517;
assign w15519 = pi335 & ~w15517;
assign w15520 = ~w15518 & ~w15519;
assign w15521 = w135 & ~w15517;
assign w15522 = pi141 & ~w135;
assign w15523 = ~w15521 & ~w15522;
assign w15524 = ~w15520 & ~w15523;
assign w15525 = w15520 & w15523;
assign w15526 = pi161 & ~w15524;
assign w15527 = ~w15525 & w15526;
assign w15528 = ~pi160 & ~w15515;
assign w15529 = ~w15527 & w15528;
assign w15530 = ~pi014 & ~pi161;
assign w15531 = pi141 & ~w15518;
assign w15532 = ~w15519 & ~w15531;
assign w15533 = ~pi336 & w15532;
assign w15534 = pi336 & ~w15532;
assign w15535 = ~w15533 & ~w15534;
assign w15536 = w135 & ~w15532;
assign w15537 = pi142 & ~w135;
assign w15538 = ~w15536 & ~w15537;
assign w15539 = ~w15535 & ~w15538;
assign w15540 = w15535 & w15538;
assign w15541 = pi161 & ~w15539;
assign w15542 = ~w15540 & w15541;
assign w15543 = ~pi160 & ~w15530;
assign w15544 = ~w15542 & w15543;
assign w15545 = ~pi015 & ~pi161;
assign w15546 = pi142 & ~w15533;
assign w15547 = ~w15534 & ~w15546;
assign w15548 = ~pi337 & w15547;
assign w15549 = pi337 & ~w15547;
assign w15550 = ~w15548 & ~w15549;
assign w15551 = w135 & ~w15547;
assign w15552 = pi143 & ~w135;
assign w15553 = ~w15551 & ~w15552;
assign w15554 = ~w15550 & ~w15553;
assign w15555 = w15550 & w15553;
assign w15556 = pi161 & ~w15554;
assign w15557 = ~w15555 & w15556;
assign w15558 = ~pi160 & ~w15545;
assign w15559 = ~w15557 & w15558;
assign w15560 = ~pi016 & ~pi161;
assign w15561 = pi143 & ~w15548;
assign w15562 = ~w15549 & ~w15561;
assign w15563 = ~pi338 & w15562;
assign w15564 = pi338 & ~w15562;
assign w15565 = ~w15563 & ~w15564;
assign w15566 = w135 & ~w15562;
assign w15567 = pi144 & ~w135;
assign w15568 = ~w15566 & ~w15567;
assign w15569 = ~w15565 & ~w15568;
assign w15570 = w15565 & w15568;
assign w15571 = pi161 & ~w15569;
assign w15572 = ~w15570 & w15571;
assign w15573 = ~pi160 & ~w15560;
assign w15574 = ~w15572 & w15573;
assign w15575 = ~pi017 & ~pi161;
assign w15576 = pi144 & ~w15563;
assign w15577 = ~w15564 & ~w15576;
assign w15578 = ~pi339 & w15577;
assign w15579 = pi339 & ~w15577;
assign w15580 = ~w15578 & ~w15579;
assign w15581 = w135 & ~w15577;
assign w15582 = pi145 & ~w135;
assign w15583 = ~w15581 & ~w15582;
assign w15584 = ~w15580 & ~w15583;
assign w15585 = w15580 & w15583;
assign w15586 = pi161 & ~w15584;
assign w15587 = ~w15585 & w15586;
assign w15588 = ~pi160 & ~w15575;
assign w15589 = ~w15587 & w15588;
assign w15590 = ~pi018 & ~pi161;
assign w15591 = pi145 & ~w15578;
assign w15592 = ~w15579 & ~w15591;
assign w15593 = ~pi340 & w15592;
assign w15594 = pi340 & ~w15592;
assign w15595 = ~w15593 & ~w15594;
assign w15596 = w135 & ~w15592;
assign w15597 = pi146 & ~w135;
assign w15598 = ~w15596 & ~w15597;
assign w15599 = ~w15595 & ~w15598;
assign w15600 = w15595 & w15598;
assign w15601 = pi161 & ~w15599;
assign w15602 = ~w15600 & w15601;
assign w15603 = ~pi160 & ~w15590;
assign w15604 = ~w15602 & w15603;
assign w15605 = ~pi019 & ~pi161;
assign w15606 = pi146 & ~w15593;
assign w15607 = ~w15594 & ~w15606;
assign w15608 = ~pi341 & w15607;
assign w15609 = pi341 & ~w15607;
assign w15610 = ~w15608 & ~w15609;
assign w15611 = w135 & ~w15607;
assign w15612 = pi147 & ~w135;
assign w15613 = ~w15611 & ~w15612;
assign w15614 = ~w15610 & ~w15613;
assign w15615 = w15610 & w15613;
assign w15616 = pi161 & ~w15614;
assign w15617 = ~w15615 & w15616;
assign w15618 = ~pi160 & ~w15605;
assign w15619 = ~w15617 & w15618;
assign w15620 = ~pi020 & ~pi161;
assign w15621 = pi147 & ~w15608;
assign w15622 = ~w15609 & ~w15621;
assign w15623 = ~pi342 & w15622;
assign w15624 = pi342 & ~w15622;
assign w15625 = ~w15623 & ~w15624;
assign w15626 = w135 & ~w15622;
assign w15627 = pi148 & ~w135;
assign w15628 = ~w15626 & ~w15627;
assign w15629 = ~w15625 & ~w15628;
assign w15630 = w15625 & w15628;
assign w15631 = pi161 & ~w15629;
assign w15632 = ~w15630 & w15631;
assign w15633 = ~pi160 & ~w15620;
assign w15634 = ~w15632 & w15633;
assign w15635 = ~pi021 & ~pi161;
assign w15636 = pi148 & ~w15623;
assign w15637 = ~w15624 & ~w15636;
assign w15638 = ~pi343 & w15637;
assign w15639 = pi343 & ~w15637;
assign w15640 = ~w15638 & ~w15639;
assign w15641 = w135 & ~w15637;
assign w15642 = pi149 & ~w135;
assign w15643 = ~w15641 & ~w15642;
assign w15644 = ~w15640 & ~w15643;
assign w15645 = w15640 & w15643;
assign w15646 = pi161 & ~w15644;
assign w15647 = ~w15645 & w15646;
assign w15648 = ~pi160 & ~w15635;
assign w15649 = ~w15647 & w15648;
assign w15650 = ~pi022 & ~pi161;
assign w15651 = pi149 & ~w15638;
assign w15652 = ~w15639 & ~w15651;
assign w15653 = ~pi344 & w15652;
assign w15654 = pi344 & ~w15652;
assign w15655 = ~w15653 & ~w15654;
assign w15656 = w135 & ~w15652;
assign w15657 = pi150 & ~w135;
assign w15658 = ~w15656 & ~w15657;
assign w15659 = ~w15655 & ~w15658;
assign w15660 = w15655 & w15658;
assign w15661 = pi161 & ~w15659;
assign w15662 = ~w15660 & w15661;
assign w15663 = ~pi160 & ~w15650;
assign w15664 = ~w15662 & w15663;
assign w15665 = ~pi023 & ~pi161;
assign w15666 = pi150 & ~w15653;
assign w15667 = ~w15654 & ~w15666;
assign w15668 = ~pi345 & w15667;
assign w15669 = pi345 & ~w15667;
assign w15670 = ~w15668 & ~w15669;
assign w15671 = w135 & ~w15667;
assign w15672 = pi151 & ~w135;
assign w15673 = ~w15671 & ~w15672;
assign w15674 = ~w15670 & ~w15673;
assign w15675 = w15670 & w15673;
assign w15676 = pi161 & ~w15674;
assign w15677 = ~w15675 & w15676;
assign w15678 = ~pi160 & ~w15665;
assign w15679 = ~w15677 & w15678;
assign w15680 = ~pi024 & ~pi161;
assign w15681 = pi151 & ~w15668;
assign w15682 = ~w15669 & ~w15681;
assign w15683 = ~pi346 & w15682;
assign w15684 = pi346 & ~w15682;
assign w15685 = ~w15683 & ~w15684;
assign w15686 = w135 & ~w15682;
assign w15687 = pi152 & ~w135;
assign w15688 = ~w15686 & ~w15687;
assign w15689 = ~w15685 & ~w15688;
assign w15690 = w15685 & w15688;
assign w15691 = pi161 & ~w15689;
assign w15692 = ~w15690 & w15691;
assign w15693 = ~pi160 & ~w15680;
assign w15694 = ~w15692 & w15693;
assign w15695 = ~pi025 & ~pi161;
assign w15696 = pi152 & ~w15683;
assign w15697 = ~w15684 & ~w15696;
assign w15698 = ~pi347 & w15697;
assign w15699 = pi347 & ~w15697;
assign w15700 = ~w15698 & ~w15699;
assign w15701 = w135 & ~w15697;
assign w15702 = pi153 & ~w135;
assign w15703 = ~w15701 & ~w15702;
assign w15704 = ~w15700 & ~w15703;
assign w15705 = w15700 & w15703;
assign w15706 = pi161 & ~w15704;
assign w15707 = ~w15705 & w15706;
assign w15708 = ~pi160 & ~w15695;
assign w15709 = ~w15707 & w15708;
assign w15710 = ~pi026 & ~pi161;
assign w15711 = pi153 & ~w15698;
assign w15712 = ~w15699 & ~w15711;
assign w15713 = ~pi348 & w15712;
assign w15714 = pi348 & ~w15712;
assign w15715 = ~w15713 & ~w15714;
assign w15716 = w135 & ~w15712;
assign w15717 = pi154 & ~w135;
assign w15718 = ~w15716 & ~w15717;
assign w15719 = ~w15715 & ~w15718;
assign w15720 = w15715 & w15718;
assign w15721 = pi161 & ~w15719;
assign w15722 = ~w15720 & w15721;
assign w15723 = ~pi160 & ~w15710;
assign w15724 = ~w15722 & w15723;
assign w15725 = ~pi027 & ~pi161;
assign w15726 = pi154 & ~w15713;
assign w15727 = ~w15714 & ~w15726;
assign w15728 = ~pi349 & w15727;
assign w15729 = pi349 & ~w15727;
assign w15730 = ~w15728 & ~w15729;
assign w15731 = w135 & ~w15727;
assign w15732 = pi155 & ~w135;
assign w15733 = ~w15731 & ~w15732;
assign w15734 = ~w15730 & ~w15733;
assign w15735 = w15730 & w15733;
assign w15736 = pi161 & ~w15734;
assign w15737 = ~w15735 & w15736;
assign w15738 = ~pi160 & ~w15725;
assign w15739 = ~w15737 & w15738;
assign w15740 = ~pi028 & ~pi161;
assign w15741 = pi155 & ~w15728;
assign w15742 = ~w15729 & ~w15741;
assign w15743 = ~pi350 & w15742;
assign w15744 = pi350 & ~w15742;
assign w15745 = ~w15743 & ~w15744;
assign w15746 = w135 & ~w15742;
assign w15747 = pi156 & ~w135;
assign w15748 = ~w15746 & ~w15747;
assign w15749 = ~w15745 & ~w15748;
assign w15750 = w15745 & w15748;
assign w15751 = pi161 & ~w15749;
assign w15752 = ~w15750 & w15751;
assign w15753 = ~pi160 & ~w15740;
assign w15754 = ~w15752 & w15753;
assign w15755 = ~pi029 & ~pi161;
assign w15756 = pi156 & ~w15743;
assign w15757 = ~w15744 & ~w15756;
assign w15758 = ~pi351 & w15757;
assign w15759 = pi351 & ~w15757;
assign w15760 = ~w15758 & ~w15759;
assign w15761 = w135 & ~w15757;
assign w15762 = pi157 & ~w135;
assign w15763 = ~w15761 & ~w15762;
assign w15764 = ~w15760 & ~w15763;
assign w15765 = w15760 & w15763;
assign w15766 = pi161 & ~w15764;
assign w15767 = ~w15765 & w15766;
assign w15768 = ~pi160 & ~w15755;
assign w15769 = ~w15767 & w15768;
assign w15770 = ~pi030 & ~pi161;
assign w15771 = pi157 & ~w15758;
assign w15772 = ~w15759 & ~w15771;
assign w15773 = pi352 & ~w15772;
assign w15774 = ~pi352 & w15772;
assign w15775 = ~w15773 & ~w15774;
assign w15776 = ~pi158 & ~w15775;
assign w15777 = pi158 & ~w15774;
assign w15778 = ~w15773 & w15777;
assign w15779 = ~w135 & ~w15776;
assign w15780 = ~w15778 & w15779;
assign w15781 = pi161 & ~w317;
assign w15782 = ~w15780 & w15781;
assign w15783 = ~pi160 & ~w15770;
assign w15784 = ~w15782 & w15783;
assign w15785 = ~pi031 & ~pi161;
assign w15786 = ~w15773 & ~w15777;
assign w15787 = pi159 & ~w15786;
assign w15788 = ~pi159 & w15786;
assign w15789 = ~w135 & ~w15787;
assign w15790 = ~w15788 & w15789;
assign w15791 = pi353 & ~w15790;
assign w15792 = ~pi353 & w15790;
assign w15793 = pi161 & ~w15791;
assign w15794 = ~w15792 & w15793;
assign w15795 = ~pi160 & ~w15785;
assign w15796 = ~w15794 & w15795;
assign w15797 = w585 & w513;
assign w15798 = ~w477 & ~pi131;
assign w15799 = w593 & ~pi259;
assign w15800 = w586 & w531;
assign w15801 = w462 & ~pi262;
assign w15802 = ~w462 & ~w753;
assign w15803 = w915 & ~w910;
assign w15804 = ~w767 & ~w746;
assign w15805 = ~w1034 & ~w908;
assign w15806 = (~w845 & w868) | (~w845 & w16053) | (w868 & w16053);
assign w15807 = ~w863 & w16054;
assign w15808 = w1039 & ~w1038;
assign w15809 = ~w1280 & ~w1512;
assign w15810 = w1280 & pi259;
assign w15811 = ~w1501 & ~w1500;
assign w15812 = ~w1314 & w1318;
assign w15813 = ~w1311 & ~w1309;
assign w15814 = w1045 & ~w1301;
assign w15815 = ~w1304 & ~w1303;
assign w15816 = ~w1045 & w1301;
assign w15817 = ~w1076 & w16330;
assign w15818 = w1519 & ~w1565;
assign w15819 = ~w1809 & ~w1812;
assign w15820 = w1830 & ~w1831;
assign w15821 = ~w1702 & w1673;
assign w15822 = ~w1976 & ~w1981;
assign w15823 = w698 & w855;
assign w15824 = w1734 & ~w1731;
assign w15825 = ~w1772 & ~w2058;
assign w15826 = w1772 & pi259;
assign w15827 = w1842 & ~w1839;
assign w15828 = w1788 & ~w1799;
assign w15829 = ~w1788 & w1799;
assign w15830 = ~w1796 & ~w1795;
assign w15831 = w1828 & w2125;
assign w15832 = ~w1828 & ~w2125;
assign w15833 = ~w1846 & ~w1850;
assign w15834 = ~pi259 & w2143;
assign w15835 = w2113 & w2277;
assign w15836 = ~w2113 & ~w2277;
assign w15837 = w2314 & ~w2317;
assign w15838 = (w1937 & ~w1966) | (w1937 & w16055) | (~w1966 & w16055);
assign w15839 = ~w2133 & w16511;
assign w15840 = (~w2113 & ~w2321) | (~w2113 & w15836) | (~w2321 & w15836);
assign w15841 = w2328 & w16620;
assign w15842 = (~w2636 & ~w2328) | (~w2636 & w16621) | (~w2328 & w16621);
assign w15843 = w3103 & ~w3102;
assign w15844 = w2267 & ~w2266;
assign w15845 = w3136 & ~w3135;
assign w15846 = ~w2363 & w2676;
assign w15847 = (w3160 & w16056) | (w3160 & w16057) | (w16056 & w16057);
assign w15848 = ~w2681 & w17712;
assign w15849 = w2742 & ~w955;
assign w15850 = (w3221 & w16331) | (w3221 & w16332) | (w16331 & w16332);
assign w15851 = ~w3220 & w17713;
assign w15852 = (~w2961 & w2897) | (~w2961 & w16058) | (w2897 & w16058);
assign w15853 = ~w2901 & ~w2957;
assign w15854 = ~w2933 & ~w2905;
assign w15855 = (~w2903 & w2904) | (~w2903 & w16059) | (w2904 & w16059);
assign w15856 = ~w466 & ~w3404;
assign w15857 = w3112 & ~w3117;
assign w15858 = w3062 & ~w3063;
assign w15859 = ~w3079 & ~w3078;
assign w15860 = w3537 & ~w3533;
assign w15861 = w3461 & ~w3514;
assign w15862 = w3493 & ~w3494;
assign w15863 = w3922 & ~w3921;
assign w15864 = w3923 & ~w3919;
assign w15865 = (w3895 & w3889) | (w3895 & w16060) | (w3889 & w16060);
assign w15866 = w3853 & ~w3912;
assign w15867 = w4109 & ~w4194;
assign w15868 = (w15866 & w16622) | (w15866 & w16623) | (w16622 & w16623);
assign w15869 = w4151 & ~w4758;
assign w15870 = ~w4151 & w4758;
assign w15871 = ~w4160 & ~w4159;
assign w15872 = w4990 & ~w4991;
assign w15873 = ~w4843 & w4241;
assign w15874 = ~w4241 & w16512;
assign w15875 = (w4241 & w16513) | (w4241 & w16514) | (w16513 & w16514);
assign w15876 = w4773 & ~w4774;
assign w15877 = (~w4733 & w4734) | (~w4733 & w16066) | (w4734 & w16066);
assign w15878 = w4786 & w5117;
assign w15879 = ~w4786 & ~w5117;
assign w15880 = ~w4820 & ~w4827;
assign w15881 = pi322 & ~w5195;
assign w15882 = ~pi322 & w5195;
assign w15883 = ~w4547 & ~w4518;
assign w15884 = w4614 & w16067;
assign w15885 = ~w5046 & ~w5045;
assign w15886 = ~w5166 & ~w5162;
assign w15887 = ~w5130 & ~w5623;
assign w15888 = w5130 & w5623;
assign w15889 = w5157 & ~w5154;
assign w15890 = ~w5537 & w16069;
assign w15891 = (pi146 & w5537) | (pi146 & w16070) | (w5537 & w16070);
assign w15892 = w5662 & ~w5663;
assign w15893 = (w5580 & w5576) | (w5580 & w16071) | (w5576 & w16071);
assign w15894 = ~w5593 & w6176;
assign w15895 = w5593 & ~w6176;
assign w15896 = ~w5599 & ~w5606;
assign w15897 = w5646 & ~w5652;
assign w15898 = ~w5721 & ~w5719;
assign w15899 = w6302 & ~w6301;
assign w15900 = w5503 & ~w6327;
assign w15901 = ~w5495 & ~w6339;
assign w15902 = w5495 & w6339;
assign w15903 = w5982 & ~w5976;
assign w15904 = w5915 & ~w6408;
assign w15905 = ~w5915 & w6408;
assign w15906 = (~w5845 & ~w5846) | (~w5845 & w16072) | (~w5846 & w16072);
assign w15907 = w5944 & ~w5941;
assign w15908 = w5947 & ~w5842;
assign w15909 = (~w5971 & w5832) | (~w5971 & w16073) | (w5832 & w16073);
assign w15910 = ~w6018 & ~w6017;
assign w15911 = w6067 & ~w2170;
assign w15912 = ~w6348 & ~w6063;
assign w15913 = w6304 & ~w6303;
assign w15914 = (w6296 & ~w6292) | (w6296 & w16075) | (~w6292 & w16075);
assign w15915 = ~w6236 & ~w6242;
assign w15916 = (~w6229 & w6232) | (~w6229 & w17616) | (w6232 & w17616);
assign w15917 = w6170 & ~w6169;
assign w15918 = w6207 & ~w7012;
assign w15919 = ~w6207 & w7012;
assign w15920 = ~w6273 & ~w7088;
assign w15921 = (~w6849 & ~w6050) | (~w6849 & w16076) | (~w6050 & w16076);
assign w15922 = w7482 & ~w7485;
assign w15923 = w6328 & ~w6329;
assign w15924 = ~w3183 & w7492;
assign w15925 = (w7156 & w16077) | (w7156 & w16078) | (w16077 & w16078);
assign w15926 = w7512 & ~w7511;
assign w15927 = ~w7554 & ~w7089;
assign w15928 = w7080 & ~w7077;
assign w15929 = w7059 & w7066;
assign w15930 = w7084 & ~w7096;
assign w15931 = ~pi322 & ~w7550;
assign w15932 = pi322 & w7550;
assign w15933 = ~w7727 & ~w8167;
assign w15934 = w7727 & pi259;
assign w15935 = w8173 & ~w8172;
assign w15936 = ~pi322 & w8162;
assign w15937 = pi322 & ~w8162;
assign w15938 = w8164 & ~w8163;
assign w15939 = w8789 & ~w8788;
assign w15940 = w9549 & w9548;
assign w15941 = ~w8607 & ~w8605;
assign w15942 = ~pi261 & w8794;
assign w15943 = (w8793 & w16515) | (w8793 & w16516) | (w16515 & w16516);
assign w15944 = ~w9750 & w8794;
assign w15945 = ~w9754 & w8794;
assign w15946 = (~w8798 & w8787) | (~w8798 & w16517) | (w8787 & w16517);
assign w15947 = (w10321 & ~w10322) | (w10321 & w16624) | (~w10322 & w16624);
assign w15948 = w10322 & w16625;
assign w15949 = w9727 & w10331;
assign w15950 = ~w9727 & ~w10331;
assign w15951 = ~w9705 & w10337;
assign w15952 = w9705 & ~w10337;
assign w15953 = ~w9680 & w10344;
assign w15954 = w9680 & ~w10344;
assign w15955 = w9639 & ~w9637;
assign w15956 = ~w8670 & w9595;
assign w15957 = ~w9581 & ~w9644;
assign w15958 = ~w9651 & ~w10420;
assign w15959 = w9651 & w10420;
assign w15960 = w10534 & w10296;
assign w15961 = w10544 & pi322;
assign w15962 = (w9802 & ~w9791) | (w9802 & w16079) | (~w9791 & w16079);
assign w15963 = w10285 & ~w10286;
assign w15964 = w9846 & ~w9847;
assign w15965 = ~w9906 & ~w9464;
assign w15966 = w10224 & w10683;
assign w15967 = (w10180 & ~w10176) | (w10180 & w16080) | (~w10176 & w16080);
assign w15968 = ~w9951 & ~w10171;
assign w15969 = ~w10677 & ~w10675;
assign w15970 = ~w10669 & ~w10667;
assign w15971 = ~w10234 & ~w10233;
assign w15972 = ~w10239 & ~w10237;
assign w15973 = ~w10244 & ~w10242;
assign w15974 = w10516 & ~w10513;
assign w15975 = (w11077 & w10499) | (w11077 & w16518) | (w10499 & w16518);
assign w15976 = ~w10499 & w16519;
assign w15977 = ~w10481 & ~w10485;
assign w15978 = w10508 & ~w10319;
assign w15979 = ~w11064 & w11073;
assign w15980 = ~w10249 & ~w10248;
assign w15981 = (w11296 & w11287) | (w11296 & w16081) | (w11287 & w16081);
assign w15982 = ~w10489 & w16082;
assign w15983 = ~w10469 & w16083;
assign w15984 = (~w11095 & w10450) | (~w11095 & w16084) | (w10450 & w16084);
assign w15985 = pi259 & w11294;
assign w15986 = ~w11297 & ~w12110;
assign w15987 = w11297 & pi259;
assign w15988 = ~pi322 & ~w11880;
assign w15989 = pi322 & w11880;
assign w15990 = ~w11336 & ~w11333;
assign w15991 = ~w11058 & ~w12157;
assign w15992 = w11058 & w12157;
assign w15993 = w3979 & w4708;
assign w15994 = ~w12211 & pi334;
assign w15995 = ~w10986 & ~w12246;
assign w15996 = w10986 & w12246;
assign w15997 = w10974 & w12268;
assign w15998 = ~w10974 & ~w12268;
assign w15999 = ~w11501 & ~w11500;
assign w16000 = ~w11718 & w11510;
assign w16001 = ~w12552 & ~w1159;
assign w16002 = ~w11738 & ~w11741;
assign w16003 = w11504 & w12593;
assign w16004 = ~w11504 & ~w12593;
assign w16005 = ~w12281 & ~w12280;
assign w16006 = w11762 & w12619;
assign w16007 = ~w11762 & ~w12619;
assign w16008 = ~w10982 & ~w10981;
assign w16009 = ~w11805 & ~w11820;
assign w16010 = w11805 & w11820;
assign w16011 = w12649 & ~w12671;
assign w16012 = ~w12673 & ~w12674;
assign w16013 = w12114 & ~w12111;
assign w16014 = ~w12038 & ~w12726;
assign w16015 = w12038 & w12726;
assign w16016 = w11961 & ~w11958;
assign w16017 = ~w11914 & ~w12003;
assign w16018 = w12022 & ~w12018;
assign w16019 = w11894 & w12927;
assign w16020 = ~w11894 & ~w12927;
assign w16021 = w11888 & w12934;
assign w16022 = ~w11888 & ~w12934;
assign w16023 = pi322 & w12974;
assign w16024 = ~pi322 & ~w12974;
assign w16025 = ~w12217 & ~w13037;
assign w16026 = w11864 & ~w11863;
assign w16027 = w11845 & ~w13078;
assign w16028 = ~w11792 & ~w13109;
assign w16029 = ~w11793 & ~w13114;
assign w16030 = ~w10974 & ~w11784;
assign w16031 = w13135 & ~w13132;
assign w16032 = ~w12930 & ~w12928;
assign w16033 = ~pi322 & w13554;
assign w16034 = pi322 & ~w13554;
assign w16035 = ~w13006 & ~w13002;
assign w16036 = w13083 & ~w13084;
assign w16037 = w12678 & ~w12677;
assign w16038 = w13677 & ~w13676;
assign w16039 = w13714 & ~w13713;
assign w16040 = ~w13141 & ~w13724;
assign w16041 = w12313 & ~w12587;
assign w16042 = ~w597 & ~pi130;
assign w16043 = ~w12606 & w16085;
assign w16044 = w13219 & w13223;
assign w16045 = w13201 & ~w13202;
assign w16046 = ~w14535 & ~w14534;
assign w16047 = w14056 & ~w14055;
assign w16048 = ~w13198 & ~w13196;
assign w16049 = ~w13760 & ~w13758;
assign w16050 = w14012 & ~w14896;
assign w16051 = ~w14012 & w14896;
assign w16052 = ~w14921 & w14925;
assign w16053 = w867 & ~w845;
assign w16054 = w698 & w479;
assign w16055 = w1964 & w1937;
assign w16056 = pi140 & w458;
assign w16057 = w2681 & w15846;
assign w16058 = ~w2896 & ~w2961;
assign w16059 = w2941 & ~w2903;
assign w16060 = w3494 & w3895;
assign w16061 = ~w4102 & w4101;
assign w16062 = ~w4319 & w16333;
assign w16063 = ~w4681 & w4914;
assign w16064 = pi259 & w5043;
assign w16065 = ~pi259 & ~w5043;
assign w16066 = w4779 & ~w4733;
assign w16067 = w4626 & ~w4620;
assign w16068 = (~w5353 & ~w4570) | (~w5353 & w16520) | (~w4570 & w16520);
assign w16069 = ~w5187 & ~pi146;
assign w16070 = w5187 & pi146;
assign w16071 = ~w5575 & w5580;
assign w16072 = ~w5934 & ~w5845;
assign w16073 = ~w5831 & ~w5971;
assign w16074 = ~w6020 & w6019;
assign w16075 = ~w6080 & w6296;
assign w16076 = w6057 & ~w6849;
assign w16077 = ~w3568 & w6329;
assign w16078 = ~w3568 & ~w15923;
assign w16079 = ~w9543 & w9802;
assign w16080 = ~w9950 & w10180;
assign w16081 = w10527 & w16521;
assign w16082 = ~w10333 & ~w11084;
assign w16083 = ~w10339 & ~w11092;
assign w16084 = w10347 & ~w11095;
assign w16085 = w5426 & pi293;
assign w16086 = w477 & pi131;
assign w16087 = w649 & ~w655;
assign w16088 = w651 & w479;
assign w16089 = ~w703 & pi320;
assign w16090 = ~w926 & ~w752;
assign w16091 = ~w928 & ~w915;
assign w16092 = w897 & w772;
assign w16093 = ~w914 & ~w920;
assign w16094 = ~w744 & pi258;
assign w16095 = w1068 & pi133;
assign w16096 = (~w1096 & w1082) | (~w1096 & w16334) | (w1082 & w16334);
assign w16097 = ~w863 & w16522;
assign w16098 = w896 & pi259;
assign w16099 = ~w1298 & ~w1038;
assign w16100 = ~w1298 & w15808;
assign w16101 = ~w1045 & w1304;
assign w16102 = w1045 & ~w1304;
assign w16103 = ~w1311 & w1310;
assign w16104 = w1311 & ~w1310;
assign w16105 = w1058 & w1314;
assign w16106 = ~w1058 & ~w1314;
assign w16107 = ~w1297 & ~w1524;
assign w16108 = (~w1297 & ~w1524) | (~w1297 & w16335) | (~w1524 & w16335);
assign w16109 = (pi130 & w1045) | (pi130 & w16523) | (w1045 & w16523);
assign w16110 = w1557 & ~w1523;
assign w16111 = ~w1511 & ~w1773;
assign w16112 = w1511 & pi259;
assign w16113 = ~w1515 & ~w1514;
assign w16114 = w1571 & ~w1570;
assign w16115 = ~w1789 & w1303;
assign w16116 = ~w1789 & ~w15815;
assign w16117 = w1548 & ~w1303;
assign w16118 = w1548 & w15815;
assign w16119 = ~w1814 & ~w1817;
assign w16120 = w1824 & ~w1783;
assign w16121 = ~w1821 & w1565;
assign w16122 = ~w1821 & w1781;
assign w16123 = w2120 & ~w2119;
assign w16124 = w2343 & ~w2348;
assign w16125 = w2659 & ~w2660;
assign w16126 = w2654 & ~w2651;
assign w16127 = w3054 & w3109;
assign w16128 = ~w3054 & ~w3109;
assign w16129 = ~w3509 & ~w3508;
assign w16130 = w4779 & ~w4174;
assign w16131 = w4779 & ~w4175;
assign w16132 = w4702 & ~w3975;
assign w16133 = pi322 & w4709;
assign w16134 = ~pi322 & ~w4709;
assign w16135 = ~w4876 & w17714;
assign w16136 = (~w4876 & ~w4270) | (~w4876 & w16336) | (~w4270 & w16336);
assign w16137 = (w4270 & w16337) | (w4270 & w16338) | (w16337 & w16338);
assign w16138 = w4270 & w16524;
assign w16139 = ~w4091 & ~w4090;
assign w16140 = ~w4325 & ~w4324;
assign w16141 = w4938 & ~w4939;
assign w16142 = w4979 & w4933;
assign w16143 = (w4979 & w4934) | (w4979 & w16142) | (w4934 & w16142);
assign w16144 = ~w4979 & ~w4933;
assign w16145 = ~w4934 & w16144;
assign w16146 = (w4923 & w16525) | (w4923 & w16526) | (w16525 & w16526);
assign w16147 = w4923 & w16339;
assign w16148 = ~w4983 & w17715;
assign w16149 = (~w4983 & ~w4923) | (~w4983 & w16340) | (~w4923 & w16340);
assign w16150 = w4988 & ~w4991;
assign w16151 = w4988 & w15872;
assign w16152 = ~w4995 & w17716;
assign w16153 = (~w4995 & ~w4910) | (~w4995 & w16341) | (~w4910 & w16341);
assign w16154 = (w4910 & w16342) | (w4910 & w16343) | (w16342 & w16343);
assign w16155 = w4910 & w16527;
assign w16156 = ~w4685 & ~w4999;
assign w16157 = w4685 & w4999;
assign w16158 = ~w4904 & ~w4689;
assign w16159 = ~w4901 & ~w4898;
assign w16160 = w3866 & ~w4126;
assign w16161 = ~w4749 & ~w4748;
assign w16162 = ~w4767 & w5092;
assign w16163 = w4767 & ~w5092;
assign w16164 = w4787 & ~w4786;
assign w16165 = w4589 & w5287;
assign w16166 = ~w4589 & ~w5287;
assign w16167 = ~w4576 & ~w4574;
assign w16168 = ~w4519 & ~w4543;
assign w16169 = w4634 & ~w4631;
assign w16170 = w4499 & ~w4641;
assign w16171 = w5042 & w5034;
assign w16172 = w5085 & w5575;
assign w16173 = ~w5085 & ~w5575;
assign w16174 = ~w5099 & w5055;
assign w16175 = w5107 & ~w5599;
assign w16176 = ~w5394 & ~w5391;
assign w16177 = ~w5354 & w5353;
assign w16178 = (~w5354 & ~w5359) | (~w5354 & w16528) | (~w5359 & w16528);
assign w16179 = ~w5773 & ~w5772;
assign w16180 = ~w5751 & ~w5749;
assign w16181 = ~w5509 & ~w5507;
assign w16182 = ~w5536 & ~w5705;
assign w16183 = w5538 & w6099;
assign w16184 = ~w6105 & ~w6100;
assign w16185 = w6101 & w6108;
assign w16186 = pi260 & ~w5538;
assign w16187 = w6266 & ~w6258;
assign w16188 = w6184 & ~w6183;
assign w16189 = ~w7090 & w7092;
assign w16190 = ~w7094 & ~w7099;
assign w16191 = w7094 & w7099;
assign w16192 = ~pi322 & ~w6908;
assign w16193 = pi322 & w6908;
assign w16194 = w8177 & ~w8171;
assign w16195 = w7525 & ~w8390;
assign w16196 = ~w7783 & ~w7781;
assign w16197 = ~w8132 & ~w8114;
assign w16198 = w8598 & w8163;
assign w16199 = w8598 & ~w15938;
assign w16200 = ~w8170 & ~w8169;
assign w16201 = ~w8161 & ~w7743;
assign w16202 = ~w8587 & ~w8585;
assign w16203 = ~w8157 & w8414;
assign w16204 = ~w8895 & ~w8898;
assign w16205 = ~w8564 & ~w8563;
assign w16206 = ~w8854 & ~w9535;
assign w16207 = w9549 & w9561;
assign w16208 = w8808 & w9775;
assign w16209 = ~w8808 & ~w9775;
assign w16210 = pi322 & ~w9785;
assign w16211 = ~pi322 & w9785;
assign w16212 = w8834 & ~w8596;
assign w16213 = ~w8596 & ~w9818;
assign w16214 = ~w8577 & ~w8575;
assign w16215 = w8808 & pi259;
assign w16216 = ~w8808 & ~w9772;
assign w16217 = ~w9771 & w10304;
assign w16218 = w9771 & ~pi154;
assign w16219 = w9761 & ~w10316;
assign w16220 = ~w9761 & w10316;
assign w16221 = ~w9748 & ~w9750;
assign w16222 = w9629 & pi133;
assign w16223 = ~w15956 & ~w10372;
assign w16224 = ~w9625 & ~w9623;
assign w16225 = ~w10406 & ~w10409;
assign w16226 = ~w10299 & ~w10297;
assign w16227 = w10541 & ~w10549;
assign w16228 = w10555 & ~w15962;
assign w16229 = w10555 & w9792;
assign w16230 = ~w9846 & ~pi330;
assign w16231 = ~w9528 & ~w9524;
assign w16232 = w10139 & ~w1420;
assign w16233 = w10139 & w1420;
assign w16234 = ~w10107 & ~w10105;
assign w16235 = w10217 & w10973;
assign w16236 = ~w10217 & ~w10973;
assign w16237 = w10988 & w10667;
assign w16238 = w10988 & ~w15970;
assign w16239 = w10992 & w10233;
assign w16240 = w10992 & ~w15971;
assign w16241 = w10997 & w10237;
assign w16242 = w10997 & ~w15972;
assign w16243 = ~w1865 & w10242;
assign w16244 = ~w1865 & ~w15973;
assign w16245 = ~w10261 & ~w11013;
assign w16246 = ~w10261 & ~w11014;
assign w16247 = w10583 & ~w10582;
assign w16248 = ~w10414 & w11168;
assign w16249 = w10414 & ~w11168;
assign w16250 = (~w10353 & ~w10429) | (~w10353 & w16344) | (~w10429 & w16344);
assign w16251 = ~w11270 & ~w10319;
assign w16252 = ~w11270 & ~w10320;
assign w16253 = w11270 & w10319;
assign w16254 = w11270 & w10320;
assign w16255 = (w11323 & w11070) | (w11323 & w16529) | (w11070 & w16529);
assign w16256 = ~w10296 & ~w11072;
assign w16257 = w10550 & ~w10557;
assign w16258 = ~w10277 & ~w11364;
assign w16259 = w10277 & w11364;
assign w16260 = ~w9883 & ~w9880;
assign w16261 = ~w11433 & ~w11432;
assign w16262 = ~w10705 & ~w11498;
assign w16263 = w10705 & ~pi129;
assign w16264 = ~w10709 & ~w10706;
assign w16265 = (w10943 & ~w10934) | (w10943 & w16530) | (~w10934 & w16530);
assign w16266 = ~w10712 & ~w10929;
assign w16267 = w10914 & ~w11707;
assign w16268 = w10914 & w11709;
assign w16269 = w10914 & w1159;
assign w16270 = ~w10914 & w11707;
assign w16271 = ~w10920 & ~w10923;
assign w16272 = (~w10710 & ~w10946) | (~w10710 & w16531) | (~w10946 & w16531);
assign w16273 = ~w10972 & ~w10971;
assign w16274 = w615 & w10983;
assign w16275 = w10977 & ~w11768;
assign w16276 = ~w615 & w793;
assign w16277 = ~w10977 & w11768;
assign w16278 = w615 & w11775;
assign w16279 = w11435 & ~w11806;
assign w16280 = ~w11435 & ~w11826;
assign w16281 = w11435 & w11826;
assign w16282 = w11411 & w3568;
assign w16283 = w11861 & ~w11860;
assign w16284 = ~w11283 & ~w11280;
assign w16285 = w11261 & ~w11258;
assign w16286 = w11201 & ~w11198;
assign w16287 = w11186 & ~w11184;
assign w16288 = (~w11097 & w11191) | (~w11097 & w16345) | (w11191 & w16345);
assign w16289 = ~w11090 & ~w11234;
assign w16290 = ~w11089 & ~w11088;
assign w16291 = w11082 & ~w11249;
assign w16292 = ~w11327 & ~w11336;
assign w16293 = w15990 | ~w11333;
assign w16294 = (~w11333 & w15990) | (~w11333 & ~w11327) | (w15990 & ~w11327);
assign w16295 = ~w11060 & w15991;
assign w16296 = w15992 & w12157;
assign w16297 = (w12157 & w15992) | (w12157 & w11060) | (w15992 & w11060);
assign w16298 = ~w11010 & ~w11009;
assign w16299 = ~w10976 & ~w10974;
assign w16300 = ~w10968 & ~w12278;
assign w16301 = w10968 & w466;
assign w16302 = w12268 & ~w11765;
assign w16303 = w12625 & ~w12623;
assign w16304 = ~w15989 & w12144;
assign w16305 = w12163 & ~w12164;
assign w16306 = (w11870 & ~w12171) | (w11870 & w16346) | (~w12171 & w16346);
assign w16307 = w12248 & ~w12247;
assign w16308 = ~w12613 & ~w13200;
assign w16309 = w12613 & w466;
assign w16310 = w13164 & ~w13165;
assign w16311 = ~w12618 & ~w12617;
assign w16312 = ~w12622 & ~w12620;
assign w16313 = ~w3183 & w12663;
assign w16314 = w13045 & ~w13267;
assign w16315 = ~w13051 & ~w13280;
assign w16316 = ~w13508 & ~w12926;
assign w16317 = w12612 & ~w13183;
assign w16318 = w14006 & ~w698;
assign w16319 = ~w14015 & w14010;
assign w16320 = w13205 & w13207;
assign w16321 = w14046 & ~w14047;
assign w16322 = w13682 & ~w13683;
assign w16323 = ~w13243 & ~w14471;
assign w16324 = ~w14539 & w14534;
assign w16325 = ~w14539 & ~w16046;
assign w16326 = w13226 & ~w13227;
assign w16327 = w13698 & ~w13691;
assign w16328 = w13731 & ~w13730;
assign w16329 = w14645 & ~w14646;
assign w16330 = (~w1285 & ~w1085) | (~w1285 & w16532) | (~w1085 & w16532);
assign w16331 = w3220 & ~w955;
assign w16332 = w3220 & w15849;
assign w16333 = ~w4070 & ~w4660;
assign w16334 = w1091 & ~w1096;
assign w16335 = ~w1039 & ~w1297;
assign w16336 = ~w4102 & ~w4876;
assign w16337 = w4876 & ~w4101;
assign w16338 = w4876 & ~w16061;
assign w16339 = ~w4661 & w4983;
assign w16340 = w4661 & ~w4983;
assign w16341 = ~w4681 & ~w4995;
assign w16342 = w4995 & ~w4914;
assign w16343 = w4995 & ~w16063;
assign w16344 = w10427 & ~w10353;
assign w16345 = ~w11189 & ~w11097;
assign w16346 = w11872 & w11870;
assign w16347 = ~w945 & w1088;
assign w16348 = w1545 & ~w1301;
assign w16349 = w1545 & w15814;
assign w16350 = ~pi263 & ~w1301;
assign w16351 = ~pi263 & w15814;
assign w16352 = ~w1544 & ~w1554;
assign w16353 = ~w1590 & w16533;
assign w16354 = w1530 & ~w16108;
assign w16355 = w1530 & ~w16107;
assign w16356 = ~w1788 & w1802;
assign w16357 = w1788 & ~w1802;
assign w16358 = ~w15829 & ~w1791;
assign w16359 = ~w2090 & w1799;
assign w16360 = ~w2090 & ~w15828;
assign w16361 = ~w1808 & ~w1807;
assign w16362 = ~w2067 & w2115;
assign w16363 = w2067 & ~w2115;
assign w16364 = w1778 & ~w1828;
assign w16365 = w2144 & w1773;
assign w16366 = w2144 & ~w16111;
assign w16367 = w16112 & w2144;
assign w16368 = w2060 & w2269;
assign w16369 = ~w2060 & ~w2269;
assign w16370 = (w1799 & w2286) | (w1799 & w16534) | (w2286 & w16534);
assign w16371 = ~w2288 & ~w15828;
assign w16372 = ~w2340 & w2335;
assign w16373 = w2340 & ~w2335;
assign w16374 = w2135 & w2343;
assign w16375 = ~w2135 & ~w2343;
assign w16376 = ~w2311 & ~w2310;
assign w16377 = ~pi259 & ~w2366;
assign w16378 = w2677 & pi139;
assign w16379 = ~w2647 & ~w2641;
assign w16380 = w2629 & ~w2630;
assign w16381 = (w2586 & w2577) | (w2586 & w16535) | (w2577 & w16535);
assign w16382 = ~w3131 & ~w3127;
assign w16383 = w3053 & ~w3107;
assign w16384 = ~w3091 & w3095;
assign w16385 = w3564 & ~w3562;
assign w16386 = w3458 & w3522;
assign w16387 = ~w3959 & ~w3955;
assign w16388 = ~w3938 & ~w3943;
assign w16389 = w3930 & ~w3927;
assign w16390 = w4105 & ~w4223;
assign w16391 = w4105 & w4223;
assign w16392 = w4200 & ~w4201;
assign w16393 = ~w4241 & w17617;
assign w16394 = (w5043 & w15874) | (w5043 & ~w4711) | (w15874 & ~w4711);
assign w16395 = w4711 & w15875;
assign w16396 = ~w4815 & ~w4813;
assign w16397 = w5646 & w5154;
assign w16398 = w5646 & w5155;
assign w16399 = ~w5646 & ~w5154;
assign w16400 = ~w5646 & ~w5155;
assign w16401 = (~w6112 & ~w5661) | (~w6112 & w16536) | (~w5661 & w16536);
assign w16402 = ~w5665 & w16537;
assign w16403 = w5661 & w16538;
assign w16404 = (w6112 & w5665) | (w6112 & w16539) | (w5665 & w16539);
assign w16405 = (w5182 & w16626) | (w5182 & w16627) | (w16626 & w16627);
assign w16406 = ~w5020 & w5524;
assign w16407 = w5020 & ~w5524;
assign w16408 = w6300 & w6301;
assign w16409 = w6300 & ~w15899;
assign w16410 = pi330 & w17717;
assign w16411 = w6326 & ~w15900;
assign w16412 = ~w5496 & w15901;
assign w16413 = w15902 & w6339;
assign w16414 = (w6339 & w15902) | (w6339 & w5496) | (w15902 & w5496);
assign w16415 = ~w5953 & ~w5952;
assign w16416 = w5331 & w5892;
assign w16417 = ~w5331 & ~w5892;
assign w16418 = w6414 & ~w4539;
assign w16419 = w6458 & w6464;
assign w16420 = w5965 & ~w6551;
assign w16421 = ~w5965 & w6551;
assign w16422 = w6557 & ~w15909;
assign w16423 = w6557 & w5834;
assign w16424 = w6573 & ~w6570;
assign w16425 = w6546 & ~w6615;
assign w16426 = ~w6546 & w6615;
assign w16427 = w6518 & ~w6621;
assign w16428 = ~w6518 & w6621;
assign w16429 = (w6405 & ~w6525) | (w6405 & w16540) | (~w6525 & w16540);
assign w16430 = w6534 & ~w6729;
assign w16431 = (w6395 & w6576) | (w6395 & w16541) | (w6576 & w16541);
assign w16432 = ~w6825 & ~w6017;
assign w16433 = ~w6825 & w15910;
assign w16434 = ~w6829 & w17718;
assign w16435 = ~w6829 & w6368;
assign w16436 = w6028 & ~w6840;
assign w16437 = ~w6135 & ~w6136;
assign w16438 = ~w6124 & ~w6177;
assign w16439 = ~w7036 & ~w6229;
assign w16440 = ~w7036 & ~w6231;
assign w16441 = w7036 & w6229;
assign w16442 = w7036 & w6231;
assign w16443 = w7182 & w7181;
assign w16444 = ~w7182 & ~w7181;
assign w16445 = ~w7190 & ~w7188;
assign w16446 = ~w6864 & ~w6863;
assign w16447 = w2373 & w7480;
assign w16448 = w7492 & w7497;
assign w16449 = w7498 & pi330;
assign w16450 = w6984 & ~w6982;
assign w16451 = (w6931 & ~w6974) | (w6931 & w16542) | (~w6974 & w16542);
assign w16452 = ~w6987 & ~w6993;
assign w16453 = w7675 & w7674;
assign w16454 = ~w7675 & ~w7674;
assign w16455 = ~w6859 & ~w6858;
assign w16456 = w7477 & w8115;
assign w16457 = ~w7477 & ~w8115;
assign w16458 = ~w8439 & ~w8438;
assign w16459 = ~w8310 & w8316;
assign w16460 = ~w8890 & ~w9507;
assign w16461 = ~w9817 & ~w9828;
assign w16462 = w9817 & w9828;
assign w16463 = w9849 & ~w8575;
assign w16464 = w9849 & w16214;
assign w16465 = w9503 & ~w9495;
assign w16466 = w10253 & w10252;
assign w16467 = ~w10253 & ~w10252;
assign w16468 = ~w9512 & ~w9510;
assign w16469 = ~w9517 & ~w9515;
assign w16470 = w9529 & ~w9838;
assign w16471 = w8847 & w9824;
assign w16472 = ~w8847 & ~w9824;
assign w16473 = ~w16218 & w10309;
assign w16474 = w8670 & ~w9595;
assign w16475 = ~w9665 & w9670;
assign w16476 = ~w9734 & ~w9739;
assign w16477 = w10581 & ~w10286;
assign w16478 = w10581 & w15963;
assign w16479 = w10723 & ~w10719;
assign w16480 = ~w9959 & ~w10112;
assign w16481 = ~w2473 & ~w10868;
assign w16482 = w10875 & w2801;
assign w16483 = ~w10148 & ~w10146;
assign w16484 = w10163 & w10914;
assign w16485 = ~w10163 & ~w10914;
assign w16486 = ~w10496 & ~w10492;
assign w16487 = w10482 & ~w11085;
assign w16488 = ~w10482 & w11085;
assign w16489 = w10410 & ~w11164;
assign w16490 = w10488 & ~w10333;
assign w16491 = pi259 & w10303;
assign w16492 = w10304 & ~w11303;
assign w16493 = ~w10304 & w11303;
assign w16494 = w10579 & ~w10578;
assign w16495 = w10644 & w9880;
assign w16496 = w10644 & ~w16260;
assign w16497 = ~w11094 & w11216;
assign w16498 = w11726 & pi298;
assign w16499 = ~w12112 & ~w12706;
assign w16500 = w12112 & w12706;
assign w16501 = ~w12087 & ~w12091;
assign w16502 = ~w11895 & w16020;
assign w16503 = w12987 & ~w12164;
assign w16504 = w12987 & w16305;
assign w16505 = ~w13000 & ~w16306;
assign w16506 = ~w13000 & w12172;
assign w16507 = w14095 & w14047;
assign w16508 = w14095 & ~w16321;
assign w16509 = w14677 & w13758;
assign w16510 = w14677 & ~w16049;
assign w16511 = w2125 & ~w2333;
assign w16512 = w4231 & w16064;
assign w16513 = w16065 | ~w5043;
assign w16514 = (~w5043 & w16065) | (~w5043 & ~w4231) | (w16065 & ~w4231);
assign w16515 = w9750 & w8788;
assign w16516 = w9750 & ~w15939;
assign w16517 = w8794 & ~w8798;
assign w16518 = pi148 & w17719;
assign w16519 = ~w10329 & ~w11077;
assign w16520 = w4513 & ~w5353;
assign w16521 = pi153 & w599;
assign w16522 = w16054 & w855;
assign w16523 = ~w1301 & pi130;
assign w16524 = pi326 & w17720;
assign w16525 = pi336 & w17721;
assign w16526 = w4983 & ~w16062;
assign w16527 = pi333 & w3819;
assign w16528 = ~w16068 & ~w5354;
assign w16529 = ~pi323 & w11323;
assign w16530 = ~w10711 & w10943;
assign w16531 = w10951 & ~w10710;
assign w16532 = ~w16098 & ~w1285;
assign w16533 = ~w1507 & ~w1594;
assign w16534 = w2079 & w1799;
assign w16535 = w2270 & w2586;
assign w16536 = w5544 & ~w6112;
assign w16537 = (~w6112 & w5169) | (~w6112 & w17618) | (w5169 & w17618);
assign w16538 = ~w5544 & w6112;
assign w16539 = ~w5169 & w17619;
assign w16540 = ~w6524 & w6405;
assign w16541 = ~w6577 & w6395;
assign w16542 = w6973 & w6931;
assign w16543 = ~w15798 & pi321;
assign w16544 = ~w658 & ~w650;
assign w16545 = ~w683 & ~w720;
assign w16546 = ~w857 & w710;
assign w16547 = w1509 & w1082;
assign w16548 = ~w1508 & ~w1082;
assign w16549 = ~w1529 & ~w1796;
assign w16550 = w1529 & w1796;
assign w16551 = ~pi322 & ~w1771;
assign w16552 = pi322 & w1771;
assign w16553 = w15830 & ~w1795;
assign w16554 = (~w1795 & w15830) | (~w1795 & ~w1529) | (w15830 & ~w1529);
assign w16555 = w2095 & ~w1799;
assign w16556 = w2095 & w15828;
assign w16557 = w15829 & w2100;
assign w16558 = w2287 & w2305;
assign w16559 = ~w2287 & ~w2305;
assign w16560 = ~w2287 & ~w2298;
assign w16561 = ~w15840 & ~w2632;
assign w16562 = w3112 & ~w2651;
assign w16563 = w3112 & ~w3048;
assign w16564 = ~w3112 & w2651;
assign w16565 = ~w3112 & w3048;
assign w16566 = ~pi259 & ~w2363;
assign w16567 = ~w3167 & ~w3451;
assign w16568 = w3167 & pi259;
assign w16569 = ~w3459 & w3518;
assign w16570 = w3459 & ~w3518;
assign w16571 = w3563 & pi322;
assign w16572 = w3563 & pi323;
assign w16573 = ~w3450 & ~w3844;
assign w16574 = w3450 & pi259;
assign w16575 = ~w3501 & ~w3500;
assign w16576 = w3963 & w3453;
assign w16577 = (w3963 & w3454) | (w3963 & w16576) | (w3454 & w16576);
assign w16578 = ~w3963 & ~w3453;
assign w16579 = ~w3454 & w16578;
assign w16580 = ~w3907 & ~w3906;
assign w16581 = ~w4179 & ~w3920;
assign w16582 = ~w3843 & ~w4232;
assign w16583 = w3843 & pi259;
assign w16584 = w4246 & pi322;
assign w16585 = ~w4231 & ~w4710;
assign w16586 = w4231 & pi259;
assign w16587 = ~w4227 & ~w4234;
assign w16588 = ~w4174 & ~w4175;
assign w16589 = w5114 & ~w5115;
assign w16590 = w5108 & ~w5107;
assign w16591 = pi146 & ~w5705;
assign w16592 = ~pi146 & w5705;
assign w16593 = ~w15881 & ~w5199;
assign w16594 = w5481 & ~w5784;
assign w16595 = ~w5480 & ~w5479;
assign w16596 = ~w5486 & ~w5485;
assign w16597 = ~w5491 & ~w5489;
assign w16598 = ~w6066 & ~w5772;
assign w16599 = ~w6066 & w16179;
assign w16600 = w6071 & w5749;
assign w16601 = w6071 & ~w16180;
assign w16602 = w6075 & w5507;
assign w16603 = w6075 & ~w16181;
assign w16604 = ~w5538 & ~w6103;
assign w16605 = ~w6237 & w6236;
assign w16606 = w6237 & ~w6236;
assign w16607 = ~w6874 & ~w6065;
assign w16608 = ~w6078 & ~w6076;
assign w16609 = ~w7488 & w7485;
assign w16610 = ~w7488 & w7161;
assign w16611 = w7056 & ~w7051;
assign w16612 = w7691 & ~w7690;
assign w16613 = ~w10984 & ~w10675;
assign w16614 = ~w10984 & w15969;
assign w16615 = w10984 & w10675;
assign w16616 = w10984 & ~w15969;
assign w16617 = ~w10987 & w15995;
assign w16618 = w15996 & w12246;
assign w16619 = (w12246 & w15996) | (w12246 & w10987) | (w15996 & w10987);
assign w16620 = w2322 & w2636;
assign w16621 = ~w2322 & ~w2636;
assign w16622 = ~w4174 & ~w3912;
assign w16623 = ~w4174 & ~w3914;
assign w16624 = w9748 & w10321;
assign w16625 = ~w9748 & ~w10321;
assign w16626 = ~w5674 & w5045;
assign w16627 = (~w5674 & w5046) | (~w5674 & w16626) | (w5046 & w16626);
assign w16628 = w14 & ~w13;
assign w16629 = ~w12 & w9;
assign w16630 = ~w6 & w29;
assign w16631 = w3 & w33;
assign w16632 = ~w108 & w109;
assign w16633 = ~w111 & w112;
assign w16634 = ~w115 & w116;
assign w16635 = w117 & ~w116;
assign w16636 = w117 & ~w16634;
assign w16637 = w118 & ~w16635;
assign w16638 = w118 & ~w16636;
assign w16639 = ~w124 & ~w82;
assign w16640 = ~w132 & ~w2;
assign w16641 = ~w136 & pi162;
assign w16642 = w136 & pi258;
assign w16643 = ~w136 & pi163;
assign w16644 = pi259 & w136;
assign w16645 = ~w136 & pi164;
assign w16646 = w136 & pi268;
assign w16647 = ~w136 & pi165;
assign w16648 = w136 & pi269;
assign w16649 = ~w136 & pi166;
assign w16650 = w136 & pi270;
assign w16651 = ~w136 & pi167;
assign w16652 = w136 & pi271;
assign w16653 = ~w136 & pi168;
assign w16654 = w136 & pi272;
assign w16655 = ~w136 & pi169;
assign w16656 = w136 & pi273;
assign w16657 = ~w136 & pi170;
assign w16658 = w136 & pi274;
assign w16659 = ~w136 & pi171;
assign w16660 = w136 & pi275;
assign w16661 = ~w136 & pi172;
assign w16662 = w136 & pi276;
assign w16663 = ~w136 & pi173;
assign w16664 = w136 & pi277;
assign w16665 = w136 & pi260;
assign w16666 = ~w136 & pi174;
assign w16667 = ~w136 & pi175;
assign w16668 = w136 & pi278;
assign w16669 = ~w136 & pi176;
assign w16670 = pi279 & w136;
assign w16671 = ~w136 & pi177;
assign w16672 = w136 & pi280;
assign w16673 = ~w136 & pi178;
assign w16674 = pi281 & w136;
assign w16675 = ~w136 & pi179;
assign w16676 = pi282 & w136;
assign w16677 = ~w136 & pi180;
assign w16678 = w136 & pi283;
assign w16679 = ~w136 & pi181;
assign w16680 = w136 & pi284;
assign w16681 = ~w136 & pi182;
assign w16682 = pi285 & w136;
assign w16683 = ~w136 & pi183;
assign w16684 = pi286 & w136;
assign w16685 = ~w136 & pi184;
assign w16686 = pi287 & w136;
assign w16687 = ~w136 & pi185;
assign w16688 = w136 & pi261;
assign w16689 = ~w136 & pi186;
assign w16690 = w136 & pi288;
assign w16691 = ~w136 & ~pi187;
assign w16692 = w136 & ~pi289;
assign w16693 = ~w136 & pi188;
assign w16694 = w136 & pi262;
assign w16695 = ~w136 & pi189;
assign w16696 = w136 & pi263;
assign w16697 = ~w136 & pi190;
assign w16698 = w136 & pi264;
assign w16699 = ~w136 & pi191;
assign w16700 = w136 & pi265;
assign w16701 = ~w136 & pi192;
assign w16702 = w136 & pi266;
assign w16703 = ~w136 & pi193;
assign w16704 = w136 & pi267;
assign w16705 = ~w136 & pi194;
assign w16706 = w136 & pi322;
assign w16707 = ~w136 & pi195;
assign w16708 = pi323 & w136;
assign w16709 = ~w136 & pi196;
assign w16710 = w136 & pi332;
assign w16711 = ~w136 & pi197;
assign w16712 = w136 & pi333;
assign w16713 = ~w136 & pi198;
assign w16714 = w136 & pi334;
assign w16715 = ~w136 & pi199;
assign w16716 = w136 & pi335;
assign w16717 = ~w136 & pi200;
assign w16718 = w136 & pi336;
assign w16719 = ~w136 & pi201;
assign w16720 = w136 & pi337;
assign w16721 = ~w136 & pi202;
assign w16722 = w136 & pi338;
assign w16723 = ~w136 & pi203;
assign w16724 = w136 & pi339;
assign w16725 = ~w136 & pi204;
assign w16726 = w136 & pi340;
assign w16727 = ~w136 & pi205;
assign w16728 = w136 & pi341;
assign w16729 = ~w136 & pi206;
assign w16730 = pi324 & w136;
assign w16731 = ~w136 & pi207;
assign w16732 = w136 & pi342;
assign w16733 = ~w136 & pi208;
assign w16734 = w136 & pi343;
assign w16735 = ~w136 & pi209;
assign w16736 = w136 & pi344;
assign w16737 = ~w136 & pi210;
assign w16738 = w136 & pi345;
assign w16739 = ~w136 & pi211;
assign w16740 = w136 & pi346;
assign w16741 = ~w136 & pi212;
assign w16742 = w136 & pi347;
assign w16743 = ~w136 & pi213;
assign w16744 = w136 & pi348;
assign w16745 = ~w136 & pi214;
assign w16746 = w136 & pi349;
assign w16747 = ~w136 & pi215;
assign w16748 = w136 & pi350;
assign w16749 = ~w136 & pi216;
assign w16750 = w136 & pi351;
assign w16751 = ~w136 & pi217;
assign w16752 = pi325 & w136;
assign w16753 = ~w136 & pi218;
assign w16754 = ~w132 & pi352;
assign w16755 = ~w136 & pi219;
assign w16756 = w136 & pi353;
assign w16757 = ~w136 & pi220;
assign w16758 = w136 & pi326;
assign w16759 = ~w136 & pi221;
assign w16760 = pi327 & w136;
assign w16761 = ~w136 & pi222;
assign w16762 = w136 & pi328;
assign w16763 = ~w136 & pi223;
assign w16764 = pi329 & w136;
assign w16765 = ~w136 & pi224;
assign w16766 = pi330 & w136;
assign w16767 = ~w136 & pi225;
assign w16768 = w136 & pi331;
assign w16769 = ~w136 & pi226;
assign w16770 = w136 & pi321;
assign w16771 = ~w136 & pi227;
assign w16772 = pi320 & w136;
assign w16773 = ~w136 & pi228;
assign w16774 = w136 & pi311;
assign w16775 = ~w136 & pi229;
assign w16776 = w136 & pi310;
assign w16777 = ~w136 & pi230;
assign w16778 = w136 & pi309;
assign w16779 = ~w136 & pi231;
assign w16780 = w136 & pi308;
assign w16781 = ~w136 & pi232;
assign w16782 = w136 & pi307;
assign w16783 = ~w136 & pi233;
assign w16784 = w136 & pi306;
assign w16785 = ~w136 & pi234;
assign w16786 = w136 & pi305;
assign w16787 = ~w136 & pi235;
assign w16788 = w136 & pi304;
assign w16789 = ~w136 & pi236;
assign w16790 = w136 & pi303;
assign w16791 = ~w136 & pi237;
assign w16792 = w136 & pi302;
assign w16793 = ~w136 & pi238;
assign w16794 = pi319 & w136;
assign w16795 = ~w136 & pi239;
assign w16796 = w136 & pi301;
assign w16797 = ~w136 & pi240;
assign w16798 = w136 & pi300;
assign w16799 = ~w136 & pi241;
assign w16800 = w136 & pi299;
assign w16801 = ~w136 & pi242;
assign w16802 = w136 & pi298;
assign w16803 = ~w136 & pi243;
assign w16804 = w136 & pi297;
assign w16805 = ~w136 & pi244;
assign w16806 = w136 & pi296;
assign w16807 = ~w136 & pi245;
assign w16808 = w136 & pi295;
assign w16809 = ~w136 & pi246;
assign w16810 = w136 & pi294;
assign w16811 = ~w136 & pi247;
assign w16812 = w136 & pi293;
assign w16813 = ~w136 & pi248;
assign w16814 = w136 & pi292;
assign w16815 = ~w136 & pi249;
assign w16816 = w136 & pi318;
assign w16817 = ~w136 & pi250;
assign w16818 = w136 & pi291;
assign w16819 = ~w136 & pi251;
assign w16820 = w136 & pi290;
assign w16821 = ~w136 & pi252;
assign w16822 = w136 & pi317;
assign w16823 = ~w136 & pi253;
assign w16824 = w136 & pi316;
assign w16825 = ~w136 & pi254;
assign w16826 = w136 & pi315;
assign w16827 = ~w136 & pi255;
assign w16828 = w136 & pi314;
assign w16829 = ~w136 & pi256;
assign w16830 = w136 & pi313;
assign w16831 = ~w136 & pi257;
assign w16832 = w136 & pi312;
assign w16833 = pi128 & ~w449;
assign w16834 = ~w16833 & pi258;
assign w16835 = ~pi258 & ~w461;
assign w16836 = ~w460 & pi322;
assign w16837 = ~pi321 & ~w477;
assign w16838 = ~pi259 & pi161;
assign w16839 = ~pi128 & pi258;
assign w16840 = ~w535 & ~w456;
assign w16841 = ~pi322 & ~w512;
assign w16842 = ~w460 & pi323;
assign w16843 = w539 & ~w512;
assign w16844 = w539 & w16841;
assign w16845 = ~w535 & ~pi324;
assign w16846 = ~pi324 & w541;
assign w16847 = ~w540 & ~w543;
assign w16848 = w481 & ~w474;
assign w16849 = ~w558 & ~w135;
assign w16850 = w491 & pi161;
assign w16851 = ~pi260 & ~w549;
assign w16852 = ~w460 & pi324;
assign w16853 = w535 & pi323;
assign w16854 = pi322 & w539;
assign w16855 = pi258 & w529;
assign w16856 = w603 & pi128;
assign w16857 = w514 & w604;
assign w16858 = ~pi322 & ~w570;
assign w16859 = ~w535 & pi322;
assign w16860 = w456 & w17722;
assign w16861 = ~w558 & ~w556;
assign w16862 = pi319 & ~w662;
assign w16863 = w670 & ~w135;
assign w16864 = ~pi261 & pi161;
assign w16865 = ~pi128 & ~w728;
assign w16866 = pi129 & w662;
assign w16867 = ~pi129 & ~w731;
assign w16868 = pi131 & pi259;
assign w16869 = pi131 & ~w15799;
assign w16870 = w783 & ~w777;
assign w16871 = ~pi322 & w743;
assign w16872 = pi322 & ~w743;
assign w16873 = ~w568 & ~w626;
assign w16874 = ~w460 & ~w512;
assign w16875 = ~w456 & ~w809;
assign w16876 = w456 & w809;
assign w16877 = pi325 & w809;
assign w16878 = pi325 & ~w16875;
assign w16879 = ~pi261 & ~w635;
assign w16880 = ~w670 & ~w642;
assign w16881 = ~w741 & ~w135;
assign w16882 = ~pi262 & pi161;
assign w16883 = ~w699 & w698;
assign w16884 = pi129 & w682;
assign w16885 = ~pi129 & w876;
assign w16886 = ~pi262 & ~w820;
assign w16887 = ~w460 & pi326;
assign w16888 = ~w805 & ~w803;
assign w16889 = w914 & ~pi130;
assign w16890 = w929 & ~w919;
assign w16891 = w789 & ~w787;
assign w16892 = ~w771 & w16891;
assign w16893 = w798 & ~w957;
assign w16894 = w798 & ~w617;
assign w16895 = ~w456 & ~w466;
assign w16896 = ~w460 & w456;
assign w16897 = w970 & ~w972;
assign w16898 = ~w537 & w972;
assign w16899 = ~w537 & ~w16897;
assign w16900 = ~w537 & pi325;
assign w16901 = w741 & ~w827;
assign w16902 = w890 & ~w135;
assign w16903 = ~pi263 & pi161;
assign w16904 = w535 & pi326;
assign w16905 = pi325 & w16898;
assign w16906 = pi325 & w16899;
assign w16907 = ~w976 & ~w1010;
assign w16908 = w1009 & w1010;
assign w16909 = w1009 & ~w16907;
assign w16910 = w894 & ~w964;
assign w16911 = ~pi262 & pi261;
assign w16912 = ~w462 & w1024;
assign w16913 = w946 & w773;
assign w16914 = ~w946 & ~w773;
assign w16915 = pi322 & ~w958;
assign w16916 = ~pi323 & ~w959;
assign w16917 = pi322 & ~w1105;
assign w16918 = ~pi322 & w1105;
assign w16919 = ~w893 & ~w980;
assign w16920 = ~w460 & ~w742;
assign w16921 = ~w456 & ~w1122;
assign w16922 = w456 & w1122;
assign w16923 = ~pi263 & ~w989;
assign w16924 = ~w995 & ~w890;
assign w16925 = w738 & ~pi129;
assign w16926 = ~w878 & ~w844;
assign w16927 = ~w846 & ~pi134;
assign w16928 = w846 & pi134;
assign w16929 = w1159 & pi321;
assign w16930 = ~w1162 & ~w1152;
assign w16931 = w1162 & w1152;
assign w16932 = ~w1169 & ~w15806;
assign w16933 = ~w1169 & w870;
assign w16934 = ~w462 & pi316;
assign w16935 = ~w1197 & ~w135;
assign w16936 = ~pi264 & pi161;
assign w16937 = ~w1185 & ~w1182;
assign w16938 = ~pi133 & ~w1155;
assign w16939 = ~w1165 & pi320;
assign w16940 = ~w1159 & pi320;
assign w16941 = ~w1171 & w1231;
assign w16942 = w1171 & ~w1231;
assign w16943 = w838 & ~pi129;
assign w16944 = ~w1191 & ~w1251;
assign w16945 = ~w462 & pi315;
assign w16946 = ~w460 & pi328;
assign w16947 = ~w1007 & ~w1270;
assign w16948 = w1007 & w466;
assign w16949 = ~w1013 & ~w1012;
assign w16950 = w1275 & w1012;
assign w16951 = w1275 & ~w16949;
assign w16952 = ~w1097 & ~w1088;
assign w16953 = ~w1097 & ~w16347;
assign w16954 = ~pi323 & ~w1103;
assign w16955 = pi322 & w1342;
assign w16956 = ~pi322 & ~w1342;
assign w16957 = ~w1018 & ~w1016;
assign w16958 = ~w1118 & ~w1116;
assign w16959 = w535 & pi327;
assign w16960 = ~w1364 & ~w466;
assign w16961 = w1366 & w1363;
assign w16962 = ~w1366 & w537;
assign w16963 = ~pi264 & ~w1134;
assign w16964 = w1197 & ~w1142;
assign w16965 = ~w1388 & w1268;
assign w16966 = w1268 & ~w135;
assign w16967 = ~pi265 & pi161;
assign w16968 = ~w1207 & ~w1246;
assign w16969 = ~w846 & ~pi135;
assign w16970 = ~w16969 & ~w1215;
assign w16971 = ~pi133 & w1215;
assign w16972 = ~pi133 & ~w16970;
assign w16973 = ~pi136 & ~pi134;
assign w16974 = w1411 & w1410;
assign w16975 = ~w1408 & ~w1414;
assign w16976 = ~w16969 & w1417;
assign w16977 = ~w1413 & pi321;
assign w16978 = w1165 & pi320;
assign w16979 = ~w1234 & w1428;
assign w16980 = w1234 & ~w1428;
assign w16981 = ~w1238 & w1209;
assign w16982 = ~w1256 & ~w1253;
assign w16983 = w1145 & ~pi129;
assign w16984 = ~w1262 & ~w1460;
assign w16985 = ~w462 & w1466;
assign w16986 = ~pi265 & ~w1382;
assign w16987 = ~w460 & pi329;
assign w16988 = ~w1269 & ~w1477;
assign w16989 = w1269 & w466;
assign w16990 = w535 & pi328;
assign w16991 = ~w1368 & ~w1483;
assign w16992 = ~w1359 & ~w1357;
assign w16993 = ~w1278 & ~w1277;
assign w16994 = w1349 & ~w1347;
assign w16995 = ~w1079 & ~w1282;
assign w16996 = w1079 & pi259;
assign w16997 = w1536 & pi130;
assign w16998 = w1536 & w16109;
assign w16999 = ~w1308 & w1557;
assign w17000 = ~w1082 & ~w1507;
assign w17001 = ~w1082 & ~w1088;
assign w17002 = ~w1082 & ~w16347;
assign w17003 = ~w1082 & pi323;
assign w17004 = ~pi322 & ~w1605;
assign w17005 = pi322 & w1605;
assign w17006 = ~w16955 & ~w1341;
assign w17007 = ~w1368 & ~w1271;
assign w17008 = ~w1474 & ~w135;
assign w17009 = ~pi266 & pi161;
assign w17010 = w1465 & w1467;
assign w17011 = ~w1404 & ~w1445;
assign w17012 = ~pi136 & ~w1676;
assign w17013 = ~pi134 & ~w1675;
assign w17014 = w846 & pi137;
assign w17015 = w1408 & pi137;
assign w17016 = w1408 & w17014;
assign w17017 = ~w1681 & ~w17015;
assign w17018 = ~w1681 & ~w17016;
assign w17019 = ~w846 & w1684;
assign w17020 = ~w17019 & ~w1685;
assign w17021 = ~w846 & w1685;
assign w17022 = ~w17021 & ~w1688;
assign w17023 = ~w1679 & pi321;
assign w17024 = w1220 & w1421;
assign w17025 = ~w1220 & ~w1420;
assign w17026 = ~w1696 & pi320;
assign w17027 = w1695 & w1694;
assign w17028 = ~w1431 & w1702;
assign w17029 = w1431 & ~w1702;
assign w17030 = ~w1435 & w1406;
assign w17031 = ~w1403 & ~w1452;
assign w17032 = w1461 & ~w1457;
assign w17033 = ~w462 & pi313;
assign w17034 = w1481 & ~w1635;
assign w17035 = ~w1489 & ~w1487;
assign w17036 = ~w1495 & ~w1619;
assign w17037 = w1497 & ~w1613;
assign w17038 = w1609 & ~w1607;
assign w17039 = w1492 & ~w1493;
assign w17040 = w535 & pi329;
assign w17041 = ~w1480 & ~w1479;
assign w17042 = ~w1896 & ~w1479;
assign w17043 = ~w1896 & w17041;
assign w17044 = ~w460 & pi330;
assign w17045 = ~w1476 & ~w1903;
assign w17046 = ~pi266 & ~w1647;
assign w17047 = w1474 & ~w1654;
assign w17048 = w1752 & ~w135;
assign w17049 = ~pi267 & pi161;
assign w17050 = ~w1413 & pi319;
assign w17051 = w15821 | w1673;
assign w17052 = (w1673 & w15821) | (w1673 & w1431) | (w15821 & w1431);
assign w17053 = w1680 & pi133;
assign w17054 = ~w1945 & ~w1947;
assign w17055 = ~pi320 & w1693;
assign w17056 = ~w1709 & w1672;
assign w17057 = w1972 & ~w1159;
assign w17058 = w1977 & ~w1670;
assign w17059 = ~w1717 & w1213;
assign w17060 = w1990 & w1936;
assign w17061 = w1997 & ~w1989;
assign w17062 = w1725 & ~w855;
assign w17063 = ~w1666 & ~w1739;
assign w17064 = w1401 & ~pi129;
assign w17065 = ~w1746 & ~w2018;
assign w17066 = ~pi267 & ~w1914;
assign w17067 = ~w460 & pi331;
assign w17068 = ~w1753 & ~w2037;
assign w17069 = w1753 & w466;
assign w17070 = ~w1899 & ~w1897;
assign w17071 = ~w1763 & ~w1762;
assign w17072 = ~w1764 & ~w1876;
assign w17073 = ~w1769 & ~w1770;
assign w17074 = ~w2079 & w1793;
assign w17075 = w1529 & w2084;
assign w17076 = ~pi131 & ~w16360;
assign w17077 = ~pi131 & ~w16359;
assign w17078 = ~w2090 & w2092;
assign w17079 = ~w2097 & ~w1791;
assign w17080 = ~w2097 & w16358;
assign w17081 = w15829 & ~pi265;
assign w17082 = w1589 & w1859;
assign w17083 = ~w2165 & ~w1859;
assign w17084 = ~w2165 & ~w17082;
assign w17085 = ~pi322 & ~w2056;
assign w17086 = pi322 & w2056;
assign w17087 = w1869 & ~w1867;
assign w17088 = ~w1886 & ~w1885;
assign w17089 = ~w1892 & ~w1756;
assign w17090 = w1905 & ~w1904;
assign w17091 = ~w2215 & w1904;
assign w17092 = ~w2215 & ~w17090;
assign w17093 = ~w1920 & ~w1752;
assign w17094 = w2034 & ~w135;
assign w17095 = ~pi268 & pi161;
assign w17096 = w535 & pi331;
assign w17097 = ~w2040 & ~w2039;
assign w17098 = w2250 & w2039;
assign w17099 = w2250 & ~w17097;
assign w17100 = ~w2041 & ~w2205;
assign w17101 = ~w2047 & ~w2046;
assign w17102 = w2257 & w2046;
assign w17103 = w2257 & ~w17101;
assign w17104 = w2049 & ~w2182;
assign w17105 = ~w2057 & ~w2265;
assign w17106 = w2057 & pi259;
assign w17107 = ~w2149 & w2143;
assign w17108 = w2078 & ~w16554;
assign w17109 = w2078 & ~w16553;
assign w17110 = ~w2077 & ~w2295;
assign w17111 = w2077 & w2295;
assign w17112 = pi129 & w2295;
assign w17113 = ~pi129 & ~w2295;
assign w17114 = pi130 & w1799;
assign w17115 = pi130 & ~w15828;
assign w17116 = ~w2090 & ~w2312;
assign w17117 = w2090 & ~w17114;
assign w17118 = w2090 & ~w17115;
assign w17119 = ~pi322 & ~w2264;
assign w17120 = pi322 & w2264;
assign w17121 = w2174 & ~w2172;
assign w17122 = ~w2177 & ~w2054;
assign w17123 = ~w2048 & ~w2188;
assign w17124 = ~w2201 & ~w2200;
assign w17125 = w537 & ~w2214;
assign w17126 = ~w537 & pi330;
assign w17127 = ~pi268 & ~w2226;
assign w17128 = ~w2233 & ~w2034;
assign w17129 = w1932 & ~pi129;
assign w17130 = ~w1932 & ~w2451;
assign w17131 = ~w1750 & ~w2026;
assign w17132 = ~w2014 & ~w2012;
assign w17133 = w1935 & ~w2004;
assign w17134 = ~w1413 & pi318;
assign w17135 = ~w1679 & pi319;
assign w17136 = w1961 & ~w1942;
assign w17137 = ~w1954 & ~w1693;
assign w17138 = ~w1954 & ~w17055;
assign w17139 = pi320 & ~w17138;
assign w17140 = pi320 & ~w17137;
assign w17141 = ~w1950 & ~w2470;
assign w17142 = w1950 & w2470;
assign w17143 = w1693 & w1955;
assign w17144 = ~w1696 & w1954;
assign w17145 = ~w2467 & w2474;
assign w17146 = w1973 & w1979;
assign w17147 = w2495 & ~w2494;
assign w17148 = ~w2495 & w2494;
assign w17149 = w1725 & ~w1936;
assign w17150 = w2019 & w653;
assign w17151 = w709 & pi313;
assign w17152 = w2541 & ~w135;
assign w17153 = ~pi269 & pi161;
assign w17154 = ~pi269 & ~w2438;
assign w17155 = w2245 & w466;
assign w17156 = ~w460 & pi333;
assign w17157 = ~w2245 & ~w2556;
assign w17158 = ~w2253 & ~w2252;
assign w17159 = w2559 & w2252;
assign w17160 = w2559 & ~w17158;
assign w17161 = ~w2261 & ~w2396;
assign w17162 = ~w2262 & ~w2389;
assign w17163 = ~w2385 & ~w2384;
assign w17164 = w2268 & ~w2578;
assign w17165 = ~w16560 & pi130;
assign w17166 = w2595 & ~pi130;
assign w17167 = w2595 & ~w17165;
assign w17168 = ~w2077 & ~w2294;
assign w17169 = ~w2293 & ~w2604;
assign w17170 = w2293 & w2604;
assign w17171 = ~w16560 & w2291;
assign w17172 = pi131 & ~w2610;
assign w17173 = w2287 & w2298;
assign w17174 = ~pi131 & w2610;
assign w17175 = ~w2364 & ~w2687;
assign w17176 = w2364 & w2687;
assign w17177 = w2368 & ~w2369;
assign w17178 = w2377 & ~w2375;
assign w17179 = ~w2260 & ~w2258;
assign w17180 = w2408 & ~w2406;
assign w17181 = ~w2254 & ~w2412;
assign w17182 = ~w2424 & ~w2421;
assign w17183 = ~w793 & w2421;
assign w17184 = ~w793 & ~w17182;
assign w17185 = pi332 & ~w537;
assign w17186 = w2248 & w2752;
assign w17187 = w2248 & ~w2246;
assign w17188 = ~w2541 & ~w2447;
assign w17189 = ~w2508 & ~w2502;
assign w17190 = ~w1413 & pi317;
assign w17191 = ~w1679 & pi318;
assign w17192 = ~w2464 & ~w2490;
assign w17193 = pi139 & ~w2469;
assign w17194 = w2789 & w2469;
assign w17195 = w2789 & ~w17193;
assign w17196 = ~pi140 & pi137;
assign w17197 = ~pi140 & ~pi138;
assign w17198 = pi139 & ~w2789;
assign w17199 = w2465 & ~w2482;
assign w17200 = ~w2463 & ~w2497;
assign w17201 = w2511 & ~w2459;
assign w17202 = w2518 & ~w2515;
assign w17203 = ~w2454 & ~w2530;
assign w17204 = ~w2453 & ~w2450;
assign w17205 = ~pi128 & ~w464;
assign w17206 = ~w2880 & ~w135;
assign w17207 = ~pi270 & pi161;
assign w17208 = ~w2845 & ~w2842;
assign w17209 = ~w2779 & ~w2837;
assign w17210 = ~w1413 & pi316;
assign w17211 = ~w1679 & pi317;
assign w17212 = ~w2783 & ~w2817;
assign w17213 = ~pi140 & ~w2909;
assign w17214 = pi138 & ~w2908;
assign w17215 = ~w2913 & ~w2912;
assign w17216 = ~pi139 & w2908;
assign w17217 = w2915 & ~pi137;
assign w17218 = ~w2788 & pi141;
assign w17219 = pi141 & pi137;
assign w17220 = pi138 & ~w2907;
assign w17221 = ~w2786 & ~w2804;
assign w17222 = ~w2808 & ~w2785;
assign w17223 = w2782 & ~w2823;
assign w17224 = ~w2780 & ~w2830;
assign w17225 = ~w2850 & ~w2777;
assign w17226 = w2860 & ~w2858;
assign w17227 = w2775 & ~w2865;
assign w17228 = w2871 & ~w2872;
assign w17229 = ~w653 & pi310;
assign w17230 = ~w2774 & ~w2999;
assign w17231 = w535 & pi333;
assign w17232 = w2555 & ~w2557;
assign w17233 = w3009 & ~w2557;
assign w17234 = w3009 & w17232;
assign w17235 = w2753 & w3014;
assign w17236 = ~w2753 & ~w3014;
assign w17237 = ~w2562 & ~w2561;
assign w17238 = w2738 & ~w2735;
assign w17239 = w2730 & ~w3024;
assign w17240 = ~w2730 & w3024;
assign w17241 = w2723 & ~w2720;
assign w17242 = ~w2716 & ~w2568;
assign w17243 = ~w2713 & ~w2711;
assign w17244 = ~w2575 & ~w2573;
assign w17245 = ~w17168 & w3059;
assign w17246 = ~w2603 & ~w3059;
assign w17247 = ~w2603 & ~w17245;
assign w17248 = ~w3062 & ~w17246;
assign w17249 = ~w3062 & ~w17247;
assign w17250 = w3066 & w17248;
assign w17251 = w3066 & w17249;
assign w17252 = w3072 & ~w2305;
assign w17253 = w3072 & ~w16558;
assign w17254 = ~w2609 & ~w17253;
assign w17255 = ~w2609 & ~w17252;
assign w17256 = ~w2619 & ~w17166;
assign w17257 = ~w2619 & ~w17167;
assign w17258 = w3085 & ~w3081;
assign w17259 = ~w3079 & ~w3081;
assign w17260 = ~w3079 & w17258;
assign w17261 = w3089 & w2630;
assign w17262 = w3089 & ~w16380;
assign w17263 = w2629 & w3091;
assign w17264 = ~w3101 & w3102;
assign w17265 = ~w3101 & ~w15843;
assign w17266 = w3101 & ~w3102;
assign w17267 = w3101 & w15843;
assign w17268 = ~w2585 & w2266;
assign w17269 = ~w2585 & ~w15844;
assign w17270 = ~w2684 & ~w2679;
assign w17271 = ~w2576 & ~w2701;
assign w17272 = ~pi322 & w3185;
assign w17273 = pi322 & ~w3185;
assign w17274 = ~w2744 & ~w15849;
assign w17275 = w15849 & ~w955;
assign w17276 = (~w955 & w15849) | (~w955 & w2744) | (w15849 & w2744);
assign w17277 = ~w955 & pi330;
assign w17278 = ~w460 & ~pi334;
assign w17279 = ~w2554 & ~w3242;
assign w17280 = w2880 & ~w2771;
assign w17281 = ~w3007 & ~w135;
assign w17282 = ~pi271 & pi161;
assign w17283 = ~w2889 & ~w3270;
assign w17284 = w2889 & ~pi129;
assign w17285 = w2980 & ~w2977;
assign w17286 = ~w1413 & pi315;
assign w17287 = w3280 & ~w15852;
assign w17288 = w3280 & w2899;
assign w17289 = ~w1679 & pi316;
assign w17290 = ~w2909 & ~w2918;
assign w17291 = ~pi138 & w3296;
assign w17292 = ~w2906 & ~w2929;
assign w17293 = w3315 & ~w15855;
assign w17294 = w3315 & w2943;
assign w17295 = ~pi317 & ~w2902;
assign w17296 = ~w2947 & ~w1693;
assign w17297 = w2947 & w1954;
assign w17298 = w3321 & w3323;
assign w17299 = w2902 & ~w1954;
assign w17300 = ~w2964 & ~w2893;
assign w17301 = ~w2967 & ~w2970;
assign w17302 = w2983 & ~w2987;
assign w17303 = ~w3384 & ~pi130;
assign w17304 = w3384 & pi130;
assign w17305 = ~pi271 & ~w3251;
assign w17306 = ~w460 & pi335;
assign w17307 = ~w537 & pi334;
assign w17308 = ~w3013 & ~w3012;
assign w17309 = ~w3410 & ~w3012;
assign w17310 = ~w3410 & w17308;
assign w17311 = ~w3017 & ~w3016;
assign w17312 = ~w3414 & w3016;
assign w17313 = ~w3414 & ~w17311;
assign w17314 = ~w3224 & w3220;
assign w17315 = w3224 & ~w3424;
assign w17316 = pi329 & ~pi330;
assign w17317 = ~w3427 & ~w3426;
assign w17318 = ~w3224 & w3424;
assign w17319 = pi330 & ~pi329;
assign w17320 = ~w3032 & ~w3031;
assign w17321 = w3438 & w3031;
assign w17322 = w3438 & ~w17320;
assign w17323 = w3033 & ~w3202;
assign w17324 = ~w3039 & ~w3037;
assign w17325 = ~w3477 & w3473;
assign w17326 = w3477 & ~w3473;
assign w17327 = ~w3071 & ~w3069;
assign w17328 = w3483 & w3069;
assign w17329 = w3483 & ~w17327;
assign w17330 = ~w3489 & ~w3078;
assign w17331 = ~w3489 & w15859;
assign w17332 = ~w3090 & w3495;
assign w17333 = w3090 & ~w3495;
assign w17334 = ~w3041 & ~w3187;
assign w17335 = w3195 & ~w3193;
assign w17336 = ~w3027 & ~w3026;
assign w17337 = w3019 & ~w3220;
assign w17338 = w3618 & ~w3617;
assign w17339 = w3007 & ~w3258;
assign w17340 = ~w3656 & ~w135;
assign w17341 = ~pi272 & pi161;
assign w17342 = ~w3269 & ~w3666;
assign w17343 = w3269 & ~pi129;
assign w17344 = ~w3273 & ~w3272;
assign w17345 = w3670 & w3272;
assign w17346 = w3670 & ~w17344;
assign w17347 = w3380 & ~w3376;
assign w17348 = ~w3275 & ~w3370;
assign w17349 = w3276 & ~w3364;
assign w17350 = ~w1413 & pi314;
assign w17351 = w3352 & ~w3349;
assign w17352 = ~w1679 & pi315;
assign w17353 = w3345 & ~w3282;
assign w17354 = w3286 & ~w3316;
assign w17355 = ~w3312 & ~w3291;
assign w17356 = ~pi141 & ~w3300;
assign w17357 = ~w3293 & ~w3308;
assign w17358 = ~w2947 & ~w3323;
assign w17359 = ~w17358 & ~w3324;
assign w17360 = ~w3735 & ~w3736;
assign w17361 = w3284 & ~w3340;
assign w17362 = ~w3278 & ~w3357;
assign w17363 = w2998 & w3777;
assign w17364 = ~w460 & pi336;
assign w17365 = ~w3402 & ~w3793;
assign w17366 = w3402 & w466;
assign w17367 = w535 & pi335;
assign w17368 = ~w3403 & ~w3638;
assign w17369 = ~w3409 & w3407;
assign w17370 = ~w615 & w3407;
assign w17371 = ~w615 & w17369;
assign w17372 = ~w3413 & ~w3412;
assign w17373 = ~w3806 & ~w3412;
assign w17374 = ~w3806 & w17372;
assign w17375 = ~w3417 & ~w3416;
assign w17376 = w3810 & ~w3416;
assign w17377 = w3810 & w17375;
assign w17378 = ~w3226 & ~w3422;
assign w17379 = ~w3815 & ~w3814;
assign w17380 = w3815 & w3814;
assign w17381 = ~w3815 & w3819;
assign w17382 = w3815 & ~w1339;
assign w17383 = ~w3610 & ~w3608;
assign w17384 = w3825 & ~w3608;
assign w17385 = w3825 & w17383;
assign w17386 = w3601 & ~w3599;
assign w17387 = ~w3441 & ~w3439;
assign w17388 = ~w3834 & ~w3439;
assign w17389 = ~w3834 & w17387;
assign w17390 = ~w3582 & ~w3581;
assign w17391 = w3839 & ~w3581;
assign w17392 = w3839 & w17390;
assign w17393 = w3090 & ~w3493;
assign w17394 = w15862 & ~w3494;
assign w17395 = (~w3494 & w15862) | (~w3494 & ~w3090) | (w15862 & ~w3090);
assign w17396 = w3476 & w3870;
assign w17397 = ~pi271 & ~w3473;
assign w17398 = ~w3474 & w3875;
assign w17399 = w3474 & w3873;
assign w17400 = w3873 & ~w3878;
assign w17401 = ~w3487 & ~w3886;
assign w17402 = w3487 & w3886;
assign w17403 = ~pi322 & ~w3571;
assign w17404 = pi322 & w3571;
assign w17405 = w3574 & ~w3572;
assign w17406 = w3447 & ~w3586;
assign w17407 = ~w3446 & ~w3444;
assign w17408 = w3997 & ~w3444;
assign w17409 = w3997 & w17407;
assign w17410 = ~w3418 & ~w3623;
assign w17411 = w3401 & ~w3647;
assign w17412 = ~w3400 & ~w3656;
assign w17413 = w3791 & ~w135;
assign w17414 = ~pi273 & pi161;
assign w17415 = ~pi273 & ~w4043;
assign w17416 = w535 & pi336;
assign w17417 = ~w3796 & ~w3795;
assign w17418 = ~w4032 & ~w3799;
assign w17419 = ~w3809 & ~w3807;
assign w17420 = ~w3813 & ~w3811;
assign w17421 = ~w3828 & ~w3827;
assign w17422 = w4006 & ~w3832;
assign w17423 = ~w3837 & ~w3836;
assign w17424 = w4097 & w3836;
assign w17425 = w4097 & ~w17423;
assign w17426 = ~w4000 & ~w3998;
assign w17427 = ~w3847 & ~w3846;
assign w17428 = ~w4124 & ~w4128;
assign w17429 = w4124 & w4128;
assign w17430 = ~w3476 & ~w3866;
assign w17431 = w3476 & w3866;
assign w17432 = w4139 & ~w4138;
assign w17433 = ~w4134 & w4138;
assign w17434 = ~w4134 & ~w17432;
assign w17435 = ~w4142 & w4118;
assign w17436 = w4142 & ~w4118;
assign w17437 = ~w3912 & ~w3914;
assign w17438 = ~w3966 & ~w3964;
assign w17439 = w3562 & ~w3564;
assign w17440 = ~w4243 & ~w3565;
assign w17441 = w3983 & ~w3981;
assign w17442 = w3563 & pi324;
assign w17443 = ~w3842 & ~w3840;
assign w17444 = w4257 & w3840;
assign w17445 = w4257 & ~w17443;
assign w17446 = w3993 & ~w3990;
assign w17447 = w4286 & w1602;
assign w17448 = ~w4286 & ~w1602;
assign w17449 = ~w4015 & ~w4018;
assign w17450 = ~w3805 & ~w3804;
assign w17451 = ~w460 & pi337;
assign w17452 = ~w3792 & ~w4322;
assign w17453 = w3792 & w466;
assign w17454 = ~w4050 & ~w3791;
assign w17455 = w3779 & ~w3775;
assign w17456 = w3770 & ~w3678;
assign w17457 = ~w1679 & pi314;
assign w17458 = ~w3747 & ~w3695;
assign w17459 = w3737 & ~w3731;
assign w17460 = ~w3724 & ~w3699;
assign w17461 = ~w3701 & ~w3720;
assign w17462 = pi143 & ~w3705;
assign w17463 = w4370 & w3705;
assign w17464 = w4370 & ~w17462;
assign w17465 = ~pi144 & pi141;
assign w17466 = ~pi144 & ~pi142;
assign w17467 = pi143 & ~w4370;
assign w17468 = ~w3703 & ~w3714;
assign w17469 = ~w3740 & ~w3697;
assign w17470 = ~w3750 & ~w3689;
assign w17471 = ~w1413 & pi313;
assign w17472 = w3758 & ~w3756;
assign w17473 = ~w3761 & ~w3684;
assign w17474 = w3680 & ~w3766;
assign w17475 = ~w3673 & ~w3671;
assign w17476 = ~w3669 & ~w3668;
assign w17477 = ~pi274 & pi161;
assign w17478 = ~w4340 & ~w4491;
assign w17479 = ~w4341 & ~w3789;
assign w17480 = ~w4342 & ~w4466;
assign w17481 = w4461 & ~w4459;
assign w17482 = ~w4435 & ~w4432;
assign w17483 = ~w1413 & pi312;
assign w17484 = ~w1679 & pi313;
assign w17485 = ~w4396 & ~w4362;
assign w17486 = ~pi144 & ~w4523;
assign w17487 = ~w4526 & ~w4527;
assign w17488 = ~w4527 & ~w4532;
assign w17489 = ~w4369 & pi145;
assign w17490 = pi145 & pi141;
assign w17491 = pi141 & ~w4520;
assign w17492 = w4538 & pi321;
assign w17493 = ~w4367 & ~w4386;
assign w17494 = ~w4365 & ~w4392;
assign w17495 = w4402 & ~w4359;
assign w17496 = ~w4407 & ~w4567;
assign w17497 = w4407 & w4567;
assign w17498 = ~w4413 & ~w4354;
assign w17499 = w4420 & ~w4417;
assign w17500 = ~w4423 & ~w4427;
assign w17501 = w4348 & ~w4440;
assign w17502 = ~w4445 & w4608;
assign w17503 = w4617 & ~w4445;
assign w17504 = w4611 & w4445;
assign w17505 = w4445 & ~w4346;
assign w17506 = ~w4344 & ~w4452;
assign w17507 = ~w4075 & w4662;
assign w17508 = w4075 & ~w4662;
assign w17509 = w4308 & w955;
assign w17510 = ~w4308 & w4668;
assign w17511 = pi333 & w4668;
assign w17512 = pi333 & w17510;
assign w17513 = ~w4308 & ~w4668;
assign w17514 = w4308 & ~w955;
assign w17515 = ~pi333 & w4668;
assign w17516 = ~pi333 & w17510;
assign w17517 = ~w4678 & ~w4677;
assign w17518 = ~w4086 & ~w4084;
assign w17519 = ~w4298 & ~w4297;
assign w17520 = ~w4096 & ~w4094;
assign w17521 = w4692 & w4094;
assign w17522 = w4692 & ~w17520;
assign w17523 = ~w4100 & ~w4099;
assign w17524 = w4696 & w4099;
assign w17525 = w4696 & ~w17523;
assign w17526 = w4267 & ~w4264;
assign w17527 = w4253 & ~w4251;
assign w17528 = w3976 & ~w4242;
assign w17529 = ~w4126 & ~w4128;
assign w17530 = ~w4126 & ~w17429;
assign w17531 = w4743 & ~w17529;
assign w17532 = w4743 & ~w17530;
assign w17533 = ~w4134 & ~w4132;
assign w17534 = w4749 & w4132;
assign w17535 = w4749 & ~w17533;
assign w17536 = ~w4145 & ~w4143;
assign w17537 = ~w4755 & ~w4143;
assign w17538 = ~w4755 & w17536;
assign w17539 = w15869 & ~w4758;
assign w17540 = (~w4758 & w15869) | (~w4758 & w4152) | (w15869 & w4152);
assign w17541 = ~w4152 & w15870;
assign w17542 = ~w4106 & w4218;
assign w17543 = ~w4260 & ~w4259;
assign w17544 = w3563 & pi325;
assign w17545 = pi324 & ~w4866;
assign w17546 = ~pi324 & w4866;
assign w17547 = w4889 & ~w4090;
assign w17548 = w4889 & w16139;
assign w17549 = w4287 & w4897;
assign w17550 = w4899 & ~w4290;
assign w17551 = ~w4081 & ~w4079;
assign w17552 = w535 & pi337;
assign w17553 = ~w971 & pi338;
assign w17554 = w4480 & ~w4338;
assign w17555 = w4955 & ~w4658;
assign w17556 = ~w4658 & ~w135;
assign w17557 = ~pi275 & pi161;
assign w17558 = w4659 & w466;
assign w17559 = ~w460 & pi339;
assign w17560 = ~w4659 & ~w4972;
assign w17561 = w537 & ~w4939;
assign w17562 = w537 & w16141;
assign w17563 = pi338 & ~w17561;
assign w17564 = pi338 & ~w17562;
assign w17565 = ~w4312 & ~w4311;
assign w17566 = w2170 & ~w4895;
assign w17567 = w4890 & w5012;
assign w17568 = ~w4890 & ~w5012;
assign w17569 = w3563 & pi326;
assign w17570 = w4861 & ~w4865;
assign w17571 = ~w4845 & w4844;
assign w17572 = w3476 & w16160;
assign w17573 = ~w5067 & ~w4741;
assign w17574 = ~w5064 & ~w4741;
assign w17575 = ~w5064 & w17573;
assign w17576 = w5070 & w5059;
assign w17577 = ~w5070 & ~w5059;
assign w17578 = (~w4748 & w16161) | (~w4748 & ~w4132) | (w16161 & ~w4132);
assign w17579 = (~w4748 & w16161) | (~w4748 & w17533) | (w16161 & w17533);
assign w17580 = w5073 & ~w17579;
assign w17581 = w5073 & ~w17578;
assign w17582 = ~w745 & w747;
assign w17583 = w4792 & ~w4793;
assign w17584 = ~w4797 & ~w4802;
assign w17585 = w5216 & ~w5213;
assign w17586 = w5139 & ~w5138;
assign w17587 = w6049 & w5479;
assign w17588 = w6049 & ~w16595;
assign w17589 = w6058 & w5485;
assign w17590 = w6058 & ~w16596;
assign w17591 = ~w6062 & ~w5489;
assign w17592 = ~w6062 & w16597;
assign w17593 = ~w5641 & ~w5639;
assign w17594 = w6854 & ~w6855;
assign w17595 = ~w6045 & ~w6847;
assign w17596 = w6322 & ~w6336;
assign w17597 = ~w6891 & ~w6303;
assign w17598 = ~w6891 & w15913;
assign w17599 = w6904 & ~w15914;
assign w17600 = w6904 & w6293;
assign w17601 = w7464 & w7188;
assign w17602 = w7464 & ~w16445;
assign w17603 = w7468 & w6863;
assign w17604 = w7468 & ~w16446;
assign w17605 = ~w2373 & w7486;
assign w17606 = ~w7041 & ~w16442;
assign w17607 = ~w7041 & ~w16441;
assign w17608 = w7803 & w6858;
assign w17609 = w7803 & ~w16455;
assign w17610 = ~w7437 & ~w7436;
assign w17611 = w8332 & ~w8328;
assign w17612 = ~w8781 & ~w8777;
assign w17613 = ~w11243 & w11899;
assign w17614 = w11243 & ~w11899;
assign w17615 = ~w11079 & w11254;
assign w17616 = w5648 & ~w6229;
assign w17617 = w16512 & w5043;
assign w17618 = w5047 & ~w6112;
assign w17619 = ~w5047 & w6112;
assign w17620 = (~w112 & ~w16633) | (~w112 & ~w110) | (~w16633 & ~w110);
assign w17621 = (w512 & ~w16841) | (w512 & ~w538) | (~w16841 & ~w538);
assign w17622 = (w649 & ~w658) | (w649 & w16544) | (~w658 & w16544);
assign w17623 = (w655 & w650) | (w655 & ~w16087) | (w650 & ~w16087);
assign w17624 = (~w772 & ~w787) | (~w772 & w16892) | (~w787 & w16892);
assign w17625 = (w617 & ~w16894) | (w617 & ~w796) | (~w16894 & ~w796);
assign w17626 = (~w1010 & w16907) | (~w1010 & ~w969) | (w16907 & ~w969);
assign w17627 = (w15806 & ~w870) | (w15806 & ~w871) | (~w870 & ~w871);
assign w17628 = (~w1012 & w16949) | (~w1012 & ~w1111) | (w16949 & ~w1111);
assign w17629 = (w1038 & ~w15808) | (w1038 & ~w1035) | (~w15808 & ~w1035);
assign w17630 = w16335 & ~w1035;
assign w17631 = (w1301 & ~w15814) | (w1301 & ~w1291) | (~w15814 & ~w1291);
assign w17632 = (~w1303 & w15815) | (~w1303 & ~w1292) | (w15815 & ~w1292);
assign w17633 = (w1675 & ~w17013) | (w1675 & ~w1677) | (~w17013 & ~w1677);
assign w17634 = (~w1297 & ~w1524) | (~w1297 & w17630) | (~w1524 & w17630);
assign w17635 = (~pi130 & ~w16109) | (~pi130 & ~w1291) | (~w16109 & ~w1291);
assign w17636 = (w1479 & ~w17041) | (w1479 & ~w1640) | (~w17041 & ~w1640);
assign w17637 = (pi137 & w17014) | (pi137 & ~w849) | (w17014 & ~w849);
assign w17638 = ~w1529 & ~w1786;
assign w17639 = (~w1795 & w15830) | (~w1795 & w17638) | (w15830 & w17638);
assign w17640 = (w2143 & w15834) | (w2143 & ~w1587) | (w15834 & ~w1587);
assign w17641 = (~w2039 & w17097) | (~w2039 & ~w2219) | (w17097 & ~w2219);
assign w17642 = (~w2046 & w17101) | (~w2046 & ~w2193) | (w17101 & ~w2193);
assign w17643 = (w17114 & w17115) | (w17114 & ~w1790) | (w17115 & ~w1790);
assign w17644 = (~w1955 & ~w17143) | (~w1955 & ~w1699) | (~w17143 & ~w1699);
assign w17645 = (~w2252 & w17158) | (~w2252 & ~w2427) | (w17158 & ~w2427);
assign w17646 = (~w2421 & w17182) | (~w2421 & ~w2417) | (w17182 & ~w2417);
assign w17647 = (~w2266 & w15844) | (~w2266 & ~w2360) | (w15844 & ~w2360);
assign w17648 = (w15852 & ~w2899) | (w15852 & ~w2900) | (~w2899 & ~w2900);
assign w17649 = (w15855 & ~w2943) | (w15855 & ~w2944) | (~w2943 & ~w2944);
assign w17650 = ~w653 & w2992;
assign w17651 = (w3012 & ~w17308) | (w3012 & ~w3235) | (~w17308 & ~w3235);
assign w17652 = (~w3016 & w17311) | (~w3016 & ~w3232) | (w17311 & ~w3232);
assign w17653 = (~w3031 & w17320) | (~w3031 & ~w3207) | (w17320 & ~w3207);
assign w17654 = (~w3063 & w15858) | (~w3063 & w17724) | (w15858 & w17724);
assign w17655 = (~w3069 & w17327) | (~w3069 & ~w3073) | (w17327 & ~w3073);
assign w17656 = (w3078 & ~w15859) | (w3078 & ~w3086) | (~w15859 & ~w3086);
assign w17657 = (~w3272 & w17344) | (~w3272 & ~w3394) | (w17344 & ~w3394);
assign w17658 = (~w3407 & ~w17369) | (~w3407 & ~w3634) | (~w17369 & ~w3634);
assign w17659 = (w3412 & ~w17372) | (w3412 & ~w3631) | (~w17372 & ~w3631);
assign w17660 = (w3416 & ~w17375) | (w3416 & ~w3628) | (~w17375 & ~w3628);
assign w17661 = (w3608 & ~w17383) | (w3608 & ~w3604) | (~w17383 & ~w3604);
assign w17662 = (w3439 & ~w17387) | (w3439 & ~w3594) | (~w17387 & ~w3594);
assign w17663 = (w3581 & ~w17390) | (w3581 & ~w3577) | (~w17390 & ~w3577);
assign w17664 = (w3444 & ~w17407) | (w3444 & ~w3591) | (~w17407 & ~w3591);
assign w17665 = (~w3836 & w17423) | (~w3836 & ~w4003) | (w17423 & ~w4003);
assign w17666 = (w3923 & ~w4179) | (w3923 & w16581) | (~w4179 & w16581);
assign w17667 = (w3919 & w3920) | (w3919 & ~w15864) | (w3920 & ~w15864);
assign w17668 = (~w3840 & w17443) | (~w3840 & ~w3986) | (w17443 & ~w3986);
assign w17669 = (~w4094 & w17520) | (~w4094 & ~w4279) | (w17520 & ~w4279);
assign w17670 = (~w4099 & w17523) | (~w4099 & ~w4276) | (w17523 & ~w4276);
assign w17671 = ~w4126 & ~w4130;
assign w17672 = (~w4132 & w17533) | (~w4132 & ~w4140) | (w17533 & ~w4140);
assign w17673 = (w4143 & ~w17536) | (w4143 & ~w4146) | (~w17536 & ~w4146);
assign w17674 = (w4174 & w4175) | (w4174 & ~w15868) | (w4175 & ~w15868);
assign w17675 = (w4090 & ~w16139) | (w4090 & ~w4282) | (~w16139 & ~w4282);
assign w17676 = (w4991 & ~w15872) | (w4991 & ~w4917) | (~w15872 & ~w4917);
assign w17677 = (w4898 & w4895) | (w4898 & ~w16159) | (w4895 & ~w16159);
assign w17678 = (~w4901 & w2170) | (~w4901 & w17566) | (w2170 & w17566);
assign w17679 = (~w4241 & ~w15873) | (~w4241 & ~w5035) | (~w15873 & ~w5035);
assign w17680 = (w4620 & ~w15884) | (w4620 & ~w4625) | (~w15884 & ~w4625);
assign w17681 = (~w5485 & w16596) | (~w5485 & ~w5779) | (w16596 & ~w5779);
assign w17682 = (w5489 & ~w16597) | (w5489 & ~w5776) | (~w16597 & ~w5776);
assign w17683 = (~w5749 & w16180) | (~w5749 & ~w5746) | (w16180 & ~w5746);
assign w17684 = (~w5507 & w16181) | (~w5507 & ~w5743) | (w16181 & ~w5743);
assign w17685 = (~w6301 & w15899) | (~w6301 & ~w5733) | (w15899 & ~w5733);
assign w17686 = (~w6327 & w15900) | (~w6327 & ~w5762) | (w15900 & ~w5762);
assign w17687 = (w15909 & ~w5834) | (w15909 & ~w5835) | (~w5834 & ~w5835);
assign w17688 = (w6017 & ~w15910) | (w6017 & ~w6372) | (~w15910 & ~w6372);
assign w17689 = (~w6348 & ~w6874) | (~w6348 & w16607) | (~w6874 & w16607);
assign w17690 = (w15914 & ~w6293) | (w15914 & ~w6295) | (~w6293 & ~w6295);
assign w17691 = (~w7188 & w16445) | (~w7188 & ~w7180) | (w16445 & ~w7180);
assign w17692 = (~w6863 & w16446) | (~w6863 & ~w7174) | (w16446 & ~w7174);
assign w17693 = (~pi330 & ~w7496) | (~pi330 & ~w16449) | (~w7496 & ~w16449);
assign w17694 = (~w6858 & w16455) | (~w6858 & ~w7177) | (w16455 & ~w7177);
assign w17695 = (~w8163 & w15938) | (~w8163 & ~w8364) | (w15938 & ~w8364);
assign w17696 = (~w9548 & ~w15940) | (~w9548 & ~w8804) | (~w15940 & ~w8804);
assign w17697 = (w8575 & ~w16214) | (w8575 & ~w8872) | (~w16214 & ~w8872);
assign w17698 = (w15962 & ~w9792) | (w15962 & ~w9794) | (~w9792 & ~w9794);
assign w17699 = (w10286 & ~w15963) | (w10286 & ~w10284) | (~w15963 & ~w10284);
assign w17700 = (~w10667 & w15970) | (~w10667 & ~w10664) | (w15970 & ~w10664);
assign w17701 = (~w10237 & w15972) | (~w10237 & ~w10658) | (w15972 & ~w10658);
assign w17702 = (~w9880 & w16260) | (~w9880 & ~w9876) | (w16260 & ~w9876);
assign w17703 = (w12164 & ~w16305) | (w12164 & ~w12156) | (~w16305 & ~w12156);
assign w17704 = (w16306 & ~w12172) | (w16306 & ~w12174) | (~w12172 & ~w12174);
assign w17705 = (w12928 & w12926) | (w12928 & ~w16032) | (w12926 & ~w16032);
assign w17706 = (~w12930 & ~w13508) | (~w12930 & w16316) | (~w13508 & w16316);
assign w17707 = (~pi293 & ~w16043) | (~pi293 & ~w14036) | (~w16043 & ~w14036);
assign w17708 = (~w14047 & w16321) | (~w14047 & ~w14044) | (w16321 & ~w14044);
assign w17709 = (~w13202 & w16045) | (~w13202 & ~w14532) | (w16045 & ~w14532);
assign w17710 = (~w14534 & w16046) | (~w14534 & ~w14532) | (w16046 & ~w14532);
assign w17711 = (~w13758 & w16049) | (~w13758 & ~w14027) | (w16049 & ~w14027);
assign w17712 = (~w2676 & ~w15846) | (~w2676 & ~w3160) | (~w15846 & ~w3160);
assign w17713 = (w955 & ~w15849) | (w955 & ~w3221) | (~w15849 & ~w3221);
assign w17714 = (w4101 & w16061) | (w4101 & ~w4270) | (w16061 & ~w4270);
assign w17715 = (~w4660 & w16062) | (~w4660 & ~w4923) | (w16062 & ~w4923);
assign w17716 = (w4914 & w16063) | (w4914 & ~w4910) | (w16063 & ~w4910);
assign w17717 = w5499 & w2698;
assign w17718 = (~w6019 & ~w16074) | (~w6019 & ~w6366) | (~w16074 & ~w6366);
assign w17719 = pi265 & pi264;
assign w17720 = ~w3183 & w2698;
assign w17721 = ~w615 & ~w793;
assign w17722 = pi324 & pi322;
assign w17723 = (~w3059 & ~w17245) | (~w3059 & ~w2285) | (~w17245 & ~w2285);
assign w17724 = ~w2603 & w17723;
assign one = 1;
assign po000 = pi194;// level 0
assign po001 = pi195;// level 0
assign po002 = pi206;// level 0
assign po003 = pi217;// level 0
assign po004 = pi220;// level 0
assign po005 = pi221;// level 0
assign po006 = pi222;// level 0
assign po007 = pi223;// level 0
assign po008 = pi224;// level 0
assign po009 = pi225;// level 0
assign po010 = pi196;// level 0
assign po011 = pi197;// level 0
assign po012 = pi198;// level 0
assign po013 = pi199;// level 0
assign po014 = pi200;// level 0
assign po015 = pi201;// level 0
assign po016 = pi202;// level 0
assign po017 = pi203;// level 0
assign po018 = pi204;// level 0
assign po019 = pi205;// level 0
assign po020 = pi207;// level 0
assign po021 = pi208;// level 0
assign po022 = pi209;// level 0
assign po023 = pi210;// level 0
assign po024 = pi211;// level 0
assign po025 = pi212;// level 0
assign po026 = pi213;// level 0
assign po027 = pi214;// level 0
assign po028 = pi215;// level 0
assign po029 = pi216;// level 0
assign po030 = pi218;// level 0
assign po031 = pi219;// level 0
assign po032 = pi226;// level 0
assign po033 = pi227;// level 0
assign po034 = pi238;// level 0
assign po035 = pi249;// level 0
assign po036 = pi252;// level 0
assign po037 = pi253;// level 0
assign po038 = pi254;// level 0
assign po039 = pi255;// level 0
assign po040 = pi256;// level 0
assign po041 = pi257;// level 0
assign po042 = pi228;// level 0
assign po043 = pi229;// level 0
assign po044 = pi230;// level 0
assign po045 = pi231;// level 0
assign po046 = pi232;// level 0
assign po047 = pi233;// level 0
assign po048 = pi234;// level 0
assign po049 = pi235;// level 0
assign po050 = pi236;// level 0
assign po051 = pi237;// level 0
assign po052 = pi239;// level 0
assign po053 = pi240;// level 0
assign po054 = pi241;// level 0
assign po055 = pi242;// level 0
assign po056 = pi243;// level 0
assign po057 = pi244;// level 0
assign po058 = pi245;// level 0
assign po059 = pi246;// level 0
assign po060 = pi247;// level 0
assign po061 = pi248;// level 0
assign po062 = pi250;// level 0
assign po063 = pi251;// level 0
assign po064 = pi162;// level 0
assign po065 = pi163;// level 0
assign po066 = pi174;// level 0
assign po067 = pi185;// level 0
assign po068 = pi188;// level 0
assign po069 = pi189;// level 0
assign po070 = pi190;// level 0
assign po071 = pi191;// level 0
assign po072 = pi192;// level 0
assign po073 = pi193;// level 0
assign po074 = pi164;// level 0
assign po075 = pi165;// level 0
assign po076 = pi166;// level 0
assign po077 = pi167;// level 0
assign po078 = pi168;// level 0
assign po079 = pi169;// level 0
assign po080 = pi170;// level 0
assign po081 = pi171;// level 0
assign po082 = pi172;// level 0
assign po083 = pi173;// level 0
assign po084 = pi175;// level 0
assign po085 = pi176;// level 0
assign po086 = pi177;// level 0
assign po087 = pi178;// level 0
assign po088 = pi179;// level 0
assign po089 = pi180;// level 0
assign po090 = pi181;// level 0
assign po091 = pi182;// level 0
assign po092 = pi183;// level 0
assign po093 = pi184;// level 0
assign po094 = pi186;// level 0
assign po095 = pi187;// level 0
assign po096 = w138;// level 13
assign po097 = ~w141;// level 13
assign po098 = ~w144;// level 13
assign po099 = ~w147;// level 13
assign po100 = ~w150;// level 13
assign po101 = ~w153;// level 13
assign po102 = ~w156;// level 13
assign po103 = ~w159;// level 13
assign po104 = ~w162;// level 13
assign po105 = ~w165;// level 13
assign po106 = ~w168;// level 13
assign po107 = ~w171;// level 13
assign po108 = ~w174;// level 13
assign po109 = ~w177;// level 13
assign po110 = ~w180;// level 13
assign po111 = ~w184;// level 13
assign po112 = ~w187;// level 13
assign po113 = ~w191;// level 13
assign po114 = ~w195;// level 13
assign po115 = ~w198;// level 13
assign po116 = ~w201;// level 13
assign po117 = ~w205;// level 13
assign po118 = ~w209;// level 13
assign po119 = ~w213;// level 13
assign po120 = ~w216;// level 13
assign po121 = ~w219;// level 13
assign po122 = w222;// level 13
assign po123 = ~w225;// level 13
assign po124 = ~w228;// level 13
assign po125 = ~w231;// level 13
assign po126 = ~w234;// level 13
assign po127 = ~w237;// level 13
assign po128 = ~w240;// level 13
assign po129 = ~w243;// level 13
assign po130 = ~w247;// level 13
assign po131 = ~w250;// level 13
assign po132 = ~w253;// level 13
assign po133 = ~w256;// level 13
assign po134 = ~w259;// level 13
assign po135 = ~w262;// level 13
assign po136 = ~w265;// level 13
assign po137 = ~w268;// level 13
assign po138 = ~w271;// level 13
assign po139 = ~w274;// level 13
assign po140 = ~w277;// level 13
assign po141 = ~w281;// level 13
assign po142 = ~w284;// level 13
assign po143 = ~w287;// level 13
assign po144 = ~w290;// level 13
assign po145 = ~w293;// level 13
assign po146 = ~w296;// level 13
assign po147 = ~w299;// level 13
assign po148 = ~w302;// level 13
assign po149 = ~w305;// level 13
assign po150 = ~w308;// level 13
assign po151 = ~w311;// level 13
assign po152 = ~w315;// level 13
assign po153 = ~w319;// level 13
assign po154 = ~w322;// level 13
assign po155 = ~w325;// level 13
assign po156 = ~w329;// level 13
assign po157 = ~w332;// level 13
assign po158 = ~w336;// level 13
assign po159 = ~w340;// level 13
assign po160 = ~w343;// level 13
assign po161 = ~w346;// level 13
assign po162 = ~w350;// level 13
assign po163 = ~w353;// level 13
assign po164 = ~w356;// level 13
assign po165 = ~w359;// level 13
assign po166 = ~w362;// level 13
assign po167 = ~w365;// level 13
assign po168 = ~w368;// level 13
assign po169 = ~w371;// level 13
assign po170 = ~w374;// level 13
assign po171 = ~w377;// level 13
assign po172 = ~w380;// level 13
assign po173 = ~w384;// level 13
assign po174 = ~w387;// level 13
assign po175 = ~w390;// level 13
assign po176 = ~w393;// level 13
assign po177 = ~w396;// level 13
assign po178 = ~w399;// level 13
assign po179 = ~w402;// level 13
assign po180 = ~w405;// level 13
assign po181 = ~w408;// level 13
assign po182 = ~w411;// level 13
assign po183 = ~w414;// level 13
assign po184 = ~w417;// level 13
assign po185 = ~w420;// level 13
assign po186 = ~w423;// level 13
assign po187 = ~w426;// level 13
assign po188 = ~w429;// level 13
assign po189 = ~w432;// level 13
assign po190 = ~w435;// level 13
assign po191 = ~w438;// level 13
assign po192 = ~w441;// level 13
assign po193 = w454;// level 15
assign po194 = w489;// level 15
assign po195 = w564;// level 20
assign po196 = w677;// level 31
assign po197 = w836;// level 36
assign po198 = w1005;// level 46
assign po199 = w1204;// level 52
assign po200 = w1399;// level 63
assign po201 = w1663;// level 73
assign po202 = w1930;// level 78
assign po203 = w2243;// level 88
assign po204 = w2548;// level 94
assign po205 = w2887;// level 98
assign po206 = w3267;// level 109
assign po207 = w3663;// level 117
assign po208 = w4060;// level 122
assign po209 = w4488;// level 126
assign po210 = w4966;// level 136
assign po211 = w5462;// level 142
assign po212 = w6011;// level 147
assign po213 = w6597;// level 158
assign po214 = w7226;// level 162
assign po215 = w7858;// level 169
assign po216 = w8521;// level 176
assign po217 = w9199;// level 182
assign po218 = w9942;// level 192
assign po219 = w10703;// level 195
assign po220 = w11494;// level 201
assign po221 = w12302;// level 206
assign po222 = w13192;// level 212
assign po223 = w14066;// level 216
assign po224 = ~w14930;// level 219
assign po225 = w15064;// level 175
assign po226 = w15073;// level 164
assign po227 = w15082;// level 156
assign po228 = w15091;// level 147
assign po229 = w15100;// level 141
assign po230 = w15109;// level 136
assign po231 = w15118;// level 132
assign po232 = w15127;// level 127
assign po233 = w15136;// level 120
assign po234 = w15145;// level 113
assign po235 = w15154;// level 107
assign po236 = w15163;// level 104
assign po237 = w15172;// level 98
assign po238 = w15181;// level 93
assign po239 = w15190;// level 89
assign po240 = w15199;// level 82
assign po241 = w15208;// level 78
assign po242 = w15217;// level 73
assign po243 = w15226;// level 67
assign po244 = w15235;// level 60
assign po245 = w15244;// level 57
assign po246 = w15253;// level 52
assign po247 = w15262;// level 48
assign po248 = w15271;// level 41
assign po249 = w15280;// level 37
assign po250 = w15289;// level 30
assign po251 = w15298;// level 28
assign po252 = w15307;// level 20
assign po253 = w15316;// level 16
assign po254 = w15324;// level 15
assign po255 = w15332;// level 15
assign po256 = w15340;// level 17
assign po257 = w15347;// level 16
assign po258 = w15359;// level 15
assign po259 = w15372;// level 15
assign po260 = w15385;// level 15
assign po261 = w15399;// level 17
assign po262 = w15413;// level 19
assign po263 = w15427;// level 22
assign po264 = w15441;// level 26
assign po265 = w15455;// level 30
assign po266 = w15469;// level 32
assign po267 = w15484;// level 35
assign po268 = w15499;// level 38
assign po269 = w15514;// level 41
assign po270 = w15529;// level 44
assign po271 = w15544;// level 47
assign po272 = w15559;// level 50
assign po273 = w15574;// level 53
assign po274 = w15589;// level 56
assign po275 = w15604;// level 59
assign po276 = w15619;// level 62
assign po277 = w15634;// level 65
assign po278 = w15649;// level 68
assign po279 = w15664;// level 71
assign po280 = w15679;// level 74
assign po281 = w15694;// level 77
assign po282 = w15709;// level 80
assign po283 = w15724;// level 83
assign po284 = w15739;// level 86
assign po285 = w15754;// level 89
assign po286 = w15769;// level 92
assign po287 = w15784;// level 96
assign po288 = w15796;// level 99
endmodule
