// Benchmark "des_perf" written by ABC on Wed Apr 29 13:47:29 2015

module des_perf ( 
    pi0000, pi0001, pi0002, pi0003, pi0004, pi0005, pi0006, pi0007, pi0008,
    pi0009, pi0010, pi0011, pi0012, pi0013, pi0014, pi0015, pi0016, pi0017,
    pi0018, pi0019, pi0020, pi0021, pi0022, pi0023, pi0024, pi0025, pi0026,
    pi0027, pi0028, pi0029, pi0030, pi0031, pi0032, pi0033, pi0034, pi0035,
    pi0036, pi0037, pi0038, pi0039, pi0040, pi0041, pi0042, pi0043, pi0044,
    pi0045, pi0046, pi0047, pi0048, pi0049, pi0050, pi0051, pi0052, pi0053,
    pi0054, pi0055, pi0056, pi0057, pi0058, pi0059, pi0060, pi0061, pi0062,
    pi0063, pi0064, pi0065, pi0066, pi0067, pi0068, pi0069, pi0070, pi0071,
    pi0072, pi0073, pi0074, pi0075, pi0076, pi0077, pi0078, pi0079, pi0080,
    pi0081, pi0082, pi0083, pi0084, pi0085, pi0086, pi0087, pi0088, pi0089,
    pi0090, pi0091, pi0092, pi0093, pi0094, pi0095, pi0096, pi0097, pi0098,
    pi0099, pi0100, pi0101, pi0102, pi0103, pi0104, pi0105, pi0106, pi0107,
    pi0108, pi0109, pi0110, pi0111, pi0112, pi0113, pi0114, pi0115, pi0116,
    pi0117, pi0118, pi0119, pi0120, pi0121, pi0122, pi0123, pi0124, pi0125,
    pi0126, pi0127, pi0128, pi0129, pi0130, pi0131, pi0132, pi0133, pi0134,
    pi0135, pi0136, pi0137, pi0138, pi0139, pi0140, pi0141, pi0142, pi0143,
    pi0144, pi0145, pi0146, pi0147, pi0148, pi0149, pi0150, pi0151, pi0152,
    pi0153, pi0154, pi0155, pi0156, pi0157, pi0158, pi0159, pi0160, pi0161,
    pi0162, pi0163, pi0164, pi0165, pi0166, pi0167, pi0168, pi0169, pi0170,
    pi0171, pi0172, pi0173, pi0174, pi0175, pi0176, pi0177, pi0178, pi0179,
    pi0180, pi0181, pi0182, pi0183, pi0184, pi0185, pi0186, pi0187, pi0188,
    pi0189, pi0190, pi0191, pi0192, pi0193, pi0194, pi0195, pi0196, pi0197,
    pi0198, pi0199, pi0200, pi0201, pi0202, pi0203, pi0204, pi0205, pi0206,
    pi0207, pi0208, pi0209, pi0210, pi0211, pi0212, pi0213, pi0214, pi0215,
    pi0216, pi0217, pi0218, pi0219, pi0220, pi0221, pi0222, pi0223, pi0224,
    pi0225, pi0226, pi0227, pi0228, pi0229, pi0230, pi0231, pi0232, pi0233,
    pi0234, pi0235, pi0236, pi0237, pi0238, pi0239, pi0240, pi0241, pi0242,
    pi0243, pi0244, pi0245, pi0246, pi0247, pi0248, pi0249, pi0250, pi0251,
    pi0252, pi0253, pi0254, pi0255, pi0256, pi0257, pi0258, pi0259, pi0260,
    pi0261, pi0262, pi0263, pi0264, pi0265, pi0266, pi0267, pi0268, pi0269,
    pi0270, pi0271, pi0272, pi0273, pi0274, pi0275, pi0276, pi0277, pi0278,
    pi0279, pi0280, pi0281, pi0282, pi0283, pi0284, pi0285, pi0286, pi0287,
    pi0288, pi0289, pi0290, pi0291, pi0292, pi0293, pi0294, pi0295, pi0296,
    pi0297, pi0298, pi0299, pi0300, pi0301, pi0302, pi0303, pi0304, pi0305,
    pi0306, pi0307, pi0308, pi0309, pi0310, pi0311, pi0312, pi0313, pi0314,
    pi0315, pi0316, pi0317, pi0318, pi0319, pi0320, pi0321, pi0322, pi0323,
    pi0324, pi0325, pi0326, pi0327, pi0328, pi0329, pi0330, pi0331, pi0332,
    pi0333, pi0334, pi0335, pi0336, pi0337, pi0338, pi0339, pi0340, pi0341,
    pi0342, pi0343, pi0344, pi0345, pi0346, pi0347, pi0348, pi0349, pi0350,
    pi0351, pi0352, pi0353, pi0354, pi0355, pi0356, pi0357, pi0358, pi0359,
    pi0360, pi0361, pi0362, pi0363, pi0364, pi0365, pi0366, pi0367, pi0368,
    pi0369, pi0370, pi0371, pi0372, pi0373, pi0374, pi0375, pi0376, pi0377,
    pi0378, pi0379, pi0380, pi0381, pi0382, pi0383, pi0384, pi0385, pi0386,
    pi0387, pi0388, pi0389, pi0390, pi0391, pi0392, pi0393, pi0394, pi0395,
    pi0396, pi0397, pi0398, pi0399, pi0400, pi0401, pi0402, pi0403, pi0404,
    pi0405, pi0406, pi0407, pi0408, pi0409, pi0410, pi0411, pi0412, pi0413,
    pi0414, pi0415, pi0416, pi0417, pi0418, pi0419, pi0420, pi0421, pi0422,
    pi0423, pi0424, pi0425, pi0426, pi0427, pi0428, pi0429, pi0430, pi0431,
    pi0432, pi0433, pi0434, pi0435, pi0436, pi0437, pi0438, pi0439, pi0440,
    pi0441, pi0442, pi0443, pi0444, pi0445, pi0446, pi0447, pi0448, pi0449,
    pi0450, pi0451, pi0452, pi0453, pi0454, pi0455, pi0456, pi0457, pi0458,
    pi0459, pi0460, pi0461, pi0462, pi0463, pi0464, pi0465, pi0466, pi0467,
    pi0468, pi0469, pi0470, pi0471, pi0472, pi0473, pi0474, pi0475, pi0476,
    pi0477, pi0478, pi0479, pi0480, pi0481, pi0482, pi0483, pi0484, pi0485,
    pi0486, pi0487, pi0488, pi0489, pi0490, pi0491, pi0492, pi0493, pi0494,
    pi0495, pi0496, pi0497, pi0498, pi0499, pi0500, pi0501, pi0502, pi0503,
    pi0504, pi0505, pi0506, pi0507, pi0508, pi0509, pi0510, pi0511, pi0512,
    pi0513, pi0514, pi0515, pi0516, pi0517, pi0518, pi0519, pi0520, pi0521,
    pi0522, pi0523, pi0524, pi0525, pi0526, pi0527, pi0528, pi0529, pi0530,
    pi0531, pi0532, pi0533, pi0534, pi0535, pi0536, pi0537, pi0538, pi0539,
    pi0540, pi0541, pi0542, pi0543, pi0544, pi0545, pi0546, pi0547, pi0548,
    pi0549, pi0550, pi0551, pi0552, pi0553, pi0554, pi0555, pi0556, pi0557,
    pi0558, pi0559, pi0560, pi0561, pi0562, pi0563, pi0564, pi0565, pi0566,
    pi0567, pi0568, pi0569, pi0570, pi0571, pi0572, pi0573, pi0574, pi0575,
    pi0576, pi0577, pi0578, pi0579, pi0580, pi0581, pi0582, pi0583, pi0584,
    pi0585, pi0586, pi0587, pi0588, pi0589, pi0590, pi0591, pi0592, pi0593,
    pi0594, pi0595, pi0596, pi0597, pi0598, pi0599, pi0600, pi0601, pi0602,
    pi0603, pi0604, pi0605, pi0606, pi0607, pi0608, pi0609, pi0610, pi0611,
    pi0612, pi0613, pi0614, pi0615, pi0616, pi0617, pi0618, pi0619, pi0620,
    pi0621, pi0622, pi0623, pi0624, pi0625, pi0626, pi0627, pi0628, pi0629,
    pi0630, pi0631, pi0632, pi0633, pi0634, pi0635, pi0636, pi0637, pi0638,
    pi0639, pi0640, pi0641, pi0642, pi0643, pi0644, pi0645, pi0646, pi0647,
    pi0648, pi0649, pi0650, pi0651, pi0652, pi0653, pi0654, pi0655, pi0656,
    pi0657, pi0658, pi0659, pi0660, pi0661, pi0662, pi0663, pi0664, pi0665,
    pi0666, pi0667, pi0668, pi0669, pi0670, pi0671, pi0672, pi0673, pi0674,
    pi0675, pi0676, pi0677, pi0678, pi0679, pi0680, pi0681, pi0682, pi0683,
    pi0684, pi0685, pi0686, pi0687, pi0688, pi0689, pi0690, pi0691, pi0692,
    pi0693, pi0694, pi0695, pi0696, pi0697, pi0698, pi0699, pi0700, pi0701,
    pi0702, pi0703, pi0704, pi0705, pi0706, pi0707, pi0708, pi0709, pi0710,
    pi0711, pi0712, pi0713, pi0714, pi0715, pi0716, pi0717, pi0718, pi0719,
    pi0720, pi0721, pi0722, pi0723, pi0724, pi0725, pi0726, pi0727, pi0728,
    pi0729, pi0730, pi0731, pi0732, pi0733, pi0734, pi0735, pi0736, pi0737,
    pi0738, pi0739, pi0740, pi0741, pi0742, pi0743, pi0744, pi0745, pi0746,
    pi0747, pi0748, pi0749, pi0750, pi0751, pi0752, pi0753, pi0754, pi0755,
    pi0756, pi0757, pi0758, pi0759, pi0760, pi0761, pi0762, pi0763, pi0764,
    pi0765, pi0766, pi0767, pi0768, pi0769, pi0770, pi0771, pi0772, pi0773,
    pi0774, pi0775, pi0776, pi0777, pi0778, pi0779, pi0780, pi0781, pi0782,
    pi0783, pi0784, pi0785, pi0786, pi0787, pi0788, pi0789, pi0790, pi0791,
    pi0792, pi0793, pi0794, pi0795, pi0796, pi0797, pi0798, pi0799, pi0800,
    pi0801, pi0802, pi0803, pi0804, pi0805, pi0806, pi0807, pi0808, pi0809,
    pi0810, pi0811, pi0812, pi0813, pi0814, pi0815, pi0816, pi0817, pi0818,
    pi0819, pi0820, pi0821, pi0822, pi0823, pi0824, pi0825, pi0826, pi0827,
    pi0828, pi0829, pi0830, pi0831, pi0832, pi0833, pi0834, pi0835, pi0836,
    pi0837, pi0838, pi0839, pi0840, pi0841, pi0842, pi0843, pi0844, pi0845,
    pi0846, pi0847, pi0848, pi0849, pi0850, pi0851, pi0852, pi0853, pi0854,
    pi0855, pi0856, pi0857, pi0858, pi0859, pi0860, pi0861, pi0862, pi0863,
    pi0864, pi0865, pi0866, pi0867, pi0868, pi0869, pi0870, pi0871, pi0872,
    pi0873, pi0874, pi0875, pi0876, pi0877, pi0878, pi0879, pi0880, pi0881,
    pi0882, pi0883, pi0884, pi0885, pi0886, pi0887, pi0888, pi0889, pi0890,
    pi0891, pi0892, pi0893, pi0894, pi0895, pi0896, pi0897, pi0898, pi0899,
    pi0900, pi0901, pi0902, pi0903, pi0904, pi0905, pi0906, pi0907, pi0908,
    pi0909, pi0910, pi0911, pi0912, pi0913, pi0914, pi0915, pi0916, pi0917,
    pi0918, pi0919, pi0920, pi0921, pi0922, pi0923, pi0924, pi0925, pi0926,
    pi0927, pi0928, pi0929, pi0930, pi0931, pi0932, pi0933, pi0934, pi0935,
    pi0936, pi0937, pi0938, pi0939, pi0940, pi0941, pi0942, pi0943, pi0944,
    pi0945, pi0946, pi0947, pi0948, pi0949, pi0950, pi0951, pi0952, pi0953,
    pi0954, pi0955, pi0956, pi0957, pi0958, pi0959, pi0960, pi0961, pi0962,
    pi0963, pi0964, pi0965, pi0966, pi0967, pi0968, pi0969, pi0970, pi0971,
    pi0972, pi0973, pi0974, pi0975, pi0976, pi0977, pi0978, pi0979, pi0980,
    pi0981, pi0982, pi0983, pi0984, pi0985, pi0986, pi0987, pi0988, pi0989,
    pi0990, pi0991, pi0992, pi0993, pi0994, pi0995, pi0996, pi0997, pi0998,
    pi0999, pi1000, pi1001, pi1002, pi1003, pi1004, pi1005, pi1006, pi1007,
    pi1008, pi1009, pi1010, pi1011, pi1012, pi1013, pi1014, pi1015, pi1016,
    pi1017, pi1018, pi1019, pi1020, pi1021, pi1022, pi1023, pi1024, pi1025,
    pi1026, pi1027, pi1028, pi1029, pi1030, pi1031, pi1032, pi1033, pi1034,
    pi1035, pi1036, pi1037, pi1038, pi1039, pi1040, pi1041, pi1042, pi1043,
    pi1044, pi1045, pi1046, pi1047, pi1048, pi1049, pi1050, pi1051, pi1052,
    pi1053, pi1054, pi1055, pi1056, pi1057, pi1058, pi1059, pi1060, pi1061,
    pi1062, pi1063, pi1064, pi1065, pi1066, pi1067, pi1068, pi1069, pi1070,
    pi1071, pi1072, pi1073, pi1074, pi1075, pi1076, pi1077, pi1078, pi1079,
    pi1080, pi1081, pi1082, pi1083, pi1084, pi1085, pi1086, pi1087, pi1088,
    pi1089, pi1090, pi1091, pi1092, pi1093, pi1094, pi1095, pi1096, pi1097,
    pi1098, pi1099, pi1100, pi1101, pi1102, pi1103, pi1104, pi1105, pi1106,
    pi1107, pi1108, pi1109, pi1110, pi1111, pi1112, pi1113, pi1114, pi1115,
    pi1116, pi1117, pi1118, pi1119, pi1120, pi1121, pi1122, pi1123, pi1124,
    pi1125, pi1126, pi1127, pi1128, pi1129, pi1130, pi1131, pi1132, pi1133,
    pi1134, pi1135, pi1136, pi1137, pi1138, pi1139, pi1140, pi1141, pi1142,
    pi1143, pi1144, pi1145, pi1146, pi1147, pi1148, pi1149, pi1150, pi1151,
    pi1152, pi1153, pi1154, pi1155, pi1156, pi1157, pi1158, pi1159, pi1160,
    pi1161, pi1162, pi1163, pi1164, pi1165, pi1166, pi1167, pi1168, pi1169,
    pi1170, pi1171, pi1172, pi1173, pi1174, pi1175, pi1176, pi1177, pi1178,
    pi1179, pi1180, pi1181, pi1182, pi1183, pi1184, pi1185, pi1186, pi1187,
    pi1188, pi1189, pi1190, pi1191, pi1192, pi1193, pi1194, pi1195, pi1196,
    pi1197, pi1198, pi1199, pi1200, pi1201, pi1202, pi1203, pi1204, pi1205,
    pi1206, pi1207, pi1208, pi1209, pi1210, pi1211, pi1212, pi1213, pi1214,
    pi1215, pi1216, pi1217, pi1218, pi1219, pi1220, pi1221, pi1222, pi1223,
    pi1224, pi1225, pi1226, pi1227, pi1228, pi1229, pi1230, pi1231, pi1232,
    pi1233, pi1234, pi1235, pi1236, pi1237, pi1238, pi1239, pi1240, pi1241,
    pi1242, pi1243, pi1244, pi1245, pi1246, pi1247, pi1248, pi1249, pi1250,
    pi1251, pi1252, pi1253, pi1254, pi1255, pi1256, pi1257, pi1258, pi1259,
    pi1260, pi1261, pi1262, pi1263, pi1264, pi1265, pi1266, pi1267, pi1268,
    pi1269, pi1270, pi1271, pi1272, pi1273, pi1274, pi1275, pi1276, pi1277,
    pi1278, pi1279, pi1280, pi1281, pi1282, pi1283, pi1284, pi1285, pi1286,
    pi1287, pi1288, pi1289, pi1290, pi1291, pi1292, pi1293, pi1294, pi1295,
    pi1296, pi1297, pi1298, pi1299, pi1300, pi1301, pi1302, pi1303, pi1304,
    pi1305, pi1306, pi1307, pi1308, pi1309, pi1310, pi1311, pi1312, pi1313,
    pi1314, pi1315, pi1316, pi1317, pi1318, pi1319, pi1320, pi1321, pi1322,
    pi1323, pi1324, pi1325, pi1326, pi1327, pi1328, pi1329, pi1330, pi1331,
    pi1332, pi1333, pi1334, pi1335, pi1336, pi1337, pi1338, pi1339, pi1340,
    pi1341, pi1342, pi1343, pi1344, pi1345, pi1346, pi1347, pi1348, pi1349,
    pi1350, pi1351, pi1352, pi1353, pi1354, pi1355, pi1356, pi1357, pi1358,
    pi1359, pi1360, pi1361, pi1362, pi1363, pi1364, pi1365, pi1366, pi1367,
    pi1368, pi1369, pi1370, pi1371, pi1372, pi1373, pi1374, pi1375, pi1376,
    pi1377, pi1378, pi1379, pi1380, pi1381, pi1382, pi1383, pi1384, pi1385,
    pi1386, pi1387, pi1388, pi1389, pi1390, pi1391, pi1392, pi1393, pi1394,
    pi1395, pi1396, pi1397, pi1398, pi1399, pi1400, pi1401, pi1402, pi1403,
    pi1404, pi1405, pi1406, pi1407, pi1408, pi1409, pi1410, pi1411, pi1412,
    pi1413, pi1414, pi1415, pi1416, pi1417, pi1418, pi1419, pi1420, pi1421,
    pi1422, pi1423, pi1424, pi1425, pi1426, pi1427, pi1428, pi1429, pi1430,
    pi1431, pi1432, pi1433, pi1434, pi1435, pi1436, pi1437, pi1438, pi1439,
    pi1440, pi1441, pi1442, pi1443, pi1444, pi1445, pi1446, pi1447, pi1448,
    pi1449, pi1450, pi1451, pi1452, pi1453, pi1454, pi1455, pi1456, pi1457,
    pi1458, pi1459, pi1460, pi1461, pi1462, pi1463, pi1464, pi1465, pi1466,
    pi1467, pi1468, pi1469, pi1470, pi1471, pi1472, pi1473, pi1474, pi1475,
    pi1476, pi1477, pi1478, pi1479, pi1480, pi1481, pi1482, pi1483, pi1484,
    pi1485, pi1486, pi1487, pi1488, pi1489, pi1490, pi1491, pi1492, pi1493,
    pi1494, pi1495, pi1496, pi1497, pi1498, pi1499, pi1500, pi1501, pi1502,
    pi1503, pi1504, pi1505, pi1506, pi1507, pi1508, pi1509, pi1510, pi1511,
    pi1512, pi1513, pi1514, pi1515, pi1516, pi1517, pi1518, pi1519, pi1520,
    pi1521, pi1522, pi1523, pi1524, pi1525, pi1526, pi1527, pi1528, pi1529,
    pi1530, pi1531, pi1532, pi1533, pi1534, pi1535, pi1536, pi1537, pi1538,
    pi1539, pi1540, pi1541, pi1542, pi1543, pi1544, pi1545, pi1546, pi1547,
    pi1548, pi1549, pi1550, pi1551, pi1552, pi1553, pi1554, pi1555, pi1556,
    pi1557, pi1558, pi1559, pi1560, pi1561, pi1562, pi1563, pi1564, pi1565,
    pi1566, pi1567, pi1568, pi1569, pi1570, pi1571, pi1572, pi1573, pi1574,
    pi1575, pi1576, pi1577, pi1578, pi1579, pi1580, pi1581, pi1582, pi1583,
    pi1584, pi1585, pi1586, pi1587, pi1588, pi1589, pi1590, pi1591, pi1592,
    pi1593, pi1594, pi1595, pi1596, pi1597, pi1598, pi1599, pi1600, pi1601,
    pi1602, pi1603, pi1604, pi1605, pi1606, pi1607, pi1608, pi1609, pi1610,
    pi1611, pi1612, pi1613, pi1614, pi1615, pi1616, pi1617, pi1618, pi1619,
    pi1620, pi1621, pi1622, pi1623, pi1624, pi1625, pi1626, pi1627, pi1628,
    pi1629, pi1630, pi1631, pi1632, pi1633, pi1634, pi1635, pi1636, pi1637,
    pi1638, pi1639, pi1640, pi1641, pi1642, pi1643, pi1644, pi1645, pi1646,
    pi1647, pi1648, pi1649, pi1650, pi1651, pi1652, pi1653, pi1654, pi1655,
    pi1656, pi1657, pi1658, pi1659, pi1660, pi1661, pi1662, pi1663, pi1664,
    pi1665, pi1666, pi1667, pi1668, pi1669, pi1670, pi1671, pi1672, pi1673,
    pi1674, pi1675, pi1676, pi1677, pi1678, pi1679, pi1680, pi1681, pi1682,
    pi1683, pi1684, pi1685, pi1686, pi1687, pi1688, pi1689, pi1690, pi1691,
    pi1692, pi1693, pi1694, pi1695, pi1696, pi1697, pi1698, pi1699, pi1700,
    pi1701, pi1702, pi1703, pi1704, pi1705, pi1706, pi1707, pi1708, pi1709,
    pi1710, pi1711, pi1712, pi1713, pi1714, pi1715, pi1716, pi1717, pi1718,
    pi1719, pi1720, pi1721, pi1722, pi1723, pi1724, pi1725, pi1726, pi1727,
    pi1728, pi1729, pi1730, pi1731, pi1732, pi1733, pi1734, pi1735, pi1736,
    pi1737, pi1738, pi1739, pi1740, pi1741, pi1742, pi1743, pi1744, pi1745,
    pi1746, pi1747, pi1748, pi1749, pi1750, pi1751, pi1752, pi1753, pi1754,
    pi1755, pi1756, pi1757, pi1758, pi1759, pi1760, pi1761, pi1762, pi1763,
    pi1764, pi1765, pi1766, pi1767, pi1768, pi1769, pi1770, pi1771, pi1772,
    pi1773, pi1774, pi1775, pi1776, pi1777, pi1778, pi1779, pi1780, pi1781,
    pi1782, pi1783, pi1784, pi1785, pi1786, pi1787, pi1788, pi1789, pi1790,
    pi1791, pi1792, pi1793, pi1794, pi1795, pi1796, pi1797, pi1798, pi1799,
    pi1800, pi1801, pi1802, pi1803, pi1804, pi1805, pi1806, pi1807, pi1808,
    pi1809, pi1810, pi1811, pi1812, pi1813, pi1814, pi1815, pi1816, pi1817,
    pi1818, pi1819, pi1820, pi1821, pi1822, pi1823, pi1824, pi1825, pi1826,
    pi1827, pi1828, pi1829, pi1830, pi1831, pi1832, pi1833, pi1834, pi1835,
    pi1836, pi1837, pi1838, pi1839, pi1840, pi1841, pi1842, pi1843, pi1844,
    pi1845, pi1846, pi1847, pi1848, pi1849, pi1850, pi1851, pi1852, pi1853,
    pi1854, pi1855, pi1856, pi1857, pi1858, pi1859, pi1860, pi1861, pi1862,
    pi1863, pi1864, pi1865, pi1866, pi1867, pi1868, pi1869, pi1870, pi1871,
    pi1872, pi1873, pi1874, pi1875, pi1876, pi1877, pi1878, pi1879, pi1880,
    pi1881, pi1882, pi1883, pi1884, pi1885, pi1886, pi1887, pi1888, pi1889,
    pi1890, pi1891, pi1892, pi1893, pi1894, pi1895, pi1896, pi1897, pi1898,
    pi1899, pi1900, pi1901, pi1902, pi1903, pi1904, pi1905, pi1906, pi1907,
    pi1908, pi1909, pi1910, pi1911, pi1912, pi1913, pi1914, pi1915, pi1916,
    pi1917, pi1918, pi1919, pi1920, pi1921, pi1922, pi1923, pi1924, pi1925,
    pi1926, pi1927, pi1928, pi1929, pi1930, pi1931, pi1932, pi1933, pi1934,
    pi1935, pi1936, pi1937, pi1938, pi1939, pi1940, pi1941, pi1942, pi1943,
    pi1944, pi1945, pi1946, pi1947, pi1948, pi1949, pi1950, pi1951, pi1952,
    pi1953, pi1954, pi1955, pi1956, pi1957, pi1958, pi1959, pi1960, pi1961,
    pi1962, pi1963, pi1964, pi1965, pi1966, pi1967, pi1968, pi1969, pi1970,
    pi1971, pi1972, pi1973, pi1974, pi1975, pi1976, pi1977, pi1978, pi1979,
    pi1980, pi1981, pi1982, pi1983, pi1984, pi1985, pi1986, pi1987, pi1988,
    pi1989, pi1990, pi1991, pi1992, pi1993, pi1994, pi1995, pi1996, pi1997,
    pi1998, pi1999, pi2000, pi2001, pi2002, pi2003, pi2004, pi2005, pi2006,
    pi2007, pi2008, pi2009, pi2010, pi2011, pi2012, pi2013, pi2014, pi2015,
    pi2016, pi2017, pi2018, pi2019, pi2020, pi2021, pi2022, pi2023, pi2024,
    pi2025, pi2026, pi2027, pi2028, pi2029, pi2030, pi2031, pi2032, pi2033,
    pi2034, pi2035, pi2036, pi2037, pi2038, pi2039, pi2040, pi2041, pi2042,
    pi2043, pi2044, pi2045, pi2046, pi2047, pi2048, pi2049, pi2050, pi2051,
    pi2052, pi2053, pi2054, pi2055, pi2056, pi2057, pi2058, pi2059, pi2060,
    pi2061, pi2062, pi2063, pi2064, pi2065, pi2066, pi2067, pi2068, pi2069,
    pi2070, pi2071, pi2072, pi2073, pi2074, pi2075, pi2076, pi2077, pi2078,
    pi2079, pi2080, pi2081, pi2082, pi2083, pi2084, pi2085, pi2086, pi2087,
    pi2088, pi2089, pi2090, pi2091, pi2092, pi2093, pi2094, pi2095, pi2096,
    pi2097, pi2098, pi2099, pi2100, pi2101, pi2102, pi2103, pi2104, pi2105,
    pi2106, pi2107, pi2108, pi2109, pi2110, pi2111, pi2112, pi2113, pi2114,
    pi2115, pi2116, pi2117, pi2118, pi2119, pi2120, pi2121, pi2122, pi2123,
    pi2124, pi2125, pi2126, pi2127, pi2128, pi2129, pi2130, pi2131, pi2132,
    pi2133, pi2134, pi2135, pi2136, pi2137, pi2138, pi2139, pi2140, pi2141,
    pi2142, pi2143, pi2144, pi2145, pi2146, pi2147, pi2148, pi2149, pi2150,
    pi2151, pi2152, pi2153, pi2154, pi2155, pi2156, pi2157, pi2158, pi2159,
    pi2160, pi2161, pi2162, pi2163, pi2164, pi2165, pi2166, pi2167, pi2168,
    pi2169, pi2170, pi2171, pi2172, pi2173, pi2174, pi2175, pi2176, pi2177,
    pi2178, pi2179, pi2180, pi2181, pi2182, pi2183, pi2184, pi2185, pi2186,
    pi2187, pi2188, pi2189, pi2190, pi2191, pi2192, pi2193, pi2194, pi2195,
    pi2196, pi2197, pi2198, pi2199, pi2200, pi2201, pi2202, pi2203, pi2204,
    pi2205, pi2206, pi2207, pi2208, pi2209, pi2210, pi2211, pi2212, pi2213,
    pi2214, pi2215, pi2216, pi2217, pi2218, pi2219, pi2220, pi2221, pi2222,
    pi2223, pi2224, pi2225, pi2226, pi2227, pi2228, pi2229, pi2230, pi2231,
    pi2232, pi2233, pi2234, pi2235, pi2236, pi2237, pi2238, pi2239, pi2240,
    pi2241, pi2242, pi2243, pi2244, pi2245, pi2246, pi2247, pi2248, pi2249,
    pi2250, pi2251, pi2252, pi2253, pi2254, pi2255, pi2256, pi2257, pi2258,
    pi2259, pi2260, pi2261, pi2262, pi2263, pi2264, pi2265, pi2266, pi2267,
    pi2268, pi2269, pi2270, pi2271, pi2272, pi2273, pi2274, pi2275, pi2276,
    pi2277, pi2278, pi2279, pi2280, pi2281, pi2282, pi2283, pi2284, pi2285,
    pi2286, pi2287, pi2288, pi2289, pi2290, pi2291, pi2292, pi2293, pi2294,
    pi2295, pi2296, pi2297, pi2298, pi2299, pi2300, pi2301, pi2302, pi2303,
    pi2304, pi2305, pi2306, pi2307, pi2308, pi2309, pi2310, pi2311, pi2312,
    pi2313, pi2314, pi2315, pi2316, pi2317, pi2318, pi2319, pi2320, pi2321,
    pi2322, pi2323, pi2324, pi2325, pi2326, pi2327, pi2328, pi2329, pi2330,
    pi2331, pi2332, pi2333, pi2334, pi2335, pi2336, pi2337, pi2338, pi2339,
    pi2340, pi2341, pi2342, pi2343, pi2344, pi2345, pi2346, pi2347, pi2348,
    pi2349, pi2350, pi2351, pi2352, pi2353, pi2354, pi2355, pi2356, pi2357,
    pi2358, pi2359, pi2360, pi2361, pi2362, pi2363, pi2364, pi2365, pi2366,
    pi2367, pi2368, pi2369, pi2370, pi2371, pi2372, pi2373, pi2374, pi2375,
    pi2376, pi2377, pi2378, pi2379, pi2380, pi2381, pi2382, pi2383, pi2384,
    pi2385, pi2386, pi2387, pi2388, pi2389, pi2390, pi2391, pi2392, pi2393,
    pi2394, pi2395, pi2396, pi2397, pi2398, pi2399, pi2400, pi2401, pi2402,
    pi2403, pi2404, pi2405, pi2406, pi2407, pi2408, pi2409, pi2410, pi2411,
    pi2412, pi2413, pi2414, pi2415, pi2416, pi2417, pi2418, pi2419, pi2420,
    pi2421, pi2422, pi2423, pi2424, pi2425, pi2426, pi2427, pi2428, pi2429,
    pi2430, pi2431, pi2432, pi2433, pi2434, pi2435, pi2436, pi2437, pi2438,
    pi2439, pi2440, pi2441, pi2442, pi2443, pi2444, pi2445, pi2446, pi2447,
    pi2448, pi2449, pi2450, pi2451, pi2452, pi2453, pi2454, pi2455, pi2456,
    pi2457, pi2458, pi2459, pi2460, pi2461, pi2462, pi2463, pi2464, pi2465,
    pi2466, pi2467, pi2468, pi2469, pi2470, pi2471, pi2472, pi2473, pi2474,
    pi2475, pi2476, pi2477, pi2478, pi2479, pi2480, pi2481, pi2482, pi2483,
    pi2484, pi2485, pi2486, pi2487, pi2488, pi2489, pi2490, pi2491, pi2492,
    pi2493, pi2494, pi2495, pi2496, pi2497, pi2498, pi2499, pi2500, pi2501,
    pi2502, pi2503, pi2504, pi2505, pi2506, pi2507, pi2508, pi2509, pi2510,
    pi2511, pi2512, pi2513, pi2514, pi2515, pi2516, pi2517, pi2518, pi2519,
    pi2520, pi2521, pi2522, pi2523, pi2524, pi2525, pi2526, pi2527, pi2528,
    pi2529, pi2530, pi2531, pi2532, pi2533, pi2534, pi2535, pi2536, pi2537,
    pi2538, pi2539, pi2540, pi2541, pi2542, pi2543, pi2544, pi2545, pi2546,
    pi2547, pi2548, pi2549, pi2550, pi2551, pi2552, pi2553, pi2554, pi2555,
    pi2556, pi2557, pi2558, pi2559, pi2560, pi2561, pi2562, pi2563, pi2564,
    pi2565, pi2566, pi2567, pi2568, pi2569, pi2570, pi2571, pi2572, pi2573,
    pi2574, pi2575, pi2576, pi2577, pi2578, pi2579, pi2580, pi2581, pi2582,
    pi2583, pi2584, pi2585, pi2586, pi2587, pi2588, pi2589, pi2590, pi2591,
    pi2592, pi2593, pi2594, pi2595, pi2596, pi2597, pi2598, pi2599, pi2600,
    pi2601, pi2602, pi2603, pi2604, pi2605, pi2606, pi2607, pi2608, pi2609,
    pi2610, pi2611, pi2612, pi2613, pi2614, pi2615, pi2616, pi2617, pi2618,
    pi2619, pi2620, pi2621, pi2622, pi2623, pi2624, pi2625, pi2626, pi2627,
    pi2628, pi2629, pi2630, pi2631, pi2632, pi2633, pi2634, pi2635, pi2636,
    pi2637, pi2638, pi2639, pi2640, pi2641, pi2642, pi2643, pi2644, pi2645,
    pi2646, pi2647, pi2648, pi2649, pi2650, pi2651, pi2652, pi2653, pi2654,
    pi2655, pi2656, pi2657, pi2658, pi2659, pi2660, pi2661, pi2662, pi2663,
    pi2664, pi2665, pi2666, pi2667, pi2668, pi2669, pi2670, pi2671, pi2672,
    pi2673, pi2674, pi2675, pi2676, pi2677, pi2678, pi2679, pi2680, pi2681,
    pi2682, pi2683, pi2684, pi2685, pi2686, pi2687, pi2688, pi2689, pi2690,
    pi2691, pi2692, pi2693, pi2694, pi2695, pi2696, pi2697, pi2698, pi2699,
    pi2700, pi2701, pi2702, pi2703, pi2704, pi2705, pi2706, pi2707, pi2708,
    pi2709, pi2710, pi2711, pi2712, pi2713, pi2714, pi2715, pi2716, pi2717,
    pi2718, pi2719, pi2720, pi2721, pi2722, pi2723, pi2724, pi2725, pi2726,
    pi2727, pi2728, pi2729, pi2730, pi2731, pi2732, pi2733, pi2734, pi2735,
    pi2736, pi2737, pi2738, pi2739, pi2740, pi2741, pi2742, pi2743, pi2744,
    pi2745, pi2746, pi2747, pi2748, pi2749, pi2750, pi2751, pi2752, pi2753,
    pi2754, pi2755, pi2756, pi2757, pi2758, pi2759, pi2760, pi2761, pi2762,
    pi2763, pi2764, pi2765, pi2766, pi2767, pi2768, pi2769, pi2770, pi2771,
    pi2772, pi2773, pi2774, pi2775, pi2776, pi2777, pi2778, pi2779, pi2780,
    pi2781, pi2782, pi2783, pi2784, pi2785, pi2786, pi2787, pi2788, pi2789,
    pi2790, pi2791, pi2792, pi2793, pi2794, pi2795, pi2796, pi2797, pi2798,
    pi2799, pi2800, pi2801, pi2802, pi2803, pi2804, pi2805, pi2806, pi2807,
    pi2808, pi2809, pi2810, pi2811, pi2812, pi2813, pi2814, pi2815, pi2816,
    pi2817, pi2818, pi2819, pi2820, pi2821, pi2822, pi2823, pi2824, pi2825,
    pi2826, pi2827, pi2828, pi2829, pi2830, pi2831, pi2832, pi2833, pi2834,
    pi2835, pi2836, pi2837, pi2838, pi2839, pi2840, pi2841, pi2842, pi2843,
    pi2844, pi2845, pi2846, pi2847, pi2848, pi2849, pi2850, pi2851, pi2852,
    pi2853, pi2854, pi2855, pi2856, pi2857, pi2858, pi2859, pi2860, pi2861,
    pi2862, pi2863, pi2864, pi2865, pi2866, pi2867, pi2868, pi2869, pi2870,
    pi2871, pi2872, pi2873, pi2874, pi2875, pi2876, pi2877, pi2878, pi2879,
    pi2880, pi2881, pi2882, pi2883, pi2884, pi2885, pi2886, pi2887, pi2888,
    pi2889, pi2890, pi2891, pi2892, pi2893, pi2894, pi2895, pi2896, pi2897,
    pi2898, pi2899, pi2900, pi2901, pi2902, pi2903, pi2904, pi2905, pi2906,
    pi2907, pi2908, pi2909, pi2910, pi2911, pi2912, pi2913, pi2914, pi2915,
    pi2916, pi2917, pi2918, pi2919, pi2920, pi2921, pi2922, pi2923, pi2924,
    pi2925, pi2926, pi2927, pi2928, pi2929, pi2930, pi2931, pi2932, pi2933,
    pi2934, pi2935, pi2936, pi2937, pi2938, pi2939, pi2940, pi2941, pi2942,
    pi2943, pi2944, pi2945, pi2946, pi2947, pi2948, pi2949, pi2950, pi2951,
    pi2952, pi2953, pi2954, pi2955, pi2956, pi2957, pi2958, pi2959, pi2960,
    pi2961, pi2962, pi2963, pi2964, pi2965, pi2966, pi2967, pi2968, pi2969,
    pi2970, pi2971, pi2972, pi2973, pi2974, pi2975, pi2976, pi2977, pi2978,
    pi2979, pi2980, pi2981, pi2982, pi2983, pi2984, pi2985, pi2986, pi2987,
    pi2988, pi2989, pi2990, pi2991, pi2992, pi2993, pi2994, pi2995, pi2996,
    pi2997, pi2998, pi2999, pi3000, pi3001, pi3002, pi3003, pi3004, pi3005,
    pi3006, pi3007, pi3008, pi3009, pi3010, pi3011, pi3012, pi3013, pi3014,
    pi3015, pi3016, pi3017, pi3018, pi3019, pi3020, pi3021, pi3022, pi3023,
    pi3024, pi3025, pi3026, pi3027, pi3028, pi3029, pi3030, pi3031, pi3032,
    pi3033, pi3034, pi3035, pi3036, pi3037, pi3038, pi3039, pi3040, pi3041,
    pi3042, pi3043, pi3044, pi3045, pi3046, pi3047, pi3048, pi3049, pi3050,
    pi3051, pi3052, pi3053, pi3054, pi3055, pi3056, pi3057, pi3058, pi3059,
    pi3060, pi3061, pi3062, pi3063, pi3064, pi3065, pi3066, pi3067, pi3068,
    pi3069, pi3070, pi3071, pi3072, pi3073, pi3074, pi3075, pi3076, pi3077,
    pi3078, pi3079, pi3080, pi3081, pi3082, pi3083, pi3084, pi3085, pi3086,
    pi3087, pi3088, pi3089, pi3090, pi3091, pi3092, pi3093, pi3094, pi3095,
    pi3096, pi3097, pi3098, pi3099, pi3100, pi3101, pi3102, pi3103, pi3104,
    pi3105, pi3106, pi3107, pi3108, pi3109, pi3110, pi3111, pi3112, pi3113,
    pi3114, pi3115, pi3116, pi3117, pi3118, pi3119, pi3120, pi3121, pi3122,
    pi3123, pi3124, pi3125, pi3126, pi3127, pi3128, pi3129, pi3130, pi3131,
    pi3132, pi3133, pi3134, pi3135, pi3136, pi3137, pi3138, pi3139, pi3140,
    pi3141, pi3142, pi3143, pi3144, pi3145, pi3146, pi3147, pi3148, pi3149,
    pi3150, pi3151, pi3152, pi3153, pi3154, pi3155, pi3156, pi3157, pi3158,
    pi3159, pi3160, pi3161, pi3162, pi3163, pi3164, pi3165, pi3166, pi3167,
    pi3168, pi3169, pi3170, pi3171, pi3172, pi3173, pi3174, pi3175, pi3176,
    pi3177, pi3178, pi3179, pi3180, pi3181, pi3182, pi3183, pi3184, pi3185,
    pi3186, pi3187, pi3188, pi3189, pi3190, pi3191, pi3192, pi3193, pi3194,
    pi3195, pi3196, pi3197, pi3198, pi3199, pi3200, pi3201, pi3202, pi3203,
    pi3204, pi3205, pi3206, pi3207, pi3208, pi3209, pi3210, pi3211, pi3212,
    pi3213, pi3214, pi3215, pi3216, pi3217, pi3218, pi3219, pi3220, pi3221,
    pi3222, pi3223, pi3224, pi3225, pi3226, pi3227, pi3228, pi3229, pi3230,
    pi3231, pi3232, pi3233, pi3234, pi3235, pi3236, pi3237, pi3238, pi3239,
    pi3240, pi3241, pi3242, pi3243, pi3244, pi3245, pi3246, pi3247, pi3248,
    pi3249, pi3250, pi3251, pi3252, pi3253, pi3254, pi3255, pi3256, pi3257,
    pi3258, pi3259, pi3260, pi3261, pi3262, pi3263, pi3264, pi3265, pi3266,
    pi3267, pi3268, pi3269, pi3270, pi3271, pi3272, pi3273, pi3274, pi3275,
    pi3276, pi3277, pi3278, pi3279, pi3280, pi3281, pi3282, pi3283, pi3284,
    pi3285, pi3286, pi3287, pi3288, pi3289, pi3290, pi3291, pi3292, pi3293,
    pi3294, pi3295, pi3296, pi3297, pi3298, pi3299, pi3300, pi3301, pi3302,
    pi3303, pi3304, pi3305, pi3306, pi3307, pi3308, pi3309, pi3310, pi3311,
    pi3312, pi3313, pi3314, pi3315, pi3316, pi3317, pi3318, pi3319, pi3320,
    pi3321, pi3322, pi3323, pi3324, pi3325, pi3326, pi3327, pi3328, pi3329,
    pi3330, pi3331, pi3332, pi3333, pi3334, pi3335, pi3336, pi3337, pi3338,
    pi3339, pi3340, pi3341, pi3342, pi3343, pi3344, pi3345, pi3346, pi3347,
    pi3348, pi3349, pi3350, pi3351, pi3352, pi3353, pi3354, pi3355, pi3356,
    pi3357, pi3358, pi3359, pi3360, pi3361, pi3362, pi3363, pi3364, pi3365,
    pi3366, pi3367, pi3368, pi3369, pi3370, pi3371, pi3372, pi3373, pi3374,
    pi3375, pi3376, pi3377, pi3378, pi3379, pi3380, pi3381, pi3382, pi3383,
    pi3384, pi3385, pi3386, pi3387, pi3388, pi3389, pi3390, pi3391, pi3392,
    pi3393, pi3394, pi3395, pi3396, pi3397, pi3398, pi3399, pi3400, pi3401,
    pi3402, pi3403, pi3404, pi3405, pi3406, pi3407, pi3408, pi3409, pi3410,
    pi3411, pi3412, pi3413, pi3414, pi3415, pi3416, pi3417, pi3418, pi3419,
    pi3420, pi3421, pi3422, pi3423, pi3424, pi3425, pi3426, pi3427, pi3428,
    pi3429, pi3430, pi3431, pi3432, pi3433, pi3434, pi3435, pi3436, pi3437,
    pi3438, pi3439, pi3440, pi3441, pi3442, pi3443, pi3444, pi3445, pi3446,
    pi3447, pi3448, pi3449, pi3450, pi3451, pi3452, pi3453, pi3454, pi3455,
    pi3456, pi3457, pi3458, pi3459, pi3460, pi3461, pi3462, pi3463, pi3464,
    pi3465, pi3466, pi3467, pi3468, pi3469, pi3470, pi3471, pi3472, pi3473,
    pi3474, pi3475, pi3476, pi3477, pi3478, pi3479, pi3480, pi3481, pi3482,
    pi3483, pi3484, pi3485, pi3486, pi3487, pi3488, pi3489, pi3490, pi3491,
    pi3492, pi3493, pi3494, pi3495, pi3496, pi3497, pi3498, pi3499, pi3500,
    pi3501, pi3502, pi3503, pi3504, pi3505, pi3506, pi3507, pi3508, pi3509,
    pi3510, pi3511, pi3512, pi3513, pi3514, pi3515, pi3516, pi3517, pi3518,
    pi3519, pi3520, pi3521, pi3522, pi3523, pi3524, pi3525, pi3526, pi3527,
    pi3528, pi3529, pi3530, pi3531, pi3532, pi3533, pi3534, pi3535, pi3536,
    pi3537, pi3538, pi3539, pi3540, pi3541, pi3542, pi3543, pi3544, pi3545,
    pi3546, pi3547, pi3548, pi3549, pi3550, pi3551, pi3552, pi3553, pi3554,
    pi3555, pi3556, pi3557, pi3558, pi3559, pi3560, pi3561, pi3562, pi3563,
    pi3564, pi3565, pi3566, pi3567, pi3568, pi3569, pi3570, pi3571, pi3572,
    pi3573, pi3574, pi3575, pi3576, pi3577, pi3578, pi3579, pi3580, pi3581,
    pi3582, pi3583, pi3584, pi3585, pi3586, pi3587, pi3588, pi3589, pi3590,
    pi3591, pi3592, pi3593, pi3594, pi3595, pi3596, pi3597, pi3598, pi3599,
    pi3600, pi3601, pi3602, pi3603, pi3604, pi3605, pi3606, pi3607, pi3608,
    pi3609, pi3610, pi3611, pi3612, pi3613, pi3614, pi3615, pi3616, pi3617,
    pi3618, pi3619, pi3620, pi3621, pi3622, pi3623, pi3624, pi3625, pi3626,
    pi3627, pi3628, pi3629, pi3630, pi3631, pi3632, pi3633, pi3634, pi3635,
    pi3636, pi3637, pi3638, pi3639, pi3640, pi3641, pi3642, pi3643, pi3644,
    pi3645, pi3646, pi3647, pi3648, pi3649, pi3650, pi3651, pi3652, pi3653,
    pi3654, pi3655, pi3656, pi3657, pi3658, pi3659, pi3660, pi3661, pi3662,
    pi3663, pi3664, pi3665, pi3666, pi3667, pi3668, pi3669, pi3670, pi3671,
    pi3672, pi3673, pi3674, pi3675, pi3676, pi3677, pi3678, pi3679, pi3680,
    pi3681, pi3682, pi3683, pi3684, pi3685, pi3686, pi3687, pi3688, pi3689,
    pi3690, pi3691, pi3692, pi3693, pi3694, pi3695, pi3696, pi3697, pi3698,
    pi3699, pi3700, pi3701, pi3702, pi3703, pi3704, pi3705, pi3706, pi3707,
    pi3708, pi3709, pi3710, pi3711, pi3712, pi3713, pi3714, pi3715, pi3716,
    pi3717, pi3718, pi3719, pi3720, pi3721, pi3722, pi3723, pi3724, pi3725,
    pi3726, pi3727, pi3728, pi3729, pi3730, pi3731, pi3732, pi3733, pi3734,
    pi3735, pi3736, pi3737, pi3738, pi3739, pi3740, pi3741, pi3742, pi3743,
    pi3744, pi3745, pi3746, pi3747, pi3748, pi3749, pi3750, pi3751, pi3752,
    pi3753, pi3754, pi3755, pi3756, pi3757, pi3758, pi3759, pi3760, pi3761,
    pi3762, pi3763, pi3764, pi3765, pi3766, pi3767, pi3768, pi3769, pi3770,
    pi3771, pi3772, pi3773, pi3774, pi3775, pi3776, pi3777, pi3778, pi3779,
    pi3780, pi3781, pi3782, pi3783, pi3784, pi3785, pi3786, pi3787, pi3788,
    pi3789, pi3790, pi3791, pi3792, pi3793, pi3794, pi3795, pi3796, pi3797,
    pi3798, pi3799, pi3800, pi3801, pi3802, pi3803, pi3804, pi3805, pi3806,
    pi3807, pi3808, pi3809, pi3810, pi3811, pi3812, pi3813, pi3814, pi3815,
    pi3816, pi3817, pi3818, pi3819, pi3820, pi3821, pi3822, pi3823, pi3824,
    pi3825, pi3826, pi3827, pi3828, pi3829, pi3830, pi3831, pi3832, pi3833,
    pi3834, pi3835, pi3836, pi3837, pi3838, pi3839, pi3840, pi3841, pi3842,
    pi3843, pi3844, pi3845, pi3846, pi3847, pi3848, pi3849, pi3850, pi3851,
    pi3852, pi3853, pi3854, pi3855, pi3856, pi3857, pi3858, pi3859, pi3860,
    pi3861, pi3862, pi3863, pi3864, pi3865, pi3866, pi3867, pi3868, pi3869,
    pi3870, pi3871, pi3872, pi3873, pi3874, pi3875, pi3876, pi3877, pi3878,
    pi3879, pi3880, pi3881, pi3882, pi3883, pi3884, pi3885, pi3886, pi3887,
    pi3888, pi3889, pi3890, pi3891, pi3892, pi3893, pi3894, pi3895, pi3896,
    pi3897, pi3898, pi3899, pi3900, pi3901, pi3902, pi3903, pi3904, pi3905,
    pi3906, pi3907, pi3908, pi3909, pi3910, pi3911, pi3912, pi3913, pi3914,
    pi3915, pi3916, pi3917, pi3918, pi3919, pi3920, pi3921, pi3922, pi3923,
    pi3924, pi3925, pi3926, pi3927, pi3928, pi3929, pi3930, pi3931, pi3932,
    pi3933, pi3934, pi3935, pi3936, pi3937, pi3938, pi3939, pi3940, pi3941,
    pi3942, pi3943, pi3944, pi3945, pi3946, pi3947, pi3948, pi3949, pi3950,
    pi3951, pi3952, pi3953, pi3954, pi3955, pi3956, pi3957, pi3958, pi3959,
    pi3960, pi3961, pi3962, pi3963, pi3964, pi3965, pi3966, pi3967, pi3968,
    pi3969, pi3970, pi3971, pi3972, pi3973, pi3974, pi3975, pi3976, pi3977,
    pi3978, pi3979, pi3980, pi3981, pi3982, pi3983, pi3984, pi3985, pi3986,
    pi3987, pi3988, pi3989, pi3990, pi3991, pi3992, pi3993, pi3994, pi3995,
    pi3996, pi3997, pi3998, pi3999, pi4000, pi4001, pi4002, pi4003, pi4004,
    pi4005, pi4006, pi4007, pi4008, pi4009, pi4010, pi4011, pi4012, pi4013,
    pi4014, pi4015, pi4016, pi4017, pi4018, pi4019, pi4020, pi4021, pi4022,
    pi4023, pi4024, pi4025, pi4026, pi4027, pi4028, pi4029, pi4030, pi4031,
    pi4032, pi4033, pi4034, pi4035, pi4036, pi4037, pi4038, pi4039, pi4040,
    pi4041, pi4042, pi4043, pi4044, pi4045, pi4046, pi4047, pi4048, pi4049,
    pi4050, pi4051, pi4052, pi4053, pi4054, pi4055, pi4056, pi4057, pi4058,
    pi4059, pi4060, pi4061, pi4062, pi4063, pi4064, pi4065, pi4066, pi4067,
    pi4068, pi4069, pi4070, pi4071, pi4072, pi4073, pi4074, pi4075, pi4076,
    pi4077, pi4078, pi4079, pi4080, pi4081, pi4082, pi4083, pi4084, pi4085,
    pi4086, pi4087, pi4088, pi4089, pi4090, pi4091, pi4092, pi4093, pi4094,
    pi4095, pi4096, pi4097, pi4098, pi4099, pi4100, pi4101, pi4102, pi4103,
    pi4104, pi4105, pi4106, pi4107, pi4108, pi4109, pi4110, pi4111, pi4112,
    pi4113, pi4114, pi4115, pi4116, pi4117, pi4118, pi4119, pi4120, pi4121,
    pi4122, pi4123, pi4124, pi4125, pi4126, pi4127, pi4128, pi4129, pi4130,
    pi4131, pi4132, pi4133, pi4134, pi4135, pi4136, pi4137, pi4138, pi4139,
    pi4140, pi4141, pi4142, pi4143, pi4144, pi4145, pi4146, pi4147, pi4148,
    pi4149, pi4150, pi4151, pi4152, pi4153, pi4154, pi4155, pi4156, pi4157,
    pi4158, pi4159, pi4160, pi4161, pi4162, pi4163, pi4164, pi4165, pi4166,
    pi4167, pi4168, pi4169, pi4170, pi4171, pi4172, pi4173, pi4174, pi4175,
    pi4176, pi4177, pi4178, pi4179, pi4180, pi4181, pi4182, pi4183, pi4184,
    pi4185, pi4186, pi4187, pi4188, pi4189, pi4190, pi4191, pi4192, pi4193,
    pi4194, pi4195, pi4196, pi4197, pi4198, pi4199, pi4200, pi4201, pi4202,
    pi4203, pi4204, pi4205, pi4206, pi4207, pi4208, pi4209, pi4210, pi4211,
    pi4212, pi4213, pi4214, pi4215, pi4216, pi4217, pi4218, pi4219, pi4220,
    pi4221, pi4222, pi4223, pi4224, pi4225, pi4226, pi4227, pi4228, pi4229,
    pi4230, pi4231, pi4232, pi4233, pi4234, pi4235, pi4236, pi4237, pi4238,
    pi4239, pi4240, pi4241, pi4242, pi4243, pi4244, pi4245, pi4246, pi4247,
    pi4248, pi4249, pi4250, pi4251, pi4252, pi4253, pi4254, pi4255, pi4256,
    pi4257, pi4258, pi4259, pi4260, pi4261, pi4262, pi4263, pi4264, pi4265,
    pi4266, pi4267, pi4268, pi4269, pi4270, pi4271, pi4272, pi4273, pi4274,
    pi4275, pi4276, pi4277, pi4278, pi4279, pi4280, pi4281, pi4282, pi4283,
    pi4284, pi4285, pi4286, pi4287, pi4288, pi4289, pi4290, pi4291, pi4292,
    pi4293, pi4294, pi4295, pi4296, pi4297, pi4298, pi4299, pi4300, pi4301,
    pi4302, pi4303, pi4304, pi4305, pi4306, pi4307, pi4308, pi4309, pi4310,
    pi4311, pi4312, pi4313, pi4314, pi4315, pi4316, pi4317, pi4318, pi4319,
    pi4320, pi4321, pi4322, pi4323, pi4324, pi4325, pi4326, pi4327, pi4328,
    pi4329, pi4330, pi4331, pi4332, pi4333, pi4334, pi4335, pi4336, pi4337,
    pi4338, pi4339, pi4340, pi4341, pi4342, pi4343, pi4344, pi4345, pi4346,
    pi4347, pi4348, pi4349, pi4350, pi4351, pi4352, pi4353, pi4354, pi4355,
    pi4356, pi4357, pi4358, pi4359, pi4360, pi4361, pi4362, pi4363, pi4364,
    pi4365, pi4366, pi4367, pi4368, pi4369, pi4370, pi4371, pi4372, pi4373,
    pi4374, pi4375, pi4376, pi4377, pi4378, pi4379, pi4380, pi4381, pi4382,
    pi4383, pi4384, pi4385, pi4386, pi4387, pi4388, pi4389, pi4390, pi4391,
    pi4392, pi4393, pi4394, pi4395, pi4396, pi4397, pi4398, pi4399, pi4400,
    pi4401, pi4402, pi4403, pi4404, pi4405, pi4406, pi4407, pi4408, pi4409,
    pi4410, pi4411, pi4412, pi4413, pi4414, pi4415, pi4416, pi4417, pi4418,
    pi4419, pi4420, pi4421, pi4422, pi4423, pi4424, pi4425, pi4426, pi4427,
    pi4428, pi4429, pi4430, pi4431, pi4432, pi4433, pi4434, pi4435, pi4436,
    pi4437, pi4438, pi4439, pi4440, pi4441, pi4442, pi4443, pi4444, pi4445,
    pi4446, pi4447, pi4448, pi4449, pi4450, pi4451, pi4452, pi4453, pi4454,
    pi4455, pi4456, pi4457, pi4458, pi4459, pi4460, pi4461, pi4462, pi4463,
    pi4464, pi4465, pi4466, pi4467, pi4468, pi4469, pi4470, pi4471, pi4472,
    pi4473, pi4474, pi4475, pi4476, pi4477, pi4478, pi4479, pi4480, pi4481,
    pi4482, pi4483, pi4484, pi4485, pi4486, pi4487, pi4488, pi4489, pi4490,
    pi4491, pi4492, pi4493, pi4494, pi4495, pi4496, pi4497, pi4498, pi4499,
    pi4500, pi4501, pi4502, pi4503, pi4504, pi4505, pi4506, pi4507, pi4508,
    pi4509, pi4510, pi4511, pi4512, pi4513, pi4514, pi4515, pi4516, pi4517,
    pi4518, pi4519, pi4520, pi4521, pi4522, pi4523, pi4524, pi4525, pi4526,
    pi4527, pi4528, pi4529, pi4530, pi4531, pi4532, pi4533, pi4534, pi4535,
    pi4536, pi4537, pi4538, pi4539, pi4540, pi4541, pi4542, pi4543, pi4544,
    pi4545, pi4546, pi4547, pi4548, pi4549, pi4550, pi4551, pi4552, pi4553,
    pi4554, pi4555, pi4556, pi4557, pi4558, pi4559, pi4560, pi4561, pi4562,
    pi4563, pi4564, pi4565, pi4566, pi4567, pi4568, pi4569, pi4570, pi4571,
    pi4572, pi4573, pi4574, pi4575, pi4576, pi4577, pi4578, pi4579, pi4580,
    pi4581, pi4582, pi4583, pi4584, pi4585, pi4586, pi4587, pi4588, pi4589,
    pi4590, pi4591, pi4592, pi4593, pi4594, pi4595, pi4596, pi4597, pi4598,
    pi4599, pi4600, pi4601, pi4602, pi4603, pi4604, pi4605, pi4606, pi4607,
    pi4608, pi4609, pi4610, pi4611, pi4612, pi4613, pi4614, pi4615, pi4616,
    pi4617, pi4618, pi4619, pi4620, pi4621, pi4622, pi4623, pi4624, pi4625,
    pi4626, pi4627, pi4628, pi4629, pi4630, pi4631, pi4632, pi4633, pi4634,
    pi4635, pi4636, pi4637, pi4638, pi4639, pi4640, pi4641, pi4642, pi4643,
    pi4644, pi4645, pi4646, pi4647, pi4648, pi4649, pi4650, pi4651, pi4652,
    pi4653, pi4654, pi4655, pi4656, pi4657, pi4658, pi4659, pi4660, pi4661,
    pi4662, pi4663, pi4664, pi4665, pi4666, pi4667, pi4668, pi4669, pi4670,
    pi4671, pi4672, pi4673, pi4674, pi4675, pi4676, pi4677, pi4678, pi4679,
    pi4680, pi4681, pi4682, pi4683, pi4684, pi4685, pi4686, pi4687, pi4688,
    pi4689, pi4690, pi4691, pi4692, pi4693, pi4694, pi4695, pi4696, pi4697,
    pi4698, pi4699, pi4700, pi4701, pi4702, pi4703, pi4704, pi4705, pi4706,
    pi4707, pi4708, pi4709, pi4710, pi4711, pi4712, pi4713, pi4714, pi4715,
    pi4716, pi4717, pi4718, pi4719, pi4720, pi4721, pi4722, pi4723, pi4724,
    pi4725, pi4726, pi4727, pi4728, pi4729, pi4730, pi4731, pi4732, pi4733,
    pi4734, pi4735, pi4736, pi4737, pi4738, pi4739, pi4740, pi4741, pi4742,
    pi4743, pi4744, pi4745, pi4746, pi4747, pi4748, pi4749, pi4750, pi4751,
    pi4752, pi4753, pi4754, pi4755, pi4756, pi4757, pi4758, pi4759, pi4760,
    pi4761, pi4762, pi4763, pi4764, pi4765, pi4766, pi4767, pi4768, pi4769,
    pi4770, pi4771, pi4772, pi4773, pi4774, pi4775, pi4776, pi4777, pi4778,
    pi4779, pi4780, pi4781, pi4782, pi4783, pi4784, pi4785, pi4786, pi4787,
    pi4788, pi4789, pi4790, pi4791, pi4792, pi4793, pi4794, pi4795, pi4796,
    pi4797, pi4798, pi4799, pi4800, pi4801, pi4802, pi4803, pi4804, pi4805,
    pi4806, pi4807, pi4808, pi4809, pi4810, pi4811, pi4812, pi4813, pi4814,
    pi4815, pi4816, pi4817, pi4818, pi4819, pi4820, pi4821, pi4822, pi4823,
    pi4824, pi4825, pi4826, pi4827, pi4828, pi4829, pi4830, pi4831, pi4832,
    pi4833, pi4834, pi4835, pi4836, pi4837, pi4838, pi4839, pi4840, pi4841,
    pi4842, pi4843, pi4844, pi4845, pi4846, pi4847, pi4848, pi4849, pi4850,
    pi4851, pi4852, pi4853, pi4854, pi4855, pi4856, pi4857, pi4858, pi4859,
    pi4860, pi4861, pi4862, pi4863, pi4864, pi4865, pi4866, pi4867, pi4868,
    pi4869, pi4870, pi4871, pi4872, pi4873, pi4874, pi4875, pi4876, pi4877,
    pi4878, pi4879, pi4880, pi4881, pi4882, pi4883, pi4884, pi4885, pi4886,
    pi4887, pi4888, pi4889, pi4890, pi4891, pi4892, pi4893, pi4894, pi4895,
    pi4896, pi4897, pi4898, pi4899, pi4900, pi4901, pi4902, pi4903, pi4904,
    pi4905, pi4906, pi4907, pi4908, pi4909, pi4910, pi4911, pi4912, pi4913,
    pi4914, pi4915, pi4916, pi4917, pi4918, pi4919, pi4920, pi4921, pi4922,
    pi4923, pi4924, pi4925, pi4926, pi4927, pi4928, pi4929, pi4930, pi4931,
    pi4932, pi4933, pi4934, pi4935, pi4936, pi4937, pi4938, pi4939, pi4940,
    pi4941, pi4942, pi4943, pi4944, pi4945, pi4946, pi4947, pi4948, pi4949,
    pi4950, pi4951, pi4952, pi4953, pi4954, pi4955, pi4956, pi4957, pi4958,
    pi4959, pi4960, pi4961, pi4962, pi4963, pi4964, pi4965, pi4966, pi4967,
    pi4968, pi4969, pi4970, pi4971, pi4972, pi4973, pi4974, pi4975, pi4976,
    pi4977, pi4978, pi4979, pi4980, pi4981, pi4982, pi4983, pi4984, pi4985,
    pi4986, pi4987, pi4988, pi4989, pi4990, pi4991, pi4992, pi4993, pi4994,
    pi4995, pi4996, pi4997, pi4998, pi4999, pi5000, pi5001, pi5002, pi5003,
    pi5004, pi5005, pi5006, pi5007, pi5008, pi5009, pi5010, pi5011, pi5012,
    pi5013, pi5014, pi5015, pi5016, pi5017, pi5018, pi5019, pi5020, pi5021,
    pi5022, pi5023, pi5024, pi5025, pi5026, pi5027, pi5028, pi5029, pi5030,
    pi5031, pi5032, pi5033, pi5034, pi5035, pi5036, pi5037, pi5038, pi5039,
    pi5040, pi5041, pi5042, pi5043, pi5044, pi5045, pi5046, pi5047, pi5048,
    pi5049, pi5050, pi5051, pi5052, pi5053, pi5054, pi5055, pi5056, pi5057,
    pi5058, pi5059, pi5060, pi5061, pi5062, pi5063, pi5064, pi5065, pi5066,
    pi5067, pi5068, pi5069, pi5070, pi5071, pi5072, pi5073, pi5074, pi5075,
    pi5076, pi5077, pi5078, pi5079, pi5080, pi5081, pi5082, pi5083, pi5084,
    pi5085, pi5086, pi5087, pi5088, pi5089, pi5090, pi5091, pi5092, pi5093,
    pi5094, pi5095, pi5096, pi5097, pi5098, pi5099, pi5100, pi5101, pi5102,
    pi5103, pi5104, pi5105, pi5106, pi5107, pi5108, pi5109, pi5110, pi5111,
    pi5112, pi5113, pi5114, pi5115, pi5116, pi5117, pi5118, pi5119, pi5120,
    pi5121, pi5122, pi5123, pi5124, pi5125, pi5126, pi5127, pi5128, pi5129,
    pi5130, pi5131, pi5132, pi5133, pi5134, pi5135, pi5136, pi5137, pi5138,
    pi5139, pi5140, pi5141, pi5142, pi5143, pi5144, pi5145, pi5146, pi5147,
    pi5148, pi5149, pi5150, pi5151, pi5152, pi5153, pi5154, pi5155, pi5156,
    pi5157, pi5158, pi5159, pi5160, pi5161, pi5162, pi5163, pi5164, pi5165,
    pi5166, pi5167, pi5168, pi5169, pi5170, pi5171, pi5172, pi5173, pi5174,
    pi5175, pi5176, pi5177, pi5178, pi5179, pi5180, pi5181, pi5182, pi5183,
    pi5184, pi5185, pi5186, pi5187, pi5188, pi5189, pi5190, pi5191, pi5192,
    pi5193, pi5194, pi5195, pi5196, pi5197, pi5198, pi5199, pi5200, pi5201,
    pi5202, pi5203, pi5204, pi5205, pi5206, pi5207, pi5208, pi5209, pi5210,
    pi5211, pi5212, pi5213, pi5214, pi5215, pi5216, pi5217, pi5218, pi5219,
    pi5220, pi5221, pi5222, pi5223, pi5224, pi5225, pi5226, pi5227, pi5228,
    pi5229, pi5230, pi5231, pi5232, pi5233, pi5234, pi5235, pi5236, pi5237,
    pi5238, pi5239, pi5240, pi5241, pi5242, pi5243, pi5244, pi5245, pi5246,
    pi5247, pi5248, pi5249, pi5250, pi5251, pi5252, pi5253, pi5254, pi5255,
    pi5256, pi5257, pi5258, pi5259, pi5260, pi5261, pi5262, pi5263, pi5264,
    pi5265, pi5266, pi5267, pi5268, pi5269, pi5270, pi5271, pi5272, pi5273,
    pi5274, pi5275, pi5276, pi5277, pi5278, pi5279, pi5280, pi5281, pi5282,
    pi5283, pi5284, pi5285, pi5286, pi5287, pi5288, pi5289, pi5290, pi5291,
    pi5292, pi5293, pi5294, pi5295, pi5296, pi5297, pi5298, pi5299, pi5300,
    pi5301, pi5302, pi5303, pi5304, pi5305, pi5306, pi5307, pi5308, pi5309,
    pi5310, pi5311, pi5312, pi5313, pi5314, pi5315, pi5316, pi5317, pi5318,
    pi5319, pi5320, pi5321, pi5322, pi5323, pi5324, pi5325, pi5326, pi5327,
    pi5328, pi5329, pi5330, pi5331, pi5332, pi5333, pi5334, pi5335, pi5336,
    pi5337, pi5338, pi5339, pi5340, pi5341, pi5342, pi5343, pi5344, pi5345,
    pi5346, pi5347, pi5348, pi5349, pi5350, pi5351, pi5352, pi5353, pi5354,
    pi5355, pi5356, pi5357, pi5358, pi5359, pi5360, pi5361, pi5362, pi5363,
    pi5364, pi5365, pi5366, pi5367, pi5368, pi5369, pi5370, pi5371, pi5372,
    pi5373, pi5374, pi5375, pi5376, pi5377, pi5378, pi5379, pi5380, pi5381,
    pi5382, pi5383, pi5384, pi5385, pi5386, pi5387, pi5388, pi5389, pi5390,
    pi5391, pi5392, pi5393, pi5394, pi5395, pi5396, pi5397, pi5398, pi5399,
    pi5400, pi5401, pi5402, pi5403, pi5404, pi5405, pi5406, pi5407, pi5408,
    pi5409, pi5410, pi5411, pi5412, pi5413, pi5414, pi5415, pi5416, pi5417,
    pi5418, pi5419, pi5420, pi5421, pi5422, pi5423, pi5424, pi5425, pi5426,
    pi5427, pi5428, pi5429, pi5430, pi5431, pi5432, pi5433, pi5434, pi5435,
    pi5436, pi5437, pi5438, pi5439, pi5440, pi5441, pi5442, pi5443, pi5444,
    pi5445, pi5446, pi5447, pi5448, pi5449, pi5450, pi5451, pi5452, pi5453,
    pi5454, pi5455, pi5456, pi5457, pi5458, pi5459, pi5460, pi5461, pi5462,
    pi5463, pi5464, pi5465, pi5466, pi5467, pi5468, pi5469, pi5470, pi5471,
    pi5472, pi5473, pi5474, pi5475, pi5476, pi5477, pi5478, pi5479, pi5480,
    pi5481, pi5482, pi5483, pi5484, pi5485, pi5486, pi5487, pi5488, pi5489,
    pi5490, pi5491, pi5492, pi5493, pi5494, pi5495, pi5496, pi5497, pi5498,
    pi5499, pi5500, pi5501, pi5502, pi5503, pi5504, pi5505, pi5506, pi5507,
    pi5508, pi5509, pi5510, pi5511, pi5512, pi5513, pi5514, pi5515, pi5516,
    pi5517, pi5518, pi5519, pi5520, pi5521, pi5522, pi5523, pi5524, pi5525,
    pi5526, pi5527, pi5528, pi5529, pi5530, pi5531, pi5532, pi5533, pi5534,
    pi5535, pi5536, pi5537, pi5538, pi5539, pi5540, pi5541, pi5542, pi5543,
    pi5544, pi5545, pi5546, pi5547, pi5548, pi5549, pi5550, pi5551, pi5552,
    pi5553, pi5554, pi5555, pi5556, pi5557, pi5558, pi5559, pi5560, pi5561,
    pi5562, pi5563, pi5564, pi5565, pi5566, pi5567, pi5568, pi5569, pi5570,
    pi5571, pi5572, pi5573, pi5574, pi5575, pi5576, pi5577, pi5578, pi5579,
    pi5580, pi5581, pi5582, pi5583, pi5584, pi5585, pi5586, pi5587, pi5588,
    pi5589, pi5590, pi5591, pi5592, pi5593, pi5594, pi5595, pi5596, pi5597,
    pi5598, pi5599, pi5600, pi5601, pi5602, pi5603, pi5604, pi5605, pi5606,
    pi5607, pi5608, pi5609, pi5610, pi5611, pi5612, pi5613, pi5614, pi5615,
    pi5616, pi5617, pi5618, pi5619, pi5620, pi5621, pi5622, pi5623, pi5624,
    pi5625, pi5626, pi5627, pi5628, pi5629, pi5630, pi5631, pi5632, pi5633,
    pi5634, pi5635, pi5636, pi5637, pi5638, pi5639, pi5640, pi5641, pi5642,
    pi5643, pi5644, pi5645, pi5646, pi5647, pi5648, pi5649, pi5650, pi5651,
    pi5652, pi5653, pi5654, pi5655, pi5656, pi5657, pi5658, pi5659, pi5660,
    pi5661, pi5662, pi5663, pi5664, pi5665, pi5666, pi5667, pi5668, pi5669,
    pi5670, pi5671, pi5672, pi5673, pi5674, pi5675, pi5676, pi5677, pi5678,
    pi5679, pi5680, pi5681, pi5682, pi5683, pi5684, pi5685, pi5686, pi5687,
    pi5688, pi5689, pi5690, pi5691, pi5692, pi5693, pi5694, pi5695, pi5696,
    pi5697, pi5698, pi5699, pi5700, pi5701, pi5702, pi5703, pi5704, pi5705,
    pi5706, pi5707, pi5708, pi5709, pi5710, pi5711, pi5712, pi5713, pi5714,
    pi5715, pi5716, pi5717, pi5718, pi5719, pi5720, pi5721, pi5722, pi5723,
    pi5724, pi5725, pi5726, pi5727, pi5728, pi5729, pi5730, pi5731, pi5732,
    pi5733, pi5734, pi5735, pi5736, pi5737, pi5738, pi5739, pi5740, pi5741,
    pi5742, pi5743, pi5744, pi5745, pi5746, pi5747, pi5748, pi5749, pi5750,
    pi5751, pi5752, pi5753, pi5754, pi5755, pi5756, pi5757, pi5758, pi5759,
    pi5760, pi5761, pi5762, pi5763, pi5764, pi5765, pi5766, pi5767, pi5768,
    pi5769, pi5770, pi5771, pi5772, pi5773, pi5774, pi5775, pi5776, pi5777,
    pi5778, pi5779, pi5780, pi5781, pi5782, pi5783, pi5784, pi5785, pi5786,
    pi5787, pi5788, pi5789, pi5790, pi5791, pi5792, pi5793, pi5794, pi5795,
    pi5796, pi5797, pi5798, pi5799, pi5800, pi5801, pi5802, pi5803, pi5804,
    pi5805, pi5806, pi5807, pi5808, pi5809, pi5810, pi5811, pi5812, pi5813,
    pi5814, pi5815, pi5816, pi5817, pi5818, pi5819, pi5820, pi5821, pi5822,
    pi5823, pi5824, pi5825, pi5826, pi5827, pi5828, pi5829, pi5830, pi5831,
    pi5832, pi5833, pi5834, pi5835, pi5836, pi5837, pi5838, pi5839, pi5840,
    pi5841, pi5842, pi5843, pi5844, pi5845, pi5846, pi5847, pi5848, pi5849,
    pi5850, pi5851, pi5852, pi5853, pi5854, pi5855, pi5856, pi5857, pi5858,
    pi5859, pi5860, pi5861, pi5862, pi5863, pi5864, pi5865, pi5866, pi5867,
    pi5868, pi5869, pi5870, pi5871, pi5872, pi5873, pi5874, pi5875, pi5876,
    pi5877, pi5878, pi5879, pi5880, pi5881, pi5882, pi5883, pi5884, pi5885,
    pi5886, pi5887, pi5888, pi5889, pi5890, pi5891, pi5892, pi5893, pi5894,
    pi5895, pi5896, pi5897, pi5898, pi5899, pi5900, pi5901, pi5902, pi5903,
    pi5904, pi5905, pi5906, pi5907, pi5908, pi5909, pi5910, pi5911, pi5912,
    pi5913, pi5914, pi5915, pi5916, pi5917, pi5918, pi5919, pi5920, pi5921,
    pi5922, pi5923, pi5924, pi5925, pi5926, pi5927, pi5928, pi5929, pi5930,
    pi5931, pi5932, pi5933, pi5934, pi5935, pi5936, pi5937, pi5938, pi5939,
    pi5940, pi5941, pi5942, pi5943, pi5944, pi5945, pi5946, pi5947, pi5948,
    pi5949, pi5950, pi5951, pi5952, pi5953, pi5954, pi5955, pi5956, pi5957,
    pi5958, pi5959, pi5960, pi5961, pi5962, pi5963, pi5964, pi5965, pi5966,
    pi5967, pi5968, pi5969, pi5970, pi5971, pi5972, pi5973, pi5974, pi5975,
    pi5976, pi5977, pi5978, pi5979, pi5980, pi5981, pi5982, pi5983, pi5984,
    pi5985, pi5986, pi5987, pi5988, pi5989, pi5990, pi5991, pi5992, pi5993,
    pi5994, pi5995, pi5996, pi5997, pi5998, pi5999, pi6000, pi6001, pi6002,
    pi6003, pi6004, pi6005, pi6006, pi6007, pi6008, pi6009, pi6010, pi6011,
    pi6012, pi6013, pi6014, pi6015, pi6016, pi6017, pi6018, pi6019, pi6020,
    pi6021, pi6022, pi6023, pi6024, pi6025, pi6026, pi6027, pi6028, pi6029,
    pi6030, pi6031, pi6032, pi6033, pi6034, pi6035, pi6036, pi6037, pi6038,
    pi6039, pi6040, pi6041, pi6042, pi6043, pi6044, pi6045, pi6046, pi6047,
    pi6048, pi6049, pi6050, pi6051, pi6052, pi6053, pi6054, pi6055, pi6056,
    pi6057, pi6058, pi6059, pi6060, pi6061, pi6062, pi6063, pi6064, pi6065,
    pi6066, pi6067, pi6068, pi6069, pi6070, pi6071, pi6072, pi6073, pi6074,
    pi6075, pi6076, pi6077, pi6078, pi6079, pi6080, pi6081, pi6082, pi6083,
    pi6084, pi6085, pi6086, pi6087, pi6088, pi6089, pi6090, pi6091, pi6092,
    pi6093, pi6094, pi6095, pi6096, pi6097, pi6098, pi6099, pi6100, pi6101,
    pi6102, pi6103, pi6104, pi6105, pi6106, pi6107, pi6108, pi6109, pi6110,
    pi6111, pi6112, pi6113, pi6114, pi6115, pi6116, pi6117, pi6118, pi6119,
    pi6120, pi6121, pi6122, pi6123, pi6124, pi6125, pi6126, pi6127, pi6128,
    pi6129, pi6130, pi6131, pi6132, pi6133, pi6134, pi6135, pi6136, pi6137,
    pi6138, pi6139, pi6140, pi6141, pi6142, pi6143, pi6144, pi6145, pi6146,
    pi6147, pi6148, pi6149, pi6150, pi6151, pi6152, pi6153, pi6154, pi6155,
    pi6156, pi6157, pi6158, pi6159, pi6160, pi6161, pi6162, pi6163, pi6164,
    pi6165, pi6166, pi6167, pi6168, pi6169, pi6170, pi6171, pi6172, pi6173,
    pi6174, pi6175, pi6176, pi6177, pi6178, pi6179, pi6180, pi6181, pi6182,
    pi6183, pi6184, pi6185, pi6186, pi6187, pi6188, pi6189, pi6190, pi6191,
    pi6192, pi6193, pi6194, pi6195, pi6196, pi6197, pi6198, pi6199, pi6200,
    pi6201, pi6202, pi6203, pi6204, pi6205, pi6206, pi6207, pi6208, pi6209,
    pi6210, pi6211, pi6212, pi6213, pi6214, pi6215, pi6216, pi6217, pi6218,
    pi6219, pi6220, pi6221, pi6222, pi6223, pi6224, pi6225, pi6226, pi6227,
    pi6228, pi6229, pi6230, pi6231, pi6232, pi6233, pi6234, pi6235, pi6236,
    pi6237, pi6238, pi6239, pi6240, pi6241, pi6242, pi6243, pi6244, pi6245,
    pi6246, pi6247, pi6248, pi6249, pi6250, pi6251, pi6252, pi6253, pi6254,
    pi6255, pi6256, pi6257, pi6258, pi6259, pi6260, pi6261, pi6262, pi6263,
    pi6264, pi6265, pi6266, pi6267, pi6268, pi6269, pi6270, pi6271, pi6272,
    pi6273, pi6274, pi6275, pi6276, pi6277, pi6278, pi6279, pi6280, pi6281,
    pi6282, pi6283, pi6284, pi6285, pi6286, pi6287, pi6288, pi6289, pi6290,
    pi6291, pi6292, pi6293, pi6294, pi6295, pi6296, pi6297, pi6298, pi6299,
    pi6300, pi6301, pi6302, pi6303, pi6304, pi6305, pi6306, pi6307, pi6308,
    pi6309, pi6310, pi6311, pi6312, pi6313, pi6314, pi6315, pi6316, pi6317,
    pi6318, pi6319, pi6320, pi6321, pi6322, pi6323, pi6324, pi6325, pi6326,
    pi6327, pi6328, pi6329, pi6330, pi6331, pi6332, pi6333, pi6334, pi6335,
    pi6336, pi6337, pi6338, pi6339, pi6340, pi6341, pi6342, pi6343, pi6344,
    pi6345, pi6346, pi6347, pi6348, pi6349, pi6350, pi6351, pi6352, pi6353,
    pi6354, pi6355, pi6356, pi6357, pi6358, pi6359, pi6360, pi6361, pi6362,
    pi6363, pi6364, pi6365, pi6366, pi6367, pi6368, pi6369, pi6370, pi6371,
    pi6372, pi6373, pi6374, pi6375, pi6376, pi6377, pi6378, pi6379, pi6380,
    pi6381, pi6382, pi6383, pi6384, pi6385, pi6386, pi6387, pi6388, pi6389,
    pi6390, pi6391, pi6392, pi6393, pi6394, pi6395, pi6396, pi6397, pi6398,
    pi6399, pi6400, pi6401, pi6402, pi6403, pi6404, pi6405, pi6406, pi6407,
    pi6408, pi6409, pi6410, pi6411, pi6412, pi6413, pi6414, pi6415, pi6416,
    pi6417, pi6418, pi6419, pi6420, pi6421, pi6422, pi6423, pi6424, pi6425,
    pi6426, pi6427, pi6428, pi6429, pi6430, pi6431, pi6432, pi6433, pi6434,
    pi6435, pi6436, pi6437, pi6438, pi6439, pi6440, pi6441, pi6442, pi6443,
    pi6444, pi6445, pi6446, pi6447, pi6448, pi6449, pi6450, pi6451, pi6452,
    pi6453, pi6454, pi6455, pi6456, pi6457, pi6458, pi6459, pi6460, pi6461,
    pi6462, pi6463, pi6464, pi6465, pi6466, pi6467, pi6468, pi6469, pi6470,
    pi6471, pi6472, pi6473, pi6474, pi6475, pi6476, pi6477, pi6478, pi6479,
    pi6480, pi6481, pi6482, pi6483, pi6484, pi6485, pi6486, pi6487, pi6488,
    pi6489, pi6490, pi6491, pi6492, pi6493, pi6494, pi6495, pi6496, pi6497,
    pi6498, pi6499, pi6500, pi6501, pi6502, pi6503, pi6504, pi6505, pi6506,
    pi6507, pi6508, pi6509, pi6510, pi6511, pi6512, pi6513, pi6514, pi6515,
    pi6516, pi6517, pi6518, pi6519, pi6520, pi6521, pi6522, pi6523, pi6524,
    pi6525, pi6526, pi6527, pi6528, pi6529, pi6530, pi6531, pi6532, pi6533,
    pi6534, pi6535, pi6536, pi6537, pi6538, pi6539, pi6540, pi6541, pi6542,
    pi6543, pi6544, pi6545, pi6546, pi6547, pi6548, pi6549, pi6550, pi6551,
    pi6552, pi6553, pi6554, pi6555, pi6556, pi6557, pi6558, pi6559, pi6560,
    pi6561, pi6562, pi6563, pi6564, pi6565, pi6566, pi6567, pi6568, pi6569,
    pi6570, pi6571, pi6572, pi6573, pi6574, pi6575, pi6576, pi6577, pi6578,
    pi6579, pi6580, pi6581, pi6582, pi6583, pi6584, pi6585, pi6586, pi6587,
    pi6588, pi6589, pi6590, pi6591, pi6592, pi6593, pi6594, pi6595, pi6596,
    pi6597, pi6598, pi6599, pi6600, pi6601, pi6602, pi6603, pi6604, pi6605,
    pi6606, pi6607, pi6608, pi6609, pi6610, pi6611, pi6612, pi6613, pi6614,
    pi6615, pi6616, pi6617, pi6618, pi6619, pi6620, pi6621, pi6622, pi6623,
    pi6624, pi6625, pi6626, pi6627, pi6628, pi6629, pi6630, pi6631, pi6632,
    pi6633, pi6634, pi6635, pi6636, pi6637, pi6638, pi6639, pi6640, pi6641,
    pi6642, pi6643, pi6644, pi6645, pi6646, pi6647, pi6648, pi6649, pi6650,
    pi6651, pi6652, pi6653, pi6654, pi6655, pi6656, pi6657, pi6658, pi6659,
    pi6660, pi6661, pi6662, pi6663, pi6664, pi6665, pi6666, pi6667, pi6668,
    pi6669, pi6670, pi6671, pi6672, pi6673, pi6674, pi6675, pi6676, pi6677,
    pi6678, pi6679, pi6680, pi6681, pi6682, pi6683, pi6684, pi6685, pi6686,
    pi6687, pi6688, pi6689, pi6690, pi6691, pi6692, pi6693, pi6694, pi6695,
    pi6696, pi6697, pi6698, pi6699, pi6700, pi6701, pi6702, pi6703, pi6704,
    pi6705, pi6706, pi6707, pi6708, pi6709, pi6710, pi6711, pi6712, pi6713,
    pi6714, pi6715, pi6716, pi6717, pi6718, pi6719, pi6720, pi6721, pi6722,
    pi6723, pi6724, pi6725, pi6726, pi6727, pi6728, pi6729, pi6730, pi6731,
    pi6732, pi6733, pi6734, pi6735, pi6736, pi6737, pi6738, pi6739, pi6740,
    pi6741, pi6742, pi6743, pi6744, pi6745, pi6746, pi6747, pi6748, pi6749,
    pi6750, pi6751, pi6752, pi6753, pi6754, pi6755, pi6756, pi6757, pi6758,
    pi6759, pi6760, pi6761, pi6762, pi6763, pi6764, pi6765, pi6766, pi6767,
    pi6768, pi6769, pi6770, pi6771, pi6772, pi6773, pi6774, pi6775, pi6776,
    pi6777, pi6778, pi6779, pi6780, pi6781, pi6782, pi6783, pi6784, pi6785,
    pi6786, pi6787, pi6788, pi6789, pi6790, pi6791, pi6792, pi6793, pi6794,
    pi6795, pi6796, pi6797, pi6798, pi6799, pi6800, pi6801, pi6802, pi6803,
    pi6804, pi6805, pi6806, pi6807, pi6808, pi6809, pi6810, pi6811, pi6812,
    pi6813, pi6814, pi6815, pi6816, pi6817, pi6818, pi6819, pi6820, pi6821,
    pi6822, pi6823, pi6824, pi6825, pi6826, pi6827, pi6828, pi6829, pi6830,
    pi6831, pi6832, pi6833, pi6834, pi6835, pi6836, pi6837, pi6838, pi6839,
    pi6840, pi6841, pi6842, pi6843, pi6844, pi6845, pi6846, pi6847, pi6848,
    pi6849, pi6850, pi6851, pi6852, pi6853, pi6854, pi6855, pi6856, pi6857,
    pi6858, pi6859, pi6860, pi6861, pi6862, pi6863, pi6864, pi6865, pi6866,
    pi6867, pi6868, pi6869, pi6870, pi6871, pi6872, pi6873, pi6874, pi6875,
    pi6876, pi6877, pi6878, pi6879, pi6880, pi6881, pi6882, pi6883, pi6884,
    pi6885, pi6886, pi6887, pi6888, pi6889, pi6890, pi6891, pi6892, pi6893,
    pi6894, pi6895, pi6896, pi6897, pi6898, pi6899, pi6900, pi6901, pi6902,
    pi6903, pi6904, pi6905, pi6906, pi6907, pi6908, pi6909, pi6910, pi6911,
    pi6912, pi6913, pi6914, pi6915, pi6916, pi6917, pi6918, pi6919, pi6920,
    pi6921, pi6922, pi6923, pi6924, pi6925, pi6926, pi6927, pi6928, pi6929,
    pi6930, pi6931, pi6932, pi6933, pi6934, pi6935, pi6936, pi6937, pi6938,
    pi6939, pi6940, pi6941, pi6942, pi6943, pi6944, pi6945, pi6946, pi6947,
    pi6948, pi6949, pi6950, pi6951, pi6952, pi6953, pi6954, pi6955, pi6956,
    pi6957, pi6958, pi6959, pi6960, pi6961, pi6962, pi6963, pi6964, pi6965,
    pi6966, pi6967, pi6968, pi6969, pi6970, pi6971, pi6972, pi6973, pi6974,
    pi6975, pi6976, pi6977, pi6978, pi6979, pi6980, pi6981, pi6982, pi6983,
    pi6984, pi6985, pi6986, pi6987, pi6988, pi6989, pi6990, pi6991, pi6992,
    pi6993, pi6994, pi6995, pi6996, pi6997, pi6998, pi6999, pi7000, pi7001,
    pi7002, pi7003, pi7004, pi7005, pi7006, pi7007, pi7008, pi7009, pi7010,
    pi7011, pi7012, pi7013, pi7014, pi7015, pi7016, pi7017, pi7018, pi7019,
    pi7020, pi7021, pi7022, pi7023, pi7024, pi7025, pi7026, pi7027, pi7028,
    pi7029, pi7030, pi7031, pi7032, pi7033, pi7034, pi7035, pi7036, pi7037,
    pi7038, pi7039, pi7040, pi7041, pi7042, pi7043, pi7044, pi7045, pi7046,
    pi7047, pi7048, pi7049, pi7050, pi7051, pi7052, pi7053, pi7054, pi7055,
    pi7056, pi7057, pi7058, pi7059, pi7060, pi7061, pi7062, pi7063, pi7064,
    pi7065, pi7066, pi7067, pi7068, pi7069, pi7070, pi7071, pi7072, pi7073,
    pi7074, pi7075, pi7076, pi7077, pi7078, pi7079, pi7080, pi7081, pi7082,
    pi7083, pi7084, pi7085, pi7086, pi7087, pi7088, pi7089, pi7090, pi7091,
    pi7092, pi7093, pi7094, pi7095, pi7096, pi7097, pi7098, pi7099, pi7100,
    pi7101, pi7102, pi7103, pi7104, pi7105, pi7106, pi7107, pi7108, pi7109,
    pi7110, pi7111, pi7112, pi7113, pi7114, pi7115, pi7116, pi7117, pi7118,
    pi7119, pi7120, pi7121, pi7122, pi7123, pi7124, pi7125, pi7126, pi7127,
    pi7128, pi7129, pi7130, pi7131, pi7132, pi7133, pi7134, pi7135, pi7136,
    pi7137, pi7138, pi7139, pi7140, pi7141, pi7142, pi7143, pi7144, pi7145,
    pi7146, pi7147, pi7148, pi7149, pi7150, pi7151, pi7152, pi7153, pi7154,
    pi7155, pi7156, pi7157, pi7158, pi7159, pi7160, pi7161, pi7162, pi7163,
    pi7164, pi7165, pi7166, pi7167, pi7168, pi7169, pi7170, pi7171, pi7172,
    pi7173, pi7174, pi7175, pi7176, pi7177, pi7178, pi7179, pi7180, pi7181,
    pi7182, pi7183, pi7184, pi7185, pi7186, pi7187, pi7188, pi7189, pi7190,
    pi7191, pi7192, pi7193, pi7194, pi7195, pi7196, pi7197, pi7198, pi7199,
    pi7200, pi7201, pi7202, pi7203, pi7204, pi7205, pi7206, pi7207, pi7208,
    pi7209, pi7210, pi7211, pi7212, pi7213, pi7214, pi7215, pi7216, pi7217,
    pi7218, pi7219, pi7220, pi7221, pi7222, pi7223, pi7224, pi7225, pi7226,
    pi7227, pi7228, pi7229, pi7230, pi7231, pi7232, pi7233, pi7234, pi7235,
    pi7236, pi7237, pi7238, pi7239, pi7240, pi7241, pi7242, pi7243, pi7244,
    pi7245, pi7246, pi7247, pi7248, pi7249, pi7250, pi7251, pi7252, pi7253,
    pi7254, pi7255, pi7256, pi7257, pi7258, pi7259, pi7260, pi7261, pi7262,
    pi7263, pi7264, pi7265, pi7266, pi7267, pi7268, pi7269, pi7270, pi7271,
    pi7272, pi7273, pi7274, pi7275, pi7276, pi7277, pi7278, pi7279, pi7280,
    pi7281, pi7282, pi7283, pi7284, pi7285, pi7286, pi7287, pi7288, pi7289,
    pi7290, pi7291, pi7292, pi7293, pi7294, pi7295, pi7296, pi7297, pi7298,
    pi7299, pi7300, pi7301, pi7302, pi7303, pi7304, pi7305, pi7306, pi7307,
    pi7308, pi7309, pi7310, pi7311, pi7312, pi7313, pi7314, pi7315, pi7316,
    pi7317, pi7318, pi7319, pi7320, pi7321, pi7322, pi7323, pi7324, pi7325,
    pi7326, pi7327, pi7328, pi7329, pi7330, pi7331, pi7332, pi7333, pi7334,
    pi7335, pi7336, pi7337, pi7338, pi7339, pi7340, pi7341, pi7342, pi7343,
    pi7344, pi7345, pi7346, pi7347, pi7348, pi7349, pi7350, pi7351, pi7352,
    pi7353, pi7354, pi7355, pi7356, pi7357, pi7358, pi7359, pi7360, pi7361,
    pi7362, pi7363, pi7364, pi7365, pi7366, pi7367, pi7368, pi7369, pi7370,
    pi7371, pi7372, pi7373, pi7374, pi7375, pi7376, pi7377, pi7378, pi7379,
    pi7380, pi7381, pi7382, pi7383, pi7384, pi7385, pi7386, pi7387, pi7388,
    pi7389, pi7390, pi7391, pi7392, pi7393, pi7394, pi7395, pi7396, pi7397,
    pi7398, pi7399, pi7400, pi7401, pi7402, pi7403, pi7404, pi7405, pi7406,
    pi7407, pi7408, pi7409, pi7410, pi7411, pi7412, pi7413, pi7414, pi7415,
    pi7416, pi7417, pi7418, pi7419, pi7420, pi7421, pi7422, pi7423, pi7424,
    pi7425, pi7426, pi7427, pi7428, pi7429, pi7430, pi7431, pi7432, pi7433,
    pi7434, pi7435, pi7436, pi7437, pi7438, pi7439, pi7440, pi7441, pi7442,
    pi7443, pi7444, pi7445, pi7446, pi7447, pi7448, pi7449, pi7450, pi7451,
    pi7452, pi7453, pi7454, pi7455, pi7456, pi7457, pi7458, pi7459, pi7460,
    pi7461, pi7462, pi7463, pi7464, pi7465, pi7466, pi7467, pi7468, pi7469,
    pi7470, pi7471, pi7472, pi7473, pi7474, pi7475, pi7476, pi7477, pi7478,
    pi7479, pi7480, pi7481, pi7482, pi7483, pi7484, pi7485, pi7486, pi7487,
    pi7488, pi7489, pi7490, pi7491, pi7492, pi7493, pi7494, pi7495, pi7496,
    pi7497, pi7498, pi7499, pi7500, pi7501, pi7502, pi7503, pi7504, pi7505,
    pi7506, pi7507, pi7508, pi7509, pi7510, pi7511, pi7512, pi7513, pi7514,
    pi7515, pi7516, pi7517, pi7518, pi7519, pi7520, pi7521, pi7522, pi7523,
    pi7524, pi7525, pi7526, pi7527, pi7528, pi7529, pi7530, pi7531, pi7532,
    pi7533, pi7534, pi7535, pi7536, pi7537, pi7538, pi7539, pi7540, pi7541,
    pi7542, pi7543, pi7544, pi7545, pi7546, pi7547, pi7548, pi7549, pi7550,
    pi7551, pi7552, pi7553, pi7554, pi7555, pi7556, pi7557, pi7558, pi7559,
    pi7560, pi7561, pi7562, pi7563, pi7564, pi7565, pi7566, pi7567, pi7568,
    pi7569, pi7570, pi7571, pi7572, pi7573, pi7574, pi7575, pi7576, pi7577,
    pi7578, pi7579, pi7580, pi7581, pi7582, pi7583, pi7584, pi7585, pi7586,
    pi7587, pi7588, pi7589, pi7590, pi7591, pi7592, pi7593, pi7594, pi7595,
    pi7596, pi7597, pi7598, pi7599, pi7600, pi7601, pi7602, pi7603, pi7604,
    pi7605, pi7606, pi7607, pi7608, pi7609, pi7610, pi7611, pi7612, pi7613,
    pi7614, pi7615, pi7616, pi7617, pi7618, pi7619, pi7620, pi7621, pi7622,
    pi7623, pi7624, pi7625, pi7626, pi7627, pi7628, pi7629, pi7630, pi7631,
    pi7632, pi7633, pi7634, pi7635, pi7636, pi7637, pi7638, pi7639, pi7640,
    pi7641, pi7642, pi7643, pi7644, pi7645, pi7646, pi7647, pi7648, pi7649,
    pi7650, pi7651, pi7652, pi7653, pi7654, pi7655, pi7656, pi7657, pi7658,
    pi7659, pi7660, pi7661, pi7662, pi7663, pi7664, pi7665, pi7666, pi7667,
    pi7668, pi7669, pi7670, pi7671, pi7672, pi7673, pi7674, pi7675, pi7676,
    pi7677, pi7678, pi7679, pi7680, pi7681, pi7682, pi7683, pi7684, pi7685,
    pi7686, pi7687, pi7688, pi7689, pi7690, pi7691, pi7692, pi7693, pi7694,
    pi7695, pi7696, pi7697, pi7698, pi7699, pi7700, pi7701, pi7702, pi7703,
    pi7704, pi7705, pi7706, pi7707, pi7708, pi7709, pi7710, pi7711, pi7712,
    pi7713, pi7714, pi7715, pi7716, pi7717, pi7718, pi7719, pi7720, pi7721,
    pi7722, pi7723, pi7724, pi7725, pi7726, pi7727, pi7728, pi7729, pi7730,
    pi7731, pi7732, pi7733, pi7734, pi7735, pi7736, pi7737, pi7738, pi7739,
    pi7740, pi7741, pi7742, pi7743, pi7744, pi7745, pi7746, pi7747, pi7748,
    pi7749, pi7750, pi7751, pi7752, pi7753, pi7754, pi7755, pi7756, pi7757,
    pi7758, pi7759, pi7760, pi7761, pi7762, pi7763, pi7764, pi7765, pi7766,
    pi7767, pi7768, pi7769, pi7770, pi7771, pi7772, pi7773, pi7774, pi7775,
    pi7776, pi7777, pi7778, pi7779, pi7780, pi7781, pi7782, pi7783, pi7784,
    pi7785, pi7786, pi7787, pi7788, pi7789, pi7790, pi7791, pi7792, pi7793,
    pi7794, pi7795, pi7796, pi7797, pi7798, pi7799, pi7800, pi7801, pi7802,
    pi7803, pi7804, pi7805, pi7806, pi7807, pi7808, pi7809, pi7810, pi7811,
    pi7812, pi7813, pi7814, pi7815, pi7816, pi7817, pi7818, pi7819, pi7820,
    pi7821, pi7822, pi7823, pi7824, pi7825, pi7826, pi7827, pi7828, pi7829,
    pi7830, pi7831, pi7832, pi7833, pi7834, pi7835, pi7836, pi7837, pi7838,
    pi7839, pi7840, pi7841, pi7842, pi7843, pi7844, pi7845, pi7846, pi7847,
    pi7848, pi7849, pi7850, pi7851, pi7852, pi7853, pi7854, pi7855, pi7856,
    pi7857, pi7858, pi7859, pi7860, pi7861, pi7862, pi7863, pi7864, pi7865,
    pi7866, pi7867, pi7868, pi7869, pi7870, pi7871, pi7872, pi7873, pi7874,
    pi7875, pi7876, pi7877, pi7878, pi7879, pi7880, pi7881, pi7882, pi7883,
    pi7884, pi7885, pi7886, pi7887, pi7888, pi7889, pi7890, pi7891, pi7892,
    pi7893, pi7894, pi7895, pi7896, pi7897, pi7898, pi7899, pi7900, pi7901,
    pi7902, pi7903, pi7904, pi7905, pi7906, pi7907, pi7908, pi7909, pi7910,
    pi7911, pi7912, pi7913, pi7914, pi7915, pi7916, pi7917, pi7918, pi7919,
    pi7920, pi7921, pi7922, pi7923, pi7924, pi7925, pi7926, pi7927, pi7928,
    pi7929, pi7930, pi7931, pi7932, pi7933, pi7934, pi7935, pi7936, pi7937,
    pi7938, pi7939, pi7940, pi7941, pi7942, pi7943, pi7944, pi7945, pi7946,
    pi7947, pi7948, pi7949, pi7950, pi7951, pi7952, pi7953, pi7954, pi7955,
    pi7956, pi7957, pi7958, pi7959, pi7960, pi7961, pi7962, pi7963, pi7964,
    pi7965, pi7966, pi7967, pi7968, pi7969, pi7970, pi7971, pi7972, pi7973,
    pi7974, pi7975, pi7976, pi7977, pi7978, pi7979, pi7980, pi7981, pi7982,
    pi7983, pi7984, pi7985, pi7986, pi7987, pi7988, pi7989, pi7990, pi7991,
    pi7992, pi7993, pi7994, pi7995, pi7996, pi7997, pi7998, pi7999, pi8000,
    pi8001, pi8002, pi8003, pi8004, pi8005, pi8006, pi8007, pi8008, pi8009,
    pi8010, pi8011, pi8012, pi8013, pi8014, pi8015, pi8016, pi8017, pi8018,
    pi8019, pi8020, pi8021, pi8022, pi8023, pi8024, pi8025, pi8026, pi8027,
    pi8028, pi8029, pi8030, pi8031, pi8032, pi8033, pi8034, pi8035, pi8036,
    pi8037, pi8038, pi8039, pi8040, pi8041, pi8042, pi8043, pi8044, pi8045,
    pi8046, pi8047, pi8048, pi8049, pi8050, pi8051, pi8052, pi8053, pi8054,
    pi8055, pi8056, pi8057, pi8058, pi8059, pi8060, pi8061, pi8062, pi8063,
    pi8064, pi8065, pi8066, pi8067, pi8068, pi8069, pi8070, pi8071, pi8072,
    pi8073, pi8074, pi8075, pi8076, pi8077, pi8078, pi8079, pi8080, pi8081,
    pi8082, pi8083, pi8084, pi8085, pi8086, pi8087, pi8088, pi8089, pi8090,
    pi8091, pi8092, pi8093, pi8094, pi8095, pi8096, pi8097, pi8098, pi8099,
    pi8100, pi8101, pi8102, pi8103, pi8104, pi8105, pi8106, pi8107, pi8108,
    pi8109, pi8110, pi8111, pi8112, pi8113, pi8114, pi8115, pi8116, pi8117,
    pi8118, pi8119, pi8120, pi8121, pi8122, pi8123, pi8124, pi8125, pi8126,
    pi8127, pi8128, pi8129, pi8130, pi8131, pi8132, pi8133, pi8134, pi8135,
    pi8136, pi8137, pi8138, pi8139, pi8140, pi8141, pi8142, pi8143, pi8144,
    pi8145, pi8146, pi8147, pi8148, pi8149, pi8150, pi8151, pi8152, pi8153,
    pi8154, pi8155, pi8156, pi8157, pi8158, pi8159, pi8160, pi8161, pi8162,
    pi8163, pi8164, pi8165, pi8166, pi8167, pi8168, pi8169, pi8170, pi8171,
    pi8172, pi8173, pi8174, pi8175, pi8176, pi8177, pi8178, pi8179, pi8180,
    pi8181, pi8182, pi8183, pi8184, pi8185, pi8186, pi8187, pi8188, pi8189,
    pi8190, pi8191, pi8192, pi8193, pi8194, pi8195, pi8196, pi8197, pi8198,
    pi8199, pi8200, pi8201, pi8202, pi8203, pi8204, pi8205, pi8206, pi8207,
    pi8208, pi8209, pi8210, pi8211, pi8212, pi8213, pi8214, pi8215, pi8216,
    pi8217, pi8218, pi8219, pi8220, pi8221, pi8222, pi8223, pi8224, pi8225,
    pi8226, pi8227, pi8228, pi8229, pi8230, pi8231, pi8232, pi8233, pi8234,
    pi8235, pi8236, pi8237, pi8238, pi8239, pi8240, pi8241, pi8242, pi8243,
    pi8244, pi8245, pi8246, pi8247, pi8248, pi8249, pi8250, pi8251, pi8252,
    pi8253, pi8254, pi8255, pi8256, pi8257, pi8258, pi8259, pi8260, pi8261,
    pi8262, pi8263, pi8264, pi8265, pi8266, pi8267, pi8268, pi8269, pi8270,
    pi8271, pi8272, pi8273, pi8274, pi8275, pi8276, pi8277, pi8278, pi8279,
    pi8280, pi8281, pi8282, pi8283, pi8284, pi8285, pi8286, pi8287, pi8288,
    pi8289, pi8290, pi8291, pi8292, pi8293, pi8294, pi8295, pi8296, pi8297,
    pi8298, pi8299, pi8300, pi8301, pi8302, pi8303, pi8304, pi8305, pi8306,
    pi8307, pi8308, pi8309, pi8310, pi8311, pi8312, pi8313, pi8314, pi8315,
    pi8316, pi8317, pi8318, pi8319, pi8320, pi8321, pi8322, pi8323, pi8324,
    pi8325, pi8326, pi8327, pi8328, pi8329, pi8330, pi8331, pi8332, pi8333,
    pi8334, pi8335, pi8336, pi8337, pi8338, pi8339, pi8340, pi8341, pi8342,
    pi8343, pi8344, pi8345, pi8346, pi8347, pi8348, pi8349, pi8350, pi8351,
    pi8352, pi8353, pi8354, pi8355, pi8356, pi8357, pi8358, pi8359, pi8360,
    pi8361, pi8362, pi8363, pi8364, pi8365, pi8366, pi8367, pi8368, pi8369,
    pi8370, pi8371, pi8372, pi8373, pi8374, pi8375, pi8376, pi8377, pi8378,
    pi8379, pi8380, pi8381, pi8382, pi8383, pi8384, pi8385, pi8386, pi8387,
    pi8388, pi8389, pi8390, pi8391, pi8392, pi8393, pi8394, pi8395, pi8396,
    pi8397, pi8398, pi8399, pi8400, pi8401, pi8402, pi8403, pi8404, pi8405,
    pi8406, pi8407, pi8408, pi8409, pi8410, pi8411, pi8412, pi8413, pi8414,
    pi8415, pi8416, pi8417, pi8418, pi8419, pi8420, pi8421, pi8422, pi8423,
    pi8424, pi8425, pi8426, pi8427, pi8428, pi8429, pi8430, pi8431, pi8432,
    pi8433, pi8434, pi8435, pi8436, pi8437, pi8438, pi8439, pi8440, pi8441,
    pi8442, pi8443, pi8444, pi8445, pi8446, pi8447, pi8448, pi8449, pi8450,
    pi8451, pi8452, pi8453, pi8454, pi8455, pi8456, pi8457, pi8458, pi8459,
    pi8460, pi8461, pi8462, pi8463, pi8464, pi8465, pi8466, pi8467, pi8468,
    pi8469, pi8470, pi8471, pi8472, pi8473, pi8474, pi8475, pi8476, pi8477,
    pi8478, pi8479, pi8480, pi8481, pi8482, pi8483, pi8484, pi8485, pi8486,
    pi8487, pi8488, pi8489, pi8490, pi8491, pi8492, pi8493, pi8494, pi8495,
    pi8496, pi8497, pi8498, pi8499, pi8500, pi8501, pi8502, pi8503, pi8504,
    pi8505, pi8506, pi8507, pi8508, pi8509, pi8510, pi8511, pi8512, pi8513,
    pi8514, pi8515, pi8516, pi8517, pi8518, pi8519, pi8520, pi8521, pi8522,
    pi8523, pi8524, pi8525, pi8526, pi8527, pi8528, pi8529, pi8530, pi8531,
    pi8532, pi8533, pi8534, pi8535, pi8536, pi8537, pi8538, pi8539, pi8540,
    pi8541, pi8542, pi8543, pi8544, pi8545, pi8546, pi8547, pi8548, pi8549,
    pi8550, pi8551, pi8552, pi8553, pi8554, pi8555, pi8556, pi8557, pi8558,
    pi8559, pi8560, pi8561, pi8562, pi8563, pi8564, pi8565, pi8566, pi8567,
    pi8568, pi8569, pi8570, pi8571, pi8572, pi8573, pi8574, pi8575, pi8576,
    pi8577, pi8578, pi8579, pi8580, pi8581, pi8582, pi8583, pi8584, pi8585,
    pi8586, pi8587, pi8588, pi8589, pi8590, pi8591, pi8592, pi8593, pi8594,
    pi8595, pi8596, pi8597, pi8598, pi8599, pi8600, pi8601, pi8602, pi8603,
    pi8604, pi8605, pi8606, pi8607, pi8608, pi8609, pi8610, pi8611, pi8612,
    pi8613, pi8614, pi8615, pi8616, pi8617, pi8618, pi8619, pi8620, pi8621,
    pi8622, pi8623, pi8624, pi8625, pi8626, pi8627, pi8628, pi8629, pi8630,
    pi8631, pi8632, pi8633, pi8634, pi8635, pi8636, pi8637, pi8638, pi8639,
    pi8640, pi8641, pi8642, pi8643, pi8644, pi8645, pi8646, pi8647, pi8648,
    pi8649, pi8650, pi8651, pi8652, pi8653, pi8654, pi8655, pi8656, pi8657,
    pi8658, pi8659, pi8660, pi8661, pi8662, pi8663, pi8664, pi8665, pi8666,
    pi8667, pi8668, pi8669, pi8670, pi8671, pi8672, pi8673, pi8674, pi8675,
    pi8676, pi8677, pi8678, pi8679, pi8680, pi8681, pi8682, pi8683, pi8684,
    pi8685, pi8686, pi8687, pi8688, pi8689, pi8690, pi8691, pi8692, pi8693,
    pi8694, pi8695, pi8696, pi8697, pi8698, pi8699, pi8700, pi8701, pi8702,
    pi8703, pi8704, pi8705, pi8706, pi8707, pi8708, pi8709, pi8710, pi8711,
    pi8712, pi8713, pi8714, pi8715, pi8716, pi8717, pi8718, pi8719, pi8720,
    pi8721, pi8722, pi8723, pi8724, pi8725, pi8726, pi8727, pi8728, pi8729,
    pi8730, pi8731, pi8732, pi8733, pi8734, pi8735, pi8736, pi8737, pi8738,
    pi8739, pi8740, pi8741, pi8742, pi8743, pi8744, pi8745, pi8746, pi8747,
    pi8748, pi8749, pi8750, pi8751, pi8752, pi8753, pi8754, pi8755, pi8756,
    pi8757, pi8758, pi8759, pi8760, pi8761, pi8762, pi8763, pi8764, pi8765,
    pi8766, pi8767, pi8768, pi8769, pi8770, pi8771, pi8772, pi8773, pi8774,
    pi8775, pi8776, pi8777, pi8778, pi8779, pi8780, pi8781, pi8782, pi8783,
    pi8784, pi8785, pi8786, pi8787, pi8788, pi8789, pi8790, pi8791, pi8792,
    pi8793, pi8794, pi8795, pi8796, pi8797, pi8798, pi8799, pi8800, pi8801,
    pi8802, pi8803, pi8804, pi8805, pi8806, pi8807, pi8808, pi8809, pi8810,
    pi8811, pi8812, pi8813, pi8814, pi8815, pi8816, pi8817, pi8818, pi8819,
    pi8820, pi8821, pi8822, pi8823, pi8824, pi8825, pi8826, pi8827, pi8828,
    pi8829, pi8830, pi8831, pi8832, pi8833, pi8834, pi8835, pi8836, pi8837,
    pi8838, pi8839, pi8840, pi8841, pi8842, pi8843, pi8844, pi8845, pi8846,
    pi8847, pi8848, pi8849, pi8850, pi8851, pi8852, pi8853, pi8854, pi8855,
    pi8856, pi8857, pi8858, pi8859, pi8860, pi8861, pi8862, pi8863, pi8864,
    pi8865, pi8866, pi8867, pi8868, pi8869, pi8870, pi8871, pi8872, pi8873,
    pi8874, pi8875, pi8876, pi8877, pi8878, pi8879, pi8880, pi8881, pi8882,
    pi8883, pi8884, pi8885, pi8886, pi8887, pi8888, pi8889, pi8890, pi8891,
    pi8892, pi8893, pi8894, pi8895, pi8896, pi8897, pi8898, pi8899, pi8900,
    pi8901, pi8902, pi8903, pi8904, pi8905, pi8906, pi8907, pi8908, pi8909,
    pi8910, pi8911, pi8912, pi8913, pi8914, pi8915, pi8916, pi8917, pi8918,
    pi8919, pi8920, pi8921, pi8922, pi8923, pi8924, pi8925, pi8926, pi8927,
    pi8928, pi8929, pi8930, pi8931, pi8932, pi8933, pi8934, pi8935, pi8936,
    pi8937, pi8938, pi8939, pi8940, pi8941, pi8942, pi8943, pi8944, pi8945,
    pi8946, pi8947, pi8948, pi8949, pi8950, pi8951, pi8952, pi8953, pi8954,
    pi8955, pi8956, pi8957, pi8958, pi8959, pi8960, pi8961, pi8962, pi8963,
    pi8964, pi8965, pi8966, pi8967, pi8968, pi8969, pi8970, pi8971, pi8972,
    pi8973, pi8974, pi8975, pi8976, pi8977, pi8978, pi8979, pi8980, pi8981,
    pi8982, pi8983, pi8984, pi8985, pi8986, pi8987, pi8988, pi8989, pi8990,
    pi8991, pi8992, pi8993, pi8994, pi8995, pi8996, pi8997, pi8998, pi8999,
    pi9000, pi9001, pi9002, pi9003, pi9004, pi9005, pi9006, pi9007, pi9008,
    pi9009, pi9010, pi9011, pi9012, pi9013, pi9014, pi9015, pi9016, pi9017,
    pi9018, pi9019, pi9020, pi9021, pi9022, pi9023, pi9024, pi9025, pi9026,
    pi9027, pi9028, pi9029, pi9030, pi9031, pi9032, pi9033, pi9034, pi9035,
    pi9036, pi9037, pi9038, pi9039, pi9040, pi9041,
    po0000, po0001, po0002, po0003, po0004, po0005, po0006, po0007, po0008,
    po0009, po0010, po0011, po0012, po0013, po0014, po0015, po0016, po0017,
    po0018, po0019, po0020, po0021, po0022, po0023, po0024, po0025, po0026,
    po0027, po0028, po0029, po0030, po0031, po0032, po0033, po0034, po0035,
    po0036, po0037, po0038, po0039, po0040, po0041, po0042, po0043, po0044,
    po0045, po0046, po0047, po0048, po0049, po0050, po0051, po0052, po0053,
    po0054, po0055, po0056, po0057, po0058, po0059, po0060, po0061, po0062,
    po0063, po0064, po0065, po0066, po0067, po0068, po0069, po0070, po0071,
    po0072, po0073, po0074, po0075, po0076, po0077, po0078, po0079, po0080,
    po0081, po0082, po0083, po0084, po0085, po0086, po0087, po0088, po0089,
    po0090, po0091, po0092, po0093, po0094, po0095, po0096, po0097, po0098,
    po0099, po0100, po0101, po0102, po0103, po0104, po0105, po0106, po0107,
    po0108, po0109, po0110, po0111, po0112, po0113, po0114, po0115, po0116,
    po0117, po0118, po0119, po0120, po0121, po0122, po0123, po0124, po0125,
    po0126, po0127, po0128, po0129, po0130, po0131, po0132, po0133, po0134,
    po0135, po0136, po0137, po0138, po0139, po0140, po0141, po0142, po0143,
    po0144, po0145, po0146, po0147, po0148, po0149, po0150, po0151, po0152,
    po0153, po0154, po0155, po0156, po0157, po0158, po0159, po0160, po0161,
    po0162, po0163, po0164, po0165, po0166, po0167, po0168, po0169, po0170,
    po0171, po0172, po0173, po0174, po0175, po0176, po0177, po0178, po0179,
    po0180, po0181, po0182, po0183, po0184, po0185, po0186, po0187, po0188,
    po0189, po0190, po0191, po0192, po0193, po0194, po0195, po0196, po0197,
    po0198, po0199, po0200, po0201, po0202, po0203, po0204, po0205, po0206,
    po0207, po0208, po0209, po0210, po0211, po0212, po0213, po0214, po0215,
    po0216, po0217, po0218, po0219, po0220, po0221, po0222, po0223, po0224,
    po0225, po0226, po0227, po0228, po0229, po0230, po0231, po0232, po0233,
    po0234, po0235, po0236, po0237, po0238, po0239, po0240, po0241, po0242,
    po0243, po0244, po0245, po0246, po0247, po0248, po0249, po0250, po0251,
    po0252, po0253, po0254, po0255, po0256, po0257, po0258, po0259, po0260,
    po0261, po0262, po0263, po0264, po0265, po0266, po0267, po0268, po0269,
    po0270, po0271, po0272, po0273, po0274, po0275, po0276, po0277, po0278,
    po0279, po0280, po0281, po0282, po0283, po0284, po0285, po0286, po0287,
    po0288, po0289, po0290, po0291, po0292, po0293, po0294, po0295, po0296,
    po0297, po0298, po0299, po0300, po0301, po0302, po0303, po0304, po0305,
    po0306, po0307, po0308, po0309, po0310, po0311, po0312, po0313, po0314,
    po0315, po0316, po0317, po0318, po0319, po0320, po0321, po0322, po0323,
    po0324, po0325, po0326, po0327, po0328, po0329, po0330, po0331, po0332,
    po0333, po0334, po0335, po0336, po0337, po0338, po0339, po0340, po0341,
    po0342, po0343, po0344, po0345, po0346, po0347, po0348, po0349, po0350,
    po0351, po0352, po0353, po0354, po0355, po0356, po0357, po0358, po0359,
    po0360, po0361, po0362, po0363, po0364, po0365, po0366, po0367, po0368,
    po0369, po0370, po0371, po0372, po0373, po0374, po0375, po0376, po0377,
    po0378, po0379, po0380, po0381, po0382, po0383, po0384, po0385, po0386,
    po0387, po0388, po0389, po0390, po0391, po0392, po0393, po0394, po0395,
    po0396, po0397, po0398, po0399, po0400, po0401, po0402, po0403, po0404,
    po0405, po0406, po0407, po0408, po0409, po0410, po0411, po0412, po0413,
    po0414, po0415, po0416, po0417, po0418, po0419, po0420, po0421, po0422,
    po0423, po0424, po0425, po0426, po0427, po0428, po0429, po0430, po0431,
    po0432, po0433, po0434, po0435, po0436, po0437, po0438, po0439, po0440,
    po0441, po0442, po0443, po0444, po0445, po0446, po0447, po0448, po0449,
    po0450, po0451, po0452, po0453, po0454, po0455, po0456, po0457, po0458,
    po0459, po0460, po0461, po0462, po0463, po0464, po0465, po0466, po0467,
    po0468, po0469, po0470, po0471, po0472, po0473, po0474, po0475, po0476,
    po0477, po0478, po0479, po0480, po0481, po0482, po0483, po0484, po0485,
    po0486, po0487, po0488, po0489, po0490, po0491, po0492, po0493, po0494,
    po0495, po0496, po0497, po0498, po0499, po0500, po0501, po0502, po0503,
    po0504, po0505, po0506, po0507, po0508, po0509, po0510, po0511, po0512,
    po0513, po0514, po0515, po0516, po0517, po0518, po0519, po0520, po0521,
    po0522, po0523, po0524, po0525, po0526, po0527, po0528, po0529, po0530,
    po0531, po0532, po0533, po0534, po0535, po0536, po0537, po0538, po0539,
    po0540, po0541, po0542, po0543, po0544, po0545, po0546, po0547, po0548,
    po0549, po0550, po0551, po0552, po0553, po0554, po0555, po0556, po0557,
    po0558, po0559, po0560, po0561, po0562, po0563, po0564, po0565, po0566,
    po0567, po0568, po0569, po0570, po0571, po0572, po0573, po0574, po0575,
    po0576, po0577, po0578, po0579, po0580, po0581, po0582, po0583, po0584,
    po0585, po0586, po0587, po0588, po0589, po0590, po0591, po0592, po0593,
    po0594, po0595, po0596, po0597, po0598, po0599, po0600, po0601, po0602,
    po0603, po0604, po0605, po0606, po0607, po0608, po0609, po0610, po0611,
    po0612, po0613, po0614, po0615, po0616, po0617, po0618, po0619, po0620,
    po0621, po0622, po0623, po0624, po0625, po0626, po0627, po0628, po0629,
    po0630, po0631, po0632, po0633, po0634, po0635, po0636, po0637, po0638,
    po0639, po0640, po0641, po0642, po0643, po0644, po0645, po0646, po0647,
    po0648, po0649, po0650, po0651, po0652, po0653, po0654, po0655, po0656,
    po0657, po0658, po0659, po0660, po0661, po0662, po0663, po0664, po0665,
    po0666, po0667, po0668, po0669, po0670, po0671, po0672, po0673, po0674,
    po0675, po0676, po0677, po0678, po0679, po0680, po0681, po0682, po0683,
    po0684, po0685, po0686, po0687, po0688, po0689, po0690, po0691, po0692,
    po0693, po0694, po0695, po0696, po0697, po0698, po0699, po0700, po0701,
    po0702, po0703, po0704, po0705, po0706, po0707, po0708, po0709, po0710,
    po0711, po0712, po0713, po0714, po0715, po0716, po0717, po0718, po0719,
    po0720, po0721, po0722, po0723, po0724, po0725, po0726, po0727, po0728,
    po0729, po0730, po0731, po0732, po0733, po0734, po0735, po0736, po0737,
    po0738, po0739, po0740, po0741, po0742, po0743, po0744, po0745, po0746,
    po0747, po0748, po0749, po0750, po0751, po0752, po0753, po0754, po0755,
    po0756, po0757, po0758, po0759, po0760, po0761, po0762, po0763, po0764,
    po0765, po0766, po0767, po0768, po0769, po0770, po0771, po0772, po0773,
    po0774, po0775, po0776, po0777, po0778, po0779, po0780, po0781, po0782,
    po0783, po0784, po0785, po0786, po0787, po0788, po0789, po0790, po0791,
    po0792, po0793, po0794, po0795, po0796, po0797, po0798, po0799, po0800,
    po0801, po0802, po0803, po0804, po0805, po0806, po0807, po0808, po0809,
    po0810, po0811, po0812, po0813, po0814, po0815, po0816, po0817, po0818,
    po0819, po0820, po0821, po0822, po0823, po0824, po0825, po0826, po0827,
    po0828, po0829, po0830, po0831, po0832, po0833, po0834, po0835, po0836,
    po0837, po0838, po0839, po0840, po0841, po0842, po0843, po0844, po0845,
    po0846, po0847, po0848, po0849, po0850, po0851, po0852, po0853, po0854,
    po0855, po0856, po0857, po0858, po0859, po0860, po0861, po0862, po0863,
    po0864, po0865, po0866, po0867, po0868, po0869, po0870, po0871, po0872,
    po0873, po0874, po0875, po0876, po0877, po0878, po0879, po0880, po0881,
    po0882, po0883, po0884, po0885, po0886, po0887, po0888, po0889, po0890,
    po0891, po0892, po0893, po0894, po0895, po0896, po0897, po0898, po0899,
    po0900, po0901, po0902, po0903, po0904, po0905, po0906, po0907, po0908,
    po0909, po0910, po0911, po0912, po0913, po0914, po0915, po0916, po0917,
    po0918, po0919, po0920, po0921, po0922, po0923, po0924, po0925, po0926,
    po0927, po0928, po0929, po0930, po0931, po0932, po0933, po0934, po0935,
    po0936, po0937, po0938, po0939, po0940, po0941, po0942, po0943, po0944,
    po0945, po0946, po0947, po0948, po0949, po0950, po0951, po0952, po0953,
    po0954, po0955, po0956, po0957, po0958, po0959, po0960, po0961, po0962,
    po0963, po0964, po0965, po0966, po0967, po0968, po0969, po0970, po0971,
    po0972, po0973, po0974, po0975, po0976, po0977, po0978, po0979, po0980,
    po0981, po0982, po0983, po0984, po0985, po0986, po0987, po0988, po0989,
    po0990, po0991, po0992, po0993, po0994, po0995, po0996, po0997, po0998,
    po0999, po1000, po1001, po1002, po1003, po1004, po1005, po1006, po1007,
    po1008, po1009, po1010, po1011, po1012, po1013, po1014, po1015, po1016,
    po1017, po1018, po1019, po1020, po1021, po1022, po1023, po1024, po1025,
    po1026, po1027, po1028, po1029, po1030, po1031, po1032, po1033, po1034,
    po1035, po1036, po1037, po1038, po1039, po1040, po1041, po1042, po1043,
    po1044, po1045, po1046, po1047, po1048, po1049, po1050, po1051, po1052,
    po1053, po1054, po1055, po1056, po1057, po1058, po1059, po1060, po1061,
    po1062, po1063, po1064, po1065, po1066, po1067, po1068, po1069, po1070,
    po1071, po1072, po1073, po1074, po1075, po1076, po1077, po1078, po1079,
    po1080, po1081, po1082, po1083, po1084, po1085, po1086, po1087, po1088,
    po1089, po1090, po1091, po1092, po1093, po1094, po1095, po1096, po1097,
    po1098, po1099, po1100, po1101, po1102, po1103, po1104, po1105, po1106,
    po1107, po1108, po1109, po1110, po1111, po1112, po1113, po1114, po1115,
    po1116, po1117, po1118, po1119, po1120, po1121, po1122, po1123, po1124,
    po1125, po1126, po1127, po1128, po1129, po1130, po1131, po1132, po1133,
    po1134, po1135, po1136, po1137, po1138, po1139, po1140, po1141, po1142,
    po1143, po1144, po1145, po1146, po1147, po1148, po1149, po1150, po1151,
    po1152, po1153, po1154, po1155, po1156, po1157, po1158, po1159, po1160,
    po1161, po1162, po1163, po1164, po1165, po1166, po1167, po1168, po1169,
    po1170, po1171, po1172, po1173, po1174, po1175, po1176, po1177, po1178,
    po1179, po1180, po1181, po1182, po1183, po1184, po1185, po1186, po1187,
    po1188, po1189, po1190, po1191, po1192, po1193, po1194, po1195, po1196,
    po1197, po1198, po1199, po1200, po1201, po1202, po1203, po1204, po1205,
    po1206, po1207, po1208, po1209, po1210, po1211, po1212, po1213, po1214,
    po1215, po1216, po1217, po1218, po1219, po1220, po1221, po1222, po1223,
    po1224, po1225, po1226, po1227, po1228, po1229, po1230, po1231, po1232,
    po1233, po1234, po1235, po1236, po1237, po1238, po1239, po1240, po1241,
    po1242, po1243, po1244, po1245, po1246, po1247, po1248, po1249, po1250,
    po1251, po1252, po1253, po1254, po1255, po1256, po1257, po1258, po1259,
    po1260, po1261, po1262, po1263, po1264, po1265, po1266, po1267, po1268,
    po1269, po1270, po1271, po1272, po1273, po1274, po1275, po1276, po1277,
    po1278, po1279, po1280, po1281, po1282, po1283, po1284, po1285, po1286,
    po1287, po1288, po1289, po1290, po1291, po1292, po1293, po1294, po1295,
    po1296, po1297, po1298, po1299, po1300, po1301, po1302, po1303, po1304,
    po1305, po1306, po1307, po1308, po1309, po1310, po1311, po1312, po1313,
    po1314, po1315, po1316, po1317, po1318, po1319, po1320, po1321, po1322,
    po1323, po1324, po1325, po1326, po1327, po1328, po1329, po1330, po1331,
    po1332, po1333, po1334, po1335, po1336, po1337, po1338, po1339, po1340,
    po1341, po1342, po1343, po1344, po1345, po1346, po1347, po1348, po1349,
    po1350, po1351, po1352, po1353, po1354, po1355, po1356, po1357, po1358,
    po1359, po1360, po1361, po1362, po1363, po1364, po1365, po1366, po1367,
    po1368, po1369, po1370, po1371, po1372, po1373, po1374, po1375, po1376,
    po1377, po1378, po1379, po1380, po1381, po1382, po1383, po1384, po1385,
    po1386, po1387, po1388, po1389, po1390, po1391, po1392, po1393, po1394,
    po1395, po1396, po1397, po1398, po1399, po1400, po1401, po1402, po1403,
    po1404, po1405, po1406, po1407, po1408, po1409, po1410, po1411, po1412,
    po1413, po1414, po1415, po1416, po1417, po1418, po1419, po1420, po1421,
    po1422, po1423, po1424, po1425, po1426, po1427, po1428, po1429, po1430,
    po1431, po1432, po1433, po1434, po1435, po1436, po1437, po1438, po1439,
    po1440, po1441, po1442, po1443, po1444, po1445, po1446, po1447, po1448,
    po1449, po1450, po1451, po1452, po1453, po1454, po1455, po1456, po1457,
    po1458, po1459, po1460, po1461, po1462, po1463, po1464, po1465, po1466,
    po1467, po1468, po1469, po1470, po1471, po1472, po1473, po1474, po1475,
    po1476, po1477, po1478, po1479, po1480, po1481, po1482, po1483, po1484,
    po1485, po1486, po1487, po1488, po1489, po1490, po1491, po1492, po1493,
    po1494, po1495, po1496, po1497, po1498, po1499, po1500, po1501, po1502,
    po1503, po1504, po1505, po1506, po1507, po1508, po1509, po1510, po1511,
    po1512, po1513, po1514, po1515, po1516, po1517, po1518, po1519, po1520,
    po1521, po1522, po1523, po1524, po1525, po1526, po1527, po1528, po1529,
    po1530, po1531, po1532, po1533, po1534, po1535, po1536, po1537, po1538,
    po1539, po1540, po1541, po1542, po1543, po1544, po1545, po1546, po1547,
    po1548, po1549, po1550, po1551, po1552, po1553, po1554, po1555, po1556,
    po1557, po1558, po1559, po1560, po1561, po1562, po1563, po1564, po1565,
    po1566, po1567, po1568, po1569, po1570, po1571, po1572, po1573, po1574,
    po1575, po1576, po1577, po1578, po1579, po1580, po1581, po1582, po1583,
    po1584, po1585, po1586, po1587, po1588, po1589, po1590, po1591, po1592,
    po1593, po1594, po1595, po1596, po1597, po1598, po1599, po1600, po1601,
    po1602, po1603, po1604, po1605, po1606, po1607, po1608, po1609, po1610,
    po1611, po1612, po1613, po1614, po1615, po1616, po1617, po1618, po1619,
    po1620, po1621, po1622, po1623, po1624, po1625, po1626, po1627, po1628,
    po1629, po1630, po1631, po1632, po1633, po1634, po1635, po1636, po1637,
    po1638, po1639, po1640, po1641, po1642, po1643, po1644, po1645, po1646,
    po1647, po1648, po1649, po1650, po1651, po1652, po1653, po1654, po1655,
    po1656, po1657, po1658, po1659, po1660, po1661, po1662, po1663, po1664,
    po1665, po1666, po1667, po1668, po1669, po1670, po1671, po1672, po1673,
    po1674, po1675, po1676, po1677, po1678, po1679, po1680, po1681, po1682,
    po1683, po1684, po1685, po1686, po1687, po1688, po1689, po1690, po1691,
    po1692, po1693, po1694, po1695, po1696, po1697, po1698, po1699, po1700,
    po1701, po1702, po1703, po1704, po1705, po1706, po1707, po1708, po1709,
    po1710, po1711, po1712, po1713, po1714, po1715, po1716, po1717, po1718,
    po1719, po1720, po1721, po1722, po1723, po1724, po1725, po1726, po1727,
    po1728, po1729, po1730, po1731, po1732, po1733, po1734, po1735, po1736,
    po1737, po1738, po1739, po1740, po1741, po1742, po1743, po1744, po1745,
    po1746, po1747, po1748, po1749, po1750, po1751, po1752, po1753, po1754,
    po1755, po1756, po1757, po1758, po1759, po1760, po1761, po1762, po1763,
    po1764, po1765, po1766, po1767, po1768, po1769, po1770, po1771, po1772,
    po1773, po1774, po1775, po1776, po1777, po1778, po1779, po1780, po1781,
    po1782, po1783, po1784, po1785, po1786, po1787, po1788, po1789, po1790,
    po1791, po1792, po1793, po1794, po1795, po1796, po1797, po1798, po1799,
    po1800, po1801, po1802, po1803, po1804, po1805, po1806, po1807, po1808,
    po1809, po1810, po1811, po1812, po1813, po1814, po1815, po1816, po1817,
    po1818, po1819, po1820, po1821, po1822, po1823, po1824, po1825, po1826,
    po1827, po1828, po1829, po1830, po1831, po1832, po1833, po1834, po1835,
    po1836, po1837, po1838, po1839, po1840, po1841, po1842, po1843, po1844,
    po1845, po1846, po1847, po1848, po1849, po1850, po1851, po1852, po1853,
    po1854, po1855, po1856, po1857, po1858, po1859, po1860, po1861, po1862,
    po1863, po1864, po1865, po1866, po1867, po1868, po1869, po1870, po1871,
    po1872, po1873, po1874, po1875, po1876, po1877, po1878, po1879, po1880,
    po1881, po1882, po1883, po1884, po1885, po1886, po1887, po1888, po1889,
    po1890, po1891, po1892, po1893, po1894, po1895, po1896, po1897, po1898,
    po1899, po1900, po1901, po1902, po1903, po1904, po1905, po1906, po1907,
    po1908, po1909, po1910, po1911, po1912, po1913, po1914, po1915, po1916,
    po1917, po1918, po1919, po1920, po1921, po1922, po1923, po1924, po1925,
    po1926, po1927, po1928, po1929, po1930, po1931, po1932, po1933, po1934,
    po1935, po1936, po1937, po1938, po1939, po1940, po1941, po1942, po1943,
    po1944, po1945, po1946, po1947, po1948, po1949, po1950, po1951, po1952,
    po1953, po1954, po1955, po1956, po1957, po1958, po1959, po1960, po1961,
    po1962, po1963, po1964, po1965, po1966, po1967, po1968, po1969, po1970,
    po1971, po1972, po1973, po1974, po1975, po1976, po1977, po1978, po1979,
    po1980, po1981, po1982, po1983, po1984, po1985, po1986, po1987, po1988,
    po1989, po1990, po1991, po1992, po1993, po1994, po1995, po1996, po1997,
    po1998, po1999, po2000, po2001, po2002, po2003, po2004, po2005, po2006,
    po2007, po2008, po2009, po2010, po2011, po2012, po2013, po2014, po2015,
    po2016, po2017, po2018, po2019, po2020, po2021, po2022, po2023, po2024,
    po2025, po2026, po2027, po2028, po2029, po2030, po2031, po2032, po2033,
    po2034, po2035, po2036, po2037, po2038, po2039, po2040, po2041, po2042,
    po2043, po2044, po2045, po2046, po2047, po2048, po2049, po2050, po2051,
    po2052, po2053, po2054, po2055, po2056, po2057, po2058, po2059, po2060,
    po2061, po2062, po2063, po2064, po2065, po2066, po2067, po2068, po2069,
    po2070, po2071, po2072, po2073, po2074, po2075, po2076, po2077, po2078,
    po2079, po2080, po2081, po2082, po2083, po2084, po2085, po2086, po2087,
    po2088, po2089, po2090, po2091, po2092, po2093, po2094, po2095, po2096,
    po2097, po2098, po2099, po2100, po2101, po2102, po2103, po2104, po2105,
    po2106, po2107, po2108, po2109, po2110, po2111, po2112, po2113, po2114,
    po2115, po2116, po2117, po2118, po2119, po2120, po2121, po2122, po2123,
    po2124, po2125, po2126, po2127, po2128, po2129, po2130, po2131, po2132,
    po2133, po2134, po2135, po2136, po2137, po2138, po2139, po2140, po2141,
    po2142, po2143, po2144, po2145, po2146, po2147, po2148, po2149, po2150,
    po2151, po2152, po2153, po2154, po2155, po2156, po2157, po2158, po2159,
    po2160, po2161, po2162, po2163, po2164, po2165, po2166, po2167, po2168,
    po2169, po2170, po2171, po2172, po2173, po2174, po2175, po2176, po2177,
    po2178, po2179, po2180, po2181, po2182, po2183, po2184, po2185, po2186,
    po2187, po2188, po2189, po2190, po2191, po2192, po2193, po2194, po2195,
    po2196, po2197, po2198, po2199, po2200, po2201, po2202, po2203, po2204,
    po2205, po2206, po2207, po2208, po2209, po2210, po2211, po2212, po2213,
    po2214, po2215, po2216, po2217, po2218, po2219, po2220, po2221, po2222,
    po2223, po2224, po2225, po2226, po2227, po2228, po2229, po2230, po2231,
    po2232, po2233, po2234, po2235, po2236, po2237, po2238, po2239, po2240,
    po2241, po2242, po2243, po2244, po2245, po2246, po2247, po2248, po2249,
    po2250, po2251, po2252, po2253, po2254, po2255, po2256, po2257, po2258,
    po2259, po2260, po2261, po2262, po2263, po2264, po2265, po2266, po2267,
    po2268, po2269, po2270, po2271, po2272, po2273, po2274, po2275, po2276,
    po2277, po2278, po2279, po2280, po2281, po2282, po2283, po2284, po2285,
    po2286, po2287, po2288, po2289, po2290, po2291, po2292, po2293, po2294,
    po2295, po2296, po2297, po2298, po2299, po2300, po2301, po2302, po2303,
    po2304, po2305, po2306, po2307, po2308, po2309, po2310, po2311, po2312,
    po2313, po2314, po2315, po2316, po2317, po2318, po2319, po2320, po2321,
    po2322, po2323, po2324, po2325, po2326, po2327, po2328, po2329, po2330,
    po2331, po2332, po2333, po2334, po2335, po2336, po2337, po2338, po2339,
    po2340, po2341, po2342, po2343, po2344, po2345, po2346, po2347, po2348,
    po2349, po2350, po2351, po2352, po2353, po2354, po2355, po2356, po2357,
    po2358, po2359, po2360, po2361, po2362, po2363, po2364, po2365, po2366,
    po2367, po2368, po2369, po2370, po2371, po2372, po2373, po2374, po2375,
    po2376, po2377, po2378, po2379, po2380, po2381, po2382, po2383, po2384,
    po2385, po2386, po2387, po2388, po2389, po2390, po2391, po2392, po2393,
    po2394, po2395, po2396, po2397, po2398, po2399, po2400, po2401, po2402,
    po2403, po2404, po2405, po2406, po2407, po2408, po2409, po2410, po2411,
    po2412, po2413, po2414, po2415, po2416, po2417, po2418, po2419, po2420,
    po2421, po2422, po2423, po2424, po2425, po2426, po2427, po2428, po2429,
    po2430, po2431, po2432, po2433, po2434, po2435, po2436, po2437, po2438,
    po2439, po2440, po2441, po2442, po2443, po2444, po2445, po2446, po2447,
    po2448, po2449, po2450, po2451, po2452, po2453, po2454, po2455, po2456,
    po2457, po2458, po2459, po2460, po2461, po2462, po2463, po2464, po2465,
    po2466, po2467, po2468, po2469, po2470, po2471, po2472, po2473, po2474,
    po2475, po2476, po2477, po2478, po2479, po2480, po2481, po2482, po2483,
    po2484, po2485, po2486, po2487, po2488, po2489, po2490, po2491, po2492,
    po2493, po2494, po2495, po2496, po2497, po2498, po2499, po2500, po2501,
    po2502, po2503, po2504, po2505, po2506, po2507, po2508, po2509, po2510,
    po2511, po2512, po2513, po2514, po2515, po2516, po2517, po2518, po2519,
    po2520, po2521, po2522, po2523, po2524, po2525, po2526, po2527, po2528,
    po2529, po2530, po2531, po2532, po2533, po2534, po2535, po2536, po2537,
    po2538, po2539, po2540, po2541, po2542, po2543, po2544, po2545, po2546,
    po2547, po2548, po2549, po2550, po2551, po2552, po2553, po2554, po2555,
    po2556, po2557, po2558, po2559, po2560, po2561, po2562, po2563, po2564,
    po2565, po2566, po2567, po2568, po2569, po2570, po2571, po2572, po2573,
    po2574, po2575, po2576, po2577, po2578, po2579, po2580, po2581, po2582,
    po2583, po2584, po2585, po2586, po2587, po2588, po2589, po2590, po2591,
    po2592, po2593, po2594, po2595, po2596, po2597, po2598, po2599, po2600,
    po2601, po2602, po2603, po2604, po2605, po2606, po2607, po2608, po2609,
    po2610, po2611, po2612, po2613, po2614, po2615, po2616, po2617, po2618,
    po2619, po2620, po2621, po2622, po2623, po2624, po2625, po2626, po2627,
    po2628, po2629, po2630, po2631, po2632, po2633, po2634, po2635, po2636,
    po2637, po2638, po2639, po2640, po2641, po2642, po2643, po2644, po2645,
    po2646, po2647, po2648, po2649, po2650, po2651, po2652, po2653, po2654,
    po2655, po2656, po2657, po2658, po2659, po2660, po2661, po2662, po2663,
    po2664, po2665, po2666, po2667, po2668, po2669, po2670, po2671, po2672,
    po2673, po2674, po2675, po2676, po2677, po2678, po2679, po2680, po2681,
    po2682, po2683, po2684, po2685, po2686, po2687, po2688, po2689, po2690,
    po2691, po2692, po2693, po2694, po2695, po2696, po2697, po2698, po2699,
    po2700, po2701, po2702, po2703, po2704, po2705, po2706, po2707, po2708,
    po2709, po2710, po2711, po2712, po2713, po2714, po2715, po2716, po2717,
    po2718, po2719, po2720, po2721, po2722, po2723, po2724, po2725, po2726,
    po2727, po2728, po2729, po2730, po2731, po2732, po2733, po2734, po2735,
    po2736, po2737, po2738, po2739, po2740, po2741, po2742, po2743, po2744,
    po2745, po2746, po2747, po2748, po2749, po2750, po2751, po2752, po2753,
    po2754, po2755, po2756, po2757, po2758, po2759, po2760, po2761, po2762,
    po2763, po2764, po2765, po2766, po2767, po2768, po2769, po2770, po2771,
    po2772, po2773, po2774, po2775, po2776, po2777, po2778, po2779, po2780,
    po2781, po2782, po2783, po2784, po2785, po2786, po2787, po2788, po2789,
    po2790, po2791, po2792, po2793, po2794, po2795, po2796, po2797, po2798,
    po2799, po2800, po2801, po2802, po2803, po2804, po2805, po2806, po2807,
    po2808, po2809, po2810, po2811, po2812, po2813, po2814, po2815, po2816,
    po2817, po2818, po2819, po2820, po2821, po2822, po2823, po2824, po2825,
    po2826, po2827, po2828, po2829, po2830, po2831, po2832, po2833, po2834,
    po2835, po2836, po2837, po2838, po2839, po2840, po2841, po2842, po2843,
    po2844, po2845, po2846, po2847, po2848, po2849, po2850, po2851, po2852,
    po2853, po2854, po2855, po2856, po2857, po2858, po2859, po2860, po2861,
    po2862, po2863, po2864, po2865, po2866, po2867, po2868, po2869, po2870,
    po2871, po2872, po2873, po2874, po2875, po2876, po2877, po2878, po2879,
    po2880, po2881, po2882, po2883, po2884, po2885, po2886, po2887, po2888,
    po2889, po2890, po2891, po2892, po2893, po2894, po2895, po2896, po2897,
    po2898, po2899, po2900, po2901, po2902, po2903, po2904, po2905, po2906,
    po2907, po2908, po2909, po2910, po2911, po2912, po2913, po2914, po2915,
    po2916, po2917, po2918, po2919, po2920, po2921, po2922, po2923, po2924,
    po2925, po2926, po2927, po2928, po2929, po2930, po2931, po2932, po2933,
    po2934, po2935, po2936, po2937, po2938, po2939, po2940, po2941, po2942,
    po2943, po2944, po2945, po2946, po2947, po2948, po2949, po2950, po2951,
    po2952, po2953, po2954, po2955, po2956, po2957, po2958, po2959, po2960,
    po2961, po2962, po2963, po2964, po2965, po2966, po2967, po2968, po2969,
    po2970, po2971, po2972, po2973, po2974, po2975, po2976, po2977, po2978,
    po2979, po2980, po2981, po2982, po2983, po2984, po2985, po2986, po2987,
    po2988, po2989, po2990, po2991, po2992, po2993, po2994, po2995, po2996,
    po2997, po2998, po2999, po3000, po3001, po3002, po3003, po3004, po3005,
    po3006, po3007, po3008, po3009, po3010, po3011, po3012, po3013, po3014,
    po3015, po3016, po3017, po3018, po3019, po3020, po3021, po3022, po3023,
    po3024, po3025, po3026, po3027, po3028, po3029, po3030, po3031, po3032,
    po3033, po3034, po3035, po3036, po3037, po3038, po3039, po3040, po3041,
    po3042, po3043, po3044, po3045, po3046, po3047, po3048, po3049, po3050,
    po3051, po3052, po3053, po3054, po3055, po3056, po3057, po3058, po3059,
    po3060, po3061, po3062, po3063, po3064, po3065, po3066, po3067, po3068,
    po3069, po3070, po3071, po3072, po3073, po3074, po3075, po3076, po3077,
    po3078, po3079, po3080, po3081, po3082, po3083, po3084, po3085, po3086,
    po3087, po3088, po3089, po3090, po3091, po3092, po3093, po3094, po3095,
    po3096, po3097, po3098, po3099, po3100, po3101, po3102, po3103, po3104,
    po3105, po3106, po3107, po3108, po3109, po3110, po3111, po3112, po3113,
    po3114, po3115, po3116, po3117, po3118, po3119, po3120, po3121, po3122,
    po3123, po3124, po3125, po3126, po3127, po3128, po3129, po3130, po3131,
    po3132, po3133, po3134, po3135, po3136, po3137, po3138, po3139, po3140,
    po3141, po3142, po3143, po3144, po3145, po3146, po3147, po3148, po3149,
    po3150, po3151, po3152, po3153, po3154, po3155, po3156, po3157, po3158,
    po3159, po3160, po3161, po3162, po3163, po3164, po3165, po3166, po3167,
    po3168, po3169, po3170, po3171, po3172, po3173, po3174, po3175, po3176,
    po3177, po3178, po3179, po3180, po3181, po3182, po3183, po3184, po3185,
    po3186, po3187, po3188, po3189, po3190, po3191, po3192, po3193, po3194,
    po3195, po3196, po3197, po3198, po3199, po3200, po3201, po3202, po3203,
    po3204, po3205, po3206, po3207, po3208, po3209, po3210, po3211, po3212,
    po3213, po3214, po3215, po3216, po3217, po3218, po3219, po3220, po3221,
    po3222, po3223, po3224, po3225, po3226, po3227, po3228, po3229, po3230,
    po3231, po3232, po3233, po3234, po3235, po3236, po3237, po3238, po3239,
    po3240, po3241, po3242, po3243, po3244, po3245, po3246, po3247, po3248,
    po3249, po3250, po3251, po3252, po3253, po3254, po3255, po3256, po3257,
    po3258, po3259, po3260, po3261, po3262, po3263, po3264, po3265, po3266,
    po3267, po3268, po3269, po3270, po3271, po3272, po3273, po3274, po3275,
    po3276, po3277, po3278, po3279, po3280, po3281, po3282, po3283, po3284,
    po3285, po3286, po3287, po3288, po3289, po3290, po3291, po3292, po3293,
    po3294, po3295, po3296, po3297, po3298, po3299, po3300, po3301, po3302,
    po3303, po3304, po3305, po3306, po3307, po3308, po3309, po3310, po3311,
    po3312, po3313, po3314, po3315, po3316, po3317, po3318, po3319, po3320,
    po3321, po3322, po3323, po3324, po3325, po3326, po3327, po3328, po3329,
    po3330, po3331, po3332, po3333, po3334, po3335, po3336, po3337, po3338,
    po3339, po3340, po3341, po3342, po3343, po3344, po3345, po3346, po3347,
    po3348, po3349, po3350, po3351, po3352, po3353, po3354, po3355, po3356,
    po3357, po3358, po3359, po3360, po3361, po3362, po3363, po3364, po3365,
    po3366, po3367, po3368, po3369, po3370, po3371, po3372, po3373, po3374,
    po3375, po3376, po3377, po3378, po3379, po3380, po3381, po3382, po3383,
    po3384, po3385, po3386, po3387, po3388, po3389, po3390, po3391, po3392,
    po3393, po3394, po3395, po3396, po3397, po3398, po3399, po3400, po3401,
    po3402, po3403, po3404, po3405, po3406, po3407, po3408, po3409, po3410,
    po3411, po3412, po3413, po3414, po3415, po3416, po3417, po3418, po3419,
    po3420, po3421, po3422, po3423, po3424, po3425, po3426, po3427, po3428,
    po3429, po3430, po3431, po3432, po3433, po3434, po3435, po3436, po3437,
    po3438, po3439, po3440, po3441, po3442, po3443, po3444, po3445, po3446,
    po3447, po3448, po3449, po3450, po3451, po3452, po3453, po3454, po3455,
    po3456, po3457, po3458, po3459, po3460, po3461, po3462, po3463, po3464,
    po3465, po3466, po3467, po3468, po3469, po3470, po3471, po3472, po3473,
    po3474, po3475, po3476, po3477, po3478, po3479, po3480, po3481, po3482,
    po3483, po3484, po3485, po3486, po3487, po3488, po3489, po3490, po3491,
    po3492, po3493, po3494, po3495, po3496, po3497, po3498, po3499, po3500,
    po3501, po3502, po3503, po3504, po3505, po3506, po3507, po3508, po3509,
    po3510, po3511, po3512, po3513, po3514, po3515, po3516, po3517, po3518,
    po3519, po3520, po3521, po3522, po3523, po3524, po3525, po3526, po3527,
    po3528, po3529, po3530, po3531, po3532, po3533, po3534, po3535, po3536,
    po3537, po3538, po3539, po3540, po3541, po3542, po3543, po3544, po3545,
    po3546, po3547, po3548, po3549, po3550, po3551, po3552, po3553, po3554,
    po3555, po3556, po3557, po3558, po3559, po3560, po3561, po3562, po3563,
    po3564, po3565, po3566, po3567, po3568, po3569, po3570, po3571, po3572,
    po3573, po3574, po3575, po3576, po3577, po3578, po3579, po3580, po3581,
    po3582, po3583, po3584, po3585, po3586, po3587, po3588, po3589, po3590,
    po3591, po3592, po3593, po3594, po3595, po3596, po3597, po3598, po3599,
    po3600, po3601, po3602, po3603, po3604, po3605, po3606, po3607, po3608,
    po3609, po3610, po3611, po3612, po3613, po3614, po3615, po3616, po3617,
    po3618, po3619, po3620, po3621, po3622, po3623, po3624, po3625, po3626,
    po3627, po3628, po3629, po3630, po3631, po3632, po3633, po3634, po3635,
    po3636, po3637, po3638, po3639, po3640, po3641, po3642, po3643, po3644,
    po3645, po3646, po3647, po3648, po3649, po3650, po3651, po3652, po3653,
    po3654, po3655, po3656, po3657, po3658, po3659, po3660, po3661, po3662,
    po3663, po3664, po3665, po3666, po3667, po3668, po3669, po3670, po3671,
    po3672, po3673, po3674, po3675, po3676, po3677, po3678, po3679, po3680,
    po3681, po3682, po3683, po3684, po3685, po3686, po3687, po3688, po3689,
    po3690, po3691, po3692, po3693, po3694, po3695, po3696, po3697, po3698,
    po3699, po3700, po3701, po3702, po3703, po3704, po3705, po3706, po3707,
    po3708, po3709, po3710, po3711, po3712, po3713, po3714, po3715, po3716,
    po3717, po3718, po3719, po3720, po3721, po3722, po3723, po3724, po3725,
    po3726, po3727, po3728, po3729, po3730, po3731, po3732, po3733, po3734,
    po3735, po3736, po3737, po3738, po3739, po3740, po3741, po3742, po3743,
    po3744, po3745, po3746, po3747, po3748, po3749, po3750, po3751, po3752,
    po3753, po3754, po3755, po3756, po3757, po3758, po3759, po3760, po3761,
    po3762, po3763, po3764, po3765, po3766, po3767, po3768, po3769, po3770,
    po3771, po3772, po3773, po3774, po3775, po3776, po3777, po3778, po3779,
    po3780, po3781, po3782, po3783, po3784, po3785, po3786, po3787, po3788,
    po3789, po3790, po3791, po3792, po3793, po3794, po3795, po3796, po3797,
    po3798, po3799, po3800, po3801, po3802, po3803, po3804, po3805, po3806,
    po3807, po3808, po3809, po3810, po3811, po3812, po3813, po3814, po3815,
    po3816, po3817, po3818, po3819, po3820, po3821, po3822, po3823, po3824,
    po3825, po3826, po3827, po3828, po3829, po3830, po3831, po3832, po3833,
    po3834, po3835, po3836, po3837, po3838, po3839, po3840, po3841, po3842,
    po3843, po3844, po3845, po3846, po3847, po3848, po3849, po3850, po3851,
    po3852, po3853, po3854, po3855, po3856, po3857, po3858, po3859, po3860,
    po3861, po3862, po3863, po3864, po3865, po3866, po3867, po3868, po3869,
    po3870, po3871, po3872, po3873, po3874, po3875, po3876, po3877, po3878,
    po3879, po3880, po3881, po3882, po3883, po3884, po3885, po3886, po3887,
    po3888, po3889, po3890, po3891, po3892, po3893, po3894, po3895, po3896,
    po3897, po3898, po3899, po3900, po3901, po3902, po3903, po3904, po3905,
    po3906, po3907, po3908, po3909, po3910, po3911, po3912, po3913, po3914,
    po3915, po3916, po3917, po3918, po3919, po3920, po3921, po3922, po3923,
    po3924, po3925, po3926, po3927, po3928, po3929, po3930, po3931, po3932,
    po3933, po3934, po3935, po3936, po3937, po3938, po3939, po3940, po3941,
    po3942, po3943, po3944, po3945, po3946, po3947, po3948, po3949, po3950,
    po3951, po3952, po3953, po3954, po3955, po3956, po3957, po3958, po3959,
    po3960, po3961, po3962, po3963, po3964, po3965, po3966, po3967, po3968,
    po3969, po3970, po3971, po3972, po3973, po3974, po3975, po3976, po3977,
    po3978, po3979, po3980, po3981, po3982, po3983, po3984, po3985, po3986,
    po3987, po3988, po3989, po3990, po3991, po3992, po3993, po3994, po3995,
    po3996, po3997, po3998, po3999, po4000, po4001, po4002, po4003, po4004,
    po4005, po4006, po4007, po4008, po4009, po4010, po4011, po4012, po4013,
    po4014, po4015, po4016, po4017, po4018, po4019, po4020, po4021, po4022,
    po4023, po4024, po4025, po4026, po4027, po4028, po4029, po4030, po4031,
    po4032, po4033, po4034, po4035, po4036, po4037, po4038, po4039, po4040,
    po4041, po4042, po4043, po4044, po4045, po4046, po4047, po4048, po4049,
    po4050, po4051, po4052, po4053, po4054, po4055, po4056, po4057, po4058,
    po4059, po4060, po4061, po4062, po4063, po4064, po4065, po4066, po4067,
    po4068, po4069, po4070, po4071, po4072, po4073, po4074, po4075, po4076,
    po4077, po4078, po4079, po4080, po4081, po4082, po4083, po4084, po4085,
    po4086, po4087, po4088, po4089, po4090, po4091, po4092, po4093, po4094,
    po4095, po4096, po4097, po4098, po4099, po4100, po4101, po4102, po4103,
    po4104, po4105, po4106, po4107, po4108, po4109, po4110, po4111, po4112,
    po4113, po4114, po4115, po4116, po4117, po4118, po4119, po4120, po4121,
    po4122, po4123, po4124, po4125, po4126, po4127, po4128, po4129, po4130,
    po4131, po4132, po4133, po4134, po4135, po4136, po4137, po4138, po4139,
    po4140, po4141, po4142, po4143, po4144, po4145, po4146, po4147, po4148,
    po4149, po4150, po4151, po4152, po4153, po4154, po4155, po4156, po4157,
    po4158, po4159, po4160, po4161, po4162, po4163, po4164, po4165, po4166,
    po4167, po4168, po4169, po4170, po4171, po4172, po4173, po4174, po4175,
    po4176, po4177, po4178, po4179, po4180, po4181, po4182, po4183, po4184,
    po4185, po4186, po4187, po4188, po4189, po4190, po4191, po4192, po4193,
    po4194, po4195, po4196, po4197, po4198, po4199, po4200, po4201, po4202,
    po4203, po4204, po4205, po4206, po4207, po4208, po4209, po4210, po4211,
    po4212, po4213, po4214, po4215, po4216, po4217, po4218, po4219, po4220,
    po4221, po4222, po4223, po4224, po4225, po4226, po4227, po4228, po4229,
    po4230, po4231, po4232, po4233, po4234, po4235, po4236, po4237, po4238,
    po4239, po4240, po4241, po4242, po4243, po4244, po4245, po4246, po4247,
    po4248, po4249, po4250, po4251, po4252, po4253, po4254, po4255, po4256,
    po4257, po4258, po4259, po4260, po4261, po4262, po4263, po4264, po4265,
    po4266, po4267, po4268, po4269, po4270, po4271, po4272, po4273, po4274,
    po4275, po4276, po4277, po4278, po4279, po4280, po4281, po4282, po4283,
    po4284, po4285, po4286, po4287, po4288, po4289, po4290, po4291, po4292,
    po4293, po4294, po4295, po4296, po4297, po4298, po4299, po4300, po4301,
    po4302, po4303, po4304, po4305, po4306, po4307, po4308, po4309, po4310,
    po4311, po4312, po4313, po4314, po4315, po4316, po4317, po4318, po4319,
    po4320, po4321, po4322, po4323, po4324, po4325, po4326, po4327, po4328,
    po4329, po4330, po4331, po4332, po4333, po4334, po4335, po4336, po4337,
    po4338, po4339, po4340, po4341, po4342, po4343, po4344, po4345, po4346,
    po4347, po4348, po4349, po4350, po4351, po4352, po4353, po4354, po4355,
    po4356, po4357, po4358, po4359, po4360, po4361, po4362, po4363, po4364,
    po4365, po4366, po4367, po4368, po4369, po4370, po4371, po4372, po4373,
    po4374, po4375, po4376, po4377, po4378, po4379, po4380, po4381, po4382,
    po4383, po4384, po4385, po4386, po4387, po4388, po4389, po4390, po4391,
    po4392, po4393, po4394, po4395, po4396, po4397, po4398, po4399, po4400,
    po4401, po4402, po4403, po4404, po4405, po4406, po4407, po4408, po4409,
    po4410, po4411, po4412, po4413, po4414, po4415, po4416, po4417, po4418,
    po4419, po4420, po4421, po4422, po4423, po4424, po4425, po4426, po4427,
    po4428, po4429, po4430, po4431, po4432, po4433, po4434, po4435, po4436,
    po4437, po4438, po4439, po4440, po4441, po4442, po4443, po4444, po4445,
    po4446, po4447, po4448, po4449, po4450, po4451, po4452, po4453, po4454,
    po4455, po4456, po4457, po4458, po4459, po4460, po4461, po4462, po4463,
    po4464, po4465, po4466, po4467, po4468, po4469, po4470, po4471, po4472,
    po4473, po4474, po4475, po4476, po4477, po4478, po4479, po4480, po4481,
    po4482, po4483, po4484, po4485, po4486, po4487, po4488, po4489, po4490,
    po4491, po4492, po4493, po4494, po4495, po4496, po4497, po4498, po4499,
    po4500, po4501, po4502, po4503, po4504, po4505, po4506, po4507, po4508,
    po4509, po4510, po4511, po4512, po4513, po4514, po4515, po4516, po4517,
    po4518, po4519, po4520, po4521, po4522, po4523, po4524, po4525, po4526,
    po4527, po4528, po4529, po4530, po4531, po4532, po4533, po4534, po4535,
    po4536, po4537, po4538, po4539, po4540, po4541, po4542, po4543, po4544,
    po4545, po4546, po4547, po4548, po4549, po4550, po4551, po4552, po4553,
    po4554, po4555, po4556, po4557, po4558, po4559, po4560, po4561, po4562,
    po4563, po4564, po4565, po4566, po4567, po4568, po4569, po4570, po4571,
    po4572, po4573, po4574, po4575, po4576, po4577, po4578, po4579, po4580,
    po4581, po4582, po4583, po4584, po4585, po4586, po4587, po4588, po4589,
    po4590, po4591, po4592, po4593, po4594, po4595, po4596, po4597, po4598,
    po4599, po4600, po4601, po4602, po4603, po4604, po4605, po4606, po4607,
    po4608, po4609, po4610, po4611, po4612, po4613, po4614, po4615, po4616,
    po4617, po4618, po4619, po4620, po4621, po4622, po4623, po4624, po4625,
    po4626, po4627, po4628, po4629, po4630, po4631, po4632, po4633, po4634,
    po4635, po4636, po4637, po4638, po4639, po4640, po4641, po4642, po4643,
    po4644, po4645, po4646, po4647, po4648, po4649, po4650, po4651, po4652,
    po4653, po4654, po4655, po4656, po4657, po4658, po4659, po4660, po4661,
    po4662, po4663, po4664, po4665, po4666, po4667, po4668, po4669, po4670,
    po4671, po4672, po4673, po4674, po4675, po4676, po4677, po4678, po4679,
    po4680, po4681, po4682, po4683, po4684, po4685, po4686, po4687, po4688,
    po4689, po4690, po4691, po4692, po4693, po4694, po4695, po4696, po4697,
    po4698, po4699, po4700, po4701, po4702, po4703, po4704, po4705, po4706,
    po4707, po4708, po4709, po4710, po4711, po4712, po4713, po4714, po4715,
    po4716, po4717, po4718, po4719, po4720, po4721, po4722, po4723, po4724,
    po4725, po4726, po4727, po4728, po4729, po4730, po4731, po4732, po4733,
    po4734, po4735, po4736, po4737, po4738, po4739, po4740, po4741, po4742,
    po4743, po4744, po4745, po4746, po4747, po4748, po4749, po4750, po4751,
    po4752, po4753, po4754, po4755, po4756, po4757, po4758, po4759, po4760,
    po4761, po4762, po4763, po4764, po4765, po4766, po4767, po4768, po4769,
    po4770, po4771, po4772, po4773, po4774, po4775, po4776, po4777, po4778,
    po4779, po4780, po4781, po4782, po4783, po4784, po4785, po4786, po4787,
    po4788, po4789, po4790, po4791, po4792, po4793, po4794, po4795, po4796,
    po4797, po4798, po4799, po4800, po4801, po4802, po4803, po4804, po4805,
    po4806, po4807, po4808, po4809, po4810, po4811, po4812, po4813, po4814,
    po4815, po4816, po4817, po4818, po4819, po4820, po4821, po4822, po4823,
    po4824, po4825, po4826, po4827, po4828, po4829, po4830, po4831, po4832,
    po4833, po4834, po4835, po4836, po4837, po4838, po4839, po4840, po4841,
    po4842, po4843, po4844, po4845, po4846, po4847, po4848, po4849, po4850,
    po4851, po4852, po4853, po4854, po4855, po4856, po4857, po4858, po4859,
    po4860, po4861, po4862, po4863, po4864, po4865, po4866, po4867, po4868,
    po4869, po4870, po4871, po4872, po4873, po4874, po4875, po4876, po4877,
    po4878, po4879, po4880, po4881, po4882, po4883, po4884, po4885, po4886,
    po4887, po4888, po4889, po4890, po4891, po4892, po4893, po4894, po4895,
    po4896, po4897, po4898, po4899, po4900, po4901, po4902, po4903, po4904,
    po4905, po4906, po4907, po4908, po4909, po4910, po4911, po4912, po4913,
    po4914, po4915, po4916, po4917, po4918, po4919, po4920, po4921, po4922,
    po4923, po4924, po4925, po4926, po4927, po4928, po4929, po4930, po4931,
    po4932, po4933, po4934, po4935, po4936, po4937, po4938, po4939, po4940,
    po4941, po4942, po4943, po4944, po4945, po4946, po4947, po4948, po4949,
    po4950, po4951, po4952, po4953, po4954, po4955, po4956, po4957, po4958,
    po4959, po4960, po4961, po4962, po4963, po4964, po4965, po4966, po4967,
    po4968, po4969, po4970, po4971, po4972, po4973, po4974, po4975, po4976,
    po4977, po4978, po4979, po4980, po4981, po4982, po4983, po4984, po4985,
    po4986, po4987, po4988, po4989, po4990, po4991, po4992, po4993, po4994,
    po4995, po4996, po4997, po4998, po4999, po5000, po5001, po5002, po5003,
    po5004, po5005, po5006, po5007, po5008, po5009, po5010, po5011, po5012,
    po5013, po5014, po5015, po5016, po5017, po5018, po5019, po5020, po5021,
    po5022, po5023, po5024, po5025, po5026, po5027, po5028, po5029, po5030,
    po5031, po5032, po5033, po5034, po5035, po5036, po5037, po5038, po5039,
    po5040, po5041, po5042, po5043, po5044, po5045, po5046, po5047, po5048,
    po5049, po5050, po5051, po5052, po5053, po5054, po5055, po5056, po5057,
    po5058, po5059, po5060, po5061, po5062, po5063, po5064, po5065, po5066,
    po5067, po5068, po5069, po5070, po5071, po5072, po5073, po5074, po5075,
    po5076, po5077, po5078, po5079, po5080, po5081, po5082, po5083, po5084,
    po5085, po5086, po5087, po5088, po5089, po5090, po5091, po5092, po5093,
    po5094, po5095, po5096, po5097, po5098, po5099, po5100, po5101, po5102,
    po5103, po5104, po5105, po5106, po5107, po5108, po5109, po5110, po5111,
    po5112, po5113, po5114, po5115, po5116, po5117, po5118, po5119, po5120,
    po5121, po5122, po5123, po5124, po5125, po5126, po5127, po5128, po5129,
    po5130, po5131, po5132, po5133, po5134, po5135, po5136, po5137, po5138,
    po5139, po5140, po5141, po5142, po5143, po5144, po5145, po5146, po5147,
    po5148, po5149, po5150, po5151, po5152, po5153, po5154, po5155, po5156,
    po5157, po5158, po5159, po5160, po5161, po5162, po5163, po5164, po5165,
    po5166, po5167, po5168, po5169, po5170, po5171, po5172, po5173, po5174,
    po5175, po5176, po5177, po5178, po5179, po5180, po5181, po5182, po5183,
    po5184, po5185, po5186, po5187, po5188, po5189, po5190, po5191, po5192,
    po5193, po5194, po5195, po5196, po5197, po5198, po5199, po5200, po5201,
    po5202, po5203, po5204, po5205, po5206, po5207, po5208, po5209, po5210,
    po5211, po5212, po5213, po5214, po5215, po5216, po5217, po5218, po5219,
    po5220, po5221, po5222, po5223, po5224, po5225, po5226, po5227, po5228,
    po5229, po5230, po5231, po5232, po5233, po5234, po5235, po5236, po5237,
    po5238, po5239, po5240, po5241, po5242, po5243, po5244, po5245, po5246,
    po5247, po5248, po5249, po5250, po5251, po5252, po5253, po5254, po5255,
    po5256, po5257, po5258, po5259, po5260, po5261, po5262, po5263, po5264,
    po5265, po5266, po5267, po5268, po5269, po5270, po5271, po5272, po5273,
    po5274, po5275, po5276, po5277, po5278, po5279, po5280, po5281, po5282,
    po5283, po5284, po5285, po5286, po5287, po5288, po5289, po5290, po5291,
    po5292, po5293, po5294, po5295, po5296, po5297, po5298, po5299, po5300,
    po5301, po5302, po5303, po5304, po5305, po5306, po5307, po5308, po5309,
    po5310, po5311, po5312, po5313, po5314, po5315, po5316, po5317, po5318,
    po5319, po5320, po5321, po5322, po5323, po5324, po5325, po5326, po5327,
    po5328, po5329, po5330, po5331, po5332, po5333, po5334, po5335, po5336,
    po5337, po5338, po5339, po5340, po5341, po5342, po5343, po5344, po5345,
    po5346, po5347, po5348, po5349, po5350, po5351, po5352, po5353, po5354,
    po5355, po5356, po5357, po5358, po5359, po5360, po5361, po5362, po5363,
    po5364, po5365, po5366, po5367, po5368, po5369, po5370, po5371, po5372,
    po5373, po5374, po5375, po5376, po5377, po5378, po5379, po5380, po5381,
    po5382, po5383, po5384, po5385, po5386, po5387, po5388, po5389, po5390,
    po5391, po5392, po5393, po5394, po5395, po5396, po5397, po5398, po5399,
    po5400, po5401, po5402, po5403, po5404, po5405, po5406, po5407, po5408,
    po5409, po5410, po5411, po5412, po5413, po5414, po5415, po5416, po5417,
    po5418, po5419, po5420, po5421, po5422, po5423, po5424, po5425, po5426,
    po5427, po5428, po5429, po5430, po5431, po5432, po5433, po5434, po5435,
    po5436, po5437, po5438, po5439, po5440, po5441, po5442, po5443, po5444,
    po5445, po5446, po5447, po5448, po5449, po5450, po5451, po5452, po5453,
    po5454, po5455, po5456, po5457, po5458, po5459, po5460, po5461, po5462,
    po5463, po5464, po5465, po5466, po5467, po5468, po5469, po5470, po5471,
    po5472, po5473, po5474, po5475, po5476, po5477, po5478, po5479, po5480,
    po5481, po5482, po5483, po5484, po5485, po5486, po5487, po5488, po5489,
    po5490, po5491, po5492, po5493, po5494, po5495, po5496, po5497, po5498,
    po5499, po5500, po5501, po5502, po5503, po5504, po5505, po5506, po5507,
    po5508, po5509, po5510, po5511, po5512, po5513, po5514, po5515, po5516,
    po5517, po5518, po5519, po5520, po5521, po5522, po5523, po5524, po5525,
    po5526, po5527, po5528, po5529, po5530, po5531, po5532, po5533, po5534,
    po5535, po5536, po5537, po5538, po5539, po5540, po5541, po5542, po5543,
    po5544, po5545, po5546, po5547, po5548, po5549, po5550, po5551, po5552,
    po5553, po5554, po5555, po5556, po5557, po5558, po5559, po5560, po5561,
    po5562, po5563, po5564, po5565, po5566, po5567, po5568, po5569, po5570,
    po5571, po5572, po5573, po5574, po5575, po5576, po5577, po5578, po5579,
    po5580, po5581, po5582, po5583, po5584, po5585, po5586, po5587, po5588,
    po5589, po5590, po5591, po5592, po5593, po5594, po5595, po5596, po5597,
    po5598, po5599, po5600, po5601, po5602, po5603, po5604, po5605, po5606,
    po5607, po5608, po5609, po5610, po5611, po5612, po5613, po5614, po5615,
    po5616, po5617, po5618, po5619, po5620, po5621, po5622, po5623, po5624,
    po5625, po5626, po5627, po5628, po5629, po5630, po5631, po5632, po5633,
    po5634, po5635, po5636, po5637, po5638, po5639, po5640, po5641, po5642,
    po5643, po5644, po5645, po5646, po5647, po5648, po5649, po5650, po5651,
    po5652, po5653, po5654, po5655, po5656, po5657, po5658, po5659, po5660,
    po5661, po5662, po5663, po5664, po5665, po5666, po5667, po5668, po5669,
    po5670, po5671, po5672, po5673, po5674, po5675, po5676, po5677, po5678,
    po5679, po5680, po5681, po5682, po5683, po5684, po5685, po5686, po5687,
    po5688, po5689, po5690, po5691, po5692, po5693, po5694, po5695, po5696,
    po5697, po5698, po5699, po5700, po5701, po5702, po5703, po5704, po5705,
    po5706, po5707, po5708, po5709, po5710, po5711, po5712, po5713, po5714,
    po5715, po5716, po5717, po5718, po5719, po5720, po5721, po5722, po5723,
    po5724, po5725, po5726, po5727, po5728, po5729, po5730, po5731, po5732,
    po5733, po5734, po5735, po5736, po5737, po5738, po5739, po5740, po5741,
    po5742, po5743, po5744, po5745, po5746, po5747, po5748, po5749, po5750,
    po5751, po5752, po5753, po5754, po5755, po5756, po5757, po5758, po5759,
    po5760, po5761, po5762, po5763, po5764, po5765, po5766, po5767, po5768,
    po5769, po5770, po5771, po5772, po5773, po5774, po5775, po5776, po5777,
    po5778, po5779, po5780, po5781, po5782, po5783, po5784, po5785, po5786,
    po5787, po5788, po5789, po5790, po5791, po5792, po5793, po5794, po5795,
    po5796, po5797, po5798, po5799, po5800, po5801, po5802, po5803, po5804,
    po5805, po5806, po5807, po5808, po5809, po5810, po5811, po5812, po5813,
    po5814, po5815, po5816, po5817, po5818, po5819, po5820, po5821, po5822,
    po5823, po5824, po5825, po5826, po5827, po5828, po5829, po5830, po5831,
    po5832, po5833, po5834, po5835, po5836, po5837, po5838, po5839, po5840,
    po5841, po5842, po5843, po5844, po5845, po5846, po5847, po5848, po5849,
    po5850, po5851, po5852, po5853, po5854, po5855, po5856, po5857, po5858,
    po5859, po5860, po5861, po5862, po5863, po5864, po5865, po5866, po5867,
    po5868, po5869, po5870, po5871, po5872, po5873, po5874, po5875, po5876,
    po5877, po5878, po5879, po5880, po5881, po5882, po5883, po5884, po5885,
    po5886, po5887, po5888, po5889, po5890, po5891, po5892, po5893, po5894,
    po5895, po5896, po5897, po5898, po5899, po5900, po5901, po5902, po5903,
    po5904, po5905, po5906, po5907, po5908, po5909, po5910, po5911, po5912,
    po5913, po5914, po5915, po5916, po5917, po5918, po5919, po5920, po5921,
    po5922, po5923, po5924, po5925, po5926, po5927, po5928, po5929, po5930,
    po5931, po5932, po5933, po5934, po5935, po5936, po5937, po5938, po5939,
    po5940, po5941, po5942, po5943, po5944, po5945, po5946, po5947, po5948,
    po5949, po5950, po5951, po5952, po5953, po5954, po5955, po5956, po5957,
    po5958, po5959, po5960, po5961, po5962, po5963, po5964, po5965, po5966,
    po5967, po5968, po5969, po5970, po5971, po5972, po5973, po5974, po5975,
    po5976, po5977, po5978, po5979, po5980, po5981, po5982, po5983, po5984,
    po5985, po5986, po5987, po5988, po5989, po5990, po5991, po5992, po5993,
    po5994, po5995, po5996, po5997, po5998, po5999, po6000, po6001, po6002,
    po6003, po6004, po6005, po6006, po6007, po6008, po6009, po6010, po6011,
    po6012, po6013, po6014, po6015, po6016, po6017, po6018, po6019, po6020,
    po6021, po6022, po6023, po6024, po6025, po6026, po6027, po6028, po6029,
    po6030, po6031, po6032, po6033, po6034, po6035, po6036, po6037, po6038,
    po6039, po6040, po6041, po6042, po6043, po6044, po6045, po6046, po6047,
    po6048, po6049, po6050, po6051, po6052, po6053, po6054, po6055, po6056,
    po6057, po6058, po6059, po6060, po6061, po6062, po6063, po6064, po6065,
    po6066, po6067, po6068, po6069, po6070, po6071, po6072, po6073, po6074,
    po6075, po6076, po6077, po6078, po6079, po6080, po6081, po6082, po6083,
    po6084, po6085, po6086, po6087, po6088, po6089, po6090, po6091, po6092,
    po6093, po6094, po6095, po6096, po6097, po6098, po6099, po6100, po6101,
    po6102, po6103, po6104, po6105, po6106, po6107, po6108, po6109, po6110,
    po6111, po6112, po6113, po6114, po6115, po6116, po6117, po6118, po6119,
    po6120, po6121, po6122, po6123, po6124, po6125, po6126, po6127, po6128,
    po6129, po6130, po6131, po6132, po6133, po6134, po6135, po6136, po6137,
    po6138, po6139, po6140, po6141, po6142, po6143, po6144, po6145, po6146,
    po6147, po6148, po6149, po6150, po6151, po6152, po6153, po6154, po6155,
    po6156, po6157, po6158, po6159, po6160, po6161, po6162, po6163, po6164,
    po6165, po6166, po6167, po6168, po6169, po6170, po6171, po6172, po6173,
    po6174, po6175, po6176, po6177, po6178, po6179, po6180, po6181, po6182,
    po6183, po6184, po6185, po6186, po6187, po6188, po6189, po6190, po6191,
    po6192, po6193, po6194, po6195, po6196, po6197, po6198, po6199, po6200,
    po6201, po6202, po6203, po6204, po6205, po6206, po6207, po6208, po6209,
    po6210, po6211, po6212, po6213, po6214, po6215, po6216, po6217, po6218,
    po6219, po6220, po6221, po6222, po6223, po6224, po6225, po6226, po6227,
    po6228, po6229, po6230, po6231, po6232, po6233, po6234, po6235, po6236,
    po6237, po6238, po6239, po6240, po6241, po6242, po6243, po6244, po6245,
    po6246, po6247, po6248, po6249, po6250, po6251, po6252, po6253, po6254,
    po6255, po6256, po6257, po6258, po6259, po6260, po6261, po6262, po6263,
    po6264, po6265, po6266, po6267, po6268, po6269, po6270, po6271, po6272,
    po6273, po6274, po6275, po6276, po6277, po6278, po6279, po6280, po6281,
    po6282, po6283, po6284, po6285, po6286, po6287, po6288, po6289, po6290,
    po6291, po6292, po6293, po6294, po6295, po6296, po6297, po6298, po6299,
    po6300, po6301, po6302, po6303, po6304, po6305, po6306, po6307, po6308,
    po6309, po6310, po6311, po6312, po6313, po6314, po6315, po6316, po6317,
    po6318, po6319, po6320, po6321, po6322, po6323, po6324, po6325, po6326,
    po6327, po6328, po6329, po6330, po6331, po6332, po6333, po6334, po6335,
    po6336, po6337, po6338, po6339, po6340, po6341, po6342, po6343, po6344,
    po6345, po6346, po6347, po6348, po6349, po6350, po6351, po6352, po6353,
    po6354, po6355, po6356, po6357, po6358, po6359, po6360, po6361, po6362,
    po6363, po6364, po6365, po6366, po6367, po6368, po6369, po6370, po6371,
    po6372, po6373, po6374, po6375, po6376, po6377, po6378, po6379, po6380,
    po6381, po6382, po6383, po6384, po6385, po6386, po6387, po6388, po6389,
    po6390, po6391, po6392, po6393, po6394, po6395, po6396, po6397, po6398,
    po6399, po6400, po6401, po6402, po6403, po6404, po6405, po6406, po6407,
    po6408, po6409, po6410, po6411, po6412, po6413, po6414, po6415, po6416,
    po6417, po6418, po6419, po6420, po6421, po6422, po6423, po6424, po6425,
    po6426, po6427, po6428, po6429, po6430, po6431, po6432, po6433, po6434,
    po6435, po6436, po6437, po6438, po6439, po6440, po6441, po6442, po6443,
    po6444, po6445, po6446, po6447, po6448, po6449, po6450, po6451, po6452,
    po6453, po6454, po6455, po6456, po6457, po6458, po6459, po6460, po6461,
    po6462, po6463, po6464, po6465, po6466, po6467, po6468, po6469, po6470,
    po6471, po6472, po6473, po6474, po6475, po6476, po6477, po6478, po6479,
    po6480, po6481, po6482, po6483, po6484, po6485, po6486, po6487, po6488,
    po6489, po6490, po6491, po6492, po6493, po6494, po6495, po6496, po6497,
    po6498, po6499, po6500, po6501, po6502, po6503, po6504, po6505, po6506,
    po6507, po6508, po6509, po6510, po6511, po6512, po6513, po6514, po6515,
    po6516, po6517, po6518, po6519, po6520, po6521, po6522, po6523, po6524,
    po6525, po6526, po6527, po6528, po6529, po6530, po6531, po6532, po6533,
    po6534, po6535, po6536, po6537, po6538, po6539, po6540, po6541, po6542,
    po6543, po6544, po6545, po6546, po6547, po6548, po6549, po6550, po6551,
    po6552, po6553, po6554, po6555, po6556, po6557, po6558, po6559, po6560,
    po6561, po6562, po6563, po6564, po6565, po6566, po6567, po6568, po6569,
    po6570, po6571, po6572, po6573, po6574, po6575, po6576, po6577, po6578,
    po6579, po6580, po6581, po6582, po6583, po6584, po6585, po6586, po6587,
    po6588, po6589, po6590, po6591, po6592, po6593, po6594, po6595, po6596,
    po6597, po6598, po6599, po6600, po6601, po6602, po6603, po6604, po6605,
    po6606, po6607, po6608, po6609, po6610, po6611, po6612, po6613, po6614,
    po6615, po6616, po6617, po6618, po6619, po6620, po6621, po6622, po6623,
    po6624, po6625, po6626, po6627, po6628, po6629, po6630, po6631, po6632,
    po6633, po6634, po6635, po6636, po6637, po6638, po6639, po6640, po6641,
    po6642, po6643, po6644, po6645, po6646, po6647, po6648, po6649, po6650,
    po6651, po6652, po6653, po6654, po6655, po6656, po6657, po6658, po6659,
    po6660, po6661, po6662, po6663, po6664, po6665, po6666, po6667, po6668,
    po6669, po6670, po6671, po6672, po6673, po6674, po6675, po6676, po6677,
    po6678, po6679, po6680, po6681, po6682, po6683, po6684, po6685, po6686,
    po6687, po6688, po6689, po6690, po6691, po6692, po6693, po6694, po6695,
    po6696, po6697, po6698, po6699, po6700, po6701, po6702, po6703, po6704,
    po6705, po6706, po6707, po6708, po6709, po6710, po6711, po6712, po6713,
    po6714, po6715, po6716, po6717, po6718, po6719, po6720, po6721, po6722,
    po6723, po6724, po6725, po6726, po6727, po6728, po6729, po6730, po6731,
    po6732, po6733, po6734, po6735, po6736, po6737, po6738, po6739, po6740,
    po6741, po6742, po6743, po6744, po6745, po6746, po6747, po6748, po6749,
    po6750, po6751, po6752, po6753, po6754, po6755, po6756, po6757, po6758,
    po6759, po6760, po6761, po6762, po6763, po6764, po6765, po6766, po6767,
    po6768, po6769, po6770, po6771, po6772, po6773, po6774, po6775, po6776,
    po6777, po6778, po6779, po6780, po6781, po6782, po6783, po6784, po6785,
    po6786, po6787, po6788, po6789, po6790, po6791, po6792, po6793, po6794,
    po6795, po6796, po6797, po6798, po6799, po6800, po6801, po6802, po6803,
    po6804, po6805, po6806, po6807, po6808, po6809, po6810, po6811, po6812,
    po6813, po6814, po6815, po6816, po6817, po6818, po6819, po6820, po6821,
    po6822, po6823, po6824, po6825, po6826, po6827, po6828, po6829, po6830,
    po6831, po6832, po6833, po6834, po6835, po6836, po6837, po6838, po6839,
    po6840, po6841, po6842, po6843, po6844, po6845, po6846, po6847, po6848,
    po6849, po6850, po6851, po6852, po6853, po6854, po6855, po6856, po6857,
    po6858, po6859, po6860, po6861, po6862, po6863, po6864, po6865, po6866,
    po6867, po6868, po6869, po6870, po6871, po6872, po6873, po6874, po6875,
    po6876, po6877, po6878, po6879, po6880, po6881, po6882, po6883, po6884,
    po6885, po6886, po6887, po6888, po6889, po6890, po6891, po6892, po6893,
    po6894, po6895, po6896, po6897, po6898, po6899, po6900, po6901, po6902,
    po6903, po6904, po6905, po6906, po6907, po6908, po6909, po6910, po6911,
    po6912, po6913, po6914, po6915, po6916, po6917, po6918, po6919, po6920,
    po6921, po6922, po6923, po6924, po6925, po6926, po6927, po6928, po6929,
    po6930, po6931, po6932, po6933, po6934, po6935, po6936, po6937, po6938,
    po6939, po6940, po6941, po6942, po6943, po6944, po6945, po6946, po6947,
    po6948, po6949, po6950, po6951, po6952, po6953, po6954, po6955, po6956,
    po6957, po6958, po6959, po6960, po6961, po6962, po6963, po6964, po6965,
    po6966, po6967, po6968, po6969, po6970, po6971, po6972, po6973, po6974,
    po6975, po6976, po6977, po6978, po6979, po6980, po6981, po6982, po6983,
    po6984, po6985, po6986, po6987, po6988, po6989, po6990, po6991, po6992,
    po6993, po6994, po6995, po6996, po6997, po6998, po6999, po7000, po7001,
    po7002, po7003, po7004, po7005, po7006, po7007, po7008, po7009, po7010,
    po7011, po7012, po7013, po7014, po7015, po7016, po7017, po7018, po7019,
    po7020, po7021, po7022, po7023, po7024, po7025, po7026, po7027, po7028,
    po7029, po7030, po7031, po7032, po7033, po7034, po7035, po7036, po7037,
    po7038, po7039, po7040, po7041, po7042, po7043, po7044, po7045, po7046,
    po7047, po7048, po7049, po7050, po7051, po7052, po7053, po7054, po7055,
    po7056, po7057, po7058, po7059, po7060, po7061, po7062, po7063, po7064,
    po7065, po7066, po7067, po7068, po7069, po7070, po7071, po7072, po7073,
    po7074, po7075, po7076, po7077, po7078, po7079, po7080, po7081, po7082,
    po7083, po7084, po7085, po7086, po7087, po7088, po7089, po7090, po7091,
    po7092, po7093, po7094, po7095, po7096, po7097, po7098, po7099, po7100,
    po7101, po7102, po7103, po7104, po7105, po7106, po7107, po7108, po7109,
    po7110, po7111, po7112, po7113, po7114, po7115, po7116, po7117, po7118,
    po7119, po7120, po7121, po7122, po7123, po7124, po7125, po7126, po7127,
    po7128, po7129, po7130, po7131, po7132, po7133, po7134, po7135, po7136,
    po7137, po7138, po7139, po7140, po7141, po7142, po7143, po7144, po7145,
    po7146, po7147, po7148, po7149, po7150, po7151, po7152, po7153, po7154,
    po7155, po7156, po7157, po7158, po7159, po7160, po7161, po7162, po7163,
    po7164, po7165, po7166, po7167, po7168, po7169, po7170, po7171, po7172,
    po7173, po7174, po7175, po7176, po7177, po7178, po7179, po7180, po7181,
    po7182, po7183, po7184, po7185, po7186, po7187, po7188, po7189, po7190,
    po7191, po7192, po7193, po7194, po7195, po7196, po7197, po7198, po7199,
    po7200, po7201, po7202, po7203, po7204, po7205, po7206, po7207, po7208,
    po7209, po7210, po7211, po7212, po7213, po7214, po7215, po7216, po7217,
    po7218, po7219, po7220, po7221, po7222, po7223, po7224, po7225, po7226,
    po7227, po7228, po7229, po7230, po7231, po7232, po7233, po7234, po7235,
    po7236, po7237, po7238, po7239, po7240, po7241, po7242, po7243, po7244,
    po7245, po7246, po7247, po7248, po7249, po7250, po7251, po7252, po7253,
    po7254, po7255, po7256, po7257, po7258, po7259, po7260, po7261, po7262,
    po7263, po7264, po7265, po7266, po7267, po7268, po7269, po7270, po7271,
    po7272, po7273, po7274, po7275, po7276, po7277, po7278, po7279, po7280,
    po7281, po7282, po7283, po7284, po7285, po7286, po7287, po7288, po7289,
    po7290, po7291, po7292, po7293, po7294, po7295, po7296, po7297, po7298,
    po7299, po7300, po7301, po7302, po7303, po7304, po7305, po7306, po7307,
    po7308, po7309, po7310, po7311, po7312, po7313, po7314, po7315, po7316,
    po7317, po7318, po7319, po7320, po7321, po7322, po7323, po7324, po7325,
    po7326, po7327, po7328, po7329, po7330, po7331, po7332, po7333, po7334,
    po7335, po7336, po7337, po7338, po7339, po7340, po7341, po7342, po7343,
    po7344, po7345, po7346, po7347, po7348, po7349, po7350, po7351, po7352,
    po7353, po7354, po7355, po7356, po7357, po7358, po7359, po7360, po7361,
    po7362, po7363, po7364, po7365, po7366, po7367, po7368, po7369, po7370,
    po7371, po7372, po7373, po7374, po7375, po7376, po7377, po7378, po7379,
    po7380, po7381, po7382, po7383, po7384, po7385, po7386, po7387, po7388,
    po7389, po7390, po7391, po7392, po7393, po7394, po7395, po7396, po7397,
    po7398, po7399, po7400, po7401, po7402, po7403, po7404, po7405, po7406,
    po7407, po7408, po7409, po7410, po7411, po7412, po7413, po7414, po7415,
    po7416, po7417, po7418, po7419, po7420, po7421, po7422, po7423, po7424,
    po7425, po7426, po7427, po7428, po7429, po7430, po7431, po7432, po7433,
    po7434, po7435, po7436, po7437, po7438, po7439, po7440, po7441, po7442,
    po7443, po7444, po7445, po7446, po7447, po7448, po7449, po7450, po7451,
    po7452, po7453, po7454, po7455, po7456, po7457, po7458, po7459, po7460,
    po7461, po7462, po7463, po7464, po7465, po7466, po7467, po7468, po7469,
    po7470, po7471, po7472, po7473, po7474, po7475, po7476, po7477, po7478,
    po7479, po7480, po7481, po7482, po7483, po7484, po7485, po7486, po7487,
    po7488, po7489, po7490, po7491, po7492, po7493, po7494, po7495, po7496,
    po7497, po7498, po7499, po7500, po7501, po7502, po7503, po7504, po7505,
    po7506, po7507, po7508, po7509, po7510, po7511, po7512, po7513, po7514,
    po7515, po7516, po7517, po7518, po7519, po7520, po7521, po7522, po7523,
    po7524, po7525, po7526, po7527, po7528, po7529, po7530, po7531, po7532,
    po7533, po7534, po7535, po7536, po7537, po7538, po7539, po7540, po7541,
    po7542, po7543, po7544, po7545, po7546, po7547, po7548, po7549, po7550,
    po7551, po7552, po7553, po7554, po7555, po7556, po7557, po7558, po7559,
    po7560, po7561, po7562, po7563, po7564, po7565, po7566, po7567, po7568,
    po7569, po7570, po7571, po7572, po7573, po7574, po7575, po7576, po7577,
    po7578, po7579, po7580, po7581, po7582, po7583, po7584, po7585, po7586,
    po7587, po7588, po7589, po7590, po7591, po7592, po7593, po7594, po7595,
    po7596, po7597, po7598, po7599, po7600, po7601, po7602, po7603, po7604,
    po7605, po7606, po7607, po7608, po7609, po7610, po7611, po7612, po7613,
    po7614, po7615, po7616, po7617, po7618, po7619, po7620, po7621, po7622,
    po7623, po7624, po7625, po7626, po7627, po7628, po7629, po7630, po7631,
    po7632, po7633, po7634, po7635, po7636, po7637, po7638, po7639, po7640,
    po7641, po7642, po7643, po7644, po7645, po7646, po7647, po7648, po7649,
    po7650, po7651, po7652, po7653, po7654, po7655, po7656, po7657, po7658,
    po7659, po7660, po7661, po7662, po7663, po7664, po7665, po7666, po7667,
    po7668, po7669, po7670, po7671, po7672, po7673, po7674, po7675, po7676,
    po7677, po7678, po7679, po7680, po7681, po7682, po7683, po7684, po7685,
    po7686, po7687, po7688, po7689, po7690, po7691, po7692, po7693, po7694,
    po7695, po7696, po7697, po7698, po7699, po7700, po7701, po7702, po7703,
    po7704, po7705, po7706, po7707, po7708, po7709, po7710, po7711, po7712,
    po7713, po7714, po7715, po7716, po7717, po7718, po7719, po7720, po7721,
    po7722, po7723, po7724, po7725, po7726, po7727, po7728, po7729, po7730,
    po7731, po7732, po7733, po7734, po7735, po7736, po7737, po7738, po7739,
    po7740, po7741, po7742, po7743, po7744, po7745, po7746, po7747, po7748,
    po7749, po7750, po7751, po7752, po7753, po7754, po7755, po7756, po7757,
    po7758, po7759, po7760, po7761, po7762, po7763, po7764, po7765, po7766,
    po7767, po7768, po7769, po7770, po7771, po7772, po7773, po7774, po7775,
    po7776, po7777, po7778, po7779, po7780, po7781, po7782, po7783, po7784,
    po7785, po7786, po7787, po7788, po7789, po7790, po7791, po7792, po7793,
    po7794, po7795, po7796, po7797, po7798, po7799, po7800, po7801, po7802,
    po7803, po7804, po7805, po7806, po7807, po7808, po7809, po7810, po7811,
    po7812, po7813, po7814, po7815, po7816, po7817, po7818, po7819, po7820,
    po7821, po7822, po7823, po7824, po7825, po7826, po7827, po7828, po7829,
    po7830, po7831, po7832, po7833, po7834, po7835, po7836, po7837, po7838,
    po7839, po7840, po7841, po7842, po7843, po7844, po7845, po7846, po7847,
    po7848, po7849, po7850, po7851, po7852, po7853, po7854, po7855, po7856,
    po7857, po7858, po7859, po7860, po7861, po7862, po7863, po7864, po7865,
    po7866, po7867, po7868, po7869, po7870, po7871, po7872, po7873, po7874,
    po7875, po7876, po7877, po7878, po7879, po7880, po7881, po7882, po7883,
    po7884, po7885, po7886, po7887, po7888, po7889, po7890, po7891, po7892,
    po7893, po7894, po7895, po7896, po7897, po7898, po7899, po7900, po7901,
    po7902, po7903, po7904, po7905, po7906, po7907, po7908, po7909, po7910,
    po7911, po7912, po7913, po7914, po7915, po7916, po7917, po7918, po7919,
    po7920, po7921, po7922, po7923, po7924, po7925, po7926, po7927, po7928,
    po7929, po7930, po7931, po7932, po7933, po7934, po7935, po7936, po7937,
    po7938, po7939, po7940, po7941, po7942, po7943, po7944, po7945, po7946,
    po7947, po7948, po7949, po7950, po7951, po7952, po7953, po7954, po7955,
    po7956, po7957, po7958, po7959, po7960, po7961, po7962, po7963, po7964,
    po7965, po7966, po7967, po7968, po7969, po7970, po7971, po7972, po7973,
    po7974, po7975, po7976, po7977, po7978, po7979, po7980, po7981, po7982,
    po7983, po7984, po7985, po7986, po7987, po7988, po7989, po7990, po7991,
    po7992, po7993, po7994, po7995, po7996, po7997, po7998, po7999, po8000,
    po8001, po8002, po8003, po8004, po8005, po8006, po8007, po8008, po8009,
    po8010, po8011, po8012, po8013, po8014, po8015, po8016, po8017, po8018,
    po8019, po8020, po8021, po8022, po8023, po8024, po8025, po8026, po8027,
    po8028, po8029, po8030, po8031, po8032, po8033, po8034, po8035, po8036,
    po8037, po8038, po8039, po8040, po8041, po8042, po8043, po8044, po8045,
    po8046, po8047, po8048, po8049, po8050, po8051, po8052, po8053, po8054,
    po8055, po8056, po8057, po8058, po8059, po8060, po8061, po8062, po8063,
    po8064, po8065, po8066, po8067, po8068, po8069, po8070, po8071, po8072,
    po8073, po8074, po8075, po8076, po8077, po8078, po8079, po8080, po8081,
    po8082, po8083, po8084, po8085, po8086, po8087, po8088, po8089, po8090,
    po8091, po8092, po8093, po8094, po8095, po8096, po8097, po8098, po8099,
    po8100, po8101, po8102, po8103, po8104, po8105, po8106, po8107, po8108,
    po8109, po8110, po8111, po8112, po8113, po8114, po8115, po8116, po8117,
    po8118, po8119, po8120, po8121, po8122, po8123, po8124, po8125, po8126,
    po8127, po8128, po8129, po8130, po8131, po8132, po8133, po8134, po8135,
    po8136, po8137, po8138, po8139, po8140, po8141, po8142, po8143, po8144,
    po8145, po8146, po8147, po8148, po8149, po8150, po8151, po8152, po8153,
    po8154, po8155, po8156, po8157, po8158, po8159, po8160, po8161, po8162,
    po8163, po8164, po8165, po8166, po8167, po8168, po8169, po8170, po8171,
    po8172, po8173, po8174, po8175, po8176, po8177, po8178, po8179, po8180,
    po8181, po8182, po8183, po8184, po8185, po8186, po8187, po8188, po8189,
    po8190, po8191, po8192, po8193, po8194, po8195, po8196, po8197, po8198,
    po8199, po8200, po8201, po8202, po8203, po8204, po8205, po8206, po8207,
    po8208, po8209, po8210, po8211, po8212, po8213, po8214, po8215, po8216,
    po8217, po8218, po8219, po8220, po8221, po8222, po8223, po8224, po8225,
    po8226, po8227, po8228, po8229, po8230, po8231, po8232, po8233, po8234,
    po8235, po8236, po8237, po8238, po8239, po8240, po8241, po8242, po8243,
    po8244, po8245, po8246, po8247, po8248, po8249, po8250, po8251, po8252,
    po8253, po8254, po8255, po8256, po8257, po8258, po8259, po8260, po8261,
    po8262, po8263, po8264, po8265, po8266, po8267, po8268, po8269, po8270,
    po8271, po8272, po8273, po8274, po8275, po8276, po8277, po8278, po8279,
    po8280, po8281, po8282, po8283, po8284, po8285, po8286, po8287, po8288,
    po8289, po8290, po8291, po8292, po8293, po8294, po8295, po8296, po8297,
    po8298, po8299, po8300, po8301, po8302, po8303, po8304, po8305, po8306,
    po8307, po8308, po8309, po8310, po8311, po8312, po8313, po8314, po8315,
    po8316, po8317, po8318, po8319, po8320, po8321, po8322, po8323, po8324,
    po8325, po8326, po8327, po8328, po8329, po8330, po8331, po8332, po8333,
    po8334, po8335, po8336, po8337, po8338, po8339, po8340, po8341, po8342,
    po8343, po8344, po8345, po8346, po8347, po8348, po8349, po8350, po8351,
    po8352, po8353, po8354, po8355, po8356, po8357, po8358, po8359, po8360,
    po8361, po8362, po8363, po8364, po8365, po8366, po8367, po8368, po8369,
    po8370, po8371, po8372, po8373, po8374, po8375, po8376, po8377, po8378,
    po8379, po8380, po8381, po8382, po8383, po8384, po8385, po8386, po8387,
    po8388, po8389, po8390, po8391, po8392, po8393, po8394, po8395, po8396,
    po8397, po8398, po8399, po8400, po8401, po8402, po8403, po8404, po8405,
    po8406, po8407, po8408, po8409, po8410, po8411, po8412, po8413, po8414,
    po8415, po8416, po8417, po8418, po8419, po8420, po8421, po8422, po8423,
    po8424, po8425, po8426, po8427, po8428, po8429, po8430, po8431, po8432,
    po8433, po8434, po8435, po8436, po8437, po8438, po8439, po8440, po8441,
    po8442, po8443, po8444, po8445, po8446, po8447, po8448, po8449, po8450,
    po8451, po8452, po8453, po8454, po8455, po8456, po8457, po8458, po8459,
    po8460, po8461, po8462, po8463, po8464, po8465, po8466, po8467, po8468,
    po8469, po8470, po8471, po8472, po8473, po8474, po8475, po8476, po8477,
    po8478, po8479, po8480, po8481, po8482, po8483, po8484, po8485, po8486,
    po8487, po8488, po8489, po8490, po8491, po8492, po8493, po8494, po8495,
    po8496, po8497, po8498, po8499, po8500, po8501, po8502, po8503, po8504,
    po8505, po8506, po8507, po8508, po8509, po8510, po8511, po8512, po8513,
    po8514, po8515, po8516, po8517, po8518, po8519, po8520, po8521, po8522,
    po8523, po8524, po8525, po8526, po8527, po8528, po8529, po8530, po8531,
    po8532, po8533, po8534, po8535, po8536, po8537, po8538, po8539, po8540,
    po8541, po8542, po8543, po8544, po8545, po8546, po8547, po8548, po8549,
    po8550, po8551, po8552, po8553, po8554, po8555, po8556, po8557, po8558,
    po8559, po8560, po8561, po8562, po8563, po8564, po8565, po8566, po8567,
    po8568, po8569, po8570, po8571, po8572, po8573, po8574, po8575, po8576,
    po8577, po8578, po8579, po8580, po8581, po8582, po8583, po8584, po8585,
    po8586, po8587, po8588, po8589, po8590, po8591, po8592, po8593, po8594,
    po8595, po8596, po8597, po8598, po8599, po8600, po8601, po8602, po8603,
    po8604, po8605, po8606, po8607, po8608, po8609, po8610, po8611, po8612,
    po8613, po8614, po8615, po8616, po8617, po8618, po8619, po8620, po8621,
    po8622, po8623, po8624, po8625, po8626, po8627, po8628, po8629, po8630,
    po8631, po8632, po8633, po8634, po8635, po8636, po8637, po8638, po8639,
    po8640, po8641, po8642, po8643, po8644, po8645, po8646, po8647, po8648,
    po8649, po8650, po8651, po8652, po8653, po8654, po8655, po8656, po8657,
    po8658, po8659, po8660, po8661, po8662, po8663, po8664, po8665, po8666,
    po8667, po8668, po8669, po8670, po8671, po8672, po8673, po8674, po8675,
    po8676, po8677, po8678, po8679, po8680, po8681, po8682, po8683, po8684,
    po8685, po8686, po8687, po8688, po8689, po8690, po8691, po8692, po8693,
    po8694, po8695, po8696, po8697, po8698, po8699, po8700, po8701, po8702,
    po8703, po8704, po8705, po8706, po8707, po8708, po8709, po8710, po8711,
    po8712, po8713, po8714, po8715, po8716, po8717, po8718, po8719, po8720,
    po8721, po8722, po8723, po8724, po8725, po8726, po8727, po8728, po8729,
    po8730, po8731, po8732, po8733, po8734, po8735, po8736, po8737, po8738,
    po8739, po8740, po8741, po8742, po8743, po8744, po8745, po8746, po8747,
    po8748, po8749, po8750, po8751, po8752, po8753, po8754, po8755, po8756,
    po8757, po8758, po8759, po8760, po8761, po8762, po8763, po8764, po8765,
    po8766, po8767, po8768, po8769, po8770, po8771, po8772, po8773, po8774,
    po8775, po8776, po8777, po8778, po8779, po8780, po8781, po8782, po8783,
    po8784, po8785, po8786, po8787, po8788, po8789, po8790, po8791, po8792,
    po8793, po8794, po8795, po8796, po8797, po8798, po8799, po8800, po8801,
    po8802, po8803, po8804, po8805, po8806, po8807, po8808, po8809, po8810,
    po8811, po8812, po8813, po8814, po8815, po8816, po8817, po8818, po8819,
    po8820, po8821, po8822, po8823, po8824, po8825, po8826, po8827, po8828,
    po8829, po8830, po8831, po8832, po8833, po8834, po8835, po8836, po8837,
    po8838, po8839, po8840, po8841, po8842, po8843, po8844, po8845, po8846,
    po8847, po8848, po8849, po8850, po8851, po8852, po8853, po8854, po8855,
    po8856, po8857, po8858, po8859, po8860, po8861, po8862, po8863, po8864,
    po8865, po8866, po8867, po8868, po8869, po8870, po8871, po8872, po8873,
    po8874, po8875, po8876, po8877, po8878, po8879, po8880, po8881, po8882,
    po8883, po8884, po8885, po8886, po8887, po8888, po8889, po8890, po8891,
    po8892, po8893, po8894, po8895, po8896, po8897, po8898, po8899, po8900,
    po8901, po8902, po8903, po8904, po8905, po8906, po8907, po8908, po8909,
    po8910, po8911, po8912, po8913, po8914, po8915, po8916, po8917, po8918,
    po8919, po8920, po8921, po8922, po8923, po8924, po8925, po8926, po8927,
    po8928, po8929, po8930, po8931, po8932, po8933, po8934, po8935, po8936,
    po8937, po8938, po8939, po8940, po8941, po8942, po8943, po8944, po8945,
    po8946, po8947, po8948, po8949, po8950, po8951, po8952, po8953, po8954,
    po8955, po8956, po8957, po8958, po8959, po8960, po8961, po8962, po8963,
    po8964, po8965, po8966, po8967, po8968, po8969, po8970, po8971, po8972,
    po8973, po8974, po8975, po8976, po8977, po8978, po8979, po8980, po8981,
    po8982, po8983, po8984, po8985, po8986, po8987, po8988, po8989, po8990,
    po8991, po8992, po8993, po8994, po8995, po8996, po8997, po8998, po8999,
    po9000, po9001, po9002, po9003, po9004, po9005, po9006, po9007, po9008,
    po9009, po9010, po9011, po9012, po9013, po9014, po9015, po9016, po9017,
    po9018, po9019, po9020, po9021, po9022, po9023, po9024, po9025, po9026,
    po9027, po9028, po9029, po9030, po9031, po9032, po9033, po9034, po9035,
    po9036, po9037  );
  input  pi0000, pi0001, pi0002, pi0003, pi0004, pi0005, pi0006, pi0007,
    pi0008, pi0009, pi0010, pi0011, pi0012, pi0013, pi0014, pi0015, pi0016,
    pi0017, pi0018, pi0019, pi0020, pi0021, pi0022, pi0023, pi0024, pi0025,
    pi0026, pi0027, pi0028, pi0029, pi0030, pi0031, pi0032, pi0033, pi0034,
    pi0035, pi0036, pi0037, pi0038, pi0039, pi0040, pi0041, pi0042, pi0043,
    pi0044, pi0045, pi0046, pi0047, pi0048, pi0049, pi0050, pi0051, pi0052,
    pi0053, pi0054, pi0055, pi0056, pi0057, pi0058, pi0059, pi0060, pi0061,
    pi0062, pi0063, pi0064, pi0065, pi0066, pi0067, pi0068, pi0069, pi0070,
    pi0071, pi0072, pi0073, pi0074, pi0075, pi0076, pi0077, pi0078, pi0079,
    pi0080, pi0081, pi0082, pi0083, pi0084, pi0085, pi0086, pi0087, pi0088,
    pi0089, pi0090, pi0091, pi0092, pi0093, pi0094, pi0095, pi0096, pi0097,
    pi0098, pi0099, pi0100, pi0101, pi0102, pi0103, pi0104, pi0105, pi0106,
    pi0107, pi0108, pi0109, pi0110, pi0111, pi0112, pi0113, pi0114, pi0115,
    pi0116, pi0117, pi0118, pi0119, pi0120, pi0121, pi0122, pi0123, pi0124,
    pi0125, pi0126, pi0127, pi0128, pi0129, pi0130, pi0131, pi0132, pi0133,
    pi0134, pi0135, pi0136, pi0137, pi0138, pi0139, pi0140, pi0141, pi0142,
    pi0143, pi0144, pi0145, pi0146, pi0147, pi0148, pi0149, pi0150, pi0151,
    pi0152, pi0153, pi0154, pi0155, pi0156, pi0157, pi0158, pi0159, pi0160,
    pi0161, pi0162, pi0163, pi0164, pi0165, pi0166, pi0167, pi0168, pi0169,
    pi0170, pi0171, pi0172, pi0173, pi0174, pi0175, pi0176, pi0177, pi0178,
    pi0179, pi0180, pi0181, pi0182, pi0183, pi0184, pi0185, pi0186, pi0187,
    pi0188, pi0189, pi0190, pi0191, pi0192, pi0193, pi0194, pi0195, pi0196,
    pi0197, pi0198, pi0199, pi0200, pi0201, pi0202, pi0203, pi0204, pi0205,
    pi0206, pi0207, pi0208, pi0209, pi0210, pi0211, pi0212, pi0213, pi0214,
    pi0215, pi0216, pi0217, pi0218, pi0219, pi0220, pi0221, pi0222, pi0223,
    pi0224, pi0225, pi0226, pi0227, pi0228, pi0229, pi0230, pi0231, pi0232,
    pi0233, pi0234, pi0235, pi0236, pi0237, pi0238, pi0239, pi0240, pi0241,
    pi0242, pi0243, pi0244, pi0245, pi0246, pi0247, pi0248, pi0249, pi0250,
    pi0251, pi0252, pi0253, pi0254, pi0255, pi0256, pi0257, pi0258, pi0259,
    pi0260, pi0261, pi0262, pi0263, pi0264, pi0265, pi0266, pi0267, pi0268,
    pi0269, pi0270, pi0271, pi0272, pi0273, pi0274, pi0275, pi0276, pi0277,
    pi0278, pi0279, pi0280, pi0281, pi0282, pi0283, pi0284, pi0285, pi0286,
    pi0287, pi0288, pi0289, pi0290, pi0291, pi0292, pi0293, pi0294, pi0295,
    pi0296, pi0297, pi0298, pi0299, pi0300, pi0301, pi0302, pi0303, pi0304,
    pi0305, pi0306, pi0307, pi0308, pi0309, pi0310, pi0311, pi0312, pi0313,
    pi0314, pi0315, pi0316, pi0317, pi0318, pi0319, pi0320, pi0321, pi0322,
    pi0323, pi0324, pi0325, pi0326, pi0327, pi0328, pi0329, pi0330, pi0331,
    pi0332, pi0333, pi0334, pi0335, pi0336, pi0337, pi0338, pi0339, pi0340,
    pi0341, pi0342, pi0343, pi0344, pi0345, pi0346, pi0347, pi0348, pi0349,
    pi0350, pi0351, pi0352, pi0353, pi0354, pi0355, pi0356, pi0357, pi0358,
    pi0359, pi0360, pi0361, pi0362, pi0363, pi0364, pi0365, pi0366, pi0367,
    pi0368, pi0369, pi0370, pi0371, pi0372, pi0373, pi0374, pi0375, pi0376,
    pi0377, pi0378, pi0379, pi0380, pi0381, pi0382, pi0383, pi0384, pi0385,
    pi0386, pi0387, pi0388, pi0389, pi0390, pi0391, pi0392, pi0393, pi0394,
    pi0395, pi0396, pi0397, pi0398, pi0399, pi0400, pi0401, pi0402, pi0403,
    pi0404, pi0405, pi0406, pi0407, pi0408, pi0409, pi0410, pi0411, pi0412,
    pi0413, pi0414, pi0415, pi0416, pi0417, pi0418, pi0419, pi0420, pi0421,
    pi0422, pi0423, pi0424, pi0425, pi0426, pi0427, pi0428, pi0429, pi0430,
    pi0431, pi0432, pi0433, pi0434, pi0435, pi0436, pi0437, pi0438, pi0439,
    pi0440, pi0441, pi0442, pi0443, pi0444, pi0445, pi0446, pi0447, pi0448,
    pi0449, pi0450, pi0451, pi0452, pi0453, pi0454, pi0455, pi0456, pi0457,
    pi0458, pi0459, pi0460, pi0461, pi0462, pi0463, pi0464, pi0465, pi0466,
    pi0467, pi0468, pi0469, pi0470, pi0471, pi0472, pi0473, pi0474, pi0475,
    pi0476, pi0477, pi0478, pi0479, pi0480, pi0481, pi0482, pi0483, pi0484,
    pi0485, pi0486, pi0487, pi0488, pi0489, pi0490, pi0491, pi0492, pi0493,
    pi0494, pi0495, pi0496, pi0497, pi0498, pi0499, pi0500, pi0501, pi0502,
    pi0503, pi0504, pi0505, pi0506, pi0507, pi0508, pi0509, pi0510, pi0511,
    pi0512, pi0513, pi0514, pi0515, pi0516, pi0517, pi0518, pi0519, pi0520,
    pi0521, pi0522, pi0523, pi0524, pi0525, pi0526, pi0527, pi0528, pi0529,
    pi0530, pi0531, pi0532, pi0533, pi0534, pi0535, pi0536, pi0537, pi0538,
    pi0539, pi0540, pi0541, pi0542, pi0543, pi0544, pi0545, pi0546, pi0547,
    pi0548, pi0549, pi0550, pi0551, pi0552, pi0553, pi0554, pi0555, pi0556,
    pi0557, pi0558, pi0559, pi0560, pi0561, pi0562, pi0563, pi0564, pi0565,
    pi0566, pi0567, pi0568, pi0569, pi0570, pi0571, pi0572, pi0573, pi0574,
    pi0575, pi0576, pi0577, pi0578, pi0579, pi0580, pi0581, pi0582, pi0583,
    pi0584, pi0585, pi0586, pi0587, pi0588, pi0589, pi0590, pi0591, pi0592,
    pi0593, pi0594, pi0595, pi0596, pi0597, pi0598, pi0599, pi0600, pi0601,
    pi0602, pi0603, pi0604, pi0605, pi0606, pi0607, pi0608, pi0609, pi0610,
    pi0611, pi0612, pi0613, pi0614, pi0615, pi0616, pi0617, pi0618, pi0619,
    pi0620, pi0621, pi0622, pi0623, pi0624, pi0625, pi0626, pi0627, pi0628,
    pi0629, pi0630, pi0631, pi0632, pi0633, pi0634, pi0635, pi0636, pi0637,
    pi0638, pi0639, pi0640, pi0641, pi0642, pi0643, pi0644, pi0645, pi0646,
    pi0647, pi0648, pi0649, pi0650, pi0651, pi0652, pi0653, pi0654, pi0655,
    pi0656, pi0657, pi0658, pi0659, pi0660, pi0661, pi0662, pi0663, pi0664,
    pi0665, pi0666, pi0667, pi0668, pi0669, pi0670, pi0671, pi0672, pi0673,
    pi0674, pi0675, pi0676, pi0677, pi0678, pi0679, pi0680, pi0681, pi0682,
    pi0683, pi0684, pi0685, pi0686, pi0687, pi0688, pi0689, pi0690, pi0691,
    pi0692, pi0693, pi0694, pi0695, pi0696, pi0697, pi0698, pi0699, pi0700,
    pi0701, pi0702, pi0703, pi0704, pi0705, pi0706, pi0707, pi0708, pi0709,
    pi0710, pi0711, pi0712, pi0713, pi0714, pi0715, pi0716, pi0717, pi0718,
    pi0719, pi0720, pi0721, pi0722, pi0723, pi0724, pi0725, pi0726, pi0727,
    pi0728, pi0729, pi0730, pi0731, pi0732, pi0733, pi0734, pi0735, pi0736,
    pi0737, pi0738, pi0739, pi0740, pi0741, pi0742, pi0743, pi0744, pi0745,
    pi0746, pi0747, pi0748, pi0749, pi0750, pi0751, pi0752, pi0753, pi0754,
    pi0755, pi0756, pi0757, pi0758, pi0759, pi0760, pi0761, pi0762, pi0763,
    pi0764, pi0765, pi0766, pi0767, pi0768, pi0769, pi0770, pi0771, pi0772,
    pi0773, pi0774, pi0775, pi0776, pi0777, pi0778, pi0779, pi0780, pi0781,
    pi0782, pi0783, pi0784, pi0785, pi0786, pi0787, pi0788, pi0789, pi0790,
    pi0791, pi0792, pi0793, pi0794, pi0795, pi0796, pi0797, pi0798, pi0799,
    pi0800, pi0801, pi0802, pi0803, pi0804, pi0805, pi0806, pi0807, pi0808,
    pi0809, pi0810, pi0811, pi0812, pi0813, pi0814, pi0815, pi0816, pi0817,
    pi0818, pi0819, pi0820, pi0821, pi0822, pi0823, pi0824, pi0825, pi0826,
    pi0827, pi0828, pi0829, pi0830, pi0831, pi0832, pi0833, pi0834, pi0835,
    pi0836, pi0837, pi0838, pi0839, pi0840, pi0841, pi0842, pi0843, pi0844,
    pi0845, pi0846, pi0847, pi0848, pi0849, pi0850, pi0851, pi0852, pi0853,
    pi0854, pi0855, pi0856, pi0857, pi0858, pi0859, pi0860, pi0861, pi0862,
    pi0863, pi0864, pi0865, pi0866, pi0867, pi0868, pi0869, pi0870, pi0871,
    pi0872, pi0873, pi0874, pi0875, pi0876, pi0877, pi0878, pi0879, pi0880,
    pi0881, pi0882, pi0883, pi0884, pi0885, pi0886, pi0887, pi0888, pi0889,
    pi0890, pi0891, pi0892, pi0893, pi0894, pi0895, pi0896, pi0897, pi0898,
    pi0899, pi0900, pi0901, pi0902, pi0903, pi0904, pi0905, pi0906, pi0907,
    pi0908, pi0909, pi0910, pi0911, pi0912, pi0913, pi0914, pi0915, pi0916,
    pi0917, pi0918, pi0919, pi0920, pi0921, pi0922, pi0923, pi0924, pi0925,
    pi0926, pi0927, pi0928, pi0929, pi0930, pi0931, pi0932, pi0933, pi0934,
    pi0935, pi0936, pi0937, pi0938, pi0939, pi0940, pi0941, pi0942, pi0943,
    pi0944, pi0945, pi0946, pi0947, pi0948, pi0949, pi0950, pi0951, pi0952,
    pi0953, pi0954, pi0955, pi0956, pi0957, pi0958, pi0959, pi0960, pi0961,
    pi0962, pi0963, pi0964, pi0965, pi0966, pi0967, pi0968, pi0969, pi0970,
    pi0971, pi0972, pi0973, pi0974, pi0975, pi0976, pi0977, pi0978, pi0979,
    pi0980, pi0981, pi0982, pi0983, pi0984, pi0985, pi0986, pi0987, pi0988,
    pi0989, pi0990, pi0991, pi0992, pi0993, pi0994, pi0995, pi0996, pi0997,
    pi0998, pi0999, pi1000, pi1001, pi1002, pi1003, pi1004, pi1005, pi1006,
    pi1007, pi1008, pi1009, pi1010, pi1011, pi1012, pi1013, pi1014, pi1015,
    pi1016, pi1017, pi1018, pi1019, pi1020, pi1021, pi1022, pi1023, pi1024,
    pi1025, pi1026, pi1027, pi1028, pi1029, pi1030, pi1031, pi1032, pi1033,
    pi1034, pi1035, pi1036, pi1037, pi1038, pi1039, pi1040, pi1041, pi1042,
    pi1043, pi1044, pi1045, pi1046, pi1047, pi1048, pi1049, pi1050, pi1051,
    pi1052, pi1053, pi1054, pi1055, pi1056, pi1057, pi1058, pi1059, pi1060,
    pi1061, pi1062, pi1063, pi1064, pi1065, pi1066, pi1067, pi1068, pi1069,
    pi1070, pi1071, pi1072, pi1073, pi1074, pi1075, pi1076, pi1077, pi1078,
    pi1079, pi1080, pi1081, pi1082, pi1083, pi1084, pi1085, pi1086, pi1087,
    pi1088, pi1089, pi1090, pi1091, pi1092, pi1093, pi1094, pi1095, pi1096,
    pi1097, pi1098, pi1099, pi1100, pi1101, pi1102, pi1103, pi1104, pi1105,
    pi1106, pi1107, pi1108, pi1109, pi1110, pi1111, pi1112, pi1113, pi1114,
    pi1115, pi1116, pi1117, pi1118, pi1119, pi1120, pi1121, pi1122, pi1123,
    pi1124, pi1125, pi1126, pi1127, pi1128, pi1129, pi1130, pi1131, pi1132,
    pi1133, pi1134, pi1135, pi1136, pi1137, pi1138, pi1139, pi1140, pi1141,
    pi1142, pi1143, pi1144, pi1145, pi1146, pi1147, pi1148, pi1149, pi1150,
    pi1151, pi1152, pi1153, pi1154, pi1155, pi1156, pi1157, pi1158, pi1159,
    pi1160, pi1161, pi1162, pi1163, pi1164, pi1165, pi1166, pi1167, pi1168,
    pi1169, pi1170, pi1171, pi1172, pi1173, pi1174, pi1175, pi1176, pi1177,
    pi1178, pi1179, pi1180, pi1181, pi1182, pi1183, pi1184, pi1185, pi1186,
    pi1187, pi1188, pi1189, pi1190, pi1191, pi1192, pi1193, pi1194, pi1195,
    pi1196, pi1197, pi1198, pi1199, pi1200, pi1201, pi1202, pi1203, pi1204,
    pi1205, pi1206, pi1207, pi1208, pi1209, pi1210, pi1211, pi1212, pi1213,
    pi1214, pi1215, pi1216, pi1217, pi1218, pi1219, pi1220, pi1221, pi1222,
    pi1223, pi1224, pi1225, pi1226, pi1227, pi1228, pi1229, pi1230, pi1231,
    pi1232, pi1233, pi1234, pi1235, pi1236, pi1237, pi1238, pi1239, pi1240,
    pi1241, pi1242, pi1243, pi1244, pi1245, pi1246, pi1247, pi1248, pi1249,
    pi1250, pi1251, pi1252, pi1253, pi1254, pi1255, pi1256, pi1257, pi1258,
    pi1259, pi1260, pi1261, pi1262, pi1263, pi1264, pi1265, pi1266, pi1267,
    pi1268, pi1269, pi1270, pi1271, pi1272, pi1273, pi1274, pi1275, pi1276,
    pi1277, pi1278, pi1279, pi1280, pi1281, pi1282, pi1283, pi1284, pi1285,
    pi1286, pi1287, pi1288, pi1289, pi1290, pi1291, pi1292, pi1293, pi1294,
    pi1295, pi1296, pi1297, pi1298, pi1299, pi1300, pi1301, pi1302, pi1303,
    pi1304, pi1305, pi1306, pi1307, pi1308, pi1309, pi1310, pi1311, pi1312,
    pi1313, pi1314, pi1315, pi1316, pi1317, pi1318, pi1319, pi1320, pi1321,
    pi1322, pi1323, pi1324, pi1325, pi1326, pi1327, pi1328, pi1329, pi1330,
    pi1331, pi1332, pi1333, pi1334, pi1335, pi1336, pi1337, pi1338, pi1339,
    pi1340, pi1341, pi1342, pi1343, pi1344, pi1345, pi1346, pi1347, pi1348,
    pi1349, pi1350, pi1351, pi1352, pi1353, pi1354, pi1355, pi1356, pi1357,
    pi1358, pi1359, pi1360, pi1361, pi1362, pi1363, pi1364, pi1365, pi1366,
    pi1367, pi1368, pi1369, pi1370, pi1371, pi1372, pi1373, pi1374, pi1375,
    pi1376, pi1377, pi1378, pi1379, pi1380, pi1381, pi1382, pi1383, pi1384,
    pi1385, pi1386, pi1387, pi1388, pi1389, pi1390, pi1391, pi1392, pi1393,
    pi1394, pi1395, pi1396, pi1397, pi1398, pi1399, pi1400, pi1401, pi1402,
    pi1403, pi1404, pi1405, pi1406, pi1407, pi1408, pi1409, pi1410, pi1411,
    pi1412, pi1413, pi1414, pi1415, pi1416, pi1417, pi1418, pi1419, pi1420,
    pi1421, pi1422, pi1423, pi1424, pi1425, pi1426, pi1427, pi1428, pi1429,
    pi1430, pi1431, pi1432, pi1433, pi1434, pi1435, pi1436, pi1437, pi1438,
    pi1439, pi1440, pi1441, pi1442, pi1443, pi1444, pi1445, pi1446, pi1447,
    pi1448, pi1449, pi1450, pi1451, pi1452, pi1453, pi1454, pi1455, pi1456,
    pi1457, pi1458, pi1459, pi1460, pi1461, pi1462, pi1463, pi1464, pi1465,
    pi1466, pi1467, pi1468, pi1469, pi1470, pi1471, pi1472, pi1473, pi1474,
    pi1475, pi1476, pi1477, pi1478, pi1479, pi1480, pi1481, pi1482, pi1483,
    pi1484, pi1485, pi1486, pi1487, pi1488, pi1489, pi1490, pi1491, pi1492,
    pi1493, pi1494, pi1495, pi1496, pi1497, pi1498, pi1499, pi1500, pi1501,
    pi1502, pi1503, pi1504, pi1505, pi1506, pi1507, pi1508, pi1509, pi1510,
    pi1511, pi1512, pi1513, pi1514, pi1515, pi1516, pi1517, pi1518, pi1519,
    pi1520, pi1521, pi1522, pi1523, pi1524, pi1525, pi1526, pi1527, pi1528,
    pi1529, pi1530, pi1531, pi1532, pi1533, pi1534, pi1535, pi1536, pi1537,
    pi1538, pi1539, pi1540, pi1541, pi1542, pi1543, pi1544, pi1545, pi1546,
    pi1547, pi1548, pi1549, pi1550, pi1551, pi1552, pi1553, pi1554, pi1555,
    pi1556, pi1557, pi1558, pi1559, pi1560, pi1561, pi1562, pi1563, pi1564,
    pi1565, pi1566, pi1567, pi1568, pi1569, pi1570, pi1571, pi1572, pi1573,
    pi1574, pi1575, pi1576, pi1577, pi1578, pi1579, pi1580, pi1581, pi1582,
    pi1583, pi1584, pi1585, pi1586, pi1587, pi1588, pi1589, pi1590, pi1591,
    pi1592, pi1593, pi1594, pi1595, pi1596, pi1597, pi1598, pi1599, pi1600,
    pi1601, pi1602, pi1603, pi1604, pi1605, pi1606, pi1607, pi1608, pi1609,
    pi1610, pi1611, pi1612, pi1613, pi1614, pi1615, pi1616, pi1617, pi1618,
    pi1619, pi1620, pi1621, pi1622, pi1623, pi1624, pi1625, pi1626, pi1627,
    pi1628, pi1629, pi1630, pi1631, pi1632, pi1633, pi1634, pi1635, pi1636,
    pi1637, pi1638, pi1639, pi1640, pi1641, pi1642, pi1643, pi1644, pi1645,
    pi1646, pi1647, pi1648, pi1649, pi1650, pi1651, pi1652, pi1653, pi1654,
    pi1655, pi1656, pi1657, pi1658, pi1659, pi1660, pi1661, pi1662, pi1663,
    pi1664, pi1665, pi1666, pi1667, pi1668, pi1669, pi1670, pi1671, pi1672,
    pi1673, pi1674, pi1675, pi1676, pi1677, pi1678, pi1679, pi1680, pi1681,
    pi1682, pi1683, pi1684, pi1685, pi1686, pi1687, pi1688, pi1689, pi1690,
    pi1691, pi1692, pi1693, pi1694, pi1695, pi1696, pi1697, pi1698, pi1699,
    pi1700, pi1701, pi1702, pi1703, pi1704, pi1705, pi1706, pi1707, pi1708,
    pi1709, pi1710, pi1711, pi1712, pi1713, pi1714, pi1715, pi1716, pi1717,
    pi1718, pi1719, pi1720, pi1721, pi1722, pi1723, pi1724, pi1725, pi1726,
    pi1727, pi1728, pi1729, pi1730, pi1731, pi1732, pi1733, pi1734, pi1735,
    pi1736, pi1737, pi1738, pi1739, pi1740, pi1741, pi1742, pi1743, pi1744,
    pi1745, pi1746, pi1747, pi1748, pi1749, pi1750, pi1751, pi1752, pi1753,
    pi1754, pi1755, pi1756, pi1757, pi1758, pi1759, pi1760, pi1761, pi1762,
    pi1763, pi1764, pi1765, pi1766, pi1767, pi1768, pi1769, pi1770, pi1771,
    pi1772, pi1773, pi1774, pi1775, pi1776, pi1777, pi1778, pi1779, pi1780,
    pi1781, pi1782, pi1783, pi1784, pi1785, pi1786, pi1787, pi1788, pi1789,
    pi1790, pi1791, pi1792, pi1793, pi1794, pi1795, pi1796, pi1797, pi1798,
    pi1799, pi1800, pi1801, pi1802, pi1803, pi1804, pi1805, pi1806, pi1807,
    pi1808, pi1809, pi1810, pi1811, pi1812, pi1813, pi1814, pi1815, pi1816,
    pi1817, pi1818, pi1819, pi1820, pi1821, pi1822, pi1823, pi1824, pi1825,
    pi1826, pi1827, pi1828, pi1829, pi1830, pi1831, pi1832, pi1833, pi1834,
    pi1835, pi1836, pi1837, pi1838, pi1839, pi1840, pi1841, pi1842, pi1843,
    pi1844, pi1845, pi1846, pi1847, pi1848, pi1849, pi1850, pi1851, pi1852,
    pi1853, pi1854, pi1855, pi1856, pi1857, pi1858, pi1859, pi1860, pi1861,
    pi1862, pi1863, pi1864, pi1865, pi1866, pi1867, pi1868, pi1869, pi1870,
    pi1871, pi1872, pi1873, pi1874, pi1875, pi1876, pi1877, pi1878, pi1879,
    pi1880, pi1881, pi1882, pi1883, pi1884, pi1885, pi1886, pi1887, pi1888,
    pi1889, pi1890, pi1891, pi1892, pi1893, pi1894, pi1895, pi1896, pi1897,
    pi1898, pi1899, pi1900, pi1901, pi1902, pi1903, pi1904, pi1905, pi1906,
    pi1907, pi1908, pi1909, pi1910, pi1911, pi1912, pi1913, pi1914, pi1915,
    pi1916, pi1917, pi1918, pi1919, pi1920, pi1921, pi1922, pi1923, pi1924,
    pi1925, pi1926, pi1927, pi1928, pi1929, pi1930, pi1931, pi1932, pi1933,
    pi1934, pi1935, pi1936, pi1937, pi1938, pi1939, pi1940, pi1941, pi1942,
    pi1943, pi1944, pi1945, pi1946, pi1947, pi1948, pi1949, pi1950, pi1951,
    pi1952, pi1953, pi1954, pi1955, pi1956, pi1957, pi1958, pi1959, pi1960,
    pi1961, pi1962, pi1963, pi1964, pi1965, pi1966, pi1967, pi1968, pi1969,
    pi1970, pi1971, pi1972, pi1973, pi1974, pi1975, pi1976, pi1977, pi1978,
    pi1979, pi1980, pi1981, pi1982, pi1983, pi1984, pi1985, pi1986, pi1987,
    pi1988, pi1989, pi1990, pi1991, pi1992, pi1993, pi1994, pi1995, pi1996,
    pi1997, pi1998, pi1999, pi2000, pi2001, pi2002, pi2003, pi2004, pi2005,
    pi2006, pi2007, pi2008, pi2009, pi2010, pi2011, pi2012, pi2013, pi2014,
    pi2015, pi2016, pi2017, pi2018, pi2019, pi2020, pi2021, pi2022, pi2023,
    pi2024, pi2025, pi2026, pi2027, pi2028, pi2029, pi2030, pi2031, pi2032,
    pi2033, pi2034, pi2035, pi2036, pi2037, pi2038, pi2039, pi2040, pi2041,
    pi2042, pi2043, pi2044, pi2045, pi2046, pi2047, pi2048, pi2049, pi2050,
    pi2051, pi2052, pi2053, pi2054, pi2055, pi2056, pi2057, pi2058, pi2059,
    pi2060, pi2061, pi2062, pi2063, pi2064, pi2065, pi2066, pi2067, pi2068,
    pi2069, pi2070, pi2071, pi2072, pi2073, pi2074, pi2075, pi2076, pi2077,
    pi2078, pi2079, pi2080, pi2081, pi2082, pi2083, pi2084, pi2085, pi2086,
    pi2087, pi2088, pi2089, pi2090, pi2091, pi2092, pi2093, pi2094, pi2095,
    pi2096, pi2097, pi2098, pi2099, pi2100, pi2101, pi2102, pi2103, pi2104,
    pi2105, pi2106, pi2107, pi2108, pi2109, pi2110, pi2111, pi2112, pi2113,
    pi2114, pi2115, pi2116, pi2117, pi2118, pi2119, pi2120, pi2121, pi2122,
    pi2123, pi2124, pi2125, pi2126, pi2127, pi2128, pi2129, pi2130, pi2131,
    pi2132, pi2133, pi2134, pi2135, pi2136, pi2137, pi2138, pi2139, pi2140,
    pi2141, pi2142, pi2143, pi2144, pi2145, pi2146, pi2147, pi2148, pi2149,
    pi2150, pi2151, pi2152, pi2153, pi2154, pi2155, pi2156, pi2157, pi2158,
    pi2159, pi2160, pi2161, pi2162, pi2163, pi2164, pi2165, pi2166, pi2167,
    pi2168, pi2169, pi2170, pi2171, pi2172, pi2173, pi2174, pi2175, pi2176,
    pi2177, pi2178, pi2179, pi2180, pi2181, pi2182, pi2183, pi2184, pi2185,
    pi2186, pi2187, pi2188, pi2189, pi2190, pi2191, pi2192, pi2193, pi2194,
    pi2195, pi2196, pi2197, pi2198, pi2199, pi2200, pi2201, pi2202, pi2203,
    pi2204, pi2205, pi2206, pi2207, pi2208, pi2209, pi2210, pi2211, pi2212,
    pi2213, pi2214, pi2215, pi2216, pi2217, pi2218, pi2219, pi2220, pi2221,
    pi2222, pi2223, pi2224, pi2225, pi2226, pi2227, pi2228, pi2229, pi2230,
    pi2231, pi2232, pi2233, pi2234, pi2235, pi2236, pi2237, pi2238, pi2239,
    pi2240, pi2241, pi2242, pi2243, pi2244, pi2245, pi2246, pi2247, pi2248,
    pi2249, pi2250, pi2251, pi2252, pi2253, pi2254, pi2255, pi2256, pi2257,
    pi2258, pi2259, pi2260, pi2261, pi2262, pi2263, pi2264, pi2265, pi2266,
    pi2267, pi2268, pi2269, pi2270, pi2271, pi2272, pi2273, pi2274, pi2275,
    pi2276, pi2277, pi2278, pi2279, pi2280, pi2281, pi2282, pi2283, pi2284,
    pi2285, pi2286, pi2287, pi2288, pi2289, pi2290, pi2291, pi2292, pi2293,
    pi2294, pi2295, pi2296, pi2297, pi2298, pi2299, pi2300, pi2301, pi2302,
    pi2303, pi2304, pi2305, pi2306, pi2307, pi2308, pi2309, pi2310, pi2311,
    pi2312, pi2313, pi2314, pi2315, pi2316, pi2317, pi2318, pi2319, pi2320,
    pi2321, pi2322, pi2323, pi2324, pi2325, pi2326, pi2327, pi2328, pi2329,
    pi2330, pi2331, pi2332, pi2333, pi2334, pi2335, pi2336, pi2337, pi2338,
    pi2339, pi2340, pi2341, pi2342, pi2343, pi2344, pi2345, pi2346, pi2347,
    pi2348, pi2349, pi2350, pi2351, pi2352, pi2353, pi2354, pi2355, pi2356,
    pi2357, pi2358, pi2359, pi2360, pi2361, pi2362, pi2363, pi2364, pi2365,
    pi2366, pi2367, pi2368, pi2369, pi2370, pi2371, pi2372, pi2373, pi2374,
    pi2375, pi2376, pi2377, pi2378, pi2379, pi2380, pi2381, pi2382, pi2383,
    pi2384, pi2385, pi2386, pi2387, pi2388, pi2389, pi2390, pi2391, pi2392,
    pi2393, pi2394, pi2395, pi2396, pi2397, pi2398, pi2399, pi2400, pi2401,
    pi2402, pi2403, pi2404, pi2405, pi2406, pi2407, pi2408, pi2409, pi2410,
    pi2411, pi2412, pi2413, pi2414, pi2415, pi2416, pi2417, pi2418, pi2419,
    pi2420, pi2421, pi2422, pi2423, pi2424, pi2425, pi2426, pi2427, pi2428,
    pi2429, pi2430, pi2431, pi2432, pi2433, pi2434, pi2435, pi2436, pi2437,
    pi2438, pi2439, pi2440, pi2441, pi2442, pi2443, pi2444, pi2445, pi2446,
    pi2447, pi2448, pi2449, pi2450, pi2451, pi2452, pi2453, pi2454, pi2455,
    pi2456, pi2457, pi2458, pi2459, pi2460, pi2461, pi2462, pi2463, pi2464,
    pi2465, pi2466, pi2467, pi2468, pi2469, pi2470, pi2471, pi2472, pi2473,
    pi2474, pi2475, pi2476, pi2477, pi2478, pi2479, pi2480, pi2481, pi2482,
    pi2483, pi2484, pi2485, pi2486, pi2487, pi2488, pi2489, pi2490, pi2491,
    pi2492, pi2493, pi2494, pi2495, pi2496, pi2497, pi2498, pi2499, pi2500,
    pi2501, pi2502, pi2503, pi2504, pi2505, pi2506, pi2507, pi2508, pi2509,
    pi2510, pi2511, pi2512, pi2513, pi2514, pi2515, pi2516, pi2517, pi2518,
    pi2519, pi2520, pi2521, pi2522, pi2523, pi2524, pi2525, pi2526, pi2527,
    pi2528, pi2529, pi2530, pi2531, pi2532, pi2533, pi2534, pi2535, pi2536,
    pi2537, pi2538, pi2539, pi2540, pi2541, pi2542, pi2543, pi2544, pi2545,
    pi2546, pi2547, pi2548, pi2549, pi2550, pi2551, pi2552, pi2553, pi2554,
    pi2555, pi2556, pi2557, pi2558, pi2559, pi2560, pi2561, pi2562, pi2563,
    pi2564, pi2565, pi2566, pi2567, pi2568, pi2569, pi2570, pi2571, pi2572,
    pi2573, pi2574, pi2575, pi2576, pi2577, pi2578, pi2579, pi2580, pi2581,
    pi2582, pi2583, pi2584, pi2585, pi2586, pi2587, pi2588, pi2589, pi2590,
    pi2591, pi2592, pi2593, pi2594, pi2595, pi2596, pi2597, pi2598, pi2599,
    pi2600, pi2601, pi2602, pi2603, pi2604, pi2605, pi2606, pi2607, pi2608,
    pi2609, pi2610, pi2611, pi2612, pi2613, pi2614, pi2615, pi2616, pi2617,
    pi2618, pi2619, pi2620, pi2621, pi2622, pi2623, pi2624, pi2625, pi2626,
    pi2627, pi2628, pi2629, pi2630, pi2631, pi2632, pi2633, pi2634, pi2635,
    pi2636, pi2637, pi2638, pi2639, pi2640, pi2641, pi2642, pi2643, pi2644,
    pi2645, pi2646, pi2647, pi2648, pi2649, pi2650, pi2651, pi2652, pi2653,
    pi2654, pi2655, pi2656, pi2657, pi2658, pi2659, pi2660, pi2661, pi2662,
    pi2663, pi2664, pi2665, pi2666, pi2667, pi2668, pi2669, pi2670, pi2671,
    pi2672, pi2673, pi2674, pi2675, pi2676, pi2677, pi2678, pi2679, pi2680,
    pi2681, pi2682, pi2683, pi2684, pi2685, pi2686, pi2687, pi2688, pi2689,
    pi2690, pi2691, pi2692, pi2693, pi2694, pi2695, pi2696, pi2697, pi2698,
    pi2699, pi2700, pi2701, pi2702, pi2703, pi2704, pi2705, pi2706, pi2707,
    pi2708, pi2709, pi2710, pi2711, pi2712, pi2713, pi2714, pi2715, pi2716,
    pi2717, pi2718, pi2719, pi2720, pi2721, pi2722, pi2723, pi2724, pi2725,
    pi2726, pi2727, pi2728, pi2729, pi2730, pi2731, pi2732, pi2733, pi2734,
    pi2735, pi2736, pi2737, pi2738, pi2739, pi2740, pi2741, pi2742, pi2743,
    pi2744, pi2745, pi2746, pi2747, pi2748, pi2749, pi2750, pi2751, pi2752,
    pi2753, pi2754, pi2755, pi2756, pi2757, pi2758, pi2759, pi2760, pi2761,
    pi2762, pi2763, pi2764, pi2765, pi2766, pi2767, pi2768, pi2769, pi2770,
    pi2771, pi2772, pi2773, pi2774, pi2775, pi2776, pi2777, pi2778, pi2779,
    pi2780, pi2781, pi2782, pi2783, pi2784, pi2785, pi2786, pi2787, pi2788,
    pi2789, pi2790, pi2791, pi2792, pi2793, pi2794, pi2795, pi2796, pi2797,
    pi2798, pi2799, pi2800, pi2801, pi2802, pi2803, pi2804, pi2805, pi2806,
    pi2807, pi2808, pi2809, pi2810, pi2811, pi2812, pi2813, pi2814, pi2815,
    pi2816, pi2817, pi2818, pi2819, pi2820, pi2821, pi2822, pi2823, pi2824,
    pi2825, pi2826, pi2827, pi2828, pi2829, pi2830, pi2831, pi2832, pi2833,
    pi2834, pi2835, pi2836, pi2837, pi2838, pi2839, pi2840, pi2841, pi2842,
    pi2843, pi2844, pi2845, pi2846, pi2847, pi2848, pi2849, pi2850, pi2851,
    pi2852, pi2853, pi2854, pi2855, pi2856, pi2857, pi2858, pi2859, pi2860,
    pi2861, pi2862, pi2863, pi2864, pi2865, pi2866, pi2867, pi2868, pi2869,
    pi2870, pi2871, pi2872, pi2873, pi2874, pi2875, pi2876, pi2877, pi2878,
    pi2879, pi2880, pi2881, pi2882, pi2883, pi2884, pi2885, pi2886, pi2887,
    pi2888, pi2889, pi2890, pi2891, pi2892, pi2893, pi2894, pi2895, pi2896,
    pi2897, pi2898, pi2899, pi2900, pi2901, pi2902, pi2903, pi2904, pi2905,
    pi2906, pi2907, pi2908, pi2909, pi2910, pi2911, pi2912, pi2913, pi2914,
    pi2915, pi2916, pi2917, pi2918, pi2919, pi2920, pi2921, pi2922, pi2923,
    pi2924, pi2925, pi2926, pi2927, pi2928, pi2929, pi2930, pi2931, pi2932,
    pi2933, pi2934, pi2935, pi2936, pi2937, pi2938, pi2939, pi2940, pi2941,
    pi2942, pi2943, pi2944, pi2945, pi2946, pi2947, pi2948, pi2949, pi2950,
    pi2951, pi2952, pi2953, pi2954, pi2955, pi2956, pi2957, pi2958, pi2959,
    pi2960, pi2961, pi2962, pi2963, pi2964, pi2965, pi2966, pi2967, pi2968,
    pi2969, pi2970, pi2971, pi2972, pi2973, pi2974, pi2975, pi2976, pi2977,
    pi2978, pi2979, pi2980, pi2981, pi2982, pi2983, pi2984, pi2985, pi2986,
    pi2987, pi2988, pi2989, pi2990, pi2991, pi2992, pi2993, pi2994, pi2995,
    pi2996, pi2997, pi2998, pi2999, pi3000, pi3001, pi3002, pi3003, pi3004,
    pi3005, pi3006, pi3007, pi3008, pi3009, pi3010, pi3011, pi3012, pi3013,
    pi3014, pi3015, pi3016, pi3017, pi3018, pi3019, pi3020, pi3021, pi3022,
    pi3023, pi3024, pi3025, pi3026, pi3027, pi3028, pi3029, pi3030, pi3031,
    pi3032, pi3033, pi3034, pi3035, pi3036, pi3037, pi3038, pi3039, pi3040,
    pi3041, pi3042, pi3043, pi3044, pi3045, pi3046, pi3047, pi3048, pi3049,
    pi3050, pi3051, pi3052, pi3053, pi3054, pi3055, pi3056, pi3057, pi3058,
    pi3059, pi3060, pi3061, pi3062, pi3063, pi3064, pi3065, pi3066, pi3067,
    pi3068, pi3069, pi3070, pi3071, pi3072, pi3073, pi3074, pi3075, pi3076,
    pi3077, pi3078, pi3079, pi3080, pi3081, pi3082, pi3083, pi3084, pi3085,
    pi3086, pi3087, pi3088, pi3089, pi3090, pi3091, pi3092, pi3093, pi3094,
    pi3095, pi3096, pi3097, pi3098, pi3099, pi3100, pi3101, pi3102, pi3103,
    pi3104, pi3105, pi3106, pi3107, pi3108, pi3109, pi3110, pi3111, pi3112,
    pi3113, pi3114, pi3115, pi3116, pi3117, pi3118, pi3119, pi3120, pi3121,
    pi3122, pi3123, pi3124, pi3125, pi3126, pi3127, pi3128, pi3129, pi3130,
    pi3131, pi3132, pi3133, pi3134, pi3135, pi3136, pi3137, pi3138, pi3139,
    pi3140, pi3141, pi3142, pi3143, pi3144, pi3145, pi3146, pi3147, pi3148,
    pi3149, pi3150, pi3151, pi3152, pi3153, pi3154, pi3155, pi3156, pi3157,
    pi3158, pi3159, pi3160, pi3161, pi3162, pi3163, pi3164, pi3165, pi3166,
    pi3167, pi3168, pi3169, pi3170, pi3171, pi3172, pi3173, pi3174, pi3175,
    pi3176, pi3177, pi3178, pi3179, pi3180, pi3181, pi3182, pi3183, pi3184,
    pi3185, pi3186, pi3187, pi3188, pi3189, pi3190, pi3191, pi3192, pi3193,
    pi3194, pi3195, pi3196, pi3197, pi3198, pi3199, pi3200, pi3201, pi3202,
    pi3203, pi3204, pi3205, pi3206, pi3207, pi3208, pi3209, pi3210, pi3211,
    pi3212, pi3213, pi3214, pi3215, pi3216, pi3217, pi3218, pi3219, pi3220,
    pi3221, pi3222, pi3223, pi3224, pi3225, pi3226, pi3227, pi3228, pi3229,
    pi3230, pi3231, pi3232, pi3233, pi3234, pi3235, pi3236, pi3237, pi3238,
    pi3239, pi3240, pi3241, pi3242, pi3243, pi3244, pi3245, pi3246, pi3247,
    pi3248, pi3249, pi3250, pi3251, pi3252, pi3253, pi3254, pi3255, pi3256,
    pi3257, pi3258, pi3259, pi3260, pi3261, pi3262, pi3263, pi3264, pi3265,
    pi3266, pi3267, pi3268, pi3269, pi3270, pi3271, pi3272, pi3273, pi3274,
    pi3275, pi3276, pi3277, pi3278, pi3279, pi3280, pi3281, pi3282, pi3283,
    pi3284, pi3285, pi3286, pi3287, pi3288, pi3289, pi3290, pi3291, pi3292,
    pi3293, pi3294, pi3295, pi3296, pi3297, pi3298, pi3299, pi3300, pi3301,
    pi3302, pi3303, pi3304, pi3305, pi3306, pi3307, pi3308, pi3309, pi3310,
    pi3311, pi3312, pi3313, pi3314, pi3315, pi3316, pi3317, pi3318, pi3319,
    pi3320, pi3321, pi3322, pi3323, pi3324, pi3325, pi3326, pi3327, pi3328,
    pi3329, pi3330, pi3331, pi3332, pi3333, pi3334, pi3335, pi3336, pi3337,
    pi3338, pi3339, pi3340, pi3341, pi3342, pi3343, pi3344, pi3345, pi3346,
    pi3347, pi3348, pi3349, pi3350, pi3351, pi3352, pi3353, pi3354, pi3355,
    pi3356, pi3357, pi3358, pi3359, pi3360, pi3361, pi3362, pi3363, pi3364,
    pi3365, pi3366, pi3367, pi3368, pi3369, pi3370, pi3371, pi3372, pi3373,
    pi3374, pi3375, pi3376, pi3377, pi3378, pi3379, pi3380, pi3381, pi3382,
    pi3383, pi3384, pi3385, pi3386, pi3387, pi3388, pi3389, pi3390, pi3391,
    pi3392, pi3393, pi3394, pi3395, pi3396, pi3397, pi3398, pi3399, pi3400,
    pi3401, pi3402, pi3403, pi3404, pi3405, pi3406, pi3407, pi3408, pi3409,
    pi3410, pi3411, pi3412, pi3413, pi3414, pi3415, pi3416, pi3417, pi3418,
    pi3419, pi3420, pi3421, pi3422, pi3423, pi3424, pi3425, pi3426, pi3427,
    pi3428, pi3429, pi3430, pi3431, pi3432, pi3433, pi3434, pi3435, pi3436,
    pi3437, pi3438, pi3439, pi3440, pi3441, pi3442, pi3443, pi3444, pi3445,
    pi3446, pi3447, pi3448, pi3449, pi3450, pi3451, pi3452, pi3453, pi3454,
    pi3455, pi3456, pi3457, pi3458, pi3459, pi3460, pi3461, pi3462, pi3463,
    pi3464, pi3465, pi3466, pi3467, pi3468, pi3469, pi3470, pi3471, pi3472,
    pi3473, pi3474, pi3475, pi3476, pi3477, pi3478, pi3479, pi3480, pi3481,
    pi3482, pi3483, pi3484, pi3485, pi3486, pi3487, pi3488, pi3489, pi3490,
    pi3491, pi3492, pi3493, pi3494, pi3495, pi3496, pi3497, pi3498, pi3499,
    pi3500, pi3501, pi3502, pi3503, pi3504, pi3505, pi3506, pi3507, pi3508,
    pi3509, pi3510, pi3511, pi3512, pi3513, pi3514, pi3515, pi3516, pi3517,
    pi3518, pi3519, pi3520, pi3521, pi3522, pi3523, pi3524, pi3525, pi3526,
    pi3527, pi3528, pi3529, pi3530, pi3531, pi3532, pi3533, pi3534, pi3535,
    pi3536, pi3537, pi3538, pi3539, pi3540, pi3541, pi3542, pi3543, pi3544,
    pi3545, pi3546, pi3547, pi3548, pi3549, pi3550, pi3551, pi3552, pi3553,
    pi3554, pi3555, pi3556, pi3557, pi3558, pi3559, pi3560, pi3561, pi3562,
    pi3563, pi3564, pi3565, pi3566, pi3567, pi3568, pi3569, pi3570, pi3571,
    pi3572, pi3573, pi3574, pi3575, pi3576, pi3577, pi3578, pi3579, pi3580,
    pi3581, pi3582, pi3583, pi3584, pi3585, pi3586, pi3587, pi3588, pi3589,
    pi3590, pi3591, pi3592, pi3593, pi3594, pi3595, pi3596, pi3597, pi3598,
    pi3599, pi3600, pi3601, pi3602, pi3603, pi3604, pi3605, pi3606, pi3607,
    pi3608, pi3609, pi3610, pi3611, pi3612, pi3613, pi3614, pi3615, pi3616,
    pi3617, pi3618, pi3619, pi3620, pi3621, pi3622, pi3623, pi3624, pi3625,
    pi3626, pi3627, pi3628, pi3629, pi3630, pi3631, pi3632, pi3633, pi3634,
    pi3635, pi3636, pi3637, pi3638, pi3639, pi3640, pi3641, pi3642, pi3643,
    pi3644, pi3645, pi3646, pi3647, pi3648, pi3649, pi3650, pi3651, pi3652,
    pi3653, pi3654, pi3655, pi3656, pi3657, pi3658, pi3659, pi3660, pi3661,
    pi3662, pi3663, pi3664, pi3665, pi3666, pi3667, pi3668, pi3669, pi3670,
    pi3671, pi3672, pi3673, pi3674, pi3675, pi3676, pi3677, pi3678, pi3679,
    pi3680, pi3681, pi3682, pi3683, pi3684, pi3685, pi3686, pi3687, pi3688,
    pi3689, pi3690, pi3691, pi3692, pi3693, pi3694, pi3695, pi3696, pi3697,
    pi3698, pi3699, pi3700, pi3701, pi3702, pi3703, pi3704, pi3705, pi3706,
    pi3707, pi3708, pi3709, pi3710, pi3711, pi3712, pi3713, pi3714, pi3715,
    pi3716, pi3717, pi3718, pi3719, pi3720, pi3721, pi3722, pi3723, pi3724,
    pi3725, pi3726, pi3727, pi3728, pi3729, pi3730, pi3731, pi3732, pi3733,
    pi3734, pi3735, pi3736, pi3737, pi3738, pi3739, pi3740, pi3741, pi3742,
    pi3743, pi3744, pi3745, pi3746, pi3747, pi3748, pi3749, pi3750, pi3751,
    pi3752, pi3753, pi3754, pi3755, pi3756, pi3757, pi3758, pi3759, pi3760,
    pi3761, pi3762, pi3763, pi3764, pi3765, pi3766, pi3767, pi3768, pi3769,
    pi3770, pi3771, pi3772, pi3773, pi3774, pi3775, pi3776, pi3777, pi3778,
    pi3779, pi3780, pi3781, pi3782, pi3783, pi3784, pi3785, pi3786, pi3787,
    pi3788, pi3789, pi3790, pi3791, pi3792, pi3793, pi3794, pi3795, pi3796,
    pi3797, pi3798, pi3799, pi3800, pi3801, pi3802, pi3803, pi3804, pi3805,
    pi3806, pi3807, pi3808, pi3809, pi3810, pi3811, pi3812, pi3813, pi3814,
    pi3815, pi3816, pi3817, pi3818, pi3819, pi3820, pi3821, pi3822, pi3823,
    pi3824, pi3825, pi3826, pi3827, pi3828, pi3829, pi3830, pi3831, pi3832,
    pi3833, pi3834, pi3835, pi3836, pi3837, pi3838, pi3839, pi3840, pi3841,
    pi3842, pi3843, pi3844, pi3845, pi3846, pi3847, pi3848, pi3849, pi3850,
    pi3851, pi3852, pi3853, pi3854, pi3855, pi3856, pi3857, pi3858, pi3859,
    pi3860, pi3861, pi3862, pi3863, pi3864, pi3865, pi3866, pi3867, pi3868,
    pi3869, pi3870, pi3871, pi3872, pi3873, pi3874, pi3875, pi3876, pi3877,
    pi3878, pi3879, pi3880, pi3881, pi3882, pi3883, pi3884, pi3885, pi3886,
    pi3887, pi3888, pi3889, pi3890, pi3891, pi3892, pi3893, pi3894, pi3895,
    pi3896, pi3897, pi3898, pi3899, pi3900, pi3901, pi3902, pi3903, pi3904,
    pi3905, pi3906, pi3907, pi3908, pi3909, pi3910, pi3911, pi3912, pi3913,
    pi3914, pi3915, pi3916, pi3917, pi3918, pi3919, pi3920, pi3921, pi3922,
    pi3923, pi3924, pi3925, pi3926, pi3927, pi3928, pi3929, pi3930, pi3931,
    pi3932, pi3933, pi3934, pi3935, pi3936, pi3937, pi3938, pi3939, pi3940,
    pi3941, pi3942, pi3943, pi3944, pi3945, pi3946, pi3947, pi3948, pi3949,
    pi3950, pi3951, pi3952, pi3953, pi3954, pi3955, pi3956, pi3957, pi3958,
    pi3959, pi3960, pi3961, pi3962, pi3963, pi3964, pi3965, pi3966, pi3967,
    pi3968, pi3969, pi3970, pi3971, pi3972, pi3973, pi3974, pi3975, pi3976,
    pi3977, pi3978, pi3979, pi3980, pi3981, pi3982, pi3983, pi3984, pi3985,
    pi3986, pi3987, pi3988, pi3989, pi3990, pi3991, pi3992, pi3993, pi3994,
    pi3995, pi3996, pi3997, pi3998, pi3999, pi4000, pi4001, pi4002, pi4003,
    pi4004, pi4005, pi4006, pi4007, pi4008, pi4009, pi4010, pi4011, pi4012,
    pi4013, pi4014, pi4015, pi4016, pi4017, pi4018, pi4019, pi4020, pi4021,
    pi4022, pi4023, pi4024, pi4025, pi4026, pi4027, pi4028, pi4029, pi4030,
    pi4031, pi4032, pi4033, pi4034, pi4035, pi4036, pi4037, pi4038, pi4039,
    pi4040, pi4041, pi4042, pi4043, pi4044, pi4045, pi4046, pi4047, pi4048,
    pi4049, pi4050, pi4051, pi4052, pi4053, pi4054, pi4055, pi4056, pi4057,
    pi4058, pi4059, pi4060, pi4061, pi4062, pi4063, pi4064, pi4065, pi4066,
    pi4067, pi4068, pi4069, pi4070, pi4071, pi4072, pi4073, pi4074, pi4075,
    pi4076, pi4077, pi4078, pi4079, pi4080, pi4081, pi4082, pi4083, pi4084,
    pi4085, pi4086, pi4087, pi4088, pi4089, pi4090, pi4091, pi4092, pi4093,
    pi4094, pi4095, pi4096, pi4097, pi4098, pi4099, pi4100, pi4101, pi4102,
    pi4103, pi4104, pi4105, pi4106, pi4107, pi4108, pi4109, pi4110, pi4111,
    pi4112, pi4113, pi4114, pi4115, pi4116, pi4117, pi4118, pi4119, pi4120,
    pi4121, pi4122, pi4123, pi4124, pi4125, pi4126, pi4127, pi4128, pi4129,
    pi4130, pi4131, pi4132, pi4133, pi4134, pi4135, pi4136, pi4137, pi4138,
    pi4139, pi4140, pi4141, pi4142, pi4143, pi4144, pi4145, pi4146, pi4147,
    pi4148, pi4149, pi4150, pi4151, pi4152, pi4153, pi4154, pi4155, pi4156,
    pi4157, pi4158, pi4159, pi4160, pi4161, pi4162, pi4163, pi4164, pi4165,
    pi4166, pi4167, pi4168, pi4169, pi4170, pi4171, pi4172, pi4173, pi4174,
    pi4175, pi4176, pi4177, pi4178, pi4179, pi4180, pi4181, pi4182, pi4183,
    pi4184, pi4185, pi4186, pi4187, pi4188, pi4189, pi4190, pi4191, pi4192,
    pi4193, pi4194, pi4195, pi4196, pi4197, pi4198, pi4199, pi4200, pi4201,
    pi4202, pi4203, pi4204, pi4205, pi4206, pi4207, pi4208, pi4209, pi4210,
    pi4211, pi4212, pi4213, pi4214, pi4215, pi4216, pi4217, pi4218, pi4219,
    pi4220, pi4221, pi4222, pi4223, pi4224, pi4225, pi4226, pi4227, pi4228,
    pi4229, pi4230, pi4231, pi4232, pi4233, pi4234, pi4235, pi4236, pi4237,
    pi4238, pi4239, pi4240, pi4241, pi4242, pi4243, pi4244, pi4245, pi4246,
    pi4247, pi4248, pi4249, pi4250, pi4251, pi4252, pi4253, pi4254, pi4255,
    pi4256, pi4257, pi4258, pi4259, pi4260, pi4261, pi4262, pi4263, pi4264,
    pi4265, pi4266, pi4267, pi4268, pi4269, pi4270, pi4271, pi4272, pi4273,
    pi4274, pi4275, pi4276, pi4277, pi4278, pi4279, pi4280, pi4281, pi4282,
    pi4283, pi4284, pi4285, pi4286, pi4287, pi4288, pi4289, pi4290, pi4291,
    pi4292, pi4293, pi4294, pi4295, pi4296, pi4297, pi4298, pi4299, pi4300,
    pi4301, pi4302, pi4303, pi4304, pi4305, pi4306, pi4307, pi4308, pi4309,
    pi4310, pi4311, pi4312, pi4313, pi4314, pi4315, pi4316, pi4317, pi4318,
    pi4319, pi4320, pi4321, pi4322, pi4323, pi4324, pi4325, pi4326, pi4327,
    pi4328, pi4329, pi4330, pi4331, pi4332, pi4333, pi4334, pi4335, pi4336,
    pi4337, pi4338, pi4339, pi4340, pi4341, pi4342, pi4343, pi4344, pi4345,
    pi4346, pi4347, pi4348, pi4349, pi4350, pi4351, pi4352, pi4353, pi4354,
    pi4355, pi4356, pi4357, pi4358, pi4359, pi4360, pi4361, pi4362, pi4363,
    pi4364, pi4365, pi4366, pi4367, pi4368, pi4369, pi4370, pi4371, pi4372,
    pi4373, pi4374, pi4375, pi4376, pi4377, pi4378, pi4379, pi4380, pi4381,
    pi4382, pi4383, pi4384, pi4385, pi4386, pi4387, pi4388, pi4389, pi4390,
    pi4391, pi4392, pi4393, pi4394, pi4395, pi4396, pi4397, pi4398, pi4399,
    pi4400, pi4401, pi4402, pi4403, pi4404, pi4405, pi4406, pi4407, pi4408,
    pi4409, pi4410, pi4411, pi4412, pi4413, pi4414, pi4415, pi4416, pi4417,
    pi4418, pi4419, pi4420, pi4421, pi4422, pi4423, pi4424, pi4425, pi4426,
    pi4427, pi4428, pi4429, pi4430, pi4431, pi4432, pi4433, pi4434, pi4435,
    pi4436, pi4437, pi4438, pi4439, pi4440, pi4441, pi4442, pi4443, pi4444,
    pi4445, pi4446, pi4447, pi4448, pi4449, pi4450, pi4451, pi4452, pi4453,
    pi4454, pi4455, pi4456, pi4457, pi4458, pi4459, pi4460, pi4461, pi4462,
    pi4463, pi4464, pi4465, pi4466, pi4467, pi4468, pi4469, pi4470, pi4471,
    pi4472, pi4473, pi4474, pi4475, pi4476, pi4477, pi4478, pi4479, pi4480,
    pi4481, pi4482, pi4483, pi4484, pi4485, pi4486, pi4487, pi4488, pi4489,
    pi4490, pi4491, pi4492, pi4493, pi4494, pi4495, pi4496, pi4497, pi4498,
    pi4499, pi4500, pi4501, pi4502, pi4503, pi4504, pi4505, pi4506, pi4507,
    pi4508, pi4509, pi4510, pi4511, pi4512, pi4513, pi4514, pi4515, pi4516,
    pi4517, pi4518, pi4519, pi4520, pi4521, pi4522, pi4523, pi4524, pi4525,
    pi4526, pi4527, pi4528, pi4529, pi4530, pi4531, pi4532, pi4533, pi4534,
    pi4535, pi4536, pi4537, pi4538, pi4539, pi4540, pi4541, pi4542, pi4543,
    pi4544, pi4545, pi4546, pi4547, pi4548, pi4549, pi4550, pi4551, pi4552,
    pi4553, pi4554, pi4555, pi4556, pi4557, pi4558, pi4559, pi4560, pi4561,
    pi4562, pi4563, pi4564, pi4565, pi4566, pi4567, pi4568, pi4569, pi4570,
    pi4571, pi4572, pi4573, pi4574, pi4575, pi4576, pi4577, pi4578, pi4579,
    pi4580, pi4581, pi4582, pi4583, pi4584, pi4585, pi4586, pi4587, pi4588,
    pi4589, pi4590, pi4591, pi4592, pi4593, pi4594, pi4595, pi4596, pi4597,
    pi4598, pi4599, pi4600, pi4601, pi4602, pi4603, pi4604, pi4605, pi4606,
    pi4607, pi4608, pi4609, pi4610, pi4611, pi4612, pi4613, pi4614, pi4615,
    pi4616, pi4617, pi4618, pi4619, pi4620, pi4621, pi4622, pi4623, pi4624,
    pi4625, pi4626, pi4627, pi4628, pi4629, pi4630, pi4631, pi4632, pi4633,
    pi4634, pi4635, pi4636, pi4637, pi4638, pi4639, pi4640, pi4641, pi4642,
    pi4643, pi4644, pi4645, pi4646, pi4647, pi4648, pi4649, pi4650, pi4651,
    pi4652, pi4653, pi4654, pi4655, pi4656, pi4657, pi4658, pi4659, pi4660,
    pi4661, pi4662, pi4663, pi4664, pi4665, pi4666, pi4667, pi4668, pi4669,
    pi4670, pi4671, pi4672, pi4673, pi4674, pi4675, pi4676, pi4677, pi4678,
    pi4679, pi4680, pi4681, pi4682, pi4683, pi4684, pi4685, pi4686, pi4687,
    pi4688, pi4689, pi4690, pi4691, pi4692, pi4693, pi4694, pi4695, pi4696,
    pi4697, pi4698, pi4699, pi4700, pi4701, pi4702, pi4703, pi4704, pi4705,
    pi4706, pi4707, pi4708, pi4709, pi4710, pi4711, pi4712, pi4713, pi4714,
    pi4715, pi4716, pi4717, pi4718, pi4719, pi4720, pi4721, pi4722, pi4723,
    pi4724, pi4725, pi4726, pi4727, pi4728, pi4729, pi4730, pi4731, pi4732,
    pi4733, pi4734, pi4735, pi4736, pi4737, pi4738, pi4739, pi4740, pi4741,
    pi4742, pi4743, pi4744, pi4745, pi4746, pi4747, pi4748, pi4749, pi4750,
    pi4751, pi4752, pi4753, pi4754, pi4755, pi4756, pi4757, pi4758, pi4759,
    pi4760, pi4761, pi4762, pi4763, pi4764, pi4765, pi4766, pi4767, pi4768,
    pi4769, pi4770, pi4771, pi4772, pi4773, pi4774, pi4775, pi4776, pi4777,
    pi4778, pi4779, pi4780, pi4781, pi4782, pi4783, pi4784, pi4785, pi4786,
    pi4787, pi4788, pi4789, pi4790, pi4791, pi4792, pi4793, pi4794, pi4795,
    pi4796, pi4797, pi4798, pi4799, pi4800, pi4801, pi4802, pi4803, pi4804,
    pi4805, pi4806, pi4807, pi4808, pi4809, pi4810, pi4811, pi4812, pi4813,
    pi4814, pi4815, pi4816, pi4817, pi4818, pi4819, pi4820, pi4821, pi4822,
    pi4823, pi4824, pi4825, pi4826, pi4827, pi4828, pi4829, pi4830, pi4831,
    pi4832, pi4833, pi4834, pi4835, pi4836, pi4837, pi4838, pi4839, pi4840,
    pi4841, pi4842, pi4843, pi4844, pi4845, pi4846, pi4847, pi4848, pi4849,
    pi4850, pi4851, pi4852, pi4853, pi4854, pi4855, pi4856, pi4857, pi4858,
    pi4859, pi4860, pi4861, pi4862, pi4863, pi4864, pi4865, pi4866, pi4867,
    pi4868, pi4869, pi4870, pi4871, pi4872, pi4873, pi4874, pi4875, pi4876,
    pi4877, pi4878, pi4879, pi4880, pi4881, pi4882, pi4883, pi4884, pi4885,
    pi4886, pi4887, pi4888, pi4889, pi4890, pi4891, pi4892, pi4893, pi4894,
    pi4895, pi4896, pi4897, pi4898, pi4899, pi4900, pi4901, pi4902, pi4903,
    pi4904, pi4905, pi4906, pi4907, pi4908, pi4909, pi4910, pi4911, pi4912,
    pi4913, pi4914, pi4915, pi4916, pi4917, pi4918, pi4919, pi4920, pi4921,
    pi4922, pi4923, pi4924, pi4925, pi4926, pi4927, pi4928, pi4929, pi4930,
    pi4931, pi4932, pi4933, pi4934, pi4935, pi4936, pi4937, pi4938, pi4939,
    pi4940, pi4941, pi4942, pi4943, pi4944, pi4945, pi4946, pi4947, pi4948,
    pi4949, pi4950, pi4951, pi4952, pi4953, pi4954, pi4955, pi4956, pi4957,
    pi4958, pi4959, pi4960, pi4961, pi4962, pi4963, pi4964, pi4965, pi4966,
    pi4967, pi4968, pi4969, pi4970, pi4971, pi4972, pi4973, pi4974, pi4975,
    pi4976, pi4977, pi4978, pi4979, pi4980, pi4981, pi4982, pi4983, pi4984,
    pi4985, pi4986, pi4987, pi4988, pi4989, pi4990, pi4991, pi4992, pi4993,
    pi4994, pi4995, pi4996, pi4997, pi4998, pi4999, pi5000, pi5001, pi5002,
    pi5003, pi5004, pi5005, pi5006, pi5007, pi5008, pi5009, pi5010, pi5011,
    pi5012, pi5013, pi5014, pi5015, pi5016, pi5017, pi5018, pi5019, pi5020,
    pi5021, pi5022, pi5023, pi5024, pi5025, pi5026, pi5027, pi5028, pi5029,
    pi5030, pi5031, pi5032, pi5033, pi5034, pi5035, pi5036, pi5037, pi5038,
    pi5039, pi5040, pi5041, pi5042, pi5043, pi5044, pi5045, pi5046, pi5047,
    pi5048, pi5049, pi5050, pi5051, pi5052, pi5053, pi5054, pi5055, pi5056,
    pi5057, pi5058, pi5059, pi5060, pi5061, pi5062, pi5063, pi5064, pi5065,
    pi5066, pi5067, pi5068, pi5069, pi5070, pi5071, pi5072, pi5073, pi5074,
    pi5075, pi5076, pi5077, pi5078, pi5079, pi5080, pi5081, pi5082, pi5083,
    pi5084, pi5085, pi5086, pi5087, pi5088, pi5089, pi5090, pi5091, pi5092,
    pi5093, pi5094, pi5095, pi5096, pi5097, pi5098, pi5099, pi5100, pi5101,
    pi5102, pi5103, pi5104, pi5105, pi5106, pi5107, pi5108, pi5109, pi5110,
    pi5111, pi5112, pi5113, pi5114, pi5115, pi5116, pi5117, pi5118, pi5119,
    pi5120, pi5121, pi5122, pi5123, pi5124, pi5125, pi5126, pi5127, pi5128,
    pi5129, pi5130, pi5131, pi5132, pi5133, pi5134, pi5135, pi5136, pi5137,
    pi5138, pi5139, pi5140, pi5141, pi5142, pi5143, pi5144, pi5145, pi5146,
    pi5147, pi5148, pi5149, pi5150, pi5151, pi5152, pi5153, pi5154, pi5155,
    pi5156, pi5157, pi5158, pi5159, pi5160, pi5161, pi5162, pi5163, pi5164,
    pi5165, pi5166, pi5167, pi5168, pi5169, pi5170, pi5171, pi5172, pi5173,
    pi5174, pi5175, pi5176, pi5177, pi5178, pi5179, pi5180, pi5181, pi5182,
    pi5183, pi5184, pi5185, pi5186, pi5187, pi5188, pi5189, pi5190, pi5191,
    pi5192, pi5193, pi5194, pi5195, pi5196, pi5197, pi5198, pi5199, pi5200,
    pi5201, pi5202, pi5203, pi5204, pi5205, pi5206, pi5207, pi5208, pi5209,
    pi5210, pi5211, pi5212, pi5213, pi5214, pi5215, pi5216, pi5217, pi5218,
    pi5219, pi5220, pi5221, pi5222, pi5223, pi5224, pi5225, pi5226, pi5227,
    pi5228, pi5229, pi5230, pi5231, pi5232, pi5233, pi5234, pi5235, pi5236,
    pi5237, pi5238, pi5239, pi5240, pi5241, pi5242, pi5243, pi5244, pi5245,
    pi5246, pi5247, pi5248, pi5249, pi5250, pi5251, pi5252, pi5253, pi5254,
    pi5255, pi5256, pi5257, pi5258, pi5259, pi5260, pi5261, pi5262, pi5263,
    pi5264, pi5265, pi5266, pi5267, pi5268, pi5269, pi5270, pi5271, pi5272,
    pi5273, pi5274, pi5275, pi5276, pi5277, pi5278, pi5279, pi5280, pi5281,
    pi5282, pi5283, pi5284, pi5285, pi5286, pi5287, pi5288, pi5289, pi5290,
    pi5291, pi5292, pi5293, pi5294, pi5295, pi5296, pi5297, pi5298, pi5299,
    pi5300, pi5301, pi5302, pi5303, pi5304, pi5305, pi5306, pi5307, pi5308,
    pi5309, pi5310, pi5311, pi5312, pi5313, pi5314, pi5315, pi5316, pi5317,
    pi5318, pi5319, pi5320, pi5321, pi5322, pi5323, pi5324, pi5325, pi5326,
    pi5327, pi5328, pi5329, pi5330, pi5331, pi5332, pi5333, pi5334, pi5335,
    pi5336, pi5337, pi5338, pi5339, pi5340, pi5341, pi5342, pi5343, pi5344,
    pi5345, pi5346, pi5347, pi5348, pi5349, pi5350, pi5351, pi5352, pi5353,
    pi5354, pi5355, pi5356, pi5357, pi5358, pi5359, pi5360, pi5361, pi5362,
    pi5363, pi5364, pi5365, pi5366, pi5367, pi5368, pi5369, pi5370, pi5371,
    pi5372, pi5373, pi5374, pi5375, pi5376, pi5377, pi5378, pi5379, pi5380,
    pi5381, pi5382, pi5383, pi5384, pi5385, pi5386, pi5387, pi5388, pi5389,
    pi5390, pi5391, pi5392, pi5393, pi5394, pi5395, pi5396, pi5397, pi5398,
    pi5399, pi5400, pi5401, pi5402, pi5403, pi5404, pi5405, pi5406, pi5407,
    pi5408, pi5409, pi5410, pi5411, pi5412, pi5413, pi5414, pi5415, pi5416,
    pi5417, pi5418, pi5419, pi5420, pi5421, pi5422, pi5423, pi5424, pi5425,
    pi5426, pi5427, pi5428, pi5429, pi5430, pi5431, pi5432, pi5433, pi5434,
    pi5435, pi5436, pi5437, pi5438, pi5439, pi5440, pi5441, pi5442, pi5443,
    pi5444, pi5445, pi5446, pi5447, pi5448, pi5449, pi5450, pi5451, pi5452,
    pi5453, pi5454, pi5455, pi5456, pi5457, pi5458, pi5459, pi5460, pi5461,
    pi5462, pi5463, pi5464, pi5465, pi5466, pi5467, pi5468, pi5469, pi5470,
    pi5471, pi5472, pi5473, pi5474, pi5475, pi5476, pi5477, pi5478, pi5479,
    pi5480, pi5481, pi5482, pi5483, pi5484, pi5485, pi5486, pi5487, pi5488,
    pi5489, pi5490, pi5491, pi5492, pi5493, pi5494, pi5495, pi5496, pi5497,
    pi5498, pi5499, pi5500, pi5501, pi5502, pi5503, pi5504, pi5505, pi5506,
    pi5507, pi5508, pi5509, pi5510, pi5511, pi5512, pi5513, pi5514, pi5515,
    pi5516, pi5517, pi5518, pi5519, pi5520, pi5521, pi5522, pi5523, pi5524,
    pi5525, pi5526, pi5527, pi5528, pi5529, pi5530, pi5531, pi5532, pi5533,
    pi5534, pi5535, pi5536, pi5537, pi5538, pi5539, pi5540, pi5541, pi5542,
    pi5543, pi5544, pi5545, pi5546, pi5547, pi5548, pi5549, pi5550, pi5551,
    pi5552, pi5553, pi5554, pi5555, pi5556, pi5557, pi5558, pi5559, pi5560,
    pi5561, pi5562, pi5563, pi5564, pi5565, pi5566, pi5567, pi5568, pi5569,
    pi5570, pi5571, pi5572, pi5573, pi5574, pi5575, pi5576, pi5577, pi5578,
    pi5579, pi5580, pi5581, pi5582, pi5583, pi5584, pi5585, pi5586, pi5587,
    pi5588, pi5589, pi5590, pi5591, pi5592, pi5593, pi5594, pi5595, pi5596,
    pi5597, pi5598, pi5599, pi5600, pi5601, pi5602, pi5603, pi5604, pi5605,
    pi5606, pi5607, pi5608, pi5609, pi5610, pi5611, pi5612, pi5613, pi5614,
    pi5615, pi5616, pi5617, pi5618, pi5619, pi5620, pi5621, pi5622, pi5623,
    pi5624, pi5625, pi5626, pi5627, pi5628, pi5629, pi5630, pi5631, pi5632,
    pi5633, pi5634, pi5635, pi5636, pi5637, pi5638, pi5639, pi5640, pi5641,
    pi5642, pi5643, pi5644, pi5645, pi5646, pi5647, pi5648, pi5649, pi5650,
    pi5651, pi5652, pi5653, pi5654, pi5655, pi5656, pi5657, pi5658, pi5659,
    pi5660, pi5661, pi5662, pi5663, pi5664, pi5665, pi5666, pi5667, pi5668,
    pi5669, pi5670, pi5671, pi5672, pi5673, pi5674, pi5675, pi5676, pi5677,
    pi5678, pi5679, pi5680, pi5681, pi5682, pi5683, pi5684, pi5685, pi5686,
    pi5687, pi5688, pi5689, pi5690, pi5691, pi5692, pi5693, pi5694, pi5695,
    pi5696, pi5697, pi5698, pi5699, pi5700, pi5701, pi5702, pi5703, pi5704,
    pi5705, pi5706, pi5707, pi5708, pi5709, pi5710, pi5711, pi5712, pi5713,
    pi5714, pi5715, pi5716, pi5717, pi5718, pi5719, pi5720, pi5721, pi5722,
    pi5723, pi5724, pi5725, pi5726, pi5727, pi5728, pi5729, pi5730, pi5731,
    pi5732, pi5733, pi5734, pi5735, pi5736, pi5737, pi5738, pi5739, pi5740,
    pi5741, pi5742, pi5743, pi5744, pi5745, pi5746, pi5747, pi5748, pi5749,
    pi5750, pi5751, pi5752, pi5753, pi5754, pi5755, pi5756, pi5757, pi5758,
    pi5759, pi5760, pi5761, pi5762, pi5763, pi5764, pi5765, pi5766, pi5767,
    pi5768, pi5769, pi5770, pi5771, pi5772, pi5773, pi5774, pi5775, pi5776,
    pi5777, pi5778, pi5779, pi5780, pi5781, pi5782, pi5783, pi5784, pi5785,
    pi5786, pi5787, pi5788, pi5789, pi5790, pi5791, pi5792, pi5793, pi5794,
    pi5795, pi5796, pi5797, pi5798, pi5799, pi5800, pi5801, pi5802, pi5803,
    pi5804, pi5805, pi5806, pi5807, pi5808, pi5809, pi5810, pi5811, pi5812,
    pi5813, pi5814, pi5815, pi5816, pi5817, pi5818, pi5819, pi5820, pi5821,
    pi5822, pi5823, pi5824, pi5825, pi5826, pi5827, pi5828, pi5829, pi5830,
    pi5831, pi5832, pi5833, pi5834, pi5835, pi5836, pi5837, pi5838, pi5839,
    pi5840, pi5841, pi5842, pi5843, pi5844, pi5845, pi5846, pi5847, pi5848,
    pi5849, pi5850, pi5851, pi5852, pi5853, pi5854, pi5855, pi5856, pi5857,
    pi5858, pi5859, pi5860, pi5861, pi5862, pi5863, pi5864, pi5865, pi5866,
    pi5867, pi5868, pi5869, pi5870, pi5871, pi5872, pi5873, pi5874, pi5875,
    pi5876, pi5877, pi5878, pi5879, pi5880, pi5881, pi5882, pi5883, pi5884,
    pi5885, pi5886, pi5887, pi5888, pi5889, pi5890, pi5891, pi5892, pi5893,
    pi5894, pi5895, pi5896, pi5897, pi5898, pi5899, pi5900, pi5901, pi5902,
    pi5903, pi5904, pi5905, pi5906, pi5907, pi5908, pi5909, pi5910, pi5911,
    pi5912, pi5913, pi5914, pi5915, pi5916, pi5917, pi5918, pi5919, pi5920,
    pi5921, pi5922, pi5923, pi5924, pi5925, pi5926, pi5927, pi5928, pi5929,
    pi5930, pi5931, pi5932, pi5933, pi5934, pi5935, pi5936, pi5937, pi5938,
    pi5939, pi5940, pi5941, pi5942, pi5943, pi5944, pi5945, pi5946, pi5947,
    pi5948, pi5949, pi5950, pi5951, pi5952, pi5953, pi5954, pi5955, pi5956,
    pi5957, pi5958, pi5959, pi5960, pi5961, pi5962, pi5963, pi5964, pi5965,
    pi5966, pi5967, pi5968, pi5969, pi5970, pi5971, pi5972, pi5973, pi5974,
    pi5975, pi5976, pi5977, pi5978, pi5979, pi5980, pi5981, pi5982, pi5983,
    pi5984, pi5985, pi5986, pi5987, pi5988, pi5989, pi5990, pi5991, pi5992,
    pi5993, pi5994, pi5995, pi5996, pi5997, pi5998, pi5999, pi6000, pi6001,
    pi6002, pi6003, pi6004, pi6005, pi6006, pi6007, pi6008, pi6009, pi6010,
    pi6011, pi6012, pi6013, pi6014, pi6015, pi6016, pi6017, pi6018, pi6019,
    pi6020, pi6021, pi6022, pi6023, pi6024, pi6025, pi6026, pi6027, pi6028,
    pi6029, pi6030, pi6031, pi6032, pi6033, pi6034, pi6035, pi6036, pi6037,
    pi6038, pi6039, pi6040, pi6041, pi6042, pi6043, pi6044, pi6045, pi6046,
    pi6047, pi6048, pi6049, pi6050, pi6051, pi6052, pi6053, pi6054, pi6055,
    pi6056, pi6057, pi6058, pi6059, pi6060, pi6061, pi6062, pi6063, pi6064,
    pi6065, pi6066, pi6067, pi6068, pi6069, pi6070, pi6071, pi6072, pi6073,
    pi6074, pi6075, pi6076, pi6077, pi6078, pi6079, pi6080, pi6081, pi6082,
    pi6083, pi6084, pi6085, pi6086, pi6087, pi6088, pi6089, pi6090, pi6091,
    pi6092, pi6093, pi6094, pi6095, pi6096, pi6097, pi6098, pi6099, pi6100,
    pi6101, pi6102, pi6103, pi6104, pi6105, pi6106, pi6107, pi6108, pi6109,
    pi6110, pi6111, pi6112, pi6113, pi6114, pi6115, pi6116, pi6117, pi6118,
    pi6119, pi6120, pi6121, pi6122, pi6123, pi6124, pi6125, pi6126, pi6127,
    pi6128, pi6129, pi6130, pi6131, pi6132, pi6133, pi6134, pi6135, pi6136,
    pi6137, pi6138, pi6139, pi6140, pi6141, pi6142, pi6143, pi6144, pi6145,
    pi6146, pi6147, pi6148, pi6149, pi6150, pi6151, pi6152, pi6153, pi6154,
    pi6155, pi6156, pi6157, pi6158, pi6159, pi6160, pi6161, pi6162, pi6163,
    pi6164, pi6165, pi6166, pi6167, pi6168, pi6169, pi6170, pi6171, pi6172,
    pi6173, pi6174, pi6175, pi6176, pi6177, pi6178, pi6179, pi6180, pi6181,
    pi6182, pi6183, pi6184, pi6185, pi6186, pi6187, pi6188, pi6189, pi6190,
    pi6191, pi6192, pi6193, pi6194, pi6195, pi6196, pi6197, pi6198, pi6199,
    pi6200, pi6201, pi6202, pi6203, pi6204, pi6205, pi6206, pi6207, pi6208,
    pi6209, pi6210, pi6211, pi6212, pi6213, pi6214, pi6215, pi6216, pi6217,
    pi6218, pi6219, pi6220, pi6221, pi6222, pi6223, pi6224, pi6225, pi6226,
    pi6227, pi6228, pi6229, pi6230, pi6231, pi6232, pi6233, pi6234, pi6235,
    pi6236, pi6237, pi6238, pi6239, pi6240, pi6241, pi6242, pi6243, pi6244,
    pi6245, pi6246, pi6247, pi6248, pi6249, pi6250, pi6251, pi6252, pi6253,
    pi6254, pi6255, pi6256, pi6257, pi6258, pi6259, pi6260, pi6261, pi6262,
    pi6263, pi6264, pi6265, pi6266, pi6267, pi6268, pi6269, pi6270, pi6271,
    pi6272, pi6273, pi6274, pi6275, pi6276, pi6277, pi6278, pi6279, pi6280,
    pi6281, pi6282, pi6283, pi6284, pi6285, pi6286, pi6287, pi6288, pi6289,
    pi6290, pi6291, pi6292, pi6293, pi6294, pi6295, pi6296, pi6297, pi6298,
    pi6299, pi6300, pi6301, pi6302, pi6303, pi6304, pi6305, pi6306, pi6307,
    pi6308, pi6309, pi6310, pi6311, pi6312, pi6313, pi6314, pi6315, pi6316,
    pi6317, pi6318, pi6319, pi6320, pi6321, pi6322, pi6323, pi6324, pi6325,
    pi6326, pi6327, pi6328, pi6329, pi6330, pi6331, pi6332, pi6333, pi6334,
    pi6335, pi6336, pi6337, pi6338, pi6339, pi6340, pi6341, pi6342, pi6343,
    pi6344, pi6345, pi6346, pi6347, pi6348, pi6349, pi6350, pi6351, pi6352,
    pi6353, pi6354, pi6355, pi6356, pi6357, pi6358, pi6359, pi6360, pi6361,
    pi6362, pi6363, pi6364, pi6365, pi6366, pi6367, pi6368, pi6369, pi6370,
    pi6371, pi6372, pi6373, pi6374, pi6375, pi6376, pi6377, pi6378, pi6379,
    pi6380, pi6381, pi6382, pi6383, pi6384, pi6385, pi6386, pi6387, pi6388,
    pi6389, pi6390, pi6391, pi6392, pi6393, pi6394, pi6395, pi6396, pi6397,
    pi6398, pi6399, pi6400, pi6401, pi6402, pi6403, pi6404, pi6405, pi6406,
    pi6407, pi6408, pi6409, pi6410, pi6411, pi6412, pi6413, pi6414, pi6415,
    pi6416, pi6417, pi6418, pi6419, pi6420, pi6421, pi6422, pi6423, pi6424,
    pi6425, pi6426, pi6427, pi6428, pi6429, pi6430, pi6431, pi6432, pi6433,
    pi6434, pi6435, pi6436, pi6437, pi6438, pi6439, pi6440, pi6441, pi6442,
    pi6443, pi6444, pi6445, pi6446, pi6447, pi6448, pi6449, pi6450, pi6451,
    pi6452, pi6453, pi6454, pi6455, pi6456, pi6457, pi6458, pi6459, pi6460,
    pi6461, pi6462, pi6463, pi6464, pi6465, pi6466, pi6467, pi6468, pi6469,
    pi6470, pi6471, pi6472, pi6473, pi6474, pi6475, pi6476, pi6477, pi6478,
    pi6479, pi6480, pi6481, pi6482, pi6483, pi6484, pi6485, pi6486, pi6487,
    pi6488, pi6489, pi6490, pi6491, pi6492, pi6493, pi6494, pi6495, pi6496,
    pi6497, pi6498, pi6499, pi6500, pi6501, pi6502, pi6503, pi6504, pi6505,
    pi6506, pi6507, pi6508, pi6509, pi6510, pi6511, pi6512, pi6513, pi6514,
    pi6515, pi6516, pi6517, pi6518, pi6519, pi6520, pi6521, pi6522, pi6523,
    pi6524, pi6525, pi6526, pi6527, pi6528, pi6529, pi6530, pi6531, pi6532,
    pi6533, pi6534, pi6535, pi6536, pi6537, pi6538, pi6539, pi6540, pi6541,
    pi6542, pi6543, pi6544, pi6545, pi6546, pi6547, pi6548, pi6549, pi6550,
    pi6551, pi6552, pi6553, pi6554, pi6555, pi6556, pi6557, pi6558, pi6559,
    pi6560, pi6561, pi6562, pi6563, pi6564, pi6565, pi6566, pi6567, pi6568,
    pi6569, pi6570, pi6571, pi6572, pi6573, pi6574, pi6575, pi6576, pi6577,
    pi6578, pi6579, pi6580, pi6581, pi6582, pi6583, pi6584, pi6585, pi6586,
    pi6587, pi6588, pi6589, pi6590, pi6591, pi6592, pi6593, pi6594, pi6595,
    pi6596, pi6597, pi6598, pi6599, pi6600, pi6601, pi6602, pi6603, pi6604,
    pi6605, pi6606, pi6607, pi6608, pi6609, pi6610, pi6611, pi6612, pi6613,
    pi6614, pi6615, pi6616, pi6617, pi6618, pi6619, pi6620, pi6621, pi6622,
    pi6623, pi6624, pi6625, pi6626, pi6627, pi6628, pi6629, pi6630, pi6631,
    pi6632, pi6633, pi6634, pi6635, pi6636, pi6637, pi6638, pi6639, pi6640,
    pi6641, pi6642, pi6643, pi6644, pi6645, pi6646, pi6647, pi6648, pi6649,
    pi6650, pi6651, pi6652, pi6653, pi6654, pi6655, pi6656, pi6657, pi6658,
    pi6659, pi6660, pi6661, pi6662, pi6663, pi6664, pi6665, pi6666, pi6667,
    pi6668, pi6669, pi6670, pi6671, pi6672, pi6673, pi6674, pi6675, pi6676,
    pi6677, pi6678, pi6679, pi6680, pi6681, pi6682, pi6683, pi6684, pi6685,
    pi6686, pi6687, pi6688, pi6689, pi6690, pi6691, pi6692, pi6693, pi6694,
    pi6695, pi6696, pi6697, pi6698, pi6699, pi6700, pi6701, pi6702, pi6703,
    pi6704, pi6705, pi6706, pi6707, pi6708, pi6709, pi6710, pi6711, pi6712,
    pi6713, pi6714, pi6715, pi6716, pi6717, pi6718, pi6719, pi6720, pi6721,
    pi6722, pi6723, pi6724, pi6725, pi6726, pi6727, pi6728, pi6729, pi6730,
    pi6731, pi6732, pi6733, pi6734, pi6735, pi6736, pi6737, pi6738, pi6739,
    pi6740, pi6741, pi6742, pi6743, pi6744, pi6745, pi6746, pi6747, pi6748,
    pi6749, pi6750, pi6751, pi6752, pi6753, pi6754, pi6755, pi6756, pi6757,
    pi6758, pi6759, pi6760, pi6761, pi6762, pi6763, pi6764, pi6765, pi6766,
    pi6767, pi6768, pi6769, pi6770, pi6771, pi6772, pi6773, pi6774, pi6775,
    pi6776, pi6777, pi6778, pi6779, pi6780, pi6781, pi6782, pi6783, pi6784,
    pi6785, pi6786, pi6787, pi6788, pi6789, pi6790, pi6791, pi6792, pi6793,
    pi6794, pi6795, pi6796, pi6797, pi6798, pi6799, pi6800, pi6801, pi6802,
    pi6803, pi6804, pi6805, pi6806, pi6807, pi6808, pi6809, pi6810, pi6811,
    pi6812, pi6813, pi6814, pi6815, pi6816, pi6817, pi6818, pi6819, pi6820,
    pi6821, pi6822, pi6823, pi6824, pi6825, pi6826, pi6827, pi6828, pi6829,
    pi6830, pi6831, pi6832, pi6833, pi6834, pi6835, pi6836, pi6837, pi6838,
    pi6839, pi6840, pi6841, pi6842, pi6843, pi6844, pi6845, pi6846, pi6847,
    pi6848, pi6849, pi6850, pi6851, pi6852, pi6853, pi6854, pi6855, pi6856,
    pi6857, pi6858, pi6859, pi6860, pi6861, pi6862, pi6863, pi6864, pi6865,
    pi6866, pi6867, pi6868, pi6869, pi6870, pi6871, pi6872, pi6873, pi6874,
    pi6875, pi6876, pi6877, pi6878, pi6879, pi6880, pi6881, pi6882, pi6883,
    pi6884, pi6885, pi6886, pi6887, pi6888, pi6889, pi6890, pi6891, pi6892,
    pi6893, pi6894, pi6895, pi6896, pi6897, pi6898, pi6899, pi6900, pi6901,
    pi6902, pi6903, pi6904, pi6905, pi6906, pi6907, pi6908, pi6909, pi6910,
    pi6911, pi6912, pi6913, pi6914, pi6915, pi6916, pi6917, pi6918, pi6919,
    pi6920, pi6921, pi6922, pi6923, pi6924, pi6925, pi6926, pi6927, pi6928,
    pi6929, pi6930, pi6931, pi6932, pi6933, pi6934, pi6935, pi6936, pi6937,
    pi6938, pi6939, pi6940, pi6941, pi6942, pi6943, pi6944, pi6945, pi6946,
    pi6947, pi6948, pi6949, pi6950, pi6951, pi6952, pi6953, pi6954, pi6955,
    pi6956, pi6957, pi6958, pi6959, pi6960, pi6961, pi6962, pi6963, pi6964,
    pi6965, pi6966, pi6967, pi6968, pi6969, pi6970, pi6971, pi6972, pi6973,
    pi6974, pi6975, pi6976, pi6977, pi6978, pi6979, pi6980, pi6981, pi6982,
    pi6983, pi6984, pi6985, pi6986, pi6987, pi6988, pi6989, pi6990, pi6991,
    pi6992, pi6993, pi6994, pi6995, pi6996, pi6997, pi6998, pi6999, pi7000,
    pi7001, pi7002, pi7003, pi7004, pi7005, pi7006, pi7007, pi7008, pi7009,
    pi7010, pi7011, pi7012, pi7013, pi7014, pi7015, pi7016, pi7017, pi7018,
    pi7019, pi7020, pi7021, pi7022, pi7023, pi7024, pi7025, pi7026, pi7027,
    pi7028, pi7029, pi7030, pi7031, pi7032, pi7033, pi7034, pi7035, pi7036,
    pi7037, pi7038, pi7039, pi7040, pi7041, pi7042, pi7043, pi7044, pi7045,
    pi7046, pi7047, pi7048, pi7049, pi7050, pi7051, pi7052, pi7053, pi7054,
    pi7055, pi7056, pi7057, pi7058, pi7059, pi7060, pi7061, pi7062, pi7063,
    pi7064, pi7065, pi7066, pi7067, pi7068, pi7069, pi7070, pi7071, pi7072,
    pi7073, pi7074, pi7075, pi7076, pi7077, pi7078, pi7079, pi7080, pi7081,
    pi7082, pi7083, pi7084, pi7085, pi7086, pi7087, pi7088, pi7089, pi7090,
    pi7091, pi7092, pi7093, pi7094, pi7095, pi7096, pi7097, pi7098, pi7099,
    pi7100, pi7101, pi7102, pi7103, pi7104, pi7105, pi7106, pi7107, pi7108,
    pi7109, pi7110, pi7111, pi7112, pi7113, pi7114, pi7115, pi7116, pi7117,
    pi7118, pi7119, pi7120, pi7121, pi7122, pi7123, pi7124, pi7125, pi7126,
    pi7127, pi7128, pi7129, pi7130, pi7131, pi7132, pi7133, pi7134, pi7135,
    pi7136, pi7137, pi7138, pi7139, pi7140, pi7141, pi7142, pi7143, pi7144,
    pi7145, pi7146, pi7147, pi7148, pi7149, pi7150, pi7151, pi7152, pi7153,
    pi7154, pi7155, pi7156, pi7157, pi7158, pi7159, pi7160, pi7161, pi7162,
    pi7163, pi7164, pi7165, pi7166, pi7167, pi7168, pi7169, pi7170, pi7171,
    pi7172, pi7173, pi7174, pi7175, pi7176, pi7177, pi7178, pi7179, pi7180,
    pi7181, pi7182, pi7183, pi7184, pi7185, pi7186, pi7187, pi7188, pi7189,
    pi7190, pi7191, pi7192, pi7193, pi7194, pi7195, pi7196, pi7197, pi7198,
    pi7199, pi7200, pi7201, pi7202, pi7203, pi7204, pi7205, pi7206, pi7207,
    pi7208, pi7209, pi7210, pi7211, pi7212, pi7213, pi7214, pi7215, pi7216,
    pi7217, pi7218, pi7219, pi7220, pi7221, pi7222, pi7223, pi7224, pi7225,
    pi7226, pi7227, pi7228, pi7229, pi7230, pi7231, pi7232, pi7233, pi7234,
    pi7235, pi7236, pi7237, pi7238, pi7239, pi7240, pi7241, pi7242, pi7243,
    pi7244, pi7245, pi7246, pi7247, pi7248, pi7249, pi7250, pi7251, pi7252,
    pi7253, pi7254, pi7255, pi7256, pi7257, pi7258, pi7259, pi7260, pi7261,
    pi7262, pi7263, pi7264, pi7265, pi7266, pi7267, pi7268, pi7269, pi7270,
    pi7271, pi7272, pi7273, pi7274, pi7275, pi7276, pi7277, pi7278, pi7279,
    pi7280, pi7281, pi7282, pi7283, pi7284, pi7285, pi7286, pi7287, pi7288,
    pi7289, pi7290, pi7291, pi7292, pi7293, pi7294, pi7295, pi7296, pi7297,
    pi7298, pi7299, pi7300, pi7301, pi7302, pi7303, pi7304, pi7305, pi7306,
    pi7307, pi7308, pi7309, pi7310, pi7311, pi7312, pi7313, pi7314, pi7315,
    pi7316, pi7317, pi7318, pi7319, pi7320, pi7321, pi7322, pi7323, pi7324,
    pi7325, pi7326, pi7327, pi7328, pi7329, pi7330, pi7331, pi7332, pi7333,
    pi7334, pi7335, pi7336, pi7337, pi7338, pi7339, pi7340, pi7341, pi7342,
    pi7343, pi7344, pi7345, pi7346, pi7347, pi7348, pi7349, pi7350, pi7351,
    pi7352, pi7353, pi7354, pi7355, pi7356, pi7357, pi7358, pi7359, pi7360,
    pi7361, pi7362, pi7363, pi7364, pi7365, pi7366, pi7367, pi7368, pi7369,
    pi7370, pi7371, pi7372, pi7373, pi7374, pi7375, pi7376, pi7377, pi7378,
    pi7379, pi7380, pi7381, pi7382, pi7383, pi7384, pi7385, pi7386, pi7387,
    pi7388, pi7389, pi7390, pi7391, pi7392, pi7393, pi7394, pi7395, pi7396,
    pi7397, pi7398, pi7399, pi7400, pi7401, pi7402, pi7403, pi7404, pi7405,
    pi7406, pi7407, pi7408, pi7409, pi7410, pi7411, pi7412, pi7413, pi7414,
    pi7415, pi7416, pi7417, pi7418, pi7419, pi7420, pi7421, pi7422, pi7423,
    pi7424, pi7425, pi7426, pi7427, pi7428, pi7429, pi7430, pi7431, pi7432,
    pi7433, pi7434, pi7435, pi7436, pi7437, pi7438, pi7439, pi7440, pi7441,
    pi7442, pi7443, pi7444, pi7445, pi7446, pi7447, pi7448, pi7449, pi7450,
    pi7451, pi7452, pi7453, pi7454, pi7455, pi7456, pi7457, pi7458, pi7459,
    pi7460, pi7461, pi7462, pi7463, pi7464, pi7465, pi7466, pi7467, pi7468,
    pi7469, pi7470, pi7471, pi7472, pi7473, pi7474, pi7475, pi7476, pi7477,
    pi7478, pi7479, pi7480, pi7481, pi7482, pi7483, pi7484, pi7485, pi7486,
    pi7487, pi7488, pi7489, pi7490, pi7491, pi7492, pi7493, pi7494, pi7495,
    pi7496, pi7497, pi7498, pi7499, pi7500, pi7501, pi7502, pi7503, pi7504,
    pi7505, pi7506, pi7507, pi7508, pi7509, pi7510, pi7511, pi7512, pi7513,
    pi7514, pi7515, pi7516, pi7517, pi7518, pi7519, pi7520, pi7521, pi7522,
    pi7523, pi7524, pi7525, pi7526, pi7527, pi7528, pi7529, pi7530, pi7531,
    pi7532, pi7533, pi7534, pi7535, pi7536, pi7537, pi7538, pi7539, pi7540,
    pi7541, pi7542, pi7543, pi7544, pi7545, pi7546, pi7547, pi7548, pi7549,
    pi7550, pi7551, pi7552, pi7553, pi7554, pi7555, pi7556, pi7557, pi7558,
    pi7559, pi7560, pi7561, pi7562, pi7563, pi7564, pi7565, pi7566, pi7567,
    pi7568, pi7569, pi7570, pi7571, pi7572, pi7573, pi7574, pi7575, pi7576,
    pi7577, pi7578, pi7579, pi7580, pi7581, pi7582, pi7583, pi7584, pi7585,
    pi7586, pi7587, pi7588, pi7589, pi7590, pi7591, pi7592, pi7593, pi7594,
    pi7595, pi7596, pi7597, pi7598, pi7599, pi7600, pi7601, pi7602, pi7603,
    pi7604, pi7605, pi7606, pi7607, pi7608, pi7609, pi7610, pi7611, pi7612,
    pi7613, pi7614, pi7615, pi7616, pi7617, pi7618, pi7619, pi7620, pi7621,
    pi7622, pi7623, pi7624, pi7625, pi7626, pi7627, pi7628, pi7629, pi7630,
    pi7631, pi7632, pi7633, pi7634, pi7635, pi7636, pi7637, pi7638, pi7639,
    pi7640, pi7641, pi7642, pi7643, pi7644, pi7645, pi7646, pi7647, pi7648,
    pi7649, pi7650, pi7651, pi7652, pi7653, pi7654, pi7655, pi7656, pi7657,
    pi7658, pi7659, pi7660, pi7661, pi7662, pi7663, pi7664, pi7665, pi7666,
    pi7667, pi7668, pi7669, pi7670, pi7671, pi7672, pi7673, pi7674, pi7675,
    pi7676, pi7677, pi7678, pi7679, pi7680, pi7681, pi7682, pi7683, pi7684,
    pi7685, pi7686, pi7687, pi7688, pi7689, pi7690, pi7691, pi7692, pi7693,
    pi7694, pi7695, pi7696, pi7697, pi7698, pi7699, pi7700, pi7701, pi7702,
    pi7703, pi7704, pi7705, pi7706, pi7707, pi7708, pi7709, pi7710, pi7711,
    pi7712, pi7713, pi7714, pi7715, pi7716, pi7717, pi7718, pi7719, pi7720,
    pi7721, pi7722, pi7723, pi7724, pi7725, pi7726, pi7727, pi7728, pi7729,
    pi7730, pi7731, pi7732, pi7733, pi7734, pi7735, pi7736, pi7737, pi7738,
    pi7739, pi7740, pi7741, pi7742, pi7743, pi7744, pi7745, pi7746, pi7747,
    pi7748, pi7749, pi7750, pi7751, pi7752, pi7753, pi7754, pi7755, pi7756,
    pi7757, pi7758, pi7759, pi7760, pi7761, pi7762, pi7763, pi7764, pi7765,
    pi7766, pi7767, pi7768, pi7769, pi7770, pi7771, pi7772, pi7773, pi7774,
    pi7775, pi7776, pi7777, pi7778, pi7779, pi7780, pi7781, pi7782, pi7783,
    pi7784, pi7785, pi7786, pi7787, pi7788, pi7789, pi7790, pi7791, pi7792,
    pi7793, pi7794, pi7795, pi7796, pi7797, pi7798, pi7799, pi7800, pi7801,
    pi7802, pi7803, pi7804, pi7805, pi7806, pi7807, pi7808, pi7809, pi7810,
    pi7811, pi7812, pi7813, pi7814, pi7815, pi7816, pi7817, pi7818, pi7819,
    pi7820, pi7821, pi7822, pi7823, pi7824, pi7825, pi7826, pi7827, pi7828,
    pi7829, pi7830, pi7831, pi7832, pi7833, pi7834, pi7835, pi7836, pi7837,
    pi7838, pi7839, pi7840, pi7841, pi7842, pi7843, pi7844, pi7845, pi7846,
    pi7847, pi7848, pi7849, pi7850, pi7851, pi7852, pi7853, pi7854, pi7855,
    pi7856, pi7857, pi7858, pi7859, pi7860, pi7861, pi7862, pi7863, pi7864,
    pi7865, pi7866, pi7867, pi7868, pi7869, pi7870, pi7871, pi7872, pi7873,
    pi7874, pi7875, pi7876, pi7877, pi7878, pi7879, pi7880, pi7881, pi7882,
    pi7883, pi7884, pi7885, pi7886, pi7887, pi7888, pi7889, pi7890, pi7891,
    pi7892, pi7893, pi7894, pi7895, pi7896, pi7897, pi7898, pi7899, pi7900,
    pi7901, pi7902, pi7903, pi7904, pi7905, pi7906, pi7907, pi7908, pi7909,
    pi7910, pi7911, pi7912, pi7913, pi7914, pi7915, pi7916, pi7917, pi7918,
    pi7919, pi7920, pi7921, pi7922, pi7923, pi7924, pi7925, pi7926, pi7927,
    pi7928, pi7929, pi7930, pi7931, pi7932, pi7933, pi7934, pi7935, pi7936,
    pi7937, pi7938, pi7939, pi7940, pi7941, pi7942, pi7943, pi7944, pi7945,
    pi7946, pi7947, pi7948, pi7949, pi7950, pi7951, pi7952, pi7953, pi7954,
    pi7955, pi7956, pi7957, pi7958, pi7959, pi7960, pi7961, pi7962, pi7963,
    pi7964, pi7965, pi7966, pi7967, pi7968, pi7969, pi7970, pi7971, pi7972,
    pi7973, pi7974, pi7975, pi7976, pi7977, pi7978, pi7979, pi7980, pi7981,
    pi7982, pi7983, pi7984, pi7985, pi7986, pi7987, pi7988, pi7989, pi7990,
    pi7991, pi7992, pi7993, pi7994, pi7995, pi7996, pi7997, pi7998, pi7999,
    pi8000, pi8001, pi8002, pi8003, pi8004, pi8005, pi8006, pi8007, pi8008,
    pi8009, pi8010, pi8011, pi8012, pi8013, pi8014, pi8015, pi8016, pi8017,
    pi8018, pi8019, pi8020, pi8021, pi8022, pi8023, pi8024, pi8025, pi8026,
    pi8027, pi8028, pi8029, pi8030, pi8031, pi8032, pi8033, pi8034, pi8035,
    pi8036, pi8037, pi8038, pi8039, pi8040, pi8041, pi8042, pi8043, pi8044,
    pi8045, pi8046, pi8047, pi8048, pi8049, pi8050, pi8051, pi8052, pi8053,
    pi8054, pi8055, pi8056, pi8057, pi8058, pi8059, pi8060, pi8061, pi8062,
    pi8063, pi8064, pi8065, pi8066, pi8067, pi8068, pi8069, pi8070, pi8071,
    pi8072, pi8073, pi8074, pi8075, pi8076, pi8077, pi8078, pi8079, pi8080,
    pi8081, pi8082, pi8083, pi8084, pi8085, pi8086, pi8087, pi8088, pi8089,
    pi8090, pi8091, pi8092, pi8093, pi8094, pi8095, pi8096, pi8097, pi8098,
    pi8099, pi8100, pi8101, pi8102, pi8103, pi8104, pi8105, pi8106, pi8107,
    pi8108, pi8109, pi8110, pi8111, pi8112, pi8113, pi8114, pi8115, pi8116,
    pi8117, pi8118, pi8119, pi8120, pi8121, pi8122, pi8123, pi8124, pi8125,
    pi8126, pi8127, pi8128, pi8129, pi8130, pi8131, pi8132, pi8133, pi8134,
    pi8135, pi8136, pi8137, pi8138, pi8139, pi8140, pi8141, pi8142, pi8143,
    pi8144, pi8145, pi8146, pi8147, pi8148, pi8149, pi8150, pi8151, pi8152,
    pi8153, pi8154, pi8155, pi8156, pi8157, pi8158, pi8159, pi8160, pi8161,
    pi8162, pi8163, pi8164, pi8165, pi8166, pi8167, pi8168, pi8169, pi8170,
    pi8171, pi8172, pi8173, pi8174, pi8175, pi8176, pi8177, pi8178, pi8179,
    pi8180, pi8181, pi8182, pi8183, pi8184, pi8185, pi8186, pi8187, pi8188,
    pi8189, pi8190, pi8191, pi8192, pi8193, pi8194, pi8195, pi8196, pi8197,
    pi8198, pi8199, pi8200, pi8201, pi8202, pi8203, pi8204, pi8205, pi8206,
    pi8207, pi8208, pi8209, pi8210, pi8211, pi8212, pi8213, pi8214, pi8215,
    pi8216, pi8217, pi8218, pi8219, pi8220, pi8221, pi8222, pi8223, pi8224,
    pi8225, pi8226, pi8227, pi8228, pi8229, pi8230, pi8231, pi8232, pi8233,
    pi8234, pi8235, pi8236, pi8237, pi8238, pi8239, pi8240, pi8241, pi8242,
    pi8243, pi8244, pi8245, pi8246, pi8247, pi8248, pi8249, pi8250, pi8251,
    pi8252, pi8253, pi8254, pi8255, pi8256, pi8257, pi8258, pi8259, pi8260,
    pi8261, pi8262, pi8263, pi8264, pi8265, pi8266, pi8267, pi8268, pi8269,
    pi8270, pi8271, pi8272, pi8273, pi8274, pi8275, pi8276, pi8277, pi8278,
    pi8279, pi8280, pi8281, pi8282, pi8283, pi8284, pi8285, pi8286, pi8287,
    pi8288, pi8289, pi8290, pi8291, pi8292, pi8293, pi8294, pi8295, pi8296,
    pi8297, pi8298, pi8299, pi8300, pi8301, pi8302, pi8303, pi8304, pi8305,
    pi8306, pi8307, pi8308, pi8309, pi8310, pi8311, pi8312, pi8313, pi8314,
    pi8315, pi8316, pi8317, pi8318, pi8319, pi8320, pi8321, pi8322, pi8323,
    pi8324, pi8325, pi8326, pi8327, pi8328, pi8329, pi8330, pi8331, pi8332,
    pi8333, pi8334, pi8335, pi8336, pi8337, pi8338, pi8339, pi8340, pi8341,
    pi8342, pi8343, pi8344, pi8345, pi8346, pi8347, pi8348, pi8349, pi8350,
    pi8351, pi8352, pi8353, pi8354, pi8355, pi8356, pi8357, pi8358, pi8359,
    pi8360, pi8361, pi8362, pi8363, pi8364, pi8365, pi8366, pi8367, pi8368,
    pi8369, pi8370, pi8371, pi8372, pi8373, pi8374, pi8375, pi8376, pi8377,
    pi8378, pi8379, pi8380, pi8381, pi8382, pi8383, pi8384, pi8385, pi8386,
    pi8387, pi8388, pi8389, pi8390, pi8391, pi8392, pi8393, pi8394, pi8395,
    pi8396, pi8397, pi8398, pi8399, pi8400, pi8401, pi8402, pi8403, pi8404,
    pi8405, pi8406, pi8407, pi8408, pi8409, pi8410, pi8411, pi8412, pi8413,
    pi8414, pi8415, pi8416, pi8417, pi8418, pi8419, pi8420, pi8421, pi8422,
    pi8423, pi8424, pi8425, pi8426, pi8427, pi8428, pi8429, pi8430, pi8431,
    pi8432, pi8433, pi8434, pi8435, pi8436, pi8437, pi8438, pi8439, pi8440,
    pi8441, pi8442, pi8443, pi8444, pi8445, pi8446, pi8447, pi8448, pi8449,
    pi8450, pi8451, pi8452, pi8453, pi8454, pi8455, pi8456, pi8457, pi8458,
    pi8459, pi8460, pi8461, pi8462, pi8463, pi8464, pi8465, pi8466, pi8467,
    pi8468, pi8469, pi8470, pi8471, pi8472, pi8473, pi8474, pi8475, pi8476,
    pi8477, pi8478, pi8479, pi8480, pi8481, pi8482, pi8483, pi8484, pi8485,
    pi8486, pi8487, pi8488, pi8489, pi8490, pi8491, pi8492, pi8493, pi8494,
    pi8495, pi8496, pi8497, pi8498, pi8499, pi8500, pi8501, pi8502, pi8503,
    pi8504, pi8505, pi8506, pi8507, pi8508, pi8509, pi8510, pi8511, pi8512,
    pi8513, pi8514, pi8515, pi8516, pi8517, pi8518, pi8519, pi8520, pi8521,
    pi8522, pi8523, pi8524, pi8525, pi8526, pi8527, pi8528, pi8529, pi8530,
    pi8531, pi8532, pi8533, pi8534, pi8535, pi8536, pi8537, pi8538, pi8539,
    pi8540, pi8541, pi8542, pi8543, pi8544, pi8545, pi8546, pi8547, pi8548,
    pi8549, pi8550, pi8551, pi8552, pi8553, pi8554, pi8555, pi8556, pi8557,
    pi8558, pi8559, pi8560, pi8561, pi8562, pi8563, pi8564, pi8565, pi8566,
    pi8567, pi8568, pi8569, pi8570, pi8571, pi8572, pi8573, pi8574, pi8575,
    pi8576, pi8577, pi8578, pi8579, pi8580, pi8581, pi8582, pi8583, pi8584,
    pi8585, pi8586, pi8587, pi8588, pi8589, pi8590, pi8591, pi8592, pi8593,
    pi8594, pi8595, pi8596, pi8597, pi8598, pi8599, pi8600, pi8601, pi8602,
    pi8603, pi8604, pi8605, pi8606, pi8607, pi8608, pi8609, pi8610, pi8611,
    pi8612, pi8613, pi8614, pi8615, pi8616, pi8617, pi8618, pi8619, pi8620,
    pi8621, pi8622, pi8623, pi8624, pi8625, pi8626, pi8627, pi8628, pi8629,
    pi8630, pi8631, pi8632, pi8633, pi8634, pi8635, pi8636, pi8637, pi8638,
    pi8639, pi8640, pi8641, pi8642, pi8643, pi8644, pi8645, pi8646, pi8647,
    pi8648, pi8649, pi8650, pi8651, pi8652, pi8653, pi8654, pi8655, pi8656,
    pi8657, pi8658, pi8659, pi8660, pi8661, pi8662, pi8663, pi8664, pi8665,
    pi8666, pi8667, pi8668, pi8669, pi8670, pi8671, pi8672, pi8673, pi8674,
    pi8675, pi8676, pi8677, pi8678, pi8679, pi8680, pi8681, pi8682, pi8683,
    pi8684, pi8685, pi8686, pi8687, pi8688, pi8689, pi8690, pi8691, pi8692,
    pi8693, pi8694, pi8695, pi8696, pi8697, pi8698, pi8699, pi8700, pi8701,
    pi8702, pi8703, pi8704, pi8705, pi8706, pi8707, pi8708, pi8709, pi8710,
    pi8711, pi8712, pi8713, pi8714, pi8715, pi8716, pi8717, pi8718, pi8719,
    pi8720, pi8721, pi8722, pi8723, pi8724, pi8725, pi8726, pi8727, pi8728,
    pi8729, pi8730, pi8731, pi8732, pi8733, pi8734, pi8735, pi8736, pi8737,
    pi8738, pi8739, pi8740, pi8741, pi8742, pi8743, pi8744, pi8745, pi8746,
    pi8747, pi8748, pi8749, pi8750, pi8751, pi8752, pi8753, pi8754, pi8755,
    pi8756, pi8757, pi8758, pi8759, pi8760, pi8761, pi8762, pi8763, pi8764,
    pi8765, pi8766, pi8767, pi8768, pi8769, pi8770, pi8771, pi8772, pi8773,
    pi8774, pi8775, pi8776, pi8777, pi8778, pi8779, pi8780, pi8781, pi8782,
    pi8783, pi8784, pi8785, pi8786, pi8787, pi8788, pi8789, pi8790, pi8791,
    pi8792, pi8793, pi8794, pi8795, pi8796, pi8797, pi8798, pi8799, pi8800,
    pi8801, pi8802, pi8803, pi8804, pi8805, pi8806, pi8807, pi8808, pi8809,
    pi8810, pi8811, pi8812, pi8813, pi8814, pi8815, pi8816, pi8817, pi8818,
    pi8819, pi8820, pi8821, pi8822, pi8823, pi8824, pi8825, pi8826, pi8827,
    pi8828, pi8829, pi8830, pi8831, pi8832, pi8833, pi8834, pi8835, pi8836,
    pi8837, pi8838, pi8839, pi8840, pi8841, pi8842, pi8843, pi8844, pi8845,
    pi8846, pi8847, pi8848, pi8849, pi8850, pi8851, pi8852, pi8853, pi8854,
    pi8855, pi8856, pi8857, pi8858, pi8859, pi8860, pi8861, pi8862, pi8863,
    pi8864, pi8865, pi8866, pi8867, pi8868, pi8869, pi8870, pi8871, pi8872,
    pi8873, pi8874, pi8875, pi8876, pi8877, pi8878, pi8879, pi8880, pi8881,
    pi8882, pi8883, pi8884, pi8885, pi8886, pi8887, pi8888, pi8889, pi8890,
    pi8891, pi8892, pi8893, pi8894, pi8895, pi8896, pi8897, pi8898, pi8899,
    pi8900, pi8901, pi8902, pi8903, pi8904, pi8905, pi8906, pi8907, pi8908,
    pi8909, pi8910, pi8911, pi8912, pi8913, pi8914, pi8915, pi8916, pi8917,
    pi8918, pi8919, pi8920, pi8921, pi8922, pi8923, pi8924, pi8925, pi8926,
    pi8927, pi8928, pi8929, pi8930, pi8931, pi8932, pi8933, pi8934, pi8935,
    pi8936, pi8937, pi8938, pi8939, pi8940, pi8941, pi8942, pi8943, pi8944,
    pi8945, pi8946, pi8947, pi8948, pi8949, pi8950, pi8951, pi8952, pi8953,
    pi8954, pi8955, pi8956, pi8957, pi8958, pi8959, pi8960, pi8961, pi8962,
    pi8963, pi8964, pi8965, pi8966, pi8967, pi8968, pi8969, pi8970, pi8971,
    pi8972, pi8973, pi8974, pi8975, pi8976, pi8977, pi8978, pi8979, pi8980,
    pi8981, pi8982, pi8983, pi8984, pi8985, pi8986, pi8987, pi8988, pi8989,
    pi8990, pi8991, pi8992, pi8993, pi8994, pi8995, pi8996, pi8997, pi8998,
    pi8999, pi9000, pi9001, pi9002, pi9003, pi9004, pi9005, pi9006, pi9007,
    pi9008, pi9009, pi9010, pi9011, pi9012, pi9013, pi9014, pi9015, pi9016,
    pi9017, pi9018, pi9019, pi9020, pi9021, pi9022, pi9023, pi9024, pi9025,
    pi9026, pi9027, pi9028, pi9029, pi9030, pi9031, pi9032, pi9033, pi9034,
    pi9035, pi9036, pi9037, pi9038, pi9039, pi9040, pi9041;
  output po0000, po0001, po0002, po0003, po0004, po0005, po0006, po0007,
    po0008, po0009, po0010, po0011, po0012, po0013, po0014, po0015, po0016,
    po0017, po0018, po0019, po0020, po0021, po0022, po0023, po0024, po0025,
    po0026, po0027, po0028, po0029, po0030, po0031, po0032, po0033, po0034,
    po0035, po0036, po0037, po0038, po0039, po0040, po0041, po0042, po0043,
    po0044, po0045, po0046, po0047, po0048, po0049, po0050, po0051, po0052,
    po0053, po0054, po0055, po0056, po0057, po0058, po0059, po0060, po0061,
    po0062, po0063, po0064, po0065, po0066, po0067, po0068, po0069, po0070,
    po0071, po0072, po0073, po0074, po0075, po0076, po0077, po0078, po0079,
    po0080, po0081, po0082, po0083, po0084, po0085, po0086, po0087, po0088,
    po0089, po0090, po0091, po0092, po0093, po0094, po0095, po0096, po0097,
    po0098, po0099, po0100, po0101, po0102, po0103, po0104, po0105, po0106,
    po0107, po0108, po0109, po0110, po0111, po0112, po0113, po0114, po0115,
    po0116, po0117, po0118, po0119, po0120, po0121, po0122, po0123, po0124,
    po0125, po0126, po0127, po0128, po0129, po0130, po0131, po0132, po0133,
    po0134, po0135, po0136, po0137, po0138, po0139, po0140, po0141, po0142,
    po0143, po0144, po0145, po0146, po0147, po0148, po0149, po0150, po0151,
    po0152, po0153, po0154, po0155, po0156, po0157, po0158, po0159, po0160,
    po0161, po0162, po0163, po0164, po0165, po0166, po0167, po0168, po0169,
    po0170, po0171, po0172, po0173, po0174, po0175, po0176, po0177, po0178,
    po0179, po0180, po0181, po0182, po0183, po0184, po0185, po0186, po0187,
    po0188, po0189, po0190, po0191, po0192, po0193, po0194, po0195, po0196,
    po0197, po0198, po0199, po0200, po0201, po0202, po0203, po0204, po0205,
    po0206, po0207, po0208, po0209, po0210, po0211, po0212, po0213, po0214,
    po0215, po0216, po0217, po0218, po0219, po0220, po0221, po0222, po0223,
    po0224, po0225, po0226, po0227, po0228, po0229, po0230, po0231, po0232,
    po0233, po0234, po0235, po0236, po0237, po0238, po0239, po0240, po0241,
    po0242, po0243, po0244, po0245, po0246, po0247, po0248, po0249, po0250,
    po0251, po0252, po0253, po0254, po0255, po0256, po0257, po0258, po0259,
    po0260, po0261, po0262, po0263, po0264, po0265, po0266, po0267, po0268,
    po0269, po0270, po0271, po0272, po0273, po0274, po0275, po0276, po0277,
    po0278, po0279, po0280, po0281, po0282, po0283, po0284, po0285, po0286,
    po0287, po0288, po0289, po0290, po0291, po0292, po0293, po0294, po0295,
    po0296, po0297, po0298, po0299, po0300, po0301, po0302, po0303, po0304,
    po0305, po0306, po0307, po0308, po0309, po0310, po0311, po0312, po0313,
    po0314, po0315, po0316, po0317, po0318, po0319, po0320, po0321, po0322,
    po0323, po0324, po0325, po0326, po0327, po0328, po0329, po0330, po0331,
    po0332, po0333, po0334, po0335, po0336, po0337, po0338, po0339, po0340,
    po0341, po0342, po0343, po0344, po0345, po0346, po0347, po0348, po0349,
    po0350, po0351, po0352, po0353, po0354, po0355, po0356, po0357, po0358,
    po0359, po0360, po0361, po0362, po0363, po0364, po0365, po0366, po0367,
    po0368, po0369, po0370, po0371, po0372, po0373, po0374, po0375, po0376,
    po0377, po0378, po0379, po0380, po0381, po0382, po0383, po0384, po0385,
    po0386, po0387, po0388, po0389, po0390, po0391, po0392, po0393, po0394,
    po0395, po0396, po0397, po0398, po0399, po0400, po0401, po0402, po0403,
    po0404, po0405, po0406, po0407, po0408, po0409, po0410, po0411, po0412,
    po0413, po0414, po0415, po0416, po0417, po0418, po0419, po0420, po0421,
    po0422, po0423, po0424, po0425, po0426, po0427, po0428, po0429, po0430,
    po0431, po0432, po0433, po0434, po0435, po0436, po0437, po0438, po0439,
    po0440, po0441, po0442, po0443, po0444, po0445, po0446, po0447, po0448,
    po0449, po0450, po0451, po0452, po0453, po0454, po0455, po0456, po0457,
    po0458, po0459, po0460, po0461, po0462, po0463, po0464, po0465, po0466,
    po0467, po0468, po0469, po0470, po0471, po0472, po0473, po0474, po0475,
    po0476, po0477, po0478, po0479, po0480, po0481, po0482, po0483, po0484,
    po0485, po0486, po0487, po0488, po0489, po0490, po0491, po0492, po0493,
    po0494, po0495, po0496, po0497, po0498, po0499, po0500, po0501, po0502,
    po0503, po0504, po0505, po0506, po0507, po0508, po0509, po0510, po0511,
    po0512, po0513, po0514, po0515, po0516, po0517, po0518, po0519, po0520,
    po0521, po0522, po0523, po0524, po0525, po0526, po0527, po0528, po0529,
    po0530, po0531, po0532, po0533, po0534, po0535, po0536, po0537, po0538,
    po0539, po0540, po0541, po0542, po0543, po0544, po0545, po0546, po0547,
    po0548, po0549, po0550, po0551, po0552, po0553, po0554, po0555, po0556,
    po0557, po0558, po0559, po0560, po0561, po0562, po0563, po0564, po0565,
    po0566, po0567, po0568, po0569, po0570, po0571, po0572, po0573, po0574,
    po0575, po0576, po0577, po0578, po0579, po0580, po0581, po0582, po0583,
    po0584, po0585, po0586, po0587, po0588, po0589, po0590, po0591, po0592,
    po0593, po0594, po0595, po0596, po0597, po0598, po0599, po0600, po0601,
    po0602, po0603, po0604, po0605, po0606, po0607, po0608, po0609, po0610,
    po0611, po0612, po0613, po0614, po0615, po0616, po0617, po0618, po0619,
    po0620, po0621, po0622, po0623, po0624, po0625, po0626, po0627, po0628,
    po0629, po0630, po0631, po0632, po0633, po0634, po0635, po0636, po0637,
    po0638, po0639, po0640, po0641, po0642, po0643, po0644, po0645, po0646,
    po0647, po0648, po0649, po0650, po0651, po0652, po0653, po0654, po0655,
    po0656, po0657, po0658, po0659, po0660, po0661, po0662, po0663, po0664,
    po0665, po0666, po0667, po0668, po0669, po0670, po0671, po0672, po0673,
    po0674, po0675, po0676, po0677, po0678, po0679, po0680, po0681, po0682,
    po0683, po0684, po0685, po0686, po0687, po0688, po0689, po0690, po0691,
    po0692, po0693, po0694, po0695, po0696, po0697, po0698, po0699, po0700,
    po0701, po0702, po0703, po0704, po0705, po0706, po0707, po0708, po0709,
    po0710, po0711, po0712, po0713, po0714, po0715, po0716, po0717, po0718,
    po0719, po0720, po0721, po0722, po0723, po0724, po0725, po0726, po0727,
    po0728, po0729, po0730, po0731, po0732, po0733, po0734, po0735, po0736,
    po0737, po0738, po0739, po0740, po0741, po0742, po0743, po0744, po0745,
    po0746, po0747, po0748, po0749, po0750, po0751, po0752, po0753, po0754,
    po0755, po0756, po0757, po0758, po0759, po0760, po0761, po0762, po0763,
    po0764, po0765, po0766, po0767, po0768, po0769, po0770, po0771, po0772,
    po0773, po0774, po0775, po0776, po0777, po0778, po0779, po0780, po0781,
    po0782, po0783, po0784, po0785, po0786, po0787, po0788, po0789, po0790,
    po0791, po0792, po0793, po0794, po0795, po0796, po0797, po0798, po0799,
    po0800, po0801, po0802, po0803, po0804, po0805, po0806, po0807, po0808,
    po0809, po0810, po0811, po0812, po0813, po0814, po0815, po0816, po0817,
    po0818, po0819, po0820, po0821, po0822, po0823, po0824, po0825, po0826,
    po0827, po0828, po0829, po0830, po0831, po0832, po0833, po0834, po0835,
    po0836, po0837, po0838, po0839, po0840, po0841, po0842, po0843, po0844,
    po0845, po0846, po0847, po0848, po0849, po0850, po0851, po0852, po0853,
    po0854, po0855, po0856, po0857, po0858, po0859, po0860, po0861, po0862,
    po0863, po0864, po0865, po0866, po0867, po0868, po0869, po0870, po0871,
    po0872, po0873, po0874, po0875, po0876, po0877, po0878, po0879, po0880,
    po0881, po0882, po0883, po0884, po0885, po0886, po0887, po0888, po0889,
    po0890, po0891, po0892, po0893, po0894, po0895, po0896, po0897, po0898,
    po0899, po0900, po0901, po0902, po0903, po0904, po0905, po0906, po0907,
    po0908, po0909, po0910, po0911, po0912, po0913, po0914, po0915, po0916,
    po0917, po0918, po0919, po0920, po0921, po0922, po0923, po0924, po0925,
    po0926, po0927, po0928, po0929, po0930, po0931, po0932, po0933, po0934,
    po0935, po0936, po0937, po0938, po0939, po0940, po0941, po0942, po0943,
    po0944, po0945, po0946, po0947, po0948, po0949, po0950, po0951, po0952,
    po0953, po0954, po0955, po0956, po0957, po0958, po0959, po0960, po0961,
    po0962, po0963, po0964, po0965, po0966, po0967, po0968, po0969, po0970,
    po0971, po0972, po0973, po0974, po0975, po0976, po0977, po0978, po0979,
    po0980, po0981, po0982, po0983, po0984, po0985, po0986, po0987, po0988,
    po0989, po0990, po0991, po0992, po0993, po0994, po0995, po0996, po0997,
    po0998, po0999, po1000, po1001, po1002, po1003, po1004, po1005, po1006,
    po1007, po1008, po1009, po1010, po1011, po1012, po1013, po1014, po1015,
    po1016, po1017, po1018, po1019, po1020, po1021, po1022, po1023, po1024,
    po1025, po1026, po1027, po1028, po1029, po1030, po1031, po1032, po1033,
    po1034, po1035, po1036, po1037, po1038, po1039, po1040, po1041, po1042,
    po1043, po1044, po1045, po1046, po1047, po1048, po1049, po1050, po1051,
    po1052, po1053, po1054, po1055, po1056, po1057, po1058, po1059, po1060,
    po1061, po1062, po1063, po1064, po1065, po1066, po1067, po1068, po1069,
    po1070, po1071, po1072, po1073, po1074, po1075, po1076, po1077, po1078,
    po1079, po1080, po1081, po1082, po1083, po1084, po1085, po1086, po1087,
    po1088, po1089, po1090, po1091, po1092, po1093, po1094, po1095, po1096,
    po1097, po1098, po1099, po1100, po1101, po1102, po1103, po1104, po1105,
    po1106, po1107, po1108, po1109, po1110, po1111, po1112, po1113, po1114,
    po1115, po1116, po1117, po1118, po1119, po1120, po1121, po1122, po1123,
    po1124, po1125, po1126, po1127, po1128, po1129, po1130, po1131, po1132,
    po1133, po1134, po1135, po1136, po1137, po1138, po1139, po1140, po1141,
    po1142, po1143, po1144, po1145, po1146, po1147, po1148, po1149, po1150,
    po1151, po1152, po1153, po1154, po1155, po1156, po1157, po1158, po1159,
    po1160, po1161, po1162, po1163, po1164, po1165, po1166, po1167, po1168,
    po1169, po1170, po1171, po1172, po1173, po1174, po1175, po1176, po1177,
    po1178, po1179, po1180, po1181, po1182, po1183, po1184, po1185, po1186,
    po1187, po1188, po1189, po1190, po1191, po1192, po1193, po1194, po1195,
    po1196, po1197, po1198, po1199, po1200, po1201, po1202, po1203, po1204,
    po1205, po1206, po1207, po1208, po1209, po1210, po1211, po1212, po1213,
    po1214, po1215, po1216, po1217, po1218, po1219, po1220, po1221, po1222,
    po1223, po1224, po1225, po1226, po1227, po1228, po1229, po1230, po1231,
    po1232, po1233, po1234, po1235, po1236, po1237, po1238, po1239, po1240,
    po1241, po1242, po1243, po1244, po1245, po1246, po1247, po1248, po1249,
    po1250, po1251, po1252, po1253, po1254, po1255, po1256, po1257, po1258,
    po1259, po1260, po1261, po1262, po1263, po1264, po1265, po1266, po1267,
    po1268, po1269, po1270, po1271, po1272, po1273, po1274, po1275, po1276,
    po1277, po1278, po1279, po1280, po1281, po1282, po1283, po1284, po1285,
    po1286, po1287, po1288, po1289, po1290, po1291, po1292, po1293, po1294,
    po1295, po1296, po1297, po1298, po1299, po1300, po1301, po1302, po1303,
    po1304, po1305, po1306, po1307, po1308, po1309, po1310, po1311, po1312,
    po1313, po1314, po1315, po1316, po1317, po1318, po1319, po1320, po1321,
    po1322, po1323, po1324, po1325, po1326, po1327, po1328, po1329, po1330,
    po1331, po1332, po1333, po1334, po1335, po1336, po1337, po1338, po1339,
    po1340, po1341, po1342, po1343, po1344, po1345, po1346, po1347, po1348,
    po1349, po1350, po1351, po1352, po1353, po1354, po1355, po1356, po1357,
    po1358, po1359, po1360, po1361, po1362, po1363, po1364, po1365, po1366,
    po1367, po1368, po1369, po1370, po1371, po1372, po1373, po1374, po1375,
    po1376, po1377, po1378, po1379, po1380, po1381, po1382, po1383, po1384,
    po1385, po1386, po1387, po1388, po1389, po1390, po1391, po1392, po1393,
    po1394, po1395, po1396, po1397, po1398, po1399, po1400, po1401, po1402,
    po1403, po1404, po1405, po1406, po1407, po1408, po1409, po1410, po1411,
    po1412, po1413, po1414, po1415, po1416, po1417, po1418, po1419, po1420,
    po1421, po1422, po1423, po1424, po1425, po1426, po1427, po1428, po1429,
    po1430, po1431, po1432, po1433, po1434, po1435, po1436, po1437, po1438,
    po1439, po1440, po1441, po1442, po1443, po1444, po1445, po1446, po1447,
    po1448, po1449, po1450, po1451, po1452, po1453, po1454, po1455, po1456,
    po1457, po1458, po1459, po1460, po1461, po1462, po1463, po1464, po1465,
    po1466, po1467, po1468, po1469, po1470, po1471, po1472, po1473, po1474,
    po1475, po1476, po1477, po1478, po1479, po1480, po1481, po1482, po1483,
    po1484, po1485, po1486, po1487, po1488, po1489, po1490, po1491, po1492,
    po1493, po1494, po1495, po1496, po1497, po1498, po1499, po1500, po1501,
    po1502, po1503, po1504, po1505, po1506, po1507, po1508, po1509, po1510,
    po1511, po1512, po1513, po1514, po1515, po1516, po1517, po1518, po1519,
    po1520, po1521, po1522, po1523, po1524, po1525, po1526, po1527, po1528,
    po1529, po1530, po1531, po1532, po1533, po1534, po1535, po1536, po1537,
    po1538, po1539, po1540, po1541, po1542, po1543, po1544, po1545, po1546,
    po1547, po1548, po1549, po1550, po1551, po1552, po1553, po1554, po1555,
    po1556, po1557, po1558, po1559, po1560, po1561, po1562, po1563, po1564,
    po1565, po1566, po1567, po1568, po1569, po1570, po1571, po1572, po1573,
    po1574, po1575, po1576, po1577, po1578, po1579, po1580, po1581, po1582,
    po1583, po1584, po1585, po1586, po1587, po1588, po1589, po1590, po1591,
    po1592, po1593, po1594, po1595, po1596, po1597, po1598, po1599, po1600,
    po1601, po1602, po1603, po1604, po1605, po1606, po1607, po1608, po1609,
    po1610, po1611, po1612, po1613, po1614, po1615, po1616, po1617, po1618,
    po1619, po1620, po1621, po1622, po1623, po1624, po1625, po1626, po1627,
    po1628, po1629, po1630, po1631, po1632, po1633, po1634, po1635, po1636,
    po1637, po1638, po1639, po1640, po1641, po1642, po1643, po1644, po1645,
    po1646, po1647, po1648, po1649, po1650, po1651, po1652, po1653, po1654,
    po1655, po1656, po1657, po1658, po1659, po1660, po1661, po1662, po1663,
    po1664, po1665, po1666, po1667, po1668, po1669, po1670, po1671, po1672,
    po1673, po1674, po1675, po1676, po1677, po1678, po1679, po1680, po1681,
    po1682, po1683, po1684, po1685, po1686, po1687, po1688, po1689, po1690,
    po1691, po1692, po1693, po1694, po1695, po1696, po1697, po1698, po1699,
    po1700, po1701, po1702, po1703, po1704, po1705, po1706, po1707, po1708,
    po1709, po1710, po1711, po1712, po1713, po1714, po1715, po1716, po1717,
    po1718, po1719, po1720, po1721, po1722, po1723, po1724, po1725, po1726,
    po1727, po1728, po1729, po1730, po1731, po1732, po1733, po1734, po1735,
    po1736, po1737, po1738, po1739, po1740, po1741, po1742, po1743, po1744,
    po1745, po1746, po1747, po1748, po1749, po1750, po1751, po1752, po1753,
    po1754, po1755, po1756, po1757, po1758, po1759, po1760, po1761, po1762,
    po1763, po1764, po1765, po1766, po1767, po1768, po1769, po1770, po1771,
    po1772, po1773, po1774, po1775, po1776, po1777, po1778, po1779, po1780,
    po1781, po1782, po1783, po1784, po1785, po1786, po1787, po1788, po1789,
    po1790, po1791, po1792, po1793, po1794, po1795, po1796, po1797, po1798,
    po1799, po1800, po1801, po1802, po1803, po1804, po1805, po1806, po1807,
    po1808, po1809, po1810, po1811, po1812, po1813, po1814, po1815, po1816,
    po1817, po1818, po1819, po1820, po1821, po1822, po1823, po1824, po1825,
    po1826, po1827, po1828, po1829, po1830, po1831, po1832, po1833, po1834,
    po1835, po1836, po1837, po1838, po1839, po1840, po1841, po1842, po1843,
    po1844, po1845, po1846, po1847, po1848, po1849, po1850, po1851, po1852,
    po1853, po1854, po1855, po1856, po1857, po1858, po1859, po1860, po1861,
    po1862, po1863, po1864, po1865, po1866, po1867, po1868, po1869, po1870,
    po1871, po1872, po1873, po1874, po1875, po1876, po1877, po1878, po1879,
    po1880, po1881, po1882, po1883, po1884, po1885, po1886, po1887, po1888,
    po1889, po1890, po1891, po1892, po1893, po1894, po1895, po1896, po1897,
    po1898, po1899, po1900, po1901, po1902, po1903, po1904, po1905, po1906,
    po1907, po1908, po1909, po1910, po1911, po1912, po1913, po1914, po1915,
    po1916, po1917, po1918, po1919, po1920, po1921, po1922, po1923, po1924,
    po1925, po1926, po1927, po1928, po1929, po1930, po1931, po1932, po1933,
    po1934, po1935, po1936, po1937, po1938, po1939, po1940, po1941, po1942,
    po1943, po1944, po1945, po1946, po1947, po1948, po1949, po1950, po1951,
    po1952, po1953, po1954, po1955, po1956, po1957, po1958, po1959, po1960,
    po1961, po1962, po1963, po1964, po1965, po1966, po1967, po1968, po1969,
    po1970, po1971, po1972, po1973, po1974, po1975, po1976, po1977, po1978,
    po1979, po1980, po1981, po1982, po1983, po1984, po1985, po1986, po1987,
    po1988, po1989, po1990, po1991, po1992, po1993, po1994, po1995, po1996,
    po1997, po1998, po1999, po2000, po2001, po2002, po2003, po2004, po2005,
    po2006, po2007, po2008, po2009, po2010, po2011, po2012, po2013, po2014,
    po2015, po2016, po2017, po2018, po2019, po2020, po2021, po2022, po2023,
    po2024, po2025, po2026, po2027, po2028, po2029, po2030, po2031, po2032,
    po2033, po2034, po2035, po2036, po2037, po2038, po2039, po2040, po2041,
    po2042, po2043, po2044, po2045, po2046, po2047, po2048, po2049, po2050,
    po2051, po2052, po2053, po2054, po2055, po2056, po2057, po2058, po2059,
    po2060, po2061, po2062, po2063, po2064, po2065, po2066, po2067, po2068,
    po2069, po2070, po2071, po2072, po2073, po2074, po2075, po2076, po2077,
    po2078, po2079, po2080, po2081, po2082, po2083, po2084, po2085, po2086,
    po2087, po2088, po2089, po2090, po2091, po2092, po2093, po2094, po2095,
    po2096, po2097, po2098, po2099, po2100, po2101, po2102, po2103, po2104,
    po2105, po2106, po2107, po2108, po2109, po2110, po2111, po2112, po2113,
    po2114, po2115, po2116, po2117, po2118, po2119, po2120, po2121, po2122,
    po2123, po2124, po2125, po2126, po2127, po2128, po2129, po2130, po2131,
    po2132, po2133, po2134, po2135, po2136, po2137, po2138, po2139, po2140,
    po2141, po2142, po2143, po2144, po2145, po2146, po2147, po2148, po2149,
    po2150, po2151, po2152, po2153, po2154, po2155, po2156, po2157, po2158,
    po2159, po2160, po2161, po2162, po2163, po2164, po2165, po2166, po2167,
    po2168, po2169, po2170, po2171, po2172, po2173, po2174, po2175, po2176,
    po2177, po2178, po2179, po2180, po2181, po2182, po2183, po2184, po2185,
    po2186, po2187, po2188, po2189, po2190, po2191, po2192, po2193, po2194,
    po2195, po2196, po2197, po2198, po2199, po2200, po2201, po2202, po2203,
    po2204, po2205, po2206, po2207, po2208, po2209, po2210, po2211, po2212,
    po2213, po2214, po2215, po2216, po2217, po2218, po2219, po2220, po2221,
    po2222, po2223, po2224, po2225, po2226, po2227, po2228, po2229, po2230,
    po2231, po2232, po2233, po2234, po2235, po2236, po2237, po2238, po2239,
    po2240, po2241, po2242, po2243, po2244, po2245, po2246, po2247, po2248,
    po2249, po2250, po2251, po2252, po2253, po2254, po2255, po2256, po2257,
    po2258, po2259, po2260, po2261, po2262, po2263, po2264, po2265, po2266,
    po2267, po2268, po2269, po2270, po2271, po2272, po2273, po2274, po2275,
    po2276, po2277, po2278, po2279, po2280, po2281, po2282, po2283, po2284,
    po2285, po2286, po2287, po2288, po2289, po2290, po2291, po2292, po2293,
    po2294, po2295, po2296, po2297, po2298, po2299, po2300, po2301, po2302,
    po2303, po2304, po2305, po2306, po2307, po2308, po2309, po2310, po2311,
    po2312, po2313, po2314, po2315, po2316, po2317, po2318, po2319, po2320,
    po2321, po2322, po2323, po2324, po2325, po2326, po2327, po2328, po2329,
    po2330, po2331, po2332, po2333, po2334, po2335, po2336, po2337, po2338,
    po2339, po2340, po2341, po2342, po2343, po2344, po2345, po2346, po2347,
    po2348, po2349, po2350, po2351, po2352, po2353, po2354, po2355, po2356,
    po2357, po2358, po2359, po2360, po2361, po2362, po2363, po2364, po2365,
    po2366, po2367, po2368, po2369, po2370, po2371, po2372, po2373, po2374,
    po2375, po2376, po2377, po2378, po2379, po2380, po2381, po2382, po2383,
    po2384, po2385, po2386, po2387, po2388, po2389, po2390, po2391, po2392,
    po2393, po2394, po2395, po2396, po2397, po2398, po2399, po2400, po2401,
    po2402, po2403, po2404, po2405, po2406, po2407, po2408, po2409, po2410,
    po2411, po2412, po2413, po2414, po2415, po2416, po2417, po2418, po2419,
    po2420, po2421, po2422, po2423, po2424, po2425, po2426, po2427, po2428,
    po2429, po2430, po2431, po2432, po2433, po2434, po2435, po2436, po2437,
    po2438, po2439, po2440, po2441, po2442, po2443, po2444, po2445, po2446,
    po2447, po2448, po2449, po2450, po2451, po2452, po2453, po2454, po2455,
    po2456, po2457, po2458, po2459, po2460, po2461, po2462, po2463, po2464,
    po2465, po2466, po2467, po2468, po2469, po2470, po2471, po2472, po2473,
    po2474, po2475, po2476, po2477, po2478, po2479, po2480, po2481, po2482,
    po2483, po2484, po2485, po2486, po2487, po2488, po2489, po2490, po2491,
    po2492, po2493, po2494, po2495, po2496, po2497, po2498, po2499, po2500,
    po2501, po2502, po2503, po2504, po2505, po2506, po2507, po2508, po2509,
    po2510, po2511, po2512, po2513, po2514, po2515, po2516, po2517, po2518,
    po2519, po2520, po2521, po2522, po2523, po2524, po2525, po2526, po2527,
    po2528, po2529, po2530, po2531, po2532, po2533, po2534, po2535, po2536,
    po2537, po2538, po2539, po2540, po2541, po2542, po2543, po2544, po2545,
    po2546, po2547, po2548, po2549, po2550, po2551, po2552, po2553, po2554,
    po2555, po2556, po2557, po2558, po2559, po2560, po2561, po2562, po2563,
    po2564, po2565, po2566, po2567, po2568, po2569, po2570, po2571, po2572,
    po2573, po2574, po2575, po2576, po2577, po2578, po2579, po2580, po2581,
    po2582, po2583, po2584, po2585, po2586, po2587, po2588, po2589, po2590,
    po2591, po2592, po2593, po2594, po2595, po2596, po2597, po2598, po2599,
    po2600, po2601, po2602, po2603, po2604, po2605, po2606, po2607, po2608,
    po2609, po2610, po2611, po2612, po2613, po2614, po2615, po2616, po2617,
    po2618, po2619, po2620, po2621, po2622, po2623, po2624, po2625, po2626,
    po2627, po2628, po2629, po2630, po2631, po2632, po2633, po2634, po2635,
    po2636, po2637, po2638, po2639, po2640, po2641, po2642, po2643, po2644,
    po2645, po2646, po2647, po2648, po2649, po2650, po2651, po2652, po2653,
    po2654, po2655, po2656, po2657, po2658, po2659, po2660, po2661, po2662,
    po2663, po2664, po2665, po2666, po2667, po2668, po2669, po2670, po2671,
    po2672, po2673, po2674, po2675, po2676, po2677, po2678, po2679, po2680,
    po2681, po2682, po2683, po2684, po2685, po2686, po2687, po2688, po2689,
    po2690, po2691, po2692, po2693, po2694, po2695, po2696, po2697, po2698,
    po2699, po2700, po2701, po2702, po2703, po2704, po2705, po2706, po2707,
    po2708, po2709, po2710, po2711, po2712, po2713, po2714, po2715, po2716,
    po2717, po2718, po2719, po2720, po2721, po2722, po2723, po2724, po2725,
    po2726, po2727, po2728, po2729, po2730, po2731, po2732, po2733, po2734,
    po2735, po2736, po2737, po2738, po2739, po2740, po2741, po2742, po2743,
    po2744, po2745, po2746, po2747, po2748, po2749, po2750, po2751, po2752,
    po2753, po2754, po2755, po2756, po2757, po2758, po2759, po2760, po2761,
    po2762, po2763, po2764, po2765, po2766, po2767, po2768, po2769, po2770,
    po2771, po2772, po2773, po2774, po2775, po2776, po2777, po2778, po2779,
    po2780, po2781, po2782, po2783, po2784, po2785, po2786, po2787, po2788,
    po2789, po2790, po2791, po2792, po2793, po2794, po2795, po2796, po2797,
    po2798, po2799, po2800, po2801, po2802, po2803, po2804, po2805, po2806,
    po2807, po2808, po2809, po2810, po2811, po2812, po2813, po2814, po2815,
    po2816, po2817, po2818, po2819, po2820, po2821, po2822, po2823, po2824,
    po2825, po2826, po2827, po2828, po2829, po2830, po2831, po2832, po2833,
    po2834, po2835, po2836, po2837, po2838, po2839, po2840, po2841, po2842,
    po2843, po2844, po2845, po2846, po2847, po2848, po2849, po2850, po2851,
    po2852, po2853, po2854, po2855, po2856, po2857, po2858, po2859, po2860,
    po2861, po2862, po2863, po2864, po2865, po2866, po2867, po2868, po2869,
    po2870, po2871, po2872, po2873, po2874, po2875, po2876, po2877, po2878,
    po2879, po2880, po2881, po2882, po2883, po2884, po2885, po2886, po2887,
    po2888, po2889, po2890, po2891, po2892, po2893, po2894, po2895, po2896,
    po2897, po2898, po2899, po2900, po2901, po2902, po2903, po2904, po2905,
    po2906, po2907, po2908, po2909, po2910, po2911, po2912, po2913, po2914,
    po2915, po2916, po2917, po2918, po2919, po2920, po2921, po2922, po2923,
    po2924, po2925, po2926, po2927, po2928, po2929, po2930, po2931, po2932,
    po2933, po2934, po2935, po2936, po2937, po2938, po2939, po2940, po2941,
    po2942, po2943, po2944, po2945, po2946, po2947, po2948, po2949, po2950,
    po2951, po2952, po2953, po2954, po2955, po2956, po2957, po2958, po2959,
    po2960, po2961, po2962, po2963, po2964, po2965, po2966, po2967, po2968,
    po2969, po2970, po2971, po2972, po2973, po2974, po2975, po2976, po2977,
    po2978, po2979, po2980, po2981, po2982, po2983, po2984, po2985, po2986,
    po2987, po2988, po2989, po2990, po2991, po2992, po2993, po2994, po2995,
    po2996, po2997, po2998, po2999, po3000, po3001, po3002, po3003, po3004,
    po3005, po3006, po3007, po3008, po3009, po3010, po3011, po3012, po3013,
    po3014, po3015, po3016, po3017, po3018, po3019, po3020, po3021, po3022,
    po3023, po3024, po3025, po3026, po3027, po3028, po3029, po3030, po3031,
    po3032, po3033, po3034, po3035, po3036, po3037, po3038, po3039, po3040,
    po3041, po3042, po3043, po3044, po3045, po3046, po3047, po3048, po3049,
    po3050, po3051, po3052, po3053, po3054, po3055, po3056, po3057, po3058,
    po3059, po3060, po3061, po3062, po3063, po3064, po3065, po3066, po3067,
    po3068, po3069, po3070, po3071, po3072, po3073, po3074, po3075, po3076,
    po3077, po3078, po3079, po3080, po3081, po3082, po3083, po3084, po3085,
    po3086, po3087, po3088, po3089, po3090, po3091, po3092, po3093, po3094,
    po3095, po3096, po3097, po3098, po3099, po3100, po3101, po3102, po3103,
    po3104, po3105, po3106, po3107, po3108, po3109, po3110, po3111, po3112,
    po3113, po3114, po3115, po3116, po3117, po3118, po3119, po3120, po3121,
    po3122, po3123, po3124, po3125, po3126, po3127, po3128, po3129, po3130,
    po3131, po3132, po3133, po3134, po3135, po3136, po3137, po3138, po3139,
    po3140, po3141, po3142, po3143, po3144, po3145, po3146, po3147, po3148,
    po3149, po3150, po3151, po3152, po3153, po3154, po3155, po3156, po3157,
    po3158, po3159, po3160, po3161, po3162, po3163, po3164, po3165, po3166,
    po3167, po3168, po3169, po3170, po3171, po3172, po3173, po3174, po3175,
    po3176, po3177, po3178, po3179, po3180, po3181, po3182, po3183, po3184,
    po3185, po3186, po3187, po3188, po3189, po3190, po3191, po3192, po3193,
    po3194, po3195, po3196, po3197, po3198, po3199, po3200, po3201, po3202,
    po3203, po3204, po3205, po3206, po3207, po3208, po3209, po3210, po3211,
    po3212, po3213, po3214, po3215, po3216, po3217, po3218, po3219, po3220,
    po3221, po3222, po3223, po3224, po3225, po3226, po3227, po3228, po3229,
    po3230, po3231, po3232, po3233, po3234, po3235, po3236, po3237, po3238,
    po3239, po3240, po3241, po3242, po3243, po3244, po3245, po3246, po3247,
    po3248, po3249, po3250, po3251, po3252, po3253, po3254, po3255, po3256,
    po3257, po3258, po3259, po3260, po3261, po3262, po3263, po3264, po3265,
    po3266, po3267, po3268, po3269, po3270, po3271, po3272, po3273, po3274,
    po3275, po3276, po3277, po3278, po3279, po3280, po3281, po3282, po3283,
    po3284, po3285, po3286, po3287, po3288, po3289, po3290, po3291, po3292,
    po3293, po3294, po3295, po3296, po3297, po3298, po3299, po3300, po3301,
    po3302, po3303, po3304, po3305, po3306, po3307, po3308, po3309, po3310,
    po3311, po3312, po3313, po3314, po3315, po3316, po3317, po3318, po3319,
    po3320, po3321, po3322, po3323, po3324, po3325, po3326, po3327, po3328,
    po3329, po3330, po3331, po3332, po3333, po3334, po3335, po3336, po3337,
    po3338, po3339, po3340, po3341, po3342, po3343, po3344, po3345, po3346,
    po3347, po3348, po3349, po3350, po3351, po3352, po3353, po3354, po3355,
    po3356, po3357, po3358, po3359, po3360, po3361, po3362, po3363, po3364,
    po3365, po3366, po3367, po3368, po3369, po3370, po3371, po3372, po3373,
    po3374, po3375, po3376, po3377, po3378, po3379, po3380, po3381, po3382,
    po3383, po3384, po3385, po3386, po3387, po3388, po3389, po3390, po3391,
    po3392, po3393, po3394, po3395, po3396, po3397, po3398, po3399, po3400,
    po3401, po3402, po3403, po3404, po3405, po3406, po3407, po3408, po3409,
    po3410, po3411, po3412, po3413, po3414, po3415, po3416, po3417, po3418,
    po3419, po3420, po3421, po3422, po3423, po3424, po3425, po3426, po3427,
    po3428, po3429, po3430, po3431, po3432, po3433, po3434, po3435, po3436,
    po3437, po3438, po3439, po3440, po3441, po3442, po3443, po3444, po3445,
    po3446, po3447, po3448, po3449, po3450, po3451, po3452, po3453, po3454,
    po3455, po3456, po3457, po3458, po3459, po3460, po3461, po3462, po3463,
    po3464, po3465, po3466, po3467, po3468, po3469, po3470, po3471, po3472,
    po3473, po3474, po3475, po3476, po3477, po3478, po3479, po3480, po3481,
    po3482, po3483, po3484, po3485, po3486, po3487, po3488, po3489, po3490,
    po3491, po3492, po3493, po3494, po3495, po3496, po3497, po3498, po3499,
    po3500, po3501, po3502, po3503, po3504, po3505, po3506, po3507, po3508,
    po3509, po3510, po3511, po3512, po3513, po3514, po3515, po3516, po3517,
    po3518, po3519, po3520, po3521, po3522, po3523, po3524, po3525, po3526,
    po3527, po3528, po3529, po3530, po3531, po3532, po3533, po3534, po3535,
    po3536, po3537, po3538, po3539, po3540, po3541, po3542, po3543, po3544,
    po3545, po3546, po3547, po3548, po3549, po3550, po3551, po3552, po3553,
    po3554, po3555, po3556, po3557, po3558, po3559, po3560, po3561, po3562,
    po3563, po3564, po3565, po3566, po3567, po3568, po3569, po3570, po3571,
    po3572, po3573, po3574, po3575, po3576, po3577, po3578, po3579, po3580,
    po3581, po3582, po3583, po3584, po3585, po3586, po3587, po3588, po3589,
    po3590, po3591, po3592, po3593, po3594, po3595, po3596, po3597, po3598,
    po3599, po3600, po3601, po3602, po3603, po3604, po3605, po3606, po3607,
    po3608, po3609, po3610, po3611, po3612, po3613, po3614, po3615, po3616,
    po3617, po3618, po3619, po3620, po3621, po3622, po3623, po3624, po3625,
    po3626, po3627, po3628, po3629, po3630, po3631, po3632, po3633, po3634,
    po3635, po3636, po3637, po3638, po3639, po3640, po3641, po3642, po3643,
    po3644, po3645, po3646, po3647, po3648, po3649, po3650, po3651, po3652,
    po3653, po3654, po3655, po3656, po3657, po3658, po3659, po3660, po3661,
    po3662, po3663, po3664, po3665, po3666, po3667, po3668, po3669, po3670,
    po3671, po3672, po3673, po3674, po3675, po3676, po3677, po3678, po3679,
    po3680, po3681, po3682, po3683, po3684, po3685, po3686, po3687, po3688,
    po3689, po3690, po3691, po3692, po3693, po3694, po3695, po3696, po3697,
    po3698, po3699, po3700, po3701, po3702, po3703, po3704, po3705, po3706,
    po3707, po3708, po3709, po3710, po3711, po3712, po3713, po3714, po3715,
    po3716, po3717, po3718, po3719, po3720, po3721, po3722, po3723, po3724,
    po3725, po3726, po3727, po3728, po3729, po3730, po3731, po3732, po3733,
    po3734, po3735, po3736, po3737, po3738, po3739, po3740, po3741, po3742,
    po3743, po3744, po3745, po3746, po3747, po3748, po3749, po3750, po3751,
    po3752, po3753, po3754, po3755, po3756, po3757, po3758, po3759, po3760,
    po3761, po3762, po3763, po3764, po3765, po3766, po3767, po3768, po3769,
    po3770, po3771, po3772, po3773, po3774, po3775, po3776, po3777, po3778,
    po3779, po3780, po3781, po3782, po3783, po3784, po3785, po3786, po3787,
    po3788, po3789, po3790, po3791, po3792, po3793, po3794, po3795, po3796,
    po3797, po3798, po3799, po3800, po3801, po3802, po3803, po3804, po3805,
    po3806, po3807, po3808, po3809, po3810, po3811, po3812, po3813, po3814,
    po3815, po3816, po3817, po3818, po3819, po3820, po3821, po3822, po3823,
    po3824, po3825, po3826, po3827, po3828, po3829, po3830, po3831, po3832,
    po3833, po3834, po3835, po3836, po3837, po3838, po3839, po3840, po3841,
    po3842, po3843, po3844, po3845, po3846, po3847, po3848, po3849, po3850,
    po3851, po3852, po3853, po3854, po3855, po3856, po3857, po3858, po3859,
    po3860, po3861, po3862, po3863, po3864, po3865, po3866, po3867, po3868,
    po3869, po3870, po3871, po3872, po3873, po3874, po3875, po3876, po3877,
    po3878, po3879, po3880, po3881, po3882, po3883, po3884, po3885, po3886,
    po3887, po3888, po3889, po3890, po3891, po3892, po3893, po3894, po3895,
    po3896, po3897, po3898, po3899, po3900, po3901, po3902, po3903, po3904,
    po3905, po3906, po3907, po3908, po3909, po3910, po3911, po3912, po3913,
    po3914, po3915, po3916, po3917, po3918, po3919, po3920, po3921, po3922,
    po3923, po3924, po3925, po3926, po3927, po3928, po3929, po3930, po3931,
    po3932, po3933, po3934, po3935, po3936, po3937, po3938, po3939, po3940,
    po3941, po3942, po3943, po3944, po3945, po3946, po3947, po3948, po3949,
    po3950, po3951, po3952, po3953, po3954, po3955, po3956, po3957, po3958,
    po3959, po3960, po3961, po3962, po3963, po3964, po3965, po3966, po3967,
    po3968, po3969, po3970, po3971, po3972, po3973, po3974, po3975, po3976,
    po3977, po3978, po3979, po3980, po3981, po3982, po3983, po3984, po3985,
    po3986, po3987, po3988, po3989, po3990, po3991, po3992, po3993, po3994,
    po3995, po3996, po3997, po3998, po3999, po4000, po4001, po4002, po4003,
    po4004, po4005, po4006, po4007, po4008, po4009, po4010, po4011, po4012,
    po4013, po4014, po4015, po4016, po4017, po4018, po4019, po4020, po4021,
    po4022, po4023, po4024, po4025, po4026, po4027, po4028, po4029, po4030,
    po4031, po4032, po4033, po4034, po4035, po4036, po4037, po4038, po4039,
    po4040, po4041, po4042, po4043, po4044, po4045, po4046, po4047, po4048,
    po4049, po4050, po4051, po4052, po4053, po4054, po4055, po4056, po4057,
    po4058, po4059, po4060, po4061, po4062, po4063, po4064, po4065, po4066,
    po4067, po4068, po4069, po4070, po4071, po4072, po4073, po4074, po4075,
    po4076, po4077, po4078, po4079, po4080, po4081, po4082, po4083, po4084,
    po4085, po4086, po4087, po4088, po4089, po4090, po4091, po4092, po4093,
    po4094, po4095, po4096, po4097, po4098, po4099, po4100, po4101, po4102,
    po4103, po4104, po4105, po4106, po4107, po4108, po4109, po4110, po4111,
    po4112, po4113, po4114, po4115, po4116, po4117, po4118, po4119, po4120,
    po4121, po4122, po4123, po4124, po4125, po4126, po4127, po4128, po4129,
    po4130, po4131, po4132, po4133, po4134, po4135, po4136, po4137, po4138,
    po4139, po4140, po4141, po4142, po4143, po4144, po4145, po4146, po4147,
    po4148, po4149, po4150, po4151, po4152, po4153, po4154, po4155, po4156,
    po4157, po4158, po4159, po4160, po4161, po4162, po4163, po4164, po4165,
    po4166, po4167, po4168, po4169, po4170, po4171, po4172, po4173, po4174,
    po4175, po4176, po4177, po4178, po4179, po4180, po4181, po4182, po4183,
    po4184, po4185, po4186, po4187, po4188, po4189, po4190, po4191, po4192,
    po4193, po4194, po4195, po4196, po4197, po4198, po4199, po4200, po4201,
    po4202, po4203, po4204, po4205, po4206, po4207, po4208, po4209, po4210,
    po4211, po4212, po4213, po4214, po4215, po4216, po4217, po4218, po4219,
    po4220, po4221, po4222, po4223, po4224, po4225, po4226, po4227, po4228,
    po4229, po4230, po4231, po4232, po4233, po4234, po4235, po4236, po4237,
    po4238, po4239, po4240, po4241, po4242, po4243, po4244, po4245, po4246,
    po4247, po4248, po4249, po4250, po4251, po4252, po4253, po4254, po4255,
    po4256, po4257, po4258, po4259, po4260, po4261, po4262, po4263, po4264,
    po4265, po4266, po4267, po4268, po4269, po4270, po4271, po4272, po4273,
    po4274, po4275, po4276, po4277, po4278, po4279, po4280, po4281, po4282,
    po4283, po4284, po4285, po4286, po4287, po4288, po4289, po4290, po4291,
    po4292, po4293, po4294, po4295, po4296, po4297, po4298, po4299, po4300,
    po4301, po4302, po4303, po4304, po4305, po4306, po4307, po4308, po4309,
    po4310, po4311, po4312, po4313, po4314, po4315, po4316, po4317, po4318,
    po4319, po4320, po4321, po4322, po4323, po4324, po4325, po4326, po4327,
    po4328, po4329, po4330, po4331, po4332, po4333, po4334, po4335, po4336,
    po4337, po4338, po4339, po4340, po4341, po4342, po4343, po4344, po4345,
    po4346, po4347, po4348, po4349, po4350, po4351, po4352, po4353, po4354,
    po4355, po4356, po4357, po4358, po4359, po4360, po4361, po4362, po4363,
    po4364, po4365, po4366, po4367, po4368, po4369, po4370, po4371, po4372,
    po4373, po4374, po4375, po4376, po4377, po4378, po4379, po4380, po4381,
    po4382, po4383, po4384, po4385, po4386, po4387, po4388, po4389, po4390,
    po4391, po4392, po4393, po4394, po4395, po4396, po4397, po4398, po4399,
    po4400, po4401, po4402, po4403, po4404, po4405, po4406, po4407, po4408,
    po4409, po4410, po4411, po4412, po4413, po4414, po4415, po4416, po4417,
    po4418, po4419, po4420, po4421, po4422, po4423, po4424, po4425, po4426,
    po4427, po4428, po4429, po4430, po4431, po4432, po4433, po4434, po4435,
    po4436, po4437, po4438, po4439, po4440, po4441, po4442, po4443, po4444,
    po4445, po4446, po4447, po4448, po4449, po4450, po4451, po4452, po4453,
    po4454, po4455, po4456, po4457, po4458, po4459, po4460, po4461, po4462,
    po4463, po4464, po4465, po4466, po4467, po4468, po4469, po4470, po4471,
    po4472, po4473, po4474, po4475, po4476, po4477, po4478, po4479, po4480,
    po4481, po4482, po4483, po4484, po4485, po4486, po4487, po4488, po4489,
    po4490, po4491, po4492, po4493, po4494, po4495, po4496, po4497, po4498,
    po4499, po4500, po4501, po4502, po4503, po4504, po4505, po4506, po4507,
    po4508, po4509, po4510, po4511, po4512, po4513, po4514, po4515, po4516,
    po4517, po4518, po4519, po4520, po4521, po4522, po4523, po4524, po4525,
    po4526, po4527, po4528, po4529, po4530, po4531, po4532, po4533, po4534,
    po4535, po4536, po4537, po4538, po4539, po4540, po4541, po4542, po4543,
    po4544, po4545, po4546, po4547, po4548, po4549, po4550, po4551, po4552,
    po4553, po4554, po4555, po4556, po4557, po4558, po4559, po4560, po4561,
    po4562, po4563, po4564, po4565, po4566, po4567, po4568, po4569, po4570,
    po4571, po4572, po4573, po4574, po4575, po4576, po4577, po4578, po4579,
    po4580, po4581, po4582, po4583, po4584, po4585, po4586, po4587, po4588,
    po4589, po4590, po4591, po4592, po4593, po4594, po4595, po4596, po4597,
    po4598, po4599, po4600, po4601, po4602, po4603, po4604, po4605, po4606,
    po4607, po4608, po4609, po4610, po4611, po4612, po4613, po4614, po4615,
    po4616, po4617, po4618, po4619, po4620, po4621, po4622, po4623, po4624,
    po4625, po4626, po4627, po4628, po4629, po4630, po4631, po4632, po4633,
    po4634, po4635, po4636, po4637, po4638, po4639, po4640, po4641, po4642,
    po4643, po4644, po4645, po4646, po4647, po4648, po4649, po4650, po4651,
    po4652, po4653, po4654, po4655, po4656, po4657, po4658, po4659, po4660,
    po4661, po4662, po4663, po4664, po4665, po4666, po4667, po4668, po4669,
    po4670, po4671, po4672, po4673, po4674, po4675, po4676, po4677, po4678,
    po4679, po4680, po4681, po4682, po4683, po4684, po4685, po4686, po4687,
    po4688, po4689, po4690, po4691, po4692, po4693, po4694, po4695, po4696,
    po4697, po4698, po4699, po4700, po4701, po4702, po4703, po4704, po4705,
    po4706, po4707, po4708, po4709, po4710, po4711, po4712, po4713, po4714,
    po4715, po4716, po4717, po4718, po4719, po4720, po4721, po4722, po4723,
    po4724, po4725, po4726, po4727, po4728, po4729, po4730, po4731, po4732,
    po4733, po4734, po4735, po4736, po4737, po4738, po4739, po4740, po4741,
    po4742, po4743, po4744, po4745, po4746, po4747, po4748, po4749, po4750,
    po4751, po4752, po4753, po4754, po4755, po4756, po4757, po4758, po4759,
    po4760, po4761, po4762, po4763, po4764, po4765, po4766, po4767, po4768,
    po4769, po4770, po4771, po4772, po4773, po4774, po4775, po4776, po4777,
    po4778, po4779, po4780, po4781, po4782, po4783, po4784, po4785, po4786,
    po4787, po4788, po4789, po4790, po4791, po4792, po4793, po4794, po4795,
    po4796, po4797, po4798, po4799, po4800, po4801, po4802, po4803, po4804,
    po4805, po4806, po4807, po4808, po4809, po4810, po4811, po4812, po4813,
    po4814, po4815, po4816, po4817, po4818, po4819, po4820, po4821, po4822,
    po4823, po4824, po4825, po4826, po4827, po4828, po4829, po4830, po4831,
    po4832, po4833, po4834, po4835, po4836, po4837, po4838, po4839, po4840,
    po4841, po4842, po4843, po4844, po4845, po4846, po4847, po4848, po4849,
    po4850, po4851, po4852, po4853, po4854, po4855, po4856, po4857, po4858,
    po4859, po4860, po4861, po4862, po4863, po4864, po4865, po4866, po4867,
    po4868, po4869, po4870, po4871, po4872, po4873, po4874, po4875, po4876,
    po4877, po4878, po4879, po4880, po4881, po4882, po4883, po4884, po4885,
    po4886, po4887, po4888, po4889, po4890, po4891, po4892, po4893, po4894,
    po4895, po4896, po4897, po4898, po4899, po4900, po4901, po4902, po4903,
    po4904, po4905, po4906, po4907, po4908, po4909, po4910, po4911, po4912,
    po4913, po4914, po4915, po4916, po4917, po4918, po4919, po4920, po4921,
    po4922, po4923, po4924, po4925, po4926, po4927, po4928, po4929, po4930,
    po4931, po4932, po4933, po4934, po4935, po4936, po4937, po4938, po4939,
    po4940, po4941, po4942, po4943, po4944, po4945, po4946, po4947, po4948,
    po4949, po4950, po4951, po4952, po4953, po4954, po4955, po4956, po4957,
    po4958, po4959, po4960, po4961, po4962, po4963, po4964, po4965, po4966,
    po4967, po4968, po4969, po4970, po4971, po4972, po4973, po4974, po4975,
    po4976, po4977, po4978, po4979, po4980, po4981, po4982, po4983, po4984,
    po4985, po4986, po4987, po4988, po4989, po4990, po4991, po4992, po4993,
    po4994, po4995, po4996, po4997, po4998, po4999, po5000, po5001, po5002,
    po5003, po5004, po5005, po5006, po5007, po5008, po5009, po5010, po5011,
    po5012, po5013, po5014, po5015, po5016, po5017, po5018, po5019, po5020,
    po5021, po5022, po5023, po5024, po5025, po5026, po5027, po5028, po5029,
    po5030, po5031, po5032, po5033, po5034, po5035, po5036, po5037, po5038,
    po5039, po5040, po5041, po5042, po5043, po5044, po5045, po5046, po5047,
    po5048, po5049, po5050, po5051, po5052, po5053, po5054, po5055, po5056,
    po5057, po5058, po5059, po5060, po5061, po5062, po5063, po5064, po5065,
    po5066, po5067, po5068, po5069, po5070, po5071, po5072, po5073, po5074,
    po5075, po5076, po5077, po5078, po5079, po5080, po5081, po5082, po5083,
    po5084, po5085, po5086, po5087, po5088, po5089, po5090, po5091, po5092,
    po5093, po5094, po5095, po5096, po5097, po5098, po5099, po5100, po5101,
    po5102, po5103, po5104, po5105, po5106, po5107, po5108, po5109, po5110,
    po5111, po5112, po5113, po5114, po5115, po5116, po5117, po5118, po5119,
    po5120, po5121, po5122, po5123, po5124, po5125, po5126, po5127, po5128,
    po5129, po5130, po5131, po5132, po5133, po5134, po5135, po5136, po5137,
    po5138, po5139, po5140, po5141, po5142, po5143, po5144, po5145, po5146,
    po5147, po5148, po5149, po5150, po5151, po5152, po5153, po5154, po5155,
    po5156, po5157, po5158, po5159, po5160, po5161, po5162, po5163, po5164,
    po5165, po5166, po5167, po5168, po5169, po5170, po5171, po5172, po5173,
    po5174, po5175, po5176, po5177, po5178, po5179, po5180, po5181, po5182,
    po5183, po5184, po5185, po5186, po5187, po5188, po5189, po5190, po5191,
    po5192, po5193, po5194, po5195, po5196, po5197, po5198, po5199, po5200,
    po5201, po5202, po5203, po5204, po5205, po5206, po5207, po5208, po5209,
    po5210, po5211, po5212, po5213, po5214, po5215, po5216, po5217, po5218,
    po5219, po5220, po5221, po5222, po5223, po5224, po5225, po5226, po5227,
    po5228, po5229, po5230, po5231, po5232, po5233, po5234, po5235, po5236,
    po5237, po5238, po5239, po5240, po5241, po5242, po5243, po5244, po5245,
    po5246, po5247, po5248, po5249, po5250, po5251, po5252, po5253, po5254,
    po5255, po5256, po5257, po5258, po5259, po5260, po5261, po5262, po5263,
    po5264, po5265, po5266, po5267, po5268, po5269, po5270, po5271, po5272,
    po5273, po5274, po5275, po5276, po5277, po5278, po5279, po5280, po5281,
    po5282, po5283, po5284, po5285, po5286, po5287, po5288, po5289, po5290,
    po5291, po5292, po5293, po5294, po5295, po5296, po5297, po5298, po5299,
    po5300, po5301, po5302, po5303, po5304, po5305, po5306, po5307, po5308,
    po5309, po5310, po5311, po5312, po5313, po5314, po5315, po5316, po5317,
    po5318, po5319, po5320, po5321, po5322, po5323, po5324, po5325, po5326,
    po5327, po5328, po5329, po5330, po5331, po5332, po5333, po5334, po5335,
    po5336, po5337, po5338, po5339, po5340, po5341, po5342, po5343, po5344,
    po5345, po5346, po5347, po5348, po5349, po5350, po5351, po5352, po5353,
    po5354, po5355, po5356, po5357, po5358, po5359, po5360, po5361, po5362,
    po5363, po5364, po5365, po5366, po5367, po5368, po5369, po5370, po5371,
    po5372, po5373, po5374, po5375, po5376, po5377, po5378, po5379, po5380,
    po5381, po5382, po5383, po5384, po5385, po5386, po5387, po5388, po5389,
    po5390, po5391, po5392, po5393, po5394, po5395, po5396, po5397, po5398,
    po5399, po5400, po5401, po5402, po5403, po5404, po5405, po5406, po5407,
    po5408, po5409, po5410, po5411, po5412, po5413, po5414, po5415, po5416,
    po5417, po5418, po5419, po5420, po5421, po5422, po5423, po5424, po5425,
    po5426, po5427, po5428, po5429, po5430, po5431, po5432, po5433, po5434,
    po5435, po5436, po5437, po5438, po5439, po5440, po5441, po5442, po5443,
    po5444, po5445, po5446, po5447, po5448, po5449, po5450, po5451, po5452,
    po5453, po5454, po5455, po5456, po5457, po5458, po5459, po5460, po5461,
    po5462, po5463, po5464, po5465, po5466, po5467, po5468, po5469, po5470,
    po5471, po5472, po5473, po5474, po5475, po5476, po5477, po5478, po5479,
    po5480, po5481, po5482, po5483, po5484, po5485, po5486, po5487, po5488,
    po5489, po5490, po5491, po5492, po5493, po5494, po5495, po5496, po5497,
    po5498, po5499, po5500, po5501, po5502, po5503, po5504, po5505, po5506,
    po5507, po5508, po5509, po5510, po5511, po5512, po5513, po5514, po5515,
    po5516, po5517, po5518, po5519, po5520, po5521, po5522, po5523, po5524,
    po5525, po5526, po5527, po5528, po5529, po5530, po5531, po5532, po5533,
    po5534, po5535, po5536, po5537, po5538, po5539, po5540, po5541, po5542,
    po5543, po5544, po5545, po5546, po5547, po5548, po5549, po5550, po5551,
    po5552, po5553, po5554, po5555, po5556, po5557, po5558, po5559, po5560,
    po5561, po5562, po5563, po5564, po5565, po5566, po5567, po5568, po5569,
    po5570, po5571, po5572, po5573, po5574, po5575, po5576, po5577, po5578,
    po5579, po5580, po5581, po5582, po5583, po5584, po5585, po5586, po5587,
    po5588, po5589, po5590, po5591, po5592, po5593, po5594, po5595, po5596,
    po5597, po5598, po5599, po5600, po5601, po5602, po5603, po5604, po5605,
    po5606, po5607, po5608, po5609, po5610, po5611, po5612, po5613, po5614,
    po5615, po5616, po5617, po5618, po5619, po5620, po5621, po5622, po5623,
    po5624, po5625, po5626, po5627, po5628, po5629, po5630, po5631, po5632,
    po5633, po5634, po5635, po5636, po5637, po5638, po5639, po5640, po5641,
    po5642, po5643, po5644, po5645, po5646, po5647, po5648, po5649, po5650,
    po5651, po5652, po5653, po5654, po5655, po5656, po5657, po5658, po5659,
    po5660, po5661, po5662, po5663, po5664, po5665, po5666, po5667, po5668,
    po5669, po5670, po5671, po5672, po5673, po5674, po5675, po5676, po5677,
    po5678, po5679, po5680, po5681, po5682, po5683, po5684, po5685, po5686,
    po5687, po5688, po5689, po5690, po5691, po5692, po5693, po5694, po5695,
    po5696, po5697, po5698, po5699, po5700, po5701, po5702, po5703, po5704,
    po5705, po5706, po5707, po5708, po5709, po5710, po5711, po5712, po5713,
    po5714, po5715, po5716, po5717, po5718, po5719, po5720, po5721, po5722,
    po5723, po5724, po5725, po5726, po5727, po5728, po5729, po5730, po5731,
    po5732, po5733, po5734, po5735, po5736, po5737, po5738, po5739, po5740,
    po5741, po5742, po5743, po5744, po5745, po5746, po5747, po5748, po5749,
    po5750, po5751, po5752, po5753, po5754, po5755, po5756, po5757, po5758,
    po5759, po5760, po5761, po5762, po5763, po5764, po5765, po5766, po5767,
    po5768, po5769, po5770, po5771, po5772, po5773, po5774, po5775, po5776,
    po5777, po5778, po5779, po5780, po5781, po5782, po5783, po5784, po5785,
    po5786, po5787, po5788, po5789, po5790, po5791, po5792, po5793, po5794,
    po5795, po5796, po5797, po5798, po5799, po5800, po5801, po5802, po5803,
    po5804, po5805, po5806, po5807, po5808, po5809, po5810, po5811, po5812,
    po5813, po5814, po5815, po5816, po5817, po5818, po5819, po5820, po5821,
    po5822, po5823, po5824, po5825, po5826, po5827, po5828, po5829, po5830,
    po5831, po5832, po5833, po5834, po5835, po5836, po5837, po5838, po5839,
    po5840, po5841, po5842, po5843, po5844, po5845, po5846, po5847, po5848,
    po5849, po5850, po5851, po5852, po5853, po5854, po5855, po5856, po5857,
    po5858, po5859, po5860, po5861, po5862, po5863, po5864, po5865, po5866,
    po5867, po5868, po5869, po5870, po5871, po5872, po5873, po5874, po5875,
    po5876, po5877, po5878, po5879, po5880, po5881, po5882, po5883, po5884,
    po5885, po5886, po5887, po5888, po5889, po5890, po5891, po5892, po5893,
    po5894, po5895, po5896, po5897, po5898, po5899, po5900, po5901, po5902,
    po5903, po5904, po5905, po5906, po5907, po5908, po5909, po5910, po5911,
    po5912, po5913, po5914, po5915, po5916, po5917, po5918, po5919, po5920,
    po5921, po5922, po5923, po5924, po5925, po5926, po5927, po5928, po5929,
    po5930, po5931, po5932, po5933, po5934, po5935, po5936, po5937, po5938,
    po5939, po5940, po5941, po5942, po5943, po5944, po5945, po5946, po5947,
    po5948, po5949, po5950, po5951, po5952, po5953, po5954, po5955, po5956,
    po5957, po5958, po5959, po5960, po5961, po5962, po5963, po5964, po5965,
    po5966, po5967, po5968, po5969, po5970, po5971, po5972, po5973, po5974,
    po5975, po5976, po5977, po5978, po5979, po5980, po5981, po5982, po5983,
    po5984, po5985, po5986, po5987, po5988, po5989, po5990, po5991, po5992,
    po5993, po5994, po5995, po5996, po5997, po5998, po5999, po6000, po6001,
    po6002, po6003, po6004, po6005, po6006, po6007, po6008, po6009, po6010,
    po6011, po6012, po6013, po6014, po6015, po6016, po6017, po6018, po6019,
    po6020, po6021, po6022, po6023, po6024, po6025, po6026, po6027, po6028,
    po6029, po6030, po6031, po6032, po6033, po6034, po6035, po6036, po6037,
    po6038, po6039, po6040, po6041, po6042, po6043, po6044, po6045, po6046,
    po6047, po6048, po6049, po6050, po6051, po6052, po6053, po6054, po6055,
    po6056, po6057, po6058, po6059, po6060, po6061, po6062, po6063, po6064,
    po6065, po6066, po6067, po6068, po6069, po6070, po6071, po6072, po6073,
    po6074, po6075, po6076, po6077, po6078, po6079, po6080, po6081, po6082,
    po6083, po6084, po6085, po6086, po6087, po6088, po6089, po6090, po6091,
    po6092, po6093, po6094, po6095, po6096, po6097, po6098, po6099, po6100,
    po6101, po6102, po6103, po6104, po6105, po6106, po6107, po6108, po6109,
    po6110, po6111, po6112, po6113, po6114, po6115, po6116, po6117, po6118,
    po6119, po6120, po6121, po6122, po6123, po6124, po6125, po6126, po6127,
    po6128, po6129, po6130, po6131, po6132, po6133, po6134, po6135, po6136,
    po6137, po6138, po6139, po6140, po6141, po6142, po6143, po6144, po6145,
    po6146, po6147, po6148, po6149, po6150, po6151, po6152, po6153, po6154,
    po6155, po6156, po6157, po6158, po6159, po6160, po6161, po6162, po6163,
    po6164, po6165, po6166, po6167, po6168, po6169, po6170, po6171, po6172,
    po6173, po6174, po6175, po6176, po6177, po6178, po6179, po6180, po6181,
    po6182, po6183, po6184, po6185, po6186, po6187, po6188, po6189, po6190,
    po6191, po6192, po6193, po6194, po6195, po6196, po6197, po6198, po6199,
    po6200, po6201, po6202, po6203, po6204, po6205, po6206, po6207, po6208,
    po6209, po6210, po6211, po6212, po6213, po6214, po6215, po6216, po6217,
    po6218, po6219, po6220, po6221, po6222, po6223, po6224, po6225, po6226,
    po6227, po6228, po6229, po6230, po6231, po6232, po6233, po6234, po6235,
    po6236, po6237, po6238, po6239, po6240, po6241, po6242, po6243, po6244,
    po6245, po6246, po6247, po6248, po6249, po6250, po6251, po6252, po6253,
    po6254, po6255, po6256, po6257, po6258, po6259, po6260, po6261, po6262,
    po6263, po6264, po6265, po6266, po6267, po6268, po6269, po6270, po6271,
    po6272, po6273, po6274, po6275, po6276, po6277, po6278, po6279, po6280,
    po6281, po6282, po6283, po6284, po6285, po6286, po6287, po6288, po6289,
    po6290, po6291, po6292, po6293, po6294, po6295, po6296, po6297, po6298,
    po6299, po6300, po6301, po6302, po6303, po6304, po6305, po6306, po6307,
    po6308, po6309, po6310, po6311, po6312, po6313, po6314, po6315, po6316,
    po6317, po6318, po6319, po6320, po6321, po6322, po6323, po6324, po6325,
    po6326, po6327, po6328, po6329, po6330, po6331, po6332, po6333, po6334,
    po6335, po6336, po6337, po6338, po6339, po6340, po6341, po6342, po6343,
    po6344, po6345, po6346, po6347, po6348, po6349, po6350, po6351, po6352,
    po6353, po6354, po6355, po6356, po6357, po6358, po6359, po6360, po6361,
    po6362, po6363, po6364, po6365, po6366, po6367, po6368, po6369, po6370,
    po6371, po6372, po6373, po6374, po6375, po6376, po6377, po6378, po6379,
    po6380, po6381, po6382, po6383, po6384, po6385, po6386, po6387, po6388,
    po6389, po6390, po6391, po6392, po6393, po6394, po6395, po6396, po6397,
    po6398, po6399, po6400, po6401, po6402, po6403, po6404, po6405, po6406,
    po6407, po6408, po6409, po6410, po6411, po6412, po6413, po6414, po6415,
    po6416, po6417, po6418, po6419, po6420, po6421, po6422, po6423, po6424,
    po6425, po6426, po6427, po6428, po6429, po6430, po6431, po6432, po6433,
    po6434, po6435, po6436, po6437, po6438, po6439, po6440, po6441, po6442,
    po6443, po6444, po6445, po6446, po6447, po6448, po6449, po6450, po6451,
    po6452, po6453, po6454, po6455, po6456, po6457, po6458, po6459, po6460,
    po6461, po6462, po6463, po6464, po6465, po6466, po6467, po6468, po6469,
    po6470, po6471, po6472, po6473, po6474, po6475, po6476, po6477, po6478,
    po6479, po6480, po6481, po6482, po6483, po6484, po6485, po6486, po6487,
    po6488, po6489, po6490, po6491, po6492, po6493, po6494, po6495, po6496,
    po6497, po6498, po6499, po6500, po6501, po6502, po6503, po6504, po6505,
    po6506, po6507, po6508, po6509, po6510, po6511, po6512, po6513, po6514,
    po6515, po6516, po6517, po6518, po6519, po6520, po6521, po6522, po6523,
    po6524, po6525, po6526, po6527, po6528, po6529, po6530, po6531, po6532,
    po6533, po6534, po6535, po6536, po6537, po6538, po6539, po6540, po6541,
    po6542, po6543, po6544, po6545, po6546, po6547, po6548, po6549, po6550,
    po6551, po6552, po6553, po6554, po6555, po6556, po6557, po6558, po6559,
    po6560, po6561, po6562, po6563, po6564, po6565, po6566, po6567, po6568,
    po6569, po6570, po6571, po6572, po6573, po6574, po6575, po6576, po6577,
    po6578, po6579, po6580, po6581, po6582, po6583, po6584, po6585, po6586,
    po6587, po6588, po6589, po6590, po6591, po6592, po6593, po6594, po6595,
    po6596, po6597, po6598, po6599, po6600, po6601, po6602, po6603, po6604,
    po6605, po6606, po6607, po6608, po6609, po6610, po6611, po6612, po6613,
    po6614, po6615, po6616, po6617, po6618, po6619, po6620, po6621, po6622,
    po6623, po6624, po6625, po6626, po6627, po6628, po6629, po6630, po6631,
    po6632, po6633, po6634, po6635, po6636, po6637, po6638, po6639, po6640,
    po6641, po6642, po6643, po6644, po6645, po6646, po6647, po6648, po6649,
    po6650, po6651, po6652, po6653, po6654, po6655, po6656, po6657, po6658,
    po6659, po6660, po6661, po6662, po6663, po6664, po6665, po6666, po6667,
    po6668, po6669, po6670, po6671, po6672, po6673, po6674, po6675, po6676,
    po6677, po6678, po6679, po6680, po6681, po6682, po6683, po6684, po6685,
    po6686, po6687, po6688, po6689, po6690, po6691, po6692, po6693, po6694,
    po6695, po6696, po6697, po6698, po6699, po6700, po6701, po6702, po6703,
    po6704, po6705, po6706, po6707, po6708, po6709, po6710, po6711, po6712,
    po6713, po6714, po6715, po6716, po6717, po6718, po6719, po6720, po6721,
    po6722, po6723, po6724, po6725, po6726, po6727, po6728, po6729, po6730,
    po6731, po6732, po6733, po6734, po6735, po6736, po6737, po6738, po6739,
    po6740, po6741, po6742, po6743, po6744, po6745, po6746, po6747, po6748,
    po6749, po6750, po6751, po6752, po6753, po6754, po6755, po6756, po6757,
    po6758, po6759, po6760, po6761, po6762, po6763, po6764, po6765, po6766,
    po6767, po6768, po6769, po6770, po6771, po6772, po6773, po6774, po6775,
    po6776, po6777, po6778, po6779, po6780, po6781, po6782, po6783, po6784,
    po6785, po6786, po6787, po6788, po6789, po6790, po6791, po6792, po6793,
    po6794, po6795, po6796, po6797, po6798, po6799, po6800, po6801, po6802,
    po6803, po6804, po6805, po6806, po6807, po6808, po6809, po6810, po6811,
    po6812, po6813, po6814, po6815, po6816, po6817, po6818, po6819, po6820,
    po6821, po6822, po6823, po6824, po6825, po6826, po6827, po6828, po6829,
    po6830, po6831, po6832, po6833, po6834, po6835, po6836, po6837, po6838,
    po6839, po6840, po6841, po6842, po6843, po6844, po6845, po6846, po6847,
    po6848, po6849, po6850, po6851, po6852, po6853, po6854, po6855, po6856,
    po6857, po6858, po6859, po6860, po6861, po6862, po6863, po6864, po6865,
    po6866, po6867, po6868, po6869, po6870, po6871, po6872, po6873, po6874,
    po6875, po6876, po6877, po6878, po6879, po6880, po6881, po6882, po6883,
    po6884, po6885, po6886, po6887, po6888, po6889, po6890, po6891, po6892,
    po6893, po6894, po6895, po6896, po6897, po6898, po6899, po6900, po6901,
    po6902, po6903, po6904, po6905, po6906, po6907, po6908, po6909, po6910,
    po6911, po6912, po6913, po6914, po6915, po6916, po6917, po6918, po6919,
    po6920, po6921, po6922, po6923, po6924, po6925, po6926, po6927, po6928,
    po6929, po6930, po6931, po6932, po6933, po6934, po6935, po6936, po6937,
    po6938, po6939, po6940, po6941, po6942, po6943, po6944, po6945, po6946,
    po6947, po6948, po6949, po6950, po6951, po6952, po6953, po6954, po6955,
    po6956, po6957, po6958, po6959, po6960, po6961, po6962, po6963, po6964,
    po6965, po6966, po6967, po6968, po6969, po6970, po6971, po6972, po6973,
    po6974, po6975, po6976, po6977, po6978, po6979, po6980, po6981, po6982,
    po6983, po6984, po6985, po6986, po6987, po6988, po6989, po6990, po6991,
    po6992, po6993, po6994, po6995, po6996, po6997, po6998, po6999, po7000,
    po7001, po7002, po7003, po7004, po7005, po7006, po7007, po7008, po7009,
    po7010, po7011, po7012, po7013, po7014, po7015, po7016, po7017, po7018,
    po7019, po7020, po7021, po7022, po7023, po7024, po7025, po7026, po7027,
    po7028, po7029, po7030, po7031, po7032, po7033, po7034, po7035, po7036,
    po7037, po7038, po7039, po7040, po7041, po7042, po7043, po7044, po7045,
    po7046, po7047, po7048, po7049, po7050, po7051, po7052, po7053, po7054,
    po7055, po7056, po7057, po7058, po7059, po7060, po7061, po7062, po7063,
    po7064, po7065, po7066, po7067, po7068, po7069, po7070, po7071, po7072,
    po7073, po7074, po7075, po7076, po7077, po7078, po7079, po7080, po7081,
    po7082, po7083, po7084, po7085, po7086, po7087, po7088, po7089, po7090,
    po7091, po7092, po7093, po7094, po7095, po7096, po7097, po7098, po7099,
    po7100, po7101, po7102, po7103, po7104, po7105, po7106, po7107, po7108,
    po7109, po7110, po7111, po7112, po7113, po7114, po7115, po7116, po7117,
    po7118, po7119, po7120, po7121, po7122, po7123, po7124, po7125, po7126,
    po7127, po7128, po7129, po7130, po7131, po7132, po7133, po7134, po7135,
    po7136, po7137, po7138, po7139, po7140, po7141, po7142, po7143, po7144,
    po7145, po7146, po7147, po7148, po7149, po7150, po7151, po7152, po7153,
    po7154, po7155, po7156, po7157, po7158, po7159, po7160, po7161, po7162,
    po7163, po7164, po7165, po7166, po7167, po7168, po7169, po7170, po7171,
    po7172, po7173, po7174, po7175, po7176, po7177, po7178, po7179, po7180,
    po7181, po7182, po7183, po7184, po7185, po7186, po7187, po7188, po7189,
    po7190, po7191, po7192, po7193, po7194, po7195, po7196, po7197, po7198,
    po7199, po7200, po7201, po7202, po7203, po7204, po7205, po7206, po7207,
    po7208, po7209, po7210, po7211, po7212, po7213, po7214, po7215, po7216,
    po7217, po7218, po7219, po7220, po7221, po7222, po7223, po7224, po7225,
    po7226, po7227, po7228, po7229, po7230, po7231, po7232, po7233, po7234,
    po7235, po7236, po7237, po7238, po7239, po7240, po7241, po7242, po7243,
    po7244, po7245, po7246, po7247, po7248, po7249, po7250, po7251, po7252,
    po7253, po7254, po7255, po7256, po7257, po7258, po7259, po7260, po7261,
    po7262, po7263, po7264, po7265, po7266, po7267, po7268, po7269, po7270,
    po7271, po7272, po7273, po7274, po7275, po7276, po7277, po7278, po7279,
    po7280, po7281, po7282, po7283, po7284, po7285, po7286, po7287, po7288,
    po7289, po7290, po7291, po7292, po7293, po7294, po7295, po7296, po7297,
    po7298, po7299, po7300, po7301, po7302, po7303, po7304, po7305, po7306,
    po7307, po7308, po7309, po7310, po7311, po7312, po7313, po7314, po7315,
    po7316, po7317, po7318, po7319, po7320, po7321, po7322, po7323, po7324,
    po7325, po7326, po7327, po7328, po7329, po7330, po7331, po7332, po7333,
    po7334, po7335, po7336, po7337, po7338, po7339, po7340, po7341, po7342,
    po7343, po7344, po7345, po7346, po7347, po7348, po7349, po7350, po7351,
    po7352, po7353, po7354, po7355, po7356, po7357, po7358, po7359, po7360,
    po7361, po7362, po7363, po7364, po7365, po7366, po7367, po7368, po7369,
    po7370, po7371, po7372, po7373, po7374, po7375, po7376, po7377, po7378,
    po7379, po7380, po7381, po7382, po7383, po7384, po7385, po7386, po7387,
    po7388, po7389, po7390, po7391, po7392, po7393, po7394, po7395, po7396,
    po7397, po7398, po7399, po7400, po7401, po7402, po7403, po7404, po7405,
    po7406, po7407, po7408, po7409, po7410, po7411, po7412, po7413, po7414,
    po7415, po7416, po7417, po7418, po7419, po7420, po7421, po7422, po7423,
    po7424, po7425, po7426, po7427, po7428, po7429, po7430, po7431, po7432,
    po7433, po7434, po7435, po7436, po7437, po7438, po7439, po7440, po7441,
    po7442, po7443, po7444, po7445, po7446, po7447, po7448, po7449, po7450,
    po7451, po7452, po7453, po7454, po7455, po7456, po7457, po7458, po7459,
    po7460, po7461, po7462, po7463, po7464, po7465, po7466, po7467, po7468,
    po7469, po7470, po7471, po7472, po7473, po7474, po7475, po7476, po7477,
    po7478, po7479, po7480, po7481, po7482, po7483, po7484, po7485, po7486,
    po7487, po7488, po7489, po7490, po7491, po7492, po7493, po7494, po7495,
    po7496, po7497, po7498, po7499, po7500, po7501, po7502, po7503, po7504,
    po7505, po7506, po7507, po7508, po7509, po7510, po7511, po7512, po7513,
    po7514, po7515, po7516, po7517, po7518, po7519, po7520, po7521, po7522,
    po7523, po7524, po7525, po7526, po7527, po7528, po7529, po7530, po7531,
    po7532, po7533, po7534, po7535, po7536, po7537, po7538, po7539, po7540,
    po7541, po7542, po7543, po7544, po7545, po7546, po7547, po7548, po7549,
    po7550, po7551, po7552, po7553, po7554, po7555, po7556, po7557, po7558,
    po7559, po7560, po7561, po7562, po7563, po7564, po7565, po7566, po7567,
    po7568, po7569, po7570, po7571, po7572, po7573, po7574, po7575, po7576,
    po7577, po7578, po7579, po7580, po7581, po7582, po7583, po7584, po7585,
    po7586, po7587, po7588, po7589, po7590, po7591, po7592, po7593, po7594,
    po7595, po7596, po7597, po7598, po7599, po7600, po7601, po7602, po7603,
    po7604, po7605, po7606, po7607, po7608, po7609, po7610, po7611, po7612,
    po7613, po7614, po7615, po7616, po7617, po7618, po7619, po7620, po7621,
    po7622, po7623, po7624, po7625, po7626, po7627, po7628, po7629, po7630,
    po7631, po7632, po7633, po7634, po7635, po7636, po7637, po7638, po7639,
    po7640, po7641, po7642, po7643, po7644, po7645, po7646, po7647, po7648,
    po7649, po7650, po7651, po7652, po7653, po7654, po7655, po7656, po7657,
    po7658, po7659, po7660, po7661, po7662, po7663, po7664, po7665, po7666,
    po7667, po7668, po7669, po7670, po7671, po7672, po7673, po7674, po7675,
    po7676, po7677, po7678, po7679, po7680, po7681, po7682, po7683, po7684,
    po7685, po7686, po7687, po7688, po7689, po7690, po7691, po7692, po7693,
    po7694, po7695, po7696, po7697, po7698, po7699, po7700, po7701, po7702,
    po7703, po7704, po7705, po7706, po7707, po7708, po7709, po7710, po7711,
    po7712, po7713, po7714, po7715, po7716, po7717, po7718, po7719, po7720,
    po7721, po7722, po7723, po7724, po7725, po7726, po7727, po7728, po7729,
    po7730, po7731, po7732, po7733, po7734, po7735, po7736, po7737, po7738,
    po7739, po7740, po7741, po7742, po7743, po7744, po7745, po7746, po7747,
    po7748, po7749, po7750, po7751, po7752, po7753, po7754, po7755, po7756,
    po7757, po7758, po7759, po7760, po7761, po7762, po7763, po7764, po7765,
    po7766, po7767, po7768, po7769, po7770, po7771, po7772, po7773, po7774,
    po7775, po7776, po7777, po7778, po7779, po7780, po7781, po7782, po7783,
    po7784, po7785, po7786, po7787, po7788, po7789, po7790, po7791, po7792,
    po7793, po7794, po7795, po7796, po7797, po7798, po7799, po7800, po7801,
    po7802, po7803, po7804, po7805, po7806, po7807, po7808, po7809, po7810,
    po7811, po7812, po7813, po7814, po7815, po7816, po7817, po7818, po7819,
    po7820, po7821, po7822, po7823, po7824, po7825, po7826, po7827, po7828,
    po7829, po7830, po7831, po7832, po7833, po7834, po7835, po7836, po7837,
    po7838, po7839, po7840, po7841, po7842, po7843, po7844, po7845, po7846,
    po7847, po7848, po7849, po7850, po7851, po7852, po7853, po7854, po7855,
    po7856, po7857, po7858, po7859, po7860, po7861, po7862, po7863, po7864,
    po7865, po7866, po7867, po7868, po7869, po7870, po7871, po7872, po7873,
    po7874, po7875, po7876, po7877, po7878, po7879, po7880, po7881, po7882,
    po7883, po7884, po7885, po7886, po7887, po7888, po7889, po7890, po7891,
    po7892, po7893, po7894, po7895, po7896, po7897, po7898, po7899, po7900,
    po7901, po7902, po7903, po7904, po7905, po7906, po7907, po7908, po7909,
    po7910, po7911, po7912, po7913, po7914, po7915, po7916, po7917, po7918,
    po7919, po7920, po7921, po7922, po7923, po7924, po7925, po7926, po7927,
    po7928, po7929, po7930, po7931, po7932, po7933, po7934, po7935, po7936,
    po7937, po7938, po7939, po7940, po7941, po7942, po7943, po7944, po7945,
    po7946, po7947, po7948, po7949, po7950, po7951, po7952, po7953, po7954,
    po7955, po7956, po7957, po7958, po7959, po7960, po7961, po7962, po7963,
    po7964, po7965, po7966, po7967, po7968, po7969, po7970, po7971, po7972,
    po7973, po7974, po7975, po7976, po7977, po7978, po7979, po7980, po7981,
    po7982, po7983, po7984, po7985, po7986, po7987, po7988, po7989, po7990,
    po7991, po7992, po7993, po7994, po7995, po7996, po7997, po7998, po7999,
    po8000, po8001, po8002, po8003, po8004, po8005, po8006, po8007, po8008,
    po8009, po8010, po8011, po8012, po8013, po8014, po8015, po8016, po8017,
    po8018, po8019, po8020, po8021, po8022, po8023, po8024, po8025, po8026,
    po8027, po8028, po8029, po8030, po8031, po8032, po8033, po8034, po8035,
    po8036, po8037, po8038, po8039, po8040, po8041, po8042, po8043, po8044,
    po8045, po8046, po8047, po8048, po8049, po8050, po8051, po8052, po8053,
    po8054, po8055, po8056, po8057, po8058, po8059, po8060, po8061, po8062,
    po8063, po8064, po8065, po8066, po8067, po8068, po8069, po8070, po8071,
    po8072, po8073, po8074, po8075, po8076, po8077, po8078, po8079, po8080,
    po8081, po8082, po8083, po8084, po8085, po8086, po8087, po8088, po8089,
    po8090, po8091, po8092, po8093, po8094, po8095, po8096, po8097, po8098,
    po8099, po8100, po8101, po8102, po8103, po8104, po8105, po8106, po8107,
    po8108, po8109, po8110, po8111, po8112, po8113, po8114, po8115, po8116,
    po8117, po8118, po8119, po8120, po8121, po8122, po8123, po8124, po8125,
    po8126, po8127, po8128, po8129, po8130, po8131, po8132, po8133, po8134,
    po8135, po8136, po8137, po8138, po8139, po8140, po8141, po8142, po8143,
    po8144, po8145, po8146, po8147, po8148, po8149, po8150, po8151, po8152,
    po8153, po8154, po8155, po8156, po8157, po8158, po8159, po8160, po8161,
    po8162, po8163, po8164, po8165, po8166, po8167, po8168, po8169, po8170,
    po8171, po8172, po8173, po8174, po8175, po8176, po8177, po8178, po8179,
    po8180, po8181, po8182, po8183, po8184, po8185, po8186, po8187, po8188,
    po8189, po8190, po8191, po8192, po8193, po8194, po8195, po8196, po8197,
    po8198, po8199, po8200, po8201, po8202, po8203, po8204, po8205, po8206,
    po8207, po8208, po8209, po8210, po8211, po8212, po8213, po8214, po8215,
    po8216, po8217, po8218, po8219, po8220, po8221, po8222, po8223, po8224,
    po8225, po8226, po8227, po8228, po8229, po8230, po8231, po8232, po8233,
    po8234, po8235, po8236, po8237, po8238, po8239, po8240, po8241, po8242,
    po8243, po8244, po8245, po8246, po8247, po8248, po8249, po8250, po8251,
    po8252, po8253, po8254, po8255, po8256, po8257, po8258, po8259, po8260,
    po8261, po8262, po8263, po8264, po8265, po8266, po8267, po8268, po8269,
    po8270, po8271, po8272, po8273, po8274, po8275, po8276, po8277, po8278,
    po8279, po8280, po8281, po8282, po8283, po8284, po8285, po8286, po8287,
    po8288, po8289, po8290, po8291, po8292, po8293, po8294, po8295, po8296,
    po8297, po8298, po8299, po8300, po8301, po8302, po8303, po8304, po8305,
    po8306, po8307, po8308, po8309, po8310, po8311, po8312, po8313, po8314,
    po8315, po8316, po8317, po8318, po8319, po8320, po8321, po8322, po8323,
    po8324, po8325, po8326, po8327, po8328, po8329, po8330, po8331, po8332,
    po8333, po8334, po8335, po8336, po8337, po8338, po8339, po8340, po8341,
    po8342, po8343, po8344, po8345, po8346, po8347, po8348, po8349, po8350,
    po8351, po8352, po8353, po8354, po8355, po8356, po8357, po8358, po8359,
    po8360, po8361, po8362, po8363, po8364, po8365, po8366, po8367, po8368,
    po8369, po8370, po8371, po8372, po8373, po8374, po8375, po8376, po8377,
    po8378, po8379, po8380, po8381, po8382, po8383, po8384, po8385, po8386,
    po8387, po8388, po8389, po8390, po8391, po8392, po8393, po8394, po8395,
    po8396, po8397, po8398, po8399, po8400, po8401, po8402, po8403, po8404,
    po8405, po8406, po8407, po8408, po8409, po8410, po8411, po8412, po8413,
    po8414, po8415, po8416, po8417, po8418, po8419, po8420, po8421, po8422,
    po8423, po8424, po8425, po8426, po8427, po8428, po8429, po8430, po8431,
    po8432, po8433, po8434, po8435, po8436, po8437, po8438, po8439, po8440,
    po8441, po8442, po8443, po8444, po8445, po8446, po8447, po8448, po8449,
    po8450, po8451, po8452, po8453, po8454, po8455, po8456, po8457, po8458,
    po8459, po8460, po8461, po8462, po8463, po8464, po8465, po8466, po8467,
    po8468, po8469, po8470, po8471, po8472, po8473, po8474, po8475, po8476,
    po8477, po8478, po8479, po8480, po8481, po8482, po8483, po8484, po8485,
    po8486, po8487, po8488, po8489, po8490, po8491, po8492, po8493, po8494,
    po8495, po8496, po8497, po8498, po8499, po8500, po8501, po8502, po8503,
    po8504, po8505, po8506, po8507, po8508, po8509, po8510, po8511, po8512,
    po8513, po8514, po8515, po8516, po8517, po8518, po8519, po8520, po8521,
    po8522, po8523, po8524, po8525, po8526, po8527, po8528, po8529, po8530,
    po8531, po8532, po8533, po8534, po8535, po8536, po8537, po8538, po8539,
    po8540, po8541, po8542, po8543, po8544, po8545, po8546, po8547, po8548,
    po8549, po8550, po8551, po8552, po8553, po8554, po8555, po8556, po8557,
    po8558, po8559, po8560, po8561, po8562, po8563, po8564, po8565, po8566,
    po8567, po8568, po8569, po8570, po8571, po8572, po8573, po8574, po8575,
    po8576, po8577, po8578, po8579, po8580, po8581, po8582, po8583, po8584,
    po8585, po8586, po8587, po8588, po8589, po8590, po8591, po8592, po8593,
    po8594, po8595, po8596, po8597, po8598, po8599, po8600, po8601, po8602,
    po8603, po8604, po8605, po8606, po8607, po8608, po8609, po8610, po8611,
    po8612, po8613, po8614, po8615, po8616, po8617, po8618, po8619, po8620,
    po8621, po8622, po8623, po8624, po8625, po8626, po8627, po8628, po8629,
    po8630, po8631, po8632, po8633, po8634, po8635, po8636, po8637, po8638,
    po8639, po8640, po8641, po8642, po8643, po8644, po8645, po8646, po8647,
    po8648, po8649, po8650, po8651, po8652, po8653, po8654, po8655, po8656,
    po8657, po8658, po8659, po8660, po8661, po8662, po8663, po8664, po8665,
    po8666, po8667, po8668, po8669, po8670, po8671, po8672, po8673, po8674,
    po8675, po8676, po8677, po8678, po8679, po8680, po8681, po8682, po8683,
    po8684, po8685, po8686, po8687, po8688, po8689, po8690, po8691, po8692,
    po8693, po8694, po8695, po8696, po8697, po8698, po8699, po8700, po8701,
    po8702, po8703, po8704, po8705, po8706, po8707, po8708, po8709, po8710,
    po8711, po8712, po8713, po8714, po8715, po8716, po8717, po8718, po8719,
    po8720, po8721, po8722, po8723, po8724, po8725, po8726, po8727, po8728,
    po8729, po8730, po8731, po8732, po8733, po8734, po8735, po8736, po8737,
    po8738, po8739, po8740, po8741, po8742, po8743, po8744, po8745, po8746,
    po8747, po8748, po8749, po8750, po8751, po8752, po8753, po8754, po8755,
    po8756, po8757, po8758, po8759, po8760, po8761, po8762, po8763, po8764,
    po8765, po8766, po8767, po8768, po8769, po8770, po8771, po8772, po8773,
    po8774, po8775, po8776, po8777, po8778, po8779, po8780, po8781, po8782,
    po8783, po8784, po8785, po8786, po8787, po8788, po8789, po8790, po8791,
    po8792, po8793, po8794, po8795, po8796, po8797, po8798, po8799, po8800,
    po8801, po8802, po8803, po8804, po8805, po8806, po8807, po8808, po8809,
    po8810, po8811, po8812, po8813, po8814, po8815, po8816, po8817, po8818,
    po8819, po8820, po8821, po8822, po8823, po8824, po8825, po8826, po8827,
    po8828, po8829, po8830, po8831, po8832, po8833, po8834, po8835, po8836,
    po8837, po8838, po8839, po8840, po8841, po8842, po8843, po8844, po8845,
    po8846, po8847, po8848, po8849, po8850, po8851, po8852, po8853, po8854,
    po8855, po8856, po8857, po8858, po8859, po8860, po8861, po8862, po8863,
    po8864, po8865, po8866, po8867, po8868, po8869, po8870, po8871, po8872,
    po8873, po8874, po8875, po8876, po8877, po8878, po8879, po8880, po8881,
    po8882, po8883, po8884, po8885, po8886, po8887, po8888, po8889, po8890,
    po8891, po8892, po8893, po8894, po8895, po8896, po8897, po8898, po8899,
    po8900, po8901, po8902, po8903, po8904, po8905, po8906, po8907, po8908,
    po8909, po8910, po8911, po8912, po8913, po8914, po8915, po8916, po8917,
    po8918, po8919, po8920, po8921, po8922, po8923, po8924, po8925, po8926,
    po8927, po8928, po8929, po8930, po8931, po8932, po8933, po8934, po8935,
    po8936, po8937, po8938, po8939, po8940, po8941, po8942, po8943, po8944,
    po8945, po8946, po8947, po8948, po8949, po8950, po8951, po8952, po8953,
    po8954, po8955, po8956, po8957, po8958, po8959, po8960, po8961, po8962,
    po8963, po8964, po8965, po8966, po8967, po8968, po8969, po8970, po8971,
    po8972, po8973, po8974, po8975, po8976, po8977, po8978, po8979, po8980,
    po8981, po8982, po8983, po8984, po8985, po8986, po8987, po8988, po8989,
    po8990, po8991, po8992, po8993, po8994, po8995, po8996, po8997, po8998,
    po8999, po9000, po9001, po9002, po9003, po9004, po9005, po9006, po9007,
    po9008, po9009, po9010, po9011, po9012, po9013, po9014, po9015, po9016,
    po9017, po9018, po9019, po9020, po9021, po9022, po9023, po9024, po9025,
    po9026, po9027, po9028, po9029, po9030, po9031, po9032, po9033, po9034,
    po9035, po9036, po9037;
  wire n18082, n18083, n18084, n18085, n18086, n18087, n18088, n18089,
    n18090, n18091, n18092, n18093, n18094, n18095, n18096, n18097, n18098,
    n18099, n18100, n18101, n18102, n18103, n18104, n18105, n18106, n18107,
    n18108, n18109, n18110, n18111, n18112, n18113, n18114, n18115, n18116,
    n18117, n18118, n18119, n18120, n18121, n18122, n18123, n18124, n18125,
    n18126, n18127, n18128, n18129, n18130, n18131, n18132, n18133, n18134,
    n18135, n18136, n18137, n18138, n18139, n18140, n18141, n18142, n18143,
    n18144, n18145, n18146, n18147, n18148, n18149, n18150, n18151, n18152,
    n18153, n18154, n18155, n18156, n18157, n18158, n18159, n18160, n18161,
    n18162, n18163, n18164, n18165, n18166, n18167, n18168, n18169, n18170,
    n18171, n18172, n18173, n18174, n18175, n18176, n18177, n18178, n18179,
    n18180, n18181, n18182, n18183, n18184, n18185, n18187, n18188, n18189,
    n18190, n18191, n18192, n18193, n18194, n18195, n18196, n18197, n18198,
    n18199, n18200, n18201, n18202, n18203, n18204, n18205, n18206, n18207,
    n18208, n18209, n18210, n18211, n18212, n18213, n18214, n18215, n18216,
    n18217, n18218, n18219, n18220, n18222, n18223, n18224, n18225, n18226,
    n18227, n18228, n18229, n18230, n18231, n18232, n18233, n18234, n18235,
    n18236, n18237, n18238, n18239, n18240, n18241, n18242, n18243, n18244,
    n18245, n18246, n18247, n18248, n18249, n18250, n18251, n18252, n18253,
    n18254, n18255, n18256, n18257, n18258, n18259, n18260, n18261, n18262,
    n18263, n18264, n18265, n18266, n18267, n18268, n18269, n18270, n18271,
    n18272, n18273, n18274, n18275, n18276, n18277, n18278, n18279, n18280,
    n18281, n18282, n18283, n18284, n18285, n18286, n18287, n18288, n18289,
    n18290, n18291, n18292, n18293, n18294, n18295, n18296, n18297, n18298,
    n18299, n18300, n18301, n18302, n18303, n18304, n18305, n18306, n18307,
    n18308, n18309, n18310, n18311, n18312, n18313, n18314, n18315, n18316,
    n18317, n18318, n18319, n18321, n18322, n18323, n18324, n18325, n18326,
    n18327, n18328, n18329, n18330, n18331, n18332, n18333, n18334, n18335,
    n18336, n18337, n18338, n18339, n18340, n18341, n18342, n18343, n18344,
    n18346, n18347, n18348, n18349, n18350, n18351, n18352, n18353, n18354,
    n18355, n18356, n18357, n18358, n18359, n18360, n18361, n18362, n18363,
    n18364, n18365, n18366, n18367, n18368, n18369, n18370, n18371, n18372,
    n18373, n18374, n18375, n18376, n18377, n18378, n18379, n18380, n18381,
    n18382, n18383, n18384, n18385, n18386, n18387, n18388, n18389, n18390,
    n18391, n18392, n18393, n18394, n18395, n18396, n18397, n18398, n18399,
    n18400, n18401, n18402, n18403, n18404, n18405, n18406, n18407, n18408,
    n18409, n18410, n18411, n18412, n18413, n18414, n18415, n18416, n18417,
    n18418, n18419, n18420, n18421, n18422, n18423, n18424, n18425, n18426,
    n18427, n18428, n18429, n18430, n18431, n18432, n18433, n18434, n18435,
    n18436, n18437, n18438, n18439, n18440, n18441, n18442, n18443, n18444,
    n18446, n18447, n18448, n18449, n18450, n18451, n18452, n18453, n18454,
    n18455, n18456, n18457, n18458, n18459, n18460, n18461, n18462, n18463,
    n18464, n18465, n18466, n18467, n18468, n18469, n18470, n18471, n18472,
    n18473, n18474, n18475, n18477, n18478, n18479, n18480, n18481, n18482,
    n18483, n18484, n18485, n18486, n18487, n18488, n18489, n18490, n18491,
    n18492, n18493, n18494, n18495, n18496, n18497, n18498, n18499, n18500,
    n18501, n18502, n18503, n18504, n18505, n18506, n18507, n18509, n18510,
    n18511, n18512, n18513, n18514, n18515, n18516, n18517, n18518, n18519,
    n18520, n18521, n18522, n18523, n18524, n18525, n18526, n18527, n18528,
    n18529, n18530, n18531, n18532, n18533, n18534, n18535, n18536, n18537,
    n18538, n18539, n18540, n18541, n18542, n18543, n18544, n18545, n18546,
    n18547, n18548, n18549, n18550, n18551, n18552, n18553, n18554, n18555,
    n18556, n18557, n18558, n18559, n18560, n18561, n18562, n18563, n18564,
    n18565, n18566, n18567, n18568, n18569, n18570, n18571, n18572, n18573,
    n18574, n18575, n18576, n18577, n18578, n18579, n18580, n18581, n18582,
    n18583, n18584, n18585, n18586, n18587, n18588, n18589, n18590, n18591,
    n18592, n18593, n18594, n18595, n18596, n18597, n18598, n18599, n18601,
    n18602, n18603, n18604, n18605, n18606, n18607, n18608, n18609, n18610,
    n18611, n18612, n18613, n18614, n18615, n18616, n18617, n18618, n18619,
    n18620, n18621, n18622, n18623, n18624, n18625, n18626, n18627, n18628,
    n18629, n18630, n18631, n18632, n18633, n18634, n18635, n18636, n18637,
    n18638, n18639, n18640, n18641, n18642, n18643, n18644, n18645, n18646,
    n18647, n18648, n18649, n18650, n18651, n18652, n18653, n18654, n18655,
    n18656, n18657, n18658, n18659, n18660, n18661, n18662, n18663, n18664,
    n18665, n18666, n18667, n18668, n18669, n18670, n18671, n18672, n18673,
    n18674, n18675, n18676, n18677, n18678, n18679, n18680, n18681, n18682,
    n18683, n18684, n18685, n18686, n18687, n18688, n18689, n18690, n18691,
    n18692, n18693, n18694, n18695, n18696, n18697, n18698, n18700, n18701,
    n18702, n18703, n18704, n18705, n18706, n18707, n18708, n18709, n18710,
    n18711, n18712, n18713, n18714, n18715, n18716, n18717, n18718, n18719,
    n18720, n18721, n18722, n18723, n18724, n18725, n18726, n18727, n18728,
    n18729, n18730, n18731, n18732, n18733, n18734, n18735, n18736, n18737,
    n18738, n18739, n18740, n18741, n18742, n18743, n18744, n18745, n18746,
    n18747, n18748, n18749, n18750, n18751, n18752, n18753, n18754, n18755,
    n18756, n18757, n18758, n18759, n18760, n18761, n18762, n18763, n18764,
    n18765, n18766, n18767, n18768, n18769, n18770, n18771, n18772, n18773,
    n18774, n18775, n18776, n18777, n18778, n18779, n18780, n18781, n18782,
    n18783, n18784, n18785, n18786, n18787, n18788, n18789, n18790, n18791,
    n18792, n18793, n18794, n18795, n18796, n18797, n18798, n18800, n18801,
    n18802, n18803, n18804, n18805, n18806, n18807, n18808, n18809, n18810,
    n18811, n18812, n18813, n18814, n18815, n18816, n18817, n18818, n18819,
    n18820, n18821, n18822, n18823, n18824, n18825, n18826, n18827, n18828,
    n18829, n18830, n18831, n18832, n18833, n18834, n18835, n18836, n18837,
    n18839, n18840, n18841, n18842, n18843, n18844, n18845, n18846, n18847,
    n18848, n18849, n18850, n18851, n18852, n18853, n18854, n18855, n18856,
    n18857, n18858, n18859, n18860, n18861, n18862, n18863, n18864, n18865,
    n18866, n18867, n18868, n18869, n18870, n18872, n18873, n18874, n18875,
    n18876, n18877, n18878, n18879, n18880, n18881, n18882, n18883, n18884,
    n18885, n18886, n18887, n18888, n18889, n18890, n18891, n18892, n18893,
    n18894, n18895, n18896, n18897, n18898, n18899, n18900, n18901, n18902,
    n18903, n18904, n18905, n18906, n18907, n18908, n18909, n18910, n18911,
    n18913, n18914, n18915, n18916, n18917, n18918, n18919, n18920, n18921,
    n18922, n18923, n18924, n18925, n18926, n18927, n18928, n18929, n18930,
    n18931, n18932, n18933, n18934, n18935, n18936, n18937, n18938, n18939,
    n18940, n18941, n18942, n18943, n18944, n18945, n18946, n18947, n18948,
    n18950, n18951, n18952, n18953, n18954, n18955, n18956, n18957, n18958,
    n18959, n18960, n18961, n18962, n18963, n18964, n18965, n18966, n18967,
    n18968, n18969, n18970, n18971, n18972, n18973, n18974, n18975, n18976,
    n18977, n18978, n18979, n18980, n18981, n18982, n18983, n18984, n18986,
    n18987, n18988, n18989, n18990, n18991, n18992, n18993, n18994, n18995,
    n18996, n18997, n18998, n18999, n19000, n19001, n19002, n19003, n19004,
    n19005, n19006, n19007, n19008, n19009, n19010, n19011, n19012, n19013,
    n19014, n19015, n19016, n19017, n19019, n19020, n19021, n19022, n19023,
    n19024, n19025, n19026, n19027, n19028, n19029, n19030, n19031, n19032,
    n19033, n19034, n19035, n19036, n19037, n19038, n19039, n19040, n19041,
    n19042, n19043, n19044, n19045, n19047, n19048, n19049, n19050, n19051,
    n19052, n19053, n19054, n19055, n19056, n19057, n19058, n19059, n19060,
    n19061, n19062, n19063, n19064, n19065, n19066, n19067, n19068, n19069,
    n19070, n19071, n19072, n19073, n19074, n19076, n19077, n19078, n19079,
    n19080, n19081, n19082, n19083, n19084, n19085, n19086, n19087, n19088,
    n19089, n19090, n19091, n19092, n19093, n19094, n19095, n19096, n19097,
    n19098, n19099, n19100, n19101, n19102, n19103, n19104, n19105, n19106,
    n19107, n19108, n19110, n19111, n19112, n19113, n19114, n19115, n19116,
    n19117, n19118, n19119, n19120, n19121, n19122, n19123, n19124, n19125,
    n19126, n19127, n19128, n19129, n19130, n19131, n19132, n19133, n19134,
    n19135, n19136, n19137, n19138, n19139, n19140, n19141, n19142, n19143,
    n19144, n19145, n19146, n19147, n19148, n19149, n19150, n19151, n19152,
    n19153, n19154, n19155, n19156, n19157, n19158, n19159, n19160, n19161,
    n19162, n19163, n19164, n19165, n19166, n19167, n19168, n19169, n19170,
    n19171, n19172, n19173, n19174, n19175, n19176, n19177, n19178, n19179,
    n19180, n19181, n19182, n19183, n19184, n19185, n19186, n19187, n19188,
    n19189, n19190, n19191, n19192, n19193, n19194, n19195, n19196, n19197,
    n19198, n19199, n19200, n19201, n19202, n19203, n19205, n19206, n19207,
    n19208, n19209, n19210, n19211, n19212, n19213, n19214, n19215, n19216,
    n19217, n19218, n19219, n19220, n19221, n19222, n19223, n19224, n19225,
    n19226, n19227, n19228, n19229, n19230, n19231, n19232, n19233, n19234,
    n19235, n19236, n19237, n19238, n19240, n19241, n19242, n19243, n19244,
    n19245, n19246, n19247, n19248, n19249, n19250, n19251, n19252, n19253,
    n19254, n19255, n19256, n19257, n19258, n19259, n19260, n19261, n19262,
    n19263, n19264, n19265, n19266, n19267, n19268, n19269, n19270, n19271,
    n19272, n19273, n19274, n19276, n19277, n19278, n19279, n19280, n19281,
    n19282, n19283, n19284, n19285, n19286, n19287, n19288, n19289, n19290,
    n19291, n19292, n19293, n19294, n19295, n19296, n19297, n19298, n19299,
    n19301, n19302, n19303, n19304, n19305, n19306, n19307, n19308, n19309,
    n19310, n19311, n19312, n19313, n19314, n19315, n19316, n19317, n19318,
    n19319, n19320, n19321, n19322, n19324, n19325, n19326, n19327, n19328,
    n19329, n19330, n19331, n19332, n19333, n19334, n19335, n19336, n19337,
    n19338, n19339, n19340, n19341, n19342, n19343, n19344, n19345, n19346,
    n19347, n19348, n19349, n19350, n19351, n19352, n19353, n19354, n19355,
    n19356, n19357, n19358, n19359, n19360, n19361, n19363, n19364, n19365,
    n19366, n19367, n19368, n19369, n19370, n19371, n19372, n19373, n19374,
    n19375, n19376, n19377, n19378, n19379, n19380, n19381, n19382, n19383,
    n19384, n19385, n19386, n19387, n19388, n19389, n19390, n19391, n19392,
    n19393, n19394, n19396, n19397, n19398, n19399, n19400, n19401, n19402,
    n19403, n19404, n19405, n19406, n19407, n19408, n19409, n19410, n19411,
    n19412, n19413, n19414, n19415, n19416, n19417, n19418, n19419, n19420,
    n19421, n19422, n19423, n19424, n19425, n19427, n19428, n19429, n19430,
    n19431, n19432, n19433, n19434, n19435, n19436, n19437, n19438, n19439,
    n19440, n19441, n19442, n19443, n19444, n19445, n19446, n19447, n19448,
    n19449, n19450, n19451, n19452, n19453, n19454, n19455, n19456, n19457,
    n19458, n19459, n19460, n19461, n19462, n19463, n19464, n19465, n19466,
    n19467, n19468, n19469, n19470, n19471, n19472, n19473, n19474, n19475,
    n19476, n19477, n19478, n19479, n19480, n19481, n19482, n19483, n19484,
    n19485, n19486, n19487, n19488, n19489, n19490, n19491, n19492, n19493,
    n19494, n19495, n19496, n19497, n19498, n19499, n19500, n19501, n19502,
    n19503, n19504, n19505, n19506, n19507, n19508, n19509, n19510, n19511,
    n19512, n19513, n19514, n19515, n19516, n19517, n19518, n19519, n19521,
    n19522, n19523, n19524, n19525, n19526, n19527, n19528, n19529, n19530,
    n19531, n19532, n19533, n19534, n19535, n19536, n19537, n19538, n19539,
    n19540, n19541, n19542, n19543, n19544, n19545, n19546, n19547, n19549,
    n19550, n19551, n19552, n19553, n19554, n19555, n19556, n19557, n19558,
    n19559, n19560, n19561, n19562, n19563, n19564, n19565, n19566, n19567,
    n19568, n19569, n19570, n19571, n19572, n19573, n19574, n19575, n19576,
    n19577, n19578, n19579, n19580, n19581, n19582, n19583, n19584, n19585,
    n19586, n19588, n19589, n19590, n19591, n19592, n19593, n19594, n19595,
    n19596, n19597, n19598, n19599, n19600, n19601, n19602, n19603, n19604,
    n19605, n19606, n19607, n19608, n19609, n19610, n19611, n19612, n19613,
    n19614, n19615, n19616, n19617, n19618, n19620, n19621, n19622, n19623,
    n19624, n19625, n19626, n19627, n19628, n19629, n19630, n19631, n19632,
    n19633, n19634, n19635, n19636, n19637, n19638, n19639, n19640, n19641,
    n19642, n19643, n19644, n19645, n19647, n19648, n19649, n19650, n19651,
    n19652, n19653, n19654, n19655, n19656, n19657, n19658, n19659, n19660,
    n19661, n19662, n19663, n19664, n19665, n19666, n19667, n19668, n19669,
    n19670, n19671, n19672, n19673, n19674, n19675, n19676, n19677, n19678,
    n19679, n19680, n19681, n19682, n19683, n19684, n19685, n19686, n19687,
    n19688, n19689, n19690, n19691, n19692, n19693, n19694, n19695, n19696,
    n19697, n19698, n19699, n19700, n19701, n19702, n19703, n19704, n19705,
    n19706, n19707, n19708, n19709, n19710, n19711, n19712, n19713, n19714,
    n19715, n19716, n19717, n19718, n19719, n19720, n19721, n19722, n19723,
    n19724, n19725, n19726, n19727, n19728, n19729, n19730, n19731, n19732,
    n19733, n19734, n19735, n19736, n19737, n19738, n19739, n19740, n19741,
    n19742, n19743, n19744, n19745, n19746, n19748, n19749, n19750, n19751,
    n19752, n19753, n19754, n19755, n19756, n19757, n19758, n19759, n19760,
    n19761, n19762, n19763, n19764, n19765, n19766, n19767, n19768, n19769,
    n19770, n19771, n19772, n19773, n19774, n19775, n19776, n19777, n19778,
    n19779, n19780, n19781, n19782, n19783, n19784, n19785, n19786, n19787,
    n19788, n19789, n19790, n19791, n19792, n19793, n19794, n19795, n19796,
    n19797, n19798, n19799, n19800, n19801, n19802, n19803, n19804, n19805,
    n19806, n19807, n19808, n19809, n19810, n19811, n19812, n19813, n19814,
    n19815, n19816, n19817, n19818, n19819, n19820, n19821, n19822, n19823,
    n19824, n19825, n19826, n19827, n19828, n19829, n19830, n19831, n19832,
    n19833, n19834, n19835, n19836, n19837, n19838, n19840, n19841, n19842,
    n19843, n19844, n19845, n19846, n19847, n19848, n19849, n19850, n19851,
    n19852, n19853, n19854, n19855, n19856, n19857, n19858, n19859, n19860,
    n19861, n19862, n19863, n19864, n19865, n19866, n19867, n19868, n19869,
    n19870, n19871, n19872, n19873, n19874, n19875, n19876, n19877, n19878,
    n19879, n19880, n19881, n19882, n19883, n19884, n19885, n19886, n19887,
    n19888, n19889, n19890, n19891, n19892, n19893, n19894, n19895, n19896,
    n19897, n19898, n19899, n19900, n19901, n19902, n19903, n19904, n19905,
    n19906, n19907, n19908, n19909, n19910, n19911, n19912, n19913, n19914,
    n19915, n19916, n19917, n19918, n19919, n19920, n19921, n19922, n19923,
    n19924, n19925, n19926, n19927, n19928, n19929, n19930, n19931, n19932,
    n19933, n19934, n19935, n19936, n19937, n19938, n19940, n19941, n19942,
    n19943, n19944, n19945, n19946, n19947, n19948, n19949, n19950, n19951,
    n19952, n19953, n19954, n19955, n19956, n19957, n19958, n19959, n19960,
    n19961, n19962, n19963, n19964, n19965, n19966, n19967, n19968, n19969,
    n19970, n19971, n19972, n19973, n19974, n19975, n19976, n19977, n19978,
    n19979, n19980, n19981, n19982, n19983, n19984, n19985, n19986, n19987,
    n19988, n19989, n19990, n19991, n19993, n19994, n19995, n19996, n19997,
    n19998, n19999, n20000, n20001, n20002, n20003, n20004, n20005, n20006,
    n20007, n20008, n20009, n20010, n20011, n20012, n20013, n20014, n20015,
    n20016, n20017, n20018, n20019, n20020, n20021, n20022, n20023, n20024,
    n20025, n20026, n20027, n20028, n20029, n20030, n20031, n20032, n20034,
    n20035, n20036, n20037, n20038, n20039, n20040, n20041, n20042, n20043,
    n20044, n20045, n20046, n20047, n20048, n20049, n20050, n20051, n20052,
    n20053, n20054, n20055, n20056, n20057, n20058, n20059, n20060, n20061,
    n20062, n20063, n20064, n20065, n20066, n20067, n20068, n20069, n20070,
    n20071, n20072, n20073, n20074, n20075, n20077, n20078, n20079, n20080,
    n20081, n20082, n20083, n20084, n20085, n20086, n20087, n20088, n20089,
    n20090, n20091, n20092, n20093, n20094, n20095, n20096, n20097, n20098,
    n20099, n20100, n20101, n20102, n20103, n20104, n20105, n20106, n20107,
    n20108, n20109, n20110, n20111, n20112, n20113, n20114, n20115, n20116,
    n20117, n20118, n20119, n20120, n20121, n20122, n20123, n20124, n20125,
    n20126, n20127, n20128, n20129, n20130, n20131, n20132, n20133, n20134,
    n20135, n20136, n20137, n20138, n20139, n20140, n20141, n20142, n20143,
    n20144, n20145, n20146, n20147, n20148, n20149, n20150, n20151, n20152,
    n20153, n20154, n20155, n20156, n20157, n20158, n20159, n20160, n20161,
    n20162, n20163, n20164, n20165, n20166, n20167, n20169, n20170, n20171,
    n20172, n20173, n20174, n20175, n20176, n20177, n20178, n20179, n20180,
    n20181, n20182, n20183, n20184, n20185, n20186, n20187, n20188, n20189,
    n20190, n20191, n20192, n20193, n20194, n20195, n20196, n20197, n20198,
    n20199, n20200, n20201, n20202, n20203, n20204, n20205, n20206, n20207,
    n20208, n20209, n20210, n20211, n20212, n20213, n20215, n20216, n20217,
    n20218, n20219, n20220, n20221, n20222, n20223, n20224, n20225, n20226,
    n20227, n20228, n20229, n20230, n20231, n20232, n20233, n20234, n20235,
    n20236, n20237, n20238, n20239, n20240, n20241, n20242, n20243, n20244,
    n20245, n20246, n20248, n20249, n20250, n20251, n20252, n20253, n20254,
    n20255, n20256, n20257, n20258, n20259, n20260, n20261, n20262, n20263,
    n20264, n20265, n20266, n20267, n20268, n20269, n20270, n20271, n20272,
    n20273, n20274, n20275, n20276, n20277, n20278, n20279, n20280, n20281,
    n20282, n20283, n20285, n20286, n20287, n20288, n20289, n20290, n20291,
    n20292, n20293, n20294, n20295, n20296, n20297, n20298, n20299, n20300,
    n20301, n20302, n20303, n20304, n20305, n20306, n20307, n20308, n20309,
    n20310, n20311, n20312, n20313, n20314, n20315, n20316, n20317, n20318,
    n20319, n20320, n20321, n20322, n20323, n20324, n20325, n20326, n20327,
    n20328, n20329, n20330, n20331, n20332, n20333, n20334, n20336, n20337,
    n20338, n20339, n20340, n20341, n20342, n20343, n20344, n20345, n20346,
    n20347, n20348, n20349, n20350, n20351, n20352, n20353, n20354, n20355,
    n20356, n20357, n20358, n20359, n20360, n20361, n20362, n20363, n20364,
    n20365, n20366, n20367, n20368, n20369, n20370, n20371, n20372, n20373,
    n20374, n20375, n20376, n20377, n20378, n20379, n20380, n20381, n20382,
    n20383, n20384, n20385, n20386, n20387, n20388, n20389, n20390, n20391,
    n20392, n20393, n20394, n20395, n20396, n20397, n20398, n20399, n20400,
    n20401, n20402, n20403, n20404, n20405, n20406, n20407, n20408, n20409,
    n20410, n20411, n20412, n20413, n20414, n20415, n20416, n20417, n20418,
    n20419, n20420, n20421, n20422, n20423, n20424, n20425, n20426, n20427,
    n20428, n20429, n20430, n20431, n20432, n20433, n20434, n20435, n20436,
    n20437, n20439, n20440, n20441, n20442, n20443, n20444, n20445, n20446,
    n20447, n20448, n20449, n20450, n20451, n20452, n20453, n20454, n20455,
    n20456, n20457, n20458, n20459, n20460, n20461, n20462, n20463, n20464,
    n20465, n20466, n20467, n20468, n20469, n20470, n20471, n20472, n20474,
    n20475, n20476, n20477, n20478, n20479, n20480, n20481, n20482, n20483,
    n20484, n20485, n20486, n20487, n20488, n20489, n20490, n20491, n20492,
    n20493, n20494, n20495, n20496, n20497, n20498, n20499, n20500, n20501,
    n20502, n20503, n20504, n20505, n20506, n20507, n20508, n20509, n20510,
    n20511, n20513, n20514, n20515, n20516, n20517, n20518, n20519, n20520,
    n20521, n20522, n20523, n20524, n20525, n20526, n20527, n20528, n20529,
    n20530, n20531, n20532, n20533, n20534, n20535, n20536, n20537, n20538,
    n20539, n20540, n20541, n20542, n20543, n20544, n20545, n20546, n20548,
    n20549, n20550, n20551, n20552, n20553, n20554, n20555, n20556, n20557,
    n20558, n20559, n20560, n20561, n20562, n20563, n20564, n20565, n20566,
    n20567, n20568, n20569, n20570, n20571, n20572, n20573, n20574, n20575,
    n20576, n20577, n20578, n20579, n20580, n20581, n20582, n20583, n20584,
    n20585, n20586, n20587, n20588, n20589, n20590, n20591, n20592, n20593,
    n20594, n20595, n20596, n20597, n20598, n20599, n20600, n20601, n20602,
    n20603, n20604, n20605, n20606, n20607, n20608, n20609, n20610, n20611,
    n20612, n20613, n20614, n20615, n20616, n20617, n20618, n20619, n20620,
    n20621, n20622, n20623, n20624, n20625, n20626, n20627, n20628, n20629,
    n20630, n20631, n20632, n20633, n20634, n20635, n20636, n20637, n20638,
    n20639, n20640, n20641, n20642, n20643, n20644, n20645, n20646, n20647,
    n20648, n20649, n20650, n20651, n20652, n20654, n20655, n20656, n20657,
    n20658, n20659, n20660, n20661, n20662, n20663, n20664, n20665, n20666,
    n20667, n20668, n20669, n20670, n20671, n20672, n20673, n20674, n20675,
    n20676, n20677, n20678, n20679, n20680, n20681, n20682, n20683, n20684,
    n20685, n20686, n20687, n20688, n20689, n20690, n20691, n20692, n20693,
    n20694, n20695, n20696, n20697, n20698, n20700, n20701, n20702, n20703,
    n20704, n20705, n20706, n20707, n20708, n20709, n20710, n20711, n20712,
    n20713, n20714, n20715, n20716, n20717, n20718, n20719, n20720, n20721,
    n20722, n20723, n20724, n20725, n20726, n20727, n20728, n20729, n20730,
    n20731, n20732, n20733, n20734, n20735, n20736, n20737, n20738, n20739,
    n20740, n20741, n20742, n20743, n20744, n20745, n20746, n20747, n20748,
    n20749, n20750, n20751, n20752, n20753, n20754, n20755, n20756, n20757,
    n20758, n20759, n20760, n20761, n20762, n20763, n20764, n20765, n20766,
    n20767, n20768, n20769, n20770, n20771, n20772, n20773, n20774, n20775,
    n20776, n20777, n20778, n20779, n20780, n20781, n20782, n20783, n20784,
    n20785, n20786, n20787, n20788, n20789, n20790, n20791, n20792, n20793,
    n20794, n20795, n20796, n20797, n20799, n20800, n20801, n20802, n20803,
    n20804, n20805, n20806, n20807, n20808, n20809, n20810, n20811, n20812,
    n20813, n20814, n20815, n20816, n20817, n20818, n20819, n20820, n20821,
    n20822, n20823, n20824, n20825, n20826, n20827, n20828, n20829, n20830,
    n20831, n20832, n20833, n20834, n20835, n20836, n20838, n20839, n20840,
    n20841, n20842, n20843, n20844, n20845, n20846, n20847, n20848, n20849,
    n20850, n20851, n20852, n20853, n20854, n20855, n20856, n20857, n20858,
    n20859, n20860, n20861, n20862, n20863, n20864, n20865, n20866, n20867,
    n20868, n20869, n20870, n20871, n20872, n20873, n20874, n20875, n20876,
    n20878, n20879, n20880, n20881, n20882, n20883, n20884, n20885, n20886,
    n20887, n20888, n20889, n20890, n20891, n20892, n20893, n20894, n20895,
    n20896, n20897, n20898, n20899, n20900, n20901, n20902, n20903, n20904,
    n20905, n20906, n20907, n20908, n20909, n20910, n20911, n20912, n20913,
    n20914, n20915, n20917, n20918, n20919, n20920, n20921, n20922, n20923,
    n20924, n20925, n20926, n20927, n20928, n20929, n20930, n20931, n20932,
    n20933, n20934, n20935, n20936, n20937, n20938, n20939, n20940, n20941,
    n20942, n20943, n20944, n20946, n20947, n20948, n20949, n20950, n20951,
    n20952, n20953, n20954, n20955, n20956, n20957, n20958, n20959, n20960,
    n20961, n20962, n20963, n20964, n20965, n20966, n20967, n20968, n20969,
    n20970, n20971, n20972, n20973, n20974, n20975, n20976, n20977, n20978,
    n20979, n20980, n20981, n20982, n20983, n20984, n20985, n20987, n20988,
    n20989, n20990, n20991, n20992, n20993, n20994, n20995, n20996, n20997,
    n20998, n20999, n21000, n21001, n21002, n21003, n21004, n21005, n21006,
    n21007, n21008, n21009, n21010, n21011, n21012, n21013, n21014, n21015,
    n21016, n21017, n21018, n21019, n21020, n21021, n21022, n21023, n21024,
    n21025, n21026, n21027, n21028, n21029, n21030, n21031, n21032, n21033,
    n21034, n21035, n21036, n21037, n21038, n21039, n21040, n21041, n21042,
    n21043, n21044, n21045, n21046, n21047, n21048, n21049, n21050, n21051,
    n21052, n21053, n21054, n21055, n21056, n21057, n21058, n21059, n21060,
    n21061, n21062, n21063, n21064, n21065, n21066, n21067, n21068, n21069,
    n21070, n21071, n21072, n21073, n21074, n21075, n21076, n21077, n21078,
    n21079, n21080, n21081, n21083, n21084, n21085, n21086, n21087, n21088,
    n21089, n21090, n21091, n21092, n21093, n21094, n21095, n21096, n21097,
    n21098, n21099, n21100, n21101, n21102, n21103, n21104, n21105, n21106,
    n21107, n21108, n21109, n21110, n21111, n21112, n21114, n21115, n21116,
    n21117, n21118, n21119, n21120, n21121, n21122, n21123, n21124, n21125,
    n21126, n21127, n21128, n21129, n21130, n21131, n21132, n21133, n21134,
    n21135, n21136, n21137, n21138, n21139, n21140, n21141, n21142, n21143,
    n21144, n21145, n21146, n21147, n21148, n21149, n21150, n21151, n21152,
    n21153, n21154, n21155, n21156, n21157, n21158, n21159, n21161, n21162,
    n21163, n21164, n21165, n21166, n21167, n21168, n21169, n21170, n21171,
    n21172, n21173, n21174, n21175, n21176, n21177, n21178, n21179, n21180,
    n21181, n21182, n21183, n21184, n21185, n21186, n21187, n21188, n21189,
    n21190, n21191, n21192, n21193, n21194, n21195, n21196, n21198, n21199,
    n21200, n21201, n21202, n21203, n21204, n21205, n21206, n21207, n21208,
    n21209, n21210, n21211, n21212, n21213, n21214, n21215, n21216, n21217,
    n21218, n21219, n21220, n21221, n21222, n21223, n21224, n21225, n21226,
    n21227, n21228, n21229, n21230, n21231, n21232, n21233, n21234, n21235,
    n21236, n21237, n21238, n21239, n21240, n21241, n21242, n21244, n21245,
    n21246, n21247, n21248, n21249, n21250, n21251, n21252, n21253, n21254,
    n21255, n21256, n21257, n21258, n21259, n21260, n21261, n21262, n21263,
    n21264, n21265, n21266, n21267, n21268, n21269, n21270, n21271, n21272,
    n21273, n21274, n21275, n21276, n21277, n21279, n21280, n21281, n21282,
    n21283, n21284, n21285, n21286, n21287, n21288, n21289, n21290, n21291,
    n21292, n21293, n21294, n21295, n21296, n21297, n21298, n21299, n21300,
    n21301, n21302, n21303, n21304, n21305, n21306, n21307, n21308, n21309,
    n21310, n21312, n21313, n21314, n21315, n21316, n21317, n21318, n21319,
    n21320, n21321, n21322, n21323, n21324, n21325, n21326, n21327, n21328,
    n21329, n21330, n21331, n21332, n21333, n21334, n21335, n21336, n21337,
    n21339, n21340, n21341, n21342, n21343, n21344, n21345, n21346, n21347,
    n21348, n21349, n21350, n21351, n21352, n21353, n21354, n21355, n21356,
    n21357, n21358, n21359, n21360, n21361, n21362, n21363, n21364, n21365,
    n21366, n21367, n21369, n21370, n21371, n21372, n21373, n21374, n21375,
    n21376, n21377, n21378, n21379, n21380, n21381, n21382, n21383, n21384,
    n21385, n21386, n21387, n21388, n21389, n21390, n21391, n21392, n21393,
    n21394, n21395, n21396, n21397, n21398, n21399, n21400, n21401, n21402,
    n21403, n21404, n21405, n21406, n21407, n21408, n21409, n21410, n21411,
    n21412, n21413, n21414, n21415, n21416, n21417, n21418, n21419, n21420,
    n21421, n21422, n21423, n21424, n21425, n21426, n21427, n21428, n21429,
    n21430, n21431, n21432, n21433, n21434, n21435, n21436, n21437, n21438,
    n21439, n21440, n21441, n21442, n21443, n21444, n21445, n21446, n21447,
    n21448, n21449, n21450, n21451, n21452, n21453, n21454, n21455, n21456,
    n21457, n21458, n21459, n21460, n21461, n21462, n21463, n21464, n21465,
    n21466, n21467, n21468, n21469, n21470, n21471, n21472, n21474, n21475,
    n21476, n21477, n21478, n21479, n21480, n21481, n21482, n21483, n21484,
    n21485, n21486, n21487, n21488, n21489, n21490, n21491, n21492, n21493,
    n21494, n21495, n21496, n21497, n21498, n21499, n21500, n21501, n21502,
    n21503, n21504, n21505, n21506, n21507, n21508, n21509, n21510, n21511,
    n21512, n21513, n21514, n21515, n21517, n21518, n21519, n21520, n21521,
    n21522, n21523, n21524, n21525, n21526, n21527, n21528, n21529, n21530,
    n21531, n21532, n21533, n21534, n21535, n21536, n21537, n21538, n21539,
    n21540, n21541, n21542, n21543, n21544, n21545, n21546, n21547, n21548,
    n21550, n21551, n21552, n21553, n21554, n21555, n21556, n21557, n21558,
    n21559, n21560, n21561, n21562, n21563, n21564, n21565, n21566, n21567,
    n21568, n21569, n21570, n21571, n21572, n21573, n21574, n21575, n21576,
    n21577, n21578, n21579, n21580, n21581, n21582, n21583, n21584, n21585,
    n21586, n21587, n21588, n21589, n21590, n21591, n21592, n21593, n21594,
    n21595, n21596, n21597, n21598, n21599, n21600, n21601, n21602, n21603,
    n21604, n21605, n21606, n21607, n21608, n21609, n21610, n21611, n21612,
    n21613, n21614, n21615, n21616, n21617, n21618, n21619, n21620, n21621,
    n21622, n21623, n21624, n21625, n21626, n21627, n21628, n21629, n21630,
    n21631, n21632, n21633, n21634, n21635, n21636, n21637, n21638, n21639,
    n21640, n21641, n21642, n21643, n21644, n21645, n21646, n21647, n21648,
    n21649, n21650, n21651, n21653, n21654, n21655, n21656, n21657, n21658,
    n21659, n21660, n21661, n21662, n21663, n21664, n21665, n21666, n21667,
    n21668, n21669, n21670, n21671, n21672, n21673, n21674, n21675, n21676,
    n21677, n21678, n21679, n21680, n21681, n21682, n21683, n21684, n21685,
    n21686, n21687, n21689, n21690, n21691, n21692, n21693, n21694, n21695,
    n21696, n21697, n21698, n21699, n21700, n21701, n21702, n21703, n21704,
    n21705, n21706, n21707, n21708, n21709, n21710, n21711, n21712, n21713,
    n21714, n21715, n21716, n21717, n21718, n21719, n21720, n21721, n21722,
    n21723, n21724, n21725, n21726, n21727, n21728, n21729, n21730, n21731,
    n21732, n21733, n21734, n21735, n21736, n21737, n21738, n21739, n21740,
    n21741, n21742, n21743, n21744, n21745, n21746, n21747, n21748, n21749,
    n21750, n21751, n21752, n21753, n21754, n21755, n21756, n21757, n21758,
    n21759, n21760, n21761, n21762, n21763, n21764, n21765, n21766, n21767,
    n21768, n21769, n21770, n21771, n21772, n21773, n21774, n21775, n21776,
    n21777, n21778, n21779, n21780, n21781, n21782, n21783, n21784, n21785,
    n21786, n21787, n21788, n21789, n21791, n21792, n21793, n21794, n21795,
    n21796, n21797, n21798, n21799, n21800, n21801, n21802, n21803, n21804,
    n21805, n21806, n21807, n21808, n21809, n21810, n21811, n21812, n21813,
    n21814, n21815, n21816, n21817, n21818, n21819, n21820, n21821, n21822,
    n21824, n21825, n21826, n21827, n21828, n21829, n21830, n21831, n21832,
    n21833, n21834, n21835, n21836, n21837, n21838, n21839, n21840, n21841,
    n21842, n21843, n21844, n21845, n21846, n21847, n21848, n21849, n21850,
    n21851, n21852, n21853, n21854, n21855, n21856, n21857, n21858, n21859,
    n21860, n21861, n21862, n21863, n21864, n21865, n21866, n21867, n21868,
    n21869, n21870, n21871, n21872, n21873, n21874, n21875, n21876, n21877,
    n21878, n21879, n21880, n21881, n21882, n21883, n21884, n21885, n21886,
    n21887, n21888, n21889, n21890, n21891, n21892, n21893, n21894, n21895,
    n21896, n21897, n21898, n21899, n21900, n21901, n21902, n21903, n21904,
    n21905, n21906, n21907, n21908, n21909, n21910, n21911, n21912, n21913,
    n21915, n21916, n21917, n21918, n21919, n21920, n21921, n21922, n21923,
    n21924, n21925, n21926, n21927, n21928, n21929, n21930, n21931, n21932,
    n21933, n21934, n21935, n21936, n21937, n21938, n21939, n21940, n21941,
    n21942, n21943, n21944, n21945, n21946, n21947, n21948, n21949, n21950,
    n21951, n21952, n21953, n21954, n21955, n21956, n21957, n21958, n21959,
    n21960, n21961, n21962, n21963, n21964, n21965, n21966, n21967, n21968,
    n21969, n21970, n21971, n21972, n21973, n21974, n21975, n21976, n21977,
    n21978, n21979, n21980, n21981, n21982, n21983, n21984, n21985, n21986,
    n21987, n21988, n21989, n21990, n21991, n21992, n21993, n21994, n21995,
    n21996, n21997, n21998, n21999, n22000, n22001, n22002, n22003, n22004,
    n22005, n22006, n22007, n22008, n22009, n22010, n22011, n22012, n22013,
    n22014, n22015, n22016, n22017, n22018, n22019, n22020, n22022, n22023,
    n22024, n22025, n22026, n22027, n22028, n22029, n22030, n22031, n22032,
    n22033, n22034, n22035, n22036, n22037, n22038, n22039, n22040, n22041,
    n22042, n22043, n22044, n22045, n22046, n22047, n22048, n22049, n22050,
    n22051, n22052, n22053, n22054, n22055, n22056, n22057, n22058, n22059,
    n22061, n22062, n22063, n22064, n22065, n22066, n22067, n22068, n22069,
    n22070, n22071, n22072, n22073, n22074, n22075, n22076, n22077, n22078,
    n22079, n22080, n22081, n22082, n22083, n22084, n22085, n22086, n22087,
    n22088, n22089, n22090, n22091, n22092, n22093, n22094, n22095, n22096,
    n22097, n22098, n22099, n22100, n22101, n22102, n22103, n22104, n22105,
    n22106, n22107, n22108, n22109, n22110, n22111, n22112, n22113, n22114,
    n22115, n22116, n22117, n22118, n22119, n22120, n22121, n22122, n22123,
    n22124, n22125, n22126, n22127, n22128, n22129, n22130, n22131, n22132,
    n22133, n22134, n22135, n22136, n22137, n22138, n22139, n22140, n22141,
    n22142, n22143, n22144, n22145, n22146, n22147, n22148, n22149, n22150,
    n22151, n22152, n22153, n22154, n22155, n22156, n22157, n22158, n22159,
    n22160, n22161, n22162, n22164, n22165, n22166, n22167, n22168, n22169,
    n22170, n22171, n22172, n22173, n22174, n22175, n22176, n22177, n22178,
    n22179, n22180, n22181, n22182, n22183, n22184, n22185, n22186, n22187,
    n22188, n22189, n22190, n22191, n22192, n22193, n22194, n22195, n22196,
    n22197, n22198, n22199, n22200, n22201, n22202, n22203, n22204, n22205,
    n22206, n22207, n22208, n22209, n22210, n22211, n22212, n22213, n22214,
    n22216, n22217, n22218, n22219, n22220, n22221, n22222, n22223, n22224,
    n22225, n22226, n22227, n22228, n22229, n22230, n22231, n22232, n22233,
    n22234, n22235, n22236, n22237, n22238, n22239, n22240, n22241, n22242,
    n22243, n22244, n22245, n22246, n22247, n22248, n22249, n22250, n22251,
    n22252, n22253, n22255, n22256, n22257, n22258, n22259, n22260, n22261,
    n22262, n22263, n22264, n22265, n22266, n22267, n22268, n22269, n22270,
    n22271, n22272, n22273, n22274, n22275, n22276, n22277, n22278, n22279,
    n22280, n22281, n22282, n22283, n22284, n22285, n22286, n22287, n22288,
    n22289, n22290, n22291, n22292, n22294, n22295, n22296, n22297, n22298,
    n22299, n22300, n22301, n22302, n22303, n22304, n22305, n22306, n22307,
    n22308, n22309, n22310, n22311, n22312, n22313, n22314, n22315, n22316,
    n22317, n22318, n22319, n22320, n22321, n22322, n22323, n22324, n22325,
    n22326, n22327, n22328, n22329, n22330, n22331, n22332, n22334, n22335,
    n22336, n22337, n22338, n22339, n22340, n22341, n22342, n22343, n22344,
    n22345, n22346, n22347, n22348, n22349, n22350, n22351, n22352, n22353,
    n22354, n22355, n22356, n22357, n22358, n22359, n22360, n22361, n22362,
    n22363, n22364, n22365, n22366, n22367, n22368, n22369, n22370, n22371,
    n22372, n22373, n22374, n22375, n22376, n22377, n22378, n22379, n22380,
    n22381, n22382, n22383, n22384, n22385, n22386, n22387, n22388, n22389,
    n22390, n22391, n22392, n22393, n22394, n22395, n22396, n22397, n22398,
    n22399, n22400, n22401, n22402, n22403, n22404, n22405, n22406, n22407,
    n22408, n22409, n22410, n22411, n22412, n22413, n22414, n22415, n22416,
    n22417, n22418, n22419, n22420, n22421, n22422, n22423, n22424, n22425,
    n22426, n22427, n22428, n22429, n22430, n22431, n22432, n22434, n22435,
    n22436, n22437, n22438, n22439, n22440, n22441, n22442, n22443, n22444,
    n22445, n22446, n22447, n22448, n22449, n22450, n22451, n22452, n22453,
    n22454, n22455, n22456, n22457, n22458, n22459, n22460, n22461, n22462,
    n22463, n22464, n22465, n22466, n22467, n22468, n22469, n22470, n22471,
    n22472, n22473, n22475, n22476, n22477, n22478, n22479, n22480, n22481,
    n22482, n22483, n22484, n22485, n22486, n22487, n22488, n22489, n22490,
    n22491, n22492, n22493, n22494, n22495, n22496, n22497, n22498, n22499,
    n22500, n22501, n22502, n22503, n22504, n22505, n22506, n22507, n22508,
    n22509, n22510, n22511, n22512, n22513, n22515, n22516, n22517, n22518,
    n22519, n22520, n22521, n22522, n22523, n22524, n22525, n22526, n22527,
    n22528, n22529, n22530, n22531, n22532, n22533, n22534, n22535, n22536,
    n22537, n22538, n22539, n22540, n22541, n22542, n22543, n22544, n22545,
    n22546, n22547, n22548, n22549, n22550, n22551, n22552, n22553, n22554,
    n22556, n22557, n22558, n22559, n22560, n22561, n22562, n22563, n22564,
    n22565, n22566, n22567, n22568, n22569, n22570, n22571, n22572, n22573,
    n22574, n22575, n22576, n22577, n22578, n22579, n22580, n22581, n22582,
    n22583, n22584, n22585, n22586, n22587, n22588, n22589, n22590, n22591,
    n22592, n22594, n22595, n22596, n22597, n22598, n22599, n22600, n22601,
    n22602, n22603, n22604, n22605, n22606, n22607, n22608, n22609, n22610,
    n22611, n22612, n22613, n22614, n22615, n22616, n22617, n22618, n22619,
    n22620, n22621, n22622, n22623, n22624, n22625, n22626, n22627, n22628,
    n22629, n22630, n22631, n22632, n22633, n22635, n22636, n22637, n22638,
    n22639, n22640, n22641, n22642, n22643, n22644, n22645, n22646, n22647,
    n22648, n22649, n22650, n22651, n22652, n22653, n22654, n22655, n22656,
    n22657, n22658, n22659, n22660, n22661, n22662, n22663, n22664, n22665,
    n22666, n22667, n22668, n22669, n22670, n22671, n22672, n22673, n22674,
    n22676, n22677, n22678, n22679, n22680, n22681, n22682, n22683, n22684,
    n22685, n22686, n22687, n22688, n22689, n22690, n22691, n22692, n22693,
    n22694, n22695, n22696, n22697, n22698, n22699, n22700, n22701, n22702,
    n22703, n22704, n22705, n22706, n22707, n22708, n22710, n22711, n22712,
    n22713, n22714, n22715, n22716, n22717, n22718, n22719, n22720, n22721,
    n22722, n22723, n22724, n22725, n22726, n22727, n22728, n22729, n22730,
    n22731, n22732, n22733, n22734, n22735, n22736, n22737, n22738, n22739,
    n22740, n22741, n22742, n22743, n22744, n22746, n22747, n22748, n22749,
    n22750, n22751, n22752, n22753, n22754, n22755, n22756, n22757, n22758,
    n22759, n22760, n22761, n22762, n22763, n22764, n22765, n22766, n22767,
    n22768, n22769, n22770, n22771, n22772, n22773, n22774, n22775, n22776,
    n22777, n22778, n22779, n22780, n22781, n22782, n22783, n22784, n22785,
    n22786, n22787, n22788, n22789, n22790, n22791, n22792, n22793, n22794,
    n22795, n22796, n22797, n22798, n22799, n22800, n22801, n22802, n22803,
    n22804, n22805, n22806, n22807, n22808, n22809, n22810, n22811, n22812,
    n22813, n22814, n22815, n22816, n22817, n22818, n22819, n22820, n22821,
    n22822, n22823, n22824, n22825, n22826, n22827, n22828, n22829, n22830,
    n22831, n22832, n22833, n22834, n22835, n22836, n22837, n22838, n22839,
    n22840, n22842, n22843, n22844, n22845, n22846, n22847, n22848, n22849,
    n22850, n22851, n22852, n22853, n22854, n22855, n22856, n22857, n22858,
    n22859, n22860, n22861, n22862, n22863, n22864, n22865, n22866, n22867,
    n22868, n22869, n22870, n22871, n22873, n22874, n22875, n22876, n22877,
    n22878, n22879, n22880, n22881, n22882, n22883, n22884, n22885, n22886,
    n22887, n22888, n22889, n22890, n22891, n22892, n22893, n22894, n22895,
    n22896, n22897, n22898, n22899, n22900, n22901, n22902, n22903, n22904,
    n22905, n22906, n22907, n22908, n22909, n22910, n22912, n22913, n22914,
    n22915, n22916, n22917, n22918, n22919, n22920, n22921, n22922, n22923,
    n22924, n22925, n22926, n22927, n22928, n22929, n22930, n22931, n22932,
    n22933, n22934, n22935, n22936, n22937, n22938, n22940, n22941, n22942,
    n22943, n22944, n22945, n22946, n22947, n22948, n22949, n22950, n22951,
    n22952, n22953, n22954, n22955, n22956, n22957, n22958, n22959, n22960,
    n22961, n22962, n22963, n22964, n22965, n22966, n22967, n22968, n22969,
    n22970, n22971, n22972, n22973, n22974, n22975, n22976, n22977, n22978,
    n22979, n22980, n22981, n22983, n22984, n22985, n22986, n22987, n22988,
    n22989, n22990, n22991, n22992, n22993, n22994, n22995, n22996, n22997,
    n22998, n22999, n23000, n23001, n23002, n23003, n23004, n23005, n23006,
    n23007, n23008, n23009, n23010, n23011, n23012, n23013, n23014, n23015,
    n23016, n23017, n23019, n23020, n23021, n23022, n23023, n23024, n23025,
    n23026, n23027, n23028, n23029, n23030, n23031, n23032, n23033, n23034,
    n23035, n23036, n23037, n23038, n23039, n23040, n23041, n23042, n23043,
    n23044, n23045, n23046, n23047, n23048, n23049, n23050, n23051, n23052,
    n23053, n23054, n23055, n23056, n23057, n23058, n23059, n23060, n23061,
    n23062, n23063, n23064, n23066, n23067, n23068, n23069, n23070, n23071,
    n23072, n23073, n23074, n23075, n23076, n23077, n23078, n23079, n23080,
    n23081, n23082, n23083, n23084, n23085, n23086, n23087, n23088, n23089,
    n23090, n23091, n23092, n23093, n23094, n23096, n23097, n23098, n23099,
    n23100, n23101, n23102, n23103, n23104, n23105, n23106, n23107, n23108,
    n23109, n23110, n23111, n23112, n23113, n23114, n23115, n23116, n23117,
    n23118, n23119, n23120, n23121, n23122, n23123, n23124, n23125, n23126,
    n23127, n23128, n23129, n23130, n23131, n23132, n23133, n23134, n23135,
    n23136, n23137, n23138, n23139, n23140, n23141, n23142, n23143, n23144,
    n23145, n23146, n23147, n23148, n23149, n23150, n23151, n23152, n23153,
    n23154, n23155, n23156, n23157, n23158, n23159, n23160, n23161, n23162,
    n23163, n23164, n23165, n23166, n23167, n23168, n23169, n23170, n23171,
    n23172, n23173, n23174, n23175, n23176, n23177, n23178, n23179, n23180,
    n23181, n23182, n23183, n23184, n23185, n23186, n23187, n23188, n23189,
    n23190, n23191, n23192, n23193, n23194, n23195, n23196, n23197, n23198,
    n23199, n23200, n23202, n23203, n23204, n23205, n23206, n23207, n23208,
    n23209, n23210, n23211, n23212, n23213, n23214, n23215, n23216, n23217,
    n23218, n23219, n23220, n23221, n23222, n23223, n23224, n23225, n23226,
    n23227, n23228, n23229, n23230, n23231, n23232, n23233, n23234, n23235,
    n23236, n23237, n23238, n23239, n23240, n23241, n23242, n23243, n23244,
    n23245, n23246, n23247, n23248, n23249, n23250, n23251, n23252, n23253,
    n23254, n23255, n23256, n23257, n23258, n23259, n23260, n23261, n23262,
    n23263, n23264, n23265, n23266, n23267, n23268, n23269, n23270, n23271,
    n23272, n23273, n23274, n23275, n23276, n23277, n23278, n23279, n23280,
    n23281, n23282, n23283, n23284, n23285, n23286, n23287, n23288, n23289,
    n23290, n23291, n23292, n23293, n23294, n23295, n23296, n23297, n23298,
    n23299, n23300, n23301, n23302, n23303, n23305, n23306, n23307, n23308,
    n23309, n23310, n23311, n23312, n23313, n23314, n23315, n23316, n23317,
    n23318, n23319, n23320, n23321, n23322, n23323, n23324, n23325, n23326,
    n23327, n23328, n23329, n23330, n23331, n23332, n23333, n23334, n23335,
    n23336, n23337, n23338, n23339, n23340, n23341, n23342, n23343, n23344,
    n23345, n23346, n23347, n23348, n23349, n23350, n23351, n23352, n23353,
    n23354, n23355, n23356, n23357, n23358, n23359, n23360, n23361, n23362,
    n23363, n23364, n23365, n23366, n23367, n23368, n23369, n23370, n23371,
    n23372, n23373, n23374, n23375, n23376, n23377, n23378, n23379, n23380,
    n23381, n23382, n23383, n23384, n23385, n23386, n23387, n23388, n23389,
    n23390, n23391, n23392, n23393, n23394, n23395, n23396, n23397, n23398,
    n23399, n23400, n23401, n23402, n23403, n23404, n23405, n23407, n23408,
    n23409, n23410, n23411, n23412, n23413, n23414, n23415, n23416, n23417,
    n23418, n23419, n23420, n23421, n23422, n23423, n23424, n23425, n23426,
    n23427, n23428, n23429, n23430, n23431, n23432, n23433, n23434, n23435,
    n23436, n23437, n23438, n23439, n23440, n23441, n23442, n23443, n23444,
    n23446, n23447, n23448, n23449, n23450, n23451, n23452, n23453, n23454,
    n23455, n23456, n23457, n23458, n23459, n23460, n23461, n23462, n23463,
    n23464, n23465, n23466, n23467, n23468, n23469, n23470, n23471, n23472,
    n23473, n23474, n23475, n23476, n23477, n23478, n23479, n23480, n23481,
    n23482, n23483, n23484, n23485, n23486, n23488, n23489, n23490, n23491,
    n23492, n23493, n23494, n23495, n23496, n23497, n23498, n23499, n23500,
    n23501, n23502, n23503, n23504, n23505, n23506, n23507, n23508, n23509,
    n23510, n23511, n23512, n23513, n23514, n23515, n23516, n23517, n23518,
    n23519, n23520, n23521, n23522, n23523, n23524, n23525, n23526, n23527,
    n23528, n23530, n23531, n23532, n23533, n23534, n23535, n23536, n23537,
    n23538, n23539, n23540, n23541, n23542, n23543, n23544, n23545, n23546,
    n23547, n23548, n23549, n23550, n23551, n23552, n23553, n23554, n23555,
    n23556, n23557, n23558, n23559, n23560, n23561, n23563, n23564, n23565,
    n23566, n23567, n23568, n23569, n23570, n23571, n23572, n23573, n23574,
    n23575, n23576, n23577, n23578, n23579, n23580, n23581, n23582, n23583,
    n23584, n23585, n23586, n23587, n23588, n23589, n23590, n23591, n23592,
    n23593, n23594, n23595, n23596, n23597, n23598, n23599, n23601, n23602,
    n23603, n23604, n23605, n23606, n23607, n23608, n23609, n23610, n23611,
    n23612, n23613, n23614, n23615, n23616, n23617, n23618, n23619, n23620,
    n23621, n23622, n23623, n23624, n23625, n23626, n23627, n23628, n23629,
    n23630, n23631, n23632, n23633, n23634, n23635, n23636, n23637, n23638,
    n23639, n23640, n23641, n23642, n23643, n23644, n23645, n23646, n23647,
    n23648, n23649, n23650, n23651, n23652, n23653, n23654, n23655, n23656,
    n23657, n23658, n23659, n23660, n23661, n23662, n23663, n23664, n23665,
    n23666, n23667, n23668, n23669, n23670, n23671, n23672, n23673, n23674,
    n23675, n23676, n23677, n23678, n23679, n23680, n23681, n23682, n23683,
    n23684, n23685, n23686, n23687, n23688, n23689, n23690, n23691, n23692,
    n23693, n23694, n23695, n23696, n23697, n23698, n23700, n23701, n23702,
    n23703, n23704, n23705, n23706, n23707, n23708, n23709, n23710, n23711,
    n23712, n23713, n23714, n23715, n23716, n23717, n23718, n23719, n23720,
    n23721, n23722, n23723, n23724, n23725, n23726, n23727, n23728, n23729,
    n23730, n23731, n23732, n23733, n23734, n23736, n23737, n23738, n23739,
    n23740, n23741, n23742, n23743, n23744, n23745, n23746, n23747, n23748,
    n23749, n23750, n23751, n23752, n23753, n23754, n23755, n23756, n23757,
    n23758, n23759, n23760, n23761, n23762, n23763, n23764, n23765, n23766,
    n23767, n23768, n23769, n23770, n23771, n23772, n23773, n23774, n23775,
    n23776, n23777, n23778, n23779, n23780, n23781, n23782, n23783, n23784,
    n23785, n23786, n23787, n23788, n23789, n23790, n23791, n23792, n23793,
    n23794, n23795, n23796, n23797, n23798, n23799, n23800, n23801, n23802,
    n23803, n23804, n23805, n23806, n23807, n23808, n23809, n23810, n23811,
    n23812, n23813, n23814, n23815, n23816, n23817, n23818, n23819, n23820,
    n23821, n23822, n23823, n23824, n23825, n23826, n23827, n23828, n23829,
    n23830, n23831, n23832, n23833, n23834, n23835, n23836, n23837, n23839,
    n23840, n23841, n23842, n23843, n23844, n23845, n23846, n23847, n23848,
    n23849, n23850, n23851, n23852, n23853, n23854, n23855, n23856, n23857,
    n23858, n23859, n23860, n23861, n23862, n23863, n23864, n23865, n23866,
    n23867, n23868, n23869, n23870, n23871, n23872, n23873, n23874, n23875,
    n23876, n23877, n23878, n23879, n23880, n23881, n23882, n23883, n23884,
    n23885, n23886, n23887, n23888, n23889, n23890, n23891, n23892, n23893,
    n23894, n23895, n23896, n23897, n23898, n23899, n23900, n23901, n23902,
    n23903, n23904, n23905, n23906, n23907, n23908, n23909, n23910, n23911,
    n23912, n23913, n23914, n23915, n23916, n23917, n23918, n23919, n23920,
    n23921, n23922, n23923, n23924, n23925, n23926, n23927, n23928, n23929,
    n23930, n23931, n23932, n23933, n23934, n23935, n23936, n23937, n23938,
    n23939, n23940, n23941, n23942, n23943, n23944, n23946, n23947, n23948,
    n23949, n23950, n23951, n23952, n23953, n23954, n23955, n23956, n23957,
    n23958, n23959, n23960, n23961, n23962, n23963, n23964, n23965, n23966,
    n23967, n23968, n23969, n23970, n23971, n23972, n23973, n23974, n23975,
    n23976, n23977, n23978, n23980, n23981, n23982, n23983, n23984, n23985,
    n23986, n23987, n23988, n23989, n23990, n23991, n23992, n23993, n23994,
    n23995, n23996, n23997, n23998, n23999, n24000, n24001, n24002, n24003,
    n24004, n24005, n24006, n24007, n24008, n24009, n24010, n24011, n24012,
    n24013, n24014, n24015, n24016, n24017, n24019, n24020, n24021, n24022,
    n24023, n24024, n24025, n24026, n24027, n24028, n24029, n24030, n24031,
    n24032, n24033, n24034, n24035, n24036, n24037, n24038, n24039, n24040,
    n24041, n24042, n24043, n24044, n24045, n24046, n24047, n24048, n24049,
    n24050, n24051, n24052, n24053, n24054, n24055, n24056, n24057, n24058,
    n24060, n24061, n24062, n24063, n24064, n24065, n24066, n24067, n24068,
    n24069, n24070, n24071, n24072, n24073, n24074, n24075, n24076, n24077,
    n24078, n24079, n24080, n24081, n24082, n24083, n24084, n24085, n24086,
    n24087, n24088, n24089, n24090, n24091, n24092, n24093, n24094, n24095,
    n24096, n24097, n24098, n24099, n24100, n24101, n24102, n24103, n24104,
    n24105, n24106, n24108, n24109, n24110, n24111, n24112, n24113, n24114,
    n24115, n24116, n24117, n24118, n24119, n24120, n24121, n24122, n24123,
    n24124, n24125, n24126, n24127, n24128, n24129, n24130, n24131, n24132,
    n24133, n24134, n24135, n24136, n24137, n24138, n24139, n24140, n24141,
    n24142, n24143, n24144, n24145, n24146, n24147, n24148, n24149, n24150,
    n24151, n24152, n24153, n24154, n24155, n24156, n24157, n24158, n24159,
    n24160, n24161, n24162, n24163, n24164, n24165, n24166, n24167, n24168,
    n24169, n24170, n24171, n24172, n24173, n24174, n24175, n24176, n24177,
    n24178, n24179, n24180, n24181, n24182, n24183, n24184, n24185, n24186,
    n24187, n24188, n24189, n24190, n24191, n24192, n24193, n24194, n24195,
    n24196, n24197, n24199, n24200, n24201, n24202, n24203, n24204, n24205,
    n24206, n24207, n24208, n24209, n24210, n24211, n24212, n24213, n24214,
    n24215, n24216, n24217, n24218, n24219, n24220, n24221, n24222, n24223,
    n24224, n24225, n24226, n24227, n24228, n24229, n24230, n24231, n24232,
    n24233, n24234, n24235, n24236, n24237, n24238, n24239, n24240, n24241,
    n24242, n24243, n24244, n24245, n24246, n24247, n24248, n24249, n24251,
    n24252, n24253, n24254, n24255, n24256, n24257, n24258, n24259, n24260,
    n24261, n24262, n24263, n24264, n24265, n24266, n24267, n24268, n24269,
    n24270, n24271, n24272, n24273, n24274, n24275, n24276, n24277, n24278,
    n24279, n24280, n24281, n24282, n24283, n24284, n24285, n24286, n24287,
    n24288, n24289, n24291, n24292, n24293, n24294, n24295, n24296, n24297,
    n24298, n24299, n24300, n24301, n24302, n24303, n24304, n24305, n24306,
    n24307, n24308, n24309, n24310, n24311, n24312, n24313, n24314, n24315,
    n24316, n24317, n24318, n24319, n24320, n24321, n24322, n24323, n24324,
    n24325, n24326, n24327, n24328, n24329, n24330, n24331, n24332, n24333,
    n24334, n24335, n24336, n24337, n24338, n24339, n24340, n24341, n24342,
    n24343, n24344, n24345, n24346, n24347, n24348, n24349, n24350, n24351,
    n24352, n24353, n24354, n24355, n24356, n24357, n24358, n24359, n24360,
    n24361, n24362, n24363, n24364, n24365, n24366, n24367, n24368, n24369,
    n24370, n24371, n24372, n24373, n24374, n24375, n24376, n24377, n24378,
    n24379, n24380, n24381, n24382, n24383, n24384, n24385, n24386, n24388,
    n24389, n24390, n24391, n24392, n24393, n24394, n24395, n24396, n24397,
    n24398, n24399, n24400, n24401, n24402, n24403, n24404, n24405, n24406,
    n24407, n24408, n24409, n24410, n24411, n24412, n24413, n24414, n24415,
    n24416, n24417, n24418, n24419, n24420, n24421, n24422, n24423, n24424,
    n24425, n24426, n24427, n24429, n24430, n24431, n24432, n24433, n24434,
    n24435, n24436, n24437, n24438, n24439, n24440, n24441, n24442, n24443,
    n24444, n24445, n24446, n24447, n24448, n24449, n24450, n24451, n24452,
    n24453, n24454, n24455, n24456, n24457, n24459, n24460, n24461, n24462,
    n24463, n24464, n24465, n24466, n24467, n24468, n24469, n24470, n24471,
    n24472, n24473, n24474, n24475, n24476, n24477, n24478, n24479, n24480,
    n24481, n24482, n24483, n24484, n24485, n24486, n24487, n24488, n24490,
    n24491, n24492, n24493, n24494, n24495, n24496, n24497, n24498, n24499,
    n24500, n24501, n24502, n24503, n24504, n24505, n24506, n24507, n24508,
    n24509, n24510, n24511, n24512, n24513, n24514, n24515, n24516, n24517,
    n24518, n24519, n24520, n24521, n24522, n24523, n24524, n24525, n24526,
    n24527, n24528, n24529, n24531, n24532, n24533, n24534, n24535, n24536,
    n24537, n24538, n24539, n24540, n24541, n24542, n24543, n24544, n24545,
    n24546, n24547, n24548, n24549, n24550, n24551, n24552, n24553, n24554,
    n24555, n24556, n24557, n24558, n24559, n24560, n24561, n24562, n24563,
    n24564, n24565, n24566, n24567, n24568, n24569, n24570, n24571, n24572,
    n24574, n24575, n24576, n24577, n24578, n24579, n24580, n24581, n24582,
    n24583, n24584, n24585, n24586, n24587, n24588, n24589, n24590, n24591,
    n24592, n24593, n24594, n24595, n24596, n24597, n24598, n24599, n24600,
    n24601, n24602, n24603, n24604, n24605, n24606, n24607, n24608, n24609,
    n24610, n24611, n24613, n24614, n24615, n24616, n24617, n24618, n24619,
    n24620, n24621, n24622, n24623, n24624, n24625, n24626, n24627, n24628,
    n24629, n24630, n24631, n24632, n24633, n24634, n24635, n24636, n24637,
    n24638, n24639, n24640, n24641, n24642, n24643, n24644, n24645, n24646,
    n24647, n24649, n24650, n24651, n24652, n24653, n24654, n24655, n24656,
    n24657, n24658, n24659, n24660, n24661, n24662, n24663, n24664, n24665,
    n24666, n24667, n24668, n24669, n24670, n24671, n24672, n24673, n24674,
    n24675, n24676, n24677, n24678, n24679, n24680, n24681, n24682, n24683,
    n24684, n24685, n24686, n24687, n24689, n24690, n24691, n24692, n24693,
    n24694, n24695, n24696, n24697, n24698, n24699, n24700, n24701, n24702,
    n24703, n24704, n24705, n24706, n24707, n24708, n24709, n24710, n24711,
    n24712, n24713, n24714, n24715, n24716, n24717, n24718, n24719, n24720,
    n24721, n24722, n24723, n24724, n24725, n24726, n24727, n24729, n24730,
    n24731, n24732, n24733, n24734, n24735, n24736, n24737, n24738, n24739,
    n24740, n24741, n24742, n24743, n24744, n24745, n24746, n24747, n24748,
    n24749, n24750, n24751, n24752, n24753, n24754, n24755, n24756, n24757,
    n24758, n24759, n24760, n24761, n24762, n24763, n24765, n24766, n24767,
    n24768, n24769, n24770, n24771, n24772, n24773, n24774, n24775, n24776,
    n24777, n24778, n24779, n24780, n24781, n24782, n24783, n24784, n24785,
    n24786, n24787, n24788, n24789, n24790, n24791, n24793, n24794, n24795,
    n24796, n24797, n24798, n24799, n24800, n24801, n24802, n24803, n24804,
    n24805, n24806, n24807, n24808, n24809, n24810, n24811, n24812, n24813,
    n24814, n24815, n24816, n24817, n24818, n24819, n24820, n24821, n24822,
    n24823, n24824, n24825, n24826, n24827, n24829, n24830, n24831, n24832,
    n24833, n24834, n24835, n24836, n24837, n24838, n24839, n24840, n24841,
    n24842, n24843, n24844, n24845, n24846, n24847, n24848, n24849, n24850,
    n24851, n24852, n24853, n24854, n24855, n24856, n24857, n24858, n24859,
    n24860, n24861, n24862, n24863, n24864, n24865, n24866, n24867, n24868,
    n24869, n24870, n24871, n24872, n24873, n24874, n24875, n24876, n24877,
    n24878, n24879, n24880, n24881, n24882, n24883, n24884, n24885, n24886,
    n24887, n24888, n24889, n24890, n24891, n24892, n24893, n24894, n24895,
    n24896, n24897, n24898, n24899, n24900, n24901, n24902, n24903, n24904,
    n24905, n24906, n24907, n24908, n24909, n24910, n24911, n24912, n24913,
    n24914, n24915, n24916, n24917, n24918, n24919, n24920, n24921, n24922,
    n24923, n24924, n24925, n24926, n24927, n24928, n24929, n24930, n24931,
    n24932, n24933, n24934, n24936, n24937, n24938, n24939, n24940, n24941,
    n24942, n24943, n24944, n24945, n24946, n24947, n24948, n24949, n24950,
    n24951, n24952, n24953, n24954, n24955, n24956, n24957, n24958, n24959,
    n24960, n24961, n24962, n24963, n24964, n24965, n24966, n24967, n24968,
    n24969, n24970, n24971, n24972, n24973, n24974, n24975, n24976, n24977,
    n24978, n24979, n24980, n24981, n24982, n24983, n24984, n24985, n24986,
    n24987, n24988, n24989, n24990, n24991, n24992, n24993, n24994, n24995,
    n24996, n24997, n24998, n24999, n25000, n25001, n25002, n25003, n25004,
    n25005, n25006, n25007, n25008, n25009, n25010, n25011, n25012, n25013,
    n25014, n25015, n25016, n25017, n25018, n25019, n25020, n25021, n25022,
    n25023, n25024, n25025, n25026, n25027, n25028, n25029, n25030, n25031,
    n25032, n25033, n25034, n25035, n25036, n25037, n25038, n25040, n25041,
    n25042, n25043, n25044, n25045, n25046, n25047, n25048, n25049, n25050,
    n25051, n25052, n25053, n25054, n25055, n25056, n25057, n25058, n25059,
    n25060, n25061, n25062, n25063, n25064, n25065, n25066, n25067, n25068,
    n25069, n25070, n25072, n25073, n25074, n25075, n25076, n25077, n25078,
    n25079, n25080, n25081, n25082, n25083, n25084, n25085, n25086, n25087,
    n25088, n25089, n25090, n25091, n25092, n25093, n25094, n25095, n25096,
    n25097, n25098, n25099, n25100, n25101, n25102, n25103, n25104, n25105,
    n25106, n25107, n25108, n25109, n25110, n25111, n25112, n25113, n25114,
    n25115, n25116, n25117, n25118, n25119, n25120, n25121, n25122, n25123,
    n25124, n25125, n25126, n25127, n25128, n25129, n25130, n25131, n25132,
    n25133, n25134, n25135, n25136, n25137, n25138, n25139, n25140, n25141,
    n25142, n25143, n25144, n25145, n25146, n25147, n25148, n25149, n25150,
    n25151, n25152, n25153, n25154, n25155, n25156, n25157, n25158, n25159,
    n25160, n25161, n25162, n25163, n25164, n25165, n25166, n25167, n25168,
    n25169, n25170, n25171, n25172, n25173, n25174, n25175, n25176, n25177,
    n25179, n25180, n25181, n25182, n25183, n25184, n25185, n25186, n25187,
    n25188, n25189, n25190, n25191, n25192, n25193, n25194, n25195, n25196,
    n25197, n25198, n25199, n25200, n25201, n25202, n25203, n25204, n25205,
    n25206, n25207, n25208, n25209, n25210, n25211, n25212, n25213, n25214,
    n25215, n25216, n25218, n25219, n25220, n25221, n25222, n25223, n25224,
    n25225, n25226, n25227, n25228, n25229, n25230, n25231, n25232, n25233,
    n25234, n25235, n25236, n25237, n25238, n25239, n25240, n25241, n25242,
    n25243, n25244, n25245, n25246, n25247, n25248, n25249, n25250, n25251,
    n25252, n25253, n25254, n25255, n25256, n25257, n25258, n25259, n25260,
    n25261, n25262, n25263, n25264, n25265, n25266, n25267, n25268, n25269,
    n25270, n25271, n25272, n25273, n25274, n25275, n25276, n25277, n25278,
    n25279, n25280, n25281, n25282, n25283, n25284, n25285, n25286, n25287,
    n25288, n25289, n25290, n25291, n25292, n25293, n25294, n25295, n25296,
    n25297, n25298, n25299, n25300, n25301, n25302, n25303, n25304, n25305,
    n25306, n25307, n25308, n25309, n25310, n25311, n25312, n25313, n25314,
    n25315, n25316, n25317, n25318, n25319, n25320, n25322, n25323, n25324,
    n25325, n25326, n25327, n25328, n25329, n25330, n25331, n25332, n25333,
    n25334, n25335, n25336, n25337, n25338, n25339, n25340, n25341, n25342,
    n25343, n25344, n25345, n25346, n25347, n25348, n25349, n25350, n25351,
    n25352, n25353, n25354, n25355, n25356, n25357, n25358, n25359, n25361,
    n25362, n25363, n25364, n25365, n25366, n25367, n25368, n25369, n25370,
    n25371, n25372, n25373, n25374, n25375, n25376, n25377, n25378, n25379,
    n25380, n25381, n25382, n25383, n25384, n25385, n25386, n25387, n25388,
    n25389, n25390, n25391, n25392, n25393, n25394, n25395, n25396, n25397,
    n25398, n25399, n25400, n25401, n25402, n25403, n25404, n25405, n25406,
    n25407, n25408, n25409, n25410, n25411, n25412, n25413, n25414, n25415,
    n25416, n25417, n25418, n25419, n25420, n25421, n25422, n25423, n25424,
    n25425, n25426, n25427, n25428, n25429, n25430, n25431, n25432, n25433,
    n25434, n25435, n25436, n25437, n25438, n25439, n25440, n25441, n25442,
    n25443, n25444, n25445, n25446, n25447, n25448, n25449, n25450, n25451,
    n25452, n25453, n25454, n25455, n25456, n25457, n25458, n25459, n25460,
    n25461, n25462, n25463, n25464, n25466, n25467, n25468, n25469, n25470,
    n25471, n25472, n25473, n25474, n25475, n25476, n25477, n25478, n25479,
    n25480, n25481, n25482, n25483, n25484, n25485, n25486, n25487, n25488,
    n25489, n25490, n25491, n25492, n25493, n25494, n25495, n25496, n25497,
    n25498, n25499, n25500, n25501, n25502, n25503, n25504, n25505, n25506,
    n25507, n25509, n25510, n25511, n25512, n25513, n25514, n25515, n25516,
    n25517, n25518, n25519, n25520, n25521, n25522, n25523, n25524, n25525,
    n25526, n25527, n25528, n25529, n25530, n25531, n25532, n25533, n25534,
    n25535, n25536, n25537, n25538, n25539, n25540, n25541, n25542, n25543,
    n25544, n25545, n25546, n25547, n25548, n25549, n25550, n25551, n25552,
    n25553, n25554, n25555, n25556, n25557, n25558, n25559, n25560, n25561,
    n25562, n25563, n25564, n25565, n25566, n25567, n25568, n25569, n25570,
    n25571, n25572, n25573, n25574, n25575, n25576, n25577, n25578, n25579,
    n25580, n25581, n25582, n25583, n25584, n25585, n25586, n25587, n25588,
    n25589, n25590, n25591, n25592, n25593, n25594, n25595, n25596, n25597,
    n25598, n25599, n25600, n25601, n25602, n25603, n25604, n25605, n25607,
    n25608, n25609, n25610, n25611, n25612, n25613, n25614, n25615, n25616,
    n25617, n25618, n25619, n25620, n25621, n25622, n25623, n25624, n25625,
    n25626, n25627, n25628, n25629, n25630, n25631, n25632, n25633, n25634,
    n25635, n25636, n25637, n25638, n25639, n25640, n25641, n25642, n25643,
    n25644, n25645, n25647, n25648, n25649, n25650, n25651, n25652, n25653,
    n25654, n25655, n25656, n25657, n25658, n25659, n25660, n25661, n25662,
    n25663, n25664, n25665, n25666, n25667, n25668, n25669, n25670, n25671,
    n25672, n25673, n25674, n25675, n25676, n25677, n25678, n25679, n25680,
    n25681, n25682, n25683, n25684, n25685, n25686, n25688, n25689, n25690,
    n25691, n25692, n25693, n25694, n25695, n25696, n25697, n25698, n25699,
    n25700, n25701, n25702, n25703, n25704, n25705, n25706, n25707, n25708,
    n25709, n25710, n25711, n25712, n25713, n25714, n25715, n25716, n25717,
    n25718, n25719, n25720, n25721, n25722, n25723, n25724, n25725, n25726,
    n25727, n25728, n25729, n25730, n25731, n25733, n25734, n25735, n25736,
    n25737, n25738, n25739, n25740, n25741, n25742, n25743, n25744, n25745,
    n25746, n25747, n25748, n25749, n25750, n25751, n25752, n25753, n25754,
    n25755, n25756, n25757, n25758, n25759, n25760, n25761, n25762, n25763,
    n25764, n25765, n25766, n25767, n25768, n25769, n25770, n25771, n25773,
    n25774, n25775, n25776, n25777, n25778, n25779, n25780, n25781, n25782,
    n25783, n25784, n25785, n25786, n25787, n25788, n25789, n25790, n25791,
    n25792, n25793, n25794, n25795, n25796, n25797, n25798, n25799, n25800,
    n25801, n25802, n25803, n25805, n25806, n25807, n25808, n25809, n25810,
    n25811, n25812, n25813, n25814, n25815, n25816, n25817, n25818, n25819,
    n25820, n25821, n25822, n25823, n25824, n25825, n25826, n25827, n25828,
    n25829, n25830, n25831, n25832, n25833, n25834, n25835, n25836, n25837,
    n25838, n25839, n25840, n25841, n25843, n25844, n25845, n25846, n25847,
    n25848, n25849, n25850, n25851, n25852, n25853, n25854, n25855, n25856,
    n25857, n25858, n25859, n25860, n25861, n25862, n25863, n25864, n25865,
    n25866, n25867, n25868, n25869, n25870, n25871, n25872, n25873, n25874,
    n25875, n25876, n25877, n25878, n25879, n25880, n25881, n25882, n25883,
    n25884, n25885, n25886, n25887, n25888, n25889, n25890, n25891, n25892,
    n25893, n25894, n25895, n25896, n25897, n25898, n25899, n25900, n25901,
    n25902, n25903, n25904, n25905, n25906, n25907, n25908, n25909, n25910,
    n25911, n25912, n25913, n25914, n25915, n25916, n25917, n25918, n25919,
    n25920, n25921, n25922, n25923, n25924, n25925, n25926, n25927, n25928,
    n25929, n25930, n25931, n25932, n25933, n25934, n25935, n25936, n25937,
    n25938, n25939, n25940, n25941, n25942, n25943, n25944, n25946, n25947,
    n25948, n25949, n25950, n25951, n25952, n25953, n25954, n25955, n25956,
    n25957, n25958, n25959, n25960, n25961, n25962, n25963, n25964, n25965,
    n25966, n25967, n25968, n25969, n25970, n25971, n25972, n25973, n25974,
    n25975, n25976, n25977, n25978, n25979, n25980, n25982, n25983, n25984,
    n25985, n25986, n25987, n25988, n25989, n25990, n25991, n25992, n25993,
    n25994, n25995, n25996, n25997, n25998, n25999, n26000, n26001, n26002,
    n26003, n26004, n26005, n26006, n26007, n26008, n26009, n26010, n26011,
    n26013, n26014, n26015, n26016, n26017, n26018, n26019, n26020, n26021,
    n26022, n26023, n26024, n26025, n26026, n26027, n26028, n26029, n26030,
    n26031, n26032, n26033, n26034, n26035, n26036, n26037, n26038, n26039,
    n26040, n26041, n26042, n26043, n26044, n26045, n26046, n26047, n26049,
    n26050, n26051, n26052, n26053, n26054, n26055, n26056, n26057, n26058,
    n26059, n26060, n26061, n26062, n26063, n26064, n26065, n26066, n26067,
    n26068, n26069, n26070, n26071, n26072, n26073, n26074, n26075, n26076,
    n26077, n26078, n26079, n26080, n26081, n26082, n26083, n26084, n26085,
    n26087, n26088, n26089, n26090, n26091, n26092, n26093, n26094, n26095,
    n26096, n26097, n26098, n26099, n26100, n26101, n26102, n26103, n26104,
    n26105, n26106, n26107, n26108, n26109, n26110, n26111, n26112, n26113,
    n26114, n26115, n26116, n26117, n26118, n26119, n26120, n26121, n26122,
    n26123, n26124, n26125, n26126, n26127, n26128, n26129, n26130, n26131,
    n26132, n26133, n26134, n26135, n26136, n26137, n26138, n26140, n26141,
    n26142, n26143, n26144, n26145, n26146, n26147, n26148, n26149, n26150,
    n26151, n26152, n26153, n26154, n26155, n26156, n26157, n26158, n26159,
    n26160, n26161, n26162, n26163, n26164, n26165, n26166, n26167, n26168,
    n26169, n26170, n26171, n26172, n26173, n26174, n26175, n26176, n26177,
    n26178, n26180, n26181, n26182, n26183, n26184, n26185, n26186, n26187,
    n26188, n26189, n26190, n26191, n26192, n26193, n26194, n26195, n26196,
    n26197, n26198, n26199, n26200, n26201, n26202, n26203, n26204, n26205,
    n26206, n26207, n26208, n26209, n26210, n26211, n26212, n26213, n26214,
    n26215, n26216, n26217, n26218, n26219, n26220, n26221, n26223, n26224,
    n26225, n26226, n26227, n26228, n26229, n26230, n26231, n26232, n26233,
    n26234, n26235, n26236, n26237, n26238, n26239, n26240, n26241, n26242,
    n26243, n26244, n26245, n26246, n26247, n26248, n26249, n26250, n26251,
    n26252, n26253, n26254, n26255, n26256, n26257, n26259, n26260, n26261,
    n26262, n26263, n26264, n26265, n26266, n26267, n26268, n26269, n26270,
    n26271, n26272, n26273, n26274, n26275, n26276, n26277, n26278, n26279,
    n26280, n26281, n26282, n26283, n26284, n26285, n26286, n26287, n26288,
    n26289, n26290, n26291, n26292, n26293, n26295, n26296, n26297, n26298,
    n26299, n26300, n26301, n26302, n26303, n26304, n26305, n26306, n26307,
    n26308, n26309, n26310, n26311, n26312, n26313, n26314, n26315, n26316,
    n26317, n26318, n26319, n26320, n26321, n26323, n26324, n26325, n26326,
    n26327, n26328, n26329, n26330, n26331, n26332, n26333, n26334, n26335,
    n26336, n26337, n26338, n26339, n26340, n26341, n26342, n26343, n26344,
    n26345, n26346, n26347, n26348, n26349, n26350, n26351, n26353, n26354,
    n26355, n26356, n26357, n26358, n26359, n26360, n26361, n26362, n26363,
    n26364, n26365, n26366, n26367, n26368, n26369, n26370, n26371, n26372,
    n26373, n26374, n26375, n26376, n26377, n26378, n26379, n26380, n26381,
    n26382, n26383, n26384, n26385, n26386, n26387, n26388, n26389, n26390,
    n26391, n26392, n26393, n26394, n26395, n26396, n26397, n26398, n26399,
    n26400, n26401, n26402, n26403, n26404, n26405, n26406, n26407, n26408,
    n26409, n26410, n26411, n26412, n26413, n26414, n26415, n26416, n26417,
    n26418, n26419, n26420, n26421, n26422, n26423, n26424, n26425, n26426,
    n26427, n26428, n26429, n26430, n26431, n26432, n26433, n26434, n26435,
    n26436, n26437, n26438, n26439, n26440, n26441, n26442, n26443, n26444,
    n26445, n26446, n26447, n26448, n26449, n26450, n26452, n26453, n26454,
    n26455, n26456, n26457, n26458, n26459, n26460, n26461, n26462, n26463,
    n26464, n26465, n26466, n26467, n26468, n26469, n26470, n26471, n26472,
    n26473, n26474, n26475, n26476, n26477, n26478, n26479, n26480, n26481,
    n26482, n26483, n26484, n26485, n26486, n26487, n26488, n26489, n26490,
    n26491, n26492, n26493, n26494, n26495, n26497, n26498, n26499, n26500,
    n26501, n26502, n26503, n26504, n26505, n26506, n26507, n26508, n26509,
    n26510, n26511, n26512, n26513, n26514, n26515, n26516, n26517, n26518,
    n26519, n26520, n26521, n26522, n26523, n26524, n26525, n26526, n26527,
    n26528, n26529, n26530, n26532, n26533, n26534, n26535, n26536, n26537,
    n26538, n26539, n26540, n26541, n26542, n26543, n26544, n26545, n26546,
    n26547, n26548, n26549, n26550, n26551, n26552, n26553, n26554, n26555,
    n26556, n26557, n26558, n26559, n26560, n26561, n26562, n26563, n26564,
    n26565, n26566, n26568, n26569, n26570, n26571, n26572, n26573, n26574,
    n26575, n26576, n26577, n26578, n26579, n26580, n26581, n26582, n26583,
    n26584, n26585, n26586, n26587, n26588, n26589, n26590, n26591, n26592,
    n26593, n26594, n26595, n26596, n26597, n26598, n26599, n26600, n26601,
    n26602, n26603, n26604, n26605, n26606, n26607, n26608, n26609, n26610,
    n26611, n26612, n26613, n26614, n26615, n26616, n26617, n26618, n26619,
    n26620, n26621, n26622, n26623, n26624, n26625, n26626, n26627, n26628,
    n26629, n26630, n26631, n26632, n26633, n26634, n26635, n26636, n26637,
    n26638, n26639, n26640, n26641, n26642, n26643, n26644, n26645, n26646,
    n26647, n26648, n26649, n26650, n26651, n26652, n26653, n26654, n26655,
    n26656, n26657, n26658, n26659, n26660, n26661, n26662, n26663, n26664,
    n26665, n26666, n26667, n26668, n26669, n26671, n26672, n26673, n26674,
    n26675, n26676, n26677, n26678, n26679, n26680, n26681, n26682, n26683,
    n26684, n26685, n26686, n26687, n26688, n26689, n26690, n26691, n26692,
    n26693, n26694, n26695, n26696, n26697, n26698, n26699, n26700, n26701,
    n26702, n26703, n26704, n26705, n26706, n26707, n26708, n26709, n26710,
    n26711, n26712, n26713, n26714, n26715, n26716, n26717, n26718, n26719,
    n26720, n26721, n26722, n26723, n26724, n26725, n26726, n26727, n26728,
    n26729, n26730, n26731, n26732, n26733, n26734, n26735, n26736, n26737,
    n26738, n26739, n26740, n26741, n26742, n26743, n26744, n26745, n26746,
    n26747, n26748, n26749, n26750, n26751, n26752, n26753, n26754, n26755,
    n26756, n26757, n26758, n26759, n26760, n26761, n26762, n26763, n26764,
    n26765, n26766, n26767, n26768, n26769, n26770, n26772, n26773, n26774,
    n26775, n26776, n26777, n26778, n26779, n26780, n26781, n26782, n26783,
    n26784, n26785, n26786, n26787, n26788, n26789, n26790, n26791, n26792,
    n26793, n26794, n26795, n26796, n26797, n26798, n26799, n26800, n26801,
    n26802, n26803, n26804, n26805, n26806, n26807, n26808, n26809, n26810,
    n26811, n26812, n26813, n26814, n26815, n26816, n26818, n26819, n26820,
    n26821, n26822, n26823, n26824, n26825, n26826, n26827, n26828, n26829,
    n26830, n26831, n26832, n26833, n26834, n26835, n26836, n26837, n26838,
    n26839, n26840, n26841, n26842, n26843, n26844, n26845, n26846, n26847,
    n26848, n26849, n26850, n26851, n26852, n26853, n26854, n26855, n26856,
    n26857, n26858, n26859, n26860, n26861, n26862, n26863, n26864, n26865,
    n26866, n26867, n26868, n26869, n26870, n26871, n26872, n26873, n26874,
    n26875, n26876, n26877, n26878, n26879, n26880, n26881, n26882, n26883,
    n26884, n26885, n26886, n26887, n26888, n26889, n26890, n26891, n26892,
    n26893, n26894, n26895, n26896, n26897, n26898, n26899, n26900, n26901,
    n26902, n26903, n26904, n26905, n26906, n26907, n26908, n26909, n26910,
    n26911, n26912, n26913, n26914, n26915, n26916, n26917, n26918, n26919,
    n26921, n26922, n26923, n26924, n26925, n26926, n26927, n26928, n26929,
    n26930, n26931, n26932, n26933, n26934, n26935, n26936, n26937, n26938,
    n26939, n26940, n26941, n26942, n26943, n26944, n26945, n26946, n26947,
    n26948, n26949, n26950, n26951, n26952, n26954, n26955, n26956, n26957,
    n26958, n26959, n26960, n26961, n26962, n26963, n26964, n26965, n26966,
    n26967, n26968, n26969, n26970, n26971, n26972, n26973, n26974, n26975,
    n26976, n26977, n26978, n26979, n26980, n26981, n26982, n26983, n26984,
    n26985, n26987, n26988, n26989, n26990, n26991, n26992, n26993, n26994,
    n26995, n26996, n26997, n26998, n26999, n27000, n27001, n27002, n27003,
    n27004, n27005, n27006, n27007, n27008, n27009, n27010, n27011, n27012,
    n27013, n27014, n27015, n27016, n27017, n27018, n27019, n27020, n27021,
    n27022, n27023, n27024, n27025, n27026, n27027, n27028, n27029, n27030,
    n27031, n27032, n27033, n27034, n27035, n27036, n27037, n27038, n27039,
    n27040, n27041, n27042, n27043, n27044, n27045, n27046, n27047, n27048,
    n27049, n27050, n27051, n27052, n27053, n27054, n27055, n27056, n27057,
    n27058, n27059, n27060, n27061, n27062, n27063, n27064, n27065, n27066,
    n27067, n27068, n27069, n27070, n27071, n27072, n27073, n27074, n27075,
    n27076, n27077, n27078, n27079, n27080, n27081, n27082, n27083, n27084,
    n27085, n27086, n27087, n27088, n27089, n27090, n27091, n27092, n27094,
    n27095, n27096, n27097, n27098, n27099, n27100, n27101, n27102, n27103,
    n27104, n27105, n27106, n27107, n27108, n27109, n27110, n27111, n27112,
    n27113, n27114, n27115, n27116, n27117, n27118, n27119, n27120, n27121,
    n27122, n27123, n27124, n27125, n27126, n27127, n27128, n27129, n27130,
    n27131, n27132, n27133, n27134, n27135, n27136, n27137, n27138, n27139,
    n27140, n27141, n27142, n27143, n27144, n27145, n27146, n27147, n27148,
    n27149, n27150, n27151, n27152, n27153, n27154, n27155, n27156, n27157,
    n27158, n27159, n27160, n27161, n27162, n27163, n27164, n27165, n27166,
    n27167, n27168, n27169, n27170, n27171, n27172, n27173, n27174, n27175,
    n27176, n27177, n27178, n27179, n27180, n27181, n27182, n27183, n27184,
    n27185, n27186, n27187, n27188, n27189, n27190, n27191, n27192, n27193,
    n27194, n27195, n27197, n27198, n27199, n27200, n27201, n27202, n27203,
    n27204, n27205, n27206, n27207, n27208, n27209, n27210, n27211, n27212,
    n27213, n27214, n27215, n27216, n27217, n27218, n27219, n27220, n27221,
    n27222, n27223, n27224, n27225, n27226, n27227, n27228, n27229, n27230,
    n27231, n27232, n27233, n27234, n27236, n27237, n27238, n27239, n27240,
    n27241, n27242, n27243, n27244, n27245, n27246, n27247, n27248, n27249,
    n27250, n27251, n27252, n27253, n27254, n27255, n27256, n27257, n27258,
    n27259, n27260, n27261, n27262, n27263, n27264, n27265, n27266, n27267,
    n27268, n27269, n27270, n27271, n27272, n27273, n27275, n27276, n27277,
    n27278, n27279, n27280, n27281, n27282, n27283, n27284, n27285, n27286,
    n27287, n27288, n27289, n27290, n27291, n27292, n27293, n27294, n27295,
    n27296, n27297, n27298, n27299, n27300, n27301, n27302, n27303, n27304,
    n27305, n27306, n27307, n27308, n27309, n27311, n27312, n27313, n27314,
    n27315, n27316, n27317, n27318, n27319, n27320, n27321, n27322, n27323,
    n27324, n27325, n27326, n27327, n27328, n27329, n27330, n27331, n27332,
    n27333, n27334, n27335, n27336, n27337, n27338, n27339, n27340, n27341,
    n27342, n27343, n27344, n27345, n27346, n27347, n27348, n27349, n27350,
    n27351, n27352, n27353, n27354, n27355, n27356, n27357, n27358, n27359,
    n27360, n27361, n27362, n27363, n27364, n27365, n27366, n27367, n27368,
    n27369, n27370, n27371, n27372, n27373, n27374, n27375, n27376, n27377,
    n27378, n27379, n27380, n27381, n27382, n27383, n27384, n27385, n27386,
    n27387, n27388, n27389, n27390, n27391, n27392, n27393, n27394, n27395,
    n27396, n27397, n27398, n27399, n27400, n27401, n27402, n27403, n27404,
    n27405, n27407, n27408, n27409, n27410, n27411, n27412, n27413, n27414,
    n27415, n27416, n27417, n27418, n27419, n27420, n27421, n27422, n27423,
    n27424, n27425, n27426, n27427, n27428, n27429, n27430, n27431, n27432,
    n27433, n27434, n27435, n27436, n27437, n27438, n27439, n27440, n27441,
    n27442, n27443, n27444, n27445, n27446, n27447, n27448, n27449, n27450,
    n27451, n27452, n27453, n27454, n27455, n27457, n27458, n27459, n27460,
    n27461, n27462, n27463, n27464, n27465, n27466, n27467, n27468, n27469,
    n27470, n27471, n27472, n27473, n27474, n27475, n27476, n27477, n27478,
    n27479, n27480, n27481, n27482, n27483, n27484, n27485, n27486, n27487,
    n27488, n27489, n27490, n27491, n27492, n27493, n27494, n27495, n27496,
    n27497, n27499, n27500, n27501, n27502, n27503, n27504, n27505, n27506,
    n27507, n27508, n27509, n27510, n27511, n27512, n27513, n27514, n27515,
    n27516, n27517, n27518, n27519, n27520, n27521, n27522, n27523, n27524,
    n27525, n27526, n27527, n27528, n27529, n27530, n27531, n27532, n27533,
    n27534, n27535, n27536, n27537, n27538, n27539, n27540, n27542, n27543,
    n27544, n27545, n27546, n27547, n27548, n27549, n27550, n27551, n27552,
    n27553, n27554, n27555, n27556, n27557, n27558, n27559, n27560, n27561,
    n27562, n27563, n27564, n27565, n27566, n27567, n27568, n27569, n27570,
    n27571, n27572, n27573, n27574, n27575, n27576, n27577, n27578, n27579,
    n27580, n27581, n27583, n27584, n27585, n27586, n27587, n27588, n27589,
    n27590, n27591, n27592, n27593, n27594, n27595, n27596, n27597, n27598,
    n27599, n27600, n27601, n27602, n27603, n27604, n27605, n27606, n27607,
    n27608, n27609, n27610, n27611, n27612, n27613, n27614, n27615, n27616,
    n27617, n27618, n27619, n27620, n27621, n27622, n27623, n27624, n27625,
    n27626, n27627, n27628, n27629, n27630, n27631, n27632, n27633, n27634,
    n27635, n27636, n27637, n27638, n27639, n27640, n27641, n27642, n27643,
    n27644, n27645, n27646, n27647, n27648, n27649, n27650, n27651, n27652,
    n27653, n27654, n27655, n27656, n27657, n27658, n27659, n27660, n27661,
    n27662, n27663, n27664, n27665, n27666, n27667, n27668, n27669, n27670,
    n27671, n27672, n27674, n27675, n27676, n27677, n27678, n27679, n27680,
    n27681, n27682, n27683, n27684, n27685, n27686, n27687, n27688, n27689,
    n27690, n27691, n27692, n27693, n27694, n27695, n27696, n27697, n27698,
    n27699, n27700, n27701, n27702, n27703, n27704, n27705, n27706, n27707,
    n27708, n27709, n27710, n27711, n27712, n27713, n27714, n27716, n27717,
    n27718, n27719, n27720, n27721, n27722, n27723, n27724, n27725, n27726,
    n27727, n27728, n27729, n27730, n27731, n27732, n27733, n27734, n27735,
    n27736, n27737, n27738, n27739, n27740, n27741, n27742, n27743, n27744,
    n27745, n27746, n27747, n27748, n27749, n27750, n27751, n27752, n27753,
    n27754, n27756, n27757, n27758, n27759, n27760, n27761, n27762, n27763,
    n27764, n27765, n27766, n27767, n27768, n27769, n27770, n27771, n27772,
    n27773, n27774, n27775, n27776, n27777, n27778, n27779, n27780, n27781,
    n27782, n27783, n27784, n27785, n27786, n27787, n27788, n27789, n27790,
    n27791, n27792, n27793, n27794, n27795, n27796, n27797, n27798, n27799,
    n27800, n27801, n27802, n27803, n27804, n27805, n27806, n27807, n27808,
    n27809, n27810, n27811, n27812, n27813, n27814, n27815, n27816, n27817,
    n27818, n27819, n27820, n27821, n27822, n27823, n27824, n27825, n27826,
    n27827, n27828, n27829, n27830, n27831, n27832, n27833, n27834, n27835,
    n27836, n27837, n27838, n27839, n27840, n27841, n27842, n27843, n27844,
    n27845, n27846, n27847, n27848, n27849, n27850, n27852, n27853, n27854,
    n27855, n27856, n27857, n27858, n27859, n27860, n27861, n27862, n27863,
    n27864, n27865, n27866, n27867, n27868, n27869, n27870, n27871, n27872,
    n27873, n27874, n27875, n27876, n27877, n27878, n27879, n27880, n27881,
    n27882, n27883, n27884, n27885, n27886, n27887, n27888, n27889, n27890,
    n27892, n27893, n27894, n27895, n27896, n27897, n27898, n27899, n27900,
    n27901, n27902, n27903, n27904, n27905, n27906, n27907, n27908, n27909,
    n27910, n27911, n27912, n27913, n27914, n27915, n27916, n27917, n27918,
    n27919, n27920, n27921, n27922, n27923, n27924, n27925, n27926, n27927,
    n27928, n27929, n27930, n27931, n27932, n27933, n27934, n27935, n27937,
    n27938, n27939, n27940, n27941, n27942, n27943, n27944, n27945, n27946,
    n27947, n27948, n27949, n27950, n27951, n27952, n27953, n27954, n27955,
    n27956, n27957, n27958, n27959, n27960, n27961, n27962, n27963, n27964,
    n27965, n27966, n27967, n27968, n27969, n27970, n27971, n27972, n27973,
    n27975, n27976, n27977, n27978, n27979, n27980, n27981, n27982, n27983,
    n27984, n27985, n27986, n27987, n27988, n27989, n27990, n27991, n27992,
    n27993, n27994, n27995, n27996, n27997, n27998, n27999, n28000, n28001,
    n28002, n28003, n28004, n28005, n28006, n28007, n28008, n28009, n28010,
    n28011, n28012, n28013, n28014, n28015, n28016, n28017, n28018, n28019,
    n28020, n28021, n28022, n28023, n28024, n28025, n28027, n28028, n28029,
    n28030, n28031, n28032, n28033, n28034, n28035, n28036, n28037, n28038,
    n28039, n28040, n28041, n28042, n28043, n28044, n28045, n28046, n28047,
    n28048, n28049, n28050, n28051, n28052, n28053, n28054, n28055, n28056,
    n28057, n28058, n28059, n28060, n28061, n28062, n28063, n28064, n28066,
    n28067, n28068, n28069, n28070, n28071, n28072, n28073, n28074, n28075,
    n28076, n28077, n28078, n28079, n28080, n28081, n28082, n28083, n28084,
    n28085, n28086, n28087, n28088, n28089, n28090, n28091, n28092, n28093,
    n28094, n28095, n28096, n28097, n28098, n28099, n28100, n28102, n28103,
    n28104, n28105, n28106, n28107, n28108, n28109, n28110, n28111, n28112,
    n28113, n28114, n28115, n28116, n28117, n28118, n28119, n28120, n28121,
    n28122, n28123, n28124, n28125, n28126, n28127, n28128, n28129, n28130,
    n28131, n28132, n28133, n28134, n28135, n28136, n28137, n28139, n28140,
    n28141, n28142, n28143, n28144, n28145, n28146, n28147, n28148, n28149,
    n28150, n28151, n28152, n28153, n28154, n28155, n28156, n28157, n28158,
    n28159, n28160, n28161, n28162, n28163, n28164, n28165, n28166, n28167,
    n28168, n28169, n28170, n28171, n28172, n28173, n28175, n28176, n28177,
    n28178, n28179, n28180, n28181, n28182, n28183, n28184, n28185, n28186,
    n28187, n28188, n28189, n28190, n28191, n28192, n28193, n28194, n28195,
    n28196, n28197, n28198, n28199, n28200, n28201, n28202, n28203, n28205,
    n28206, n28207, n28208, n28209, n28210, n28211, n28212, n28213, n28214,
    n28215, n28216, n28217, n28218, n28219, n28220, n28221, n28222, n28223,
    n28224, n28225, n28226, n28227, n28228, n28229, n28230, n28231, n28232,
    n28233, n28234, n28236, n28237, n28238, n28239, n28240, n28241, n28242,
    n28243, n28244, n28245, n28246, n28247, n28248, n28249, n28250, n28251,
    n28252, n28253, n28254, n28255, n28256, n28257, n28258, n28259, n28260,
    n28261, n28262, n28263, n28264, n28265, n28266, n28267, n28268, n28269,
    n28270, n28272, n28273, n28274, n28275, n28276, n28277, n28278, n28279,
    n28280, n28281, n28282, n28283, n28284, n28285, n28286, n28287, n28288,
    n28289, n28290, n28291, n28292, n28293, n28294, n28295, n28296, n28297,
    n28298, n28300, n28301, n28302, n28303, n28304, n28305, n28306, n28307,
    n28308, n28309, n28310, n28311, n28312, n28313, n28314, n28315, n28316,
    n28317, n28318, n28319, n28320, n28321, n28322, n28323, n28324, n28325,
    n28326, n28327, n28328, n28329, n28330, n28331, n28332, n28333, n28334,
    n28335, n28336, n28337, n28338, n28339, n28340, n28341, n28342, n28343,
    n28344, n28345, n28346, n28347, n28348, n28349, n28350, n28351, n28352,
    n28353, n28354, n28355, n28356, n28357, n28358, n28359, n28360, n28361,
    n28362, n28363, n28364, n28365, n28366, n28367, n28368, n28369, n28370,
    n28371, n28372, n28373, n28374, n28375, n28376, n28377, n28378, n28379,
    n28380, n28381, n28382, n28383, n28384, n28385, n28386, n28387, n28388,
    n28389, n28390, n28391, n28392, n28393, n28394, n28395, n28396, n28397,
    n28398, n28399, n28401, n28402, n28403, n28404, n28405, n28406, n28407,
    n28408, n28409, n28410, n28411, n28412, n28413, n28414, n28415, n28416,
    n28417, n28418, n28419, n28420, n28421, n28422, n28423, n28424, n28425,
    n28426, n28427, n28428, n28429, n28430, n28431, n28432, n28433, n28434,
    n28435, n28436, n28437, n28438, n28439, n28440, n28441, n28442, n28443,
    n28444, n28445, n28446, n28447, n28448, n28449, n28450, n28451, n28452,
    n28453, n28454, n28455, n28456, n28457, n28458, n28459, n28460, n28461,
    n28462, n28463, n28464, n28465, n28466, n28467, n28468, n28469, n28470,
    n28471, n28472, n28473, n28474, n28475, n28476, n28477, n28478, n28479,
    n28480, n28481, n28482, n28483, n28484, n28485, n28486, n28487, n28488,
    n28489, n28490, n28491, n28492, n28493, n28494, n28495, n28496, n28497,
    n28498, n28499, n28500, n28502, n28503, n28504, n28505, n28506, n28507,
    n28508, n28509, n28510, n28511, n28512, n28513, n28514, n28515, n28516,
    n28517, n28518, n28519, n28520, n28521, n28522, n28523, n28524, n28525,
    n28526, n28527, n28528, n28529, n28530, n28531, n28532, n28533, n28534,
    n28535, n28536, n28537, n28538, n28539, n28540, n28541, n28542, n28543,
    n28544, n28545, n28546, n28547, n28548, n28549, n28550, n28551, n28552,
    n28553, n28554, n28555, n28556, n28557, n28558, n28559, n28560, n28561,
    n28562, n28563, n28564, n28565, n28566, n28567, n28568, n28569, n28570,
    n28571, n28572, n28573, n28574, n28575, n28576, n28577, n28578, n28579,
    n28580, n28581, n28582, n28583, n28584, n28585, n28586, n28587, n28588,
    n28589, n28590, n28591, n28592, n28593, n28594, n28595, n28596, n28597,
    n28598, n28599, n28601, n28602, n28603, n28604, n28605, n28606, n28607,
    n28608, n28609, n28610, n28611, n28612, n28613, n28614, n28615, n28616,
    n28617, n28618, n28619, n28620, n28621, n28622, n28623, n28624, n28625,
    n28626, n28627, n28628, n28629, n28630, n28631, n28632, n28633, n28634,
    n28635, n28636, n28637, n28638, n28639, n28640, n28641, n28642, n28643,
    n28644, n28645, n28646, n28647, n28648, n28649, n28650, n28651, n28652,
    n28653, n28654, n28655, n28656, n28657, n28658, n28659, n28660, n28661,
    n28662, n28663, n28664, n28665, n28666, n28667, n28668, n28669, n28670,
    n28671, n28672, n28673, n28674, n28675, n28676, n28677, n28678, n28679,
    n28680, n28681, n28682, n28683, n28684, n28685, n28686, n28687, n28688,
    n28689, n28690, n28691, n28692, n28693, n28694, n28695, n28696, n28697,
    n28698, n28699, n28700, n28701, n28702, n28704, n28705, n28706, n28707,
    n28708, n28709, n28710, n28711, n28712, n28713, n28714, n28715, n28716,
    n28717, n28718, n28719, n28720, n28721, n28722, n28723, n28724, n28725,
    n28726, n28727, n28728, n28729, n28730, n28731, n28732, n28733, n28734,
    n28735, n28736, n28737, n28738, n28739, n28740, n28741, n28742, n28743,
    n28744, n28745, n28747, n28748, n28749, n28750, n28751, n28752, n28753,
    n28754, n28755, n28756, n28757, n28758, n28759, n28760, n28761, n28762,
    n28763, n28764, n28765, n28766, n28767, n28768, n28769, n28770, n28771,
    n28772, n28773, n28774, n28775, n28776, n28777, n28778, n28779, n28780,
    n28781, n28782, n28783, n28784, n28785, n28786, n28787, n28788, n28789,
    n28790, n28791, n28792, n28793, n28794, n28795, n28796, n28797, n28798,
    n28799, n28800, n28801, n28802, n28803, n28804, n28805, n28806, n28807,
    n28808, n28809, n28810, n28811, n28812, n28813, n28814, n28815, n28816,
    n28817, n28818, n28819, n28820, n28821, n28822, n28823, n28824, n28825,
    n28826, n28827, n28828, n28829, n28830, n28831, n28832, n28833, n28834,
    n28835, n28836, n28837, n28838, n28839, n28840, n28841, n28842, n28843,
    n28844, n28845, n28846, n28847, n28848, n28849, n28850, n28852, n28853,
    n28854, n28855, n28856, n28857, n28858, n28859, n28860, n28861, n28862,
    n28863, n28864, n28865, n28866, n28867, n28868, n28869, n28870, n28871,
    n28872, n28873, n28874, n28875, n28876, n28877, n28878, n28879, n28880,
    n28881, n28882, n28883, n28884, n28885, n28886, n28887, n28888, n28889,
    n28890, n28891, n28892, n28893, n28894, n28895, n28896, n28898, n28899,
    n28900, n28901, n28902, n28903, n28904, n28905, n28906, n28907, n28908,
    n28909, n28910, n28911, n28912, n28913, n28914, n28915, n28916, n28917,
    n28918, n28919, n28920, n28921, n28922, n28923, n28924, n28925, n28926,
    n28927, n28928, n28929, n28930, n28931, n28932, n28933, n28934, n28935,
    n28936, n28937, n28938, n28939, n28940, n28941, n28942, n28943, n28944,
    n28945, n28946, n28947, n28948, n28949, n28950, n28951, n28952, n28953,
    n28954, n28955, n28956, n28957, n28958, n28959, n28960, n28961, n28962,
    n28963, n28964, n28965, n28966, n28967, n28968, n28969, n28970, n28971,
    n28972, n28973, n28974, n28975, n28976, n28977, n28978, n28979, n28980,
    n28981, n28982, n28983, n28984, n28985, n28986, n28987, n28988, n28990,
    n28991, n28992, n28993, n28994, n28995, n28996, n28997, n28998, n28999,
    n29000, n29001, n29002, n29003, n29004, n29005, n29006, n29007, n29008,
    n29009, n29010, n29011, n29012, n29013, n29014, n29015, n29016, n29017,
    n29018, n29019, n29020, n29021, n29022, n29023, n29024, n29025, n29026,
    n29027, n29028, n29029, n29030, n29031, n29032, n29033, n29034, n29035,
    n29036, n29038, n29039, n29040, n29041, n29042, n29043, n29044, n29045,
    n29046, n29047, n29048, n29049, n29050, n29051, n29052, n29053, n29054,
    n29055, n29056, n29057, n29058, n29059, n29060, n29061, n29062, n29063,
    n29064, n29065, n29066, n29067, n29068, n29069, n29070, n29071, n29072,
    n29073, n29074, n29075, n29076, n29077, n29078, n29079, n29080, n29081,
    n29082, n29083, n29084, n29085, n29086, n29087, n29088, n29089, n29091,
    n29092, n29093, n29094, n29095, n29096, n29097, n29098, n29099, n29100,
    n29101, n29102, n29103, n29104, n29105, n29106, n29107, n29108, n29109,
    n29110, n29111, n29112, n29113, n29114, n29115, n29116, n29117, n29118,
    n29119, n29120, n29121, n29122, n29124, n29125, n29126, n29127, n29128,
    n29129, n29130, n29131, n29132, n29133, n29134, n29135, n29136, n29137,
    n29138, n29139, n29140, n29141, n29142, n29143, n29144, n29145, n29146,
    n29147, n29148, n29149, n29150, n29151, n29152, n29153, n29154, n29155,
    n29156, n29157, n29158, n29159, n29160, n29161, n29162, n29163, n29164,
    n29165, n29166, n29167, n29168, n29169, n29171, n29172, n29173, n29174,
    n29175, n29176, n29177, n29178, n29179, n29180, n29181, n29182, n29183,
    n29184, n29185, n29186, n29187, n29188, n29189, n29190, n29191, n29192,
    n29193, n29194, n29195, n29196, n29197, n29198, n29199, n29200, n29201,
    n29203, n29204, n29205, n29206, n29207, n29208, n29209, n29210, n29211,
    n29212, n29213, n29214, n29215, n29216, n29217, n29218, n29219, n29220,
    n29221, n29222, n29223, n29224, n29225, n29226, n29227, n29228, n29229,
    n29230, n29231, n29232, n29233, n29234, n29236, n29237, n29238, n29239,
    n29240, n29241, n29242, n29243, n29244, n29245, n29246, n29247, n29248,
    n29249, n29250, n29251, n29252, n29253, n29254, n29255, n29256, n29257,
    n29258, n29259, n29260, n29261, n29262, n29263, n29264, n29265, n29266,
    n29267, n29268, n29269, n29270, n29271, n29272, n29273, n29274, n29275,
    n29276, n29277, n29278, n29279, n29280, n29282, n29283, n29284, n29285,
    n29286, n29287, n29288, n29289, n29290, n29291, n29292, n29293, n29294,
    n29295, n29296, n29297, n29298, n29299, n29300, n29301, n29302, n29303,
    n29304, n29305, n29306, n29307, n29308, n29309, n29310, n29311, n29312,
    n29313, n29314, n29315, n29316, n29317, n29318, n29319, n29320, n29321,
    n29322, n29323, n29324, n29325, n29326, n29327, n29328, n29329, n29330,
    n29331, n29332, n29333, n29334, n29335, n29336, n29337, n29338, n29339,
    n29340, n29341, n29342, n29343, n29344, n29345, n29346, n29347, n29348,
    n29349, n29350, n29351, n29352, n29353, n29354, n29355, n29356, n29357,
    n29358, n29359, n29360, n29361, n29362, n29363, n29364, n29365, n29366,
    n29367, n29368, n29369, n29370, n29371, n29372, n29373, n29374, n29375,
    n29376, n29377, n29378, n29379, n29381, n29382, n29383, n29384, n29385,
    n29386, n29387, n29388, n29389, n29390, n29391, n29392, n29393, n29394,
    n29395, n29396, n29397, n29398, n29399, n29400, n29401, n29402, n29403,
    n29404, n29405, n29406, n29407, n29408, n29409, n29410, n29411, n29412,
    n29413, n29414, n29415, n29416, n29417, n29418, n29419, n29420, n29421,
    n29422, n29423, n29424, n29426, n29427, n29428, n29429, n29430, n29431,
    n29432, n29433, n29434, n29435, n29436, n29437, n29438, n29439, n29440,
    n29441, n29442, n29443, n29444, n29445, n29446, n29447, n29448, n29449,
    n29450, n29451, n29452, n29453, n29454, n29455, n29456, n29457, n29458,
    n29459, n29460, n29461, n29463, n29464, n29465, n29466, n29467, n29468,
    n29469, n29470, n29471, n29472, n29473, n29474, n29475, n29476, n29477,
    n29478, n29479, n29480, n29481, n29482, n29483, n29484, n29485, n29486,
    n29487, n29488, n29489, n29490, n29491, n29492, n29493, n29494, n29495,
    n29496, n29497, n29498, n29499, n29500, n29501, n29502, n29503, n29504,
    n29505, n29506, n29507, n29508, n29509, n29510, n29511, n29512, n29513,
    n29514, n29515, n29516, n29517, n29518, n29519, n29520, n29521, n29522,
    n29523, n29524, n29525, n29526, n29527, n29528, n29529, n29530, n29531,
    n29532, n29533, n29534, n29535, n29536, n29537, n29538, n29539, n29540,
    n29541, n29542, n29543, n29544, n29545, n29546, n29547, n29548, n29549,
    n29550, n29551, n29552, n29553, n29554, n29555, n29556, n29557, n29558,
    n29559, n29560, n29561, n29562, n29563, n29564, n29565, n29566, n29567,
    n29568, n29570, n29571, n29572, n29573, n29574, n29575, n29576, n29577,
    n29578, n29579, n29580, n29581, n29582, n29583, n29584, n29585, n29586,
    n29587, n29588, n29589, n29590, n29591, n29592, n29593, n29594, n29595,
    n29596, n29597, n29598, n29599, n29600, n29601, n29602, n29603, n29604,
    n29605, n29606, n29607, n29609, n29610, n29611, n29612, n29613, n29614,
    n29615, n29616, n29617, n29618, n29619, n29620, n29621, n29622, n29623,
    n29624, n29625, n29626, n29627, n29628, n29629, n29630, n29631, n29632,
    n29633, n29634, n29635, n29636, n29637, n29638, n29639, n29640, n29641,
    n29642, n29643, n29645, n29646, n29647, n29648, n29649, n29650, n29651,
    n29652, n29653, n29654, n29655, n29656, n29657, n29658, n29659, n29660,
    n29661, n29662, n29663, n29664, n29665, n29666, n29667, n29668, n29669,
    n29670, n29671, n29672, n29673, n29674, n29675, n29676, n29677, n29678,
    n29679, n29680, n29682, n29683, n29684, n29685, n29686, n29687, n29688,
    n29689, n29690, n29691, n29692, n29693, n29694, n29695, n29696, n29697,
    n29698, n29699, n29700, n29701, n29702, n29703, n29704, n29705, n29706,
    n29707, n29708, n29709, n29710, n29711, n29712, n29713, n29714, n29715,
    n29716, n29717, n29719, n29720, n29721, n29722, n29723, n29724, n29725,
    n29726, n29727, n29728, n29729, n29730, n29731, n29732, n29733, n29734,
    n29735, n29736, n29737, n29738, n29739, n29740, n29741, n29742, n29743,
    n29744, n29745, n29746, n29747, n29749, n29750, n29751, n29752, n29753,
    n29754, n29755, n29756, n29757, n29758, n29759, n29760, n29761, n29762,
    n29763, n29764, n29765, n29766, n29767, n29768, n29769, n29770, n29771,
    n29772, n29773, n29774, n29775, n29776, n29777, n29778, n29779, n29780,
    n29781, n29783, n29784, n29785, n29786, n29787, n29788, n29789, n29790,
    n29791, n29792, n29793, n29794, n29795, n29796, n29797, n29798, n29799,
    n29800, n29801, n29802, n29803, n29804, n29805, n29806, n29807, n29808,
    n29809, n29810, n29811, n29812, n29813, n29814, n29815, n29816, n29817,
    n29818, n29819, n29820, n29822, n29823, n29824, n29825, n29826, n29827,
    n29828, n29829, n29830, n29831, n29832, n29833, n29834, n29835, n29836,
    n29837, n29838, n29839, n29840, n29841, n29842, n29843, n29844, n29845,
    n29846, n29847, n29848, n29849, n29850, n29851, n29852, n29853, n29854,
    n29855, n29856, n29858, n29859, n29860, n29861, n29862, n29863, n29864,
    n29865, n29866, n29867, n29868, n29869, n29870, n29871, n29872, n29873,
    n29874, n29875, n29876, n29877, n29878, n29879, n29880, n29881, n29882,
    n29883, n29884, n29885, n29886, n29887, n29888, n29889, n29890, n29891,
    n29892, n29893, n29894, n29895, n29897, n29898, n29899, n29900, n29901,
    n29902, n29903, n29904, n29905, n29906, n29907, n29908, n29909, n29910,
    n29911, n29912, n29913, n29914, n29915, n29916, n29917, n29918, n29919,
    n29920, n29921, n29922, n29923, n29924, n29925, n29926, n29927, n29928,
    n29929, n29930, n29931, n29932, n29933, n29934, n29935, n29937, n29938,
    n29939, n29940, n29941, n29942, n29943, n29944, n29945, n29946, n29947,
    n29948, n29949, n29950, n29951, n29952, n29953, n29954, n29955, n29956,
    n29957, n29958, n29959, n29960, n29961, n29962, n29963, n29964, n29965,
    n29966, n29968, n29969, n29970, n29971, n29972, n29973, n29974, n29975,
    n29976, n29977, n29978, n29979, n29980, n29981, n29982, n29983, n29984,
    n29985, n29986, n29987, n29988, n29989, n29990, n29991, n29992, n29993,
    n29994, n29996, n29997, n29998, n29999, n30000, n30001, n30002, n30003,
    n30004, n30005, n30006, n30007, n30008, n30009, n30010, n30011, n30012,
    n30013, n30014, n30015, n30016, n30017, n30018, n30019, n30020, n30021,
    n30022, n30023, n30024, n30025, n30026, n30027, n30028, n30029, n30030,
    n30032, n30033, n30034, n30035, n30036, n30037, n30038, n30039, n30040,
    n30041, n30042, n30043, n30044, n30045, n30046, n30047, n30048, n30049,
    n30050, n30051, n30052, n30053, n30054, n30055, n30056, n30057, n30058,
    n30059, n30060, n30061, n30062, n30063, n30064, n30065, n30066, n30067,
    n30068, n30069, n30070, n30071, n30072, n30073, n30074, n30075, n30076,
    n30077, n30078, n30079, n30080, n30081, n30082, n30083, n30084, n30085,
    n30086, n30087, n30088, n30089, n30090, n30091, n30092, n30093, n30094,
    n30095, n30096, n30097, n30098, n30099, n30100, n30101, n30102, n30103,
    n30104, n30105, n30106, n30107, n30108, n30109, n30110, n30111, n30112,
    n30113, n30114, n30115, n30116, n30117, n30118, n30119, n30120, n30121,
    n30122, n30123, n30124, n30125, n30126, n30127, n30128, n30129, n30130,
    n30131, n30132, n30133, n30134, n30135, n30137, n30138, n30139, n30140,
    n30141, n30142, n30143, n30144, n30145, n30146, n30147, n30148, n30149,
    n30150, n30151, n30152, n30153, n30154, n30155, n30156, n30157, n30158,
    n30159, n30160, n30161, n30162, n30163, n30164, n30165, n30166, n30167,
    n30168, n30169, n30170, n30171, n30172, n30173, n30174, n30175, n30176,
    n30178, n30179, n30180, n30181, n30182, n30183, n30184, n30185, n30186,
    n30187, n30188, n30189, n30190, n30191, n30192, n30193, n30194, n30195,
    n30196, n30197, n30198, n30199, n30200, n30201, n30202, n30203, n30204,
    n30205, n30206, n30207, n30208, n30209, n30210, n30211, n30212, n30213,
    n30214, n30215, n30216, n30217, n30218, n30219, n30220, n30221, n30222,
    n30223, n30224, n30225, n30226, n30227, n30228, n30229, n30230, n30231,
    n30232, n30233, n30234, n30235, n30236, n30237, n30238, n30239, n30240,
    n30241, n30242, n30243, n30244, n30245, n30246, n30247, n30248, n30249,
    n30250, n30251, n30252, n30253, n30254, n30255, n30256, n30257, n30258,
    n30259, n30260, n30261, n30262, n30263, n30264, n30265, n30266, n30267,
    n30269, n30270, n30271, n30272, n30273, n30274, n30275, n30276, n30277,
    n30278, n30279, n30280, n30281, n30282, n30283, n30284, n30285, n30286,
    n30287, n30288, n30289, n30290, n30291, n30292, n30293, n30294, n30295,
    n30296, n30297, n30298, n30299, n30300, n30301, n30302, n30303, n30304,
    n30305, n30306, n30307, n30308, n30309, n30310, n30311, n30312, n30313,
    n30314, n30315, n30316, n30317, n30318, n30319, n30320, n30321, n30322,
    n30323, n30324, n30325, n30326, n30327, n30328, n30329, n30330, n30331,
    n30332, n30333, n30334, n30335, n30336, n30337, n30338, n30339, n30340,
    n30341, n30342, n30343, n30344, n30345, n30346, n30347, n30348, n30349,
    n30350, n30351, n30352, n30353, n30354, n30355, n30356, n30357, n30358,
    n30359, n30360, n30361, n30362, n30363, n30364, n30365, n30366, n30367,
    n30368, n30369, n30370, n30371, n30372, n30374, n30375, n30376, n30377,
    n30378, n30379, n30380, n30381, n30382, n30383, n30384, n30385, n30386,
    n30387, n30388, n30389, n30390, n30391, n30392, n30393, n30394, n30395,
    n30396, n30397, n30398, n30399, n30400, n30401, n30402, n30403, n30404,
    n30405, n30406, n30407, n30408, n30409, n30410, n30411, n30412, n30413,
    n30414, n30415, n30416, n30417, n30418, n30419, n30420, n30421, n30422,
    n30423, n30424, n30425, n30426, n30427, n30428, n30429, n30430, n30431,
    n30432, n30433, n30434, n30435, n30436, n30437, n30438, n30439, n30440,
    n30441, n30442, n30443, n30444, n30445, n30446, n30447, n30448, n30449,
    n30450, n30451, n30452, n30453, n30454, n30455, n30456, n30457, n30458,
    n30459, n30460, n30461, n30462, n30463, n30464, n30465, n30466, n30467,
    n30468, n30469, n30470, n30471, n30472, n30473, n30474, n30476, n30477,
    n30478, n30479, n30480, n30481, n30482, n30483, n30484, n30485, n30486,
    n30487, n30488, n30489, n30490, n30491, n30492, n30493, n30494, n30495,
    n30496, n30497, n30498, n30499, n30500, n30501, n30502, n30503, n30504,
    n30505, n30506, n30507, n30508, n30509, n30510, n30511, n30512, n30513,
    n30514, n30515, n30517, n30518, n30519, n30520, n30521, n30522, n30523,
    n30524, n30525, n30526, n30527, n30528, n30529, n30530, n30531, n30532,
    n30533, n30534, n30535, n30536, n30537, n30538, n30539, n30540, n30541,
    n30542, n30543, n30544, n30545, n30546, n30547, n30548, n30549, n30550,
    n30551, n30552, n30553, n30554, n30555, n30556, n30557, n30558, n30559,
    n30560, n30561, n30562, n30563, n30564, n30565, n30566, n30567, n30569,
    n30570, n30571, n30572, n30573, n30574, n30575, n30576, n30577, n30578,
    n30579, n30580, n30581, n30582, n30583, n30584, n30585, n30586, n30587,
    n30588, n30589, n30590, n30591, n30592, n30593, n30594, n30595, n30596,
    n30597, n30598, n30599, n30600, n30601, n30602, n30603, n30604, n30605,
    n30606, n30607, n30609, n30610, n30611, n30612, n30613, n30614, n30615,
    n30616, n30617, n30618, n30619, n30620, n30621, n30622, n30623, n30624,
    n30625, n30626, n30627, n30628, n30629, n30630, n30631, n30632, n30633,
    n30634, n30635, n30636, n30637, n30638, n30640, n30641, n30642, n30643,
    n30644, n30645, n30646, n30647, n30648, n30649, n30650, n30651, n30652,
    n30653, n30654, n30655, n30656, n30657, n30658, n30659, n30660, n30661,
    n30662, n30663, n30664, n30665, n30666, n30667, n30668, n30669, n30670,
    n30671, n30672, n30673, n30674, n30675, n30676, n30677, n30678, n30679,
    n30680, n30681, n30682, n30683, n30684, n30685, n30686, n30687, n30688,
    n30689, n30690, n30691, n30692, n30693, n30694, n30695, n30696, n30697,
    n30698, n30699, n30700, n30701, n30702, n30703, n30704, n30705, n30706,
    n30707, n30708, n30709, n30710, n30711, n30712, n30713, n30714, n30715,
    n30716, n30717, n30718, n30719, n30720, n30721, n30722, n30723, n30724,
    n30725, n30726, n30727, n30728, n30729, n30730, n30731, n30732, n30733,
    n30734, n30735, n30736, n30737, n30738, n30739, n30740, n30741, n30743,
    n30744, n30745, n30746, n30747, n30748, n30749, n30750, n30751, n30752,
    n30753, n30754, n30755, n30756, n30757, n30758, n30759, n30760, n30761,
    n30762, n30763, n30764, n30765, n30766, n30767, n30768, n30769, n30770,
    n30771, n30772, n30773, n30774, n30775, n30776, n30777, n30778, n30779,
    n30780, n30781, n30782, n30783, n30784, n30785, n30786, n30787, n30788,
    n30789, n30790, n30791, n30792, n30793, n30794, n30795, n30796, n30797,
    n30798, n30799, n30800, n30801, n30802, n30803, n30804, n30805, n30806,
    n30807, n30808, n30809, n30810, n30811, n30812, n30813, n30814, n30815,
    n30816, n30817, n30818, n30819, n30820, n30821, n30822, n30823, n30824,
    n30825, n30826, n30827, n30828, n30829, n30830, n30831, n30832, n30833,
    n30834, n30835, n30836, n30837, n30838, n30839, n30840, n30841, n30842,
    n30844, n30845, n30846, n30847, n30848, n30849, n30850, n30851, n30852,
    n30853, n30854, n30855, n30856, n30857, n30858, n30859, n30860, n30861,
    n30862, n30863, n30864, n30865, n30866, n30867, n30868, n30869, n30870,
    n30871, n30872, n30873, n30874, n30876, n30877, n30878, n30879, n30880,
    n30881, n30882, n30883, n30884, n30885, n30886, n30887, n30888, n30889,
    n30890, n30891, n30892, n30893, n30894, n30895, n30896, n30897, n30898,
    n30899, n30900, n30901, n30902, n30903, n30904, n30905, n30906, n30907,
    n30908, n30909, n30910, n30911, n30912, n30913, n30914, n30915, n30917,
    n30918, n30919, n30920, n30921, n30922, n30923, n30924, n30925, n30926,
    n30927, n30928, n30929, n30930, n30931, n30932, n30933, n30934, n30935,
    n30936, n30937, n30938, n30939, n30940, n30941, n30942, n30943, n30944,
    n30945, n30946, n30947, n30948, n30949, n30950, n30951, n30952, n30953,
    n30954, n30955, n30956, n30957, n30958, n30959, n30960, n30961, n30962,
    n30963, n30964, n30965, n30966, n30967, n30968, n30969, n30970, n30971,
    n30972, n30973, n30974, n30975, n30976, n30977, n30978, n30979, n30980,
    n30981, n30982, n30983, n30984, n30985, n30986, n30987, n30988, n30989,
    n30990, n30991, n30992, n30993, n30994, n30995, n30996, n30997, n30998,
    n30999, n31000, n31001, n31002, n31003, n31004, n31005, n31006, n31007,
    n31008, n31009, n31010, n31011, n31012, n31014, n31015, n31016, n31017,
    n31018, n31019, n31020, n31021, n31022, n31023, n31024, n31025, n31026,
    n31027, n31028, n31029, n31030, n31031, n31032, n31033, n31034, n31035,
    n31036, n31037, n31038, n31039, n31040, n31041, n31042, n31043, n31044,
    n31045, n31046, n31047, n31048, n31049, n31050, n31051, n31052, n31053,
    n31054, n31055, n31056, n31057, n31058, n31059, n31060, n31061, n31062,
    n31063, n31064, n31065, n31066, n31067, n31068, n31069, n31070, n31071,
    n31072, n31073, n31074, n31075, n31076, n31077, n31078, n31079, n31080,
    n31081, n31082, n31083, n31084, n31085, n31086, n31087, n31088, n31089,
    n31090, n31091, n31092, n31093, n31094, n31095, n31096, n31097, n31098,
    n31099, n31100, n31101, n31102, n31103, n31104, n31105, n31106, n31107,
    n31108, n31109, n31110, n31111, n31112, n31113, n31114, n31115, n31116,
    n31117, n31119, n31120, n31121, n31122, n31123, n31124, n31125, n31126,
    n31127, n31128, n31129, n31130, n31131, n31132, n31133, n31134, n31135,
    n31136, n31137, n31138, n31139, n31140, n31141, n31142, n31143, n31144,
    n31145, n31146, n31147, n31148, n31149, n31150, n31151, n31152, n31153,
    n31154, n31155, n31156, n31157, n31158, n31159, n31160, n31161, n31162,
    n31163, n31164, n31166, n31167, n31168, n31169, n31170, n31171, n31172,
    n31173, n31174, n31175, n31176, n31177, n31178, n31179, n31180, n31181,
    n31182, n31183, n31184, n31185, n31186, n31187, n31188, n31189, n31190,
    n31191, n31192, n31193, n31194, n31195, n31196, n31197, n31199, n31200,
    n31201, n31202, n31203, n31204, n31205, n31206, n31207, n31208, n31209,
    n31210, n31211, n31212, n31213, n31214, n31215, n31216, n31217, n31218,
    n31219, n31220, n31221, n31222, n31223, n31224, n31225, n31226, n31227,
    n31228, n31229, n31230, n31231, n31232, n31233, n31234, n31235, n31236,
    n31237, n31238, n31239, n31240, n31241, n31242, n31243, n31244, n31246,
    n31247, n31248, n31249, n31250, n31251, n31252, n31253, n31254, n31255,
    n31256, n31257, n31258, n31259, n31260, n31261, n31262, n31263, n31264,
    n31265, n31266, n31267, n31268, n31269, n31270, n31271, n31272, n31273,
    n31274, n31275, n31276, n31277, n31278, n31279, n31280, n31281, n31283,
    n31284, n31285, n31286, n31287, n31288, n31289, n31290, n31291, n31292,
    n31293, n31294, n31295, n31296, n31297, n31298, n31299, n31300, n31301,
    n31302, n31303, n31304, n31305, n31306, n31307, n31308, n31309, n31310,
    n31311, n31312, n31313, n31314, n31315, n31316, n31317, n31318, n31319,
    n31320, n31322, n31323, n31324, n31325, n31326, n31327, n31328, n31329,
    n31330, n31331, n31332, n31333, n31334, n31335, n31336, n31337, n31338,
    n31339, n31340, n31341, n31342, n31343, n31344, n31345, n31346, n31347,
    n31348, n31349, n31350, n31351, n31352, n31353, n31354, n31355, n31356,
    n31357, n31358, n31359, n31360, n31361, n31362, n31364, n31365, n31366,
    n31367, n31368, n31369, n31370, n31371, n31372, n31373, n31374, n31375,
    n31376, n31377, n31378, n31379, n31380, n31381, n31382, n31383, n31384,
    n31385, n31386, n31387, n31388, n31389, n31390, n31391, n31392, n31393,
    n31394, n31395, n31396, n31397, n31398, n31399, n31401, n31402, n31403,
    n31404, n31405, n31406, n31407, n31408, n31409, n31410, n31411, n31412,
    n31413, n31414, n31415, n31416, n31417, n31418, n31419, n31420, n31421,
    n31422, n31423, n31424, n31425, n31426, n31427, n31428, n31429, n31431,
    n31432, n31433, n31434, n31435, n31436, n31437, n31438, n31439, n31440,
    n31441, n31442, n31443, n31444, n31445, n31446, n31447, n31448, n31449,
    n31450, n31451, n31452, n31453, n31454, n31455, n31456, n31457, n31459,
    n31460, n31461, n31462, n31463, n31464, n31465, n31466, n31467, n31468,
    n31469, n31470, n31471, n31472, n31473, n31474, n31475, n31476, n31477,
    n31478, n31479, n31480, n31481, n31482, n31483, n31484, n31485, n31486,
    n31487, n31488, n31489, n31490, n31492, n31493, n31494, n31495, n31496,
    n31497, n31498, n31499, n31500, n31501, n31502, n31503, n31504, n31505,
    n31506, n31507, n31508, n31509, n31510, n31511, n31512, n31513, n31514,
    n31515, n31516, n31517, n31518, n31519, n31520, n31521, n31522, n31523,
    n31524, n31525, n31526, n31527, n31529, n31530, n31531, n31532, n31533,
    n31534, n31535, n31536, n31537, n31538, n31539, n31540, n31541, n31542,
    n31543, n31544, n31545, n31546, n31547, n31548, n31549, n31550, n31551,
    n31552, n31553, n31554, n31555, n31556, n31557, n31558, n31559, n31560,
    n31561, n31562, n31564, n31565, n31566, n31567, n31568, n31569, n31570,
    n31571, n31572, n31573, n31574, n31575, n31576, n31577, n31578, n31579,
    n31580, n31581, n31582, n31583, n31584, n31585, n31586, n31587, n31588,
    n31589, n31590, n31591, n31592, n31593, n31594, n31595, n31596, n31597,
    n31598, n31599, n31600, n31601, n31602, n31603, n31605, n31606, n31607,
    n31608, n31609, n31610, n31611, n31612, n31613, n31614, n31615, n31616,
    n31617, n31618, n31619, n31620, n31621, n31622, n31623, n31624, n31625,
    n31626, n31627, n31628, n31629, n31630, n31631, n31632, n31633, n31634,
    n31635, n31636, n31637, n31638, n31639, n31640, n31641, n31642, n31643,
    n31644, n31645, n31646, n31648, n31649, n31650, n31651, n31652, n31653,
    n31654, n31655, n31656, n31657, n31658, n31659, n31660, n31661, n31662,
    n31663, n31664, n31665, n31666, n31667, n31668, n31669, n31670, n31671,
    n31672, n31673, n31674, n31675, n31676, n31677, n31678, n31679, n31680,
    n31681, n31682, n31684, n31685, n31686, n31687, n31688, n31689, n31690,
    n31691, n31692, n31693, n31694, n31695, n31696, n31697, n31698, n31699,
    n31700, n31701, n31702, n31703, n31704, n31705, n31706, n31707, n31708,
    n31709, n31710, n31711, n31712, n31713, n31714, n31715, n31716, n31717,
    n31718, n31719, n31720, n31721, n31722, n31724, n31725, n31726, n31727,
    n31728, n31729, n31730, n31731, n31732, n31733, n31734, n31735, n31736,
    n31737, n31738, n31739, n31740, n31741, n31742, n31743, n31744, n31745,
    n31746, n31747, n31748, n31749, n31750, n31751, n31752, n31753, n31754,
    n31755, n31756, n31757, n31758, n31760, n31761, n31762, n31763, n31764,
    n31765, n31766, n31767, n31768, n31769, n31770, n31771, n31772, n31773,
    n31774, n31775, n31776, n31777, n31778, n31779, n31780, n31781, n31782,
    n31783, n31784, n31785, n31786, n31787, n31788, n31789, n31790, n31791,
    n31792, n31793, n31794, n31795, n31796, n31797, n31798, n31799, n31800,
    n31801, n31802, n31803, n31804, n31805, n31806, n31807, n31808, n31809,
    n31810, n31811, n31812, n31813, n31814, n31815, n31816, n31817, n31818,
    n31819, n31820, n31821, n31822, n31823, n31824, n31825, n31826, n31827,
    n31828, n31829, n31830, n31831, n31832, n31833, n31834, n31835, n31836,
    n31837, n31838, n31839, n31840, n31841, n31842, n31843, n31844, n31845,
    n31846, n31847, n31848, n31849, n31850, n31851, n31852, n31853, n31854,
    n31855, n31856, n31857, n31858, n31859, n31860, n31861, n31863, n31864,
    n31865, n31866, n31867, n31868, n31869, n31870, n31871, n31872, n31873,
    n31874, n31875, n31876, n31877, n31878, n31879, n31880, n31881, n31882,
    n31883, n31884, n31885, n31886, n31887, n31888, n31889, n31890, n31891,
    n31892, n31893, n31894, n31895, n31896, n31897, n31898, n31899, n31900,
    n31901, n31902, n31903, n31904, n31905, n31906, n31907, n31908, n31909,
    n31910, n31911, n31912, n31913, n31914, n31915, n31916, n31917, n31918,
    n31919, n31920, n31921, n31922, n31923, n31924, n31925, n31926, n31927,
    n31928, n31929, n31930, n31931, n31932, n31933, n31934, n31935, n31936,
    n31937, n31938, n31939, n31940, n31941, n31942, n31943, n31944, n31945,
    n31946, n31947, n31948, n31949, n31950, n31951, n31952, n31953, n31954,
    n31955, n31956, n31957, n31958, n31959, n31960, n31961, n31962, n31963,
    n31964, n31965, n31966, n31967, n31968, n31969, n31971, n31972, n31973,
    n31974, n31975, n31976, n31977, n31978, n31979, n31980, n31981, n31982,
    n31983, n31984, n31985, n31986, n31987, n31988, n31989, n31990, n31991,
    n31992, n31993, n31994, n31995, n31996, n31997, n31998, n31999, n32000,
    n32001, n32002, n32003, n32004, n32005, n32006, n32007, n32008, n32009,
    n32010, n32011, n32012, n32013, n32014, n32015, n32016, n32017, n32018,
    n32019, n32020, n32021, n32022, n32023, n32024, n32025, n32026, n32027,
    n32028, n32029, n32030, n32031, n32032, n32033, n32034, n32035, n32036,
    n32037, n32038, n32039, n32040, n32041, n32042, n32043, n32044, n32045,
    n32046, n32047, n32048, n32049, n32050, n32051, n32052, n32053, n32054,
    n32055, n32056, n32057, n32058, n32059, n32060, n32061, n32062, n32063,
    n32064, n32065, n32066, n32067, n32068, n32069, n32070, n32071, n32072,
    n32073, n32074, n32076, n32077, n32078, n32079, n32080, n32081, n32082,
    n32083, n32084, n32085, n32086, n32087, n32088, n32089, n32090, n32091,
    n32092, n32093, n32094, n32095, n32096, n32097, n32098, n32099, n32100,
    n32101, n32102, n32103, n32104, n32105, n32106, n32107, n32108, n32109,
    n32110, n32111, n32112, n32113, n32114, n32115, n32117, n32118, n32119,
    n32120, n32121, n32122, n32123, n32124, n32125, n32126, n32127, n32128,
    n32129, n32130, n32131, n32132, n32133, n32134, n32135, n32136, n32137,
    n32138, n32139, n32140, n32141, n32142, n32143, n32144, n32145, n32146,
    n32147, n32148, n32149, n32150, n32151, n32152, n32153, n32154, n32156,
    n32157, n32158, n32159, n32160, n32161, n32162, n32163, n32164, n32165,
    n32166, n32167, n32168, n32169, n32170, n32171, n32172, n32173, n32174,
    n32175, n32176, n32177, n32178, n32179, n32180, n32181, n32182, n32183,
    n32184, n32185, n32186, n32187, n32188, n32189, n32190, n32191, n32192,
    n32193, n32194, n32195, n32196, n32197, n32198, n32199, n32200, n32201,
    n32202, n32203, n32204, n32205, n32206, n32207, n32208, n32209, n32210,
    n32211, n32212, n32213, n32214, n32215, n32216, n32217, n32218, n32219,
    n32220, n32221, n32222, n32223, n32224, n32225, n32226, n32227, n32228,
    n32229, n32230, n32231, n32232, n32233, n32234, n32235, n32236, n32237,
    n32238, n32239, n32240, n32241, n32242, n32243, n32244, n32245, n32246,
    n32247, n32248, n32249, n32250, n32251, n32252, n32253, n32254, n32255,
    n32256, n32258, n32259, n32260, n32261, n32262, n32263, n32264, n32265,
    n32266, n32267, n32268, n32269, n32270, n32271, n32272, n32273, n32274,
    n32275, n32276, n32277, n32278, n32279, n32280, n32281, n32282, n32283,
    n32284, n32285, n32286, n32287, n32288, n32289, n32290, n32291, n32292,
    n32293, n32294, n32295, n32296, n32297, n32298, n32299, n32300, n32301,
    n32302, n32303, n32304, n32305, n32306, n32307, n32308, n32309, n32310,
    n32311, n32312, n32313, n32314, n32315, n32316, n32317, n32318, n32319,
    n32320, n32321, n32322, n32323, n32324, n32325, n32326, n32327, n32328,
    n32329, n32330, n32331, n32332, n32333, n32334, n32335, n32336, n32337,
    n32338, n32339, n32340, n32341, n32342, n32343, n32344, n32345, n32346,
    n32347, n32348, n32350, n32351, n32352, n32353, n32354, n32355, n32356,
    n32357, n32358, n32359, n32360, n32361, n32362, n32363, n32364, n32365,
    n32366, n32367, n32368, n32369, n32370, n32371, n32372, n32373, n32374,
    n32375, n32376, n32377, n32378, n32379, n32380, n32381, n32382, n32383,
    n32384, n32385, n32386, n32387, n32388, n32389, n32390, n32391, n32392,
    n32393, n32394, n32395, n32396, n32397, n32398, n32400, n32401, n32402,
    n32403, n32404, n32405, n32406, n32407, n32408, n32409, n32410, n32411,
    n32412, n32413, n32414, n32415, n32416, n32417, n32418, n32419, n32420,
    n32421, n32422, n32423, n32424, n32425, n32426, n32427, n32428, n32429,
    n32430, n32431, n32432, n32433, n32434, n32435, n32436, n32437, n32438,
    n32439, n32440, n32441, n32442, n32443, n32444, n32445, n32446, n32447,
    n32448, n32449, n32450, n32451, n32452, n32453, n32454, n32455, n32456,
    n32457, n32458, n32459, n32460, n32461, n32462, n32463, n32464, n32465,
    n32466, n32467, n32468, n32469, n32470, n32471, n32472, n32473, n32474,
    n32475, n32476, n32477, n32478, n32479, n32480, n32481, n32482, n32483,
    n32484, n32485, n32486, n32487, n32488, n32489, n32490, n32491, n32492,
    n32493, n32494, n32495, n32496, n32497, n32498, n32499, n32500, n32502,
    n32503, n32504, n32505, n32506, n32507, n32508, n32509, n32510, n32511,
    n32512, n32513, n32514, n32515, n32516, n32517, n32518, n32519, n32520,
    n32521, n32522, n32523, n32524, n32525, n32526, n32527, n32528, n32529,
    n32530, n32531, n32532, n32533, n32534, n32535, n32536, n32537, n32538,
    n32539, n32540, n32541, n32542, n32543, n32544, n32545, n32546, n32547,
    n32548, n32549, n32550, n32551, n32552, n32554, n32555, n32556, n32557,
    n32558, n32559, n32560, n32561, n32562, n32563, n32564, n32565, n32566,
    n32567, n32568, n32569, n32570, n32571, n32572, n32573, n32574, n32575,
    n32576, n32577, n32578, n32579, n32580, n32581, n32582, n32583, n32584,
    n32585, n32587, n32588, n32589, n32590, n32591, n32592, n32593, n32594,
    n32595, n32596, n32597, n32598, n32599, n32600, n32601, n32602, n32603,
    n32604, n32605, n32606, n32607, n32608, n32609, n32610, n32611, n32612,
    n32613, n32614, n32615, n32616, n32617, n32618, n32619, n32620, n32621,
    n32622, n32623, n32624, n32625, n32626, n32627, n32628, n32629, n32630,
    n32631, n32633, n32634, n32635, n32636, n32637, n32638, n32639, n32640,
    n32641, n32642, n32643, n32644, n32645, n32646, n32647, n32648, n32649,
    n32650, n32651, n32652, n32653, n32654, n32655, n32656, n32657, n32658,
    n32659, n32660, n32661, n32663, n32664, n32665, n32666, n32667, n32668,
    n32669, n32670, n32671, n32672, n32673, n32674, n32675, n32676, n32677,
    n32678, n32679, n32680, n32681, n32682, n32683, n32684, n32685, n32686,
    n32687, n32688, n32689, n32690, n32691, n32692, n32693, n32694, n32695,
    n32696, n32697, n32698, n32699, n32700, n32701, n32702, n32703, n32704,
    n32705, n32706, n32707, n32709, n32710, n32711, n32712, n32713, n32714,
    n32715, n32716, n32717, n32718, n32719, n32720, n32721, n32722, n32723,
    n32724, n32725, n32726, n32727, n32728, n32729, n32730, n32731, n32732,
    n32733, n32734, n32735, n32736, n32737, n32738, n32739, n32740, n32741,
    n32742, n32743, n32744, n32746, n32747, n32748, n32749, n32750, n32751,
    n32752, n32753, n32754, n32755, n32756, n32757, n32758, n32759, n32760,
    n32761, n32762, n32763, n32764, n32765, n32766, n32767, n32768, n32769,
    n32770, n32771, n32772, n32773, n32774, n32775, n32776, n32777, n32778,
    n32779, n32780, n32781, n32782, n32783, n32784, n32785, n32786, n32787,
    n32788, n32789, n32790, n32791, n32792, n32793, n32794, n32795, n32796,
    n32797, n32798, n32799, n32800, n32801, n32802, n32803, n32804, n32805,
    n32806, n32807, n32808, n32809, n32810, n32811, n32812, n32813, n32814,
    n32815, n32816, n32817, n32818, n32819, n32820, n32821, n32822, n32823,
    n32824, n32825, n32826, n32827, n32828, n32829, n32830, n32831, n32832,
    n32833, n32834, n32835, n32836, n32837, n32838, n32839, n32840, n32841,
    n32842, n32843, n32845, n32846, n32847, n32848, n32849, n32850, n32851,
    n32852, n32853, n32854, n32855, n32856, n32857, n32858, n32859, n32860,
    n32861, n32862, n32863, n32864, n32865, n32866, n32867, n32868, n32869,
    n32870, n32871, n32872, n32873, n32874, n32875, n32876, n32877, n32878,
    n32879, n32880, n32881, n32882, n32883, n32884, n32885, n32886, n32888,
    n32889, n32890, n32891, n32892, n32893, n32894, n32895, n32896, n32897,
    n32898, n32899, n32900, n32901, n32902, n32903, n32904, n32905, n32906,
    n32907, n32908, n32909, n32910, n32911, n32912, n32913, n32914, n32915,
    n32916, n32917, n32918, n32919, n32920, n32921, n32922, n32924, n32925,
    n32926, n32927, n32928, n32929, n32930, n32931, n32932, n32933, n32934,
    n32935, n32936, n32937, n32938, n32939, n32940, n32941, n32942, n32943,
    n32944, n32945, n32946, n32947, n32948, n32949, n32950, n32951, n32952,
    n32953, n32954, n32955, n32956, n32957, n32958, n32959, n32960, n32961,
    n32962, n32963, n32964, n32965, n32966, n32967, n32968, n32969, n32970,
    n32971, n32972, n32973, n32974, n32975, n32976, n32977, n32978, n32979,
    n32980, n32981, n32982, n32983, n32984, n32985, n32986, n32987, n32988,
    n32989, n32990, n32991, n32992, n32993, n32994, n32995, n32996, n32997,
    n32998, n32999, n33000, n33001, n33002, n33003, n33004, n33005, n33006,
    n33007, n33008, n33009, n33010, n33011, n33012, n33013, n33014, n33015,
    n33016, n33017, n33018, n33019, n33020, n33021, n33023, n33024, n33025,
    n33026, n33027, n33028, n33029, n33030, n33031, n33032, n33033, n33034,
    n33035, n33036, n33037, n33038, n33039, n33040, n33041, n33042, n33043,
    n33044, n33045, n33046, n33047, n33048, n33049, n33050, n33051, n33052,
    n33053, n33054, n33055, n33056, n33057, n33058, n33059, n33060, n33061,
    n33062, n33063, n33064, n33065, n33066, n33068, n33069, n33070, n33071,
    n33072, n33073, n33074, n33075, n33076, n33077, n33078, n33079, n33080,
    n33081, n33082, n33083, n33084, n33085, n33086, n33087, n33088, n33089,
    n33090, n33091, n33092, n33093, n33094, n33095, n33096, n33097, n33098,
    n33099, n33100, n33101, n33102, n33103, n33104, n33105, n33106, n33108,
    n33109, n33110, n33111, n33112, n33113, n33114, n33115, n33116, n33117,
    n33118, n33119, n33120, n33121, n33122, n33123, n33124, n33125, n33126,
    n33127, n33128, n33129, n33130, n33131, n33132, n33133, n33134, n33135,
    n33136, n33137, n33138, n33139, n33141, n33142, n33143, n33144, n33145,
    n33146, n33147, n33148, n33149, n33150, n33151, n33152, n33153, n33154,
    n33155, n33156, n33157, n33158, n33159, n33160, n33161, n33162, n33163,
    n33164, n33165, n33166, n33167, n33168, n33169, n33170, n33171, n33172,
    n33174, n33175, n33176, n33177, n33178, n33179, n33180, n33181, n33182,
    n33183, n33184, n33185, n33186, n33187, n33188, n33189, n33190, n33191,
    n33192, n33193, n33194, n33195, n33196, n33197, n33198, n33199, n33200,
    n33201, n33202, n33203, n33204, n33205, n33206, n33207, n33208, n33210,
    n33211, n33212, n33213, n33214, n33215, n33216, n33217, n33218, n33219,
    n33220, n33221, n33222, n33223, n33224, n33225, n33226, n33227, n33228,
    n33229, n33230, n33231, n33232, n33233, n33234, n33235, n33236, n33237,
    n33238, n33239, n33240, n33241, n33242, n33243, n33244, n33245, n33246,
    n33247, n33248, n33250, n33251, n33252, n33253, n33254, n33255, n33256,
    n33257, n33258, n33259, n33260, n33261, n33262, n33263, n33264, n33265,
    n33266, n33267, n33268, n33269, n33270, n33271, n33272, n33273, n33274,
    n33275, n33276, n33277, n33278, n33279, n33280, n33281, n33282, n33283,
    n33285, n33286, n33287, n33288, n33289, n33290, n33291, n33292, n33293,
    n33294, n33295, n33296, n33297, n33298, n33299, n33300, n33301, n33302,
    n33303, n33304, n33305, n33306, n33307, n33308, n33309, n33310, n33311,
    n33313, n33314, n33315, n33316, n33317, n33318, n33319, n33320, n33321,
    n33322, n33323, n33324, n33325, n33326, n33327, n33328, n33329, n33330,
    n33331, n33332, n33333, n33334, n33335, n33336, n33337, n33338, n33339,
    n33340, n33341, n33342, n33343, n33344, n33345, n33346, n33347, n33349,
    n33350, n33351, n33352, n33353, n33354, n33355, n33356, n33357, n33358,
    n33359, n33360, n33361, n33362, n33363, n33364, n33365, n33366, n33367,
    n33368, n33369, n33370, n33371, n33372, n33373, n33374, n33375, n33376,
    n33377, n33378, n33379, n33380, n33381, n33382, n33383, n33385, n33386,
    n33387, n33388, n33389, n33390, n33391, n33392, n33393, n33394, n33395,
    n33396, n33397, n33398, n33399, n33400, n33401, n33402, n33403, n33404,
    n33405, n33406, n33407, n33408, n33409, n33410, n33411, n33412, n33413,
    n33414, n33415, n33416, n33417, n33418, n33419, n33420, n33421, n33422,
    n33423, n33424, n33425, n33426, n33427, n33428, n33429, n33431, n33432,
    n33433, n33434, n33435, n33436, n33437, n33438, n33439, n33440, n33441,
    n33442, n33443, n33444, n33445, n33446, n33447, n33448, n33449, n33450,
    n33451, n33452, n33453, n33454, n33455, n33456, n33457, n33458, n33459,
    n33460, n33461, n33462, n33463, n33464, n33465, n33467, n33468, n33469,
    n33470, n33471, n33472, n33473, n33474, n33475, n33476, n33477, n33478,
    n33479, n33480, n33481, n33482, n33483, n33484, n33485, n33486, n33487,
    n33488, n33489, n33490, n33491, n33492, n33493, n33494, n33495, n33497,
    n33498, n33499, n33500, n33501, n33502, n33503, n33504, n33505, n33506,
    n33507, n33508, n33509, n33510, n33511, n33512, n33513, n33514, n33515,
    n33516, n33517, n33518, n33519, n33520, n33521, n33522, n33523, n33524,
    n33525, n33526, n33527, n33528, n33529, n33530, n33531, n33532, n33533,
    n33534, n33535, n33536, n33537, n33538, n33539, n33540, n33541, n33542,
    n33543, n33544, n33545, n33546, n33547, n33548, n33549, n33550, n33551,
    n33552, n33553, n33554, n33555, n33556, n33557, n33558, n33559, n33560,
    n33561, n33562, n33563, n33564, n33565, n33566, n33567, n33568, n33569,
    n33570, n33571, n33572, n33573, n33574, n33575, n33576, n33577, n33578,
    n33579, n33580, n33581, n33582, n33583, n33584, n33585, n33586, n33587,
    n33588, n33589, n33590, n33591, n33592, n33593, n33594, n33595, n33596,
    n33597, n33599, n33600, n33601, n33602, n33603, n33604, n33605, n33606,
    n33607, n33608, n33609, n33610, n33611, n33612, n33613, n33614, n33615,
    n33616, n33617, n33618, n33619, n33620, n33621, n33622, n33623, n33624,
    n33625, n33626, n33627, n33628, n33629, n33630, n33631, n33632, n33633,
    n33634, n33635, n33636, n33637, n33638, n33639, n33640, n33641, n33642,
    n33643, n33644, n33645, n33646, n33647, n33648, n33649, n33650, n33651,
    n33652, n33653, n33654, n33655, n33656, n33657, n33658, n33659, n33660,
    n33661, n33662, n33663, n33664, n33665, n33666, n33667, n33668, n33669,
    n33670, n33671, n33672, n33673, n33674, n33675, n33676, n33677, n33678,
    n33679, n33680, n33681, n33682, n33683, n33684, n33685, n33686, n33687,
    n33688, n33689, n33690, n33691, n33692, n33693, n33694, n33695, n33696,
    n33697, n33698, n33700, n33701, n33702, n33703, n33704, n33705, n33706,
    n33707, n33708, n33709, n33710, n33711, n33712, n33713, n33714, n33715,
    n33716, n33717, n33718, n33719, n33720, n33721, n33722, n33723, n33724,
    n33725, n33726, n33727, n33728, n33729, n33730, n33731, n33732, n33733,
    n33734, n33735, n33736, n33737, n33738, n33739, n33740, n33741, n33742,
    n33743, n33744, n33745, n33746, n33747, n33748, n33749, n33750, n33751,
    n33752, n33753, n33754, n33755, n33756, n33757, n33758, n33759, n33760,
    n33761, n33762, n33763, n33764, n33765, n33766, n33767, n33768, n33769,
    n33770, n33771, n33772, n33773, n33774, n33775, n33776, n33777, n33778,
    n33779, n33780, n33781, n33782, n33783, n33784, n33785, n33786, n33787,
    n33788, n33789, n33790, n33791, n33792, n33793, n33794, n33795, n33796,
    n33797, n33799, n33800, n33801, n33802, n33803, n33804, n33805, n33806,
    n33807, n33808, n33809, n33810, n33811, n33812, n33813, n33814, n33815,
    n33816, n33817, n33818, n33819, n33820, n33821, n33822, n33823, n33824,
    n33825, n33826, n33827, n33828, n33829, n33830, n33831, n33832, n33833,
    n33834, n33835, n33836, n33837, n33838, n33839, n33840, n33841, n33842,
    n33843, n33844, n33845, n33846, n33847, n33848, n33849, n33850, n33851,
    n33852, n33853, n33854, n33855, n33856, n33857, n33858, n33859, n33860,
    n33861, n33862, n33863, n33864, n33865, n33866, n33867, n33868, n33869,
    n33870, n33871, n33872, n33873, n33874, n33875, n33876, n33877, n33878,
    n33879, n33880, n33881, n33882, n33883, n33884, n33885, n33886, n33887,
    n33888, n33889, n33890, n33891, n33892, n33893, n33894, n33895, n33896,
    n33897, n33898, n33899, n33900, n33901, n33903, n33904, n33905, n33906,
    n33907, n33908, n33909, n33910, n33911, n33912, n33913, n33914, n33915,
    n33916, n33917, n33918, n33919, n33920, n33921, n33922, n33923, n33924,
    n33925, n33926, n33927, n33928, n33929, n33930, n33931, n33932, n33933,
    n33934, n33935, n33936, n33937, n33938, n33939, n33940, n33941, n33942,
    n33943, n33944, n33945, n33946, n33947, n33949, n33950, n33951, n33952,
    n33953, n33954, n33955, n33956, n33957, n33958, n33959, n33960, n33961,
    n33962, n33963, n33964, n33965, n33966, n33967, n33968, n33969, n33970,
    n33971, n33972, n33973, n33974, n33975, n33976, n33977, n33978, n33979,
    n33980, n33981, n33982, n33983, n33984, n33985, n33986, n33987, n33988,
    n33989, n33990, n33991, n33992, n33993, n33995, n33996, n33997, n33998,
    n33999, n34000, n34001, n34002, n34003, n34004, n34005, n34006, n34007,
    n34008, n34009, n34010, n34011, n34012, n34013, n34014, n34015, n34016,
    n34017, n34018, n34019, n34020, n34021, n34022, n34023, n34024, n34025,
    n34026, n34027, n34028, n34029, n34030, n34031, n34032, n34033, n34034,
    n34035, n34036, n34037, n34038, n34039, n34040, n34041, n34042, n34043,
    n34044, n34045, n34046, n34047, n34048, n34049, n34050, n34051, n34052,
    n34053, n34054, n34055, n34056, n34057, n34058, n34059, n34060, n34061,
    n34062, n34063, n34064, n34065, n34066, n34067, n34068, n34069, n34070,
    n34071, n34072, n34073, n34074, n34075, n34076, n34077, n34078, n34079,
    n34080, n34081, n34082, n34083, n34084, n34085, n34086, n34087, n34088,
    n34089, n34090, n34091, n34092, n34093, n34094, n34095, n34096, n34097,
    n34098, n34100, n34101, n34102, n34103, n34104, n34105, n34106, n34107,
    n34108, n34109, n34110, n34111, n34112, n34113, n34114, n34115, n34116,
    n34117, n34118, n34119, n34120, n34121, n34122, n34123, n34124, n34125,
    n34126, n34127, n34128, n34129, n34130, n34131, n34133, n34134, n34135,
    n34136, n34137, n34138, n34139, n34140, n34141, n34142, n34143, n34144,
    n34145, n34146, n34147, n34148, n34149, n34150, n34151, n34152, n34153,
    n34154, n34155, n34156, n34157, n34158, n34159, n34160, n34161, n34162,
    n34163, n34164, n34165, n34166, n34167, n34168, n34169, n34170, n34171,
    n34172, n34174, n34175, n34176, n34177, n34178, n34179, n34180, n34181,
    n34182, n34183, n34184, n34185, n34186, n34187, n34188, n34189, n34190,
    n34191, n34192, n34193, n34194, n34195, n34196, n34197, n34198, n34199,
    n34200, n34201, n34202, n34203, n34204, n34205, n34206, n34207, n34208,
    n34209, n34210, n34211, n34212, n34213, n34214, n34215, n34216, n34217,
    n34218, n34219, n34220, n34221, n34222, n34223, n34224, n34225, n34226,
    n34227, n34228, n34229, n34230, n34231, n34232, n34233, n34234, n34235,
    n34236, n34237, n34238, n34239, n34240, n34241, n34242, n34243, n34244,
    n34245, n34246, n34247, n34248, n34249, n34250, n34251, n34252, n34253,
    n34254, n34255, n34256, n34257, n34258, n34259, n34260, n34261, n34262,
    n34263, n34264, n34265, n34267, n34268, n34269, n34270, n34271, n34272,
    n34273, n34274, n34275, n34276, n34277, n34278, n34279, n34280, n34281,
    n34282, n34283, n34284, n34285, n34286, n34287, n34288, n34289, n34290,
    n34291, n34292, n34293, n34294, n34295, n34296, n34297, n34298, n34299,
    n34300, n34301, n34302, n34303, n34304, n34305, n34306, n34307, n34308,
    n34309, n34311, n34312, n34313, n34314, n34315, n34316, n34317, n34318,
    n34319, n34320, n34321, n34322, n34323, n34324, n34325, n34326, n34327,
    n34328, n34329, n34330, n34331, n34332, n34333, n34334, n34335, n34336,
    n34337, n34338, n34339, n34340, n34341, n34342, n34343, n34344, n34345,
    n34346, n34347, n34348, n34349, n34350, n34351, n34352, n34353, n34354,
    n34355, n34356, n34357, n34358, n34359, n34360, n34361, n34362, n34363,
    n34364, n34365, n34366, n34367, n34368, n34369, n34370, n34371, n34372,
    n34373, n34374, n34375, n34376, n34377, n34378, n34379, n34380, n34381,
    n34382, n34383, n34384, n34385, n34386, n34387, n34388, n34389, n34390,
    n34391, n34392, n34393, n34394, n34395, n34396, n34397, n34398, n34399,
    n34400, n34401, n34402, n34403, n34404, n34405, n34406, n34407, n34408,
    n34409, n34410, n34411, n34413, n34414, n34415, n34416, n34417, n34418,
    n34419, n34420, n34421, n34422, n34423, n34424, n34425, n34426, n34427,
    n34428, n34429, n34430, n34431, n34432, n34433, n34434, n34435, n34436,
    n34437, n34438, n34439, n34440, n34441, n34442, n34443, n34444, n34446,
    n34447, n34448, n34449, n34450, n34451, n34452, n34453, n34454, n34455,
    n34456, n34457, n34458, n34459, n34460, n34461, n34462, n34463, n34464,
    n34465, n34466, n34467, n34468, n34469, n34470, n34471, n34472, n34473,
    n34474, n34475, n34476, n34477, n34478, n34479, n34480, n34481, n34482,
    n34483, n34484, n34485, n34487, n34488, n34489, n34490, n34491, n34492,
    n34493, n34494, n34495, n34496, n34497, n34498, n34499, n34500, n34501,
    n34502, n34503, n34504, n34505, n34506, n34507, n34508, n34509, n34510,
    n34511, n34512, n34513, n34514, n34515, n34516, n34517, n34518, n34519,
    n34520, n34521, n34522, n34523, n34524, n34525, n34526, n34527, n34528,
    n34529, n34530, n34531, n34532, n34533, n34534, n34536, n34537, n34538,
    n34539, n34540, n34541, n34542, n34543, n34544, n34545, n34546, n34547,
    n34548, n34549, n34550, n34551, n34552, n34553, n34554, n34555, n34556,
    n34557, n34558, n34559, n34560, n34561, n34562, n34563, n34564, n34565,
    n34566, n34567, n34568, n34569, n34570, n34571, n34572, n34573, n34574,
    n34575, n34576, n34577, n34578, n34579, n34580, n34581, n34582, n34583,
    n34584, n34585, n34586, n34588, n34589, n34590, n34591, n34592, n34593,
    n34594, n34595, n34596, n34597, n34598, n34599, n34600, n34601, n34602,
    n34603, n34604, n34605, n34606, n34607, n34608, n34609, n34610, n34611,
    n34612, n34613, n34614, n34615, n34616, n34617, n34618, n34619, n34620,
    n34621, n34622, n34624, n34625, n34626, n34627, n34628, n34629, n34630,
    n34631, n34632, n34633, n34634, n34635, n34636, n34637, n34638, n34639,
    n34640, n34641, n34642, n34643, n34644, n34645, n34646, n34647, n34648,
    n34649, n34650, n34651, n34652, n34653, n34654, n34655, n34656, n34657,
    n34658, n34659, n34660, n34661, n34662, n34664, n34665, n34666, n34667,
    n34668, n34669, n34670, n34671, n34672, n34673, n34674, n34675, n34676,
    n34677, n34678, n34679, n34680, n34681, n34682, n34683, n34684, n34685,
    n34686, n34687, n34688, n34689, n34690, n34691, n34692, n34693, n34694,
    n34695, n34696, n34697, n34698, n34699, n34701, n34702, n34703, n34704,
    n34705, n34706, n34707, n34708, n34709, n34710, n34711, n34712, n34713,
    n34714, n34715, n34716, n34717, n34718, n34719, n34720, n34721, n34722,
    n34723, n34724, n34725, n34726, n34727, n34728, n34729, n34731, n34732,
    n34733, n34734, n34735, n34736, n34737, n34738, n34739, n34740, n34741,
    n34742, n34743, n34744, n34745, n34746, n34747, n34748, n34749, n34750,
    n34751, n34752, n34753, n34754, n34755, n34756, n34757, n34758, n34759,
    n34760, n34761, n34762, n34763, n34764, n34765, n34766, n34767, n34768,
    n34769, n34770, n34771, n34772, n34773, n34774, n34775, n34776, n34778,
    n34779, n34780, n34781, n34782, n34783, n34784, n34785, n34786, n34787,
    n34788, n34789, n34790, n34791, n34792, n34793, n34794, n34795, n34796,
    n34797, n34798, n34799, n34800, n34801, n34802, n34803, n34804, n34805,
    n34806, n34807, n34808, n34809, n34810, n34812, n34813, n34814, n34815,
    n34816, n34817, n34818, n34819, n34820, n34821, n34822, n34823, n34824,
    n34825, n34826, n34827, n34828, n34829, n34830, n34831, n34832, n34833,
    n34834, n34835, n34836, n34837, n34838, n34839, n34840, n34841, n34842,
    n34843, n34844, n34845, n34846, n34848, n34849, n34850, n34851, n34852,
    n34853, n34854, n34855, n34856, n34857, n34858, n34859, n34860, n34861,
    n34862, n34863, n34864, n34865, n34866, n34867, n34868, n34869, n34870,
    n34871, n34872, n34873, n34874, n34875, n34876, n34877, n34878, n34879,
    n34880, n34881, n34882, n34883, n34885, n34886, n34887, n34888, n34889,
    n34890, n34891, n34892, n34893, n34894, n34895, n34896, n34897, n34898,
    n34899, n34900, n34901, n34902, n34903, n34904, n34905, n34906, n34907,
    n34908, n34909, n34910, n34911, n34912, n34913, n34914, n34915, n34916,
    n34917, n34918, n34919, n34920, n34921, n34922, n34923, n34924, n34925,
    n34926, n34927, n34928, n34929, n34930, n34931, n34932, n34933, n34934,
    n34935, n34936, n34937, n34938, n34939, n34940, n34941, n34942, n34943,
    n34944, n34945, n34946, n34947, n34948, n34949, n34950, n34951, n34952,
    n34953, n34954, n34955, n34956, n34957, n34958, n34959, n34960, n34961,
    n34962, n34963, n34964, n34965, n34966, n34967, n34968, n34969, n34970,
    n34971, n34972, n34973, n34974, n34975, n34976, n34977, n34978, n34979,
    n34981, n34982, n34983, n34984, n34985, n34986, n34987, n34988, n34989,
    n34990, n34991, n34992, n34993, n34994, n34995, n34996, n34997, n34998,
    n34999, n35000, n35001, n35002, n35003, n35004, n35005, n35006, n35007,
    n35008, n35009, n35010, n35011, n35012, n35013, n35014, n35015, n35016,
    n35017, n35018, n35019, n35020, n35021, n35022, n35023, n35024, n35026,
    n35027, n35028, n35029, n35030, n35031, n35032, n35033, n35034, n35035,
    n35036, n35037, n35038, n35039, n35040, n35041, n35042, n35043, n35044,
    n35045, n35046, n35047, n35048, n35049, n35050, n35051, n35052, n35053,
    n35054, n35055, n35057, n35058, n35059, n35060, n35061, n35062, n35063,
    n35064, n35065, n35066, n35067, n35068, n35069, n35070, n35071, n35072,
    n35073, n35074, n35075, n35076, n35077, n35078, n35079, n35080, n35081,
    n35082, n35083, n35084, n35085, n35087, n35088, n35089, n35090, n35091,
    n35092, n35093, n35094, n35095, n35096, n35097, n35098, n35099, n35100,
    n35101, n35102, n35103, n35104, n35105, n35106, n35107, n35108, n35109,
    n35110, n35111, n35112, n35113, n35114, n35115, n35116, n35117, n35118,
    n35119, n35120, n35121, n35123, n35124, n35125, n35126, n35127, n35128,
    n35129, n35130, n35131, n35132, n35133, n35134, n35135, n35136, n35137,
    n35138, n35139, n35140, n35141, n35142, n35143, n35144, n35145, n35146,
    n35147, n35148, n35149, n35150, n35151, n35152, n35153, n35154, n35155,
    n35156, n35157, n35158, n35160, n35161, n35162, n35163, n35164, n35165,
    n35166, n35167, n35168, n35169, n35170, n35171, n35172, n35173, n35174,
    n35175, n35176, n35177, n35178, n35179, n35180, n35181, n35182, n35183,
    n35184, n35185, n35186, n35187, n35188, n35189, n35190, n35191, n35192,
    n35193, n35194, n35195, n35197, n35198, n35199, n35200, n35201, n35202,
    n35203, n35204, n35205, n35206, n35207, n35208, n35209, n35210, n35211,
    n35212, n35213, n35214, n35215, n35216, n35217, n35218, n35219, n35220,
    n35221, n35222, n35223, n35224, n35225, n35226, n35227, n35228, n35229,
    n35230, n35231, n35233, n35234, n35235, n35236, n35237, n35238, n35239,
    n35240, n35241, n35242, n35243, n35244, n35245, n35246, n35247, n35248,
    n35249, n35250, n35251, n35252, n35253, n35254, n35255, n35256, n35257,
    n35258, n35259, n35260, n35261, n35262, n35263, n35264, n35265, n35266,
    n35267, n35268, n35269, n35270, n35271, n35272, n35273, n35274, n35275,
    n35276, n35277, n35278, n35279, n35280, n35281, n35282, n35283, n35284,
    n35285, n35286, n35287, n35288, n35289, n35290, n35291, n35292, n35293,
    n35294, n35295, n35296, n35297, n35298, n35299, n35300, n35301, n35302,
    n35303, n35304, n35305, n35306, n35307, n35308, n35309, n35310, n35311,
    n35312, n35313, n35314, n35315, n35316, n35317, n35318, n35319, n35320,
    n35321, n35322, n35323, n35324, n35325, n35326, n35327, n35328, n35329,
    n35330, n35331, n35332, n35333, n35334, n35336, n35337, n35338, n35339,
    n35340, n35341, n35342, n35343, n35344, n35345, n35346, n35347, n35348,
    n35349, n35350, n35351, n35352, n35353, n35354, n35355, n35356, n35357,
    n35358, n35359, n35360, n35361, n35362, n35363, n35364, n35365, n35366,
    n35367, n35368, n35369, n35370, n35371, n35372, n35373, n35374, n35375,
    n35376, n35377, n35378, n35379, n35380, n35381, n35382, n35383, n35384,
    n35385, n35386, n35387, n35388, n35389, n35390, n35391, n35392, n35393,
    n35394, n35395, n35396, n35397, n35398, n35399, n35400, n35401, n35402,
    n35403, n35404, n35405, n35406, n35407, n35408, n35409, n35410, n35411,
    n35412, n35413, n35414, n35415, n35416, n35417, n35418, n35419, n35420,
    n35421, n35422, n35423, n35424, n35425, n35426, n35427, n35428, n35429,
    n35430, n35431, n35432, n35433, n35434, n35435, n35436, n35437, n35438,
    n35439, n35440, n35441, n35442, n35444, n35445, n35446, n35447, n35448,
    n35449, n35450, n35451, n35452, n35453, n35454, n35455, n35456, n35457,
    n35458, n35459, n35460, n35461, n35462, n35463, n35464, n35465, n35466,
    n35467, n35468, n35469, n35470, n35471, n35472, n35473, n35474, n35475,
    n35476, n35477, n35478, n35479, n35480, n35481, n35482, n35483, n35485,
    n35486, n35487, n35488, n35489, n35490, n35491, n35492, n35493, n35494,
    n35495, n35496, n35497, n35498, n35499, n35500, n35501, n35502, n35503,
    n35504, n35505, n35506, n35507, n35508, n35509, n35510, n35511, n35512,
    n35513, n35514, n35515, n35516, n35517, n35518, n35519, n35520, n35521,
    n35522, n35523, n35524, n35525, n35526, n35527, n35528, n35529, n35530,
    n35531, n35532, n35533, n35534, n35535, n35536, n35537, n35538, n35539,
    n35540, n35541, n35542, n35543, n35544, n35545, n35546, n35547, n35548,
    n35549, n35550, n35551, n35552, n35553, n35554, n35555, n35556, n35557,
    n35558, n35559, n35560, n35561, n35562, n35563, n35564, n35565, n35566,
    n35567, n35568, n35569, n35570, n35571, n35572, n35573, n35574, n35575,
    n35576, n35578, n35579, n35580, n35581, n35582, n35583, n35584, n35585,
    n35586, n35587, n35588, n35589, n35590, n35591, n35592, n35593, n35594,
    n35595, n35596, n35597, n35598, n35599, n35600, n35601, n35602, n35603,
    n35604, n35605, n35606, n35607, n35608, n35609, n35610, n35611, n35612,
    n35613, n35614, n35615, n35616, n35617, n35618, n35619, n35620, n35621,
    n35622, n35623, n35624, n35625, n35626, n35627, n35628, n35629, n35630,
    n35631, n35632, n35633, n35634, n35635, n35636, n35637, n35638, n35639,
    n35640, n35641, n35642, n35643, n35644, n35645, n35646, n35647, n35648,
    n35649, n35650, n35651, n35652, n35653, n35654, n35655, n35656, n35657,
    n35658, n35659, n35660, n35661, n35662, n35663, n35664, n35665, n35666,
    n35667, n35668, n35669, n35670, n35671, n35672, n35673, n35674, n35675,
    n35676, n35677, n35678, n35679, n35680, n35681, n35682, n35683, n35685,
    n35686, n35687, n35688, n35689, n35690, n35691, n35692, n35693, n35694,
    n35695, n35696, n35697, n35698, n35699, n35700, n35701, n35702, n35703,
    n35704, n35705, n35706, n35707, n35708, n35709, n35710, n35711, n35712,
    n35713, n35714, n35715, n35716, n35717, n35718, n35719, n35720, n35721,
    n35722, n35723, n35725, n35726, n35727, n35728, n35729, n35730, n35731,
    n35732, n35733, n35734, n35735, n35736, n35737, n35738, n35739, n35740,
    n35741, n35742, n35743, n35744, n35745, n35746, n35747, n35748, n35749,
    n35750, n35751, n35752, n35753, n35754, n35755, n35756, n35757, n35758,
    n35759, n35760, n35761, n35762, n35763, n35764, n35765, n35766, n35767,
    n35768, n35769, n35770, n35771, n35772, n35773, n35774, n35775, n35777,
    n35778, n35779, n35780, n35781, n35782, n35783, n35784, n35785, n35786,
    n35787, n35788, n35789, n35790, n35791, n35792, n35793, n35794, n35795,
    n35796, n35797, n35798, n35799, n35800, n35801, n35802, n35803, n35804,
    n35805, n35806, n35807, n35808, n35810, n35811, n35812, n35813, n35814,
    n35815, n35816, n35817, n35818, n35819, n35820, n35821, n35822, n35823,
    n35824, n35825, n35826, n35827, n35828, n35829, n35830, n35831, n35832,
    n35833, n35834, n35835, n35836, n35837, n35838, n35839, n35840, n35841,
    n35842, n35843, n35844, n35845, n35846, n35847, n35848, n35849, n35850,
    n35851, n35852, n35853, n35854, n35855, n35856, n35857, n35858, n35859,
    n35860, n35861, n35862, n35863, n35864, n35865, n35866, n35867, n35868,
    n35869, n35870, n35871, n35872, n35873, n35874, n35875, n35876, n35877,
    n35878, n35879, n35880, n35881, n35882, n35883, n35884, n35885, n35886,
    n35887, n35888, n35889, n35890, n35891, n35892, n35893, n35894, n35895,
    n35896, n35897, n35898, n35899, n35900, n35901, n35902, n35903, n35904,
    n35905, n35906, n35907, n35909, n35910, n35911, n35912, n35913, n35914,
    n35915, n35916, n35917, n35918, n35919, n35920, n35921, n35922, n35923,
    n35924, n35925, n35926, n35927, n35928, n35929, n35930, n35931, n35932,
    n35933, n35934, n35935, n35936, n35937, n35938, n35939, n35940, n35941,
    n35942, n35943, n35944, n35945, n35946, n35947, n35948, n35949, n35950,
    n35951, n35952, n35953, n35954, n35955, n35956, n35957, n35958, n35959,
    n35960, n35961, n35962, n35963, n35964, n35965, n35966, n35967, n35968,
    n35969, n35970, n35971, n35972, n35973, n35974, n35975, n35976, n35977,
    n35978, n35979, n35980, n35981, n35982, n35983, n35984, n35985, n35986,
    n35987, n35988, n35989, n35990, n35991, n35992, n35993, n35994, n35995,
    n35996, n35997, n35998, n35999, n36000, n36001, n36002, n36003, n36004,
    n36005, n36006, n36007, n36008, n36009, n36010, n36012, n36013, n36014,
    n36015, n36016, n36017, n36018, n36019, n36020, n36021, n36022, n36023,
    n36024, n36025, n36026, n36027, n36028, n36029, n36030, n36031, n36032,
    n36033, n36034, n36035, n36036, n36037, n36038, n36039, n36040, n36041,
    n36042, n36043, n36044, n36045, n36046, n36047, n36048, n36049, n36050,
    n36051, n36052, n36053, n36055, n36056, n36057, n36058, n36059, n36060,
    n36061, n36062, n36063, n36064, n36065, n36066, n36067, n36068, n36069,
    n36070, n36071, n36072, n36073, n36074, n36075, n36076, n36077, n36078,
    n36079, n36080, n36081, n36082, n36083, n36084, n36085, n36086, n36087,
    n36088, n36089, n36090, n36091, n36092, n36093, n36094, n36095, n36096,
    n36097, n36098, n36099, n36100, n36101, n36102, n36103, n36104, n36105,
    n36106, n36107, n36108, n36109, n36110, n36111, n36112, n36113, n36114,
    n36115, n36116, n36117, n36118, n36119, n36120, n36121, n36122, n36123,
    n36124, n36125, n36126, n36127, n36128, n36129, n36130, n36131, n36132,
    n36133, n36134, n36135, n36136, n36137, n36138, n36139, n36140, n36141,
    n36142, n36143, n36144, n36145, n36146, n36147, n36148, n36149, n36150,
    n36151, n36152, n36153, n36155, n36156, n36157, n36158, n36159, n36160,
    n36161, n36162, n36163, n36164, n36165, n36166, n36167, n36168, n36169,
    n36170, n36171, n36172, n36173, n36174, n36175, n36176, n36177, n36178,
    n36179, n36180, n36181, n36182, n36183, n36184, n36185, n36186, n36187,
    n36188, n36189, n36190, n36191, n36193, n36194, n36195, n36196, n36197,
    n36198, n36199, n36200, n36201, n36202, n36203, n36204, n36205, n36206,
    n36207, n36208, n36209, n36210, n36211, n36212, n36213, n36214, n36215,
    n36216, n36217, n36218, n36219, n36220, n36221, n36222, n36223, n36224,
    n36225, n36226, n36227, n36228, n36229, n36230, n36231, n36232, n36233,
    n36234, n36235, n36236, n36237, n36238, n36239, n36240, n36241, n36242,
    n36243, n36244, n36245, n36246, n36247, n36248, n36249, n36250, n36251,
    n36252, n36253, n36254, n36255, n36256, n36257, n36258, n36259, n36260,
    n36261, n36262, n36263, n36264, n36265, n36266, n36267, n36268, n36269,
    n36270, n36271, n36272, n36273, n36274, n36275, n36276, n36277, n36278,
    n36279, n36280, n36281, n36282, n36283, n36284, n36285, n36286, n36287,
    n36288, n36289, n36290, n36291, n36292, n36293, n36294, n36296, n36297,
    n36298, n36299, n36300, n36301, n36302, n36303, n36304, n36305, n36306,
    n36307, n36308, n36309, n36310, n36311, n36312, n36313, n36314, n36315,
    n36316, n36317, n36318, n36319, n36320, n36321, n36322, n36323, n36324,
    n36325, n36326, n36327, n36328, n36329, n36330, n36331, n36332, n36333,
    n36334, n36335, n36336, n36337, n36338, n36339, n36340, n36342, n36343,
    n36344, n36345, n36346, n36347, n36348, n36349, n36350, n36351, n36352,
    n36353, n36354, n36355, n36356, n36357, n36358, n36359, n36360, n36361,
    n36362, n36363, n36364, n36365, n36366, n36367, n36368, n36369, n36370,
    n36371, n36372, n36373, n36374, n36375, n36376, n36378, n36379, n36380,
    n36381, n36382, n36383, n36384, n36385, n36386, n36387, n36388, n36389,
    n36390, n36391, n36392, n36393, n36394, n36395, n36396, n36397, n36398,
    n36399, n36400, n36401, n36402, n36403, n36404, n36405, n36406, n36407,
    n36408, n36409, n36410, n36411, n36412, n36413, n36414, n36415, n36417,
    n36418, n36419, n36420, n36421, n36422, n36423, n36424, n36425, n36426,
    n36427, n36428, n36429, n36430, n36431, n36432, n36433, n36434, n36435,
    n36436, n36437, n36438, n36439, n36440, n36441, n36442, n36443, n36444,
    n36445, n36446, n36447, n36448, n36449, n36451, n36452, n36453, n36454,
    n36455, n36456, n36457, n36458, n36459, n36460, n36461, n36462, n36463,
    n36464, n36465, n36466, n36467, n36468, n36469, n36470, n36471, n36472,
    n36473, n36474, n36475, n36476, n36477, n36478, n36479, n36480, n36481,
    n36482, n36483, n36484, n36485, n36486, n36487, n36488, n36489, n36490,
    n36491, n36492, n36493, n36494, n36495, n36496, n36498, n36499, n36500,
    n36501, n36502, n36503, n36504, n36505, n36506, n36507, n36508, n36509,
    n36510, n36511, n36512, n36513, n36514, n36515, n36516, n36517, n36518,
    n36519, n36520, n36521, n36522, n36523, n36524, n36525, n36526, n36527,
    n36528, n36529, n36530, n36531, n36532, n36533, n36534, n36535, n36536,
    n36538, n36539, n36540, n36541, n36542, n36543, n36544, n36545, n36546,
    n36547, n36548, n36549, n36550, n36551, n36552, n36553, n36554, n36555,
    n36556, n36557, n36558, n36559, n36560, n36561, n36562, n36563, n36564,
    n36565, n36566, n36567, n36568, n36569, n36570, n36571, n36572, n36573,
    n36574, n36575, n36576, n36577, n36578, n36579, n36581, n36582, n36583,
    n36584, n36585, n36586, n36587, n36588, n36589, n36590, n36591, n36592,
    n36593, n36594, n36595, n36596, n36597, n36598, n36599, n36600, n36601,
    n36602, n36603, n36604, n36605, n36606, n36607, n36608, n36609, n36610,
    n36611, n36612, n36614, n36615, n36616, n36617, n36618, n36619, n36620,
    n36621, n36622, n36623, n36624, n36625, n36626, n36627, n36628, n36629,
    n36630, n36631, n36632, n36633, n36634, n36635, n36636, n36637, n36638,
    n36639, n36640, n36641, n36642, n36643, n36644, n36645, n36646, n36647,
    n36648, n36649, n36650, n36651, n36652, n36653, n36654, n36655, n36656,
    n36657, n36658, n36660, n36661, n36662, n36663, n36664, n36665, n36666,
    n36667, n36668, n36669, n36670, n36671, n36672, n36673, n36674, n36675,
    n36676, n36677, n36678, n36679, n36680, n36681, n36682, n36683, n36684,
    n36685, n36686, n36687, n36688, n36689, n36690, n36691, n36692, n36693,
    n36694, n36695, n36697, n36698, n36699, n36700, n36701, n36702, n36703,
    n36704, n36705, n36706, n36707, n36708, n36709, n36710, n36711, n36712,
    n36713, n36714, n36715, n36716, n36717, n36718, n36719, n36720, n36721,
    n36722, n36723, n36724, n36725, n36726, n36728, n36729, n36730, n36731,
    n36732, n36733, n36734, n36735, n36736, n36737, n36738, n36739, n36740,
    n36741, n36742, n36743, n36744, n36745, n36746, n36747, n36748, n36749,
    n36750, n36751, n36752, n36753, n36754, n36756, n36757, n36758, n36759,
    n36760, n36761, n36762, n36763, n36764, n36765, n36766, n36767, n36768,
    n36769, n36770, n36771, n36772, n36773, n36774, n36775, n36776, n36777,
    n36778, n36779, n36780, n36781, n36782, n36783, n36784, n36785, n36786,
    n36787, n36789, n36790, n36791, n36792, n36793, n36794, n36795, n36796,
    n36797, n36798, n36799, n36800, n36801, n36802, n36803, n36804, n36805,
    n36806, n36807, n36808, n36809, n36810, n36811, n36812, n36813, n36814,
    n36815, n36816, n36817, n36818, n36819, n36820, n36821, n36822, n36823,
    n36825, n36826, n36827, n36828, n36829, n36830, n36831, n36832, n36833,
    n36834, n36835, n36836, n36837, n36838, n36839, n36840, n36841, n36842,
    n36843, n36844, n36845, n36846, n36847, n36848, n36849, n36850, n36851,
    n36852, n36853, n36854, n36855, n36856, n36857, n36858, n36859, n36860,
    n36862, n36863, n36864, n36865, n36866, n36867, n36868, n36869, n36870,
    n36871, n36872, n36873, n36874, n36875, n36876, n36877, n36878, n36879,
    n36880, n36881, n36882, n36883, n36884, n36885, n36886, n36887, n36888,
    n36889, n36890, n36892, n36893, n36894, n36895, n36896, n36897, n36898,
    n36899, n36900, n36901, n36902, n36903, n36904, n36905, n36906, n36907,
    n36908, n36909, n36910, n36911, n36912, n36913, n36914, n36915, n36916,
    n36917, n36918, n36919, n36920, n36921, n36922, n36923, n36924, n36925,
    n36926, n36927, n36928, n36929, n36930, n36932, n36933, n36934, n36935,
    n36936, n36937, n36938, n36939, n36940, n36941, n36942, n36943, n36944,
    n36945, n36946, n36947, n36948, n36949, n36950, n36951, n36952, n36953,
    n36954, n36955, n36956, n36957, n36958, n36959, n36960, n36961, n36962,
    n36963, n36964, n36965, n36966, n36968, n36969, n36970, n36971, n36972,
    n36973, n36974, n36975, n36976, n36977, n36978, n36979, n36980, n36981,
    n36982, n36983, n36984, n36985, n36986, n36987, n36988, n36989, n36990,
    n36991, n36992, n36993, n36994, n36995, n36996, n36997, n36998, n36999,
    n37000, n37001, n37002, n37003, n37004, n37005, n37006, n37007, n37008,
    n37009, n37010, n37011, n37012, n37013, n37014, n37015, n37016, n37017,
    n37018, n37019, n37020, n37021, n37022, n37023, n37024, n37025, n37026,
    n37027, n37028, n37029, n37030, n37031, n37032, n37033, n37034, n37035,
    n37036, n37037, n37038, n37039, n37040, n37041, n37042, n37043, n37044,
    n37045, n37046, n37047, n37048, n37049, n37050, n37051, n37052, n37053,
    n37054, n37055, n37056, n37057, n37058, n37059, n37060, n37061, n37062,
    n37063, n37064, n37065, n37066, n37067, n37068, n37070, n37071, n37072,
    n37073, n37074, n37075, n37076, n37077, n37078, n37079, n37080, n37081,
    n37082, n37083, n37084, n37085, n37086, n37087, n37088, n37089, n37090,
    n37091, n37092, n37093, n37094, n37095, n37096, n37097, n37098, n37099,
    n37100, n37101, n37102, n37103, n37104, n37105, n37106, n37107, n37108,
    n37109, n37110, n37111, n37112, n37113, n37114, n37115, n37116, n37117,
    n37118, n37119, n37120, n37121, n37122, n37123, n37124, n37125, n37126,
    n37127, n37128, n37129, n37130, n37131, n37132, n37133, n37134, n37135,
    n37136, n37137, n37138, n37139, n37140, n37141, n37142, n37143, n37144,
    n37145, n37146, n37147, n37148, n37149, n37150, n37151, n37152, n37153,
    n37154, n37155, n37156, n37157, n37158, n37159, n37160, n37161, n37163,
    n37164, n37165, n37166, n37167, n37168, n37169, n37170, n37171, n37172,
    n37173, n37174, n37175, n37176, n37177, n37178, n37179, n37180, n37181,
    n37182, n37183, n37184, n37185, n37186, n37187, n37188, n37189, n37190,
    n37191, n37192, n37193, n37194, n37195, n37196, n37197, n37198, n37199,
    n37200, n37201, n37202, n37203, n37204, n37205, n37206, n37207, n37208,
    n37209, n37210, n37211, n37212, n37213, n37214, n37215, n37216, n37217,
    n37218, n37219, n37220, n37221, n37222, n37223, n37224, n37225, n37226,
    n37227, n37228, n37229, n37230, n37231, n37232, n37233, n37234, n37235,
    n37236, n37237, n37238, n37239, n37240, n37241, n37242, n37243, n37244,
    n37245, n37246, n37247, n37248, n37249, n37250, n37251, n37252, n37253,
    n37254, n37255, n37256, n37257, n37258, n37259, n37260, n37261, n37262,
    n37263, n37264, n37265, n37266, n37267, n37268, n37270, n37271, n37272,
    n37273, n37274, n37275, n37276, n37277, n37278, n37279, n37280, n37281,
    n37282, n37283, n37284, n37285, n37286, n37287, n37288, n37289, n37290,
    n37291, n37292, n37293, n37294, n37295, n37296, n37297, n37298, n37299,
    n37300, n37301, n37302, n37303, n37304, n37305, n37306, n37307, n37308,
    n37310, n37311, n37312, n37313, n37314, n37315, n37316, n37317, n37318,
    n37319, n37320, n37321, n37322, n37323, n37324, n37325, n37326, n37327,
    n37328, n37329, n37330, n37331, n37332, n37333, n37334, n37335, n37336,
    n37337, n37338, n37339, n37340, n37341, n37342, n37343, n37344, n37345,
    n37346, n37347, n37348, n37349, n37350, n37351, n37352, n37353, n37354,
    n37355, n37356, n37357, n37358, n37359, n37360, n37362, n37363, n37364,
    n37365, n37366, n37367, n37368, n37369, n37370, n37371, n37372, n37373,
    n37374, n37375, n37376, n37377, n37378, n37379, n37380, n37381, n37382,
    n37383, n37384, n37385, n37386, n37387, n37388, n37389, n37390, n37391,
    n37392, n37393, n37394, n37395, n37396, n37397, n37398, n37399, n37400,
    n37401, n37402, n37403, n37404, n37405, n37406, n37407, n37408, n37409,
    n37410, n37411, n37412, n37413, n37414, n37415, n37416, n37417, n37418,
    n37419, n37420, n37421, n37422, n37423, n37424, n37425, n37426, n37427,
    n37428, n37429, n37430, n37431, n37432, n37433, n37434, n37435, n37436,
    n37437, n37438, n37439, n37440, n37441, n37442, n37443, n37444, n37445,
    n37446, n37447, n37448, n37449, n37450, n37451, n37452, n37453, n37454,
    n37455, n37456, n37457, n37458, n37459, n37460, n37461, n37462, n37463,
    n37464, n37465, n37466, n37468, n37469, n37470, n37471, n37472, n37473,
    n37474, n37475, n37476, n37477, n37478, n37479, n37480, n37481, n37482,
    n37483, n37484, n37485, n37486, n37487, n37488, n37489, n37490, n37491,
    n37492, n37493, n37494, n37495, n37496, n37497, n37498, n37499, n37500,
    n37501, n37502, n37503, n37504, n37505, n37506, n37507, n37508, n37509,
    n37510, n37511, n37512, n37513, n37514, n37515, n37516, n37517, n37518,
    n37519, n37520, n37521, n37522, n37523, n37524, n37525, n37526, n37527,
    n37528, n37529, n37530, n37531, n37532, n37533, n37534, n37535, n37536,
    n37537, n37538, n37539, n37540, n37541, n37542, n37543, n37544, n37545,
    n37546, n37547, n37548, n37549, n37550, n37551, n37552, n37553, n37554,
    n37555, n37556, n37557, n37558, n37559, n37560, n37561, n37562, n37563,
    n37564, n37565, n37566, n37567, n37568, n37569, n37570, n37571, n37572,
    n37573, n37574, n37576, n37577, n37578, n37579, n37580, n37581, n37582,
    n37583, n37584, n37585, n37586, n37587, n37588, n37589, n37590, n37591,
    n37592, n37593, n37594, n37595, n37596, n37597, n37598, n37599, n37600,
    n37601, n37602, n37603, n37604, n37605, n37606, n37607, n37608, n37609,
    n37610, n37611, n37612, n37613, n37614, n37615, n37616, n37617, n37618,
    n37619, n37620, n37621, n37622, n37623, n37624, n37625, n37626, n37627,
    n37628, n37629, n37630, n37631, n37632, n37633, n37634, n37635, n37636,
    n37637, n37638, n37639, n37640, n37641, n37642, n37643, n37644, n37645,
    n37646, n37647, n37648, n37649, n37650, n37651, n37652, n37653, n37654,
    n37655, n37656, n37657, n37658, n37659, n37660, n37661, n37662, n37663,
    n37664, n37665, n37666, n37667, n37668, n37669, n37670, n37671, n37672,
    n37673, n37674, n37675, n37676, n37677, n37679, n37680, n37681, n37682,
    n37683, n37684, n37685, n37686, n37687, n37688, n37689, n37690, n37691,
    n37692, n37693, n37694, n37695, n37696, n37697, n37698, n37699, n37700,
    n37701, n37702, n37703, n37704, n37705, n37706, n37707, n37708, n37709,
    n37710, n37711, n37712, n37713, n37714, n37715, n37716, n37717, n37719,
    n37720, n37721, n37722, n37723, n37724, n37725, n37726, n37727, n37728,
    n37729, n37730, n37731, n37732, n37733, n37734, n37735, n37736, n37737,
    n37738, n37739, n37740, n37741, n37742, n37743, n37744, n37745, n37746,
    n37747, n37748, n37749, n37750, n37751, n37752, n37753, n37754, n37755,
    n37756, n37757, n37758, n37759, n37760, n37761, n37762, n37763, n37764,
    n37765, n37766, n37767, n37768, n37769, n37770, n37771, n37772, n37773,
    n37774, n37775, n37776, n37777, n37778, n37779, n37780, n37781, n37782,
    n37783, n37784, n37785, n37786, n37787, n37788, n37789, n37790, n37791,
    n37792, n37793, n37794, n37795, n37796, n37797, n37798, n37799, n37800,
    n37801, n37802, n37803, n37804, n37805, n37806, n37807, n37808, n37809,
    n37810, n37811, n37812, n37813, n37814, n37815, n37816, n37817, n37818,
    n37820, n37821, n37822, n37823, n37824, n37825, n37826, n37827, n37828,
    n37829, n37830, n37831, n37832, n37833, n37834, n37835, n37836, n37837,
    n37838, n37839, n37840, n37841, n37842, n37843, n37844, n37845, n37846,
    n37847, n37848, n37849, n37850, n37851, n37852, n37853, n37854, n37855,
    n37856, n37857, n37858, n37859, n37861, n37862, n37863, n37864, n37865,
    n37866, n37867, n37868, n37869, n37870, n37871, n37872, n37873, n37874,
    n37875, n37876, n37877, n37878, n37879, n37880, n37881, n37882, n37883,
    n37884, n37885, n37886, n37887, n37888, n37889, n37890, n37891, n37892,
    n37893, n37894, n37895, n37896, n37897, n37898, n37900, n37901, n37902,
    n37903, n37904, n37905, n37906, n37907, n37908, n37909, n37910, n37911,
    n37912, n37913, n37914, n37915, n37916, n37917, n37918, n37919, n37920,
    n37921, n37922, n37923, n37924, n37925, n37926, n37927, n37928, n37929,
    n37930, n37931, n37932, n37933, n37934, n37935, n37936, n37937, n37938,
    n37940, n37941, n37942, n37943, n37944, n37945, n37946, n37947, n37948,
    n37949, n37950, n37951, n37952, n37953, n37954, n37955, n37956, n37957,
    n37958, n37959, n37960, n37961, n37962, n37963, n37964, n37965, n37966,
    n37967, n37968, n37969, n37970, n37971, n37972, n37973, n37974, n37975,
    n37976, n37977, n37978, n37979, n37981, n37982, n37983, n37984, n37985,
    n37986, n37987, n37988, n37989, n37990, n37991, n37992, n37993, n37994,
    n37995, n37996, n37997, n37998, n37999, n38000, n38001, n38002, n38003,
    n38004, n38005, n38006, n38007, n38008, n38009, n38010, n38011, n38013,
    n38014, n38015, n38016, n38017, n38018, n38019, n38020, n38021, n38022,
    n38023, n38024, n38025, n38026, n38027, n38028, n38029, n38030, n38031,
    n38032, n38033, n38034, n38035, n38036, n38037, n38038, n38039, n38040,
    n38041, n38042, n38043, n38044, n38045, n38046, n38047, n38048, n38049,
    n38050, n38051, n38052, n38053, n38054, n38055, n38056, n38057, n38058,
    n38060, n38061, n38062, n38063, n38064, n38065, n38066, n38067, n38068,
    n38069, n38070, n38071, n38072, n38073, n38074, n38075, n38076, n38077,
    n38078, n38079, n38080, n38081, n38082, n38083, n38084, n38085, n38086,
    n38087, n38088, n38089, n38090, n38091, n38092, n38093, n38094, n38095,
    n38096, n38097, n38098, n38099, n38100, n38101, n38103, n38104, n38105,
    n38106, n38107, n38108, n38109, n38110, n38111, n38112, n38113, n38114,
    n38115, n38116, n38117, n38118, n38119, n38120, n38121, n38122, n38123,
    n38124, n38125, n38126, n38127, n38128, n38129, n38130, n38131, n38132,
    n38133, n38134, n38136, n38137, n38138, n38139, n38140, n38141, n38142,
    n38143, n38144, n38145, n38146, n38147, n38148, n38149, n38150, n38151,
    n38152, n38153, n38154, n38155, n38156, n38157, n38158, n38159, n38160,
    n38161, n38162, n38163, n38164, n38166, n38167, n38168, n38169, n38170,
    n38171, n38172, n38173, n38174, n38175, n38176, n38177, n38178, n38179,
    n38180, n38181, n38182, n38183, n38184, n38185, n38186, n38187, n38188,
    n38189, n38190, n38191, n38192, n38193, n38194, n38195, n38197, n38198,
    n38199, n38200, n38201, n38202, n38203, n38204, n38205, n38206, n38207,
    n38208, n38209, n38210, n38211, n38212, n38213, n38214, n38215, n38216,
    n38217, n38218, n38219, n38220, n38221, n38222, n38223, n38225, n38226,
    n38227, n38228, n38229, n38230, n38231, n38232, n38233, n38234, n38235,
    n38236, n38237, n38238, n38239, n38240, n38241, n38242, n38243, n38244,
    n38245, n38246, n38247, n38248, n38249, n38250, n38251, n38252, n38253,
    n38254, n38255, n38256, n38257, n38258, n38259, n38260, n38261, n38262,
    n38263, n38264, n38265, n38267, n38268, n38269, n38270, n38271, n38272,
    n38273, n38274, n38275, n38276, n38277, n38278, n38279, n38280, n38281,
    n38282, n38283, n38284, n38285, n38286, n38287, n38288, n38289, n38290,
    n38291, n38292, n38293, n38294, n38295, n38296, n38297, n38298, n38299,
    n38300, n38301, n38302, n38304, n38305, n38306, n38307, n38308, n38309,
    n38310, n38311, n38312, n38313, n38314, n38315, n38316, n38317, n38318,
    n38319, n38320, n38321, n38322, n38323, n38324, n38325, n38326, n38327,
    n38328, n38329, n38330, n38331, n38332, n38333, n38334, n38335, n38336,
    n38337, n38338, n38339, n38340, n38341, n38342, n38343, n38344, n38346,
    n38347, n38348, n38349, n38350, n38351, n38352, n38353, n38354, n38355,
    n38356, n38357, n38358, n38359, n38360, n38361, n38362, n38363, n38364,
    n38365, n38366, n38367, n38368, n38369, n38370, n38371, n38372, n38373,
    n38374, n38375, n38376, n38377, n38378, n38379, n38380, n38382, n38383,
    n38384, n38385, n38386, n38387, n38388, n38389, n38390, n38391, n38392,
    n38393, n38394, n38395, n38396, n38397, n38398, n38399, n38400, n38401,
    n38402, n38403, n38404, n38405, n38406, n38407, n38408, n38409, n38410,
    n38411, n38412, n38413, n38414, n38415, n38416, n38418, n38419, n38420,
    n38421, n38422, n38423, n38424, n38425, n38426, n38427, n38428, n38429,
    n38430, n38431, n38432, n38433, n38434, n38435, n38436, n38437, n38438,
    n38439, n38440, n38441, n38442, n38443, n38444, n38445, n38446, n38447,
    n38448, n38449, n38450, n38451, n38452, n38453, n38454, n38455, n38456,
    n38457, n38459, n38460, n38461, n38462, n38463, n38464, n38465, n38466,
    n38467, n38468, n38469, n38470, n38471, n38472, n38473, n38474, n38475,
    n38476, n38477, n38478, n38479, n38480, n38481, n38482, n38483, n38484,
    n38485, n38486, n38487, n38488, n38489, n38490, n38491, n38492, n38493,
    n38495, n38496, n38497, n38498, n38499, n38500, n38501, n38502, n38503,
    n38504, n38505, n38506, n38507, n38508, n38509, n38510, n38511, n38512,
    n38513, n38514, n38515, n38516, n38517, n38518, n38519, n38520, n38521,
    n38522, n38523, n38524, n38525, n38526, n38527, n38528, n38529, n38530,
    n38531, n38532, n38533, n38534, n38535, n38536, n38537, n38538, n38539,
    n38540, n38541, n38542, n38543, n38544, n38545, n38546, n38547, n38548,
    n38549, n38550, n38551, n38552, n38553, n38554, n38555, n38556, n38557,
    n38558, n38559, n38560, n38561, n38562, n38563, n38564, n38565, n38566,
    n38567, n38568, n38569, n38570, n38571, n38572, n38573, n38574, n38575,
    n38576, n38577, n38578, n38579, n38580, n38581, n38582, n38583, n38584,
    n38585, n38586, n38588, n38589, n38590, n38591, n38592, n38593, n38594,
    n38595, n38596, n38597, n38598, n38599, n38600, n38601, n38602, n38603,
    n38604, n38605, n38606, n38607, n38608, n38609, n38610, n38611, n38612,
    n38613, n38614, n38615, n38616, n38617, n38618, n38619, n38620, n38621,
    n38622, n38623, n38624, n38625, n38626, n38627, n38628, n38629, n38630,
    n38631, n38632, n38633, n38635, n38636, n38637, n38638, n38639, n38640,
    n38641, n38642, n38643, n38644, n38645, n38646, n38647, n38648, n38649,
    n38650, n38651, n38652, n38653, n38654, n38655, n38656, n38657, n38658,
    n38659, n38660, n38661, n38662, n38663, n38664, n38665, n38666, n38667,
    n38668, n38669, n38671, n38672, n38673, n38674, n38675, n38676, n38677,
    n38678, n38679, n38680, n38681, n38682, n38683, n38684, n38685, n38686,
    n38687, n38688, n38689, n38690, n38691, n38692, n38693, n38694, n38695,
    n38696, n38697, n38698, n38699, n38700, n38701, n38702, n38703, n38704,
    n38705, n38706, n38707, n38709, n38710, n38711, n38712, n38713, n38714,
    n38715, n38716, n38717, n38718, n38719, n38720, n38721, n38722, n38723,
    n38724, n38725, n38726, n38727, n38728, n38729, n38730, n38731, n38732,
    n38733, n38734, n38735, n38736, n38737, n38738, n38739, n38740, n38741,
    n38742, n38743, n38744, n38745, n38746, n38747, n38748, n38749, n38750,
    n38751, n38752, n38753, n38754, n38755, n38756, n38757, n38758, n38759,
    n38760, n38761, n38762, n38763, n38764, n38765, n38766, n38767, n38768,
    n38769, n38770, n38771, n38772, n38773, n38774, n38775, n38776, n38777,
    n38778, n38779, n38780, n38781, n38782, n38783, n38784, n38785, n38786,
    n38787, n38788, n38789, n38790, n38791, n38792, n38793, n38794, n38795,
    n38796, n38797, n38798, n38799, n38800, n38801, n38802, n38803, n38804,
    n38805, n38806, n38807, n38808, n38809, n38810, n38811, n38813, n38814,
    n38815, n38816, n38817, n38818, n38819, n38820, n38821, n38822, n38823,
    n38824, n38825, n38826, n38827, n38828, n38829, n38830, n38831, n38832,
    n38833, n38834, n38835, n38836, n38837, n38838, n38839, n38840, n38841,
    n38842, n38843, n38844, n38845, n38846, n38847, n38848, n38849, n38850,
    n38851, n38852, n38853, n38854, n38855, n38856, n38857, n38858, n38859,
    n38860, n38861, n38862, n38863, n38864, n38865, n38866, n38867, n38868,
    n38869, n38870, n38871, n38872, n38873, n38874, n38875, n38876, n38877,
    n38878, n38879, n38880, n38881, n38882, n38883, n38884, n38885, n38886,
    n38887, n38888, n38889, n38890, n38891, n38892, n38893, n38894, n38895,
    n38896, n38897, n38898, n38899, n38900, n38901, n38902, n38903, n38904,
    n38905, n38906, n38907, n38908, n38909, n38910, n38911, n38912, n38913,
    n38914, n38915, n38917, n38918, n38919, n38920, n38921, n38922, n38923,
    n38924, n38925, n38926, n38927, n38928, n38929, n38930, n38931, n38932,
    n38933, n38934, n38935, n38936, n38937, n38938, n38939, n38940, n38941,
    n38942, n38943, n38944, n38945, n38946, n38947, n38948, n38949, n38950,
    n38951, n38952, n38953, n38954, n38955, n38956, n38957, n38958, n38959,
    n38960, n38961, n38962, n38963, n38964, n38965, n38966, n38967, n38968,
    n38969, n38970, n38971, n38972, n38973, n38974, n38975, n38976, n38977,
    n38978, n38979, n38980, n38981, n38982, n38983, n38984, n38985, n38986,
    n38987, n38988, n38989, n38990, n38991, n38992, n38993, n38994, n38995,
    n38996, n38997, n38998, n38999, n39000, n39001, n39002, n39003, n39004,
    n39005, n39006, n39007, n39008, n39009, n39010, n39011, n39012, n39013,
    n39014, n39015, n39017, n39018, n39019, n39020, n39021, n39022, n39023,
    n39024, n39025, n39026, n39027, n39028, n39029, n39030, n39031, n39032,
    n39033, n39034, n39035, n39036, n39037, n39038, n39039, n39040, n39041,
    n39042, n39043, n39044, n39045, n39046, n39047, n39048, n39049, n39050,
    n39051, n39052, n39053, n39054, n39055, n39056, n39057, n39058, n39059,
    n39060, n39061, n39062, n39063, n39064, n39065, n39066, n39067, n39068,
    n39069, n39070, n39071, n39072, n39073, n39074, n39075, n39076, n39077,
    n39078, n39079, n39080, n39081, n39082, n39083, n39084, n39085, n39086,
    n39087, n39088, n39089, n39090, n39091, n39092, n39093, n39094, n39095,
    n39096, n39097, n39098, n39099, n39100, n39101, n39102, n39103, n39104,
    n39105, n39106, n39107, n39108, n39109, n39110, n39111, n39112, n39113,
    n39114, n39115, n39116, n39117, n39118, n39119, n39120, n39121, n39123,
    n39124, n39125, n39126, n39127, n39128, n39129, n39130, n39131, n39132,
    n39133, n39134, n39135, n39136, n39137, n39138, n39139, n39140, n39141,
    n39142, n39143, n39144, n39145, n39146, n39147, n39148, n39149, n39150,
    n39151, n39152, n39153, n39154, n39156, n39157, n39158, n39159, n39160,
    n39161, n39162, n39163, n39164, n39165, n39166, n39167, n39168, n39169,
    n39170, n39171, n39172, n39173, n39174, n39175, n39176, n39177, n39178,
    n39179, n39180, n39181, n39182, n39183, n39184, n39185, n39186, n39187,
    n39188, n39189, n39190, n39191, n39192, n39193, n39194, n39195, n39196,
    n39197, n39198, n39199, n39200, n39201, n39202, n39203, n39205, n39206,
    n39207, n39208, n39209, n39210, n39211, n39212, n39213, n39214, n39215,
    n39216, n39217, n39218, n39219, n39220, n39221, n39222, n39223, n39224,
    n39225, n39226, n39227, n39228, n39229, n39230, n39231, n39232, n39233,
    n39234, n39235, n39236, n39237, n39238, n39239, n39240, n39241, n39242,
    n39243, n39244, n39245, n39246, n39247, n39248, n39249, n39250, n39251,
    n39252, n39253, n39254, n39255, n39256, n39257, n39258, n39259, n39260,
    n39261, n39262, n39263, n39264, n39265, n39266, n39267, n39268, n39269,
    n39270, n39271, n39272, n39273, n39274, n39275, n39276, n39277, n39278,
    n39279, n39280, n39281, n39282, n39283, n39284, n39285, n39286, n39287,
    n39288, n39289, n39290, n39291, n39292, n39293, n39294, n39296, n39297,
    n39298, n39299, n39300, n39301, n39302, n39303, n39304, n39305, n39306,
    n39307, n39308, n39309, n39310, n39311, n39312, n39313, n39314, n39315,
    n39316, n39317, n39318, n39319, n39320, n39321, n39322, n39323, n39324,
    n39325, n39326, n39327, n39328, n39329, n39330, n39331, n39333, n39334,
    n39335, n39336, n39337, n39338, n39339, n39340, n39341, n39342, n39343,
    n39344, n39345, n39346, n39347, n39348, n39349, n39350, n39351, n39352,
    n39353, n39354, n39355, n39356, n39357, n39358, n39359, n39360, n39361,
    n39362, n39363, n39364, n39365, n39366, n39367, n39368, n39369, n39370,
    n39371, n39372, n39373, n39374, n39375, n39377, n39378, n39379, n39380,
    n39381, n39382, n39383, n39384, n39385, n39386, n39387, n39388, n39389,
    n39390, n39391, n39392, n39393, n39394, n39395, n39396, n39397, n39398,
    n39399, n39400, n39401, n39402, n39403, n39404, n39405, n39406, n39407,
    n39408, n39409, n39410, n39411, n39412, n39413, n39414, n39415, n39416,
    n39418, n39419, n39420, n39421, n39422, n39423, n39424, n39425, n39426,
    n39427, n39428, n39429, n39430, n39431, n39432, n39433, n39434, n39435,
    n39436, n39437, n39438, n39439, n39440, n39441, n39442, n39443, n39444,
    n39445, n39446, n39447, n39448, n39449, n39450, n39451, n39452, n39453,
    n39454, n39455, n39456, n39457, n39458, n39459, n39460, n39461, n39462,
    n39463, n39464, n39465, n39466, n39467, n39468, n39469, n39470, n39471,
    n39472, n39473, n39474, n39475, n39476, n39477, n39478, n39479, n39480,
    n39481, n39482, n39483, n39484, n39485, n39486, n39487, n39488, n39489,
    n39490, n39491, n39492, n39493, n39494, n39495, n39496, n39497, n39498,
    n39499, n39500, n39501, n39502, n39503, n39504, n39505, n39506, n39507,
    n39508, n39509, n39510, n39511, n39512, n39513, n39514, n39515, n39516,
    n39517, n39518, n39519, n39520, n39522, n39523, n39524, n39525, n39526,
    n39527, n39528, n39529, n39530, n39531, n39532, n39533, n39534, n39535,
    n39536, n39537, n39538, n39539, n39540, n39541, n39542, n39543, n39544,
    n39545, n39546, n39547, n39548, n39549, n39550, n39551, n39552, n39553,
    n39554, n39555, n39556, n39557, n39558, n39559, n39560, n39561, n39562,
    n39563, n39564, n39565, n39566, n39567, n39568, n39569, n39570, n39571,
    n39572, n39574, n39575, n39576, n39577, n39578, n39579, n39580, n39581,
    n39582, n39583, n39584, n39585, n39586, n39587, n39588, n39589, n39590,
    n39591, n39592, n39593, n39594, n39595, n39596, n39597, n39598, n39599,
    n39600, n39601, n39602, n39603, n39604, n39605, n39606, n39607, n39608,
    n39609, n39611, n39612, n39613, n39614, n39615, n39616, n39617, n39618,
    n39619, n39620, n39621, n39622, n39623, n39624, n39625, n39626, n39627,
    n39628, n39629, n39630, n39631, n39632, n39633, n39634, n39635, n39636,
    n39637, n39638, n39639, n39640, n39641, n39642, n39643, n39644, n39645,
    n39646, n39648, n39649, n39650, n39651, n39652, n39653, n39654, n39655,
    n39656, n39657, n39658, n39659, n39660, n39661, n39662, n39663, n39664,
    n39665, n39666, n39667, n39668, n39669, n39670, n39671, n39672, n39673,
    n39674, n39675, n39676, n39677, n39678, n39679, n39680, n39681, n39682,
    n39683, n39684, n39685, n39686, n39687, n39688, n39689, n39690, n39691,
    n39692, n39693, n39694, n39695, n39696, n39697, n39698, n39699, n39700,
    n39701, n39702, n39703, n39704, n39705, n39706, n39707, n39708, n39709,
    n39710, n39711, n39712, n39713, n39714, n39715, n39716, n39717, n39718,
    n39719, n39720, n39721, n39722, n39723, n39724, n39725, n39726, n39727,
    n39728, n39729, n39730, n39731, n39732, n39733, n39734, n39735, n39736,
    n39737, n39738, n39739, n39740, n39741, n39742, n39744, n39745, n39746,
    n39747, n39748, n39749, n39750, n39751, n39752, n39753, n39754, n39755,
    n39756, n39757, n39758, n39759, n39760, n39761, n39762, n39763, n39764,
    n39765, n39766, n39767, n39768, n39769, n39770, n39771, n39772, n39774,
    n39775, n39776, n39777, n39778, n39779, n39780, n39781, n39782, n39783,
    n39784, n39785, n39786, n39787, n39788, n39789, n39790, n39791, n39792,
    n39793, n39794, n39795, n39796, n39797, n39798, n39799, n39800, n39801,
    n39802, n39803, n39804, n39805, n39806, n39807, n39808, n39809, n39810,
    n39811, n39812, n39813, n39814, n39815, n39816, n39817, n39818, n39819,
    n39820, n39821, n39823, n39824, n39825, n39826, n39827, n39828, n39829,
    n39830, n39831, n39832, n39833, n39834, n39835, n39836, n39837, n39838,
    n39839, n39840, n39841, n39842, n39843, n39844, n39845, n39846, n39847,
    n39848, n39849, n39850, n39851, n39852, n39853, n39854, n39855, n39856,
    n39857, n39858, n39859, n39861, n39862, n39863, n39864, n39865, n39866,
    n39867, n39868, n39869, n39870, n39871, n39872, n39873, n39874, n39875,
    n39876, n39877, n39878, n39879, n39880, n39881, n39882, n39883, n39884,
    n39885, n39886, n39887, n39888, n39889, n39890, n39891, n39892, n39893,
    n39894, n39895, n39896, n39897, n39898, n39899, n39900, n39901, n39902,
    n39904, n39905, n39906, n39907, n39908, n39909, n39910, n39911, n39912,
    n39913, n39914, n39915, n39916, n39917, n39918, n39919, n39920, n39921,
    n39922, n39923, n39924, n39925, n39926, n39927, n39928, n39929, n39930,
    n39931, n39932, n39933, n39934, n39935, n39936, n39937, n39938, n39939,
    n39940, n39941, n39942, n39943, n39944, n39945, n39946, n39947, n39948,
    n39949, n39951, n39952, n39953, n39954, n39955, n39956, n39957, n39958,
    n39959, n39960, n39961, n39962, n39963, n39964, n39965, n39966, n39967,
    n39968, n39969, n39970, n39971, n39972, n39973, n39974, n39975, n39976,
    n39977, n39978, n39979, n39980, n39981, n39982, n39983, n39984, n39985,
    n39987, n39988, n39989, n39990, n39991, n39992, n39993, n39994, n39995,
    n39996, n39997, n39998, n39999, n40000, n40001, n40002, n40003, n40004,
    n40005, n40006, n40007, n40008, n40009, n40010, n40011, n40012, n40013,
    n40014, n40015, n40016, n40017, n40018, n40019, n40020, n40021, n40022,
    n40023, n40024, n40025, n40026, n40027, n40028, n40029, n40030, n40031,
    n40032, n40033, n40034, n40035, n40036, n40037, n40038, n40039, n40040,
    n40041, n40042, n40043, n40044, n40045, n40046, n40047, n40048, n40049,
    n40050, n40051, n40052, n40053, n40054, n40055, n40056, n40057, n40058,
    n40059, n40060, n40061, n40062, n40063, n40064, n40065, n40066, n40067,
    n40068, n40069, n40070, n40071, n40072, n40073, n40074, n40075, n40076,
    n40077, n40078, n40079, n40080, n40081, n40082, n40083, n40084, n40086,
    n40087, n40088, n40089, n40090, n40091, n40092, n40093, n40094, n40095,
    n40096, n40097, n40098, n40099, n40100, n40101, n40102, n40103, n40104,
    n40105, n40106, n40107, n40108, n40109, n40110, n40111, n40112, n40113,
    n40114, n40115, n40116, n40117, n40118, n40119, n40120, n40121, n40122,
    n40123, n40124, n40126, n40127, n40128, n40129, n40130, n40131, n40132,
    n40133, n40134, n40135, n40136, n40137, n40138, n40139, n40140, n40141,
    n40142, n40143, n40144, n40145, n40146, n40147, n40148, n40149, n40150,
    n40151, n40152, n40153, n40154, n40155, n40157, n40158, n40159, n40160,
    n40161, n40162, n40163, n40164, n40165, n40166, n40167, n40168, n40169,
    n40170, n40171, n40172, n40173, n40174, n40175, n40176, n40177, n40178,
    n40179, n40180, n40181, n40182, n40183, n40184, n40185, n40186, n40187,
    n40188, n40189, n40190, n40191, n40192, n40193, n40194, n40195, n40196,
    n40197, n40198, n40199, n40200, n40202, n40203, n40204, n40205, n40206,
    n40207, n40208, n40209, n40210, n40211, n40212, n40213, n40214, n40215,
    n40216, n40217, n40218, n40219, n40220, n40221, n40222, n40223, n40224,
    n40225, n40226, n40227, n40228, n40229, n40230, n40231, n40232, n40233,
    n40234, n40235, n40236, n40237, n40239, n40240, n40241, n40242, n40243,
    n40244, n40245, n40246, n40247, n40248, n40249, n40250, n40251, n40252,
    n40253, n40254, n40255, n40256, n40257, n40258, n40259, n40260, n40261,
    n40262, n40263, n40264, n40265, n40266, n40267, n40268, n40269, n40270,
    n40272, n40273, n40274, n40275, n40276, n40277, n40278, n40279, n40280,
    n40281, n40282, n40283, n40284, n40285, n40286, n40287, n40288, n40289,
    n40290, n40291, n40292, n40293, n40294, n40295, n40296, n40297, n40298,
    n40299, n40300, n40301, n40302, n40303, n40304, n40305, n40306, n40308,
    n40309, n40310, n40311, n40312, n40313, n40314, n40315, n40316, n40317,
    n40318, n40319, n40320, n40321, n40322, n40323, n40324, n40325, n40326,
    n40327, n40328, n40329, n40330, n40331, n40332, n40333, n40334, n40335,
    n40336, n40337, n40338, n40339, n40340, n40341, n40342, n40344, n40345,
    n40346, n40347, n40348, n40349, n40350, n40351, n40352, n40353, n40354,
    n40355, n40356, n40357, n40358, n40359, n40360, n40361, n40362, n40363,
    n40364, n40365, n40366, n40367, n40368, n40369, n40370, n40371, n40372,
    n40373, n40374, n40375, n40376, n40377, n40379, n40380, n40381, n40382,
    n40383, n40384, n40385, n40386, n40387, n40388, n40389, n40390, n40391,
    n40392, n40393, n40394, n40395, n40396, n40397, n40398, n40399, n40400,
    n40401, n40402, n40403, n40404, n40405, n40406, n40407, n40408, n40409,
    n40410, n40411, n40412, n40413, n40415, n40416, n40417, n40418, n40419,
    n40420, n40421, n40422, n40423, n40424, n40425, n40426, n40427, n40428,
    n40429, n40430, n40431, n40432, n40433, n40434, n40435, n40436, n40437,
    n40438, n40439, n40440, n40441, n40442, n40443, n40445, n40446, n40447,
    n40448, n40449, n40450, n40451, n40452, n40453, n40454, n40455, n40456,
    n40457, n40458, n40459, n40460, n40461, n40462, n40463, n40464, n40465,
    n40466, n40467, n40468, n40469, n40470, n40471, n40472, n40473, n40474,
    n40475, n40476, n40477, n40478, n40479, n40480, n40481, n40482, n40483,
    n40484, n40485, n40486, n40487, n40488, n40489, n40490, n40491, n40492,
    n40493, n40494, n40495, n40496, n40497, n40498, n40499, n40500, n40501,
    n40502, n40503, n40504, n40505, n40506, n40507, n40508, n40509, n40510,
    n40511, n40512, n40513, n40514, n40515, n40516, n40517, n40518, n40519,
    n40520, n40521, n40522, n40523, n40524, n40525, n40526, n40527, n40528,
    n40529, n40530, n40531, n40532, n40533, n40534, n40535, n40536, n40537,
    n40538, n40539, n40540, n40541, n40542, n40543, n40544, n40546, n40547,
    n40548, n40549, n40550, n40551, n40552, n40553, n40554, n40555, n40556,
    n40557, n40558, n40559, n40560, n40561, n40562, n40563, n40564, n40565,
    n40566, n40567, n40568, n40569, n40570, n40571, n40572, n40573, n40574,
    n40575, n40576, n40577, n40578, n40579, n40580, n40581, n40582, n40583,
    n40584, n40585, n40586, n40587, n40588, n40589, n40590, n40591, n40592,
    n40593, n40594, n40595, n40596, n40597, n40598, n40599, n40600, n40601,
    n40602, n40603, n40604, n40605, n40606, n40607, n40608, n40609, n40610,
    n40611, n40612, n40613, n40614, n40615, n40616, n40617, n40618, n40619,
    n40620, n40621, n40622, n40623, n40624, n40625, n40626, n40627, n40628,
    n40629, n40630, n40631, n40632, n40633, n40634, n40635, n40636, n40637,
    n40638, n40639, n40640, n40641, n40642, n40643, n40644, n40645, n40646,
    n40647, n40648, n40650, n40651, n40652, n40653, n40654, n40655, n40656,
    n40657, n40658, n40659, n40660, n40661, n40662, n40663, n40664, n40665,
    n40666, n40667, n40668, n40669, n40670, n40671, n40672, n40673, n40674,
    n40675, n40676, n40677, n40678, n40679, n40680, n40681, n40682, n40683,
    n40684, n40685, n40686, n40687, n40688, n40689, n40690, n40691, n40693,
    n40694, n40695, n40696, n40697, n40698, n40699, n40700, n40701, n40702,
    n40703, n40704, n40705, n40706, n40707, n40708, n40709, n40710, n40711,
    n40712, n40713, n40714, n40715, n40716, n40717, n40718, n40719, n40720,
    n40721, n40722, n40723, n40724, n40725, n40726, n40727, n40728, n40729,
    n40730, n40731, n40732, n40733, n40734, n40735, n40736, n40737, n40738,
    n40739, n40740, n40741, n40742, n40743, n40744, n40745, n40746, n40747,
    n40748, n40749, n40750, n40751, n40752, n40753, n40754, n40755, n40756,
    n40757, n40758, n40759, n40760, n40761, n40762, n40763, n40764, n40765,
    n40766, n40767, n40768, n40769, n40770, n40771, n40772, n40773, n40774,
    n40775, n40776, n40777, n40778, n40779, n40780, n40781, n40782, n40783,
    n40784, n40785, n40786, n40787, n40788, n40789, n40790, n40791, n40792,
    n40793, n40794, n40795, n40796, n40798, n40799, n40800, n40801, n40802,
    n40803, n40804, n40805, n40806, n40807, n40808, n40809, n40810, n40811,
    n40812, n40813, n40814, n40815, n40816, n40817, n40818, n40819, n40820,
    n40821, n40822, n40823, n40824, n40825, n40826, n40827, n40828, n40829,
    n40830, n40831, n40832, n40833, n40834, n40835, n40836, n40837, n40838,
    n40839, n40840, n40841, n40842, n40843, n40844, n40845, n40846, n40847,
    n40848, n40849, n40850, n40851, n40852, n40853, n40854, n40855, n40856,
    n40857, n40858, n40859, n40860, n40861, n40862, n40863, n40864, n40865,
    n40866, n40867, n40868, n40869, n40870, n40871, n40872, n40873, n40874,
    n40875, n40876, n40877, n40878, n40879, n40880, n40881, n40882, n40883,
    n40884, n40885, n40886, n40887, n40888, n40890, n40891, n40892, n40893,
    n40894, n40895, n40896, n40897, n40898, n40899, n40900, n40901, n40902,
    n40903, n40904, n40905, n40906, n40907, n40908, n40909, n40910, n40911,
    n40912, n40913, n40914, n40915, n40916, n40917, n40918, n40919, n40920,
    n40921, n40923, n40924, n40925, n40926, n40927, n40928, n40929, n40930,
    n40931, n40932, n40933, n40934, n40935, n40936, n40937, n40938, n40939,
    n40940, n40941, n40942, n40943, n40944, n40945, n40946, n40947, n40948,
    n40949, n40950, n40951, n40952, n40953, n40954, n40955, n40956, n40957,
    n40958, n40959, n40960, n40961, n40962, n40963, n40964, n40965, n40966,
    n40967, n40968, n40969, n40970, n40971, n40972, n40973, n40974, n40975,
    n40976, n40977, n40978, n40979, n40980, n40981, n40982, n40983, n40984,
    n40985, n40986, n40987, n40988, n40989, n40990, n40991, n40992, n40993,
    n40994, n40995, n40996, n40997, n40998, n40999, n41000, n41001, n41002,
    n41003, n41004, n41005, n41006, n41007, n41008, n41009, n41010, n41011,
    n41012, n41013, n41014, n41015, n41016, n41017, n41018, n41019, n41020,
    n41022, n41023, n41024, n41025, n41026, n41027, n41028, n41029, n41030,
    n41031, n41032, n41033, n41034, n41035, n41036, n41037, n41038, n41039,
    n41040, n41041, n41042, n41043, n41044, n41045, n41046, n41047, n41048,
    n41049, n41050, n41051, n41052, n41053, n41054, n41055, n41056, n41057,
    n41058, n41059, n41060, n41061, n41062, n41063, n41064, n41065, n41066,
    n41067, n41068, n41069, n41070, n41071, n41072, n41073, n41074, n41075,
    n41076, n41077, n41078, n41079, n41080, n41081, n41082, n41083, n41084,
    n41085, n41086, n41087, n41088, n41089, n41090, n41091, n41092, n41093,
    n41094, n41095, n41096, n41097, n41098, n41099, n41100, n41101, n41102,
    n41103, n41104, n41105, n41106, n41107, n41108, n41109, n41110, n41111,
    n41112, n41113, n41114, n41115, n41116, n41117, n41118, n41119, n41120,
    n41121, n41122, n41123, n41124, n41125, n41126, n41128, n41129, n41130,
    n41131, n41132, n41133, n41134, n41135, n41136, n41137, n41138, n41139,
    n41140, n41141, n41142, n41143, n41144, n41145, n41146, n41147, n41148,
    n41149, n41150, n41151, n41152, n41153, n41154, n41155, n41156, n41157,
    n41158, n41159, n41161, n41162, n41163, n41164, n41165, n41166, n41167,
    n41168, n41169, n41170, n41171, n41172, n41173, n41174, n41175, n41176,
    n41177, n41178, n41179, n41180, n41181, n41182, n41183, n41184, n41185,
    n41186, n41187, n41188, n41189, n41190, n41191, n41192, n41193, n41194,
    n41195, n41196, n41197, n41198, n41199, n41200, n41201, n41202, n41203,
    n41204, n41205, n41206, n41207, n41208, n41209, n41210, n41211, n41212,
    n41213, n41214, n41215, n41216, n41217, n41218, n41219, n41220, n41221,
    n41222, n41223, n41224, n41225, n41226, n41227, n41228, n41229, n41230,
    n41231, n41232, n41233, n41234, n41235, n41236, n41237, n41238, n41239,
    n41240, n41241, n41242, n41243, n41244, n41245, n41246, n41247, n41248,
    n41249, n41250, n41251, n41252, n41253, n41254, n41255, n41256, n41257,
    n41258, n41259, n41260, n41261, n41262, n41263, n41264, n41266, n41267,
    n41268, n41269, n41270, n41271, n41272, n41273, n41274, n41275, n41276,
    n41277, n41278, n41279, n41280, n41281, n41282, n41283, n41284, n41285,
    n41286, n41287, n41288, n41289, n41290, n41291, n41292, n41293, n41294,
    n41295, n41296, n41297, n41298, n41299, n41300, n41301, n41302, n41303,
    n41304, n41305, n41306, n41307, n41308, n41309, n41310, n41311, n41312,
    n41313, n41314, n41315, n41317, n41318, n41319, n41320, n41321, n41322,
    n41323, n41324, n41325, n41326, n41327, n41328, n41329, n41330, n41331,
    n41332, n41333, n41334, n41335, n41336, n41337, n41338, n41339, n41340,
    n41341, n41342, n41343, n41344, n41345, n41346, n41347, n41348, n41349,
    n41350, n41351, n41353, n41354, n41355, n41356, n41357, n41358, n41359,
    n41360, n41361, n41362, n41363, n41364, n41365, n41366, n41367, n41368,
    n41369, n41370, n41371, n41372, n41373, n41374, n41375, n41376, n41377,
    n41378, n41379, n41380, n41381, n41382, n41383, n41384, n41385, n41386,
    n41387, n41388, n41389, n41390, n41392, n41393, n41394, n41395, n41396,
    n41397, n41398, n41399, n41400, n41401, n41402, n41403, n41404, n41405,
    n41406, n41407, n41408, n41409, n41410, n41411, n41412, n41413, n41414,
    n41415, n41416, n41417, n41418, n41419, n41420, n41421, n41422, n41423,
    n41424, n41425, n41426, n41427, n41428, n41429, n41430, n41431, n41432,
    n41433, n41435, n41436, n41437, n41438, n41439, n41440, n41441, n41442,
    n41443, n41444, n41445, n41446, n41447, n41448, n41449, n41450, n41451,
    n41452, n41453, n41454, n41455, n41456, n41457, n41458, n41459, n41460,
    n41461, n41462, n41463, n41464, n41465, n41466, n41467, n41468, n41469,
    n41470, n41471, n41472, n41473, n41474, n41476, n41477, n41478, n41479,
    n41480, n41481, n41482, n41483, n41484, n41485, n41486, n41487, n41488,
    n41489, n41490, n41491, n41492, n41493, n41494, n41495, n41496, n41497,
    n41498, n41499, n41500, n41501, n41502, n41503, n41504, n41505, n41506,
    n41507, n41508, n41509, n41510, n41511, n41512, n41513, n41514, n41515,
    n41517, n41518, n41519, n41520, n41521, n41522, n41523, n41524, n41525,
    n41526, n41527, n41528, n41529, n41530, n41531, n41532, n41533, n41534,
    n41535, n41536, n41537, n41538, n41539, n41540, n41541, n41542, n41543,
    n41544, n41545, n41546, n41547, n41548, n41549, n41550, n41551, n41552,
    n41553, n41554, n41556, n41557, n41558, n41559, n41560, n41561, n41562,
    n41563, n41564, n41565, n41566, n41567, n41568, n41569, n41570, n41571,
    n41572, n41573, n41574, n41575, n41576, n41577, n41578, n41579, n41580,
    n41581, n41582, n41583, n41584, n41585, n41586, n41587, n41588, n41589,
    n41590, n41591, n41592, n41593, n41594, n41595, n41596, n41597, n41598,
    n41599, n41600, n41601, n41602, n41604, n41605, n41606, n41607, n41608,
    n41609, n41610, n41611, n41612, n41613, n41614, n41615, n41616, n41617,
    n41618, n41619, n41620, n41621, n41622, n41623, n41624, n41625, n41626,
    n41627, n41628, n41629, n41630, n41631, n41632, n41633, n41634, n41635,
    n41636, n41637, n41638, n41639, n41640, n41642, n41643, n41644, n41645,
    n41646, n41647, n41648, n41649, n41650, n41651, n41652, n41653, n41654,
    n41655, n41656, n41657, n41658, n41659, n41660, n41661, n41662, n41663,
    n41664, n41665, n41666, n41667, n41668, n41669, n41670, n41671, n41672,
    n41673, n41674, n41675, n41676, n41677, n41678, n41679, n41680, n41681,
    n41682, n41683, n41684, n41685, n41686, n41687, n41688, n41690, n41691,
    n41692, n41693, n41694, n41695, n41696, n41697, n41698, n41699, n41700,
    n41701, n41702, n41703, n41704, n41705, n41706, n41707, n41708, n41709,
    n41710, n41711, n41712, n41713, n41714, n41715, n41716, n41717, n41718,
    n41719, n41720, n41721, n41722, n41723, n41724, n41725, n41727, n41728,
    n41729, n41730, n41731, n41732, n41733, n41734, n41735, n41736, n41737,
    n41738, n41739, n41740, n41741, n41742, n41743, n41744, n41745, n41746,
    n41747, n41748, n41749, n41750, n41751, n41752, n41753, n41754, n41755,
    n41756, n41757, n41758, n41759, n41760, n41761, n41762, n41763, n41764,
    n41765, n41767, n41768, n41769, n41770, n41771, n41772, n41773, n41774,
    n41775, n41776, n41777, n41778, n41779, n41780, n41781, n41782, n41783,
    n41784, n41785, n41786, n41787, n41788, n41789, n41790, n41791, n41792,
    n41793, n41794, n41795, n41796, n41797, n41798, n41799, n41800, n41801,
    n41802, n41803, n41804, n41805, n41806, n41807, n41808, n41809, n41810,
    n41811, n41812, n41813, n41814, n41815, n41816, n41817, n41818, n41819,
    n41820, n41821, n41822, n41823, n41824, n41825, n41826, n41827, n41828,
    n41829, n41830, n41831, n41832, n41833, n41834, n41835, n41836, n41837,
    n41838, n41839, n41840, n41841, n41842, n41843, n41844, n41845, n41846,
    n41847, n41848, n41849, n41850, n41851, n41852, n41853, n41854, n41855,
    n41856, n41857, n41858, n41860, n41861, n41862, n41863, n41864, n41865,
    n41866, n41867, n41868, n41869, n41870, n41871, n41872, n41873, n41874,
    n41875, n41876, n41877, n41878, n41879, n41880, n41881, n41882, n41883,
    n41884, n41885, n41886, n41887, n41888, n41889, n41890, n41891, n41892,
    n41893, n41894, n41896, n41897, n41898, n41899, n41900, n41901, n41902,
    n41903, n41904, n41905, n41906, n41907, n41908, n41909, n41910, n41911,
    n41912, n41913, n41914, n41915, n41916, n41917, n41918, n41919, n41920,
    n41921, n41922, n41923, n41924, n41925, n41926, n41927, n41928, n41929,
    n41930, n41931, n41932, n41933, n41934, n41936, n41937, n41938, n41939,
    n41940, n41941, n41942, n41943, n41944, n41945, n41946, n41947, n41948,
    n41949, n41950, n41951, n41952, n41953, n41954, n41955, n41956, n41957,
    n41958, n41959, n41960, n41961, n41962, n41963, n41964, n41965, n41966,
    n41967, n41968, n41969, n41970, n41971, n41972, n41973, n41974, n41975,
    n41976, n41977, n41978, n41979, n41980, n41981, n41983, n41984, n41985,
    n41986, n41987, n41988, n41989, n41990, n41991, n41992, n41993, n41994,
    n41995, n41996, n41997, n41998, n41999, n42000, n42001, n42002, n42003,
    n42004, n42005, n42006, n42007, n42008, n42009, n42010, n42011, n42012,
    n42013, n42014, n42015, n42016, n42017, n42019, n42020, n42021, n42022,
    n42023, n42024, n42025, n42026, n42027, n42028, n42029, n42030, n42031,
    n42032, n42033, n42034, n42035, n42036, n42037, n42038, n42039, n42040,
    n42041, n42042, n42043, n42044, n42045, n42046, n42047, n42048, n42049,
    n42050, n42051, n42052, n42053, n42054, n42055, n42057, n42058, n42059,
    n42060, n42061, n42062, n42063, n42064, n42065, n42066, n42067, n42068,
    n42069, n42070, n42071, n42072, n42073, n42074, n42075, n42076, n42077,
    n42078, n42079, n42080, n42081, n42082, n42083, n42084, n42085, n42087,
    n42088, n42089, n42090, n42091, n42092, n42093, n42094, n42095, n42096,
    n42097, n42098, n42099, n42100, n42101, n42102, n42103, n42104, n42105,
    n42106, n42107, n42108, n42109, n42110, n42111, n42112, n42113, n42114,
    n42115, n42116, n42118, n42119, n42120, n42121, n42122, n42123, n42124,
    n42125, n42126, n42127, n42128, n42129, n42130, n42131, n42132, n42133,
    n42134, n42135, n42136, n42137, n42138, n42139, n42140, n42141, n42142,
    n42143, n42144, n42146, n42147, n42148, n42149, n42150, n42151, n42152,
    n42153, n42154, n42155, n42156, n42157, n42158, n42159, n42160, n42161,
    n42162, n42163, n42164, n42165, n42166, n42167, n42168, n42169, n42170,
    n42171, n42172, n42173, n42174, n42175, n42176, n42177, n42178, n42179,
    n42180, n42182, n42183, n42184, n42185, n42186, n42187, n42188, n42189,
    n42190, n42191, n42192, n42193, n42194, n42195, n42196, n42197, n42198,
    n42199, n42200, n42201, n42202, n42203, n42204, n42205, n42206, n42207,
    n42208, n42209, n42210, n42211, n42212, n42213, n42214, n42215, n42216,
    n42217, n42218, n42219, n42220, n42221, n42222, n42223, n42224, n42225,
    n42226, n42227, n42228, n42229, n42230, n42231, n42232, n42233, n42234,
    n42235, n42236, n42237, n42238, n42239, n42240, n42241, n42242, n42243,
    n42244, n42245, n42246, n42247, n42248, n42249, n42250, n42251, n42252,
    n42253, n42254, n42255, n42256, n42257, n42258, n42259, n42260, n42261,
    n42262, n42263, n42264, n42265, n42266, n42267, n42268, n42269, n42270,
    n42271, n42272, n42273, n42274, n42275, n42276, n42277, n42278, n42279,
    n42280, n42281, n42282, n42283, n42285, n42286, n42287, n42288, n42289,
    n42290, n42291, n42292, n42293, n42294, n42295, n42296, n42297, n42298,
    n42299, n42300, n42301, n42302, n42303, n42304, n42305, n42306, n42307,
    n42308, n42309, n42310, n42311, n42312, n42313, n42314, n42315, n42316,
    n42317, n42318, n42319, n42320, n42321, n42322, n42323, n42324, n42325,
    n42326, n42327, n42328, n42329, n42330, n42331, n42332, n42333, n42334,
    n42335, n42336, n42337, n42338, n42339, n42340, n42341, n42342, n42343,
    n42344, n42345, n42346, n42347, n42348, n42349, n42350, n42351, n42352,
    n42353, n42354, n42355, n42356, n42357, n42358, n42359, n42360, n42361,
    n42362, n42363, n42364, n42365, n42366, n42367, n42368, n42369, n42370,
    n42371, n42372, n42373, n42374, n42376, n42377, n42378, n42379, n42380,
    n42381, n42382, n42383, n42384, n42385, n42386, n42387, n42388, n42389,
    n42390, n42391, n42392, n42393, n42394, n42395, n42396, n42397, n42398,
    n42399, n42400, n42401, n42402, n42403, n42404, n42405, n42406, n42407,
    n42408, n42409, n42410, n42411, n42412, n42413, n42414, n42415, n42416,
    n42417, n42418, n42419, n42420, n42421, n42422, n42423, n42424, n42425,
    n42426, n42427, n42428, n42429, n42430, n42431, n42432, n42433, n42434,
    n42435, n42436, n42437, n42438, n42439, n42440, n42441, n42442, n42443,
    n42444, n42445, n42446, n42447, n42448, n42449, n42450, n42451, n42452,
    n42453, n42454, n42455, n42456, n42457, n42458, n42459, n42460, n42461,
    n42462, n42463, n42464, n42465, n42466, n42467, n42468, n42469, n42470,
    n42471, n42472, n42473, n42474, n42475, n42476, n42477, n42478, n42479,
    n42480, n42481, n42482, n42484, n42485, n42486, n42487, n42488, n42489,
    n42490, n42491, n42492, n42493, n42494, n42495, n42496, n42497, n42498,
    n42499, n42500, n42501, n42502, n42503, n42504, n42505, n42506, n42507,
    n42508, n42509, n42510, n42511, n42512, n42513, n42514, n42515, n42516,
    n42517, n42518, n42519, n42520, n42521, n42522, n42523, n42524, n42525,
    n42526, n42527, n42528, n42529, n42530, n42531, n42532, n42533, n42534,
    n42535, n42536, n42537, n42538, n42539, n42540, n42541, n42542, n42543,
    n42544, n42545, n42546, n42547, n42548, n42549, n42550, n42551, n42552,
    n42553, n42554, n42555, n42556, n42557, n42558, n42559, n42560, n42561,
    n42562, n42563, n42564, n42565, n42566, n42567, n42568, n42569, n42570,
    n42571, n42572, n42573, n42574, n42575, n42576, n42577, n42578, n42579,
    n42580, n42581, n42582, n42583, n42585, n42586, n42587, n42588, n42589,
    n42590, n42591, n42592, n42593, n42594, n42595, n42596, n42597, n42598,
    n42599, n42600, n42601, n42602, n42603, n42604, n42605, n42606, n42607,
    n42608, n42609, n42610, n42611, n42612, n42613, n42614, n42615, n42616,
    n42617, n42618, n42619, n42620, n42621, n42622, n42623, n42625, n42626,
    n42627, n42628, n42629, n42630, n42631, n42632, n42633, n42634, n42635,
    n42636, n42637, n42638, n42639, n42640, n42641, n42642, n42643, n42644,
    n42645, n42646, n42647, n42648, n42649, n42650, n42651, n42652, n42653,
    n42654, n42655, n42656, n42657, n42658, n42659, n42660, n42662, n42663,
    n42664, n42665, n42666, n42667, n42668, n42669, n42670, n42671, n42672,
    n42673, n42674, n42675, n42676, n42677, n42678, n42679, n42680, n42681,
    n42682, n42683, n42684, n42685, n42686, n42687, n42688, n42689, n42690,
    n42691, n42692, n42693, n42694, n42695, n42696, n42697, n42698, n42699,
    n42700, n42701, n42702, n42703, n42704, n42705, n42706, n42707, n42708,
    n42709, n42710, n42711, n42712, n42713, n42714, n42715, n42716, n42717,
    n42718, n42719, n42720, n42721, n42722, n42723, n42724, n42725, n42726,
    n42727, n42728, n42729, n42730, n42731, n42732, n42733, n42734, n42735,
    n42736, n42737, n42738, n42739, n42740, n42741, n42742, n42743, n42744,
    n42745, n42746, n42747, n42748, n42749, n42750, n42751, n42752, n42753,
    n42754, n42755, n42756, n42757, n42758, n42759, n42761, n42762, n42763,
    n42764, n42765, n42766, n42767, n42768, n42769, n42770, n42771, n42772,
    n42773, n42774, n42775, n42776, n42777, n42778, n42779, n42780, n42781,
    n42782, n42783, n42784, n42785, n42786, n42787, n42788, n42789, n42790,
    n42791, n42792, n42793, n42794, n42795, n42796, n42797, n42798, n42799,
    n42800, n42801, n42802, n42803, n42804, n42805, n42806, n42807, n42808,
    n42809, n42810, n42811, n42812, n42813, n42814, n42815, n42816, n42817,
    n42818, n42819, n42820, n42821, n42822, n42823, n42824, n42825, n42826,
    n42827, n42828, n42829, n42830, n42831, n42832, n42833, n42834, n42835,
    n42836, n42837, n42838, n42839, n42840, n42841, n42842, n42843, n42844,
    n42845, n42846, n42847, n42848, n42849, n42850, n42851, n42852, n42853,
    n42854, n42855, n42856, n42857, n42858, n42859, n42860, n42861, n42862,
    n42864, n42865, n42866, n42867, n42868, n42869, n42870, n42871, n42872,
    n42873, n42874, n42875, n42876, n42877, n42878, n42879, n42880, n42881,
    n42882, n42883, n42884, n42885, n42886, n42887, n42888, n42889, n42890,
    n42891, n42892, n42893, n42894, n42895, n42896, n42897, n42898, n42899,
    n42900, n42901, n42902, n42903, n42904, n42905, n42906, n42907, n42908,
    n42909, n42910, n42911, n42912, n42913, n42914, n42916, n42917, n42918,
    n42919, n42920, n42921, n42922, n42923, n42924, n42925, n42926, n42927,
    n42928, n42929, n42930, n42931, n42932, n42933, n42934, n42935, n42936,
    n42937, n42938, n42939, n42940, n42941, n42942, n42943, n42944, n42945,
    n42946, n42947, n42948, n42949, n42950, n42951, n42952, n42953, n42954,
    n42955, n42956, n42957, n42959, n42960, n42961, n42962, n42963, n42964,
    n42965, n42966, n42967, n42968, n42969, n42970, n42971, n42972, n42973,
    n42974, n42975, n42976, n42977, n42978, n42979, n42980, n42981, n42982,
    n42983, n42984, n42985, n42986, n42987, n42988, n42989, n42990, n42991,
    n42992, n42993, n42994, n42995, n42996, n42997, n42998, n42999, n43000,
    n43001, n43002, n43003, n43004, n43006, n43007, n43008, n43009, n43010,
    n43011, n43012, n43013, n43014, n43015, n43016, n43017, n43018, n43019,
    n43020, n43021, n43022, n43023, n43024, n43025, n43026, n43027, n43028,
    n43029, n43030, n43031, n43032, n43033, n43034, n43035, n43036, n43037,
    n43038, n43039, n43040, n43041, n43043, n43044, n43045, n43046, n43047,
    n43048, n43049, n43050, n43051, n43052, n43053, n43054, n43055, n43056,
    n43057, n43058, n43059, n43060, n43061, n43062, n43063, n43064, n43065,
    n43066, n43067, n43068, n43069, n43070, n43071, n43072, n43073, n43074,
    n43075, n43076, n43077, n43078, n43079, n43080, n43081, n43082, n43083,
    n43084, n43085, n43086, n43087, n43088, n43089, n43090, n43091, n43092,
    n43093, n43094, n43096, n43097, n43098, n43099, n43100, n43101, n43102,
    n43103, n43104, n43105, n43106, n43107, n43108, n43109, n43110, n43111,
    n43112, n43113, n43114, n43115, n43116, n43117, n43118, n43119, n43120,
    n43121, n43122, n43123, n43124, n43125, n43126, n43127, n43128, n43129,
    n43131, n43132, n43133, n43134, n43135, n43136, n43137, n43138, n43139,
    n43140, n43141, n43142, n43143, n43144, n43145, n43146, n43147, n43148,
    n43149, n43150, n43151, n43152, n43153, n43154, n43155, n43156, n43157,
    n43158, n43159, n43160, n43161, n43162, n43163, n43164, n43165, n43167,
    n43168, n43169, n43170, n43171, n43172, n43173, n43174, n43175, n43176,
    n43177, n43178, n43179, n43180, n43181, n43182, n43183, n43184, n43185,
    n43186, n43187, n43188, n43189, n43190, n43191, n43192, n43193, n43194,
    n43195, n43196, n43197, n43198, n43199, n43200, n43201, n43202, n43203,
    n43204, n43205, n43207, n43208, n43209, n43210, n43211, n43212, n43213,
    n43214, n43215, n43216, n43217, n43218, n43219, n43220, n43221, n43222,
    n43223, n43224, n43225, n43226, n43227, n43228, n43229, n43230, n43231,
    n43232, n43233, n43234, n43235, n43236, n43237, n43238, n43239, n43240,
    n43241, n43242, n43243, n43244, n43245, n43246, n43247, n43248, n43249,
    n43250, n43251, n43252, n43253, n43254, n43255, n43256, n43257, n43258,
    n43259, n43260, n43261, n43262, n43263, n43264, n43265, n43266, n43267,
    n43268, n43269, n43270, n43271, n43272, n43273, n43274, n43275, n43276,
    n43277, n43278, n43279, n43280, n43281, n43282, n43283, n43284, n43285,
    n43286, n43287, n43288, n43289, n43290, n43291, n43292, n43293, n43294,
    n43295, n43296, n43297, n43298, n43300, n43301, n43302, n43303, n43304,
    n43305, n43306, n43307, n43308, n43309, n43310, n43311, n43312, n43313,
    n43314, n43315, n43316, n43317, n43318, n43319, n43320, n43321, n43322,
    n43323, n43324, n43325, n43326, n43327, n43328, n43329, n43330, n43331,
    n43332, n43333, n43334, n43335, n43336, n43337, n43338, n43339, n43340,
    n43341, n43342, n43343, n43344, n43345, n43346, n43347, n43348, n43349,
    n43350, n43351, n43352, n43353, n43354, n43355, n43356, n43357, n43358,
    n43359, n43360, n43361, n43362, n43363, n43364, n43365, n43366, n43367,
    n43368, n43369, n43370, n43371, n43372, n43373, n43374, n43375, n43376,
    n43377, n43378, n43379, n43380, n43381, n43382, n43383, n43384, n43385,
    n43386, n43387, n43388, n43389, n43390, n43391, n43392, n43393, n43394,
    n43395, n43396, n43397, n43398, n43399, n43400, n43401, n43402, n43403,
    n43405, n43406, n43407, n43408, n43409, n43410, n43411, n43412, n43413,
    n43414, n43415, n43416, n43417, n43418, n43419, n43420, n43421, n43422,
    n43423, n43424, n43425, n43426, n43427, n43428, n43429, n43430, n43431,
    n43432, n43433, n43434, n43435, n43436, n43437, n43438, n43439, n43440,
    n43441, n43442, n43444, n43445, n43446, n43447, n43448, n43449, n43450,
    n43451, n43452, n43453, n43454, n43455, n43456, n43457, n43458, n43459,
    n43460, n43461, n43462, n43463, n43464, n43465, n43466, n43467, n43468,
    n43469, n43470, n43471, n43472, n43473, n43474, n43475, n43476, n43477,
    n43478, n43479, n43480, n43481, n43482, n43483, n43484, n43485, n43486,
    n43487, n43488, n43489, n43491, n43492, n43493, n43494, n43495, n43496,
    n43497, n43498, n43499, n43500, n43501, n43502, n43503, n43504, n43505,
    n43506, n43507, n43508, n43509, n43510, n43511, n43512, n43513, n43514,
    n43515, n43516, n43517, n43518, n43519, n43520, n43521, n43522, n43523,
    n43524, n43525, n43527, n43528, n43529, n43530, n43531, n43532, n43533,
    n43534, n43535, n43536, n43537, n43538, n43539, n43540, n43541, n43542,
    n43543, n43544, n43545, n43546, n43547, n43548, n43549, n43550, n43551,
    n43552, n43553, n43554, n43555, n43556, n43557, n43558, n43559, n43560,
    n43561, n43562, n43563, n43565, n43566, n43567, n43568, n43569, n43570,
    n43571, n43572, n43573, n43574, n43575, n43576, n43577, n43578, n43579,
    n43580, n43581, n43582, n43583, n43584, n43585, n43586, n43587, n43588,
    n43589, n43590, n43591, n43592, n43593, n43594, n43596, n43597, n43598,
    n43599, n43600, n43601, n43602, n43603, n43604, n43605, n43606, n43607,
    n43608, n43609, n43610, n43611, n43612, n43613, n43614, n43615, n43616,
    n43617, n43618, n43619, n43620, n43621, n43622, n43624, n43625, n43626,
    n43627, n43628, n43629, n43630, n43631, n43632, n43633, n43634, n43635,
    n43636, n43637, n43638, n43639, n43640, n43641, n43642, n43643, n43644,
    n43645, n43646, n43647, n43648, n43649, n43650, n43651, n43652, n43653,
    n43654, n43656, n43657, n43658, n43659, n43660, n43661, n43662, n43663,
    n43664, n43665, n43666, n43667, n43668, n43669, n43670, n43671, n43672,
    n43673, n43674, n43675, n43676, n43677, n43678, n43679, n43680, n43681,
    n43682, n43683, n43684, n43685, n43686, n43687, n43688, n43689, n43690,
    n43692, n43693, n43694, n43695, n43696, n43697, n43698, n43699, n43700,
    n43701, n43702, n43703, n43704, n43705, n43706, n43707, n43708, n43709,
    n43710, n43711, n43712, n43713, n43714, n43715, n43716, n43717, n43718,
    n43719, n43720, n43721, n43722, n43723, n43724, n43725, n43726, n43727,
    n43728, n43729, n43730, n43731, n43732, n43733, n43734, n43735, n43736,
    n43737, n43739, n43740, n43741, n43742, n43743, n43744, n43745, n43746,
    n43747, n43748, n43749, n43750, n43751, n43752, n43753, n43754, n43755,
    n43756, n43757, n43758, n43759, n43760, n43761, n43762, n43763, n43764,
    n43765, n43766, n43767, n43769, n43770, n43771, n43772, n43773, n43774,
    n43775, n43776, n43777, n43778, n43779, n43780, n43781, n43782, n43783,
    n43784, n43785, n43786, n43787, n43788, n43789, n43790, n43791, n43792,
    n43793, n43794, n43795, n43796, n43797, n43798, n43799, n43800, n43801,
    n43802, n43803, n43804, n43806, n43807, n43808, n43809, n43810, n43811,
    n43812, n43813, n43814, n43815, n43816, n43817, n43818, n43819, n43820,
    n43821, n43822, n43823, n43824, n43825, n43826, n43827, n43828, n43829,
    n43830, n43831, n43832, n43833, n43834, n43835, n43836, n43837, n43838,
    n43839, n43840, n43842, n43843, n43844, n43845, n43846, n43847, n43848,
    n43849, n43850, n43851, n43852, n43853, n43854, n43855, n43856, n43857,
    n43858, n43859, n43860, n43861, n43862, n43863, n43864, n43865, n43866,
    n43867, n43868, n43869, n43870, n43871, n43872, n43873, n43874, n43875,
    n43876, n43877, n43878, n43879, n43880, n43882, n43883, n43884, n43885,
    n43886, n43887, n43888, n43889, n43890, n43891, n43892, n43893, n43894,
    n43895, n43896, n43897, n43898, n43899, n43900, n43901, n43902, n43903,
    n43904, n43905, n43906, n43907, n43908, n43909, n43910, n43911, n43912,
    n43913, n43914, n43915, n43916, n43918, n43919, n43920, n43921, n43922,
    n43923, n43924, n43925, n43926, n43927, n43928, n43929, n43930, n43931,
    n43932, n43933, n43934, n43935, n43936, n43937, n43938, n43939, n43940,
    n43941, n43942, n43943, n43944, n43945, n43946, n43947, n43948, n43949,
    n43950, n43951, n43952, n43953, n43954, n43955, n43956, n43957, n43958,
    n43959, n43960, n43961, n43962, n43963, n43964, n43965, n43966, n43967,
    n43968, n43969, n43970, n43971, n43972, n43973, n43974, n43975, n43976,
    n43977, n43978, n43979, n43980, n43981, n43982, n43983, n43984, n43985,
    n43986, n43987, n43988, n43989, n43990, n43991, n43992, n43993, n43994,
    n43995, n43996, n43997, n43998, n43999, n44000, n44001, n44002, n44003,
    n44004, n44005, n44006, n44007, n44008, n44009, n44010, n44011, n44012,
    n44013, n44014, n44015, n44016, n44017, n44018, n44020, n44021, n44022,
    n44023, n44024, n44025, n44026, n44027, n44028, n44029, n44030, n44031,
    n44032, n44033, n44034, n44035, n44036, n44037, n44038, n44039, n44040,
    n44041, n44042, n44043, n44044, n44045, n44046, n44047, n44048, n44049,
    n44050, n44051, n44052, n44053, n44054, n44055, n44056, n44057, n44058,
    n44059, n44060, n44061, n44062, n44063, n44064, n44065, n44066, n44067,
    n44068, n44069, n44070, n44071, n44072, n44073, n44074, n44075, n44076,
    n44077, n44078, n44079, n44080, n44081, n44082, n44083, n44084, n44085,
    n44086, n44087, n44088, n44089, n44090, n44091, n44092, n44093, n44094,
    n44095, n44096, n44097, n44098, n44099, n44100, n44101, n44102, n44103,
    n44104, n44105, n44106, n44107, n44108, n44109, n44110, n44111, n44112,
    n44113, n44114, n44115, n44116, n44117, n44118, n44119, n44120, n44121,
    n44122, n44123, n44125, n44126, n44127, n44128, n44129, n44130, n44131,
    n44132, n44133, n44134, n44135, n44136, n44137, n44138, n44139, n44140,
    n44141, n44142, n44143, n44144, n44145, n44146, n44147, n44148, n44149,
    n44150, n44151, n44152, n44153, n44154, n44155, n44156, n44157, n44158,
    n44159, n44160, n44161, n44162, n44163, n44164, n44165, n44166, n44167,
    n44168, n44169, n44170, n44171, n44172, n44173, n44174, n44175, n44176,
    n44177, n44178, n44179, n44180, n44181, n44182, n44183, n44184, n44185,
    n44186, n44187, n44188, n44189, n44190, n44191, n44192, n44193, n44194,
    n44195, n44196, n44197, n44198, n44199, n44200, n44201, n44202, n44203,
    n44204, n44205, n44206, n44207, n44208, n44209, n44210, n44211, n44212,
    n44213, n44214, n44215, n44216, n44217, n44218, n44219, n44220, n44221,
    n44222, n44223, n44224, n44225, n44226, n44227, n44228, n44229, n44230,
    n44232, n44233, n44234, n44235, n44236, n44237, n44238, n44239, n44240,
    n44241, n44242, n44243, n44244, n44245, n44246, n44247, n44248, n44249,
    n44250, n44251, n44252, n44253, n44254, n44255, n44256, n44257, n44258,
    n44259, n44260, n44261, n44262, n44263, n44264, n44265, n44266, n44267,
    n44268, n44269, n44270, n44271, n44272, n44273, n44274, n44275, n44276,
    n44277, n44278, n44279, n44280, n44281, n44282, n44283, n44284, n44285,
    n44286, n44287, n44288, n44289, n44290, n44291, n44292, n44293, n44294,
    n44295, n44296, n44297, n44298, n44299, n44300, n44301, n44302, n44303,
    n44304, n44305, n44306, n44307, n44308, n44309, n44310, n44311, n44312,
    n44313, n44314, n44315, n44316, n44317, n44318, n44319, n44320, n44321,
    n44322, n44323, n44324, n44325, n44326, n44327, n44328, n44329, n44330,
    n44331, n44332, n44333, n44334, n44335, n44336, n44338, n44339, n44340,
    n44341, n44342, n44343, n44344, n44345, n44346, n44347, n44348, n44349,
    n44350, n44351, n44352, n44353, n44354, n44355, n44356, n44357, n44358,
    n44359, n44360, n44361, n44362, n44363, n44364, n44365, n44366, n44367,
    n44368, n44369, n44370, n44371, n44372, n44373, n44374, n44375, n44376,
    n44377, n44378, n44379, n44380, n44381, n44382, n44384, n44385, n44386,
    n44387, n44388, n44389, n44390, n44391, n44392, n44393, n44394, n44395,
    n44396, n44397, n44398, n44399, n44400, n44401, n44402, n44403, n44404,
    n44405, n44406, n44407, n44408, n44409, n44410, n44411, n44412, n44413,
    n44414, n44415, n44416, n44417, n44419, n44420, n44421, n44422, n44423,
    n44424, n44425, n44426, n44427, n44428, n44429, n44430, n44431, n44432,
    n44433, n44434, n44435, n44436, n44437, n44438, n44439, n44440, n44441,
    n44442, n44443, n44444, n44445, n44446, n44447, n44448, n44449, n44450,
    n44451, n44452, n44453, n44454, n44455, n44456, n44457, n44459, n44460,
    n44461, n44462, n44463, n44464, n44465, n44466, n44467, n44468, n44469,
    n44470, n44471, n44472, n44473, n44474, n44475, n44476, n44477, n44478,
    n44479, n44480, n44481, n44482, n44483, n44484, n44485, n44486, n44487,
    n44488, n44489, n44490, n44491, n44492, n44493, n44494, n44495, n44496,
    n44497, n44499, n44500, n44501, n44502, n44503, n44504, n44505, n44506,
    n44507, n44508, n44509, n44510, n44511, n44512, n44513, n44514, n44515,
    n44516, n44517, n44518, n44519, n44520, n44521, n44522, n44523, n44524,
    n44525, n44526, n44527, n44528, n44530, n44531, n44532, n44533, n44534,
    n44535, n44536, n44537, n44538, n44539, n44540, n44541, n44542, n44543,
    n44544, n44545, n44546, n44547, n44548, n44549, n44550, n44551, n44552,
    n44553, n44554, n44555, n44556, n44557, n44558, n44559, n44560, n44561,
    n44563, n44564, n44565, n44566, n44567, n44568, n44569, n44570, n44571,
    n44572, n44573, n44574, n44575, n44576, n44577, n44578, n44579, n44580,
    n44581, n44582, n44583, n44584, n44585, n44586, n44587, n44588, n44589,
    n44590, n44591, n44592, n44593, n44594, n44595, n44596, n44597, n44598,
    n44599, n44600, n44601, n44602, n44603, n44605, n44606, n44607, n44608,
    n44609, n44610, n44611, n44612, n44613, n44614, n44615, n44616, n44617,
    n44618, n44619, n44620, n44621, n44622, n44623, n44624, n44625, n44626,
    n44627, n44628, n44629, n44630, n44631, n44632, n44633, n44634, n44635,
    n44636, n44637, n44638, n44639, n44640, n44641, n44642, n44643, n44644,
    n44645, n44646, n44647, n44648, n44649, n44650, n44651, n44652, n44653,
    n44654, n44655, n44656, n44657, n44658, n44659, n44660, n44661, n44662,
    n44663, n44664, n44665, n44666, n44667, n44668, n44669, n44670, n44671,
    n44672, n44673, n44674, n44675, n44676, n44677, n44678, n44679, n44680,
    n44681, n44682, n44683, n44684, n44685, n44686, n44687, n44688, n44689,
    n44690, n44691, n44692, n44693, n44694, n44696, n44697, n44698, n44699,
    n44700, n44701, n44702, n44703, n44704, n44705, n44706, n44707, n44708,
    n44709, n44710, n44711, n44712, n44713, n44714, n44715, n44716, n44717,
    n44718, n44719, n44720, n44721, n44722, n44723, n44724, n44725, n44726,
    n44727, n44728, n44729, n44730, n44731, n44732, n44733, n44734, n44735,
    n44736, n44738, n44739, n44740, n44741, n44742, n44743, n44744, n44745,
    n44746, n44747, n44748, n44749, n44750, n44751, n44752, n44753, n44754,
    n44755, n44756, n44757, n44758, n44759, n44760, n44761, n44762, n44763,
    n44764, n44765, n44766, n44767, n44768, n44769, n44770, n44771, n44772,
    n44773, n44774, n44775, n44776, n44777, n44778, n44779, n44780, n44781,
    n44782, n44783, n44784, n44785, n44786, n44787, n44788, n44789, n44790,
    n44791, n44792, n44793, n44794, n44795, n44796, n44797, n44798, n44799,
    n44800, n44801, n44802, n44803, n44804, n44805, n44806, n44807, n44808,
    n44809, n44810, n44811, n44812, n44813, n44814, n44815, n44816, n44817,
    n44818, n44819, n44820, n44821, n44822, n44823, n44824, n44825, n44826,
    n44827, n44829, n44830, n44831, n44832, n44833, n44834, n44835, n44836,
    n44837, n44838, n44839, n44840, n44841, n44842, n44843, n44844, n44845,
    n44846, n44847, n44848, n44849, n44850, n44851, n44852, n44853, n44854,
    n44855, n44856, n44857, n44858, n44859, n44860, n44861, n44862, n44863,
    n44864, n44865, n44866, n44867, n44868, n44869, n44870, n44871, n44872,
    n44873, n44875, n44876, n44877, n44878, n44879, n44880, n44881, n44882,
    n44883, n44884, n44885, n44886, n44887, n44888, n44889, n44890, n44891,
    n44892, n44893, n44894, n44895, n44896, n44897, n44898, n44899, n44900,
    n44901, n44902, n44903, n44904, n44905, n44906, n44907, n44908, n44909,
    n44910, n44911, n44912, n44913, n44914, n44915, n44916, n44918, n44919,
    n44920, n44921, n44922, n44923, n44924, n44925, n44926, n44927, n44928,
    n44929, n44930, n44931, n44932, n44933, n44934, n44935, n44936, n44937,
    n44938, n44939, n44940, n44941, n44942, n44943, n44944, n44945, n44946,
    n44947, n44948, n44949, n44950, n44951, n44952, n44953, n44954, n44956,
    n44957, n44958, n44959, n44960, n44961, n44962, n44963, n44964, n44965,
    n44966, n44967, n44968, n44969, n44970, n44971, n44972, n44973, n44974,
    n44975, n44976, n44977, n44978, n44979, n44980, n44981, n44982, n44983,
    n44984, n44985, n44986, n44987, n44988, n44989, n44990, n44991, n44992,
    n44993, n44994, n44995, n44996, n44997, n44998, n44999, n45000, n45001,
    n45002, n45003, n45004, n45005, n45006, n45008, n45009, n45010, n45011,
    n45012, n45013, n45014, n45015, n45016, n45017, n45018, n45019, n45020,
    n45021, n45022, n45023, n45024, n45025, n45026, n45027, n45028, n45029,
    n45030, n45031, n45032, n45033, n45034, n45035, n45036, n45037, n45038,
    n45039, n45040, n45041, n45042, n45043, n45045, n45046, n45047, n45048,
    n45049, n45050, n45051, n45052, n45053, n45054, n45055, n45056, n45057,
    n45058, n45059, n45060, n45061, n45062, n45063, n45064, n45065, n45066,
    n45067, n45068, n45069, n45070, n45071, n45072, n45073, n45074, n45075,
    n45076, n45077, n45078, n45079, n45080, n45081, n45082, n45083, n45085,
    n45086, n45087, n45088, n45089, n45090, n45091, n45092, n45093, n45094,
    n45095, n45096, n45097, n45098, n45099, n45100, n45101, n45102, n45103,
    n45104, n45105, n45106, n45107, n45108, n45109, n45110, n45111, n45112,
    n45113, n45114, n45115, n45116, n45117, n45118, n45119, n45120, n45121,
    n45122, n45123, n45124, n45125, n45126, n45127, n45128, n45129, n45130,
    n45131, n45132, n45133, n45134, n45135, n45136, n45137, n45138, n45139,
    n45140, n45141, n45142, n45143, n45144, n45145, n45146, n45147, n45148,
    n45149, n45150, n45151, n45152, n45153, n45154, n45155, n45156, n45157,
    n45158, n45159, n45160, n45161, n45162, n45163, n45164, n45165, n45166,
    n45167, n45168, n45169, n45170, n45171, n45172, n45173, n45174, n45175,
    n45176, n45177, n45178, n45179, n45181, n45182, n45183, n45184, n45185,
    n45186, n45187, n45188, n45189, n45190, n45191, n45192, n45193, n45194,
    n45195, n45196, n45197, n45198, n45199, n45200, n45201, n45202, n45203,
    n45204, n45205, n45206, n45207, n45208, n45209, n45210, n45211, n45212,
    n45213, n45214, n45215, n45217, n45218, n45219, n45220, n45221, n45222,
    n45223, n45224, n45225, n45226, n45227, n45228, n45229, n45230, n45231,
    n45232, n45233, n45234, n45235, n45236, n45237, n45238, n45239, n45240,
    n45241, n45242, n45243, n45244, n45245, n45246, n45247, n45248, n45249,
    n45250, n45251, n45252, n45253, n45254, n45255, n45256, n45257, n45258,
    n45259, n45260, n45261, n45262, n45263, n45264, n45266, n45267, n45268,
    n45269, n45270, n45271, n45272, n45273, n45274, n45275, n45276, n45277,
    n45278, n45279, n45280, n45281, n45282, n45283, n45284, n45285, n45286,
    n45287, n45288, n45289, n45290, n45291, n45292, n45293, n45294, n45295,
    n45296, n45297, n45298, n45299, n45300, n45301, n45302, n45303, n45304,
    n45305, n45306, n45307, n45309, n45310, n45311, n45312, n45313, n45314,
    n45315, n45316, n45317, n45318, n45319, n45320, n45321, n45322, n45323,
    n45324, n45325, n45326, n45327, n45328, n45329, n45330, n45331, n45332,
    n45333, n45334, n45335, n45336, n45337, n45338, n45339, n45340, n45341,
    n45342, n45343, n45344, n45345, n45346, n45348, n45349, n45350, n45351,
    n45352, n45353, n45354, n45355, n45356, n45357, n45358, n45359, n45360,
    n45361, n45362, n45363, n45364, n45365, n45366, n45367, n45368, n45369,
    n45370, n45371, n45372, n45373, n45374, n45375, n45376, n45377, n45378,
    n45379, n45380, n45381, n45382, n45384, n45385, n45386, n45387, n45388,
    n45389, n45390, n45391, n45392, n45393, n45394, n45395, n45396, n45397,
    n45398, n45399, n45400, n45401, n45402, n45403, n45404, n45405, n45406,
    n45407, n45408, n45409, n45410, n45411, n45412, n45413, n45414, n45415,
    n45416, n45417, n45418, n45419, n45420, n45421, n45422, n45423, n45424,
    n45425, n45426, n45427, n45428, n45429, n45430, n45431, n45432, n45433,
    n45434, n45435, n45436, n45437, n45438, n45439, n45440, n45441, n45442,
    n45443, n45444, n45445, n45446, n45447, n45448, n45449, n45450, n45451,
    n45452, n45453, n45454, n45455, n45456, n45457, n45458, n45459, n45460,
    n45461, n45462, n45463, n45464, n45465, n45466, n45467, n45468, n45469,
    n45470, n45471, n45472, n45473, n45474, n45475, n45476, n45477, n45478,
    n45480, n45481, n45482, n45483, n45484, n45485, n45486, n45487, n45488,
    n45489, n45490, n45491, n45492, n45493, n45494, n45495, n45496, n45497,
    n45498, n45499, n45500, n45501, n45502, n45503, n45504, n45505, n45506,
    n45507, n45508, n45510, n45511, n45512, n45513, n45514, n45515, n45516,
    n45517, n45518, n45519, n45520, n45521, n45522, n45523, n45524, n45525,
    n45526, n45527, n45528, n45529, n45530, n45531, n45532, n45533, n45534,
    n45535, n45536, n45537, n45538, n45539, n45540, n45541, n45542, n45543,
    n45544, n45545, n45546, n45547, n45549, n45550, n45551, n45552, n45553,
    n45554, n45555, n45556, n45557, n45558, n45559, n45560, n45561, n45562,
    n45563, n45564, n45565, n45566, n45567, n45568, n45569, n45570, n45571,
    n45572, n45573, n45574, n45575, n45576, n45577, n45578, n45579, n45580,
    n45581, n45582, n45583, n45584, n45585, n45586, n45587, n45588, n45589,
    n45590, n45592, n45593, n45594, n45595, n45596, n45597, n45598, n45599,
    n45600, n45601, n45602, n45603, n45604, n45605, n45606, n45607, n45608,
    n45609, n45610, n45611, n45612, n45613, n45614, n45615, n45616, n45617,
    n45618, n45619, n45620, n45621, n45622, n45623, n45624, n45625, n45626,
    n45628, n45629, n45630, n45631, n45632, n45633, n45634, n45635, n45636,
    n45637, n45638, n45639, n45640, n45641, n45642, n45643, n45644, n45645,
    n45646, n45647, n45648, n45649, n45650, n45651, n45652, n45653, n45654,
    n45656, n45657, n45658, n45659, n45660, n45661, n45662, n45663, n45664,
    n45665, n45666, n45667, n45668, n45669, n45670, n45671, n45672, n45673,
    n45674, n45675, n45676, n45677, n45678, n45679, n45680, n45681, n45682,
    n45683, n45684, n45685, n45686, n45687, n45688, n45689, n45690, n45691,
    n45692, n45693, n45694, n45695, n45696, n45697, n45698, n45699, n45700,
    n45701, n45702, n45703, n45704, n45705, n45706, n45707, n45708, n45709,
    n45710, n45711, n45712, n45713, n45714, n45715, n45716, n45717, n45718,
    n45719, n45720, n45721, n45722, n45723, n45724, n45725, n45726, n45727,
    n45728, n45729, n45730, n45731, n45732, n45733, n45734, n45735, n45736,
    n45737, n45738, n45739, n45740, n45741, n45742, n45743, n45744, n45745,
    n45746, n45747, n45748, n45749, n45750, n45751, n45752, n45753, n45754,
    n45755, n45756, n45757, n45758, n45760, n45761, n45762, n45763, n45764,
    n45765, n45766, n45767, n45768, n45769, n45770, n45771, n45772, n45773,
    n45774, n45775, n45776, n45777, n45778, n45779, n45780, n45781, n45782,
    n45783, n45784, n45785, n45786, n45787, n45788, n45789, n45790, n45791,
    n45792, n45793, n45794, n45795, n45796, n45797, n45798, n45799, n45800,
    n45801, n45802, n45803, n45804, n45805, n45806, n45807, n45808, n45809,
    n45810, n45811, n45812, n45813, n45814, n45815, n45816, n45817, n45818,
    n45819, n45820, n45821, n45822, n45823, n45824, n45825, n45826, n45827,
    n45828, n45829, n45830, n45831, n45832, n45833, n45834, n45835, n45836,
    n45837, n45838, n45839, n45840, n45841, n45842, n45843, n45844, n45845,
    n45846, n45847, n45848, n45849, n45850, n45851, n45852, n45853, n45854,
    n45855, n45856, n45857, n45858, n45860, n45861, n45862, n45863, n45864,
    n45865, n45866, n45867, n45868, n45869, n45870, n45871, n45872, n45873,
    n45874, n45875, n45876, n45877, n45878, n45879, n45880, n45881, n45882,
    n45883, n45884, n45885, n45886, n45887, n45888, n45889, n45890, n45891,
    n45892, n45893, n45894, n45895, n45896, n45897, n45898, n45899, n45900,
    n45901, n45902, n45903, n45904, n45905, n45906, n45907, n45908, n45909,
    n45910, n45911, n45912, n45913, n45914, n45915, n45916, n45917, n45918,
    n45919, n45920, n45921, n45922, n45923, n45924, n45925, n45926, n45927,
    n45928, n45929, n45930, n45931, n45932, n45933, n45934, n45935, n45936,
    n45937, n45938, n45939, n45940, n45941, n45942, n45943, n45944, n45945,
    n45946, n45947, n45948, n45949, n45950, n45951, n45952, n45953, n45955,
    n45956, n45957, n45958, n45959, n45960, n45961, n45962, n45963, n45964,
    n45965, n45966, n45967, n45968, n45969, n45970, n45971, n45972, n45973,
    n45974, n45975, n45976, n45977, n45978, n45979, n45980, n45981, n45982,
    n45983, n45984, n45985, n45986, n45987, n45988, n45989, n45991, n45992,
    n45993, n45994, n45995, n45996, n45997, n45998, n45999, n46000, n46001,
    n46002, n46003, n46004, n46005, n46006, n46007, n46008, n46009, n46010,
    n46011, n46012, n46013, n46014, n46015, n46016, n46017, n46018, n46019,
    n46020, n46021, n46022, n46023, n46024, n46026, n46027, n46028, n46029,
    n46030, n46031, n46032, n46033, n46034, n46035, n46036, n46037, n46038,
    n46039, n46040, n46041, n46042, n46043, n46044, n46045, n46046, n46047,
    n46048, n46049, n46051, n46052, n46053, n46054, n46055, n46056, n46057,
    n46058, n46059, n46060, n46061, n46062, n46063, n46064, n46065, n46066,
    n46067, n46068, n46069, n46070, n46071, n46072, n46073, n46074, n46075,
    n46076, n46077, n46078, n46079, n46080, n46081, n46082, n46083, n46084,
    n46085, n46086, n46087, n46088, n46089, n46090, n46091, n46092, n46093,
    n46094, n46095, n46096, n46097, n46098, n46099, n46100, n46101, n46102,
    n46103, n46104, n46105, n46106, n46107, n46108, n46109, n46110, n46111,
    n46112, n46113, n46114, n46115, n46116, n46117, n46118, n46119, n46120,
    n46121, n46122, n46123, n46124, n46125, n46126, n46127, n46128, n46129,
    n46130, n46131, n46132, n46133, n46134, n46135, n46136, n46137, n46138,
    n46139, n46140, n46141, n46142, n46143, n46144, n46145, n46146, n46147,
    n46148, n46149, n46150, n46151, n46152, n46153, n46155, n46156, n46157,
    n46158, n46159, n46160, n46161, n46162, n46163, n46164, n46165, n46166,
    n46167, n46168, n46169, n46170, n46171, n46172, n46173, n46174, n46175,
    n46176, n46177, n46178, n46179, n46180, n46181, n46182, n46183, n46184,
    n46185, n46186, n46187, n46188, n46189, n46190, n46191, n46192, n46193,
    n46195, n46196, n46197, n46198, n46199, n46200, n46201, n46202, n46203,
    n46204, n46205, n46206, n46207, n46208, n46209, n46210, n46211, n46212,
    n46213, n46214, n46215, n46216, n46217, n46218, n46219, n46220, n46221,
    n46222, n46223, n46224, n46225, n46227, n46228, n46229, n46230, n46231,
    n46232, n46233, n46234, n46235, n46236, n46237, n46238, n46239, n46240,
    n46241, n46242, n46243, n46244, n46245, n46246, n46247, n46248, n46249,
    n46250, n46251, n46252, n46253, n46254, n46255, n46256, n46257, n46258,
    n46259, n46260, n46261, n46262, n46263, n46264, n46265, n46266, n46267,
    n46268, n46269, n46270, n46271, n46272, n46273, n46274, n46275, n46276,
    n46277, n46278, n46279, n46280, n46281, n46282, n46283, n46284, n46285,
    n46286, n46287, n46288, n46289, n46290, n46291, n46292, n46293, n46294,
    n46295, n46296, n46297, n46298, n46299, n46300, n46301, n46302, n46303,
    n46304, n46305, n46306, n46307, n46308, n46309, n46310, n46311, n46312,
    n46313, n46314, n46315, n46316, n46317, n46318, n46319, n46320, n46321,
    n46322, n46324, n46325, n46326, n46327, n46328, n46329, n46330, n46331,
    n46332, n46333, n46334, n46335, n46336, n46337, n46338, n46339, n46340,
    n46341, n46342, n46343, n46344, n46345, n46346, n46347, n46348, n46349,
    n46351, n46352, n46353, n46354, n46355, n46356, n46357, n46358, n46359,
    n46360, n46361, n46362, n46363, n46364, n46365, n46366, n46367, n46368,
    n46369, n46370, n46371, n46372, n46373, n46374, n46375, n46376, n46377,
    n46378, n46379, n46380, n46381, n46382, n46383, n46384, n46385, n46386,
    n46387, n46388, n46389, n46390, n46391, n46392, n46393, n46394, n46395,
    n46396, n46397, n46398, n46399, n46400, n46401, n46402, n46403, n46404,
    n46405, n46406, n46407, n46408, n46409, n46410, n46411, n46412, n46413,
    n46414, n46415, n46416, n46417, n46418, n46419, n46420, n46421, n46422,
    n46423, n46424, n46425, n46426, n46427, n46428, n46429, n46430, n46431,
    n46432, n46433, n46434, n46435, n46437, n46438, n46439, n46440, n46441,
    n46442, n46443, n46444, n46445, n46446, n46447, n46448, n46449, n46450,
    n46451, n46452, n46453, n46454, n46455, n46456, n46457, n46458, n46459,
    n46460, n46461, n46462, n46463, n46464, n46465, n46466, n46467, n46468,
    n46469, n46470, n46471, n46473, n46474, n46475, n46476, n46477, n46478,
    n46479, n46480, n46481, n46482, n46483, n46484, n46485, n46486, n46487,
    n46488, n46489, n46490, n46491, n46492, n46493, n46494, n46495, n46496,
    n46497, n46498, n46499, n46501, n46502, n46503, n46504, n46505, n46506,
    n46507, n46508, n46509, n46510, n46511, n46512, n46513, n46514, n46515,
    n46516, n46517, n46518, n46519, n46520, n46521, n46522, n46523, n46524,
    n46525, n46526, n46527, n46528, n46529, n46530, n46531, n46532, n46533,
    n46534, n46535, n46536, n46537, n46538, n46539, n46540, n46541, n46542,
    n46543, n46544, n46546, n46547, n46548, n46549, n46550, n46551, n46552,
    n46553, n46554, n46555, n46556, n46557, n46558, n46559, n46560, n46561,
    n46562, n46563, n46564, n46565, n46566, n46567, n46568, n46569, n46570,
    n46571, n46572, n46573, n46574, n46575, n46576, n46577, n46578, n46579,
    n46580, n46582, n46583, n46584, n46585, n46586, n46587, n46588, n46589,
    n46590, n46591, n46592, n46593, n46594, n46595, n46596, n46597, n46598,
    n46599, n46600, n46601, n46602, n46603, n46604, n46605, n46606, n46607,
    n46608, n46609, n46610, n46611, n46612, n46614, n46615, n46616, n46617,
    n46618, n46619, n46620, n46621, n46622, n46623, n46624, n46625, n46626,
    n46627, n46628, n46629, n46630, n46631, n46632, n46633, n46634, n46635,
    n46636, n46637, n46638, n46639, n46640, n46641, n46642, n46644, n46645,
    n46646, n46647, n46648, n46649, n46650, n46651, n46652, n46653, n46654,
    n46655, n46656, n46657, n46658, n46659, n46660, n46661, n46662, n46663,
    n46664, n46665, n46666, n46667, n46668, n46669, n46670, n46671, n46672,
    n46673, n46674, n46675, n46676, n46677, n46678, n46679, n46680, n46681,
    n46682, n46683, n46684, n46685, n46686, n46687, n46688, n46689, n46690,
    n46691, n46692, n46693, n46694, n46695, n46696, n46697, n46698, n46699,
    n46700, n46701, n46702, n46703, n46704, n46705, n46706, n46707, n46708,
    n46709, n46710, n46711, n46712, n46713, n46714, n46715, n46716, n46717,
    n46718, n46719, n46720, n46721, n46722, n46723, n46724, n46725, n46726,
    n46727, n46728, n46729, n46730, n46731, n46732, n46733, n46734, n46735,
    n46737, n46738, n46739, n46740, n46741, n46742, n46743, n46744, n46745,
    n46746, n46747, n46748, n46749, n46750, n46751, n46752, n46753, n46754,
    n46755, n46756, n46757, n46758, n46759, n46760, n46761, n46762, n46763,
    n46764, n46765, n46766, n46767, n46768, n46769, n46770, n46771, n46772,
    n46773, n46775, n46776, n46777, n46778, n46779, n46780, n46781, n46782,
    n46783, n46784, n46785, n46786, n46787, n46788, n46789, n46790, n46791,
    n46792, n46793, n46794, n46795, n46796, n46797, n46798, n46799, n46800,
    n46801, n46802, n46803, n46804, n46805, n46806, n46807, n46808, n46809,
    n46811, n46812, n46813, n46814, n46815, n46816, n46817, n46818, n46819,
    n46820, n46821, n46822, n46823, n46824, n46825, n46826, n46827, n46828,
    n46829, n46830, n46831, n46832, n46833, n46834, n46835, n46836, n46837,
    n46838, n46839, n46840, n46842, n46843, n46844, n46845, n46846, n46847,
    n46848, n46849, n46850, n46851, n46852, n46853, n46854, n46855, n46856,
    n46857, n46858, n46859, n46860, n46861, n46862, n46863, n46864, n46865,
    n46866, n46867, n46868, n46869, n46870, n46871, n46872, n46873, n46874,
    n46875, n46876, n46877, n46878, n46879, n46880, n46881, n46882, n46883,
    n46884, n46885, n46886, n46887, n46889, n46890, n46891, n46892, n46893,
    n46894, n46895, n46896, n46897, n46898, n46899, n46900, n46901, n46902,
    n46903, n46904, n46905, n46906, n46907, n46908, n46909, n46910, n46911,
    n46912, n46913, n46914, n46915, n46916, n46917, n46918, n46919, n46920,
    n46921, n46922, n46923, n46924, n46925, n46926, n46927, n46928, n46929,
    n46930, n46931, n46932, n46933, n46934, n46935, n46936, n46937, n46938,
    n46939, n46940, n46941, n46942, n46943, n46944, n46945, n46946, n46947,
    n46948, n46949, n46950, n46951, n46952, n46953, n46954, n46955, n46956,
    n46957, n46958, n46959, n46960, n46961, n46962, n46963, n46964, n46965,
    n46966, n46967, n46968, n46969, n46970, n46971, n46972, n46973, n46974,
    n46975, n46976, n46977, n46978, n46979, n46980, n46982, n46983, n46984,
    n46985, n46986, n46987, n46988, n46989, n46990, n46991, n46992, n46993,
    n46994, n46995, n46996, n46997, n46998, n46999, n47000, n47001, n47002,
    n47003, n47004, n47005, n47006, n47007, n47008, n47009, n47011, n47012,
    n47013, n47014, n47015, n47016, n47017, n47018, n47019, n47020, n47021,
    n47022, n47023, n47024, n47025, n47026, n47027, n47028, n47029, n47030,
    n47031, n47032, n47033, n47034, n47035, n47036, n47037, n47038, n47039,
    n47040, n47041, n47042, n47043, n47044, n47045, n47046, n47048, n47049,
    n47050, n47051, n47052, n47053, n47054, n47055, n47056, n47057, n47058,
    n47059, n47060, n47061, n47062, n47063, n47064, n47065, n47066, n47067,
    n47068, n47069, n47070, n47071, n47072, n47073, n47074, n47075, n47076,
    n47077, n47078, n47079, n47080, n47081, n47082, n47083, n47084, n47085,
    n47086, n47087, n47089, n47090, n47091, n47092, n47093, n47094, n47095,
    n47096, n47097, n47098, n47099, n47100, n47101, n47102, n47103, n47104,
    n47105, n47106, n47107, n47108, n47109, n47110, n47111, n47112, n47113,
    n47114, n47115, n47116, n47117, n47118, n47120, n47121, n47122, n47123,
    n47124, n47125, n47126, n47127, n47128, n47129, n47130, n47131, n47132,
    n47133, n47134, n47135, n47136, n47137, n47138, n47139, n47140, n47141,
    n47142, n47143, n47144, n47145, n47147, n47148, n47149, n47150, n47151,
    n47152, n47153, n47154, n47155, n47156, n47157, n47158, n47159, n47160,
    n47161, n47162, n47163, n47164, n47165, n47166, n47167, n47168, n47169,
    n47170, n47171, n47173, n47174, n47175, n47176, n47177, n47178, n47179,
    n47180, n47181, n47182, n47183, n47184, n47185, n47186, n47187, n47188,
    n47189, n47190, n47191, n47192, n47193, n47194, n47195, n47196, n47197,
    n47198, n47199, n47200, n47201, n47202, n47203, n47205, n47206, n47207,
    n47208, n47209, n47210, n47211, n47212, n47213, n47214, n47215, n47216,
    n47217, n47218, n47219, n47220, n47221, n47222, n47223, n47224, n47225,
    n47226, n47227, n47228, n47230, n47231, n47232, n47233, n47234, n47235,
    n47236, n47237, n47238, n47239, n47240, n47241, n47242, n47243, n47244,
    n47245, n47246, n47247, n47248, n47249, n47250, n47251, n47252, n47253,
    n47254, n47255, n47256, n47257, n47258, n47259, n47260, n47261, n47262,
    n47263, n47264, n47265, n47266, n47267, n47268, n47269, n47270, n47271,
    n47272, n47273, n47274, n47275, n47276, n47277, n47278, n47279, n47280,
    n47281, n47282, n47283, n47284, n47285, n47286, n47287, n47288, n47289,
    n47290, n47291, n47292, n47293, n47294, n47295, n47296, n47297, n47298,
    n47299, n47300, n47301, n47302, n47303, n47304, n47305, n47306, n47307,
    n47308, n47309, n47310, n47311, n47312, n47313, n47314, n47315, n47316,
    n47317, n47318, n47319, n47320, n47321, n47322, n47323, n47324, n47325,
    n47326, n47327, n47328, n47329, n47330, n47332, n47333, n47334, n47335,
    n47336, n47337, n47338, n47339, n47340, n47341, n47342, n47343, n47344,
    n47345, n47346, n47347, n47348, n47349, n47350, n47351, n47352, n47353,
    n47354, n47355, n47356, n47357, n47358, n47359, n47360, n47361, n47362,
    n47363, n47364, n47365, n47366, n47367, n47368, n47369, n47370, n47371,
    n47372, n47373, n47374, n47375, n47376, n47377, n47378, n47379, n47380,
    n47381, n47382, n47383, n47384, n47385, n47386, n47387, n47388, n47389,
    n47390, n47391, n47392, n47393, n47394, n47395, n47396, n47397, n47398,
    n47399, n47400, n47401, n47402, n47403, n47404, n47405, n47406, n47407,
    n47408, n47409, n47410, n47411, n47412, n47413, n47414, n47415, n47416,
    n47417, n47418, n47419, n47420, n47421, n47422, n47423, n47424, n47425,
    n47426, n47427, n47428, n47429, n47430, n47431, n47432, n47433, n47435,
    n47436, n47437, n47438, n47439, n47440, n47441, n47442, n47443, n47444,
    n47445, n47446, n47447, n47448, n47449, n47450, n47451, n47452, n47453,
    n47454, n47455, n47456, n47457, n47458, n47459, n47460, n47461, n47462,
    n47463, n47464, n47465, n47466, n47467, n47468, n47469, n47470, n47471,
    n47472, n47473, n47474, n47475, n47476, n47477, n47478, n47479, n47481,
    n47482, n47483, n47484, n47485, n47486, n47487, n47488, n47489, n47490,
    n47491, n47492, n47493, n47494, n47495, n47496, n47497, n47498, n47499,
    n47500, n47501, n47502, n47503, n47504, n47505, n47506, n47507, n47508,
    n47509, n47510, n47511, n47512, n47513, n47514, n47515, n47516, n47517,
    n47518, n47519, n47521, n47522, n47523, n47524, n47525, n47526, n47527,
    n47528, n47529, n47530, n47531, n47532, n47533, n47534, n47535, n47536,
    n47537, n47538, n47539, n47540, n47541, n47542, n47543, n47544, n47545,
    n47546, n47547, n47548, n47549, n47550, n47551, n47552, n47553, n47554,
    n47555, n47556, n47557, n47558, n47559, n47560, n47561, n47562, n47563,
    n47564, n47565, n47566, n47567, n47568, n47569, n47570, n47571, n47572,
    n47573, n47574, n47575, n47576, n47577, n47578, n47579, n47580, n47581,
    n47582, n47583, n47584, n47585, n47586, n47587, n47588, n47589, n47590,
    n47591, n47592, n47593, n47594, n47595, n47596, n47597, n47598, n47599,
    n47600, n47601, n47602, n47603, n47604, n47605, n47606, n47607, n47608,
    n47609, n47610, n47611, n47612, n47613, n47614, n47615, n47616, n47617,
    n47618, n47620, n47621, n47622, n47623, n47624, n47625, n47626, n47627,
    n47628, n47629, n47630, n47631, n47632, n47633, n47634, n47635, n47636,
    n47637, n47638, n47639, n47640, n47641, n47642, n47643, n47644, n47645,
    n47646, n47647, n47648, n47649, n47650, n47651, n47652, n47653, n47654,
    n47655, n47656, n47657, n47658, n47659, n47660, n47661, n47662, n47663,
    n47664, n47665, n47666, n47667, n47668, n47669, n47670, n47671, n47672,
    n47673, n47674, n47675, n47676, n47677, n47678, n47679, n47680, n47681,
    n47682, n47683, n47684, n47685, n47686, n47687, n47688, n47689, n47690,
    n47691, n47692, n47693, n47694, n47695, n47696, n47697, n47698, n47699,
    n47700, n47701, n47702, n47703, n47704, n47705, n47706, n47707, n47708,
    n47709, n47710, n47711, n47712, n47713, n47714, n47715, n47716, n47717,
    n47718, n47719, n47720, n47721, n47722, n47723, n47724, n47726, n47727,
    n47728, n47729, n47730, n47731, n47732, n47733, n47734, n47735, n47736,
    n47737, n47738, n47739, n47740, n47741, n47742, n47743, n47744, n47745,
    n47746, n47747, n47748, n47749, n47750, n47751, n47752, n47753, n47754,
    n47755, n47756, n47757, n47758, n47759, n47760, n47761, n47762, n47763,
    n47764, n47765, n47766, n47767, n47768, n47769, n47770, n47771, n47772,
    n47773, n47774, n47775, n47776, n47777, n47778, n47779, n47780, n47781,
    n47782, n47783, n47784, n47785, n47786, n47787, n47788, n47789, n47790,
    n47791, n47792, n47793, n47794, n47795, n47796, n47797, n47798, n47799,
    n47800, n47801, n47802, n47803, n47804, n47805, n47806, n47807, n47808,
    n47809, n47810, n47811, n47812, n47813, n47814, n47815, n47816, n47817,
    n47818, n47819, n47820, n47821, n47822, n47823, n47824, n47825, n47826,
    n47827, n47829, n47830, n47831, n47832, n47833, n47834, n47835, n47836,
    n47837, n47838, n47839, n47840, n47841, n47842, n47843, n47844, n47845,
    n47846, n47847, n47848, n47849, n47850, n47851, n47852, n47853, n47854,
    n47855, n47856, n47857, n47858, n47859, n47860, n47861, n47862, n47863,
    n47864, n47865, n47866, n47867, n47868, n47869, n47870, n47871, n47872,
    n47873, n47874, n47875, n47876, n47877, n47878, n47879, n47880, n47881,
    n47882, n47883, n47884, n47885, n47886, n47887, n47888, n47889, n47890,
    n47891, n47892, n47893, n47894, n47895, n47896, n47897, n47898, n47899,
    n47900, n47901, n47902, n47903, n47904, n47905, n47906, n47907, n47908,
    n47909, n47910, n47911, n47912, n47913, n47914, n47915, n47916, n47917,
    n47918, n47919, n47920, n47921, n47922, n47923, n47924, n47925, n47926,
    n47927, n47929, n47930, n47931, n47932, n47933, n47934, n47935, n47936,
    n47937, n47938, n47939, n47940, n47941, n47942, n47943, n47944, n47945,
    n47946, n47947, n47948, n47949, n47950, n47951, n47952, n47953, n47954,
    n47956, n47957, n47958, n47959, n47960, n47961, n47962, n47963, n47964,
    n47965, n47966, n47967, n47968, n47969, n47970, n47971, n47972, n47973,
    n47974, n47975, n47976, n47977, n47978, n47979, n47980, n47981, n47982,
    n47983, n47984, n47985, n47986, n47987, n47988, n47989, n47990, n47991,
    n47992, n47993, n47994, n47995, n47996, n47998, n47999, n48000, n48001,
    n48002, n48003, n48004, n48005, n48006, n48007, n48008, n48009, n48010,
    n48011, n48012, n48013, n48014, n48015, n48016, n48017, n48018, n48019,
    n48020, n48021, n48022, n48023, n48024, n48025, n48026, n48027, n48028,
    n48029, n48031, n48032, n48033, n48034, n48035, n48036, n48037, n48038,
    n48039, n48040, n48041, n48042, n48043, n48044, n48045, n48046, n48047,
    n48048, n48049, n48050, n48051, n48052, n48053, n48054, n48055, n48056,
    n48057, n48058, n48059, n48060, n48061, n48062, n48063, n48064, n48065,
    n48066, n48067, n48068, n48069, n48070, n48071, n48072, n48073, n48074,
    n48075, n48076, n48077, n48078, n48080, n48081, n48082, n48083, n48084,
    n48085, n48086, n48087, n48088, n48089, n48090, n48091, n48092, n48093,
    n48094, n48095, n48096, n48097, n48098, n48099, n48100, n48101, n48102,
    n48103, n48104, n48105, n48106, n48107, n48108, n48109, n48110, n48111,
    n48112, n48113, n48114, n48115, n48116, n48117, n48118, n48119, n48120,
    n48121, n48122, n48123, n48124, n48125, n48126, n48127, n48128, n48129,
    n48130, n48131, n48132, n48133, n48134, n48135, n48136, n48137, n48138,
    n48139, n48140, n48141, n48142, n48143, n48144, n48145, n48146, n48147,
    n48148, n48149, n48150, n48151, n48152, n48153, n48154, n48155, n48156,
    n48157, n48158, n48159, n48160, n48161, n48162, n48163, n48164, n48165,
    n48166, n48167, n48168, n48169, n48171, n48172, n48173, n48174, n48175,
    n48176, n48177, n48178, n48179, n48180, n48181, n48182, n48183, n48184,
    n48185, n48186, n48187, n48188, n48189, n48190, n48191, n48192, n48193,
    n48194, n48195, n48196, n48197, n48198, n48199, n48200, n48201, n48202,
    n48203, n48204, n48205, n48206, n48207, n48209, n48210, n48211, n48212,
    n48213, n48214, n48215, n48216, n48217, n48218, n48219, n48220, n48221,
    n48222, n48223, n48224, n48225, n48226, n48227, n48228, n48229, n48230,
    n48231, n48232, n48233, n48234, n48235, n48236, n48237, n48238, n48239,
    n48240, n48241, n48242, n48243, n48244, n48245, n48246, n48247, n48248,
    n48249, n48250, n48251, n48252, n48253, n48254, n48255, n48256, n48257,
    n48258, n48259, n48260, n48261, n48262, n48263, n48264, n48265, n48266,
    n48267, n48268, n48269, n48270, n48271, n48272, n48273, n48274, n48275,
    n48276, n48277, n48278, n48279, n48280, n48281, n48282, n48283, n48284,
    n48285, n48286, n48287, n48288, n48289, n48290, n48291, n48292, n48293,
    n48294, n48295, n48296, n48297, n48298, n48299, n48300, n48301, n48302,
    n48303, n48304, n48305, n48307, n48308, n48309, n48310, n48311, n48312,
    n48313, n48314, n48315, n48316, n48317, n48318, n48319, n48320, n48321,
    n48322, n48323, n48324, n48325, n48326, n48327, n48328, n48329, n48330,
    n48331, n48332, n48333, n48334, n48335, n48336, n48337, n48338, n48339,
    n48340, n48341, n48342, n48343, n48345, n48346, n48347, n48348, n48349,
    n48350, n48351, n48352, n48353, n48354, n48355, n48356, n48357, n48358,
    n48359, n48360, n48361, n48362, n48363, n48364, n48365, n48366, n48367,
    n48368, n48369, n48370, n48371, n48372, n48373, n48374, n48375, n48376,
    n48377, n48378, n48379, n48380, n48381, n48382, n48383, n48384, n48385,
    n48386, n48387, n48388, n48390, n48391, n48392, n48393, n48394, n48395,
    n48396, n48397, n48398, n48399, n48400, n48401, n48402, n48403, n48404,
    n48405, n48406, n48407, n48408, n48409, n48410, n48411, n48412, n48413,
    n48414, n48415, n48416, n48417, n48418, n48419, n48420, n48421, n48422,
    n48423, n48424, n48425, n48426, n48427, n48428, n48429, n48430, n48431,
    n48432, n48433, n48434, n48435, n48436, n48437, n48438, n48439, n48440,
    n48442, n48443, n48444, n48445, n48446, n48447, n48448, n48449, n48450,
    n48451, n48452, n48453, n48454, n48455, n48456, n48457, n48458, n48459,
    n48460, n48461, n48462, n48463, n48464, n48465, n48466, n48467, n48468,
    n48469, n48470, n48471, n48472, n48473, n48474, n48476, n48477, n48478,
    n48479, n48480, n48481, n48482, n48483, n48484, n48485, n48486, n48487,
    n48488, n48489, n48490, n48491, n48492, n48493, n48494, n48495, n48496,
    n48497, n48498, n48499, n48500, n48501, n48502, n48503, n48504, n48505,
    n48506, n48507, n48508, n48509, n48510, n48511, n48512, n48513, n48514,
    n48515, n48516, n48517, n48518, n48520, n48521, n48522, n48523, n48524,
    n48525, n48526, n48527, n48528, n48529, n48530, n48531, n48532, n48533,
    n48534, n48535, n48536, n48537, n48538, n48539, n48540, n48541, n48542,
    n48543, n48544, n48545, n48546, n48547, n48548, n48549, n48550, n48551,
    n48552, n48553, n48554, n48555, n48557, n48558, n48559, n48560, n48561,
    n48562, n48563, n48564, n48565, n48566, n48567, n48568, n48569, n48570,
    n48571, n48572, n48573, n48574, n48575, n48576, n48577, n48578, n48579,
    n48580, n48581, n48582, n48583, n48584, n48585, n48586, n48587, n48588,
    n48589, n48590, n48592, n48593, n48594, n48595, n48596, n48597, n48598,
    n48599, n48600, n48601, n48602, n48603, n48604, n48605, n48606, n48607,
    n48608, n48609, n48610, n48611, n48612, n48613, n48614, n48615, n48616,
    n48617, n48618, n48619, n48620, n48621, n48622, n48623, n48624, n48625,
    n48626, n48627, n48628, n48629, n48630, n48631, n48633, n48634, n48635,
    n48636, n48637, n48638, n48639, n48640, n48641, n48642, n48643, n48644,
    n48645, n48646, n48647, n48648, n48649, n48650, n48651, n48652, n48653,
    n48654, n48655, n48656, n48657, n48658, n48659, n48660, n48661, n48662,
    n48663, n48664, n48665, n48666, n48668, n48669, n48670, n48671, n48672,
    n48673, n48674, n48675, n48676, n48677, n48678, n48679, n48680, n48681,
    n48682, n48683, n48684, n48685, n48686, n48687, n48688, n48689, n48690,
    n48691, n48692, n48693, n48694, n48695, n48696, n48697, n48698, n48699,
    n48700, n48701, n48702, n48703, n48705, n48706, n48707, n48708, n48709,
    n48710, n48711, n48712, n48713, n48714, n48715, n48716, n48717, n48718,
    n48719, n48720, n48721, n48722, n48723, n48724, n48725, n48726, n48727,
    n48728, n48729, n48730, n48731, n48732, n48733, n48734, n48735, n48736,
    n48737, n48738, n48739, n48740, n48741, n48742, n48743, n48744, n48745,
    n48746, n48747, n48748, n48749, n48751, n48752, n48753, n48754, n48755,
    n48756, n48757, n48758, n48759, n48760, n48761, n48762, n48763, n48764,
    n48765, n48766, n48767, n48768, n48769, n48770, n48771, n48772, n48773,
    n48774, n48775, n48776, n48777, n48778, n48779, n48780, n48781, n48782,
    n48783, n48784, n48785, n48786, n48788, n48789, n48790, n48791, n48792,
    n48793, n48794, n48795, n48796, n48797, n48798, n48799, n48800, n48801,
    n48802, n48803, n48804, n48805, n48806, n48807, n48808, n48809, n48810,
    n48811, n48812, n48813, n48814, n48815, n48816, n48818, n48819, n48820,
    n48821, n48822, n48823, n48824, n48825, n48826, n48827, n48828, n48829,
    n48830, n48831, n48832, n48833, n48834, n48835, n48836, n48837, n48838,
    n48839, n48840, n48841, n48842, n48843, n48844, n48845, n48846, n48847,
    n48848, n48849, n48850, n48851, n48852, n48853, n48854, n48855, n48856,
    n48858, n48859, n48860, n48861, n48862, n48863, n48864, n48865, n48866,
    n48867, n48868, n48869, n48870, n48871, n48872, n48873, n48874, n48875,
    n48876, n48877, n48878, n48879, n48880, n48881, n48882, n48883, n48884,
    n48885, n48886, n48887, n48888, n48889, n48890, n48891, n48893, n48894,
    n48895, n48896, n48897, n48898, n48899, n48900, n48901, n48902, n48903,
    n48904, n48905, n48906, n48907, n48908, n48909, n48910, n48911, n48912,
    n48913, n48914, n48915, n48916, n48917, n48918, n48919, n48920, n48921,
    n48923, n48924, n48925, n48926, n48927, n48928, n48929, n48930, n48931,
    n48932, n48933, n48934, n48935, n48936, n48937, n48938, n48939, n48940,
    n48941, n48942, n48943, n48944, n48945, n48946, n48947, n48948, n48949,
    n48951, n48952, n48953, n48954, n48955, n48956, n48957, n48958, n48959,
    n48960, n48961, n48962, n48963, n48964, n48965, n48966, n48967, n48968,
    n48969, n48970, n48971, n48972, n48973, n48974, n48975, n48976, n48977,
    n48978, n48979, n48980, n48981, n48982, n48983, n48984, n48985, n48986,
    n48987, n48988, n48989, n48990, n48991, n48992, n48993, n48994, n48995,
    n48996, n48997, n48998, n48999, n49000, n49001, n49002, n49003, n49004,
    n49005, n49006, n49007, n49008, n49009, n49010, n49011, n49012, n49013,
    n49014, n49015, n49016, n49017, n49018, n49019, n49020, n49021, n49022,
    n49023, n49024, n49025, n49026, n49027, n49028, n49029, n49030, n49031,
    n49032, n49033, n49034, n49035, n49036, n49037, n49038, n49039, n49040,
    n49041, n49042, n49043, n49044, n49045, n49046, n49047, n49048, n49049,
    n49050, n49051, n49053, n49054, n49055, n49056, n49057, n49058, n49059,
    n49060, n49061, n49062, n49063, n49064, n49065, n49066, n49067, n49068,
    n49069, n49070, n49071, n49072, n49073, n49074, n49075, n49076, n49077,
    n49078, n49079, n49080, n49081, n49082, n49083, n49084, n49085, n49086,
    n49087, n49088, n49089, n49090, n49091, n49092, n49093, n49094, n49095,
    n49096, n49097, n49098, n49099, n49100, n49102, n49103, n49104, n49105,
    n49106, n49107, n49108, n49109, n49110, n49111, n49112, n49113, n49114,
    n49115, n49116, n49117, n49118, n49119, n49120, n49121, n49122, n49123,
    n49124, n49125, n49126, n49127, n49128, n49129, n49130, n49131, n49132,
    n49133, n49135, n49136, n49137, n49138, n49139, n49140, n49141, n49142,
    n49143, n49144, n49145, n49146, n49147, n49148, n49149, n49150, n49151,
    n49152, n49153, n49154, n49155, n49156, n49157, n49158, n49159, n49160,
    n49161, n49162, n49163, n49164, n49165, n49166, n49167, n49168, n49169,
    n49170, n49171, n49172, n49173, n49174, n49175, n49176, n49177, n49178,
    n49179, n49180, n49181, n49182, n49183, n49184, n49185, n49186, n49187,
    n49188, n49189, n49190, n49191, n49192, n49193, n49194, n49195, n49196,
    n49197, n49198, n49199, n49200, n49201, n49202, n49203, n49204, n49205,
    n49206, n49207, n49208, n49209, n49210, n49211, n49212, n49213, n49214,
    n49215, n49216, n49217, n49218, n49219, n49220, n49221, n49222, n49223,
    n49224, n49226, n49227, n49228, n49229, n49230, n49231, n49232, n49233,
    n49234, n49235, n49236, n49237, n49238, n49239, n49240, n49241, n49242,
    n49243, n49244, n49245, n49246, n49247, n49248, n49249, n49250, n49251,
    n49252, n49253, n49254, n49255, n49256, n49257, n49258, n49259, n49260,
    n49261, n49262, n49263, n49264, n49265, n49266, n49267, n49268, n49269,
    n49270, n49271, n49272, n49273, n49274, n49275, n49276, n49277, n49278,
    n49279, n49280, n49281, n49282, n49283, n49284, n49285, n49286, n49287,
    n49288, n49289, n49290, n49291, n49292, n49293, n49294, n49295, n49296,
    n49297, n49298, n49299, n49300, n49301, n49302, n49303, n49304, n49305,
    n49306, n49307, n49308, n49309, n49310, n49311, n49312, n49313, n49314,
    n49315, n49316, n49317, n49318, n49319, n49320, n49321, n49322, n49323,
    n49324, n49326, n49327, n49328, n49329, n49330, n49331, n49332, n49333,
    n49334, n49335, n49336, n49337, n49338, n49339, n49340, n49341, n49342,
    n49343, n49344, n49345, n49346, n49347, n49348, n49349, n49350, n49351,
    n49352, n49353, n49354, n49355, n49356, n49357, n49358, n49359, n49360,
    n49361, n49362, n49363, n49364, n49365, n49366, n49367, n49368, n49369,
    n49370, n49371, n49372, n49373, n49374, n49375, n49376, n49377, n49378,
    n49379, n49380, n49381, n49382, n49383, n49384, n49385, n49386, n49387,
    n49388, n49389, n49390, n49391, n49392, n49393, n49394, n49395, n49396,
    n49397, n49398, n49399, n49400, n49401, n49402, n49403, n49404, n49405,
    n49406, n49407, n49408, n49409, n49410, n49411, n49412, n49413, n49414,
    n49415, n49416, n49417, n49418, n49419, n49420, n49421, n49422, n49423,
    n49424, n49425, n49426, n49427, n49428, n49429, n49431, n49432, n49433,
    n49434, n49435, n49436, n49437, n49438, n49439, n49440, n49441, n49442,
    n49443, n49444, n49445, n49446, n49447, n49448, n49449, n49450, n49451,
    n49452, n49453, n49454, n49455, n49456, n49457, n49458, n49459, n49460,
    n49461, n49462, n49463, n49464, n49465, n49466, n49467, n49468, n49469,
    n49470, n49471, n49472, n49473, n49474, n49475, n49476, n49477, n49478,
    n49479, n49480, n49481, n49482, n49483, n49484, n49485, n49486, n49487,
    n49488, n49489, n49490, n49491, n49492, n49493, n49494, n49495, n49496,
    n49497, n49498, n49499, n49500, n49501, n49502, n49503, n49504, n49505,
    n49506, n49507, n49508, n49509, n49510, n49511, n49512, n49513, n49514,
    n49515, n49516, n49517, n49518, n49519, n49520, n49521, n49522, n49523,
    n49524, n49525, n49526, n49527, n49528, n49529, n49530, n49531, n49533,
    n49534, n49535, n49536, n49537, n49538, n49539, n49540, n49541, n49542,
    n49543, n49544, n49545, n49546, n49547, n49548, n49549, n49550, n49551,
    n49552, n49553, n49554, n49555, n49556, n49557, n49558, n49559, n49560,
    n49561, n49562, n49563, n49564, n49565, n49566, n49567, n49568, n49569,
    n49570, n49571, n49572, n49573, n49574, n49575, n49576, n49577, n49578,
    n49579, n49580, n49581, n49582, n49583, n49585, n49586, n49587, n49588,
    n49589, n49590, n49591, n49592, n49593, n49594, n49595, n49596, n49597,
    n49598, n49599, n49600, n49601, n49602, n49603, n49604, n49605, n49606,
    n49607, n49608, n49609, n49610, n49611, n49612, n49613, n49614, n49615,
    n49616, n49617, n49618, n49619, n49620, n49621, n49622, n49624, n49625,
    n49626, n49627, n49628, n49629, n49630, n49631, n49632, n49633, n49634,
    n49635, n49636, n49637, n49638, n49639, n49640, n49641, n49642, n49643,
    n49644, n49645, n49646, n49647, n49648, n49649, n49650, n49651, n49652,
    n49653, n49654, n49655, n49656, n49657, n49658, n49659, n49660, n49661,
    n49662, n49663, n49665, n49666, n49667, n49668, n49669, n49670, n49671,
    n49672, n49673, n49674, n49675, n49676, n49677, n49678, n49679, n49680,
    n49681, n49682, n49683, n49684, n49685, n49686, n49687, n49688, n49689,
    n49690, n49691, n49692, n49693, n49694, n49695, n49696, n49697, n49698,
    n49699, n49700, n49701, n49702, n49703, n49704, n49705, n49706, n49707,
    n49708, n49709, n49710, n49711, n49712, n49713, n49714, n49715, n49716,
    n49717, n49718, n49719, n49720, n49721, n49722, n49723, n49724, n49725,
    n49726, n49727, n49728, n49729, n49730, n49731, n49732, n49733, n49734,
    n49735, n49736, n49737, n49738, n49739, n49740, n49741, n49742, n49743,
    n49744, n49745, n49746, n49747, n49748, n49749, n49750, n49751, n49752,
    n49753, n49754, n49755, n49756, n49757, n49758, n49759, n49760, n49761,
    n49762, n49763, n49764, n49765, n49766, n49767, n49768, n49769, n49771,
    n49772, n49773, n49774, n49775, n49776, n49777, n49778, n49779, n49780,
    n49781, n49782, n49783, n49784, n49785, n49786, n49787, n49788, n49789,
    n49790, n49791, n49792, n49793, n49794, n49795, n49796, n49797, n49798,
    n49799, n49800, n49801, n49802, n49803, n49804, n49805, n49806, n49807,
    n49808, n49810, n49811, n49812, n49813, n49814, n49815, n49816, n49817,
    n49818, n49819, n49820, n49821, n49822, n49823, n49824, n49825, n49826,
    n49827, n49828, n49829, n49830, n49831, n49832, n49833, n49834, n49835,
    n49836, n49837, n49838, n49839, n49840, n49841, n49843, n49844, n49845,
    n49846, n49847, n49848, n49849, n49850, n49851, n49852, n49853, n49854,
    n49855, n49856, n49857, n49858, n49859, n49860, n49861, n49862, n49863,
    n49864, n49865, n49866, n49867, n49868, n49869, n49870, n49871, n49872,
    n49873, n49874, n49875, n49876, n49877, n49878, n49879, n49880, n49881,
    n49882, n49884, n49885, n49886, n49887, n49888, n49889, n49890, n49891,
    n49892, n49893, n49894, n49895, n49896, n49897, n49898, n49899, n49900,
    n49901, n49902, n49903, n49904, n49905, n49906, n49907, n49908, n49909,
    n49910, n49911, n49912, n49913, n49914, n49915, n49916, n49917, n49918,
    n49920, n49921, n49922, n49923, n49924, n49925, n49926, n49927, n49928,
    n49929, n49930, n49931, n49932, n49933, n49934, n49935, n49936, n49937,
    n49938, n49939, n49940, n49941, n49942, n49943, n49944, n49945, n49946,
    n49947, n49948, n49949, n49950, n49951, n49952, n49953, n49955, n49956,
    n49957, n49958, n49959, n49960, n49961, n49962, n49963, n49964, n49965,
    n49966, n49967, n49968, n49969, n49970, n49971, n49972, n49973, n49974,
    n49975, n49976, n49977, n49978, n49979, n49980, n49981, n49982, n49983,
    n49985, n49986, n49987, n49988, n49989, n49990, n49991, n49992, n49993,
    n49994, n49995, n49996, n49997, n49998, n49999, n50000, n50001, n50002,
    n50003, n50004, n50005, n50006, n50007, n50008, n50009, n50010, n50011,
    n50013, n50014, n50015, n50016, n50017, n50018, n50019, n50020, n50021,
    n50022, n50023, n50024, n50025, n50026, n50027, n50028, n50029, n50030,
    n50031, n50032, n50033, n50034, n50035, n50036, n50037, n50038, n50039,
    n50040, n50041, n50042, n50043, n50044, n50045, n50046, n50047, n50048,
    n50049, n50050, n50051, n50052, n50053, n50054, n50055, n50056, n50057,
    n50058, n50059, n50060, n50061, n50062, n50063, n50064, n50065, n50066,
    n50067, n50068, n50069, n50070, n50071, n50072, n50073, n50074, n50075,
    n50076, n50077, n50078, n50079, n50080, n50081, n50082, n50083, n50084,
    n50085, n50086, n50087, n50088, n50089, n50090, n50091, n50092, n50093,
    n50094, n50095, n50096, n50097, n50098, n50099, n50100, n50101, n50102,
    n50103, n50104, n50105, n50106, n50107, n50108, n50109, n50110, n50112,
    n50113, n50114, n50115, n50116, n50117, n50118, n50119, n50120, n50121,
    n50122, n50123, n50124, n50125, n50126, n50127, n50128, n50129, n50130,
    n50131, n50132, n50133, n50134, n50135, n50136, n50137, n50138, n50139,
    n50140, n50141, n50142, n50143, n50144, n50145, n50146, n50147, n50148,
    n50149, n50151, n50152, n50153, n50154, n50155, n50156, n50157, n50158,
    n50159, n50160, n50161, n50162, n50163, n50164, n50165, n50166, n50167,
    n50168, n50169, n50170, n50171, n50172, n50173, n50174, n50175, n50176,
    n50177, n50178, n50179, n50180, n50181, n50182, n50183, n50184, n50185,
    n50186, n50187, n50188, n50189, n50190, n50191, n50192, n50194, n50195,
    n50196, n50197, n50198, n50199, n50200, n50201, n50202, n50203, n50204,
    n50205, n50206, n50207, n50208, n50209, n50210, n50211, n50212, n50213,
    n50214, n50215, n50216, n50217, n50218, n50219, n50220, n50221, n50222,
    n50223, n50224, n50225, n50226, n50227, n50228, n50230, n50231, n50232,
    n50233, n50234, n50235, n50236, n50237, n50238, n50239, n50240, n50241,
    n50242, n50243, n50244, n50245, n50246, n50247, n50248, n50249, n50250,
    n50251, n50252, n50253, n50254, n50255, n50256, n50257, n50258, n50259,
    n50260, n50261, n50262, n50263, n50264, n50265, n50266, n50267, n50268,
    n50269, n50270, n50271, n50272, n50273, n50274, n50275, n50276, n50277,
    n50278, n50279, n50280, n50281, n50282, n50283, n50284, n50285, n50286,
    n50287, n50288, n50289, n50290, n50291, n50292, n50293, n50294, n50295,
    n50296, n50297, n50298, n50299, n50300, n50301, n50302, n50303, n50304,
    n50305, n50306, n50307, n50308, n50309, n50310, n50311, n50312, n50313,
    n50314, n50315, n50316, n50317, n50318, n50319, n50320, n50321, n50322,
    n50323, n50324, n50325, n50326, n50327, n50328, n50329, n50330, n50331,
    n50332, n50333, n50334, n50335, n50337, n50338, n50339, n50340, n50341,
    n50342, n50343, n50344, n50345, n50346, n50347, n50348, n50349, n50350,
    n50351, n50352, n50353, n50354, n50355, n50356, n50357, n50358, n50359,
    n50360, n50361, n50362, n50363, n50364, n50365, n50366, n50367, n50368,
    n50369, n50370, n50371, n50372, n50373, n50374, n50375, n50376, n50377,
    n50378, n50379, n50380, n50381, n50382, n50384, n50385, n50386, n50387,
    n50388, n50389, n50390, n50391, n50392, n50393, n50394, n50395, n50396,
    n50397, n50398, n50399, n50400, n50401, n50402, n50403, n50404, n50405,
    n50406, n50407, n50408, n50409, n50410, n50411, n50412, n50413, n50414,
    n50415, n50416, n50417, n50419, n50420, n50421, n50422, n50423, n50424,
    n50425, n50426, n50427, n50428, n50429, n50430, n50431, n50432, n50433,
    n50434, n50435, n50436, n50437, n50438, n50439, n50440, n50441, n50442,
    n50443, n50444, n50445, n50446, n50447, n50448, n50449, n50450, n50451,
    n50452, n50453, n50454, n50455, n50456, n50458, n50459, n50460, n50461,
    n50462, n50463, n50464, n50465, n50466, n50467, n50468, n50469, n50470,
    n50471, n50472, n50473, n50474, n50475, n50476, n50477, n50478, n50479,
    n50480, n50481, n50482, n50483, n50484, n50485, n50486, n50487, n50488,
    n50489, n50490, n50491, n50492, n50493, n50494, n50495, n50496, n50498,
    n50499, n50500, n50501, n50502, n50503, n50504, n50505, n50506, n50507,
    n50508, n50509, n50510, n50511, n50512, n50513, n50514, n50515, n50516,
    n50517, n50518, n50519, n50520, n50521, n50522, n50523, n50524, n50525,
    n50526, n50527, n50528, n50529, n50530, n50531, n50532, n50534, n50535,
    n50536, n50537, n50538, n50539, n50540, n50541, n50542, n50543, n50544,
    n50545, n50546, n50547, n50548, n50549, n50550, n50551, n50552, n50553,
    n50554, n50555, n50556, n50557, n50558, n50559, n50560, n50561, n50562,
    n50563, n50564, n50565, n50566, n50567, n50568, n50569, n50570, n50571,
    n50572, n50574, n50575, n50576, n50577, n50578, n50579, n50580, n50581,
    n50582, n50583, n50584, n50585, n50586, n50587, n50588, n50589, n50590,
    n50591, n50592, n50593, n50594, n50595, n50596, n50597, n50598, n50599,
    n50600, n50601, n50602, n50603, n50604, n50605, n50606, n50607, n50608,
    n50609, n50610, n50612, n50613, n50614, n50615, n50616, n50617, n50618,
    n50619, n50620, n50621, n50622, n50623, n50624, n50625, n50626, n50627,
    n50628, n50629, n50630, n50631, n50632, n50633, n50634, n50635, n50636,
    n50637, n50638, n50639, n50640, n50641, n50642, n50643, n50644, n50645,
    n50647, n50648, n50649, n50650, n50651, n50652, n50653, n50654, n50655,
    n50656, n50657, n50658, n50659, n50660, n50661, n50662, n50663, n50664,
    n50665, n50666, n50667, n50668, n50669, n50670, n50671, n50672, n50673,
    n50674, n50675, n50677, n50678, n50679, n50680, n50681, n50682, n50683,
    n50684, n50685, n50686, n50687, n50688, n50689, n50690, n50691, n50692,
    n50693, n50694, n50695, n50696, n50697, n50698, n50699, n50700, n50701,
    n50702, n50703, n50704, n50705, n50706, n50707, n50708, n50709, n50710,
    n50711, n50712, n50713, n50714, n50715, n50716, n50717, n50718, n50719,
    n50720, n50721, n50722, n50723, n50724, n50725, n50726, n50727, n50728,
    n50729, n50730, n50731, n50732, n50733, n50734, n50735, n50736, n50737,
    n50738, n50739, n50740, n50741, n50742, n50743, n50744, n50745, n50746,
    n50747, n50748, n50749, n50750, n50751, n50752, n50753, n50754, n50755,
    n50756, n50757, n50758, n50759, n50760, n50761, n50762, n50763, n50764,
    n50765, n50766, n50767, n50768, n50769, n50770, n50771, n50772, n50773,
    n50774, n50775, n50776, n50778, n50779, n50780, n50781, n50782, n50783,
    n50784, n50785, n50786, n50787, n50788, n50789, n50790, n50791, n50792,
    n50793, n50794, n50795, n50796, n50797, n50798, n50799, n50800, n50801,
    n50802, n50803, n50804, n50805, n50806, n50807, n50808, n50809, n50810,
    n50811, n50812, n50813, n50814, n50815, n50816, n50817, n50818, n50819,
    n50820, n50821, n50822, n50823, n50824, n50825, n50826, n50827, n50828,
    n50829, n50830, n50831, n50832, n50833, n50834, n50835, n50836, n50837,
    n50838, n50839, n50840, n50841, n50842, n50843, n50844, n50845, n50846,
    n50847, n50848, n50849, n50850, n50851, n50852, n50853, n50854, n50855,
    n50856, n50857, n50858, n50859, n50860, n50861, n50862, n50863, n50864,
    n50865, n50866, n50867, n50868, n50869, n50870, n50871, n50872, n50873,
    n50874, n50875, n50876, n50877, n50878, n50879, n50880, n50882, n50883,
    n50884, n50885, n50886, n50887, n50888, n50889, n50890, n50891, n50892,
    n50893, n50894, n50895, n50896, n50897, n50898, n50899, n50900, n50901,
    n50902, n50903, n50904, n50905, n50906, n50907, n50908, n50909, n50910,
    n50911, n50912, n50914, n50915, n50916, n50917, n50918, n50919, n50920,
    n50921, n50922, n50923, n50924, n50925, n50926, n50927, n50928, n50929,
    n50930, n50931, n50932, n50933, n50934, n50935, n50936, n50937, n50938,
    n50939, n50940, n50941, n50942, n50943, n50944, n50945, n50946, n50947,
    n50948, n50949, n50950, n50951, n50952, n50953, n50954, n50955, n50956,
    n50957, n50958, n50959, n50960, n50961, n50962, n50963, n50964, n50965,
    n50966, n50967, n50968, n50969, n50970, n50971, n50972, n50973, n50974,
    n50975, n50976, n50977, n50978, n50979, n50980, n50981, n50982, n50983,
    n50984, n50985, n50986, n50987, n50988, n50989, n50990, n50991, n50992,
    n50993, n50994, n50995, n50996, n50997, n50998, n50999, n51000, n51001,
    n51002, n51003, n51004, n51005, n51006, n51007, n51008, n51009, n51010,
    n51011, n51012, n51013, n51014, n51015, n51016, n51017, n51018, n51019,
    n51020, n51021, n51022, n51023, n51024, n51025, n51026, n51028, n51029,
    n51030, n51031, n51032, n51033, n51034, n51035, n51036, n51037, n51038,
    n51039, n51040, n51041, n51042, n51043, n51044, n51045, n51046, n51047,
    n51048, n51049, n51050, n51051, n51052, n51053, n51054, n51055, n51056,
    n51057, n51058, n51059, n51060, n51061, n51062, n51063, n51064, n51065,
    n51066, n51067, n51068, n51069, n51070, n51071, n51072, n51073, n51074,
    n51075, n51076, n51077, n51078, n51079, n51080, n51081, n51082, n51083,
    n51084, n51085, n51086, n51087, n51088, n51089, n51090, n51091, n51092,
    n51093, n51094, n51095, n51096, n51097, n51098, n51099, n51100, n51101,
    n51102, n51103, n51104, n51105, n51106, n51107, n51108, n51109, n51110,
    n51111, n51112, n51113, n51114, n51115, n51116, n51117, n51118, n51119,
    n51120, n51121, n51122, n51123, n51124, n51125, n51126, n51127, n51128,
    n51129, n51130, n51131, n51133, n51134, n51135, n51136, n51137, n51138,
    n51139, n51140, n51141, n51142, n51143, n51144, n51145, n51146, n51147,
    n51148, n51149, n51150, n51151, n51152, n51153, n51154, n51155, n51156,
    n51157, n51158, n51159, n51160, n51161, n51162, n51163, n51164, n51165,
    n51166, n51167, n51168, n51169, n51170, n51171, n51172, n51173, n51174,
    n51175, n51176, n51177, n51178, n51179, n51180, n51181, n51182, n51183,
    n51184, n51185, n51186, n51187, n51188, n51189, n51190, n51191, n51192,
    n51193, n51194, n51195, n51196, n51197, n51198, n51199, n51200, n51201,
    n51202, n51203, n51204, n51205, n51206, n51207, n51208, n51209, n51210,
    n51211, n51212, n51213, n51214, n51215, n51216, n51217, n51218, n51219,
    n51220, n51221, n51222, n51223, n51224, n51225, n51226, n51227, n51228,
    n51229, n51230, n51231, n51232, n51233, n51234, n51235, n51237, n51238,
    n51239, n51240, n51241, n51242, n51243, n51244, n51245, n51246, n51247,
    n51248, n51249, n51250, n51251, n51252, n51253, n51254, n51255, n51256,
    n51257, n51258, n51259, n51260, n51261, n51262, n51263, n51264, n51265,
    n51266, n51267, n51268, n51269, n51270, n51271, n51272, n51273, n51274,
    n51275, n51276, n51277, n51278, n51279, n51280, n51281, n51282, n51283,
    n51284, n51285, n51286, n51287, n51288, n51289, n51290, n51291, n51292,
    n51293, n51294, n51295, n51296, n51297, n51298, n51299, n51300, n51301,
    n51302, n51303, n51304, n51305, n51306, n51307, n51308, n51309, n51310,
    n51311, n51312, n51313, n51314, n51315, n51316, n51317, n51318, n51319,
    n51320, n51321, n51322, n51323, n51324, n51325, n51326, n51327, n51328,
    n51329, n51330, n51331, n51332, n51333, n51334, n51336, n51337, n51338,
    n51339, n51340, n51341, n51342, n51343, n51344, n51345, n51346, n51347,
    n51348, n51349, n51350, n51351, n51352, n51353, n51354, n51355, n51356,
    n51357, n51358, n51359, n51360, n51361, n51362, n51363, n51364, n51365,
    n51366, n51367, n51368, n51369, n51370, n51371, n51372, n51373, n51374,
    n51375, n51376, n51377, n51378, n51379, n51380, n51381, n51383, n51384,
    n51385, n51386, n51387, n51388, n51389, n51390, n51391, n51392, n51393,
    n51394, n51395, n51396, n51397, n51398, n51399, n51400, n51401, n51402,
    n51403, n51404, n51405, n51406, n51407, n51408, n51409, n51410, n51411,
    n51412, n51413, n51414, n51415, n51416, n51417, n51418, n51419, n51420,
    n51421, n51422, n51423, n51425, n51426, n51427, n51428, n51429, n51430,
    n51431, n51432, n51433, n51434, n51435, n51436, n51437, n51438, n51439,
    n51440, n51441, n51442, n51443, n51444, n51445, n51446, n51447, n51448,
    n51449, n51450, n51451, n51452, n51453, n51454, n51455, n51456, n51457,
    n51458, n51459, n51460, n51461, n51462, n51463, n51464, n51465, n51466,
    n51468, n51469, n51470, n51471, n51472, n51473, n51474, n51475, n51476,
    n51477, n51478, n51479, n51480, n51481, n51482, n51483, n51484, n51485,
    n51486, n51487, n51488, n51489, n51490, n51491, n51492, n51493, n51494,
    n51495, n51496, n51497, n51498, n51499, n51500, n51501, n51502, n51503,
    n51504, n51505, n51506, n51507, n51508, n51510, n51511, n51512, n51513,
    n51514, n51515, n51516, n51517, n51518, n51519, n51520, n51521, n51522,
    n51523, n51524, n51525, n51526, n51527, n51528, n51529, n51530, n51531,
    n51532, n51533, n51534, n51535, n51536, n51537, n51538, n51539, n51540,
    n51541, n51542, n51543, n51544, n51545, n51546, n51547, n51548, n51549,
    n51550, n51551, n51552, n51553, n51554, n51555, n51556, n51557, n51558,
    n51559, n51560, n51561, n51562, n51563, n51564, n51565, n51566, n51567,
    n51568, n51569, n51570, n51571, n51572, n51573, n51574, n51575, n51576,
    n51577, n51578, n51579, n51580, n51581, n51582, n51583, n51584, n51585,
    n51586, n51587, n51588, n51589, n51590, n51591, n51592, n51593, n51594,
    n51595, n51596, n51597, n51598, n51599, n51600, n51602, n51603, n51604,
    n51605, n51606, n51607, n51608, n51609, n51610, n51611, n51612, n51613,
    n51614, n51615, n51616, n51617, n51618, n51619, n51620, n51621, n51622,
    n51623, n51624, n51625, n51626, n51627, n51628, n51629, n51630, n51631,
    n51632, n51633, n51634, n51635, n51636, n51637, n51638, n51639, n51640,
    n51642, n51643, n51644, n51645, n51646, n51647, n51648, n51649, n51650,
    n51651, n51652, n51653, n51654, n51655, n51656, n51657, n51658, n51659,
    n51660, n51661, n51662, n51663, n51664, n51665, n51666, n51667, n51668,
    n51669, n51670, n51671, n51672, n51673, n51674, n51675, n51676, n51677,
    n51679, n51680, n51681, n51682, n51683, n51684, n51685, n51686, n51687,
    n51688, n51689, n51690, n51691, n51692, n51693, n51694, n51695, n51696,
    n51697, n51698, n51699, n51700, n51701, n51702, n51703, n51704, n51705,
    n51706, n51707, n51708, n51709, n51710, n51711, n51712, n51713, n51714,
    n51715, n51716, n51717, n51719, n51720, n51721, n51722, n51723, n51724,
    n51725, n51726, n51727, n51728, n51729, n51730, n51731, n51732, n51733,
    n51734, n51735, n51736, n51737, n51738, n51739, n51740, n51741, n51742,
    n51743, n51744, n51745, n51746, n51747, n51748, n51749, n51750, n51751,
    n51752, n51753, n51754, n51755, n51756, n51757, n51758, n51759, n51760,
    n51761, n51762, n51763, n51764, n51765, n51766, n51767, n51768, n51770,
    n51771, n51772, n51773, n51774, n51775, n51776, n51777, n51778, n51779,
    n51780, n51781, n51782, n51783, n51784, n51785, n51786, n51787, n51788,
    n51789, n51790, n51791, n51792, n51793, n51794, n51795, n51796, n51797,
    n51798, n51799, n51800, n51801, n51802, n51803, n51804, n51805, n51807,
    n51808, n51809, n51810, n51811, n51812, n51813, n51814, n51815, n51816,
    n51817, n51818, n51819, n51820, n51821, n51822, n51823, n51824, n51825,
    n51826, n51827, n51828, n51829, n51830, n51831, n51832, n51833, n51834,
    n51835, n51836, n51837, n51838, n51839, n51841, n51842, n51843, n51844,
    n51845, n51846, n51847, n51848, n51849, n51850, n51851, n51852, n51853,
    n51854, n51855, n51856, n51857, n51858, n51859, n51860, n51861, n51862,
    n51863, n51864, n51865, n51866, n51867, n51868, n51869, n51870, n51871,
    n51872, n51873, n51874, n51876, n51877, n51878, n51879, n51880, n51881,
    n51882, n51883, n51884, n51885, n51886, n51887, n51888, n51889, n51890,
    n51891, n51892, n51893, n51894, n51895, n51896, n51897, n51898, n51899,
    n51900, n51901, n51902, n51903, n51904, n51905, n51906, n51907, n51908,
    n51909, n51910, n51911, n51913, n51914, n51915, n51916, n51917, n51918,
    n51919, n51920, n51921, n51922, n51923, n51924, n51925, n51926, n51927,
    n51928, n51929, n51930, n51931, n51932, n51933, n51934, n51935, n51936,
    n51937, n51938, n51939, n51940, n51941, n51942, n51943, n51944, n51945,
    n51946, n51947, n51948, n51949, n51950, n51951, n51952, n51953, n51954,
    n51955, n51956, n51957, n51958, n51959, n51960, n51961, n51962, n51963,
    n51964, n51965, n51966, n51967, n51968, n51969, n51970, n51971, n51972,
    n51973, n51974, n51975, n51976, n51977, n51978, n51979, n51980, n51981,
    n51982, n51983, n51984, n51985, n51986, n51987, n51988, n51989, n51990,
    n51991, n51992, n51993, n51994, n51995, n51996, n51997, n51998, n51999,
    n52000, n52001, n52002, n52003, n52004, n52005, n52006, n52007, n52008,
    n52010, n52011, n52012, n52013, n52014, n52015, n52016, n52017, n52018,
    n52019, n52020, n52021, n52022, n52023, n52024, n52025, n52026, n52027,
    n52028, n52029, n52030, n52031, n52032, n52033, n52034, n52035, n52036,
    n52037, n52039, n52040, n52041, n52042, n52043, n52044, n52045, n52046,
    n52047, n52048, n52049, n52050, n52051, n52052, n52053, n52054, n52055,
    n52056, n52057, n52058, n52059, n52060, n52061, n52062, n52063, n52064,
    n52065, n52066, n52067, n52068, n52069, n52070, n52071, n52072, n52073,
    n52074, n52075, n52076, n52077, n52078, n52079, n52080, n52081, n52082,
    n52083, n52084, n52086, n52087, n52088, n52089, n52090, n52091, n52092,
    n52093, n52094, n52095, n52096, n52097, n52098, n52099, n52100, n52101,
    n52102, n52103, n52104, n52105, n52106, n52107, n52108, n52109, n52110,
    n52111, n52112, n52113, n52114, n52115, n52116, n52117, n52118, n52119,
    n52120, n52121, n52122, n52123, n52124, n52125, n52126, n52127, n52129,
    n52130, n52131, n52132, n52133, n52134, n52135, n52136, n52137, n52138,
    n52139, n52140, n52141, n52142, n52143, n52144, n52145, n52146, n52147,
    n52148, n52149, n52150, n52151, n52152, n52153, n52154, n52155, n52156,
    n52157, n52158, n52159, n52160, n52161, n52162, n52163, n52164, n52165,
    n52166, n52167, n52168, n52169, n52170, n52171, n52172, n52173, n52175,
    n52176, n52177, n52178, n52179, n52180, n52181, n52182, n52183, n52184,
    n52185, n52186, n52187, n52188, n52189, n52190, n52191, n52192, n52193,
    n52194, n52195, n52196, n52197, n52198, n52199, n52200, n52201, n52202,
    n52203, n52204, n52205, n52206, n52207, n52209, n52210, n52211, n52212,
    n52213, n52214, n52215, n52216, n52217, n52218, n52219, n52220, n52221,
    n52222, n52223, n52224, n52225, n52226, n52227, n52228, n52229, n52230,
    n52231, n52232, n52233, n52234, n52235, n52236, n52237, n52238, n52239,
    n52240, n52241, n52242, n52244, n52245, n52246, n52247, n52248, n52249,
    n52250, n52251, n52252, n52253, n52254, n52255, n52256, n52257, n52258,
    n52259, n52260, n52261, n52262, n52263, n52264, n52265, n52266, n52267,
    n52268, n52269, n52270, n52271, n52272, n52273, n52274, n52275, n52276,
    n52277, n52278, n52279, n52280, n52281, n52282, n52283, n52285, n52286,
    n52287, n52288, n52289, n52290, n52291, n52292, n52293, n52294, n52295,
    n52296, n52297, n52298, n52299, n52300, n52301, n52302, n52303, n52304,
    n52305, n52306, n52307, n52308, n52309, n52310, n52311, n52312, n52313,
    n52315, n52316, n52317, n52318, n52319, n52320, n52321, n52322, n52323,
    n52324, n52325, n52326, n52327, n52328, n52329, n52330, n52331, n52332,
    n52333, n52334, n52335, n52336, n52337, n52338, n52339, n52340, n52341,
    n52342, n52343, n52344, n52346, n52347, n52348, n52349, n52350, n52351,
    n52352, n52353, n52354, n52355, n52356, n52357, n52358, n52359, n52360,
    n52361, n52362, n52363, n52364, n52365, n52366, n52367, n52368, n52369,
    n52370, n52371, n52372, n52373, n52374, n52375, n52376, n52377, n52378,
    n52379, n52381, n52382, n52383, n52384, n52385, n52386, n52387, n52388,
    n52389, n52390, n52391, n52392, n52393, n52394, n52395, n52396, n52397,
    n52398, n52399, n52400, n52401, n52402, n52403, n52404, n52405, n52407,
    n52408, n52409, n52410, n52411, n52412, n52413, n52414, n52415, n52416,
    n52417, n52418, n52419, n52420, n52421, n52422, n52423, n52424, n52425,
    n52426, n52427, n52428, n52429, n52430, n52431, n52432, n52433, n52434,
    n52435, n52436, n52437, n52438, n52439, n52440, n52441, n52442, n52443,
    n52444, n52445, n52446, n52447, n52448, n52449, n52450, n52451, n52452,
    n52453, n52454, n52455, n52456, n52457, n52458, n52459, n52460, n52461,
    n52462, n52463, n52464, n52465, n52466, n52467, n52468, n52469, n52470,
    n52471, n52472, n52473, n52474, n52475, n52476, n52477, n52478, n52479,
    n52480, n52481, n52482, n52483, n52484, n52485, n52486, n52487, n52488,
    n52489, n52490, n52491, n52492, n52493, n52494, n52495, n52496, n52497,
    n52498, n52499, n52500, n52501, n52502, n52503, n52504, n52505, n52506,
    n52507, n52508, n52510, n52511, n52512, n52513, n52514, n52515, n52516,
    n52517, n52518, n52519, n52520, n52521, n52522, n52523, n52524, n52525,
    n52526, n52527, n52528, n52529, n52530, n52531, n52532, n52533, n52534,
    n52535, n52536, n52537, n52538, n52539, n52540, n52541, n52542, n52543,
    n52544, n52545, n52546, n52547, n52548, n52549, n52550, n52551, n52552,
    n52553, n52554, n52555, n52556, n52557, n52558, n52559, n52560, n52561,
    n52562, n52563, n52564, n52565, n52566, n52567, n52568, n52569, n52570,
    n52571, n52572, n52573, n52574, n52575, n52576, n52577, n52578, n52579,
    n52580, n52581, n52582, n52583, n52584, n52585, n52586, n52587, n52588,
    n52589, n52590, n52591, n52592, n52593, n52594, n52595, n52596, n52597,
    n52598, n52599, n52600, n52601, n52602, n52603, n52604, n52605, n52606,
    n52607, n52608, n52609, n52610, n52611, n52612, n52613, n52614, n52615,
    n52616, n52617, n52619, n52620, n52621, n52622, n52623, n52624, n52625,
    n52626, n52627, n52628, n52629, n52630, n52631, n52632, n52633, n52634,
    n52635, n52636, n52637, n52638, n52639, n52640, n52641, n52642, n52643,
    n52644, n52645, n52646, n52647, n52648, n52649, n52650, n52651, n52652,
    n52653, n52654, n52655, n52656, n52657, n52658, n52659, n52660, n52661,
    n52662, n52663, n52664, n52665, n52666, n52667, n52668, n52669, n52670,
    n52671, n52672, n52673, n52674, n52675, n52676, n52677, n52678, n52679,
    n52680, n52681, n52682, n52683, n52684, n52685, n52686, n52687, n52688,
    n52689, n52690, n52691, n52692, n52693, n52694, n52695, n52696, n52697,
    n52698, n52699, n52700, n52701, n52702, n52703, n52704, n52705, n52706,
    n52707, n52708, n52709, n52710, n52711, n52712, n52713, n52714, n52715,
    n52716, n52717, n52718, n52720, n52721, n52722, n52723, n52724, n52725,
    n52726, n52727, n52728, n52729, n52730, n52731, n52732, n52733, n52734,
    n52735, n52736, n52737, n52738, n52739, n52740, n52741, n52742, n52743,
    n52744, n52745, n52746, n52747, n52748, n52749, n52750, n52751, n52752,
    n52753, n52754, n52755, n52756, n52757, n52758, n52759, n52760, n52761,
    n52762, n52763, n52764, n52765, n52766, n52767, n52768, n52769, n52770,
    n52771, n52772, n52773, n52774, n52775, n52776, n52777, n52778, n52779,
    n52780, n52781, n52782, n52783, n52784, n52785, n52786, n52787, n52788,
    n52789, n52790, n52791, n52792, n52793, n52794, n52795, n52796, n52797,
    n52798, n52799, n52800, n52801, n52802, n52803, n52804, n52805, n52806,
    n52807, n52808, n52809, n52810, n52811, n52812, n52813, n52814, n52815,
    n52816, n52817, n52818, n52820, n52821, n52822, n52823, n52824, n52825,
    n52826, n52827, n52828, n52829, n52830, n52831, n52832, n52833, n52834,
    n52835, n52836, n52837, n52838, n52839, n52840, n52841, n52842, n52843,
    n52844, n52845, n52846, n52847, n52848, n52849, n52850, n52851, n52852,
    n52853, n52854, n52855, n52856, n52857, n52858, n52859, n52860, n52861,
    n52862, n52863, n52864, n52865, n52867, n52868, n52869, n52870, n52871,
    n52872, n52873, n52874, n52875, n52876, n52877, n52878, n52879, n52880,
    n52881, n52882, n52883, n52884, n52885, n52886, n52887, n52888, n52889,
    n52890, n52891, n52892, n52893, n52894, n52895, n52896, n52897, n52898,
    n52899, n52900, n52901, n52902, n52903, n52904, n52905, n52906, n52907,
    n52908, n52909, n52910, n52911, n52912, n52913, n52914, n52915, n52916,
    n52917, n52918, n52919, n52920, n52921, n52922, n52923, n52924, n52925,
    n52926, n52927, n52928, n52929, n52930, n52931, n52932, n52933, n52934,
    n52935, n52936, n52937, n52938, n52939, n52940, n52941, n52942, n52943,
    n52944, n52945, n52946, n52947, n52948, n52949, n52950, n52951, n52952,
    n52953, n52954, n52955, n52956, n52957, n52958, n52959, n52960, n52961,
    n52962, n52963, n52964, n52965, n52966, n52967, n52969, n52970, n52971,
    n52972, n52973, n52974, n52975, n52976, n52977, n52978, n52979, n52980,
    n52981, n52982, n52983, n52984, n52985, n52986, n52987, n52988, n52989,
    n52990, n52991, n52992, n52993, n52994, n52995, n52996, n52997, n52998,
    n52999, n53000, n53001, n53002, n53003, n53004, n53005, n53006, n53007,
    n53008, n53009, n53010, n53011, n53012, n53013, n53014, n53015, n53016,
    n53017, n53018, n53019, n53020, n53021, n53022, n53023, n53024, n53025,
    n53026, n53027, n53028, n53029, n53030, n53031, n53032, n53033, n53034,
    n53035, n53036, n53037, n53038, n53039, n53040, n53041, n53042, n53043,
    n53044, n53045, n53046, n53047, n53048, n53049, n53050, n53051, n53052,
    n53053, n53054, n53055, n53056, n53057, n53058, n53060, n53061, n53062,
    n53063, n53064, n53065, n53066, n53067, n53068, n53069, n53070, n53071,
    n53072, n53073, n53074, n53075, n53076, n53077, n53078, n53079, n53080,
    n53081, n53082, n53083, n53084, n53085, n53086, n53087, n53088, n53089,
    n53090, n53091, n53092, n53093, n53094, n53095, n53096, n53097, n53098,
    n53099, n53100, n53101, n53102, n53103, n53104, n53105, n53107, n53108,
    n53109, n53110, n53111, n53112, n53113, n53114, n53115, n53116, n53117,
    n53118, n53119, n53120, n53121, n53122, n53123, n53124, n53125, n53126,
    n53127, n53128, n53129, n53130, n53131, n53132, n53133, n53134, n53135,
    n53136, n53137, n53138, n53139, n53140, n53142, n53143, n53144, n53145,
    n53146, n53147, n53148, n53149, n53150, n53151, n53152, n53153, n53154,
    n53155, n53156, n53157, n53158, n53159, n53160, n53161, n53162, n53163,
    n53164, n53165, n53166, n53167, n53168, n53169, n53170, n53171, n53172,
    n53173, n53175, n53176, n53177, n53178, n53179, n53180, n53181, n53182,
    n53183, n53184, n53185, n53186, n53187, n53188, n53189, n53190, n53191,
    n53192, n53193, n53194, n53195, n53196, n53197, n53198, n53199, n53200,
    n53201, n53202, n53203, n53204, n53205, n53206, n53207, n53208, n53209,
    n53210, n53211, n53212, n53213, n53215, n53216, n53217, n53218, n53219,
    n53220, n53221, n53222, n53223, n53224, n53225, n53226, n53227, n53228,
    n53229, n53230, n53231, n53232, n53233, n53234, n53235, n53236, n53237,
    n53238, n53239, n53240, n53241, n53242, n53243, n53244, n53245, n53246,
    n53247, n53248, n53249, n53250, n53251, n53252, n53253, n53254, n53255,
    n53256, n53257, n53258, n53259, n53260, n53261, n53262, n53263, n53265,
    n53266, n53267, n53268, n53269, n53270, n53271, n53272, n53273, n53274,
    n53275, n53276, n53277, n53278, n53279, n53280, n53281, n53282, n53283,
    n53284, n53285, n53286, n53287, n53288, n53289, n53290, n53291, n53292,
    n53293, n53294, n53295, n53296, n53297, n53298, n53299, n53300, n53301,
    n53303, n53304, n53305, n53306, n53307, n53308, n53309, n53310, n53311,
    n53312, n53313, n53314, n53315, n53316, n53317, n53318, n53319, n53320,
    n53321, n53322, n53323, n53324, n53325, n53326, n53327, n53328, n53329,
    n53330, n53331, n53332, n53333, n53334, n53335, n53336, n53337, n53338,
    n53339, n53340, n53341, n53342, n53343, n53344, n53345, n53346, n53347,
    n53348, n53349, n53350, n53351, n53352, n53353, n53354, n53355, n53356,
    n53357, n53358, n53359, n53360, n53361, n53362, n53363, n53364, n53365,
    n53366, n53367, n53368, n53369, n53370, n53371, n53372, n53373, n53374,
    n53375, n53376, n53377, n53378, n53379, n53380, n53381, n53382, n53383,
    n53384, n53385, n53386, n53387, n53388, n53389, n53390, n53391, n53392,
    n53393, n53394, n53395, n53396, n53398, n53399, n53400, n53401, n53402,
    n53403, n53404, n53405, n53406, n53407, n53408, n53409, n53410, n53411,
    n53412, n53413, n53414, n53415, n53416, n53417, n53418, n53419, n53420,
    n53421, n53422, n53423, n53424, n53425, n53426, n53427, n53428, n53429,
    n53430, n53431, n53432, n53433, n53434, n53435, n53436, n53437, n53438,
    n53439, n53440, n53441, n53442, n53444, n53445, n53446, n53447, n53448,
    n53449, n53450, n53451, n53452, n53453, n53454, n53455, n53456, n53457,
    n53458, n53459, n53460, n53461, n53462, n53463, n53464, n53465, n53466,
    n53467, n53468, n53469, n53470, n53471, n53472, n53473, n53474, n53475,
    n53476, n53477, n53478, n53479, n53480, n53481, n53482, n53483, n53484,
    n53485, n53486, n53487, n53488, n53489, n53490, n53491, n53492, n53493,
    n53494, n53495, n53496, n53497, n53498, n53499, n53500, n53501, n53502,
    n53503, n53504, n53505, n53506, n53507, n53508, n53509, n53510, n53511,
    n53512, n53513, n53514, n53515, n53516, n53517, n53518, n53519, n53520,
    n53521, n53522, n53523, n53524, n53525, n53526, n53527, n53528, n53529,
    n53530, n53531, n53532, n53533, n53534, n53535, n53536, n53537, n53538,
    n53540, n53541, n53542, n53543, n53544, n53545, n53546, n53547, n53548,
    n53549, n53550, n53551, n53552, n53553, n53554, n53555, n53556, n53557,
    n53558, n53559, n53560, n53561, n53562, n53563, n53564, n53565, n53566,
    n53567, n53569, n53570, n53571, n53572, n53573, n53574, n53575, n53576,
    n53577, n53578, n53579, n53580, n53581, n53582, n53583, n53584, n53585,
    n53586, n53587, n53588, n53589, n53590, n53591, n53592, n53593, n53594,
    n53595, n53596, n53597, n53598, n53599, n53600, n53601, n53602, n53603,
    n53604, n53605, n53607, n53608, n53609, n53610, n53611, n53612, n53613,
    n53614, n53615, n53616, n53617, n53618, n53619, n53620, n53621, n53622,
    n53623, n53624, n53625, n53626, n53627, n53628, n53629, n53630, n53631,
    n53632, n53633, n53634, n53635, n53636, n53637, n53638, n53639, n53640,
    n53641, n53642, n53643, n53644, n53645, n53647, n53648, n53649, n53650,
    n53651, n53652, n53653, n53654, n53655, n53656, n53657, n53658, n53659,
    n53660, n53661, n53662, n53663, n53664, n53665, n53666, n53667, n53668,
    n53669, n53670, n53671, n53672, n53673, n53674, n53675, n53676, n53677,
    n53678, n53679, n53680, n53681, n53682, n53683, n53684, n53685, n53686,
    n53687, n53688, n53689, n53690, n53692, n53693, n53694, n53695, n53696,
    n53697, n53698, n53699, n53700, n53701, n53702, n53703, n53704, n53705,
    n53706, n53707, n53708, n53709, n53710, n53711, n53712, n53713, n53714,
    n53715, n53716, n53717, n53718, n53719, n53720, n53722, n53723, n53724,
    n53725, n53726, n53727, n53728, n53729, n53730, n53731, n53732, n53733,
    n53734, n53735, n53736, n53737, n53738, n53739, n53740, n53741, n53742,
    n53743, n53744, n53745, n53746, n53747, n53748, n53749, n53750, n53751,
    n53752, n53753, n53754, n53755, n53756, n53757, n53758, n53759, n53760,
    n53761, n53762, n53763, n53764, n53765, n53766, n53767, n53769, n53770,
    n53771, n53772, n53773, n53774, n53775, n53776, n53777, n53778, n53779,
    n53780, n53781, n53782, n53783, n53784, n53785, n53786, n53787, n53788,
    n53789, n53790, n53791, n53792, n53793, n53794, n53795, n53796, n53797,
    n53798, n53799, n53800, n53801, n53802, n53803, n53804, n53805, n53806,
    n53807, n53808, n53809, n53811, n53812, n53813, n53814, n53815, n53816,
    n53817, n53818, n53819, n53820, n53821, n53822, n53823, n53824, n53825,
    n53826, n53827, n53828, n53829, n53830, n53831, n53832, n53833, n53834,
    n53835, n53836, n53837, n53838, n53839, n53840, n53841, n53842, n53843,
    n53844, n53846, n53847, n53848, n53849, n53850, n53851, n53852, n53853,
    n53854, n53855, n53856, n53857, n53858, n53859, n53860, n53861, n53862,
    n53863, n53864, n53865, n53866, n53867, n53868, n53869, n53870, n53871,
    n53872, n53873, n53874, n53875, n53876, n53877, n53878, n53879, n53880,
    n53881, n53882, n53883, n53884, n53885, n53886, n53887, n53889, n53890,
    n53891, n53892, n53893, n53894, n53895, n53896, n53897, n53898, n53899,
    n53900, n53901, n53902, n53903, n53904, n53905, n53906, n53907, n53908,
    n53909, n53910, n53911, n53912, n53913, n53914, n53915, n53916, n53917,
    n53918, n53919, n53920, n53921, n53922, n53923, n53924, n53925, n53926,
    n53928, n53929, n53930, n53931, n53932, n53933, n53934, n53935, n53936,
    n53937, n53938, n53939, n53940, n53941, n53942, n53943, n53944, n53945,
    n53946, n53947, n53948, n53949, n53950, n53951, n53952, n53953, n53954,
    n53955, n53956, n53957, n53958, n53959, n53960, n53961, n53962, n53963,
    n53965, n53966, n53967, n53968, n53969, n53970, n53971, n53972, n53973,
    n53974, n53975, n53976, n53977, n53978, n53979, n53980, n53981, n53982,
    n53983, n53984, n53985, n53986, n53987, n53988, n53989, n53990, n53991,
    n53992, n53993, n53994, n53995, n53996, n53997, n53998, n53999, n54000,
    n54002, n54003, n54004, n54005, n54006, n54007, n54008, n54009, n54010,
    n54011, n54012, n54013, n54014, n54015, n54016, n54017, n54018, n54019,
    n54020, n54021, n54022, n54023, n54024, n54025, n54026, n54027, n54028,
    n54029, n54030, n54031, n54032, n54033, n54034, n54035, n54036, n54037,
    n54039, n54040, n54041, n54042, n54043, n54044, n54045, n54046, n54047,
    n54048, n54049, n54050, n54051, n54052, n54053, n54054, n54055, n54056,
    n54057, n54058, n54059, n54060, n54061, n54062, n54063, n54064, n54065,
    n54066, n54067, n54068, n54069, n54070, n54071, n54073, n54074, n54075,
    n54076, n54077, n54078, n54079, n54080, n54081, n54082, n54083, n54084,
    n54085, n54086, n54087, n54088, n54089, n54090, n54091, n54092, n54093,
    n54094, n54095, n54096, n54097, n54098, n54099, n54100, n54101, n54103,
    n54104, n54105, n54106, n54107, n54108, n54109, n54110, n54111, n54112,
    n54113, n54114, n54115, n54116, n54117, n54118, n54119, n54120, n54121,
    n54122, n54123, n54124, n54125, n54126, n54127, n54129, n54130, n54131,
    n54132, n54133, n54134, n54135, n54136, n54137, n54138, n54139, n54140,
    n54141, n54142, n54143, n54144, n54145, n54146, n54147, n54148, n54149,
    n54150, n54151, n54152, n54153, n54154, n54155, n54156, n54157, n54158,
    n54159, n54160, n54161, n54162, n54163, n54164, n54165, n54166, n54167,
    n54168, n54169, n54170, n54171, n54172, n54173, n54174, n54175, n54176,
    n54177, n54178, n54179, n54180, n54181, n54182, n54183, n54184, n54185,
    n54186, n54187, n54188, n54189, n54190, n54191, n54192, n54193, n54194,
    n54195, n54196, n54197, n54198, n54199, n54200, n54201, n54202, n54203,
    n54204, n54205, n54206, n54207, n54208, n54209, n54210, n54211, n54212,
    n54213, n54214, n54215, n54216, n54217, n54218, n54219, n54220, n54221,
    n54222, n54223, n54224, n54225, n54226, n54227, n54228, n54229, n54230,
    n54231, n54232, n54233, n54235, n54236, n54237, n54238, n54239, n54240,
    n54241, n54242, n54243, n54244, n54245, n54246, n54247, n54248, n54249,
    n54250, n54251, n54252, n54253, n54254, n54255, n54256, n54257, n54258,
    n54259, n54260, n54261, n54262, n54263, n54264, n54265, n54266, n54267,
    n54268, n54269, n54270, n54271, n54272, n54273, n54274, n54275, n54276,
    n54277, n54278, n54279, n54280, n54281, n54282, n54283, n54284, n54285,
    n54286, n54287, n54288, n54289, n54290, n54291, n54292, n54293, n54294,
    n54295, n54296, n54297, n54298, n54299, n54300, n54301, n54302, n54303,
    n54304, n54305, n54306, n54307, n54308, n54309, n54310, n54311, n54312,
    n54313, n54314, n54315, n54316, n54317, n54318, n54319, n54320, n54321,
    n54322, n54323, n54324, n54325, n54326, n54327, n54328, n54329, n54330,
    n54331, n54332, n54333, n54334, n54335, n54337, n54338, n54339, n54340,
    n54341, n54342, n54343, n54344, n54345, n54346, n54347, n54348, n54349,
    n54350, n54351, n54352, n54353, n54354, n54355, n54356, n54357, n54358,
    n54359, n54360, n54361, n54362, n54363, n54364, n54365, n54366, n54367,
    n54368, n54369, n54370, n54371, n54372, n54373, n54374, n54375, n54376,
    n54377, n54379, n54380, n54381, n54382, n54383, n54384, n54385, n54386,
    n54387, n54388, n54389, n54390, n54391, n54392, n54393, n54394, n54395,
    n54396, n54397, n54398, n54399, n54400, n54401, n54402, n54403, n54404,
    n54405, n54406, n54407, n54408, n54410, n54411, n54412, n54413, n54414,
    n54415, n54416, n54417, n54418, n54419, n54420, n54421, n54422, n54423,
    n54424, n54425, n54426, n54427, n54428, n54429, n54430, n54431, n54432,
    n54433, n54434, n54435, n54436, n54437, n54438, n54439, n54440, n54441,
    n54442, n54443, n54444, n54445, n54446, n54447, n54448, n54449, n54450,
    n54451, n54452, n54453, n54454, n54455, n54456, n54457, n54458, n54459,
    n54460, n54461, n54462, n54463, n54464, n54465, n54466, n54467, n54468,
    n54469, n54470, n54471, n54472, n54473, n54474, n54475, n54476, n54477,
    n54478, n54479, n54480, n54481, n54482, n54483, n54484, n54485, n54486,
    n54487, n54488, n54489, n54490, n54491, n54492, n54493, n54494, n54495,
    n54496, n54497, n54498, n54499, n54500, n54501, n54502, n54503, n54504,
    n54505, n54506, n54508, n54509, n54510, n54511, n54512, n54513, n54514,
    n54515, n54516, n54517, n54518, n54519, n54520, n54521, n54522, n54523,
    n54524, n54525, n54526, n54527, n54528, n54529, n54530, n54531, n54532,
    n54533, n54534, n54535, n54536, n54537, n54538, n54539, n54540, n54541,
    n54542, n54543, n54544, n54545, n54546, n54547, n54548, n54549, n54550,
    n54551, n54552, n54553, n54554, n54555, n54556, n54557, n54558, n54559,
    n54560, n54561, n54562, n54563, n54564, n54565, n54566, n54567, n54568,
    n54569, n54570, n54571, n54572, n54573, n54574, n54575, n54576, n54577,
    n54578, n54579, n54580, n54581, n54582, n54583, n54584, n54585, n54586,
    n54587, n54588, n54589, n54590, n54591, n54592, n54593, n54594, n54595,
    n54596, n54597, n54598, n54599, n54600, n54601, n54602, n54603, n54604,
    n54605, n54606, n54607, n54608, n54609, n54610, n54611, n54612, n54613,
    n54615, n54616, n54617, n54618, n54619, n54620, n54621, n54622, n54623,
    n54624, n54625, n54626, n54627, n54628, n54629, n54630, n54631, n54632,
    n54633, n54634, n54635, n54636, n54637, n54638, n54639, n54640, n54641,
    n54642, n54643, n54644, n54645, n54646, n54647, n54648, n54649, n54650,
    n54651, n54652, n54653, n54654, n54655, n54656, n54657, n54658, n54659,
    n54660, n54661, n54662, n54663, n54664, n54665, n54666, n54667, n54668,
    n54669, n54670, n54671, n54672, n54673, n54674, n54675, n54676, n54677,
    n54678, n54679, n54680, n54681, n54682, n54683, n54684, n54685, n54686,
    n54687, n54688, n54689, n54690, n54691, n54692, n54693, n54694, n54695,
    n54696, n54697, n54698, n54699, n54700, n54701, n54702, n54703, n54704,
    n54705, n54706, n54707, n54708, n54709, n54710, n54711, n54712, n54713,
    n54714, n54715, n54716, n54717, n54718, n54720, n54721, n54722, n54723,
    n54724, n54725, n54726, n54727, n54728, n54729, n54730, n54731, n54732,
    n54733, n54734, n54735, n54736, n54737, n54738, n54739, n54740, n54741,
    n54742, n54743, n54744, n54745, n54746, n54747, n54748, n54749, n54750,
    n54751, n54752, n54753, n54754, n54756, n54757, n54758, n54759, n54760,
    n54761, n54762, n54763, n54764, n54765, n54766, n54767, n54768, n54769,
    n54770, n54771, n54772, n54773, n54774, n54775, n54776, n54777, n54778,
    n54779, n54780, n54781, n54782, n54783, n54784, n54785, n54786, n54787,
    n54788, n54789, n54790, n54791, n54792, n54793, n54794, n54795, n54796,
    n54797, n54798, n54799, n54800, n54801, n54802, n54803, n54804, n54805,
    n54806, n54807, n54808, n54809, n54810, n54811, n54812, n54813, n54814,
    n54815, n54816, n54817, n54818, n54819, n54820, n54821, n54822, n54823,
    n54824, n54825, n54826, n54827, n54828, n54829, n54830, n54831, n54832,
    n54833, n54834, n54835, n54836, n54837, n54838, n54839, n54840, n54841,
    n54842, n54843, n54844, n54845, n54846, n54847, n54848, n54849, n54850,
    n54851, n54852, n54853, n54854, n54855, n54856, n54857, n54858, n54860,
    n54861, n54862, n54863, n54864, n54865, n54866, n54867, n54868, n54869,
    n54870, n54871, n54872, n54873, n54874, n54875, n54876, n54877, n54878,
    n54879, n54880, n54881, n54882, n54883, n54884, n54885, n54886, n54887,
    n54888, n54889, n54890, n54891, n54892, n54893, n54894, n54895, n54896,
    n54897, n54898, n54899, n54900, n54901, n54902, n54903, n54904, n54905,
    n54906, n54907, n54909, n54910, n54911, n54912, n54913, n54914, n54915,
    n54916, n54917, n54918, n54919, n54920, n54921, n54922, n54923, n54924,
    n54925, n54926, n54927, n54928, n54929, n54930, n54931, n54932, n54933,
    n54934, n54935, n54936, n54937, n54938, n54939, n54940, n54941, n54942,
    n54943, n54944, n54945, n54946, n54947, n54949, n54950, n54951, n54952,
    n54953, n54954, n54955, n54956, n54957, n54958, n54959, n54960, n54961,
    n54962, n54963, n54964, n54965, n54966, n54967, n54968, n54969, n54970,
    n54971, n54972, n54973, n54974, n54975, n54976, n54977, n54978, n54979,
    n54980, n54981, n54982, n54983, n54984, n54985, n54986, n54987, n54988,
    n54989, n54990, n54992, n54993, n54994, n54995, n54996, n54997, n54998,
    n54999, n55000, n55001, n55002, n55003, n55004, n55005, n55006, n55007,
    n55008, n55009, n55010, n55011, n55012, n55013, n55014, n55015, n55016,
    n55017, n55018, n55019, n55020, n55021, n55022, n55023, n55024, n55025,
    n55026, n55027, n55028, n55029, n55030, n55032, n55033, n55034, n55035,
    n55036, n55037, n55038, n55039, n55040, n55041, n55042, n55043, n55044,
    n55045, n55046, n55047, n55048, n55049, n55050, n55051, n55052, n55053,
    n55054, n55055, n55056, n55057, n55058, n55059, n55060, n55061, n55062,
    n55063, n55064, n55065, n55066, n55067, n55068, n55069, n55070, n55071,
    n55072, n55073, n55074, n55075, n55076, n55077, n55078, n55079, n55080,
    n55081, n55082, n55083, n55084, n55085, n55086, n55087, n55088, n55089,
    n55090, n55091, n55092, n55093, n55094, n55095, n55096, n55097, n55098,
    n55099, n55100, n55101, n55102, n55103, n55104, n55105, n55106, n55107,
    n55108, n55109, n55110, n55111, n55112, n55113, n55114, n55115, n55116,
    n55117, n55118, n55119, n55120, n55121, n55122, n55123, n55124, n55125,
    n55126, n55128, n55129, n55130, n55131, n55132, n55133, n55134, n55135,
    n55136, n55137, n55138, n55139, n55140, n55141, n55142, n55143, n55144,
    n55145, n55146, n55147, n55148, n55149, n55150, n55151, n55152, n55153,
    n55154, n55155, n55156, n55158, n55159, n55160, n55161, n55162, n55163,
    n55164, n55165, n55166, n55167, n55168, n55169, n55170, n55171, n55172,
    n55173, n55174, n55175, n55176, n55177, n55178, n55179, n55180, n55181,
    n55182, n55183, n55184, n55185, n55186, n55187, n55188, n55189, n55190,
    n55191, n55192, n55193, n55194, n55195, n55196, n55197, n55198, n55199,
    n55200, n55201, n55202, n55204, n55205, n55206, n55207, n55208, n55209,
    n55210, n55211, n55212, n55213, n55214, n55215, n55216, n55217, n55218,
    n55219, n55220, n55221, n55222, n55223, n55224, n55225, n55226, n55227,
    n55228, n55229, n55230, n55231, n55232, n55233, n55234, n55235, n55236,
    n55238, n55239, n55240, n55241, n55242, n55243, n55244, n55245, n55246,
    n55247, n55248, n55249, n55250, n55251, n55252, n55253, n55254, n55255,
    n55256, n55257, n55258, n55259, n55260, n55261, n55262, n55263, n55264,
    n55265, n55266, n55267, n55268, n55269, n55270, n55271, n55272, n55273,
    n55274, n55275, n55276, n55277, n55278, n55279, n55280, n55281, n55283,
    n55284, n55285, n55286, n55287, n55288, n55289, n55290, n55291, n55292,
    n55293, n55294, n55295, n55296, n55297, n55298, n55299, n55300, n55301,
    n55302, n55303, n55304, n55305, n55306, n55307, n55308, n55309, n55310,
    n55311, n55312, n55313, n55314, n55315, n55316, n55317, n55318, n55319,
    n55321, n55322, n55323, n55324, n55325, n55326, n55327, n55328, n55329,
    n55330, n55331, n55332, n55333, n55334, n55335, n55336, n55337, n55338,
    n55339, n55340, n55341, n55342, n55343, n55344, n55345, n55346, n55347,
    n55348, n55349, n55350, n55352, n55353, n55354, n55355, n55356, n55357,
    n55358, n55359, n55360, n55361, n55362, n55363, n55364, n55365, n55366,
    n55367, n55368, n55369, n55370, n55371, n55372, n55373, n55374, n55375,
    n55376, n55377, n55378, n55379, n55380, n55381, n55382, n55383, n55384,
    n55385, n55386, n55387, n55388, n55389, n55390, n55391, n55392, n55393,
    n55394, n55395, n55396, n55397, n55398, n55399, n55400, n55401, n55402,
    n55403, n55404, n55405, n55406, n55407, n55408, n55409, n55410, n55411,
    n55412, n55413, n55414, n55415, n55416, n55417, n55418, n55419, n55420,
    n55421, n55422, n55423, n55424, n55425, n55426, n55427, n55428, n55429,
    n55430, n55431, n55432, n55433, n55434, n55435, n55436, n55437, n55438,
    n55439, n55440, n55441, n55442, n55443, n55444, n55445, n55446, n55447,
    n55448, n55450, n55451, n55452, n55453, n55454, n55455, n55456, n55457,
    n55458, n55459, n55460, n55461, n55462, n55463, n55464, n55465, n55466,
    n55467, n55468, n55469, n55470, n55471, n55472, n55473, n55474, n55475,
    n55476, n55477, n55478, n55479, n55480, n55481, n55482, n55483, n55484,
    n55485, n55486, n55487, n55489, n55490, n55491, n55492, n55493, n55494,
    n55495, n55496, n55497, n55498, n55499, n55500, n55501, n55502, n55503,
    n55504, n55505, n55506, n55507, n55508, n55509, n55510, n55511, n55512,
    n55513, n55514, n55515, n55516, n55517, n55518, n55519, n55520, n55521,
    n55522, n55523, n55524, n55525, n55526, n55528, n55529, n55530, n55531,
    n55532, n55533, n55534, n55535, n55536, n55537, n55538, n55539, n55540,
    n55541, n55542, n55543, n55544, n55545, n55546, n55547, n55548, n55549,
    n55550, n55551, n55552, n55553, n55554, n55555, n55556, n55557, n55558,
    n55559, n55560, n55561, n55562, n55563, n55564, n55565, n55566, n55567,
    n55569, n55570, n55571, n55572, n55573, n55574, n55575, n55576, n55577,
    n55578, n55579, n55580, n55581, n55582, n55583, n55584, n55585, n55586,
    n55587, n55588, n55589, n55590, n55591, n55592, n55593, n55594, n55595,
    n55596, n55597, n55598, n55599, n55600, n55601, n55602, n55604, n55605,
    n55606, n55607, n55608, n55609, n55610, n55611, n55612, n55613, n55614,
    n55615, n55616, n55617, n55618, n55619, n55620, n55621, n55622, n55623,
    n55624, n55625, n55626, n55627, n55628, n55629, n55630, n55631, n55632,
    n55633, n55634, n55635, n55636, n55637, n55638, n55639, n55640, n55641,
    n55642, n55643, n55644, n55646, n55647, n55648, n55649, n55650, n55651,
    n55652, n55653, n55654, n55655, n55656, n55657, n55658, n55659, n55660,
    n55661, n55662, n55663, n55664, n55665, n55666, n55667, n55668, n55669,
    n55670, n55671, n55672, n55673, n55674, n55675, n55676, n55677, n55678,
    n55679, n55680, n55681, n55683, n55684, n55685, n55686, n55687, n55688,
    n55689, n55690, n55691, n55692, n55693, n55694, n55695, n55696, n55697,
    n55698, n55699, n55700, n55701, n55702, n55703, n55704, n55705, n55706,
    n55707, n55708, n55709, n55710, n55711, n55713, n55714, n55715, n55716,
    n55717, n55718, n55719, n55720, n55721, n55722, n55723, n55724, n55725,
    n55726, n55727, n55728, n55729, n55730, n55731, n55732, n55733, n55734,
    n55735, n55736, n55737, n55738, n55739, n55740, n55741, n55742, n55743,
    n55744, n55745, n55746, n55747, n55748, n55749, n55750, n55751, n55753,
    n55754, n55755, n55756, n55757, n55758, n55759, n55760, n55761, n55762,
    n55763, n55764, n55765, n55766, n55767, n55768, n55769, n55770, n55771,
    n55772, n55773, n55774, n55775, n55776, n55777, n55778, n55779, n55780,
    n55781, n55782, n55783, n55784, n55785, n55786, n55787, n55789, n55790,
    n55791, n55792, n55793, n55794, n55795, n55796, n55797, n55798, n55799,
    n55800, n55801, n55802, n55803, n55804, n55805, n55806, n55807, n55808,
    n55809, n55810, n55811, n55812, n55813, n55814, n55815, n55816, n55817,
    n55818, n55819, n55820, n55821, n55822, n55823, n55824, n55826, n55827,
    n55828, n55829, n55830, n55831, n55832, n55833, n55834, n55835, n55836,
    n55837, n55838, n55839, n55840, n55841, n55842, n55843, n55844, n55845,
    n55846, n55847, n55848, n55849, n55850, n55852, n55853, n55854, n55855,
    n55856, n55857, n55858, n55859, n55860, n55861, n55862, n55863, n55864,
    n55865, n55866, n55867, n55868, n55869, n55870, n55871, n55872, n55873,
    n55874, n55875, n55876, n55877, n55878, n55879, n55880, n55881, n55882,
    n55883, n55884, n55885, n55886, n55887, n55888, n55889, n55890, n55891,
    n55892, n55893, n55894, n55895, n55896, n55897, n55898, n55899, n55900,
    n55901, n55902, n55903, n55904, n55905, n55906, n55907, n55908, n55909,
    n55910, n55911, n55912, n55913, n55914, n55915, n55916, n55917, n55918,
    n55919, n55920, n55921, n55922, n55923, n55924, n55925, n55926, n55927,
    n55928, n55929, n55930, n55931, n55932, n55933, n55934, n55935, n55936,
    n55937, n55938, n55939, n55940, n55941, n55942, n55943, n55944, n55945,
    n55946, n55947, n55948, n55949, n55950, n55951, n55952, n55953, n55955,
    n55956, n55957, n55958, n55959, n55960, n55961, n55962, n55963, n55964,
    n55965, n55966, n55967, n55968, n55969, n55970, n55971, n55972, n55973,
    n55974, n55975, n55976, n55977, n55978, n55979, n55980, n55981, n55982,
    n55983, n55984, n55985, n55986, n55987, n55988, n55989, n55990, n55991,
    n55992, n55993, n55994, n55995, n55996, n55997, n55998, n55999, n56000,
    n56001, n56002, n56003, n56004, n56005, n56006, n56007, n56008, n56009,
    n56010, n56011, n56012, n56013, n56014, n56015, n56016, n56017, n56018,
    n56019, n56020, n56021, n56022, n56023, n56024, n56025, n56026, n56027,
    n56028, n56029, n56030, n56031, n56032, n56033, n56034, n56035, n56036,
    n56037, n56038, n56039, n56040, n56041, n56042, n56043, n56044, n56045,
    n56046, n56047, n56048, n56049, n56050, n56051, n56052, n56053, n56054,
    n56055, n56056, n56057, n56058, n56059, n56060, n56061, n56062, n56063,
    n56064, n56066, n56067, n56068, n56069, n56070, n56071, n56072, n56073,
    n56074, n56075, n56076, n56077, n56078, n56079, n56080, n56081, n56082,
    n56083, n56084, n56085, n56086, n56087, n56088, n56089, n56090, n56091,
    n56092, n56093, n56094, n56095, n56096, n56097, n56098, n56099, n56100,
    n56101, n56102, n56103, n56104, n56105, n56106, n56107, n56108, n56109,
    n56110, n56111, n56112, n56113, n56114, n56115, n56116, n56117, n56118,
    n56119, n56120, n56121, n56122, n56123, n56124, n56125, n56126, n56127,
    n56128, n56129, n56130, n56131, n56132, n56133, n56134, n56135, n56136,
    n56137, n56138, n56139, n56140, n56141, n56142, n56143, n56144, n56145,
    n56146, n56147, n56148, n56149, n56150, n56151, n56152, n56153, n56154,
    n56155, n56156, n56157, n56158, n56159, n56160, n56161, n56162, n56163,
    n56164, n56166, n56167, n56168, n56169, n56170, n56171, n56172, n56173,
    n56174, n56175, n56176, n56177, n56178, n56179, n56180, n56181, n56182,
    n56183, n56184, n56185, n56186, n56187, n56188, n56189, n56190, n56191,
    n56192, n56193, n56194, n56195, n56196, n56197, n56198, n56199, n56200,
    n56201, n56202, n56203, n56204, n56205, n56206, n56207, n56208, n56209,
    n56210, n56211, n56212, n56213, n56214, n56215, n56216, n56217, n56218,
    n56219, n56220, n56221, n56222, n56223, n56224, n56225, n56226, n56227,
    n56228, n56229, n56230, n56231, n56232, n56233, n56234, n56235, n56236,
    n56237, n56238, n56239, n56240, n56241, n56242, n56243, n56244, n56245,
    n56246, n56247, n56248, n56249, n56250, n56251, n56252, n56253, n56254,
    n56255, n56256, n56257, n56258, n56259, n56260, n56261, n56262, n56263,
    n56264, n56266, n56267, n56268, n56269, n56270, n56271, n56272, n56273,
    n56274, n56275, n56276, n56277, n56278, n56279, n56280, n56281, n56282,
    n56283, n56284, n56285, n56286, n56287, n56288, n56289, n56290, n56291,
    n56292, n56293, n56294, n56295, n56296, n56297, n56298, n56299, n56300,
    n56301, n56302, n56303, n56304, n56305, n56306, n56307, n56308, n56309,
    n56310, n56311, n56312, n56313, n56314, n56315, n56316, n56317, n56318,
    n56319, n56320, n56321, n56322, n56323, n56324, n56325, n56326, n56327,
    n56328, n56329, n56330, n56331, n56332, n56333, n56334, n56335, n56336,
    n56337, n56338, n56339, n56340, n56341, n56342, n56343, n56344, n56345,
    n56346, n56347, n56348, n56349, n56350, n56351, n56352, n56353, n56354,
    n56355, n56356, n56357, n56358, n56359, n56360, n56361, n56362, n56363,
    n56364, n56365, n56366, n56368, n56369, n56370, n56371, n56372, n56373,
    n56374, n56375, n56376, n56377, n56378, n56379, n56380, n56381, n56382,
    n56383, n56384, n56385, n56386, n56387, n56388, n56389, n56390, n56391,
    n56392, n56393, n56394, n56395, n56396, n56397, n56398, n56400, n56401,
    n56402, n56403, n56404, n56405, n56406, n56407, n56408, n56409, n56410,
    n56411, n56412, n56413, n56414, n56415, n56416, n56417, n56418, n56419,
    n56420, n56421, n56422, n56423, n56424, n56425, n56426, n56427, n56428,
    n56429, n56430, n56431, n56432, n56433, n56434, n56435, n56436, n56437,
    n56438, n56439, n56440, n56441, n56442, n56443, n56444, n56445, n56446,
    n56447, n56448, n56449, n56450, n56451, n56452, n56453, n56454, n56455,
    n56456, n56457, n56458, n56459, n56460, n56461, n56462, n56463, n56464,
    n56465, n56466, n56467, n56468, n56469, n56470, n56471, n56472, n56473,
    n56474, n56475, n56476, n56477, n56478, n56479, n56480, n56481, n56482,
    n56483, n56484, n56485, n56486, n56487, n56488, n56489, n56490, n56491,
    n56492, n56493, n56494, n56495, n56496, n56497, n56498, n56499, n56500,
    n56501, n56502, n56503, n56505, n56506, n56507, n56508, n56509, n56510,
    n56511, n56512, n56513, n56514, n56515, n56516, n56517, n56518, n56519,
    n56520, n56521, n56522, n56523, n56524, n56525, n56526, n56527, n56528,
    n56529, n56530, n56531, n56532, n56533, n56534, n56535, n56536, n56537,
    n56538, n56539, n56540, n56541, n56542, n56543, n56544, n56545, n56546,
    n56547, n56548, n56549, n56550, n56551, n56552, n56554, n56555, n56556,
    n56557, n56558, n56559, n56560, n56561, n56562, n56563, n56564, n56565,
    n56566, n56567, n56568, n56569, n56570, n56571, n56572, n56573, n56574,
    n56575, n56576, n56577, n56578, n56579, n56580, n56581, n56582, n56583,
    n56584, n56585, n56586, n56588, n56589, n56590, n56591, n56592, n56593,
    n56594, n56595, n56596, n56597, n56598, n56599, n56600, n56601, n56602,
    n56603, n56604, n56605, n56606, n56607, n56608, n56609, n56610, n56611,
    n56612, n56613, n56614, n56615, n56616, n56617, n56618, n56619, n56620,
    n56621, n56622, n56623, n56624, n56625, n56626, n56628, n56629, n56630,
    n56631, n56632, n56633, n56634, n56635, n56636, n56637, n56638, n56639,
    n56640, n56641, n56642, n56643, n56644, n56645, n56646, n56647, n56648,
    n56649, n56650, n56651, n56652, n56653, n56654, n56655, n56656, n56657,
    n56658, n56659, n56660, n56661, n56662, n56663, n56664, n56665, n56666,
    n56667, n56668, n56669, n56670, n56671, n56672, n56673, n56674, n56675,
    n56676, n56677, n56678, n56679, n56680, n56681, n56682, n56683, n56684,
    n56685, n56686, n56687, n56688, n56689, n56690, n56691, n56692, n56693,
    n56694, n56695, n56696, n56697, n56698, n56699, n56700, n56701, n56702,
    n56703, n56704, n56705, n56706, n56707, n56708, n56709, n56710, n56711,
    n56712, n56713, n56714, n56715, n56716, n56718, n56719, n56720, n56721,
    n56722, n56723, n56724, n56725, n56726, n56727, n56728, n56729, n56730,
    n56731, n56732, n56733, n56734, n56735, n56736, n56737, n56738, n56739,
    n56740, n56741, n56742, n56743, n56744, n56745, n56746, n56747, n56748,
    n56749, n56750, n56751, n56752, n56753, n56754, n56755, n56756, n56757,
    n56758, n56760, n56761, n56762, n56763, n56764, n56765, n56766, n56767,
    n56768, n56769, n56770, n56771, n56772, n56773, n56774, n56775, n56776,
    n56777, n56778, n56779, n56780, n56781, n56782, n56783, n56784, n56785,
    n56786, n56787, n56788, n56789, n56790, n56791, n56792, n56793, n56794,
    n56795, n56796, n56797, n56798, n56799, n56801, n56802, n56803, n56804,
    n56805, n56806, n56807, n56808, n56809, n56810, n56811, n56812, n56813,
    n56814, n56815, n56816, n56817, n56818, n56819, n56820, n56821, n56822,
    n56823, n56824, n56825, n56826, n56827, n56828, n56829, n56830, n56831,
    n56832, n56833, n56834, n56835, n56836, n56837, n56838, n56839, n56840,
    n56841, n56842, n56843, n56844, n56845, n56846, n56847, n56848, n56849,
    n56850, n56851, n56852, n56853, n56854, n56855, n56856, n56857, n56858,
    n56859, n56860, n56861, n56862, n56863, n56864, n56865, n56866, n56867,
    n56868, n56869, n56870, n56871, n56872, n56873, n56874, n56875, n56876,
    n56877, n56878, n56879, n56880, n56881, n56882, n56883, n56884, n56885,
    n56886, n56887, n56889, n56890, n56891, n56892, n56893, n56894, n56895,
    n56896, n56897, n56898, n56899, n56900, n56901, n56902, n56903, n56904,
    n56905, n56906, n56907, n56908, n56909, n56910, n56911, n56912, n56913,
    n56914, n56915, n56916, n56917, n56918, n56919, n56920, n56921, n56922,
    n56923, n56924, n56925, n56926, n56927, n56928, n56929, n56930, n56931,
    n56932, n56933, n56934, n56935, n56936, n56937, n56939, n56940, n56941,
    n56942, n56943, n56944, n56945, n56946, n56947, n56948, n56949, n56950,
    n56951, n56952, n56953, n56954, n56955, n56956, n56957, n56958, n56959,
    n56960, n56961, n56962, n56963, n56964, n56965, n56966, n56967, n56968,
    n56969, n56970, n56971, n56972, n56973, n56974, n56976, n56977, n56978,
    n56979, n56980, n56981, n56982, n56983, n56984, n56985, n56986, n56987,
    n56988, n56989, n56990, n56991, n56992, n56993, n56994, n56995, n56996,
    n56997, n56998, n56999, n57000, n57001, n57002, n57003, n57004, n57005,
    n57006, n57007, n57008, n57009, n57010, n57011, n57012, n57013, n57014,
    n57015, n57016, n57017, n57018, n57019, n57021, n57022, n57023, n57024,
    n57025, n57026, n57027, n57028, n57029, n57030, n57031, n57032, n57033,
    n57034, n57035, n57036, n57037, n57038, n57039, n57040, n57041, n57042,
    n57043, n57044, n57045, n57046, n57047, n57048, n57049, n57050, n57051,
    n57052, n57053, n57054, n57056, n57057, n57058, n57059, n57060, n57061,
    n57062, n57063, n57064, n57065, n57066, n57067, n57068, n57069, n57070,
    n57071, n57072, n57073, n57074, n57075, n57076, n57077, n57078, n57079,
    n57080, n57081, n57082, n57083, n57084, n57085, n57086, n57087, n57088,
    n57089, n57090, n57091, n57092, n57093, n57094, n57095, n57096, n57097,
    n57098, n57099, n57100, n57101, n57102, n57103, n57104, n57105, n57106,
    n57108, n57109, n57110, n57111, n57112, n57113, n57114, n57115, n57116,
    n57117, n57118, n57119, n57120, n57121, n57122, n57123, n57124, n57125,
    n57126, n57127, n57128, n57129, n57130, n57131, n57132, n57133, n57134,
    n57135, n57136, n57137, n57138, n57139, n57140, n57141, n57142, n57143,
    n57144, n57146, n57147, n57148, n57149, n57150, n57151, n57152, n57153,
    n57154, n57155, n57156, n57157, n57158, n57159, n57160, n57161, n57162,
    n57163, n57164, n57165, n57166, n57167, n57168, n57169, n57170, n57171,
    n57172, n57173, n57174, n57175, n57176, n57177, n57178, n57180, n57181,
    n57182, n57183, n57184, n57185, n57186, n57187, n57188, n57189, n57190,
    n57191, n57192, n57193, n57194, n57195, n57196, n57197, n57198, n57199,
    n57200, n57201, n57202, n57203, n57204, n57205, n57206, n57207, n57208,
    n57209, n57210, n57211, n57212, n57213, n57214, n57215, n57216, n57217,
    n57218, n57220, n57221, n57222, n57223, n57224, n57225, n57226, n57227,
    n57228, n57229, n57230, n57231, n57232, n57233, n57234, n57235, n57236,
    n57237, n57238, n57239, n57240, n57241, n57242, n57243, n57244, n57245,
    n57246, n57247, n57248, n57249, n57250, n57251, n57252, n57253, n57254,
    n57255, n57256, n57257, n57258, n57259, n57260, n57261, n57262, n57263,
    n57264, n57265, n57266, n57267, n57268, n57270, n57271, n57272, n57273,
    n57274, n57275, n57276, n57277, n57278, n57279, n57280, n57281, n57282,
    n57283, n57284, n57285, n57286, n57287, n57288, n57289, n57290, n57291,
    n57292, n57293, n57294, n57295, n57296, n57297, n57298, n57299, n57300,
    n57301, n57302, n57303, n57304, n57305, n57307, n57308, n57309, n57310,
    n57311, n57312, n57313, n57314, n57315, n57316, n57317, n57318, n57319,
    n57320, n57321, n57322, n57323, n57324, n57325, n57326, n57327, n57328,
    n57329, n57330, n57331, n57332, n57333, n57334, n57336, n57337, n57338,
    n57339, n57340, n57341, n57342, n57343, n57344, n57345, n57346, n57347,
    n57348, n57349, n57350, n57351, n57352, n57353, n57354, n57355, n57356,
    n57357, n57358, n57359, n57360, n57361, n57362, n57363, n57364, n57365,
    n57366, n57367, n57368, n57369, n57370, n57371, n57372, n57374, n57375,
    n57376, n57377, n57378, n57379, n57380, n57381, n57382, n57383, n57384,
    n57385, n57386, n57387, n57388, n57389, n57390, n57391, n57392, n57393,
    n57394, n57395, n57396, n57397, n57398, n57399, n57400, n57401, n57402,
    n57403, n57404, n57405, n57406, n57407, n57408, n57409, n57411, n57412,
    n57413, n57414, n57415, n57416, n57417, n57418, n57419, n57420, n57421,
    n57422, n57423, n57424, n57425, n57426, n57427, n57428, n57429, n57430,
    n57431, n57432, n57433, n57434, n57435, n57436, n57437, n57438, n57439,
    n57441, n57442, n57443, n57444, n57445, n57446, n57447, n57448, n57449,
    n57450, n57451, n57452, n57453, n57454, n57455, n57456, n57457, n57458,
    n57459, n57460, n57461, n57462, n57463, n57464, n57465, n57466, n57467,
    n57468, n57469, n57470, n57471, n57472, n57473, n57474, n57475, n57476,
    n57477, n57479, n57480, n57481, n57482, n57483, n57484, n57485, n57486,
    n57487, n57488, n57489, n57490, n57491, n57492, n57493, n57494, n57495,
    n57496, n57497, n57498, n57499, n57500, n57501, n57502, n57503, n57504,
    n57505, n57506, n57507, n57509, n57510, n57511, n57512, n57513, n57514,
    n57515, n57516, n57517, n57518, n57519, n57520, n57521, n57522, n57523,
    n57524, n57525, n57526, n57527, n57528, n57529, n57530, n57531, n57532,
    n57533, n57534, n57535, n57536, n57537, n57538, n57539, n57540, n57542,
    n57543, n57544, n57545, n57546, n57547, n57548, n57549, n57550, n57551,
    n57552, n57553, n57554, n57555, n57556, n57557, n57558, n57559, n57560,
    n57561, n57562, n57563, n57564, n57565, n57566, n57568, n57569, n57570,
    n57571, n57572, n57573, n57574, n57575, n57576, n57577, n57578, n57579,
    n57580, n57581, n57582, n57583, n57584, n57585, n57586, n57587, n57588,
    n57589, n57590, n57591, n57592, n57593, n57594, n57595, n57596, n57597,
    n57598, n57599, n57600, n57601, n57602, n57603, n57604, n57605, n57606,
    n57607, n57608, n57609, n57610, n57611, n57612, n57613, n57614, n57615,
    n57616, n57617, n57618, n57619, n57620, n57621, n57622, n57623, n57624,
    n57625, n57626, n57627, n57628, n57629, n57630, n57631, n57632, n57633,
    n57634, n57635, n57636, n57637, n57638, n57639, n57640, n57641, n57642,
    n57643, n57644, n57645, n57646, n57647, n57648, n57649, n57650, n57651,
    n57652, n57653, n57654, n57655, n57656, n57657, n57658, n57659, n57660,
    n57661, n57662, n57663, n57664, n57665, n57666, n57667, n57668, n57669,
    n57670, n57671, n57673, n57674, n57675, n57676, n57677, n57678, n57679,
    n57680, n57681, n57682, n57683, n57684, n57685, n57686, n57687, n57688,
    n57689, n57690, n57691, n57692, n57693, n57694, n57695, n57696, n57697,
    n57698, n57699, n57700, n57701, n57702, n57703, n57704, n57705, n57706,
    n57707, n57708, n57709, n57710, n57711, n57712, n57713, n57714, n57716,
    n57717, n57718, n57719, n57720, n57721, n57722, n57723, n57724, n57725,
    n57726, n57727, n57728, n57729, n57730, n57731, n57732, n57733, n57734,
    n57735, n57736, n57737, n57738, n57739, n57740, n57741, n57742, n57743,
    n57744, n57745, n57746, n57747, n57748, n57749, n57750, n57751, n57752,
    n57753, n57754, n57755, n57756, n57757, n57758, n57759, n57760, n57761,
    n57762, n57763, n57764, n57765, n57766, n57767, n57768, n57769, n57770,
    n57771, n57772, n57773, n57774, n57775, n57776, n57777, n57778, n57779,
    n57780, n57781, n57782, n57783, n57784, n57785, n57786, n57787, n57788,
    n57789, n57790, n57791, n57792, n57793, n57794, n57795, n57796, n57797,
    n57798, n57799, n57800, n57801, n57802, n57803, n57804, n57805, n57806,
    n57807, n57808, n57809, n57810, n57811, n57812, n57813, n57814, n57815,
    n57816, n57817, n57818, n57820, n57821, n57822, n57823, n57824, n57825,
    n57826, n57827, n57828, n57829, n57830, n57831, n57832, n57833, n57834,
    n57835, n57836, n57837, n57838, n57839, n57840, n57841, n57842, n57843,
    n57844, n57845, n57846, n57847, n57848, n57849, n57850, n57851, n57852,
    n57853, n57854, n57855, n57856, n57857, n57858, n57859, n57860, n57861,
    n57862, n57863, n57864, n57865, n57866, n57867, n57868, n57869, n57870,
    n57871, n57872, n57873, n57874, n57875, n57876, n57877, n57878, n57879,
    n57880, n57881, n57882, n57883, n57884, n57885, n57886, n57887, n57888,
    n57889, n57890, n57891, n57892, n57893, n57894, n57895, n57896, n57897,
    n57898, n57899, n57900, n57901, n57902, n57903, n57904, n57905, n57906,
    n57907, n57908, n57909, n57910, n57911, n57912, n57913, n57914, n57915,
    n57916, n57917, n57918, n57919, n57920, n57921, n57922, n57923, n57924,
    n57925, n57927, n57928, n57929, n57930, n57931, n57932, n57933, n57934,
    n57935, n57936, n57937, n57938, n57939, n57940, n57941, n57942, n57943,
    n57944, n57945, n57946, n57947, n57948, n57949, n57950, n57951, n57952,
    n57953, n57954, n57955, n57956, n57957, n57958, n57959, n57960, n57961,
    n57962, n57963, n57964, n57965, n57966, n57967, n57968, n57969, n57970,
    n57971, n57972, n57973, n57974, n57975, n57976, n57977, n57978, n57979,
    n57980, n57981, n57982, n57983, n57984, n57985, n57986, n57987, n57988,
    n57989, n57990, n57991, n57992, n57993, n57994, n57995, n57996, n57997,
    n57998, n57999, n58000, n58001, n58002, n58003, n58004, n58005, n58006,
    n58007, n58008, n58009, n58010, n58011, n58012, n58013, n58014, n58015,
    n58016, n58017, n58018, n58019, n58020, n58021, n58022, n58023, n58024,
    n58025, n58026, n58027, n58029, n58030, n58031, n58032, n58033, n58034,
    n58035, n58036, n58037, n58038, n58039, n58040, n58041, n58042, n58043,
    n58044, n58045, n58046, n58047, n58048, n58049, n58050, n58051, n58052,
    n58053, n58054, n58055, n58056, n58057, n58058, n58059, n58060, n58061,
    n58062, n58063, n58064, n58065, n58066, n58067, n58068, n58070, n58071,
    n58072, n58073, n58074, n58075, n58076, n58077, n58078, n58079, n58080,
    n58081, n58082, n58083, n58084, n58085, n58086, n58087, n58088, n58089,
    n58090, n58091, n58092, n58093, n58094, n58095, n58096, n58097, n58098,
    n58099, n58100, n58102, n58103, n58104, n58105, n58106, n58107, n58108,
    n58109, n58110, n58111, n58112, n58113, n58114, n58115, n58116, n58117,
    n58118, n58119, n58120, n58121, n58122, n58123, n58124, n58125, n58126,
    n58127, n58128, n58129, n58130, n58131, n58132, n58133, n58134, n58135,
    n58136, n58137, n58138, n58139, n58140, n58141, n58142, n58143, n58144,
    n58145, n58146, n58147, n58148, n58149, n58150, n58151, n58152, n58153,
    n58154, n58155, n58156, n58157, n58158, n58159, n58160, n58161, n58162,
    n58163, n58164, n58165, n58166, n58167, n58168, n58169, n58170, n58171,
    n58172, n58173, n58174, n58175, n58176, n58177, n58178, n58179, n58180,
    n58181, n58182, n58183, n58184, n58185, n58186, n58187, n58188, n58189,
    n58190, n58191, n58192, n58193, n58194, n58195, n58196, n58197, n58198,
    n58200, n58201, n58202, n58203, n58204, n58205, n58206, n58207, n58208,
    n58209, n58210, n58211, n58212, n58213, n58214, n58215, n58216, n58217,
    n58218, n58219, n58220, n58221, n58222, n58223, n58224, n58225, n58226,
    n58227, n58228, n58229, n58230, n58231, n58232, n58233, n58234, n58235,
    n58236, n58237, n58239, n58240, n58241, n58242, n58243, n58244, n58245,
    n58246, n58247, n58248, n58249, n58250, n58251, n58252, n58253, n58254,
    n58255, n58256, n58257, n58258, n58259, n58260, n58261, n58262, n58263,
    n58264, n58265, n58266, n58267, n58268, n58269, n58270, n58271, n58272,
    n58273, n58274, n58275, n58276, n58277, n58278, n58279, n58280, n58281,
    n58282, n58283, n58284, n58285, n58286, n58287, n58288, n58289, n58290,
    n58291, n58292, n58293, n58294, n58295, n58296, n58297, n58298, n58299,
    n58300, n58301, n58302, n58303, n58304, n58305, n58306, n58307, n58308,
    n58309, n58310, n58311, n58312, n58313, n58314, n58315, n58316, n58317,
    n58318, n58319, n58320, n58321, n58322, n58323, n58324, n58325, n58326,
    n58327, n58328, n58329, n58330, n58331, n58332, n58333, n58334, n58335,
    n58336, n58337, n58338, n58339, n58340, n58341, n58342, n58344, n58345,
    n58346, n58347, n58348, n58349, n58350, n58351, n58352, n58353, n58354,
    n58355, n58356, n58357, n58358, n58359, n58360, n58361, n58362, n58363,
    n58364, n58365, n58366, n58367, n58368, n58369, n58370, n58371, n58372,
    n58373, n58374, n58375, n58376, n58377, n58378, n58379, n58380, n58381,
    n58382, n58383, n58385, n58386, n58387, n58388, n58389, n58390, n58391,
    n58392, n58393, n58394, n58395, n58396, n58397, n58398, n58399, n58400,
    n58401, n58402, n58403, n58404, n58405, n58406, n58407, n58408, n58409,
    n58410, n58411, n58412, n58413, n58415, n58416, n58417, n58418, n58419,
    n58420, n58421, n58422, n58423, n58424, n58425, n58426, n58427, n58428,
    n58429, n58430, n58431, n58432, n58433, n58434, n58435, n58436, n58437,
    n58438, n58439, n58440, n58441, n58442, n58443, n58444, n58445, n58446,
    n58447, n58448, n58449, n58450, n58451, n58452, n58453, n58454, n58455,
    n58456, n58457, n58458, n58459, n58460, n58461, n58463, n58464, n58465,
    n58466, n58467, n58468, n58469, n58470, n58471, n58472, n58473, n58474,
    n58475, n58476, n58477, n58478, n58479, n58480, n58481, n58482, n58483,
    n58484, n58485, n58486, n58487, n58488, n58489, n58490, n58491, n58492,
    n58493, n58494, n58495, n58496, n58497, n58498, n58499, n58500, n58501,
    n58502, n58503, n58504, n58505, n58506, n58507, n58508, n58509, n58510,
    n58511, n58512, n58513, n58514, n58515, n58516, n58517, n58518, n58519,
    n58520, n58521, n58522, n58523, n58524, n58525, n58526, n58527, n58528,
    n58529, n58530, n58531, n58532, n58533, n58534, n58535, n58536, n58537,
    n58538, n58539, n58540, n58541, n58542, n58543, n58544, n58545, n58546,
    n58547, n58548, n58549, n58550, n58551, n58552, n58553, n58554, n58555,
    n58556, n58557, n58559, n58560, n58561, n58562, n58563, n58564, n58565,
    n58566, n58567, n58568, n58569, n58570, n58571, n58572, n58573, n58574,
    n58575, n58576, n58577, n58578, n58579, n58580, n58581, n58582, n58583,
    n58584, n58585, n58586, n58587, n58588, n58589, n58590, n58591, n58592,
    n58593, n58595, n58596, n58597, n58598, n58599, n58600, n58601, n58602,
    n58603, n58604, n58605, n58606, n58607, n58608, n58609, n58610, n58611,
    n58612, n58613, n58614, n58615, n58616, n58617, n58618, n58619, n58620,
    n58621, n58622, n58623, n58624, n58625, n58626, n58628, n58629, n58630,
    n58631, n58632, n58633, n58634, n58635, n58636, n58637, n58638, n58639,
    n58640, n58641, n58642, n58643, n58644, n58645, n58646, n58647, n58648,
    n58649, n58650, n58651, n58652, n58653, n58654, n58655, n58656, n58657,
    n58658, n58659, n58660, n58661, n58662, n58663, n58664, n58665, n58666,
    n58667, n58668, n58669, n58670, n58671, n58672, n58673, n58675, n58676,
    n58677, n58678, n58679, n58680, n58681, n58682, n58683, n58684, n58685,
    n58686, n58687, n58688, n58689, n58690, n58691, n58692, n58693, n58694,
    n58695, n58696, n58697, n58698, n58699, n58700, n58701, n58702, n58703,
    n58704, n58705, n58706, n58707, n58708, n58709, n58710, n58711, n58712,
    n58713, n58714, n58715, n58716, n58717, n58718, n58720, n58721, n58722,
    n58723, n58724, n58725, n58726, n58727, n58728, n58729, n58730, n58731,
    n58732, n58733, n58734, n58735, n58736, n58737, n58738, n58739, n58740,
    n58741, n58742, n58743, n58744, n58745, n58746, n58747, n58748, n58749,
    n58750, n58751, n58752, n58753, n58754, n58755, n58756, n58757, n58758,
    n58760, n58761, n58762, n58763, n58764, n58765, n58766, n58767, n58768,
    n58769, n58770, n58771, n58772, n58773, n58774, n58775, n58776, n58777,
    n58778, n58779, n58780, n58781, n58782, n58783, n58784, n58785, n58786,
    n58787, n58788, n58789, n58790, n58791, n58792, n58793, n58794, n58795,
    n58796, n58797, n58799, n58800, n58801, n58802, n58803, n58804, n58805,
    n58806, n58807, n58808, n58809, n58810, n58811, n58812, n58813, n58814,
    n58815, n58816, n58817, n58818, n58819, n58820, n58821, n58822, n58823,
    n58824, n58825, n58826, n58827, n58828, n58829, n58830, n58831, n58833,
    n58834, n58835, n58836, n58837, n58838, n58839, n58840, n58841, n58842,
    n58843, n58844, n58845, n58846, n58847, n58848, n58849, n58850, n58851,
    n58852, n58853, n58854, n58855, n58856, n58857, n58858, n58859, n58860,
    n58861, n58862, n58863, n58864, n58865, n58866, n58867, n58868, n58869,
    n58870, n58871, n58872, n58873, n58874, n58875, n58876, n58878, n58879,
    n58880, n58881, n58882, n58883, n58884, n58885, n58886, n58887, n58888,
    n58889, n58890, n58891, n58892, n58893, n58894, n58895, n58896, n58897,
    n58898, n58899, n58900, n58901, n58902, n58903, n58904, n58905, n58906,
    n58907, n58908, n58909, n58910, n58911, n58912, n58913, n58914, n58915,
    n58917, n58918, n58919, n58920, n58921, n58922, n58923, n58924, n58925,
    n58926, n58927, n58928, n58929, n58930, n58931, n58932, n58933, n58934,
    n58935, n58936, n58937, n58938, n58939, n58940, n58941, n58942, n58943,
    n58944, n58945, n58946, n58947, n58948, n58949, n58950, n58951, n58952,
    n58953, n58954, n58955, n58956, n58957, n58958, n58959, n58960, n58961,
    n58962, n58963, n58964, n58965, n58966, n58967, n58968, n58969, n58970,
    n58971, n58972, n58973, n58974, n58975, n58976, n58977, n58978, n58979,
    n58980, n58981, n58982, n58983, n58984, n58985, n58986, n58987, n58988,
    n58989, n58990, n58991, n58992, n58993, n58994, n58995, n58996, n58997,
    n58998, n58999, n59000, n59001, n59002, n59003, n59004, n59005, n59006,
    n59007, n59008, n59009, n59010, n59011, n59013, n59014, n59015, n59016,
    n59017, n59018, n59019, n59020, n59021, n59022, n59023, n59024, n59025,
    n59026, n59027, n59028, n59029, n59030, n59031, n59032, n59033, n59034,
    n59035, n59036, n59037, n59038, n59039, n59040, n59041, n59042, n59043,
    n59044, n59045, n59046, n59047, n59048, n59049, n59050, n59051, n59052,
    n59053, n59054, n59055, n59056, n59057, n59059, n59060, n59061, n59062,
    n59063, n59064, n59065, n59066, n59067, n59068, n59069, n59070, n59071,
    n59072, n59073, n59074, n59075, n59076, n59077, n59078, n59079, n59080,
    n59081, n59082, n59083, n59084, n59085, n59086, n59087, n59088, n59089,
    n59090, n59091, n59092, n59094, n59095, n59096, n59097, n59098, n59099,
    n59100, n59101, n59102, n59103, n59104, n59105, n59106, n59107, n59108,
    n59109, n59110, n59111, n59112, n59113, n59114, n59115, n59116, n59117,
    n59118, n59119, n59120, n59121, n59122, n59123, n59124, n59125, n59126,
    n59127, n59128, n59130, n59131, n59132, n59133, n59134, n59135, n59136,
    n59137, n59138, n59139, n59140, n59141, n59142, n59143, n59144, n59145,
    n59146, n59147, n59148, n59149, n59150, n59151, n59152, n59153, n59154,
    n59155, n59156, n59157, n59158, n59160, n59161, n59162, n59163, n59164,
    n59165, n59166, n59167, n59168, n59169, n59170, n59171, n59172, n59173,
    n59174, n59175, n59176, n59177, n59178, n59179, n59180, n59181, n59182,
    n59183, n59184, n59185, n59186, n59187, n59188, n59189, n59190, n59191,
    n59192, n59193, n59194, n59195, n59197, n59198, n59199, n59200, n59201,
    n59202, n59203, n59204, n59205, n59206, n59207, n59208, n59209, n59210,
    n59211, n59212, n59213, n59214, n59215, n59216, n59217, n59218, n59219,
    n59220, n59221, n59222, n59223, n59224, n59225, n59226, n59227, n59228,
    n59229, n59230, n59231, n59233, n59234, n59235, n59236, n59237, n59238,
    n59239, n59240, n59241, n59242, n59243, n59244, n59245, n59246, n59247,
    n59248, n59249, n59250, n59251, n59252, n59253, n59254, n59255, n59256,
    n59257, n59258, n59259, n59260, n59261, n59262, n59263, n59264, n59265,
    n59267, n59268, n59269, n59270, n59271, n59272, n59273, n59274, n59275,
    n59276, n59277, n59278, n59279, n59280, n59281, n59282, n59283, n59284,
    n59285, n59286, n59287, n59288, n59289, n59290, n59291, n59293, n59294,
    n59295, n59296, n59297, n59298, n59299, n59300, n59301, n59302, n59303,
    n59304, n59305, n59306, n59307, n59308, n59309, n59310, n59311, n59312,
    n59313, n59314, n59315, n59316, n59317, n59318, n59319, n59320, n59321,
    n59322, n59323, n59324, n59325, n59326, n59327, n59328, n59329, n59330,
    n59331, n59332, n59333, n59334, n59335, n59336, n59337, n59338, n59339,
    n59340, n59341, n59342, n59343, n59344, n59345, n59346, n59347, n59348,
    n59349, n59350, n59351, n59352, n59353, n59354, n59355, n59356, n59357,
    n59358, n59359, n59360, n59361, n59362, n59363, n59364, n59365, n59366,
    n59367, n59368, n59369, n59370, n59371, n59372, n59373, n59374, n59375,
    n59376, n59377, n59378, n59379, n59380, n59381, n59382, n59383, n59384,
    n59385, n59386, n59387, n59388, n59389, n59390, n59391, n59392, n59394,
    n59395, n59396, n59397, n59398, n59399, n59400, n59401, n59402, n59403,
    n59404, n59405, n59406, n59407, n59408, n59409, n59410, n59411, n59412,
    n59413, n59414, n59415, n59416, n59417, n59418, n59419, n59420, n59421,
    n59422, n59423, n59424, n59425, n59426, n59427, n59428, n59429, n59430,
    n59431, n59432, n59433, n59434, n59435, n59436, n59437, n59438, n59439,
    n59440, n59441, n59442, n59443, n59444, n59445, n59446, n59447, n59448,
    n59449, n59450, n59451, n59452, n59453, n59454, n59455, n59456, n59457,
    n59458, n59459, n59460, n59461, n59462, n59463, n59464, n59465, n59466,
    n59467, n59468, n59469, n59470, n59471, n59472, n59473, n59474, n59475,
    n59476, n59477, n59478, n59479, n59480, n59481, n59482, n59483, n59484,
    n59485, n59486, n59487, n59488, n59489, n59490, n59491, n59492, n59494,
    n59495, n59496, n59497, n59498, n59499, n59500, n59501, n59502, n59503,
    n59504, n59505, n59506, n59507, n59508, n59509, n59510, n59511, n59512,
    n59513, n59514, n59515, n59516, n59517, n59518, n59519, n59520, n59521,
    n59522, n59523, n59524, n59525, n59526, n59527, n59528, n59529, n59530,
    n59531, n59532, n59533, n59534, n59535, n59536, n59537, n59538, n59539,
    n59540, n59541, n59542, n59543, n59544, n59545, n59546, n59547, n59548,
    n59549, n59550, n59551, n59552, n59553, n59554, n59555, n59556, n59557,
    n59558, n59559, n59560, n59561, n59562, n59563, n59564, n59565, n59566,
    n59567, n59568, n59569, n59570, n59571, n59572, n59573, n59574, n59575,
    n59576, n59577, n59578, n59579, n59580, n59581, n59582, n59583, n59584,
    n59585, n59586, n59587, n59588, n59589, n59590, n59591, n59592, n59593,
    n59595, n59596, n59597, n59598, n59599, n59600, n59601, n59602, n59603,
    n59604, n59605, n59606, n59607, n59608, n59609, n59610, n59611, n59612,
    n59613, n59614, n59615, n59616, n59617, n59618, n59619, n59620, n59621,
    n59622, n59623, n59624, n59625, n59626, n59627, n59628, n59629, n59630,
    n59631, n59632, n59633, n59634, n59635, n59636, n59637, n59638, n59639,
    n59640, n59641, n59642, n59643, n59644, n59645, n59646, n59647, n59648,
    n59649, n59650, n59651, n59652, n59653, n59654, n59655, n59656, n59657,
    n59658, n59659, n59660, n59661, n59662, n59663, n59664, n59665, n59666,
    n59667, n59668, n59669, n59670, n59671, n59672, n59673, n59674, n59675,
    n59676, n59677, n59678, n59679, n59680, n59681, n59682, n59683, n59684,
    n59685, n59686, n59687, n59688, n59689, n59690, n59691, n59692, n59693,
    n59694, n59695, n59696, n59697, n59698, n59700, n59701, n59702, n59703,
    n59704, n59705, n59706, n59707, n59708, n59709, n59710, n59711, n59712,
    n59713, n59714, n59715, n59716, n59717, n59718, n59719, n59720, n59721,
    n59722, n59723, n59724, n59725, n59726, n59727, n59728, n59729, n59730,
    n59731, n59732, n59733, n59734, n59735, n59736, n59737, n59738, n59739,
    n59740, n59741, n59742, n59743, n59744, n59745, n59746, n59747, n59748,
    n59749, n59750, n59751, n59752, n59753, n59754, n59755, n59756, n59757,
    n59758, n59759, n59760, n59761, n59762, n59763, n59764, n59765, n59766,
    n59767, n59768, n59769, n59770, n59771, n59772, n59773, n59774, n59775,
    n59776, n59777, n59778, n59779, n59780, n59781, n59782, n59783, n59784,
    n59785, n59786, n59787, n59788, n59790, n59791, n59792, n59793, n59794,
    n59795, n59796, n59797, n59798, n59799, n59800, n59801, n59802, n59803,
    n59804, n59805, n59806, n59807, n59808, n59809, n59810, n59811, n59812,
    n59813, n59814, n59815, n59816, n59817, n59818, n59819, n59820, n59821,
    n59822, n59823, n59824, n59825, n59826, n59827, n59828, n59829, n59830,
    n59831, n59832, n59833, n59834, n59835, n59836, n59837, n59838, n59839,
    n59840, n59841, n59842, n59843, n59844, n59845, n59846, n59847, n59848,
    n59849, n59850, n59851, n59852, n59853, n59854, n59855, n59856, n59857,
    n59858, n59859, n59860, n59861, n59862, n59863, n59864, n59865, n59866,
    n59867, n59868, n59869, n59870, n59871, n59872, n59873, n59874, n59875,
    n59876, n59877, n59878, n59879, n59880, n59881, n59882, n59883, n59884,
    n59885, n59886, n59887, n59888, n59889, n59890, n59891, n59892, n59893,
    n59894, n59896, n59897, n59898, n59899, n59900, n59901, n59902, n59903,
    n59904, n59905, n59906, n59907, n59908, n59909, n59910, n59911, n59912,
    n59913, n59914, n59915, n59916, n59917, n59918, n59919, n59920, n59921,
    n59922, n59923, n59924, n59925, n59926, n59927, n59928, n59929, n59930,
    n59931, n59932, n59933, n59934, n59935, n59936, n59937, n59938, n59939,
    n59940, n59941, n59942, n59943, n59944, n59945, n59946, n59947, n59948,
    n59949, n59950, n59951, n59952, n59953, n59954, n59955, n59956, n59957,
    n59958, n59959, n59960, n59961, n59962, n59963, n59964, n59965, n59966,
    n59967, n59968, n59969, n59970, n59971, n59972, n59973, n59974, n59975,
    n59976, n59977, n59978, n59979, n59980, n59981, n59982, n59983, n59984,
    n59985, n59986, n59987, n59988, n59989, n59990, n59991, n59992, n59993,
    n59994, n59995, n59996, n59997, n59998, n59999, n60001, n60002, n60003,
    n60004, n60005, n60006, n60007, n60008, n60009, n60010, n60011, n60012,
    n60013, n60014, n60015, n60016, n60017, n60018, n60019, n60020, n60021,
    n60022, n60023, n60024, n60025, n60026, n60027, n60028, n60029, n60030,
    n60031, n60032, n60033, n60034, n60035, n60036, n60037, n60038, n60039,
    n60040, n60042, n60043, n60044, n60045, n60046, n60047, n60048, n60049,
    n60050, n60051, n60052, n60053, n60054, n60055, n60056, n60057, n60058,
    n60059, n60060, n60061, n60062, n60063, n60064, n60065, n60066, n60067,
    n60068, n60069, n60070, n60071, n60072, n60073, n60074, n60075, n60076,
    n60077, n60078, n60079, n60080, n60081, n60082, n60083, n60084, n60085,
    n60086, n60087, n60088, n60089, n60090, n60092, n60093, n60094, n60095,
    n60096, n60097, n60098, n60099, n60100, n60101, n60102, n60103, n60104,
    n60105, n60106, n60107, n60108, n60109, n60110, n60111, n60112, n60113,
    n60114, n60115, n60116, n60117, n60118, n60119, n60120, n60121, n60122,
    n60123, n60124, n60125, n60126, n60127, n60128, n60129, n60130, n60131,
    n60132, n60134, n60135, n60136, n60137, n60138, n60139, n60140, n60141,
    n60142, n60143, n60144, n60145, n60146, n60147, n60148, n60149, n60150,
    n60151, n60152, n60153, n60154, n60155, n60156, n60157, n60158, n60159,
    n60160, n60161, n60162, n60163, n60164, n60165, n60166, n60167, n60168,
    n60169, n60170, n60171, n60173, n60174, n60175, n60176, n60177, n60178,
    n60179, n60180, n60181, n60182, n60183, n60184, n60185, n60186, n60187,
    n60188, n60189, n60190, n60191, n60192, n60193, n60194, n60195, n60196,
    n60197, n60198, n60199, n60200, n60201, n60202, n60203, n60204, n60205,
    n60206, n60207, n60208, n60209, n60210, n60211, n60212, n60214, n60215,
    n60216, n60217, n60218, n60219, n60220, n60221, n60222, n60223, n60224,
    n60225, n60226, n60227, n60228, n60229, n60230, n60231, n60232, n60233,
    n60234, n60235, n60236, n60237, n60238, n60239, n60240, n60241, n60242,
    n60243, n60244, n60245, n60246, n60247, n60248, n60249, n60250, n60251,
    n60252, n60253, n60254, n60255, n60256, n60257, n60258, n60259, n60260,
    n60261, n60262, n60263, n60264, n60265, n60266, n60267, n60268, n60269,
    n60270, n60271, n60272, n60273, n60274, n60275, n60276, n60277, n60278,
    n60279, n60280, n60281, n60282, n60283, n60284, n60285, n60286, n60287,
    n60288, n60289, n60290, n60291, n60292, n60293, n60294, n60295, n60296,
    n60297, n60298, n60299, n60300, n60301, n60302, n60303, n60304, n60305,
    n60306, n60307, n60308, n60309, n60311, n60312, n60313, n60314, n60315,
    n60316, n60317, n60318, n60319, n60320, n60321, n60322, n60323, n60324,
    n60325, n60326, n60327, n60328, n60329, n60330, n60331, n60332, n60333,
    n60334, n60335, n60336, n60337, n60338, n60339, n60340, n60341, n60342,
    n60343, n60344, n60345, n60346, n60347, n60348, n60349, n60350, n60351,
    n60352, n60353, n60354, n60355, n60356, n60357, n60358, n60360, n60361,
    n60362, n60363, n60364, n60365, n60366, n60367, n60368, n60369, n60370,
    n60371, n60372, n60373, n60374, n60375, n60376, n60377, n60378, n60379,
    n60380, n60381, n60382, n60383, n60384, n60385, n60386, n60387, n60388,
    n60389, n60390, n60391, n60392, n60394, n60395, n60396, n60397, n60398,
    n60399, n60400, n60401, n60402, n60403, n60404, n60405, n60406, n60407,
    n60408, n60409, n60410, n60411, n60412, n60413, n60414, n60415, n60416,
    n60417, n60418, n60419, n60420, n60421, n60422, n60423, n60424, n60425,
    n60427, n60428, n60429, n60430, n60431, n60432, n60433, n60434, n60435,
    n60436, n60437, n60438, n60439, n60440, n60441, n60442, n60443, n60444,
    n60445, n60446, n60447, n60448, n60449, n60450, n60451, n60452, n60453,
    n60454, n60455, n60456, n60457, n60458, n60459, n60460, n60461, n60462,
    n60463, n60464, n60465, n60466, n60467, n60468, n60469, n60470, n60472,
    n60473, n60474, n60475, n60476, n60477, n60478, n60479, n60480, n60481,
    n60482, n60483, n60484, n60485, n60486, n60487, n60488, n60489, n60490,
    n60491, n60492, n60493, n60494, n60495, n60496, n60497, n60498, n60499,
    n60500, n60501, n60502, n60503, n60504, n60505, n60506, n60507, n60508,
    n60509, n60510, n60511, n60512, n60513, n60514, n60515, n60517, n60518,
    n60519, n60520, n60521, n60522, n60523, n60524, n60525, n60526, n60527,
    n60528, n60529, n60530, n60531, n60532, n60533, n60534, n60535, n60536,
    n60537, n60538, n60539, n60540, n60541, n60542, n60543, n60544, n60545,
    n60546, n60547, n60548, n60549, n60551, n60552, n60553, n60554, n60555,
    n60556, n60557, n60558, n60559, n60560, n60561, n60562, n60563, n60564,
    n60565, n60566, n60567, n60568, n60569, n60570, n60571, n60572, n60573,
    n60574, n60575, n60576, n60577, n60578, n60579, n60581, n60582, n60583,
    n60584, n60585, n60586, n60587, n60588, n60589, n60590, n60591, n60592,
    n60593, n60594, n60595, n60596, n60597, n60598, n60599, n60600, n60601,
    n60602, n60603, n60604, n60605, n60606, n60607, n60608, n60609, n60610,
    n60611, n60612, n60613, n60614, n60616, n60617, n60618, n60619, n60620,
    n60621, n60622, n60623, n60624, n60625, n60626, n60627, n60628, n60629,
    n60630, n60631, n60632, n60633, n60634, n60635, n60636, n60637, n60638,
    n60639, n60640, n60641, n60642, n60643, n60644, n60645, n60646, n60647,
    n60648, n60649, n60650, n60651, n60652, n60653, n60654, n60655, n60656,
    n60657, n60658, n60659, n60660, n60661, n60663, n60664, n60665, n60666,
    n60667, n60668, n60669, n60670, n60671, n60672, n60673, n60674, n60675,
    n60676, n60677, n60678, n60679, n60680, n60681, n60682, n60683, n60684,
    n60685, n60686, n60687, n60688, n60689, n60690, n60691, n60692, n60693,
    n60694, n60695, n60696, n60697, n60698, n60700, n60701, n60702, n60703,
    n60704, n60705, n60706, n60707, n60708, n60709, n60710, n60711, n60712,
    n60713, n60714, n60715, n60716, n60717, n60718, n60719, n60720, n60721,
    n60722, n60723, n60724, n60725, n60726, n60727, n60729, n60730, n60731,
    n60732, n60733, n60734, n60735, n60736, n60737, n60738, n60739, n60740,
    n60741, n60742, n60743, n60744, n60745, n60746, n60747, n60748, n60749,
    n60750, n60751, n60752, n60753, n60754, n60755, n60756, n60757, n60758,
    n60759, n60760, n60761, n60762, n60763, n60764, n60765, n60767, n60768,
    n60769, n60770, n60771, n60772, n60773, n60774, n60775, n60776, n60777,
    n60778, n60779, n60780, n60781, n60782, n60783, n60784, n60785, n60786,
    n60787, n60788, n60789, n60790, n60791, n60792, n60793, n60794, n60795,
    n60796, n60797, n60798, n60799, n60800, n60801, n60802, n60803, n60805,
    n60806, n60807, n60808, n60809, n60810, n60811, n60812, n60813, n60814,
    n60815, n60816, n60817, n60818, n60819, n60820, n60821, n60822, n60823,
    n60824, n60825, n60826, n60827, n60828, n60829, n60830, n60831, n60832,
    n60833, n60834, n60835, n60836, n60837, n60838, n60839, n60840, n60841,
    n60842, n60843, n60845, n60846, n60847, n60848, n60849, n60850, n60851,
    n60852, n60853, n60854, n60855, n60856, n60857, n60858, n60859, n60860,
    n60861, n60862, n60863, n60864, n60865, n60866, n60867, n60868, n60869,
    n60870, n60871, n60872, n60873, n60874, n60875, n60876, n60877, n60878,
    n60880, n60881, n60882, n60883, n60884, n60885, n60886, n60887, n60888,
    n60889, n60890, n60891, n60892, n60893, n60894, n60895, n60896, n60897,
    n60898, n60899, n60900, n60901, n60902, n60903, n60904, n60905, n60906,
    n60907, n60908, n60909, n60910, n60911, n60912, n60913, n60914, n60915,
    n60917, n60918, n60919, n60920, n60921, n60922, n60923, n60924, n60925,
    n60926, n60927, n60928, n60929, n60930, n60931, n60932, n60933, n60934,
    n60935, n60936, n60937, n60938, n60939, n60940, n60941, n60942, n60943,
    n60944, n60945, n60947, n60948, n60949, n60950, n60951, n60952, n60953,
    n60954, n60955, n60956, n60957, n60958, n60959, n60960, n60961, n60962,
    n60963, n60964, n60965, n60966, n60967, n60968, n60969, n60970, n60971,
    n60972, n60974, n60975, n60976, n60977, n60978, n60979, n60980, n60981,
    n60982, n60983, n60984, n60985, n60986, n60987, n60988, n60989, n60990,
    n60991, n60992, n60993, n60994, n60995, n60996, n60997, n60998, n60999,
    n61000, n61001, n61002, n61003, n61004, n61005, n61006, n61008, n61009,
    n61010, n61011, n61012, n61013, n61014, n61015, n61016, n61017, n61018,
    n61019, n61020, n61021, n61022, n61023, n61024, n61025, n61026, n61027,
    n61028, n61029, n61030, n61031, n61032, n61033, n61034, n61035, n61036,
    n61037, n61038, n61039, n61040, n61041, n61042, n61043, n61044, n61045,
    n61046, n61047, n61048, n61049, n61050, n61051, n61052, n61053, n61054,
    n61055, n61056, n61057, n61058, n61059, n61060, n61061, n61062, n61063,
    n61064, n61065, n61066, n61067, n61068, n61069, n61070, n61071, n61072,
    n61073, n61074, n61075, n61076, n61077, n61078, n61079, n61080, n61081,
    n61082, n61083, n61084, n61085, n61086, n61087, n61088, n61089, n61090,
    n61091, n61092, n61093, n61094, n61095, n61096, n61097, n61098, n61099,
    n61100, n61101, n61102, n61103, n61104, n61105, n61107, n61108, n61109,
    n61110, n61111, n61112, n61113, n61114, n61115, n61116, n61117, n61118,
    n61119, n61120, n61121, n61122, n61123, n61124, n61125, n61126, n61127,
    n61128, n61129, n61130, n61131, n61132, n61133, n61134, n61135, n61136,
    n61137, n61138, n61139, n61140, n61141, n61142, n61143, n61144, n61145,
    n61146, n61147, n61148, n61149, n61150, n61151, n61152, n61153, n61154,
    n61155, n61156, n61157, n61158, n61159, n61160, n61161, n61162, n61163,
    n61164, n61165, n61166, n61167, n61168, n61169, n61170, n61171, n61172,
    n61173, n61174, n61175, n61176, n61177, n61178, n61179, n61180, n61181,
    n61182, n61183, n61184, n61185, n61186, n61187, n61188, n61189, n61190,
    n61191, n61192, n61193, n61194, n61195, n61196, n61197, n61198, n61199,
    n61200, n61201, n61202, n61203, n61204, n61205, n61206, n61207, n61208,
    n61209, n61210, n61211, n61212, n61214, n61215, n61216, n61217, n61218,
    n61219, n61220, n61221, n61222, n61223, n61224, n61225, n61226, n61227,
    n61228, n61229, n61230, n61231, n61232, n61233, n61234, n61235, n61236,
    n61237, n61238, n61239, n61240, n61241, n61242, n61243, n61244, n61245,
    n61246, n61247, n61248, n61249, n61250, n61251, n61252, n61253, n61255,
    n61256, n61257, n61258, n61259, n61260, n61261, n61262, n61263, n61264,
    n61265, n61266, n61267, n61268, n61269, n61270, n61271, n61272, n61273,
    n61274, n61275, n61276, n61277, n61278, n61279, n61280, n61281, n61282,
    n61283, n61284, n61285, n61286, n61287, n61288, n61289, n61290, n61291,
    n61292, n61293, n61294, n61295, n61296, n61297, n61298, n61299, n61300,
    n61301, n61302, n61303, n61304, n61305, n61306, n61307, n61308, n61309,
    n61310, n61311, n61312, n61313, n61314, n61315, n61316, n61317, n61318,
    n61319, n61320, n61321, n61322, n61323, n61324, n61325, n61326, n61327,
    n61328, n61329, n61330, n61331, n61332, n61333, n61334, n61335, n61336,
    n61337, n61338, n61339, n61340, n61341, n61342, n61343, n61344, n61345,
    n61346, n61347, n61348, n61349, n61350, n61352, n61353, n61354, n61355,
    n61356, n61357, n61358, n61359, n61360, n61361, n61362, n61363, n61364,
    n61365, n61366, n61367, n61368, n61369, n61370, n61371, n61372, n61373,
    n61374, n61375, n61376, n61377, n61378, n61379, n61380, n61381, n61382,
    n61383, n61384, n61385, n61386, n61387, n61388, n61389, n61390, n61391,
    n61392, n61393, n61394, n61395, n61396, n61397, n61398, n61399, n61400,
    n61401, n61402, n61403, n61404, n61405, n61406, n61407, n61408, n61409,
    n61410, n61411, n61412, n61413, n61414, n61415, n61416, n61417, n61418,
    n61419, n61420, n61421, n61422, n61423, n61424, n61425, n61426, n61427,
    n61428, n61429, n61430, n61431, n61432, n61433, n61434, n61435, n61436,
    n61437, n61438, n61439, n61440, n61441, n61442, n61443, n61444, n61445,
    n61447, n61448, n61449, n61450, n61451, n61452, n61453, n61454, n61455,
    n61456, n61457, n61458, n61459, n61460, n61461, n61462, n61463, n61464,
    n61465, n61466, n61467, n61468, n61469, n61470, n61471, n61472, n61473,
    n61474, n61475, n61476, n61477, n61478, n61479, n61480, n61481, n61482,
    n61483, n61484, n61485, n61486, n61487, n61488, n61489, n61490, n61491,
    n61492, n61493, n61494, n61496, n61497, n61498, n61499, n61500, n61501,
    n61502, n61503, n61504, n61505, n61506, n61507, n61508, n61509, n61510,
    n61511, n61512, n61513, n61514, n61515, n61516, n61517, n61518, n61519,
    n61520, n61521, n61522, n61523, n61524, n61525, n61526, n61527, n61528,
    n61529, n61530, n61531, n61532, n61533, n61534, n61535, n61536, n61537,
    n61539, n61540, n61541, n61542, n61543, n61544, n61545, n61546, n61547,
    n61548, n61549, n61550, n61551, n61552, n61553, n61554, n61555, n61556,
    n61557, n61558, n61559, n61560, n61561, n61562, n61563, n61564, n61565,
    n61566, n61567, n61568, n61569, n61570, n61571, n61572, n61573, n61574,
    n61575, n61576, n61577, n61578, n61579, n61580, n61581, n61582, n61584,
    n61585, n61586, n61587, n61588, n61589, n61590, n61591, n61592, n61593,
    n61594, n61595, n61596, n61597, n61598, n61599, n61600, n61601, n61602,
    n61603, n61604, n61605, n61606, n61607, n61608, n61609, n61610, n61611,
    n61612, n61613, n61614, n61615, n61616, n61617, n61618, n61619, n61620,
    n61621, n61622, n61623, n61624, n61625, n61626, n61627, n61628, n61629,
    n61630, n61631, n61632, n61633, n61634, n61635, n61636, n61637, n61638,
    n61639, n61640, n61641, n61642, n61643, n61644, n61645, n61646, n61647,
    n61648, n61649, n61650, n61651, n61652, n61653, n61654, n61655, n61656,
    n61657, n61658, n61659, n61660, n61661, n61662, n61663, n61664, n61665,
    n61666, n61667, n61668, n61669, n61670, n61671, n61672, n61673, n61674,
    n61675, n61676, n61677, n61678, n61679, n61680, n61681, n61682, n61683,
    n61684, n61686, n61687, n61688, n61689, n61690, n61691, n61692, n61693,
    n61694, n61695, n61696, n61697, n61698, n61699, n61700, n61701, n61702,
    n61703, n61704, n61705, n61706, n61707, n61708, n61709, n61710, n61711,
    n61712, n61713, n61714, n61715, n61716, n61717, n61718, n61719, n61720,
    n61721, n61722, n61723, n61724, n61725, n61726, n61727, n61728, n61729,
    n61730, n61731, n61732, n61733, n61734, n61735, n61736, n61737, n61738,
    n61739, n61740, n61741, n61742, n61743, n61744, n61745, n61746, n61747,
    n61748, n61749, n61750, n61751, n61752, n61753, n61754, n61755, n61756,
    n61757, n61758, n61759, n61760, n61761, n61762, n61763, n61764, n61765,
    n61766, n61767, n61768, n61769, n61770, n61771, n61772, n61773, n61774,
    n61775, n61776, n61777, n61778, n61779, n61780, n61781, n61782, n61783,
    n61785, n61786, n61787, n61788, n61789, n61790, n61791, n61792, n61793,
    n61794, n61795, n61796, n61797, n61798, n61799, n61800, n61801, n61802,
    n61803, n61804, n61805, n61806, n61807, n61808, n61809, n61810, n61811,
    n61812, n61813, n61814, n61815, n61816, n61817, n61818, n61819, n61820,
    n61821, n61823, n61824, n61825, n61826, n61827, n61828, n61829, n61830,
    n61831, n61832, n61833, n61834, n61835, n61836, n61837, n61838, n61839,
    n61840, n61841, n61842, n61843, n61844, n61845, n61846, n61847, n61848,
    n61849, n61850, n61851, n61852, n61853, n61854, n61855, n61856, n61857,
    n61858, n61859, n61860, n61861, n61862, n61863, n61864, n61865, n61866,
    n61867, n61868, n61869, n61870, n61871, n61872, n61873, n61874, n61875,
    n61876, n61877, n61878, n61879, n61880, n61881, n61882, n61883, n61884,
    n61885, n61886, n61887, n61888, n61889, n61890, n61891, n61892, n61893,
    n61894, n61895, n61896, n61897, n61898, n61899, n61900, n61901, n61902,
    n61903, n61904, n61905, n61906, n61907, n61908, n61909, n61910, n61911,
    n61912, n61913, n61914, n61915, n61916, n61917, n61918, n61919, n61920,
    n61921, n61922, n61923, n61925, n61926, n61927, n61928, n61929, n61930,
    n61931, n61932, n61933, n61934, n61935, n61936, n61937, n61938, n61939,
    n61940, n61941, n61942, n61943, n61944, n61945, n61946, n61947, n61948,
    n61949, n61950, n61951, n61952, n61953, n61955, n61956, n61957, n61958,
    n61959, n61960, n61961, n61962, n61963, n61964, n61965, n61966, n61967,
    n61968, n61969, n61970, n61971, n61972, n61973, n61974, n61975, n61976,
    n61977, n61978, n61979, n61980, n61981, n61982, n61983, n61984, n61985,
    n61986, n61987, n61988, n61989, n61990, n61991, n61992, n61993, n61994,
    n61995, n61996, n61997, n61998, n61999, n62000, n62001, n62003, n62004,
    n62005, n62006, n62007, n62008, n62009, n62010, n62011, n62012, n62013,
    n62014, n62015, n62016, n62017, n62018, n62019, n62020, n62021, n62022,
    n62023, n62024, n62025, n62026, n62027, n62028, n62029, n62030, n62031,
    n62032, n62033, n62034, n62035, n62036, n62037, n62038, n62039, n62040,
    n62041, n62042, n62043, n62044, n62045, n62046, n62047, n62048, n62049,
    n62050, n62052, n62053, n62054, n62055, n62056, n62057, n62058, n62059,
    n62060, n62061, n62062, n62063, n62064, n62065, n62066, n62067, n62068,
    n62069, n62070, n62071, n62072, n62073, n62074, n62075, n62076, n62077,
    n62078, n62079, n62080, n62081, n62082, n62083, n62085, n62086, n62087,
    n62088, n62089, n62090, n62091, n62092, n62093, n62094, n62095, n62096,
    n62097, n62098, n62099, n62100, n62101, n62102, n62103, n62104, n62105,
    n62106, n62107, n62108, n62109, n62110, n62111, n62112, n62113, n62114,
    n62115, n62116, n62117, n62118, n62119, n62120, n62121, n62122, n62124,
    n62125, n62126, n62127, n62128, n62129, n62130, n62131, n62132, n62133,
    n62134, n62135, n62136, n62137, n62138, n62139, n62140, n62141, n62142,
    n62143, n62144, n62145, n62146, n62147, n62148, n62149, n62150, n62151,
    n62152, n62153, n62154, n62155, n62156, n62158, n62159, n62160, n62161,
    n62162, n62163, n62164, n62165, n62166, n62167, n62168, n62169, n62170,
    n62171, n62172, n62173, n62174, n62175, n62176, n62177, n62178, n62179,
    n62180, n62181, n62182, n62183, n62184, n62185, n62186, n62187, n62188,
    n62190, n62191, n62192, n62193, n62194, n62195, n62196, n62197, n62198,
    n62199, n62200, n62201, n62202, n62203, n62204, n62205, n62206, n62207,
    n62208, n62209, n62210, n62211, n62212, n62213, n62214, n62215, n62216,
    n62217, n62218, n62219, n62220, n62221, n62222, n62223, n62225, n62226,
    n62227, n62228, n62229, n62230, n62231, n62232, n62233, n62234, n62235,
    n62236, n62237, n62238, n62239, n62240, n62241, n62242, n62243, n62244,
    n62245, n62246, n62247, n62248, n62249, n62250, n62251, n62252, n62253,
    n62254, n62255, n62256, n62257, n62258, n62260, n62261, n62262, n62263,
    n62264, n62265, n62266, n62267, n62268, n62269, n62270, n62271, n62272,
    n62273, n62274, n62275, n62276, n62277, n62278, n62279, n62280, n62281,
    n62282, n62283, n62284, n62285, n62286, n62287, n62288, n62289, n62290,
    n62291, n62292, n62293, n62294, n62295, n62296, n62297, n62298, n62299,
    n62300, n62301, n62302, n62303, n62304, n62305, n62306, n62307, n62309,
    n62310, n62311, n62312, n62313, n62314, n62315, n62316, n62317, n62318,
    n62319, n62320, n62321, n62322, n62323, n62324, n62325, n62326, n62327,
    n62328, n62329, n62330, n62331, n62332, n62333, n62334, n62335, n62336,
    n62337, n62338, n62339, n62340, n62341, n62342, n62343, n62344, n62345,
    n62347, n62348, n62349, n62350, n62351, n62352, n62353, n62354, n62355,
    n62356, n62357, n62358, n62359, n62360, n62361, n62362, n62363, n62364,
    n62365, n62366, n62367, n62368, n62369, n62370, n62371, n62372, n62373,
    n62374, n62375, n62377, n62378, n62379, n62380, n62381, n62382, n62383,
    n62384, n62385, n62386, n62387, n62388, n62389, n62390, n62391, n62392,
    n62393, n62394, n62395, n62396, n62397, n62398, n62399, n62400, n62401,
    n62402, n62403, n62404, n62405, n62406, n62407, n62408, n62409, n62410,
    n62411, n62412, n62413, n62414, n62415, n62417, n62418, n62419, n62420,
    n62421, n62422, n62423, n62424, n62425, n62426, n62427, n62428, n62429,
    n62430, n62431, n62432, n62433, n62434, n62435, n62436, n62437, n62438,
    n62439, n62440, n62441, n62442, n62443, n62444, n62445, n62446, n62447,
    n62448, n62449, n62450, n62451, n62452, n62454, n62455, n62456, n62457,
    n62458, n62459, n62460, n62461, n62462, n62463, n62464, n62465, n62466,
    n62467, n62468, n62469, n62470, n62471, n62472, n62473, n62474, n62475,
    n62476, n62477, n62478, n62479, n62480, n62481, n62482, n62483, n62484,
    n62485, n62486, n62487, n62488, n62489, n62490, n62491, n62492, n62493,
    n62494, n62495, n62496, n62497, n62498, n62499, n62500, n62501, n62502,
    n62503, n62504, n62505, n62506, n62507, n62508, n62509, n62510, n62511,
    n62512, n62513, n62514, n62515, n62516, n62517, n62518, n62519, n62520,
    n62521, n62522, n62523, n62524, n62525, n62526, n62527, n62528, n62529,
    n62530, n62531, n62532, n62533, n62534, n62535, n62536, n62537, n62538,
    n62539, n62541, n62542, n62543, n62544, n62545, n62546, n62547, n62548,
    n62549, n62550, n62551, n62552, n62553, n62554, n62555, n62556, n62557,
    n62558, n62559, n62560, n62561, n62562, n62563, n62564, n62565, n62567,
    n62568, n62569, n62570, n62571, n62572, n62573, n62574, n62575, n62576,
    n62577, n62578, n62579, n62580, n62581, n62582, n62583, n62584, n62585,
    n62586, n62587, n62588, n62589, n62590, n62591, n62592, n62593, n62594,
    n62595, n62596, n62597, n62598, n62600, n62601, n62602, n62603, n62604,
    n62605, n62606, n62607, n62608, n62609, n62610, n62611, n62612, n62613,
    n62614, n62615, n62616, n62617, n62618, n62619, n62620, n62621, n62622,
    n62623, n62624, n62625, n62626, n62627, n62628, n62629, n62630, n62631,
    n62632, n62633, n62634, n62635, n62636, n62637, n62638, n62639, n62640,
    n62641, n62642, n62643, n62644, n62645, n62646, n62647, n62648, n62649,
    n62650, n62652, n62653, n62654, n62655, n62656, n62657, n62658, n62659,
    n62660, n62661, n62662, n62663, n62664, n62665, n62666, n62667, n62668,
    n62669, n62670, n62671, n62672, n62673, n62674, n62675, n62676, n62677,
    n62678, n62679, n62680, n62681, n62682, n62683, n62684, n62685, n62686,
    n62687, n62688, n62690, n62691, n62692, n62693, n62694, n62695, n62696,
    n62697, n62698, n62699, n62700, n62701, n62702, n62703, n62704, n62705,
    n62706, n62707, n62708, n62709, n62710, n62711, n62712, n62713, n62714,
    n62715, n62716, n62717, n62718, n62719, n62720, n62721, n62722, n62723,
    n62725, n62726, n62727, n62728, n62729, n62730, n62731, n62732, n62733,
    n62734, n62735, n62736, n62737, n62738, n62739, n62740, n62741, n62742,
    n62743, n62744, n62745, n62746, n62747, n62748, n62749, n62750, n62751,
    n62752, n62753, n62754, n62755, n62756, n62757, n62758, n62759, n62760,
    n62761, n62762, n62763, n62764, n62765, n62766, n62767, n62768, n62769,
    n62770, n62771, n62772, n62773, n62774, n62775, n62776, n62777, n62778,
    n62779, n62780, n62781, n62782, n62783, n62784, n62785, n62786, n62787,
    n62788, n62789, n62790, n62791, n62792, n62793, n62794, n62795, n62796,
    n62797, n62798, n62799, n62800, n62801, n62802, n62803, n62804, n62805,
    n62806, n62807, n62808, n62809, n62810, n62811, n62812, n62813, n62814,
    n62815, n62816, n62817, n62818, n62819, n62820, n62821, n62822, n62823,
    n62824, n62826, n62827, n62828, n62829, n62830, n62831, n62832, n62833,
    n62834, n62835, n62836, n62837, n62838, n62839, n62840, n62841, n62842,
    n62843, n62844, n62845, n62846, n62847, n62848, n62849, n62850, n62851,
    n62852, n62853, n62854, n62855, n62856, n62857, n62858, n62859, n62860,
    n62861, n62862, n62863, n62864, n62865, n62866, n62867, n62868, n62869,
    n62870, n62871, n62872, n62873, n62874, n62875, n62876, n62877, n62878,
    n62879, n62880, n62881, n62882, n62883, n62884, n62885, n62886, n62887,
    n62888, n62889, n62890, n62891, n62892, n62893, n62894, n62895, n62896,
    n62897, n62898, n62899, n62900, n62901, n62902, n62903, n62904, n62905,
    n62906, n62907, n62908, n62909, n62910, n62911, n62912, n62913, n62914,
    n62915, n62916, n62917, n62918, n62919, n62920, n62921, n62922, n62923,
    n62924, n62925, n62926, n62928, n62929, n62930, n62931, n62932, n62933,
    n62934, n62935, n62936, n62937, n62938, n62939, n62940, n62941, n62942,
    n62943, n62944, n62945, n62946, n62947, n62948, n62949, n62950, n62951,
    n62952, n62953, n62954, n62955, n62956, n62957, n62958, n62959, n62961,
    n62962, n62963, n62964, n62965, n62966, n62967, n62968, n62969, n62970,
    n62971, n62972, n62973, n62974, n62975, n62976, n62977, n62978, n62979,
    n62980, n62981, n62982, n62983, n62984, n62985, n62986, n62987, n62988,
    n62989, n62990, n62991, n62992, n62993, n62994, n62995, n62996, n62997,
    n62998, n62999, n63000, n63001, n63002, n63003, n63004, n63005, n63006,
    n63008, n63009, n63010, n63011, n63012, n63013, n63014, n63015, n63016,
    n63017, n63018, n63019, n63020, n63021, n63022, n63023, n63024, n63025,
    n63026, n63027, n63028, n63029, n63030, n63031, n63032, n63033, n63034,
    n63035, n63036, n63037, n63038, n63039, n63040, n63041, n63042, n63043,
    n63044, n63045, n63046, n63047, n63048, n63049, n63050, n63051, n63052,
    n63053, n63054, n63055, n63056, n63057, n63058, n63059, n63060, n63061,
    n63062, n63063, n63064, n63065, n63066, n63067, n63068, n63069, n63070,
    n63071, n63072, n63073, n63074, n63075, n63076, n63077, n63078, n63079,
    n63080, n63081, n63082, n63083, n63084, n63085, n63086, n63087, n63088,
    n63089, n63090, n63091, n63092, n63093, n63094, n63095, n63096, n63097,
    n63098, n63099, n63100, n63101, n63102, n63103, n63104, n63105, n63106,
    n63108, n63109, n63110, n63111, n63112, n63113, n63114, n63115, n63116,
    n63117, n63118, n63119, n63120, n63121, n63122, n63123, n63124, n63125,
    n63126, n63127, n63128, n63129, n63130, n63131, n63132, n63133, n63134,
    n63135, n63136, n63137, n63138, n63139, n63140, n63141, n63142, n63143,
    n63144, n63146, n63147, n63148, n63149, n63150, n63151, n63152, n63153,
    n63154, n63155, n63156, n63157, n63158, n63159, n63160, n63161, n63162,
    n63163, n63164, n63165, n63166, n63167, n63168, n63169, n63170, n63171,
    n63172, n63173, n63174, n63175, n63176, n63177, n63178, n63179, n63180,
    n63181, n63182, n63183, n63184, n63185, n63186, n63187, n63188, n63189,
    n63190, n63191, n63192, n63193, n63194, n63195, n63196, n63197, n63198,
    n63199, n63200, n63201, n63202, n63203, n63204, n63205, n63206, n63207,
    n63208, n63209, n63210, n63211, n63212, n63213, n63214, n63215, n63216,
    n63217, n63218, n63219, n63220, n63221, n63222, n63223, n63224, n63225,
    n63226, n63227, n63228, n63229, n63230, n63231, n63232, n63233, n63234,
    n63235, n63236, n63237, n63238, n63239, n63240, n63241, n63242, n63243,
    n63245, n63246, n63247, n63248, n63249, n63250, n63251, n63252, n63253,
    n63254, n63255, n63256, n63257, n63258, n63259, n63260, n63261, n63262,
    n63263, n63264, n63265, n63266, n63267, n63268, n63269, n63270, n63271,
    n63272, n63273, n63274, n63275, n63276, n63277, n63278, n63279, n63280,
    n63281, n63282, n63283, n63284, n63285, n63286, n63287, n63288, n63289,
    n63290, n63291, n63292, n63293, n63294, n63295, n63296, n63297, n63298,
    n63299, n63300, n63301, n63302, n63303, n63304, n63305, n63306, n63307,
    n63308, n63309, n63310, n63311, n63312, n63313, n63314, n63315, n63316,
    n63317, n63318, n63319, n63320, n63321, n63322, n63323, n63324, n63325,
    n63326, n63327, n63328, n63329, n63330, n63331, n63332, n63333, n63335,
    n63336, n63337, n63338, n63339, n63340, n63341, n63342, n63343, n63344,
    n63345, n63346, n63347, n63348, n63349, n63350, n63351, n63352, n63353,
    n63354, n63355, n63356, n63357, n63358, n63359, n63360, n63361, n63362,
    n63363, n63364, n63365, n63366, n63367, n63368, n63369, n63370, n63371,
    n63372, n63373, n63375, n63376, n63377, n63378, n63379, n63380, n63381,
    n63382, n63383, n63384, n63385, n63386, n63387, n63388, n63389, n63390,
    n63391, n63392, n63393, n63394, n63395, n63396, n63397, n63398, n63399,
    n63400, n63401, n63402, n63403, n63404, n63405, n63406, n63407, n63408,
    n63409, n63410, n63411, n63412, n63413, n63415, n63416, n63417, n63418,
    n63419, n63420, n63421, n63422, n63423, n63424, n63425, n63426, n63427,
    n63428, n63429, n63430, n63431, n63432, n63433, n63434, n63435, n63436,
    n63437, n63438, n63439, n63440, n63441, n63442, n63443, n63444, n63445,
    n63446, n63447, n63448, n63449, n63450, n63451, n63452, n63453, n63454,
    n63455, n63456, n63457, n63458, n63459, n63460, n63461, n63462, n63463,
    n63464, n63465, n63466, n63467, n63468, n63469, n63470, n63471, n63472,
    n63473, n63474, n63475, n63476, n63477, n63478, n63479, n63480, n63481,
    n63482, n63483, n63484, n63485, n63486, n63487, n63488, n63489, n63490,
    n63491, n63492, n63493, n63494, n63495, n63496, n63497, n63498, n63499,
    n63500, n63501, n63502, n63503, n63504, n63505, n63506, n63507, n63508,
    n63509, n63510, n63511, n63512, n63513, n63514, n63515, n63516, n63517,
    n63518, n63519, n63520, n63522, n63523, n63524, n63525, n63526, n63527,
    n63528, n63529, n63530, n63531, n63532, n63533, n63534, n63535, n63536,
    n63537, n63538, n63539, n63540, n63541, n63542, n63543, n63544, n63545,
    n63546, n63547, n63548, n63549, n63550, n63551, n63552, n63553, n63554,
    n63555, n63556, n63557, n63558, n63559, n63561, n63562, n63563, n63564,
    n63565, n63566, n63567, n63568, n63569, n63570, n63571, n63572, n63573,
    n63574, n63575, n63576, n63577, n63578, n63579, n63580, n63581, n63582,
    n63583, n63584, n63585, n63586, n63587, n63588, n63589, n63590, n63591,
    n63592, n63593, n63595, n63596, n63597, n63598, n63599, n63600, n63601,
    n63602, n63603, n63604, n63605, n63606, n63607, n63608, n63609, n63610,
    n63611, n63612, n63613, n63614, n63615, n63616, n63617, n63618, n63619,
    n63620, n63621, n63622, n63623, n63624, n63625, n63626, n63627, n63628,
    n63629, n63630, n63631, n63632, n63633, n63634, n63635, n63636, n63637,
    n63638, n63639, n63640, n63641, n63642, n63643, n63644, n63645, n63646,
    n63647, n63648, n63649, n63650, n63651, n63652, n63653, n63654, n63655,
    n63656, n63657, n63658, n63659, n63660, n63661, n63662, n63663, n63664,
    n63665, n63666, n63667, n63668, n63669, n63670, n63671, n63672, n63673,
    n63674, n63675, n63676, n63677, n63678, n63679, n63680, n63681, n63682,
    n63683, n63684, n63685, n63686, n63687, n63688, n63689, n63690, n63691,
    n63692, n63693, n63694, n63695, n63696, n63697, n63698, n63700, n63701,
    n63702, n63703, n63704, n63705, n63706, n63707, n63708, n63709, n63710,
    n63711, n63712, n63713, n63714, n63715, n63716, n63717, n63718, n63719,
    n63720, n63721, n63722, n63723, n63724, n63725, n63726, n63727, n63728,
    n63729, n63730, n63731, n63732, n63733, n63734, n63735, n63737, n63738,
    n63739, n63740, n63741, n63742, n63743, n63744, n63745, n63746, n63747,
    n63748, n63749, n63750, n63751, n63752, n63753, n63754, n63755, n63756,
    n63757, n63758, n63759, n63760, n63761, n63762, n63763, n63764, n63765,
    n63766, n63767, n63768, n63769, n63770, n63771, n63772, n63773, n63774,
    n63776, n63777, n63778, n63779, n63780, n63781, n63782, n63783, n63784,
    n63785, n63786, n63787, n63788, n63789, n63790, n63791, n63792, n63793,
    n63794, n63795, n63796, n63797, n63798, n63799, n63800, n63801, n63802,
    n63803, n63804, n63805, n63806, n63807, n63808, n63809, n63810, n63811,
    n63812, n63813, n63814, n63815, n63816, n63817, n63818, n63819, n63820,
    n63821, n63822, n63823, n63825, n63826, n63827, n63828, n63829, n63830,
    n63831, n63832, n63833, n63834, n63835, n63836, n63837, n63838, n63839,
    n63840, n63841, n63842, n63843, n63844, n63845, n63846, n63847, n63848,
    n63849, n63850, n63851, n63852, n63853, n63854, n63855, n63856, n63857,
    n63858, n63859, n63860, n63861, n63862, n63863, n63864, n63865, n63866,
    n63867, n63868, n63869, n63870, n63872, n63873, n63874, n63875, n63876,
    n63877, n63878, n63879, n63880, n63881, n63882, n63883, n63884, n63885,
    n63886, n63887, n63888, n63889, n63890, n63891, n63892, n63893, n63894,
    n63895, n63896, n63897, n63898, n63899, n63900, n63901, n63902, n63903,
    n63904, n63905, n63906, n63907, n63908, n63909, n63910, n63911, n63913,
    n63914, n63915, n63916, n63917, n63918, n63919, n63920, n63921, n63922,
    n63923, n63924, n63925, n63926, n63927, n63928, n63929, n63930, n63931,
    n63932, n63933, n63934, n63935, n63936, n63937, n63938, n63939, n63940,
    n63941, n63942, n63943, n63944, n63945, n63946, n63947, n63948, n63949,
    n63950, n63951, n63952, n63953, n63954, n63955, n63956, n63957, n63958,
    n63959, n63960, n63961, n63962, n63964, n63965, n63966, n63967, n63968,
    n63969, n63970, n63971, n63972, n63973, n63974, n63975, n63976, n63977,
    n63978, n63979, n63980, n63981, n63982, n63983, n63984, n63985, n63986,
    n63987, n63988, n63989, n63990, n63991, n63992, n63993, n63994, n63995,
    n63996, n63997, n63998, n64000, n64001, n64002, n64003, n64004, n64005,
    n64006, n64007, n64008, n64009, n64010, n64011, n64012, n64013, n64014,
    n64015, n64016, n64017, n64018, n64019, n64020, n64021, n64022, n64023,
    n64024, n64025, n64026, n64027, n64028, n64029, n64030, n64031, n64032,
    n64033, n64034, n64035, n64036, n64038, n64039, n64040, n64041, n64042,
    n64043, n64044, n64045, n64046, n64047, n64048, n64049, n64050, n64051,
    n64052, n64053, n64054, n64055, n64056, n64057, n64058, n64059, n64060,
    n64061, n64062, n64063, n64064, n64065, n64066, n64067, n64068, n64069,
    n64070, n64072, n64073, n64074, n64075, n64076, n64077, n64078, n64079,
    n64080, n64081, n64082, n64083, n64084, n64085, n64086, n64087, n64088,
    n64089, n64090, n64091, n64092, n64093, n64094, n64095, n64096, n64097,
    n64098, n64099, n64100, n64101, n64102, n64103, n64104, n64105, n64106,
    n64107, n64108, n64109, n64111, n64112, n64113, n64114, n64115, n64116,
    n64117, n64118, n64119, n64120, n64121, n64122, n64123, n64124, n64125,
    n64126, n64127, n64128, n64129, n64130, n64131, n64132, n64133, n64134,
    n64135, n64136, n64137, n64138, n64139, n64140, n64141, n64142, n64143,
    n64144, n64145, n64146, n64147, n64148, n64149, n64150, n64151, n64152,
    n64153, n64154, n64155, n64156, n64157, n64158, n64159, n64160, n64161,
    n64162, n64163, n64164, n64165, n64166, n64167, n64168, n64169, n64170,
    n64171, n64172, n64173, n64174, n64175, n64176, n64177, n64178, n64179,
    n64180, n64181, n64182, n64183, n64184, n64185, n64186, n64187, n64188,
    n64189, n64190, n64191, n64192, n64193, n64194, n64195, n64196, n64197,
    n64198, n64199, n64200, n64201, n64202, n64203, n64204, n64206, n64207,
    n64208, n64209, n64210, n64211, n64212, n64213, n64214, n64215, n64216,
    n64217, n64218, n64219, n64220, n64221, n64222, n64223, n64224, n64225,
    n64226, n64227, n64228, n64229, n64230, n64231, n64232, n64233, n64234,
    n64235, n64236, n64237, n64238, n64239, n64240, n64241, n64242, n64243,
    n64244, n64245, n64246, n64247, n64248, n64249, n64250, n64251, n64253,
    n64254, n64255, n64256, n64257, n64258, n64259, n64260, n64261, n64262,
    n64263, n64264, n64265, n64266, n64267, n64268, n64269, n64270, n64271,
    n64272, n64273, n64274, n64275, n64276, n64277, n64278, n64279, n64280,
    n64281, n64282, n64283, n64284, n64285, n64286, n64288, n64289, n64290,
    n64291, n64292, n64293, n64294, n64295, n64296, n64297, n64298, n64299,
    n64300, n64301, n64302, n64303, n64304, n64305, n64306, n64307, n64308,
    n64309, n64310, n64311, n64312, n64313, n64314, n64315, n64316, n64317,
    n64319, n64320, n64321, n64322, n64323, n64324, n64325, n64326, n64327,
    n64328, n64329, n64330, n64331, n64332, n64333, n64334, n64335, n64336,
    n64337, n64338, n64339, n64340, n64341, n64342, n64343, n64344, n64345,
    n64346, n64347, n64348, n64349, n64350, n64351, n64352, n64354, n64355,
    n64356, n64357, n64358, n64359, n64360, n64361, n64362, n64363, n64364,
    n64365, n64366, n64367, n64368, n64369, n64370, n64371, n64372, n64373,
    n64374, n64375, n64376, n64377, n64378, n64379, n64380, n64381, n64382,
    n64383, n64384, n64385, n64386, n64387, n64388, n64390, n64391, n64392,
    n64393, n64394, n64395, n64396, n64397, n64398, n64399, n64400, n64401,
    n64402, n64403, n64404, n64405, n64406, n64407, n64408, n64409, n64410,
    n64411, n64412, n64413, n64414, n64415, n64416, n64417, n64418, n64420,
    n64421, n64422, n64423, n64424, n64425, n64426, n64427, n64428, n64429,
    n64430, n64431, n64432, n64433, n64434, n64435, n64436, n64437, n64438,
    n64439, n64440, n64441, n64442, n64443, n64444, n64446, n64447, n64448,
    n64449, n64450, n64451, n64452, n64453, n64454, n64455, n64456, n64457,
    n64458, n64459, n64460, n64461, n64462, n64463, n64464, n64465, n64466,
    n64467, n64468, n64469, n64470, n64471, n64472, n64473, n64474, n64475,
    n64476, n64477, n64478, n64479, n64480, n64481, n64482, n64483, n64484,
    n64485, n64486, n64487, n64488, n64489, n64490, n64491, n64492, n64493,
    n64494, n64495, n64496, n64497, n64498, n64499, n64500, n64501, n64502,
    n64503, n64504, n64505, n64506, n64507, n64508, n64509, n64510, n64511,
    n64512, n64513, n64514, n64515, n64516, n64517, n64518, n64519, n64520,
    n64521, n64522, n64523, n64524, n64525, n64526, n64527, n64528, n64529,
    n64530, n64531, n64532, n64533, n64534, n64535, n64536, n64537, n64538,
    n64539, n64540, n64541, n64542, n64543, n64545, n64546, n64547, n64548,
    n64549, n64550, n64551, n64552, n64553, n64554, n64555, n64556, n64557,
    n64558, n64559, n64560, n64561, n64562, n64563, n64564, n64565, n64566,
    n64567, n64568, n64569, n64570, n64571, n64572, n64573, n64574, n64575,
    n64576, n64577, n64578, n64579, n64580, n64581, n64582, n64583, n64584,
    n64585, n64586, n64587, n64588, n64589, n64590, n64591, n64592, n64593,
    n64594, n64595, n64596, n64597, n64598, n64599, n64600, n64601, n64602,
    n64603, n64604, n64605, n64606, n64607, n64608, n64609, n64610, n64611,
    n64612, n64613, n64614, n64615, n64616, n64617, n64618, n64619, n64620,
    n64621, n64622, n64623, n64624, n64625, n64626, n64627, n64628, n64629,
    n64630, n64631, n64632, n64633, n64634, n64635, n64636, n64637, n64638,
    n64639, n64640, n64641, n64642, n64644, n64645, n64646, n64647, n64648,
    n64649, n64650, n64651, n64652, n64653, n64654, n64655, n64656, n64657,
    n64658, n64659, n64660, n64661, n64662, n64663, n64664, n64665, n64666,
    n64667, n64668, n64669, n64670, n64671, n64672, n64673, n64674, n64675,
    n64676, n64677, n64678, n64679, n64680, n64681, n64682, n64684, n64685,
    n64686, n64687, n64688, n64689, n64690, n64691, n64692, n64693, n64694,
    n64695, n64696, n64697, n64698, n64699, n64700, n64701, n64702, n64703,
    n64704, n64705, n64706, n64707, n64708, n64709, n64710, n64711, n64712,
    n64713, n64714, n64715, n64716, n64717, n64718, n64719, n64720, n64721,
    n64722, n64723, n64724, n64725, n64726, n64727, n64728, n64729, n64730,
    n64731, n64732, n64733, n64734, n64735, n64736, n64737, n64738, n64739,
    n64740, n64741, n64742, n64743, n64744, n64745, n64746, n64747, n64748,
    n64749, n64750, n64751, n64752, n64753, n64754, n64755, n64756, n64757,
    n64758, n64759, n64760, n64761, n64762, n64763, n64764, n64765, n64766,
    n64767, n64768, n64769, n64770, n64771, n64772, n64773, n64774, n64775,
    n64776, n64777, n64778, n64779, n64780, n64781, n64783, n64784, n64785,
    n64786, n64787, n64788, n64789, n64790, n64791, n64792, n64793, n64794,
    n64795, n64796, n64797, n64798, n64799, n64800, n64801, n64802, n64803,
    n64804, n64805, n64806, n64807, n64808, n64809, n64810, n64811, n64812,
    n64813, n64814, n64815, n64816, n64817, n64818, n64819, n64820, n64821,
    n64822, n64823, n64824, n64825, n64826, n64827, n64828, n64829, n64830,
    n64831, n64832, n64833, n64834, n64835, n64836, n64837, n64838, n64839,
    n64840, n64841, n64842, n64843, n64844, n64845, n64846, n64847, n64848,
    n64849, n64850, n64851, n64852, n64853, n64854, n64855, n64856, n64857,
    n64858, n64859, n64860, n64861, n64862, n64863, n64864, n64865, n64866,
    n64867, n64868, n64869, n64870, n64871, n64872, n64873, n64874, n64875,
    n64876, n64877, n64878, n64879, n64880, n64881, n64882, n64883, n64884,
    n64885, n64886, n64887, n64888, n64890, n64891, n64892, n64893, n64894,
    n64895, n64896, n64897, n64898, n64899, n64900, n64901, n64902, n64903,
    n64904, n64905, n64906, n64907, n64908, n64909, n64910, n64911, n64912,
    n64913, n64914, n64915, n64916, n64917, n64918, n64919, n64920, n64921,
    n64922, n64923, n64924, n64925, n64926, n64927, n64928, n64929, n64930,
    n64931, n64932, n64933, n64934, n64935, n64936, n64937, n64938, n64939,
    n64940, n64941, n64942, n64943, n64944, n64945, n64946, n64947, n64948,
    n64949, n64950, n64951, n64952, n64953, n64954, n64955, n64956, n64957,
    n64958, n64959, n64960, n64961, n64962, n64963, n64964, n64965, n64966,
    n64967, n64968, n64969, n64970, n64971, n64972, n64973, n64974, n64975,
    n64976, n64977, n64978, n64979, n64980, n64981, n64982, n64983, n64984,
    n64985, n64986, n64987, n64988, n64989, n64990, n64992, n64993, n64994,
    n64995, n64996, n64997, n64998, n64999, n65000, n65001, n65002, n65003,
    n65004, n65005, n65006, n65007, n65008, n65009, n65010, n65011, n65012,
    n65013, n65014, n65015, n65016, n65017, n65018, n65019, n65020, n65021,
    n65022, n65023, n65024, n65025, n65026, n65027, n65028, n65030, n65031,
    n65032, n65033, n65034, n65035, n65036, n65037, n65038, n65039, n65040,
    n65041, n65042, n65043, n65044, n65045, n65046, n65047, n65048, n65049,
    n65050, n65051, n65052, n65053, n65054, n65055, n65056, n65057, n65058,
    n65059, n65060, n65061, n65062, n65063, n65064, n65065, n65067, n65068,
    n65069, n65070, n65071, n65072, n65073, n65074, n65075, n65076, n65077,
    n65078, n65079, n65080, n65081, n65082, n65083, n65084, n65085, n65086,
    n65087, n65088, n65089, n65090, n65091, n65092, n65093, n65094, n65095,
    n65096, n65097, n65098, n65099, n65100, n65101, n65102, n65103, n65104,
    n65105, n65106, n65108, n65109, n65110, n65111, n65112, n65113, n65114,
    n65115, n65116, n65117, n65118, n65119, n65120, n65121, n65122, n65123,
    n65124, n65125, n65126, n65127, n65128, n65129, n65130, n65131, n65132,
    n65133, n65134, n65135, n65136, n65137, n65138, n65139, n65140, n65141,
    n65142, n65143, n65144, n65145, n65146, n65147, n65148, n65149, n65150,
    n65151, n65152, n65153, n65154, n65155, n65156, n65157, n65158, n65159,
    n65160, n65161, n65162, n65163, n65164, n65165, n65166, n65167, n65168,
    n65169, n65170, n65171, n65172, n65173, n65174, n65175, n65176, n65177,
    n65178, n65179, n65180, n65181, n65182, n65183, n65184, n65185, n65186,
    n65187, n65188, n65189, n65190, n65191, n65192, n65193, n65194, n65195,
    n65196, n65197, n65198, n65199, n65200, n65201, n65202, n65203, n65204,
    n65205, n65206, n65207, n65208, n65210, n65211, n65212, n65213, n65214,
    n65215, n65216, n65217, n65218, n65219, n65220, n65221, n65222, n65223,
    n65224, n65225, n65226, n65227, n65228, n65229, n65230, n65231, n65232,
    n65233, n65234, n65235, n65236, n65237, n65238, n65239, n65240, n65241,
    n65242, n65243, n65244, n65245, n65246, n65247, n65248, n65249, n65250,
    n65251, n65252, n65253, n65254, n65255, n65256, n65257, n65258, n65259,
    n65260, n65261, n65262, n65263, n65264, n65265, n65266, n65267, n65268,
    n65269, n65270, n65271, n65272, n65273, n65274, n65275, n65276, n65277,
    n65278, n65279, n65280, n65281, n65282, n65283, n65284, n65285, n65286,
    n65287, n65288, n65289, n65290, n65291, n65292, n65293, n65294, n65295,
    n65296, n65297, n65298, n65299, n65300, n65301, n65302, n65303, n65304,
    n65306, n65307, n65308, n65309, n65310, n65311, n65312, n65313, n65314,
    n65315, n65316, n65317, n65318, n65319, n65320, n65321, n65322, n65323,
    n65324, n65325, n65326, n65327, n65328, n65329, n65330, n65331, n65332,
    n65333, n65334, n65335, n65336, n65337, n65338, n65339, n65340, n65341,
    n65342, n65343, n65344, n65346, n65347, n65348, n65349, n65350, n65351,
    n65352, n65353, n65354, n65355, n65356, n65357, n65358, n65359, n65360,
    n65361, n65362, n65363, n65364, n65365, n65366, n65367, n65368, n65369,
    n65370, n65371, n65372, n65373, n65374, n65375, n65376, n65377, n65378,
    n65379, n65380, n65381, n65382, n65383, n65384, n65385, n65386, n65387,
    n65389, n65390, n65391, n65392, n65393, n65394, n65395, n65396, n65397,
    n65398, n65399, n65400, n65401, n65402, n65403, n65404, n65405, n65406,
    n65407, n65408, n65409, n65410, n65411, n65412, n65413, n65414, n65415,
    n65416, n65417, n65418, n65419, n65420, n65421, n65422, n65423, n65424,
    n65425, n65426, n65427, n65428, n65429, n65430, n65431, n65432, n65434,
    n65435, n65436, n65437, n65438, n65439, n65440, n65441, n65442, n65443,
    n65444, n65445, n65446, n65447, n65448, n65449, n65450, n65451, n65452,
    n65453, n65454, n65455, n65456, n65457, n65458, n65459, n65460, n65461,
    n65462, n65463, n65464, n65465, n65466, n65467, n65468, n65469, n65470,
    n65471, n65472, n65473, n65475, n65476, n65477, n65478, n65479, n65480,
    n65481, n65482, n65483, n65484, n65485, n65486, n65487, n65488, n65489,
    n65490, n65491, n65492, n65493, n65494, n65495, n65496, n65497, n65498,
    n65499, n65500, n65501, n65502, n65503, n65504, n65505, n65506, n65507,
    n65508, n65509, n65510, n65511, n65512, n65513, n65514, n65515, n65516,
    n65517, n65518, n65519, n65520, n65521, n65522, n65523, n65524, n65525,
    n65526, n65527, n65528, n65529, n65530, n65531, n65532, n65533, n65534,
    n65535, n65536, n65537, n65538, n65539, n65540, n65541, n65542, n65543,
    n65544, n65545, n65546, n65547, n65548, n65549, n65550, n65551, n65552,
    n65553, n65554, n65555, n65556, n65557, n65558, n65559, n65560, n65561,
    n65562, n65564, n65565, n65566, n65567, n65568, n65569, n65570, n65571,
    n65572, n65573, n65574, n65575, n65576, n65577, n65578, n65579, n65580,
    n65581, n65582, n65583, n65584, n65585, n65586, n65587, n65588, n65589,
    n65590, n65591, n65592, n65593, n65594, n65595, n65597, n65598, n65599,
    n65600, n65601, n65602, n65603, n65604, n65605, n65606, n65607, n65608,
    n65609, n65610, n65611, n65612, n65613, n65614, n65615, n65616, n65617,
    n65618, n65619, n65620, n65621, n65622, n65623, n65624, n65625, n65626,
    n65627, n65628, n65629, n65630, n65631, n65632, n65633, n65634, n65636,
    n65637, n65638, n65639, n65640, n65641, n65642, n65643, n65644, n65645,
    n65646, n65647, n65648, n65649, n65650, n65651, n65652, n65653, n65654,
    n65655, n65656, n65657, n65658, n65659, n65660, n65661, n65662, n65663,
    n65664, n65665, n65666, n65667, n65668, n65669, n65670, n65671, n65672,
    n65673, n65674, n65675, n65676, n65677, n65678, n65679, n65680, n65681,
    n65683, n65684, n65685, n65686, n65687, n65688, n65689, n65690, n65691,
    n65692, n65693, n65694, n65695, n65696, n65697, n65698, n65699, n65700,
    n65701, n65702, n65703, n65704, n65705, n65706, n65707, n65708, n65709,
    n65710, n65711, n65712, n65713, n65714, n65715, n65716, n65717, n65718,
    n65719, n65721, n65722, n65723, n65724, n65725, n65726, n65727, n65728,
    n65729, n65730, n65731, n65732, n65733, n65734, n65735, n65736, n65737,
    n65738, n65739, n65740, n65741, n65742, n65743, n65744, n65745, n65746,
    n65747, n65748, n65749, n65750, n65751, n65752, n65753, n65754, n65755,
    n65756, n65757, n65758, n65759, n65760, n65761, n65762, n65763, n65765,
    n65766, n65767, n65768, n65769, n65770, n65771, n65772, n65773, n65774,
    n65775, n65776, n65777, n65778, n65779, n65780, n65781, n65782, n65783,
    n65784, n65785, n65786, n65787, n65788, n65789, n65790, n65791, n65792,
    n65793, n65795, n65796, n65797, n65798, n65799, n65800, n65801, n65802,
    n65803, n65804, n65805, n65806, n65807, n65808, n65809, n65810, n65811,
    n65812, n65813, n65814, n65815, n65816, n65817, n65818, n65819, n65820,
    n65821, n65822, n65823, n65824, n65825, n65826, n65827, n65828, n65829,
    n65830, n65831, n65832, n65833, n65834, n65835, n65836, n65837, n65838,
    n65840, n65841, n65842, n65843, n65844, n65845, n65846, n65847, n65848,
    n65849, n65850, n65851, n65852, n65853, n65854, n65855, n65856, n65857,
    n65858, n65859, n65860, n65861, n65862, n65863, n65864, n65865, n65866,
    n65867, n65868, n65869, n65870, n65871, n65872, n65873, n65875, n65876,
    n65877, n65878, n65879, n65880, n65881, n65882, n65883, n65884, n65885,
    n65886, n65887, n65888, n65889, n65890, n65891, n65892, n65893, n65894,
    n65895, n65896, n65897, n65898, n65899, n65900, n65901, n65902, n65903,
    n65904, n65905, n65906, n65907, n65908, n65909, n65910, n65911, n65912,
    n65913, n65915, n65916, n65917, n65918, n65919, n65920, n65921, n65922,
    n65923, n65924, n65925, n65926, n65927, n65928, n65929, n65930, n65931,
    n65932, n65933, n65934, n65935, n65936, n65937, n65938, n65939, n65940,
    n65941, n65942, n65943, n65944, n65945, n65946, n65948, n65949, n65950,
    n65951, n65952, n65953, n65954, n65955, n65956, n65957, n65958, n65959,
    n65960, n65961, n65962, n65963, n65964, n65965, n65966, n65967, n65968,
    n65969, n65970, n65971, n65972, n65973, n65974, n65975, n65976, n65977,
    n65978, n65979, n65980, n65981, n65982, n65983, n65984, n65985, n65986,
    n65987, n65988, n65989, n65990, n65991, n65992, n65993, n65995, n65996,
    n65997, n65998, n65999, n66000, n66001, n66002, n66003, n66004, n66005,
    n66006, n66007, n66008, n66009, n66010, n66011, n66012, n66013, n66014,
    n66015, n66016, n66017, n66018, n66019, n66020, n66021, n66022, n66023,
    n66024, n66025, n66026, n66027, n66028, n66029, n66030, n66031, n66033,
    n66034, n66035, n66036, n66037, n66038, n66039, n66040, n66041, n66042,
    n66043, n66044, n66045, n66046, n66047, n66048, n66049, n66050, n66051,
    n66052, n66053, n66054, n66055, n66056, n66057, n66058, n66059, n66060,
    n66061, n66062, n66063, n66064, n66065, n66066, n66067, n66068, n66070,
    n66071, n66072, n66073, n66074, n66075, n66076, n66077, n66078, n66079,
    n66080, n66081, n66082, n66083, n66084, n66085, n66086, n66087, n66088,
    n66089, n66090, n66091, n66092, n66093, n66094, n66095, n66096, n66097,
    n66098, n66100, n66101, n66102, n66103, n66104, n66105, n66106, n66107,
    n66108, n66109, n66110, n66111, n66112, n66113, n66114, n66115, n66116,
    n66117, n66118, n66119, n66120, n66121, n66122, n66123, n66124, n66126,
    n66127, n66128, n66129, n66130, n66131, n66132, n66133, n66134, n66135,
    n66136, n66137, n66138, n66139, n66140, n66141, n66142, n66143, n66144,
    n66145, n66146, n66147, n66148, n66149, n66150, n66151, n66152, n66153,
    n66154, n66155, n66156, n66157, n66159, n66160, n66161, n66162, n66163,
    n66164, n66165, n66166, n66167, n66168, n66169, n66170, n66171, n66172,
    n66173, n66174, n66175, n66176, n66177, n66178, n66179, n66180, n66181,
    n66182, n66183, n66184, n66185, n66186, n66187, n66188, n66189, n66190,
    n66191, n66192, n66193, n66194, n66195, n66196, n66197, n66198, n66199,
    n66200, n66201, n66202, n66203, n66204, n66205, n66206, n66207, n66208,
    n66209, n66210, n66211, n66212, n66213, n66214, n66215, n66216, n66217,
    n66218, n66219, n66220, n66221, n66222, n66223, n66224, n66225, n66226,
    n66227, n66228, n66229, n66230, n66231, n66232, n66233, n66234, n66235,
    n66236, n66237, n66238, n66239, n66240, n66241, n66242, n66243, n66244,
    n66245, n66246, n66247, n66248, n66249, n66250, n66251, n66252, n66253,
    n66254, n66255, n66256, n66258, n66259, n66260, n66261, n66262, n66263,
    n66264, n66265, n66266, n66267, n66268, n66269, n66270, n66271, n66272,
    n66273, n66274, n66275, n66276, n66277, n66278, n66279, n66280, n66281,
    n66282, n66283, n66284, n66285, n66286, n66287, n66288, n66289, n66290,
    n66291, n66292, n66293, n66294, n66295, n66296, n66297, n66298, n66299,
    n66300, n66301, n66302, n66303, n66304, n66305, n66306, n66307, n66308,
    n66309, n66310, n66311, n66312, n66313, n66314, n66315, n66316, n66317,
    n66318, n66319, n66320, n66321, n66322, n66323, n66324, n66325, n66326,
    n66327, n66328, n66329, n66330, n66331, n66332, n66333, n66334, n66335,
    n66336, n66337, n66338, n66339, n66340, n66341, n66342, n66343, n66344,
    n66345, n66346, n66347, n66348, n66349, n66350, n66351, n66352, n66353,
    n66354, n66355, n66356, n66357, n66358, n66360, n66361, n66362, n66363,
    n66364, n66365, n66366, n66367, n66368, n66369, n66370, n66371, n66372,
    n66373, n66374, n66375, n66376, n66377, n66378, n66379, n66380, n66381,
    n66382, n66383, n66384, n66385, n66386, n66387, n66388, n66389, n66390,
    n66391, n66392, n66393, n66394, n66395, n66396, n66397, n66398, n66399,
    n66400, n66401, n66402, n66403, n66404, n66405, n66406, n66407, n66408,
    n66409, n66410, n66411, n66412, n66413, n66414, n66415, n66416, n66417,
    n66418, n66419, n66420, n66421, n66422, n66423, n66424, n66425, n66426,
    n66427, n66428, n66429, n66430, n66431, n66432, n66433, n66434, n66435,
    n66436, n66437, n66438, n66439, n66440, n66441, n66442, n66443, n66444,
    n66445, n66446, n66447, n66448, n66449, n66450, n66451, n66452, n66453,
    n66454, n66455, n66456, n66457, n66458, n66459, n66460, n66461, n66462,
    n66463, n66464, n66465, n66467, n66468, n66469, n66470, n66471, n66472,
    n66473, n66474, n66475, n66476, n66477, n66478, n66479, n66480, n66481,
    n66482, n66483, n66484, n66485, n66486, n66487, n66488, n66489, n66490,
    n66491, n66492, n66493, n66494, n66495, n66496, n66497, n66498, n66499,
    n66500, n66501, n66502, n66503, n66504, n66505, n66506, n66507, n66508,
    n66509, n66510, n66511, n66512, n66513, n66514, n66515, n66516, n66517,
    n66518, n66519, n66520, n66521, n66522, n66523, n66524, n66525, n66526,
    n66527, n66528, n66529, n66530, n66531, n66532, n66533, n66534, n66535,
    n66536, n66537, n66538, n66539, n66540, n66541, n66542, n66543, n66544,
    n66545, n66546, n66547, n66548, n66549, n66550, n66551, n66552, n66553,
    n66554, n66555, n66556, n66557, n66558, n66559, n66560, n66561, n66562,
    n66563, n66564, n66565, n66566, n66567, n66568, n66569, n66570, n66572,
    n66573, n66574, n66575, n66576, n66577, n66578, n66579, n66580, n66581,
    n66582, n66583, n66584, n66585, n66586, n66587, n66588, n66589, n66590,
    n66591, n66592, n66593, n66594, n66595, n66596, n66597, n66598, n66599,
    n66600, n66601, n66602, n66603, n66604, n66605, n66606, n66607, n66608,
    n66609, n66610, n66611, n66612, n66613, n66614, n66615, n66616, n66617,
    n66618, n66619, n66620, n66621, n66622, n66623, n66624, n66625, n66626,
    n66627, n66628, n66629, n66630, n66631, n66632, n66633, n66634, n66635,
    n66636, n66637, n66638, n66639, n66640, n66641, n66642, n66643, n66644,
    n66645, n66646, n66647, n66648, n66649, n66650, n66651, n66652, n66653,
    n66654, n66655, n66656, n66657, n66658, n66659, n66660, n66661, n66662,
    n66663, n66664, n66665, n66666, n66667, n66668, n66669, n66670, n66671,
    n66672, n66673, n66674, n66676, n66677, n66678, n66679, n66680, n66681,
    n66682, n66683, n66684, n66685, n66686, n66687, n66688, n66689, n66690,
    n66691, n66692, n66693, n66694, n66695, n66696, n66697, n66698, n66699,
    n66700, n66701, n66702, n66703, n66704, n66705, n66706, n66707, n66708,
    n66709, n66710, n66711, n66712, n66713, n66714, n66715, n66717, n66718,
    n66719, n66720, n66721, n66722, n66723, n66724, n66725, n66726, n66727,
    n66728, n66729, n66730, n66731, n66732, n66733, n66734, n66735, n66736,
    n66737, n66738, n66739, n66740, n66741, n66742, n66743, n66744, n66745,
    n66746, n66747, n66748, n66749, n66750, n66751, n66752, n66753, n66754,
    n66755, n66756, n66757, n66758, n66759, n66760, n66761, n66762, n66763,
    n66764, n66765, n66766, n66767, n66768, n66769, n66770, n66771, n66772,
    n66773, n66774, n66775, n66776, n66777, n66778, n66779, n66780, n66781,
    n66782, n66783, n66784, n66785, n66786, n66787, n66788, n66789, n66790,
    n66791, n66792, n66793, n66794, n66795, n66796, n66797, n66798, n66799,
    n66800, n66801, n66802, n66803, n66804, n66805, n66807, n66808, n66809,
    n66810, n66811, n66812, n66813, n66814, n66815, n66816, n66817, n66818,
    n66819, n66820, n66821, n66822, n66823, n66824, n66825, n66826, n66827,
    n66828, n66829, n66830, n66831, n66832, n66833, n66834, n66835, n66836,
    n66837, n66838, n66839, n66840, n66841, n66842, n66843, n66844, n66845,
    n66846, n66847, n66848, n66849, n66850, n66851, n66852, n66853, n66854,
    n66855, n66856, n66858, n66859, n66860, n66861, n66862, n66863, n66864,
    n66865, n66866, n66867, n66868, n66869, n66870, n66871, n66872, n66873,
    n66874, n66875, n66876, n66877, n66878, n66879, n66880, n66881, n66882,
    n66883, n66884, n66885, n66886, n66887, n66888, n66889, n66891, n66892,
    n66893, n66894, n66895, n66896, n66897, n66898, n66899, n66900, n66901,
    n66902, n66903, n66904, n66905, n66906, n66907, n66908, n66909, n66910,
    n66911, n66912, n66913, n66914, n66915, n66916, n66917, n66918, n66919,
    n66920, n66921, n66922, n66923, n66924, n66925, n66926, n66927, n66928,
    n66929, n66930, n66931, n66932, n66933, n66934, n66935, n66936, n66937,
    n66938, n66939, n66940, n66941, n66942, n66943, n66944, n66945, n66946,
    n66947, n66948, n66949, n66950, n66951, n66952, n66953, n66954, n66955,
    n66956, n66957, n66958, n66959, n66960, n66961, n66962, n66963, n66964,
    n66965, n66966, n66967, n66968, n66969, n66970, n66971, n66972, n66973,
    n66974, n66975, n66976, n66977, n66978, n66979, n66980, n66981, n66982,
    n66983, n66984, n66985, n66986, n66987, n66988, n66990, n66991, n66992,
    n66993, n66994, n66995, n66996, n66997, n66998, n66999, n67000, n67001,
    n67002, n67003, n67004, n67005, n67006, n67007, n67008, n67009, n67010,
    n67011, n67012, n67013, n67014, n67015, n67016, n67017, n67018, n67019,
    n67020, n67021, n67022, n67023, n67024, n67025, n67026, n67027, n67028,
    n67029, n67030, n67031, n67032, n67033, n67034, n67035, n67037, n67038,
    n67039, n67040, n67041, n67042, n67043, n67044, n67045, n67046, n67047,
    n67048, n67049, n67050, n67051, n67052, n67053, n67054, n67055, n67056,
    n67057, n67058, n67059, n67060, n67061, n67062, n67063, n67064, n67065,
    n67066, n67067, n67068, n67069, n67070, n67071, n67072, n67073, n67074,
    n67075, n67076, n67077, n67079, n67080, n67081, n67082, n67083, n67084,
    n67085, n67086, n67087, n67088, n67089, n67090, n67091, n67092, n67093,
    n67094, n67095, n67096, n67097, n67098, n67099, n67100, n67101, n67102,
    n67103, n67104, n67105, n67106, n67107, n67108, n67109, n67110, n67111,
    n67112, n67113, n67114, n67115, n67117, n67118, n67119, n67120, n67121,
    n67122, n67123, n67124, n67125, n67126, n67127, n67128, n67129, n67130,
    n67131, n67132, n67133, n67134, n67135, n67136, n67137, n67138, n67139,
    n67140, n67141, n67142, n67143, n67144, n67145, n67146, n67147, n67148,
    n67149, n67150, n67151, n67152, n67153, n67154, n67156, n67157, n67158,
    n67159, n67160, n67161, n67162, n67163, n67164, n67165, n67166, n67167,
    n67168, n67169, n67170, n67171, n67172, n67173, n67174, n67175, n67176,
    n67177, n67178, n67179, n67180, n67181, n67182, n67183, n67184, n67186,
    n67187, n67188, n67189, n67190, n67191, n67192, n67193, n67194, n67195,
    n67196, n67197, n67198, n67199, n67200, n67201, n67202, n67203, n67204,
    n67205, n67206, n67207, n67208, n67209, n67210, n67211, n67212, n67213,
    n67214, n67215, n67216, n67217, n67218, n67220, n67221, n67222, n67223,
    n67224, n67225, n67226, n67227, n67228, n67229, n67230, n67231, n67232,
    n67233, n67234, n67235, n67236, n67237, n67238, n67239, n67240, n67241,
    n67242, n67243, n67244, n67245, n67246, n67247, n67248, n67249, n67250,
    n67251, n67252, n67253, n67254, n67255, n67256, n67257, n67258, n67259,
    n67260, n67261, n67262, n67263, n67264, n67265, n67267, n67268, n67269,
    n67270, n67271, n67272, n67273, n67274, n67275, n67276, n67277, n67278,
    n67279, n67280, n67281, n67282, n67283, n67284, n67285, n67286, n67287,
    n67288, n67289, n67290, n67291, n67292, n67293, n67294, n67295, n67296,
    n67297, n67298, n67299, n67300, n67302, n67303, n67304, n67305, n67306,
    n67307, n67308, n67309, n67310, n67311, n67312, n67313, n67314, n67315,
    n67316, n67317, n67318, n67319, n67320, n67321, n67322, n67323, n67324,
    n67325, n67326, n67327, n67328, n67329, n67330, n67331, n67332, n67333,
    n67334, n67335, n67336, n67337, n67339, n67340, n67341, n67342, n67343,
    n67344, n67345, n67346, n67347, n67348, n67349, n67350, n67351, n67352,
    n67353, n67354, n67355, n67356, n67357, n67358, n67359, n67360, n67361,
    n67362, n67363, n67364, n67365, n67366, n67367, n67368, n67369, n67370,
    n67371, n67372, n67373, n67374, n67375, n67376, n67378, n67379, n67380,
    n67381, n67382, n67383, n67384, n67385, n67386, n67387, n67388, n67389,
    n67390, n67391, n67392, n67393, n67394, n67395, n67396, n67397, n67398,
    n67399, n67400, n67401, n67402, n67403, n67404, n67405, n67407, n67408,
    n67409, n67410, n67411, n67412, n67413, n67414, n67415, n67416, n67417,
    n67418, n67419, n67420, n67421, n67422, n67423, n67424, n67425, n67426,
    n67427, n67428, n67429, n67430, n67431, n67432, n67433, n67434, n67435,
    n67436, n67437, n67438, n67439, n67440, n67441, n67442, n67443, n67444,
    n67445, n67447, n67448, n67449, n67450, n67451, n67452, n67453, n67454,
    n67455, n67456, n67457, n67458, n67459, n67460, n67461, n67462, n67463,
    n67464, n67465, n67466, n67467, n67468, n67469, n67470, n67471, n67472,
    n67473, n67474, n67475, n67477, n67478, n67479, n67480, n67481, n67482,
    n67483, n67484, n67485, n67486, n67487, n67488, n67489, n67490, n67491,
    n67492, n67493, n67494, n67495, n67496, n67497, n67498, n67499, n67500,
    n67501, n67502, n67503, n67504, n67505, n67506, n67507, n67508, n67509,
    n67510, n67511, n67512, n67513, n67514, n67515, n67516, n67517, n67518,
    n67519, n67520, n67521, n67522, n67523, n67524, n67525, n67526, n67528,
    n67529, n67530, n67531, n67532, n67533, n67534, n67535, n67536, n67537,
    n67538, n67539, n67540, n67541, n67542, n67543, n67544, n67545, n67546,
    n67547, n67548, n67549, n67550, n67551, n67552, n67553, n67554, n67555,
    n67556, n67557, n67558, n67559, n67560, n67561, n67562, n67563, n67564,
    n67566, n67567, n67568, n67569, n67570, n67571, n67572, n67573, n67574,
    n67575, n67576, n67577, n67578, n67579, n67580, n67581, n67582, n67583,
    n67584, n67585, n67586, n67587, n67588, n67589, n67590, n67591, n67592,
    n67593, n67594, n67595, n67596, n67597, n67598, n67599, n67600, n67601,
    n67603, n67604, n67605, n67606, n67607, n67608, n67609, n67610, n67611,
    n67612, n67613, n67614, n67615, n67616, n67617, n67618, n67619, n67620,
    n67621, n67622, n67623, n67624, n67625, n67626, n67627, n67628, n67629,
    n67630, n67631, n67632, n67633, n67634, n67635, n67636, n67637, n67638,
    n67639, n67640, n67641, n67642, n67643, n67644, n67645, n67646, n67647,
    n67648, n67649, n67650, n67651, n67652, n67653, n67654, n67655, n67656,
    n67657, n67658, n67659, n67660, n67661, n67662, n67663, n67664, n67665,
    n67666, n67667, n67668, n67669, n67670, n67671, n67672, n67673, n67674,
    n67675, n67676, n67677, n67678, n67679, n67680, n67681, n67682, n67683,
    n67684, n67685, n67686, n67687, n67688, n67690, n67691, n67692, n67693,
    n67694, n67695, n67696, n67697, n67698, n67699, n67700, n67701, n67702,
    n67703, n67704, n67705, n67706, n67707, n67708, n67709, n67710, n67711,
    n67712, n67713, n67714, n67716, n67717, n67718, n67719, n67720, n67721,
    n67722, n67723, n67724, n67725, n67726, n67727, n67728, n67729, n67730,
    n67731, n67732, n67733, n67734, n67735, n67736, n67737, n67738, n67739,
    n67740, n67741, n67742, n67743, n67744, n67745, n67746, n67747, n67749,
    n67750, n67751, n67752, n67753, n67754, n67755, n67756, n67757, n67758,
    n67759, n67760, n67761, n67762, n67763, n67764, n67765, n67766, n67767,
    n67768, n67769, n67770, n67771, n67772, n67773, n67774, n67775, n67776,
    n67777, n67778, n67779, n67780, n67781, n67782, n67783, n67784, n67785,
    n67786, n67787, n67788, n67789, n67790, n67791, n67792, n67793, n67794,
    n67795, n67796, n67797, n67798, n67799, n67800, n67802, n67803, n67804,
    n67805, n67806, n67807, n67808, n67809, n67810, n67811, n67812, n67813,
    n67814, n67815, n67816, n67817, n67818, n67819, n67820, n67821, n67822,
    n67823, n67824, n67825, n67826, n67827, n67828, n67829, n67830, n67831,
    n67832, n67833, n67834, n67835, n67836, n67837, n67838, n67839, n67841,
    n67842, n67843, n67844, n67845, n67846, n67847, n67848, n67849, n67850,
    n67851, n67852, n67853, n67854, n67855, n67856, n67857, n67858, n67859,
    n67860, n67861, n67862, n67863, n67864, n67865, n67866, n67867, n67868,
    n67869, n67870, n67871, n67872, n67873, n67875, n67876, n67877, n67878,
    n67879, n67880, n67881, n67882, n67883, n67884, n67885, n67886, n67887,
    n67888, n67889, n67890, n67891, n67892, n67893, n67894, n67895, n67896,
    n67897, n67898, n67899, n67900, n67901, n67902, n67903, n67904, n67905,
    n67906, n67907, n67908, n67909, n67910, n67911, n67912, n67913, n67914,
    n67915, n67916, n67917, n67918, n67919, n67920, n67921, n67922, n67923,
    n67924, n67925, n67926, n67927, n67928, n67929, n67930, n67931, n67932,
    n67933, n67934, n67935, n67936, n67937, n67938, n67939, n67940, n67941,
    n67942, n67943, n67944, n67945, n67946, n67947, n67948, n67949, n67950,
    n67951, n67952, n67953, n67954, n67955, n67956, n67957, n67958, n67959,
    n67960, n67961, n67962, n67963, n67964, n67965, n67966, n67967, n67968,
    n67969, n67970, n67971, n67972, n67973, n67975, n67976, n67977, n67978,
    n67979, n67980, n67981, n67982, n67983, n67984, n67985, n67986, n67987,
    n67988, n67989, n67990, n67991, n67992, n67993, n67994, n67995, n67996,
    n67997, n67998, n67999, n68000, n68001, n68002, n68003, n68004, n68005,
    n68006, n68007, n68008, n68009, n68010, n68011, n68012, n68013, n68014,
    n68015, n68016, n68017, n68018, n68019, n68020, n68021, n68022, n68023,
    n68024, n68025, n68026, n68027, n68028, n68029, n68030, n68031, n68032,
    n68033, n68034, n68035, n68036, n68037, n68038, n68039, n68040, n68041,
    n68042, n68043, n68044, n68045, n68046, n68047, n68048, n68049, n68050,
    n68051, n68052, n68053, n68054, n68055, n68056, n68057, n68058, n68059,
    n68060, n68061, n68062, n68063, n68064, n68065, n68066, n68067, n68068,
    n68069, n68070, n68071, n68072, n68073, n68074, n68075, n68077, n68078,
    n68079, n68080, n68081, n68082, n68083, n68084, n68085, n68086, n68087,
    n68088, n68089, n68090, n68091, n68092, n68093, n68094, n68095, n68096,
    n68097, n68098, n68099, n68100, n68101, n68102, n68103, n68104, n68105,
    n68106, n68107, n68108, n68109, n68110, n68111, n68112, n68113, n68114,
    n68115, n68116, n68117, n68118, n68119, n68120, n68121, n68122, n68123,
    n68124, n68125, n68126, n68127, n68128, n68129, n68130, n68131, n68132,
    n68133, n68134, n68135, n68136, n68137, n68138, n68139, n68140, n68141,
    n68142, n68143, n68144, n68145, n68146, n68147, n68148, n68149, n68150,
    n68151, n68152, n68153, n68154, n68155, n68156, n68157, n68158, n68159,
    n68160, n68161, n68162, n68163, n68164, n68165, n68166, n68167, n68168,
    n68169, n68170, n68171, n68172, n68173, n68174, n68175, n68176, n68177,
    n68178, n68179, n68180, n68182, n68183, n68184, n68185, n68186, n68187,
    n68188, n68189, n68190, n68191, n68192, n68193, n68194, n68195, n68196,
    n68197, n68198, n68199, n68200, n68201, n68202, n68203, n68204, n68205,
    n68206, n68207, n68208, n68209, n68210, n68211, n68212, n68213, n68214,
    n68215, n68216, n68217, n68218, n68219, n68220, n68221, n68222, n68223,
    n68225, n68226, n68227, n68228, n68229, n68230, n68231, n68232, n68233,
    n68234, n68235, n68236, n68237, n68238, n68239, n68240, n68241, n68242,
    n68243, n68244, n68245, n68246, n68247, n68248, n68249, n68250, n68251,
    n68252, n68253, n68254, n68255, n68256, n68258, n68259, n68260, n68261,
    n68262, n68263, n68264, n68265, n68266, n68267, n68268, n68269, n68270,
    n68271, n68272, n68273, n68274, n68275, n68276, n68277, n68278, n68279,
    n68280, n68281, n68282, n68283, n68284, n68285, n68286, n68287, n68288,
    n68289, n68290, n68291, n68292, n68293, n68294, n68295, n68296, n68297,
    n68298, n68299, n68300, n68301, n68302, n68303, n68304, n68305, n68306,
    n68307, n68308, n68309, n68310, n68311, n68312, n68313, n68314, n68315,
    n68316, n68317, n68318, n68319, n68320, n68321, n68322, n68323, n68324,
    n68325, n68326, n68327, n68328, n68329, n68330, n68331, n68332, n68333,
    n68334, n68335, n68336, n68337, n68338, n68339, n68340, n68341, n68342,
    n68343, n68344, n68345, n68346, n68347, n68348, n68349, n68350, n68351,
    n68352, n68353, n68354, n68355, n68356, n68358, n68359, n68360, n68361,
    n68362, n68363, n68364, n68365, n68366, n68367, n68368, n68369, n68370,
    n68371, n68372, n68373, n68374, n68375, n68376, n68377, n68378, n68379,
    n68380, n68381, n68382, n68383, n68384, n68385, n68386, n68387, n68388,
    n68389, n68390, n68391, n68392, n68393, n68394, n68395, n68396, n68397,
    n68398, n68399, n68400, n68401, n68402, n68403, n68404, n68405, n68406,
    n68407, n68408, n68409, n68410, n68411, n68412, n68413, n68414, n68415,
    n68416, n68417, n68418, n68419, n68420, n68421, n68422, n68423, n68424,
    n68425, n68426, n68427, n68428, n68429, n68430, n68431, n68432, n68433,
    n68434, n68435, n68436, n68437, n68438, n68439, n68440, n68441, n68442,
    n68443, n68444, n68445, n68446, n68447, n68448, n68449, n68450, n68451,
    n68452, n68453, n68454, n68455, n68456, n68457, n68458, n68460, n68461,
    n68462, n68463, n68464, n68465, n68466, n68467, n68468, n68469, n68470,
    n68471, n68472, n68473, n68474, n68475, n68476, n68477, n68478, n68479,
    n68480, n68481, n68482, n68483, n68484, n68485, n68486, n68487, n68488,
    n68489, n68490, n68491, n68492, n68493, n68494, n68495, n68496, n68497,
    n68498, n68499, n68500, n68501, n68502, n68503, n68504, n68505, n68506,
    n68507, n68508, n68509, n68510, n68511, n68512, n68513, n68514, n68515,
    n68516, n68517, n68518, n68519, n68520, n68521, n68522, n68523, n68524,
    n68525, n68526, n68527, n68528, n68529, n68530, n68531, n68532, n68533,
    n68534, n68535, n68536, n68537, n68538, n68539, n68540, n68541, n68542,
    n68543, n68544, n68545, n68546, n68547, n68548, n68549, n68550, n68551,
    n68552, n68553, n68554, n68555, n68556, n68557, n68558, n68559, n68560,
    n68561, n68562, n68563, n68564, n68565, n68567, n68568, n68569, n68570,
    n68571, n68572, n68573, n68574, n68575, n68576, n68577, n68578, n68579,
    n68580, n68581, n68582, n68583, n68584, n68585, n68586, n68587, n68588,
    n68589, n68590, n68591, n68592, n68593, n68594, n68595, n68596, n68597,
    n68598, n68599, n68600, n68601, n68602, n68603, n68604, n68605, n68606,
    n68607, n68608, n68609, n68610, n68611, n68613, n68614, n68615, n68616,
    n68617, n68618, n68619, n68620, n68621, n68622, n68623, n68624, n68625,
    n68626, n68627, n68628, n68629, n68630, n68631, n68632, n68633, n68634,
    n68635, n68636, n68637, n68638, n68639, n68640, n68641, n68642, n68643,
    n68644, n68645, n68646, n68647, n68648, n68650, n68651, n68652, n68653,
    n68654, n68655, n68656, n68657, n68658, n68659, n68660, n68661, n68662,
    n68663, n68664, n68665, n68666, n68667, n68668, n68669, n68670, n68671,
    n68672, n68673, n68674, n68675, n68676, n68677, n68678, n68679, n68680,
    n68681, n68682, n68683, n68684, n68685, n68686, n68687, n68688, n68689,
    n68690, n68691, n68692, n68693, n68694, n68695, n68696, n68697, n68698,
    n68699, n68700, n68701, n68702, n68703, n68704, n68705, n68706, n68707,
    n68708, n68709, n68710, n68711, n68712, n68713, n68714, n68715, n68716,
    n68717, n68718, n68719, n68720, n68721, n68722, n68723, n68724, n68725,
    n68726, n68727, n68728, n68729, n68730, n68731, n68732, n68733, n68734,
    n68735, n68736, n68737, n68738, n68739, n68741, n68742, n68743, n68744,
    n68745, n68746, n68747, n68748, n68749, n68750, n68751, n68752, n68753,
    n68754, n68755, n68756, n68757, n68758, n68759, n68760, n68761, n68762,
    n68763, n68764, n68765, n68766, n68767, n68768, n68769, n68770, n68771,
    n68772, n68773, n68774, n68776, n68777, n68778, n68779, n68780, n68781,
    n68782, n68783, n68784, n68785, n68786, n68787, n68788, n68789, n68790,
    n68791, n68792, n68793, n68794, n68795, n68796, n68797, n68798, n68799,
    n68800, n68801, n68802, n68803, n68804, n68805, n68806, n68807, n68808,
    n68809, n68810, n68811, n68812, n68813, n68814, n68815, n68816, n68817,
    n68818, n68819, n68820, n68821, n68822, n68824, n68825, n68826, n68827,
    n68828, n68829, n68830, n68831, n68832, n68833, n68834, n68835, n68836,
    n68837, n68838, n68839, n68840, n68841, n68842, n68843, n68844, n68845,
    n68846, n68847, n68848, n68849, n68850, n68851, n68852, n68853, n68854,
    n68855, n68856, n68857, n68858, n68859, n68861, n68862, n68863, n68864,
    n68865, n68866, n68867, n68868, n68869, n68870, n68871, n68872, n68873,
    n68874, n68875, n68876, n68877, n68878, n68879, n68880, n68881, n68882,
    n68883, n68884, n68885, n68886, n68887, n68888, n68889, n68890, n68891,
    n68892, n68893, n68894, n68895, n68896, n68897, n68898, n68899, n68901,
    n68902, n68903, n68904, n68905, n68906, n68907, n68908, n68909, n68910,
    n68911, n68912, n68913, n68914, n68915, n68916, n68917, n68918, n68919,
    n68920, n68921, n68922, n68923, n68924, n68925, n68926, n68927, n68928,
    n68929, n68930, n68931, n68932, n68933, n68934, n68935, n68936, n68937,
    n68938, n68939, n68940, n68942, n68943, n68944, n68945, n68946, n68947,
    n68948, n68949, n68950, n68951, n68952, n68953, n68954, n68955, n68956,
    n68957, n68958, n68959, n68960, n68961, n68962, n68963, n68964, n68965,
    n68966, n68967, n68968, n68969, n68970, n68972, n68973, n68974, n68975,
    n68976, n68977, n68978, n68979, n68980, n68981, n68982, n68983, n68984,
    n68985, n68986, n68987, n68988, n68989, n68990, n68991, n68992, n68993,
    n68994, n68995, n68996, n68997, n68998, n68999, n69000, n69001, n69002,
    n69003, n69004, n69005, n69006, n69007, n69008, n69009, n69010, n69012,
    n69013, n69014, n69015, n69016, n69017, n69018, n69019, n69020, n69021,
    n69022, n69023, n69024, n69025, n69026, n69027, n69028, n69029, n69030,
    n69031, n69032, n69033, n69034, n69035, n69036, n69037, n69038, n69039,
    n69040, n69041, n69042, n69043, n69044, n69045, n69046, n69047, n69049,
    n69050, n69051, n69052, n69053, n69054, n69055, n69056, n69057, n69058,
    n69059, n69060, n69061, n69062, n69063, n69064, n69065, n69066, n69067,
    n69068, n69069, n69070, n69071, n69072, n69073, n69074, n69075, n69076,
    n69077, n69078, n69079, n69080, n69081, n69082, n69083, n69084, n69085,
    n69086, n69087, n69088, n69089, n69090, n69091, n69092, n69093, n69094,
    n69095, n69096, n69097, n69098, n69099, n69100, n69101, n69102, n69103,
    n69104, n69105, n69106, n69107, n69108, n69109, n69110, n69111, n69112,
    n69113, n69114, n69115, n69116, n69117, n69118, n69119, n69120, n69121,
    n69122, n69123, n69124, n69125, n69126, n69127, n69128, n69129, n69130,
    n69131, n69132, n69133, n69134, n69135, n69136, n69137, n69138, n69139,
    n69140, n69141, n69142, n69143, n69144, n69145, n69147, n69148, n69149,
    n69150, n69151, n69152, n69153, n69154, n69155, n69156, n69157, n69158,
    n69159, n69160, n69161, n69162, n69163, n69164, n69165, n69166, n69167,
    n69168, n69169, n69170, n69171, n69172, n69173, n69174, n69175, n69176,
    n69177, n69178, n69179, n69180, n69181, n69182, n69183, n69184, n69186,
    n69187, n69188, n69189, n69190, n69191, n69192, n69193, n69194, n69195,
    n69196, n69197, n69198, n69199, n69200, n69201, n69202, n69203, n69204,
    n69205, n69206, n69207, n69208, n69209, n69210, n69211, n69212, n69213,
    n69214, n69215, n69216, n69217, n69218, n69219, n69220, n69221, n69222,
    n69223, n69224, n69225, n69226, n69227, n69228, n69229, n69230, n69231,
    n69232, n69233, n69234, n69236, n69237, n69238, n69239, n69240, n69241,
    n69242, n69243, n69244, n69245, n69246, n69247, n69248, n69249, n69250,
    n69251, n69252, n69253, n69254, n69255, n69256, n69257, n69258, n69259,
    n69260, n69261, n69262, n69263, n69264, n69265, n69266, n69267, n69268,
    n69269, n69270, n69271, n69272, n69273, n69274, n69275, n69276, n69277,
    n69278, n69279, n69280, n69282, n69283, n69284, n69285, n69286, n69287,
    n69288, n69289, n69290, n69291, n69292, n69293, n69294, n69295, n69296,
    n69297, n69298, n69299, n69300, n69301, n69302, n69303, n69304, n69305,
    n69306, n69307, n69308, n69309, n69310, n69311, n69312, n69313, n69314,
    n69315, n69317, n69318, n69319, n69320, n69321, n69322, n69323, n69324,
    n69325, n69326, n69327, n69328, n69329, n69330, n69331, n69332, n69333,
    n69334, n69335, n69336, n69337, n69338, n69339, n69340, n69341, n69342,
    n69343, n69344, n69345, n69346, n69347, n69348, n69349, n69350, n69351,
    n69352, n69353, n69355, n69356, n69357, n69358, n69359, n69360, n69361,
    n69362, n69363, n69364, n69365, n69366, n69367, n69368, n69369, n69370,
    n69371, n69372, n69373, n69374, n69375, n69376, n69377, n69378, n69379,
    n69380, n69381, n69382, n69383, n69384, n69385, n69386, n69388, n69389,
    n69390, n69391, n69392, n69393, n69394, n69395, n69396, n69397, n69398,
    n69399, n69400, n69401, n69402, n69403, n69404, n69405, n69406, n69407,
    n69408, n69409, n69410, n69411, n69412, n69413, n69414, n69415, n69416,
    n69417, n69418, n69419, n69420, n69421, n69422, n69423, n69424, n69425,
    n69426, n69428, n69429, n69430, n69431, n69432, n69433, n69434, n69435,
    n69436, n69437, n69438, n69439, n69440, n69441, n69442, n69443, n69444,
    n69445, n69446, n69447, n69448, n69449, n69450, n69451, n69452, n69453,
    n69454, n69455, n69456, n69458, n69459, n69460, n69461, n69462, n69463,
    n69464, n69465, n69466, n69467, n69468, n69469, n69470, n69471, n69472,
    n69473, n69474, n69475, n69476, n69477, n69478, n69479, n69480, n69481,
    n69482, n69483, n69484, n69485, n69486, n69487, n69488, n69489, n69490,
    n69491, n69492, n69494, n69495, n69496, n69497, n69498, n69499, n69500,
    n69501, n69502, n69503, n69504, n69505, n69506, n69507, n69508, n69509,
    n69510, n69511, n69512, n69513, n69514, n69515, n69516, n69517, n69518,
    n69519, n69520, n69521, n69522, n69523, n69524, n69525, n69526, n69527,
    n69528, n69529, n69530, n69531, n69532, n69533, n69535, n69536, n69537,
    n69538, n69539, n69540, n69541, n69542, n69543, n69544, n69545, n69546,
    n69547, n69548, n69549, n69550, n69551, n69552, n69553, n69554, n69555,
    n69556, n69557, n69558, n69559, n69560, n69561, n69562, n69563, n69565,
    n69566, n69567, n69568, n69569, n69570, n69571, n69572, n69573, n69574,
    n69575, n69576, n69577, n69578, n69579, n69580, n69581, n69582, n69583,
    n69584, n69585, n69586, n69587, n69588, n69589, n69591, n69592, n69593,
    n69594, n69595, n69596, n69597, n69598, n69599, n69600, n69601, n69602,
    n69603, n69604, n69605, n69606, n69607, n69608, n69609, n69610, n69611,
    n69612, n69613, n69614, n69615, n69616, n69617, n69618, n69619, n69620,
    n69621, n69622, n69623, n69624, n69625, n69626, n69627, n69628, n69629,
    n69630, n69631, n69632, n69633, n69634, n69635, n69636, n69637, n69638,
    n69639, n69640, n69641, n69642, n69643, n69644, n69645, n69646, n69647,
    n69648, n69649, n69650, n69651, n69652, n69653, n69654, n69655, n69656,
    n69657, n69658, n69659, n69660, n69661, n69662, n69663, n69664, n69665,
    n69666, n69667, n69668, n69669, n69670, n69671, n69672, n69673, n69674,
    n69675, n69676, n69677, n69678, n69679, n69680, n69681, n69682, n69683,
    n69684, n69685, n69686, n69687, n69688, n69689, n69690, n69692, n69693,
    n69694, n69695, n69696, n69697, n69698, n69699, n69700, n69701, n69702,
    n69703, n69704, n69705, n69706, n69707, n69708, n69709, n69710, n69711,
    n69712, n69713, n69714, n69715, n69716, n69717, n69718, n69719, n69720,
    n69721, n69722, n69723, n69724, n69725, n69726, n69727, n69728, n69729,
    n69730, n69731, n69732, n69733, n69734, n69735, n69736, n69737, n69738,
    n69739, n69740, n69741, n69742, n69743, n69744, n69745, n69746, n69747,
    n69748, n69749, n69750, n69751, n69752, n69753, n69754, n69755, n69756,
    n69757, n69758, n69759, n69760, n69761, n69762, n69763, n69764, n69765,
    n69766, n69767, n69768, n69769, n69770, n69771, n69772, n69773, n69774,
    n69775, n69776, n69777, n69778, n69779, n69780, n69781, n69782, n69783,
    n69784, n69785, n69786, n69787, n69788, n69789, n69791, n69792, n69793,
    n69794, n69795, n69796, n69797, n69798, n69799, n69800, n69801, n69802,
    n69803, n69804, n69805, n69806, n69807, n69808, n69809, n69810, n69811,
    n69812, n69813, n69814, n69815, n69816, n69817, n69818, n69819, n69820,
    n69821, n69822, n69823, n69824, n69825, n69826, n69827, n69828, n69829,
    n69830, n69831, n69832, n69833, n69834, n69835, n69836, n69837, n69838,
    n69839, n69840, n69841, n69842, n69843, n69844, n69845, n69846, n69847,
    n69848, n69849, n69850, n69851, n69852, n69853, n69854, n69855, n69856,
    n69857, n69858, n69859, n69860, n69861, n69862, n69863, n69864, n69865,
    n69866, n69867, n69868, n69869, n69870, n69871, n69872, n69873, n69874,
    n69875, n69876, n69877, n69878, n69879, n69880, n69881, n69882, n69883,
    n69884, n69885, n69886, n69887, n69888, n69889, n69890, n69891, n69892,
    n69893, n69894, n69896, n69897, n69898, n69899, n69900, n69901, n69902,
    n69903, n69904, n69905, n69906, n69907, n69908, n69909, n69910, n69911,
    n69912, n69913, n69914, n69915, n69916, n69917, n69918, n69919, n69920,
    n69921, n69922, n69923, n69924, n69925, n69926, n69927, n69928, n69929,
    n69930, n69931, n69932, n69933, n69934, n69935, n69936, n69937, n69938,
    n69939, n69940, n69942, n69943, n69944, n69945, n69946, n69947, n69948,
    n69949, n69950, n69951, n69952, n69953, n69954, n69955, n69956, n69957,
    n69958, n69959, n69960, n69961, n69962, n69963, n69964, n69965, n69966,
    n69967, n69968, n69969, n69970, n69971, n69972, n69974, n69975, n69976,
    n69977, n69978, n69979, n69980, n69981, n69982, n69983, n69984, n69985,
    n69986, n69987, n69988, n69989, n69990, n69991, n69992, n69993, n69994,
    n69995, n69996, n69997, n69998, n69999, n70000, n70001, n70002, n70003,
    n70004, n70005, n70006, n70007, n70008, n70009, n70010, n70011, n70012,
    n70013, n70014, n70015, n70016, n70017, n70018, n70019, n70020, n70021,
    n70022, n70023, n70024, n70025, n70026, n70027, n70028, n70029, n70030,
    n70031, n70032, n70033, n70034, n70035, n70036, n70037, n70038, n70039,
    n70040, n70041, n70042, n70043, n70044, n70045, n70046, n70047, n70048,
    n70049, n70050, n70051, n70052, n70053, n70054, n70055, n70056, n70057,
    n70058, n70059, n70060, n70061, n70062, n70063, n70064, n70065, n70066,
    n70067, n70068, n70069, n70070, n70071, n70072, n70073, n70074, n70075,
    n70077, n70078, n70079, n70080, n70081, n70082, n70083, n70084, n70085,
    n70086, n70087, n70088, n70089, n70090, n70091, n70092, n70093, n70094,
    n70095, n70096, n70097, n70098, n70099, n70100, n70101, n70102, n70103,
    n70104, n70105, n70106, n70107, n70108, n70109, n70110, n70111, n70112,
    n70113, n70114, n70115, n70116, n70117, n70118, n70119, n70120, n70121,
    n70122, n70123, n70124, n70126, n70127, n70128, n70129, n70130, n70131,
    n70132, n70133, n70134, n70135, n70136, n70137, n70138, n70139, n70140,
    n70141, n70142, n70143, n70144, n70145, n70146, n70147, n70148, n70149,
    n70150, n70151, n70152, n70153, n70154, n70155, n70156, n70157, n70158,
    n70159, n70160, n70161, n70162, n70163, n70164, n70165, n70166, n70167,
    n70168, n70169, n70170, n70171, n70172, n70173, n70174, n70175, n70176,
    n70177, n70178, n70179, n70180, n70181, n70182, n70183, n70184, n70185,
    n70186, n70187, n70188, n70189, n70190, n70191, n70192, n70193, n70194,
    n70195, n70196, n70197, n70198, n70199, n70200, n70201, n70202, n70203,
    n70204, n70205, n70206, n70207, n70208, n70209, n70210, n70211, n70212,
    n70213, n70214, n70215, n70216, n70217, n70218, n70219, n70220, n70221,
    n70222, n70223, n70224, n70225, n70226, n70227, n70228, n70229, n70230,
    n70231, n70233, n70234, n70235, n70236, n70237, n70238, n70239, n70240,
    n70241, n70242, n70243, n70244, n70245, n70246, n70247, n70248, n70249,
    n70250, n70251, n70252, n70253, n70254, n70255, n70256, n70257, n70258,
    n70259, n70260, n70261, n70262, n70263, n70264, n70265, n70266, n70267,
    n70269, n70270, n70271, n70272, n70273, n70274, n70275, n70276, n70277,
    n70278, n70279, n70280, n70281, n70282, n70283, n70284, n70285, n70286,
    n70287, n70288, n70289, n70290, n70291, n70292, n70293, n70294, n70295,
    n70296, n70297, n70298, n70299, n70300, n70302, n70303, n70304, n70305,
    n70306, n70307, n70308, n70309, n70310, n70311, n70312, n70313, n70314,
    n70315, n70316, n70317, n70318, n70319, n70320, n70321, n70322, n70323,
    n70324, n70325, n70326, n70327, n70328, n70329, n70330, n70331, n70332,
    n70333, n70334, n70335, n70336, n70337, n70338, n70339, n70340, n70341,
    n70342, n70343, n70344, n70345, n70346, n70347, n70348, n70349, n70350,
    n70351, n70352, n70353, n70354, n70355, n70356, n70357, n70358, n70359,
    n70360, n70361, n70362, n70363, n70364, n70365, n70366, n70367, n70368,
    n70369, n70370, n70371, n70372, n70373, n70374, n70375, n70376, n70377,
    n70378, n70379, n70380, n70381, n70382, n70383, n70384, n70385, n70386,
    n70387, n70388, n70389, n70390, n70391, n70393, n70394, n70395, n70396,
    n70397, n70398, n70399, n70400, n70401, n70402, n70403, n70404, n70405,
    n70406, n70407, n70408, n70409, n70410, n70411, n70412, n70413, n70414,
    n70415, n70416, n70417, n70418, n70419, n70420, n70421, n70422, n70423,
    n70424, n70425, n70426, n70427, n70428, n70429, n70430, n70431, n70432,
    n70434, n70435, n70436, n70437, n70438, n70439, n70440, n70441, n70442,
    n70443, n70444, n70445, n70446, n70447, n70448, n70449, n70450, n70451,
    n70452, n70453, n70454, n70455, n70456, n70457, n70458, n70459, n70460,
    n70461, n70462, n70463, n70464, n70465, n70466, n70468, n70469, n70470,
    n70471, n70472, n70473, n70474, n70475, n70476, n70477, n70478, n70479,
    n70480, n70481, n70482, n70483, n70484, n70485, n70486, n70487, n70488,
    n70489, n70490, n70491, n70492, n70493, n70494, n70495, n70496, n70497,
    n70499, n70500, n70501, n70502, n70503, n70504, n70505, n70506, n70507,
    n70508, n70509, n70510, n70511, n70512, n70513, n70514, n70515, n70516,
    n70517, n70518, n70519, n70520, n70521, n70522, n70523, n70524, n70525,
    n70526, n70527, n70528, n70529, n70530, n70531, n70532, n70533, n70534,
    n70535, n70536, n70537, n70538, n70539, n70540, n70541, n70542, n70543,
    n70544, n70545, n70546, n70547, n70549, n70550, n70551, n70552, n70553,
    n70554, n70555, n70556, n70557, n70558, n70559, n70560, n70561, n70562,
    n70563, n70564, n70565, n70566, n70567, n70568, n70569, n70570, n70571,
    n70572, n70573, n70574, n70575, n70576, n70577, n70578, n70579, n70580,
    n70581, n70582, n70583, n70584, n70585, n70586, n70587, n70588, n70589,
    n70590, n70591, n70592, n70593, n70594, n70595, n70596, n70597, n70598,
    n70599, n70600, n70601, n70602, n70603, n70604, n70605, n70606, n70607,
    n70608, n70609, n70610, n70611, n70612, n70613, n70614, n70615, n70616,
    n70617, n70618, n70619, n70620, n70621, n70622, n70623, n70624, n70625,
    n70626, n70627, n70628, n70629, n70630, n70631, n70632, n70633, n70634,
    n70635, n70636, n70637, n70638, n70639, n70640, n70641, n70642, n70643,
    n70644, n70645, n70646, n70648, n70649, n70650, n70651, n70652, n70653,
    n70654, n70655, n70656, n70657, n70658, n70659, n70660, n70661, n70662,
    n70663, n70664, n70665, n70666, n70667, n70668, n70669, n70670, n70671,
    n70672, n70673, n70674, n70675, n70676, n70677, n70678, n70679, n70680,
    n70681, n70682, n70683, n70684, n70685, n70686, n70687, n70689, n70690,
    n70691, n70692, n70693, n70694, n70695, n70696, n70697, n70698, n70699,
    n70700, n70701, n70702, n70703, n70704, n70705, n70706, n70707, n70708,
    n70709, n70710, n70711, n70712, n70713, n70714, n70715, n70716, n70717,
    n70718, n70719, n70720, n70721, n70722, n70723, n70724, n70725, n70726,
    n70727, n70728, n70729, n70730, n70731, n70732, n70734, n70735, n70736,
    n70737, n70738, n70739, n70740, n70741, n70742, n70743, n70744, n70745,
    n70746, n70747, n70748, n70749, n70750, n70751, n70752, n70753, n70754,
    n70755, n70756, n70757, n70758, n70759, n70760, n70761, n70762, n70763,
    n70764, n70765, n70766, n70767, n70768, n70769, n70770, n70772, n70773,
    n70774, n70775, n70776, n70777, n70778, n70779, n70780, n70781, n70782,
    n70783, n70784, n70785, n70786, n70787, n70788, n70789, n70790, n70791,
    n70792, n70793, n70794, n70795, n70796, n70797, n70798, n70799, n70800,
    n70801, n70802, n70803, n70804, n70805, n70807, n70808, n70809, n70810,
    n70811, n70812, n70813, n70814, n70815, n70816, n70817, n70818, n70819,
    n70820, n70821, n70822, n70823, n70824, n70825, n70826, n70827, n70828,
    n70829, n70830, n70831, n70832, n70833, n70834, n70835, n70836, n70837,
    n70838, n70839, n70840, n70841, n70842, n70843, n70844, n70845, n70846,
    n70847, n70848, n70849, n70850, n70851, n70852, n70853, n70854, n70855,
    n70856, n70857, n70858, n70859, n70860, n70861, n70862, n70863, n70864,
    n70865, n70866, n70867, n70868, n70869, n70870, n70871, n70872, n70873,
    n70874, n70875, n70876, n70877, n70878, n70879, n70880, n70881, n70882,
    n70883, n70884, n70885, n70886, n70887, n70888, n70889, n70890, n70891,
    n70892, n70893, n70894, n70895, n70896, n70897, n70898, n70899, n70900,
    n70901, n70903, n70904, n70905, n70906, n70907, n70908, n70909, n70910,
    n70911, n70912, n70913, n70914, n70915, n70916, n70917, n70918, n70919,
    n70920, n70921, n70922, n70923, n70924, n70925, n70926, n70927, n70928,
    n70929, n70930, n70931, n70932, n70933, n70934, n70935, n70936, n70937,
    n70938, n70939, n70940, n70941, n70943, n70944, n70945, n70946, n70947,
    n70948, n70949, n70950, n70951, n70952, n70953, n70954, n70955, n70956,
    n70957, n70958, n70959, n70960, n70961, n70962, n70963, n70964, n70965,
    n70966, n70967, n70968, n70969, n70970, n70971, n70972, n70973, n70974,
    n70975, n70976, n70977, n70978, n70979, n70980, n70981, n70982, n70983,
    n70984, n70985, n70986, n70988, n70989, n70990, n70991, n70992, n70993,
    n70994, n70995, n70996, n70997, n70998, n70999, n71000, n71001, n71002,
    n71003, n71004, n71005, n71006, n71007, n71008, n71009, n71010, n71011,
    n71012, n71013, n71014, n71015, n71016, n71018, n71019, n71020, n71021,
    n71022, n71023, n71024, n71025, n71026, n71027, n71028, n71029, n71030,
    n71031, n71032, n71033, n71034, n71035, n71036, n71037, n71038, n71039,
    n71040, n71041, n71042, n71043, n71044, n71045, n71046, n71047, n71048,
    n71049, n71050, n71051, n71053, n71054, n71055, n71056, n71057, n71058,
    n71059, n71060, n71061, n71062, n71063, n71064, n71065, n71066, n71067,
    n71068, n71069, n71070, n71071, n71072, n71073, n71074, n71075, n71076,
    n71077, n71078, n71079, n71080, n71081, n71082, n71083, n71084, n71085,
    n71086, n71087, n71088, n71089, n71090, n71091, n71092, n71094, n71095,
    n71096, n71097, n71098, n71099, n71100, n71101, n71102, n71103, n71104,
    n71105, n71106, n71107, n71108, n71109, n71110, n71111, n71112, n71113,
    n71114, n71115, n71116, n71117, n71118, n71119, n71120, n71121, n71122,
    n71123, n71124, n71125, n71126, n71127, n71128, n71129, n71130, n71131,
    n71132, n71133, n71134, n71135, n71136, n71137, n71138, n71139, n71140,
    n71142, n71143, n71144, n71145, n71146, n71147, n71148, n71149, n71150,
    n71151, n71152, n71153, n71154, n71155, n71156, n71157, n71158, n71159,
    n71160, n71161, n71162, n71163, n71164, n71165, n71166, n71167, n71168,
    n71169, n71170, n71171, n71172, n71173, n71174, n71175, n71176, n71177,
    n71178, n71179, n71181, n71182, n71183, n71184, n71185, n71186, n71187,
    n71188, n71189, n71190, n71191, n71192, n71193, n71194, n71195, n71196,
    n71197, n71198, n71199, n71200, n71201, n71202, n71203, n71204, n71205,
    n71206, n71207, n71208, n71209, n71210, n71211, n71212, n71213, n71214,
    n71216, n71217, n71218, n71219, n71220, n71221, n71222, n71223, n71224,
    n71225, n71226, n71227, n71228, n71229, n71230, n71231, n71232, n71233,
    n71234, n71235, n71236, n71237, n71238, n71239, n71240, n71241, n71242,
    n71243, n71244, n71245, n71246, n71247, n71248, n71249, n71250, n71251,
    n71253, n71254, n71255, n71256, n71257, n71258, n71259, n71260, n71261,
    n71262, n71263, n71264, n71265, n71266, n71267, n71268, n71269, n71270,
    n71271, n71272, n71273, n71274, n71275, n71276, n71277, n71279, n71280,
    n71281, n71282, n71283, n71284, n71285, n71286, n71287, n71288, n71289,
    n71290, n71291, n71292, n71293, n71294, n71295, n71296, n71297, n71298,
    n71299, n71300, n71301, n71302, n71303, n71304, n71305, n71306, n71307,
    n71308, n71309, n71310, n71312, n71313, n71314, n71315, n71316, n71317,
    n71318, n71319, n71320, n71321, n71322, n71323, n71324, n71325, n71326,
    n71327, n71328, n71329, n71330, n71331, n71332, n71333, n71334, n71335,
    n71336, n71337, n71338, n71339, n71340, n71341, n71342, n71343, n71344,
    n71345, n71346, n71347, n71348, n71349, n71350, n71351, n71352, n71353,
    n71354, n71355, n71356, n71357, n71358, n71359, n71360, n71361, n71362,
    n71363, n71364, n71365, n71366, n71367, n71368, n71369, n71370, n71371,
    n71372, n71373, n71374, n71375, n71376, n71377, n71378, n71379, n71380,
    n71381, n71382, n71383, n71384, n71385, n71386, n71387, n71388, n71389,
    n71390, n71391, n71392, n71393, n71394, n71395, n71396, n71397, n71398,
    n71399, n71400, n71401, n71402, n71403, n71404, n71405, n71406, n71407,
    n71408, n71409, n71410, n71411, n71412, n71413, n71414, n71415, n71416,
    n71418, n71419, n71420, n71421, n71422, n71423, n71424, n71425, n71426,
    n71427, n71428, n71429, n71430, n71431, n71432, n71433, n71434, n71435,
    n71436, n71437, n71438, n71439, n71440, n71441, n71442, n71443, n71444,
    n71445, n71446, n71447, n71448, n71449, n71450, n71451, n71452, n71453,
    n71454, n71455, n71456, n71457, n71458, n71459, n71460, n71461, n71462,
    n71463, n71464, n71465, n71466, n71467, n71468, n71469, n71470, n71471,
    n71472, n71473, n71474, n71475, n71476, n71477, n71478, n71479, n71480,
    n71481, n71482, n71483, n71484, n71485, n71486, n71487, n71488, n71489,
    n71490, n71491, n71492, n71493, n71494, n71495, n71496, n71497, n71498,
    n71499, n71500, n71501, n71502, n71503, n71504, n71505, n71506, n71507,
    n71508, n71509, n71510, n71511, n71512, n71513, n71514, n71515, n71517,
    n71518, n71519, n71520, n71521, n71522, n71523, n71524, n71525, n71526,
    n71527, n71528, n71529, n71530, n71531, n71532, n71533, n71534, n71535,
    n71536, n71537, n71538, n71539, n71540, n71541, n71542, n71543, n71544,
    n71545, n71546, n71547, n71548, n71549, n71550, n71551, n71552, n71553,
    n71554, n71555, n71556, n71557, n71558, n71559, n71560, n71562, n71563,
    n71564, n71565, n71566, n71567, n71568, n71569, n71570, n71571, n71572,
    n71573, n71574, n71575, n71576, n71577, n71578, n71579, n71580, n71581,
    n71582, n71583, n71584, n71585, n71586, n71587, n71588, n71589, n71590,
    n71591, n71592, n71593, n71594, n71595, n71596, n71597, n71598, n71599,
    n71600, n71601, n71602, n71603, n71604, n71605, n71606, n71607, n71608,
    n71609, n71610, n71611, n71612, n71613, n71614, n71615, n71616, n71617,
    n71618, n71619, n71620, n71621, n71622, n71623, n71624, n71625, n71626,
    n71627, n71628, n71629, n71630, n71631, n71632, n71633, n71634, n71635,
    n71636, n71637, n71638, n71639, n71640, n71641, n71642, n71643, n71644,
    n71645, n71646, n71647, n71648, n71649, n71650, n71651, n71652, n71653,
    n71654, n71655, n71656, n71657, n71658, n71659, n71660, n71661, n71662,
    n71663, n71664, n71665, n71667, n71668, n71669, n71670, n71671, n71672,
    n71673, n71674, n71675, n71676, n71677, n71678, n71679, n71680, n71681,
    n71682, n71683, n71684, n71685, n71686, n71687, n71688, n71689, n71690,
    n71691, n71692, n71693, n71694, n71695, n71696, n71697, n71698, n71699,
    n71700, n71701, n71702, n71703, n71704, n71705, n71706, n71707, n71708,
    n71709, n71710, n71711, n71712, n71714, n71715, n71716, n71717, n71718,
    n71719, n71720, n71721, n71722, n71723, n71724, n71725, n71726, n71727,
    n71728, n71729, n71730, n71731, n71732, n71733, n71734, n71735, n71736,
    n71737, n71738, n71739, n71740, n71741, n71742, n71743, n71744, n71745,
    n71746, n71747, n71748, n71749, n71750, n71751, n71752, n71753, n71754,
    n71755, n71756, n71757, n71758, n71759, n71760, n71761, n71762, n71763,
    n71764, n71765, n71766, n71767, n71768, n71769, n71770, n71771, n71772,
    n71773, n71774, n71775, n71776, n71777, n71778, n71779, n71780, n71781,
    n71782, n71783, n71784, n71785, n71786, n71787, n71788, n71789, n71790,
    n71791, n71792, n71793, n71794, n71795, n71796, n71797, n71798, n71799,
    n71800, n71801, n71802, n71803, n71804, n71805, n71806, n71807, n71808,
    n71809, n71810, n71811, n71812, n71814, n71815, n71816, n71817, n71818,
    n71819, n71820, n71821, n71822, n71823, n71824, n71825, n71826, n71827,
    n71828, n71829, n71830, n71831, n71832, n71833, n71834, n71835, n71836,
    n71837, n71838, n71839, n71840, n71841, n71842, n71843, n71844, n71845,
    n71846, n71847, n71849, n71850, n71851, n71852, n71853, n71854, n71855,
    n71856, n71857, n71858, n71859, n71860, n71861, n71862, n71863, n71864,
    n71865, n71866, n71867, n71868, n71869, n71870, n71871, n71872, n71873,
    n71874, n71875, n71876, n71877, n71878, n71879, n71880, n71881, n71882,
    n71883, n71884, n71885, n71886, n71887, n71888, n71889, n71890, n71891,
    n71892, n71893, n71894, n71895, n71896, n71898, n71899, n71900, n71901,
    n71902, n71903, n71904, n71905, n71906, n71907, n71908, n71909, n71910,
    n71911, n71912, n71913, n71914, n71915, n71916, n71917, n71918, n71919,
    n71920, n71921, n71922, n71923, n71924, n71925, n71926, n71927, n71928,
    n71929, n71930, n71931, n71933, n71934, n71935, n71936, n71937, n71938,
    n71939, n71940, n71941, n71942, n71943, n71944, n71945, n71946, n71947,
    n71948, n71949, n71950, n71951, n71952, n71953, n71954, n71955, n71956,
    n71957, n71958, n71959, n71960, n71961, n71962, n71963, n71964, n71965,
    n71966, n71967, n71968, n71969, n71970, n71971, n71972, n71973, n71974,
    n71975, n71976, n71977, n71978, n71979, n71980, n71981, n71982, n71983,
    n71984, n71985, n71986, n71987, n71988, n71989, n71990, n71991, n71992,
    n71993, n71994, n71995, n71996, n71997, n71998, n71999, n72000, n72001,
    n72002, n72003, n72004, n72005, n72006, n72007, n72008, n72009, n72010,
    n72011, n72012, n72013, n72014, n72015, n72016, n72017, n72018, n72019,
    n72020, n72021, n72023, n72024, n72025, n72026, n72027, n72028, n72029,
    n72030, n72031, n72032, n72033, n72034, n72035, n72036, n72037, n72038,
    n72039, n72040, n72041, n72042, n72043, n72044, n72045, n72046, n72047,
    n72048, n72049, n72050, n72052, n72053, n72054, n72055, n72056, n72057,
    n72058, n72059, n72060, n72061, n72062, n72063, n72064, n72065, n72066,
    n72067, n72068, n72069, n72070, n72071, n72072, n72073, n72074, n72075,
    n72076, n72077, n72078, n72079, n72080, n72081, n72082, n72083, n72084,
    n72085, n72086, n72087, n72089, n72090, n72091, n72092, n72093, n72094,
    n72095, n72096, n72097, n72098, n72099, n72100, n72101, n72102, n72103,
    n72104, n72105, n72106, n72107, n72108, n72109, n72110, n72111, n72112,
    n72113, n72114, n72115, n72116, n72117, n72118, n72119, n72120, n72121,
    n72122, n72123, n72124, n72125, n72126, n72127, n72128, n72129, n72130,
    n72131, n72132, n72133, n72134, n72135, n72136, n72137, n72138, n72140,
    n72141, n72142, n72143, n72144, n72145, n72146, n72147, n72148, n72149,
    n72150, n72151, n72152, n72153, n72154, n72155, n72156, n72157, n72158,
    n72159, n72160, n72161, n72162, n72163, n72164, n72165, n72166, n72167,
    n72168, n72169, n72170, n72171, n72172, n72173, n72175, n72176, n72177,
    n72178, n72179, n72180, n72181, n72182, n72183, n72184, n72185, n72186,
    n72187, n72188, n72189, n72190, n72191, n72192, n72193, n72194, n72195,
    n72196, n72197, n72198, n72199, n72200, n72201, n72202, n72203, n72204,
    n72205, n72206, n72207, n72208, n72209, n72210, n72211, n72212, n72213,
    n72214, n72215, n72216, n72217, n72218, n72219, n72220, n72221, n72222,
    n72223, n72224, n72225, n72226, n72227, n72228, n72229, n72230, n72231,
    n72232, n72233, n72234, n72235, n72236, n72237, n72238, n72239, n72240,
    n72241, n72242, n72243, n72244, n72245, n72246, n72247, n72248, n72249,
    n72250, n72251, n72252, n72253, n72254, n72255, n72256, n72257, n72258,
    n72259, n72260, n72261, n72262, n72263, n72264, n72265, n72266, n72267,
    n72268, n72269, n72270, n72271, n72272, n72273, n72274, n72275, n72277,
    n72278, n72279, n72280, n72281, n72282, n72283, n72284, n72285, n72286,
    n72287, n72288, n72289, n72290, n72291, n72292, n72293, n72294, n72295,
    n72296, n72297, n72298, n72299, n72300, n72301, n72302, n72303, n72304,
    n72305, n72306, n72307, n72308, n72309, n72310, n72311, n72312, n72313,
    n72314, n72315, n72317, n72318, n72319, n72320, n72321, n72322, n72323,
    n72324, n72325, n72326, n72327, n72328, n72329, n72330, n72331, n72332,
    n72333, n72334, n72335, n72336, n72337, n72338, n72339, n72340, n72341,
    n72342, n72343, n72344, n72345, n72347, n72348, n72349, n72350, n72351,
    n72352, n72353, n72354, n72355, n72356, n72357, n72358, n72359, n72360,
    n72361, n72362, n72363, n72364, n72365, n72366, n72367, n72368, n72369,
    n72370, n72371, n72372, n72373, n72374, n72375, n72376, n72377, n72378,
    n72379, n72380, n72381, n72382, n72383, n72384, n72385, n72386, n72387,
    n72388, n72389, n72390, n72391, n72392, n72394, n72395, n72396, n72397,
    n72398, n72399, n72400, n72401, n72402, n72403, n72404, n72405, n72406,
    n72407, n72408, n72409, n72410, n72411, n72412, n72413, n72414, n72415,
    n72416, n72417, n72418, n72419, n72420, n72421, n72422, n72423, n72424,
    n72425, n72426, n72427, n72428, n72429, n72430, n72431, n72432, n72433,
    n72434, n72435, n72436, n72437, n72438, n72439, n72440, n72441, n72442,
    n72443, n72444, n72445, n72446, n72447, n72448, n72449, n72450, n72451,
    n72452, n72453, n72454, n72455, n72456, n72457, n72458, n72459, n72460,
    n72461, n72462, n72463, n72464, n72465, n72466, n72467, n72468, n72469,
    n72470, n72471, n72472, n72473, n72474, n72475, n72476, n72477, n72478,
    n72479, n72480, n72481, n72482, n72483, n72484, n72485, n72486, n72487,
    n72488, n72489, n72490, n72491, n72492, n72493, n72494, n72495, n72496,
    n72497, n72498, n72499, n72501, n72502, n72503, n72504, n72505, n72506,
    n72507, n72508, n72509, n72510, n72511, n72512, n72513, n72514, n72515,
    n72516, n72517, n72518, n72519, n72520, n72521, n72522, n72523, n72524,
    n72525, n72526, n72527, n72528, n72529, n72530, n72531, n72532, n72533,
    n72534, n72535, n72536, n72537, n72538, n72540, n72541, n72542, n72543,
    n72544, n72545, n72546, n72547, n72548, n72549, n72550, n72551, n72552,
    n72553, n72554, n72555, n72556, n72557, n72558, n72559, n72560, n72561,
    n72562, n72563, n72564, n72565, n72566, n72567, n72568, n72569, n72570,
    n72571, n72572, n72573, n72574, n72575, n72576, n72577, n72578, n72579,
    n72580, n72581, n72582, n72583, n72584, n72585, n72586, n72587, n72588,
    n72589, n72590, n72591, n72592, n72593, n72594, n72595, n72596, n72597,
    n72598, n72599, n72600, n72601, n72602, n72603, n72604, n72605, n72606,
    n72607, n72608, n72609, n72610, n72611, n72612, n72613, n72614, n72615,
    n72616, n72617, n72618, n72619, n72620, n72621, n72622, n72623, n72624,
    n72625, n72626, n72627, n72628, n72629, n72630, n72631, n72632, n72633,
    n72634, n72635, n72637, n72638, n72639, n72640, n72641, n72642, n72643,
    n72644, n72645, n72646, n72647, n72648, n72649, n72650, n72651, n72652,
    n72653, n72654, n72655, n72656, n72657, n72658, n72659, n72660, n72661,
    n72662, n72663, n72664, n72665, n72666, n72667, n72668, n72669, n72670,
    n72671, n72672, n72674, n72675, n72676, n72677, n72678, n72679, n72680,
    n72681, n72682, n72683, n72684, n72685, n72686, n72687, n72688, n72689,
    n72690, n72691, n72692, n72693, n72694, n72695, n72696, n72697, n72698,
    n72699, n72700, n72701, n72702, n72703, n72704, n72705, n72706, n72707,
    n72708, n72709, n72710, n72711, n72712, n72713, n72715, n72716, n72717,
    n72718, n72719, n72720, n72721, n72722, n72723, n72724, n72725, n72726,
    n72727, n72728, n72729, n72730, n72731, n72732, n72733, n72734, n72735,
    n72736, n72737, n72738, n72739, n72740, n72741, n72742, n72743, n72744,
    n72745, n72746, n72748, n72749, n72750, n72751, n72752, n72753, n72754,
    n72755, n72756, n72757, n72758, n72759, n72760, n72761, n72762, n72763,
    n72764, n72765, n72766, n72767, n72768, n72769, n72770, n72771, n72772,
    n72773, n72774, n72775, n72776, n72778, n72779, n72780, n72781, n72782,
    n72783, n72784, n72785, n72786, n72787, n72788, n72789, n72790, n72791,
    n72792, n72793, n72794, n72795, n72796, n72797, n72798, n72799, n72800,
    n72801, n72802, n72803, n72804, n72805, n72806, n72807, n72808, n72809,
    n72811, n72812, n72813, n72814, n72815, n72816, n72817, n72818, n72819,
    n72820, n72821, n72822, n72823, n72824, n72825, n72826, n72827, n72828,
    n72829, n72830, n72831, n72832, n72833, n72834, n72835, n72836, n72837,
    n72838, n72839, n72840, n72841, n72842, n72843, n72844, n72845, n72846,
    n72847, n72848, n72849, n72850, n72851, n72852, n72853, n72854, n72856,
    n72857, n72858, n72859, n72860, n72861, n72862, n72863, n72864, n72865,
    n72866, n72867, n72868, n72869, n72870, n72871, n72872, n72873, n72874,
    n72875, n72876, n72877, n72878, n72879, n72880, n72881, n72882, n72883,
    n72884, n72885, n72886, n72887, n72889, n72890, n72891, n72892, n72893,
    n72894, n72895, n72896, n72897, n72898, n72899, n72900, n72901, n72902,
    n72903, n72904, n72905, n72906, n72907, n72908, n72909, n72910, n72911,
    n72912, n72913, n72914, n72915, n72916, n72917, n72918, n72919, n72920,
    n72921, n72922, n72923, n72924, n72925, n72927, n72928, n72929, n72930,
    n72931, n72932, n72933, n72934, n72935, n72936, n72937, n72938, n72939,
    n72940, n72941, n72942, n72943, n72944, n72945, n72946, n72947, n72948,
    n72949, n72950, n72951, n72952, n72953, n72954, n72955, n72956, n72957,
    n72958, n72959, n72960, n72961, n72962, n72963, n72964, n72965, n72967,
    n72968, n72969, n72970, n72971, n72972, n72973, n72974, n72975, n72976,
    n72977, n72978, n72979, n72980, n72981, n72982, n72983, n72984, n72985,
    n72986, n72987, n72988, n72989, n72990, n72991, n72992, n72993, n72994,
    n72995, n72996, n72997, n72998, n72999, n73000, n73001, n73002, n73004,
    n73005, n73006, n73007, n73008, n73009, n73010, n73011, n73012, n73013,
    n73014, n73015, n73016, n73017, n73018, n73019, n73020, n73021, n73022,
    n73023, n73024, n73025, n73026, n73027, n73028, n73030, n73031, n73032,
    n73033, n73034, n73035, n73036, n73037, n73038, n73039, n73040, n73041,
    n73042, n73043, n73044, n73045, n73046, n73047, n73048, n73049, n73050,
    n73051, n73052, n73053, n73054, n73055, n73056, n73057, n73058, n73059,
    n73060, n73061, n73062, n73063, n73064, n73065, n73066, n73067, n73068,
    n73069, n73070, n73071, n73072, n73073, n73074, n73075, n73076, n73077,
    n73078, n73079, n73080, n73081, n73082, n73083, n73084, n73085, n73086,
    n73087, n73088, n73089, n73090, n73091, n73092, n73093, n73094, n73095,
    n73096, n73097, n73098, n73099, n73100, n73101, n73102, n73103, n73104,
    n73105, n73106, n73107, n73108, n73109, n73110, n73111, n73112, n73113,
    n73114, n73115, n73116, n73117, n73118, n73119, n73120, n73121, n73122,
    n73123, n73124, n73125, n73126, n73127, n73128, n73129, n73131, n73132,
    n73133, n73134, n73135, n73136, n73137, n73138, n73139, n73140, n73141,
    n73142, n73143, n73144, n73145, n73146, n73147, n73148, n73149, n73150,
    n73151, n73152, n73153, n73154, n73155, n73156, n73157, n73158, n73159,
    n73160, n73161, n73162, n73163, n73164, n73165, n73166, n73167, n73168,
    n73170, n73171, n73172, n73173, n73174, n73175, n73176, n73177, n73178,
    n73179, n73180, n73181, n73182, n73183, n73184, n73185, n73186, n73187,
    n73188, n73189, n73190, n73191, n73192, n73193, n73194, n73195, n73196,
    n73197, n73198, n73199, n73200, n73201, n73202, n73203, n73204, n73205,
    n73206, n73207, n73208, n73209, n73210, n73211, n73212, n73213, n73214,
    n73215, n73216, n73217, n73218, n73219, n73220, n73221, n73222, n73223,
    n73224, n73225, n73226, n73227, n73228, n73229, n73230, n73231, n73232,
    n73233, n73234, n73235, n73236, n73237, n73238, n73239, n73240, n73241,
    n73242, n73243, n73244, n73245, n73246, n73247, n73248, n73249, n73250,
    n73251, n73252, n73253, n73254, n73255, n73256, n73257, n73258, n73259,
    n73260, n73261, n73262, n73263, n73264, n73265, n73266, n73267, n73269,
    n73270, n73271, n73272, n73273, n73274, n73275, n73276, n73277, n73278,
    n73279, n73280, n73281, n73282, n73283, n73284, n73285, n73286, n73287,
    n73288, n73289, n73290, n73291, n73292, n73293, n73294, n73295, n73296,
    n73297, n73298, n73299, n73300, n73301, n73302, n73303, n73304, n73305,
    n73306, n73307, n73308, n73309, n73310, n73311, n73312, n73313, n73314,
    n73315, n73316, n73317, n73318, n73319, n73320, n73321, n73322, n73323,
    n73324, n73325, n73326, n73327, n73328, n73329, n73330, n73331, n73332,
    n73333, n73334, n73335, n73336, n73337, n73338, n73339, n73340, n73341,
    n73342, n73343, n73344, n73345, n73346, n73347, n73348, n73349, n73350,
    n73351, n73352, n73353, n73354, n73355, n73356, n73357, n73358, n73359,
    n73360, n73362, n73363, n73364, n73365, n73366, n73367, n73368, n73369,
    n73370, n73371, n73372, n73373, n73374, n73375, n73376, n73377, n73378,
    n73379, n73380, n73381, n73382, n73383, n73384, n73385, n73386, n73387,
    n73388, n73389, n73390, n73391, n73392, n73393, n73394, n73395, n73397,
    n73398, n73399, n73400, n73401, n73402, n73403, n73404, n73405, n73406,
    n73407, n73408, n73409, n73410, n73411, n73412, n73413, n73414, n73415,
    n73416, n73417, n73418, n73419, n73420, n73421, n73422, n73423, n73424,
    n73425, n73426, n73427, n73428, n73429, n73430, n73431, n73433, n73434,
    n73435, n73436, n73437, n73438, n73439, n73440, n73441, n73442, n73443,
    n73444, n73445, n73446, n73447, n73448, n73449, n73450, n73451, n73452,
    n73453, n73454, n73455, n73456, n73457, n73458, n73459, n73460, n73462,
    n73463, n73464, n73465, n73466, n73467, n73468, n73469, n73470, n73471,
    n73472, n73473, n73474, n73475, n73476, n73477, n73478, n73479, n73480,
    n73481, n73482, n73483, n73484, n73485, n73486, n73487, n73489, n73490,
    n73491, n73492, n73493, n73494, n73495, n73496, n73497, n73498, n73499,
    n73500, n73501, n73502, n73503, n73504, n73505, n73506, n73507, n73508,
    n73509, n73510, n73511, n73512, n73513, n73514, n73515, n73516, n73517,
    n73518, n73519, n73520, n73521, n73522, n73523, n73524, n73525, n73526,
    n73527, n73528, n73529, n73530, n73531, n73532, n73533, n73534, n73535,
    n73536, n73537, n73538, n73539, n73540, n73541, n73542, n73543, n73544,
    n73545, n73546, n73547, n73548, n73549, n73550, n73551, n73552, n73553,
    n73554, n73555, n73556, n73557, n73558, n73559, n73560, n73561, n73562,
    n73563, n73564, n73565, n73566, n73567, n73568, n73569, n73570, n73571,
    n73572, n73573, n73574, n73575, n73576, n73577, n73578, n73579, n73580,
    n73581, n73582, n73583, n73584, n73586, n73587, n73588, n73589, n73590,
    n73591, n73592, n73593, n73594, n73595, n73596, n73597, n73598, n73599,
    n73600, n73601, n73602, n73603, n73604, n73605, n73606, n73607, n73608,
    n73609, n73610, n73611, n73612, n73613, n73614, n73615, n73616, n73617,
    n73618, n73619, n73621, n73622, n73623, n73624, n73625, n73626, n73627,
    n73628, n73629, n73630, n73631, n73632, n73633, n73634, n73635, n73636,
    n73637, n73638, n73639, n73640, n73641, n73642, n73643, n73644, n73645,
    n73646, n73647, n73648, n73649, n73650, n73651, n73652, n73653, n73654,
    n73655, n73656, n73657, n73658, n73659, n73660, n73661, n73662, n73663,
    n73664, n73665, n73666, n73667, n73668, n73669, n73670, n73671, n73672,
    n73673, n73674, n73675, n73676, n73677, n73678, n73679, n73680, n73681,
    n73682, n73683, n73684, n73685, n73686, n73687, n73688, n73689, n73690,
    n73691, n73692, n73693, n73694, n73695, n73696, n73697, n73698, n73699,
    n73700, n73701, n73702, n73703, n73704, n73705, n73706, n73707, n73708,
    n73709, n73710, n73711, n73712, n73713, n73714, n73715, n73717, n73718,
    n73719, n73720, n73721, n73722, n73723, n73724, n73725, n73726, n73727,
    n73728, n73729, n73730, n73731, n73732, n73733, n73734, n73735, n73736,
    n73737, n73738, n73739, n73740, n73741, n73742, n73743, n73744, n73745,
    n73746, n73747, n73748, n73749, n73750, n73751, n73752, n73754, n73755,
    n73756, n73757, n73758, n73759, n73760, n73761, n73762, n73763, n73764,
    n73765, n73766, n73767, n73768, n73769, n73770, n73771, n73772, n73773,
    n73774, n73775, n73776, n73777, n73778, n73779, n73780, n73781, n73782,
    n73783, n73784, n73785, n73786, n73787, n73788, n73789, n73790, n73791,
    n73792, n73793, n73794, n73795, n73796, n73797, n73798, n73799, n73800,
    n73801, n73802, n73803, n73804, n73805, n73806, n73807, n73808, n73809,
    n73810, n73811, n73812, n73813, n73814, n73815, n73816, n73817, n73818,
    n73819, n73820, n73821, n73822, n73823, n73824, n73825, n73826, n73827,
    n73828, n73829, n73830, n73831, n73832, n73833, n73834, n73835, n73836,
    n73837, n73838, n73839, n73840, n73841, n73842, n73843, n73844, n73845,
    n73846, n73847, n73848, n73849, n73850, n73851, n73852, n73853, n73854,
    n73855, n73857, n73858, n73859, n73860, n73861, n73862, n73863, n73864,
    n73865, n73866, n73867, n73868, n73869, n73870, n73871, n73872, n73873,
    n73874, n73875, n73876, n73877, n73878, n73879, n73880, n73881, n73882,
    n73883, n73884, n73885, n73886, n73887, n73888, n73889, n73890, n73891,
    n73892, n73893, n73894, n73895, n73896, n73897, n73898, n73899, n73900,
    n73901, n73902, n73903, n73904, n73905, n73906, n73907, n73908, n73909,
    n73910, n73911, n73912, n73913, n73914, n73915, n73916, n73917, n73918,
    n73919, n73920, n73921, n73922, n73923, n73924, n73925, n73926, n73927,
    n73928, n73929, n73930, n73931, n73932, n73933, n73934, n73935, n73936,
    n73937, n73938, n73939, n73940, n73941, n73942, n73943, n73944, n73945,
    n73946, n73947, n73948, n73949, n73950, n73951, n73952, n73953, n73955,
    n73956, n73957, n73958, n73959, n73960, n73961, n73962, n73963, n73964,
    n73965, n73966, n73967, n73968, n73969, n73970, n73971, n73972, n73973,
    n73974, n73975, n73976, n73977, n73978, n73979, n73980, n73981, n73982,
    n73983, n73984, n73985, n73986, n73988, n73989, n73990, n73991, n73992,
    n73993, n73994, n73995, n73996, n73997, n73998, n73999, n74000, n74001,
    n74002, n74003, n74004, n74005, n74006, n74007, n74008, n74009, n74010,
    n74011, n74012, n74013, n74014, n74015, n74016, n74017, n74018, n74019,
    n74020, n74021, n74022, n74023, n74024, n74025, n74027, n74028, n74029,
    n74030, n74031, n74032, n74033, n74034, n74035, n74036, n74037, n74038,
    n74039, n74040, n74041, n74042, n74043, n74044, n74045, n74046, n74047,
    n74048, n74049, n74050, n74051, n74052, n74053, n74054, n74055, n74056,
    n74057, n74058, n74059, n74060, n74061, n74062, n74063, n74064, n74065,
    n74066, n74067, n74069, n74070, n74071, n74072, n74073, n74074, n74075,
    n74076, n74077, n74078, n74079, n74080, n74081, n74082, n74083, n74084,
    n74085, n74086, n74087, n74088, n74089, n74090, n74091, n74092, n74093,
    n74094, n74095, n74096, n74097, n74098, n74099, n74100, n74101, n74103,
    n74104, n74105, n74106, n74107, n74108, n74109, n74110, n74111, n74112,
    n74113, n74114, n74115, n74116, n74117, n74118, n74119, n74120, n74121,
    n74122, n74123, n74124, n74125, n74126, n74127, n74128, n74129, n74130,
    n74131, n74132, n74133, n74134, n74135, n74137, n74138, n74139, n74140,
    n74141, n74142, n74143, n74144, n74145, n74146, n74147, n74148, n74149,
    n74150, n74151, n74152, n74153, n74154, n74155, n74156, n74157, n74158,
    n74159, n74160, n74161, n74162, n74163, n74164, n74165, n74166, n74167,
    n74168, n74170, n74171, n74172, n74173, n74174, n74175, n74176, n74177,
    n74178, n74179, n74180, n74181, n74182, n74183, n74184, n74185, n74186,
    n74187, n74188, n74189, n74190, n74191, n74192, n74193, n74194, n74195,
    n74196, n74197, n74198, n74199, n74201, n74202, n74203, n74204, n74205,
    n74206, n74207, n74208, n74209, n74210, n74211, n74212, n74213, n74214,
    n74215, n74216, n74217, n74218, n74219, n74220, n74221, n74222, n74223,
    n74224, n74225, n74226, n74227, n74228, n74229, n74230, n74231, n74232,
    n74233, n74234, n74235, n74236, n74237, n74238, n74239, n74240, n74241,
    n74242, n74243, n74244, n74245, n74246, n74247, n74248, n74249, n74250,
    n74251, n74252, n74253, n74254, n74255, n74256, n74257, n74258, n74259,
    n74260, n74261, n74262, n74263, n74264, n74265, n74266, n74267, n74268,
    n74269, n74270, n74271, n74272, n74273, n74274, n74275, n74276, n74277,
    n74278, n74279, n74280, n74281, n74282, n74283, n74284, n74285, n74286,
    n74287, n74288, n74289, n74290, n74291, n74292, n74293, n74295, n74296,
    n74297, n74298, n74299, n74300, n74301, n74302, n74303, n74304, n74305,
    n74306, n74307, n74308, n74309, n74310, n74311, n74312, n74313, n74314,
    n74315, n74316, n74317, n74318, n74319, n74320, n74321, n74323, n74324,
    n74325, n74326, n74327, n74328, n74329, n74330, n74331, n74332, n74333,
    n74334, n74335, n74336, n74337, n74338, n74339, n74340, n74341, n74342,
    n74343, n74344, n74345, n74346, n74347, n74348, n74349, n74350, n74351,
    n74352, n74353, n74354, n74355, n74356, n74357, n74358, n74360, n74361,
    n74362, n74363, n74364, n74365, n74366, n74367, n74368, n74369, n74370,
    n74371, n74372, n74373, n74374, n74375, n74376, n74377, n74378, n74379,
    n74380, n74381, n74382, n74383, n74384, n74385, n74386, n74387, n74389,
    n74390, n74391, n74392, n74393, n74394, n74395, n74396, n74397, n74398,
    n74399, n74400, n74401, n74402, n74403, n74404, n74405, n74406, n74407,
    n74408, n74409, n74410, n74411, n74412, n74413, n74414, n74415, n74416,
    n74417, n74418, n74419, n74420, n74421, n74422, n74423, n74425, n74426,
    n74427, n74428, n74429, n74430, n74431, n74432, n74433, n74434, n74435,
    n74436, n74437, n74438, n74439, n74440, n74441, n74442, n74443, n74444,
    n74445, n74446, n74447, n74448, n74449, n74451, n74452, n74453, n74454,
    n74455, n74456, n74457, n74458, n74459, n74460, n74461, n74462, n74463,
    n74464, n74465, n74466, n74467, n74468, n74469, n74470, n74471, n74472,
    n74473, n74474, n74475, n74476, n74477, n74478, n74479, n74480, n74481,
    n74482, n74483, n74484, n74485, n74486, n74487, n74488, n74489, n74490,
    n74492, n74493, n74494, n74495, n74496, n74497, n74498, n74499, n74500,
    n74501, n74502, n74503, n74504, n74505, n74506, n74507, n74508, n74509,
    n74510, n74511, n74512, n74513, n74514, n74515, n74516, n74517, n74518,
    n74519, n74520, n74521, n74522, n74523, n74524, n74525, n74526, n74528,
    n74529, n74530, n74531, n74532, n74533, n74534, n74535, n74536, n74537,
    n74538, n74539, n74540, n74541, n74542, n74543, n74544, n74545, n74546,
    n74547, n74548, n74549, n74550, n74551, n74552, n74553, n74554, n74555,
    n74556, n74558, n74559, n74560, n74561, n74562, n74563, n74564, n74565,
    n74566, n74567, n74568, n74569, n74570, n74571, n74572, n74573, n74574,
    n74575, n74576, n74577, n74578, n74579, n74580, n74581, n74582, n74583,
    n74584, n74585, n74586, n74587, n74588, n74589, n74590, n74591, n74593,
    n74594, n74595, n74596, n74597, n74598, n74599, n74600, n74601, n74602,
    n74603, n74604, n74605, n74606, n74607, n74608, n74609, n74610, n74611,
    n74612, n74613, n74614, n74615, n74616, n74617, n74618, n74619, n74620,
    n74621, n74622, n74623, n74624, n74626, n74627, n74628, n74629, n74630,
    n74631, n74632, n74633, n74634, n74635, n74636, n74637, n74638, n74639,
    n74640, n74641, n74642, n74643, n74644, n74645, n74646, n74647, n74648,
    n74649, n74650, n74651, n74652, n74653, n74654, n74655, n74656, n74657,
    n74658, n74659, n74660, n74661, n74662, n74663, n74664, n74665, n74666,
    n74667, n74668, n74669, n74670, n74671, n74672, n74673, n74674, n74675,
    n74676, n74677, n74678, n74679, n74680, n74681, n74682, n74683, n74684,
    n74685, n74686, n74687, n74688, n74689, n74690, n74691, n74692, n74693,
    n74694, n74695, n74696, n74697, n74698, n74699, n74700, n74701, n74702,
    n74703, n74704, n74705, n74706, n74707, n74708, n74709, n74710, n74711,
    n74712, n74713, n74714, n74715, n74716, n74717, n74718, n74719, n74720,
    n74721, n74722, n74723, n74724, n74725, n74726, n74727, n74728, n74729,
    n74730, n74732, n74733, n74734, n74735, n74736, n74737, n74738, n74739,
    n74740, n74741, n74742, n74743, n74744, n74745, n74746, n74747, n74748,
    n74749, n74750, n74751, n74752, n74753, n74754, n74755, n74756, n74757,
    n74758, n74759, n74760, n74761, n74762, n74763, n74764, n74765, n74766,
    n74767, n74768, n74769, n74770, n74771, n74773, n74774, n74775, n74776,
    n74777, n74778, n74779, n74780, n74781, n74782, n74783, n74784, n74785,
    n74786, n74787, n74788, n74789, n74790, n74791, n74792, n74793, n74794,
    n74795, n74796, n74797, n74798, n74799, n74800, n74801, n74802, n74803,
    n74804, n74805, n74806, n74807, n74808, n74809, n74811, n74812, n74813,
    n74814, n74815, n74816, n74817, n74818, n74819, n74820, n74821, n74822,
    n74823, n74824, n74825, n74826, n74827, n74828, n74829, n74830, n74831,
    n74832, n74833, n74834, n74835, n74836, n74837, n74838, n74839, n74841,
    n74842, n74843, n74844, n74845, n74846, n74847, n74848, n74849, n74850,
    n74851, n74852, n74853, n74854, n74855, n74856, n74857, n74858, n74859,
    n74860, n74861, n74862, n74863, n74864, n74865, n74866, n74867, n74868,
    n74869, n74870, n74871, n74872, n74873, n74874, n74875, n74876, n74877,
    n74878, n74879, n74880, n74881, n74882, n74883, n74884, n74885, n74886,
    n74887, n74888, n74889, n74890, n74891, n74892, n74893, n74894, n74895,
    n74896, n74897, n74898, n74899, n74900, n74901, n74902, n74903, n74904,
    n74905, n74906, n74907, n74908, n74909, n74910, n74911, n74912, n74913,
    n74914, n74915, n74916, n74917, n74918, n74919, n74920, n74921, n74922,
    n74923, n74924, n74925, n74926, n74927, n74928, n74929, n74931, n74932,
    n74933, n74934, n74935, n74936, n74937, n74938, n74939, n74940, n74941,
    n74942, n74943, n74944, n74945, n74946, n74947, n74948, n74949, n74950,
    n74951, n74952, n74953, n74954, n74955, n74956, n74957, n74958, n74959,
    n74960, n74961, n74962, n74963, n74964, n74965, n74966, n74967, n74968,
    n74969, n74970, n74971, n74972, n74973, n74974, n74975, n74976, n74977,
    n74978, n74979, n74980, n74982, n74983, n74984, n74985, n74986, n74987,
    n74988, n74989, n74990, n74991, n74992, n74993, n74994, n74995, n74996,
    n74997, n74998, n74999, n75000, n75001, n75002, n75003, n75004, n75005,
    n75006, n75007, n75008, n75009, n75010, n75011, n75012, n75013, n75014,
    n75015, n75016, n75017, n75018, n75019, n75020, n75021, n75022, n75023,
    n75024, n75025, n75026, n75027, n75028, n75029, n75030, n75031, n75032,
    n75033, n75034, n75035, n75036, n75037, n75038, n75039, n75040, n75041,
    n75042, n75043, n75044, n75045, n75046, n75047, n75048, n75049, n75050,
    n75051, n75052, n75053, n75054, n75055, n75056, n75057, n75058, n75059,
    n75060, n75061, n75062, n75063, n75064, n75065, n75066, n75067, n75068,
    n75069, n75070, n75071, n75072, n75073, n75074, n75075, n75076, n75077,
    n75078, n75079, n75080, n75081, n75082, n75083, n75085, n75086, n75087,
    n75088, n75089, n75090, n75091, n75092, n75093, n75094, n75095, n75096,
    n75097, n75098, n75099, n75100, n75101, n75102, n75103, n75104, n75105,
    n75106, n75107, n75108, n75109, n75110, n75111, n75112, n75113, n75114,
    n75115, n75116, n75117, n75118, n75119, n75120, n75121, n75122, n75123,
    n75124, n75125, n75126, n75127, n75128, n75129, n75130, n75131, n75132,
    n75133, n75134, n75135, n75136, n75137, n75138, n75139, n75140, n75141,
    n75142, n75143, n75144, n75145, n75146, n75147, n75148, n75149, n75150,
    n75151, n75152, n75153, n75154, n75155, n75156, n75157, n75158, n75159,
    n75160, n75161, n75162, n75163, n75164, n75165, n75166, n75167, n75168,
    n75169, n75170, n75171, n75172, n75173, n75174, n75175, n75176, n75177,
    n75178, n75179, n75180, n75181, n75182, n75183, n75184, n75185, n75187,
    n75188, n75189, n75190, n75191, n75192, n75193, n75194, n75195, n75196,
    n75197, n75198, n75199, n75200, n75201, n75202, n75203, n75204, n75205,
    n75206, n75207, n75208, n75209, n75210, n75211, n75212, n75213, n75214,
    n75215, n75216, n75217, n75218, n75219, n75220, n75221, n75222, n75223,
    n75224, n75225, n75226, n75227, n75228, n75229, n75230, n75231, n75232,
    n75233, n75234, n75235, n75236, n75237, n75238, n75239, n75240, n75241,
    n75242, n75243, n75244, n75245, n75246, n75247, n75248, n75249, n75250,
    n75251, n75252, n75253, n75254, n75255, n75256, n75257, n75258, n75259,
    n75260, n75261, n75262, n75263, n75264, n75265, n75266, n75267, n75268,
    n75269, n75270, n75271, n75272, n75273, n75274, n75275, n75276, n75277,
    n75278, n75279, n75280, n75281, n75282, n75283, n75284, n75285, n75286,
    n75287, n75289, n75290, n75291, n75292, n75293, n75294, n75295, n75296,
    n75297, n75298, n75299, n75300, n75301, n75302, n75303, n75304, n75305,
    n75306, n75307, n75308, n75309, n75310, n75311, n75312, n75313, n75314,
    n75315, n75316, n75317, n75318, n75319, n75320, n75321, n75322, n75323,
    n75324, n75325, n75326, n75327, n75328, n75329, n75330, n75331, n75332,
    n75333, n75334, n75335, n75336, n75337, n75338, n75339, n75340, n75341,
    n75342, n75343, n75344, n75345, n75346, n75347, n75348, n75349, n75350,
    n75351, n75352, n75353, n75354, n75355, n75356, n75357, n75358, n75359,
    n75360, n75361, n75362, n75363, n75364, n75365, n75366, n75367, n75368,
    n75369, n75370, n75371, n75372, n75373, n75374, n75375, n75376, n75377,
    n75378, n75379, n75380, n75381, n75382, n75384, n75385, n75386, n75387,
    n75388, n75389, n75390, n75391, n75392, n75393, n75394, n75395, n75396,
    n75397, n75398, n75399, n75400, n75401, n75402, n75403, n75404, n75405,
    n75406, n75407, n75408, n75409, n75410, n75411, n75412, n75413, n75414,
    n75415, n75416, n75417, n75418, n75419, n75420, n75421, n75423, n75424,
    n75425, n75426, n75427, n75428, n75429, n75430, n75431, n75432, n75433,
    n75434, n75435, n75436, n75437, n75438, n75439, n75440, n75441, n75442,
    n75443, n75444, n75445, n75446, n75447, n75448, n75449, n75450, n75451,
    n75452, n75453, n75454, n75455, n75456, n75457, n75458, n75459, n75460,
    n75461, n75462, n75463, n75464, n75465, n75466, n75467, n75469, n75470,
    n75471, n75472, n75473, n75474, n75475, n75476, n75477, n75478, n75479,
    n75480, n75481, n75482, n75483, n75484, n75485, n75486, n75487, n75488,
    n75489, n75490, n75491, n75492, n75493, n75494, n75495, n75496, n75497,
    n75498, n75499, n75500, n75501, n75502, n75503, n75504, n75505, n75506,
    n75507, n75508, n75509, n75510, n75511, n75512, n75513, n75514, n75516,
    n75517, n75518, n75519, n75520, n75521, n75522, n75523, n75524, n75525,
    n75526, n75527, n75528, n75529, n75530, n75531, n75532, n75533, n75534,
    n75535, n75536, n75537, n75538, n75539, n75540, n75541, n75542, n75543,
    n75544, n75545, n75546, n75547, n75548, n75549, n75550, n75551, n75552,
    n75553, n75554, n75555, n75557, n75558, n75559, n75560, n75561, n75562,
    n75563, n75564, n75565, n75566, n75567, n75568, n75569, n75570, n75571,
    n75572, n75573, n75574, n75575, n75576, n75577, n75578, n75579, n75580,
    n75581, n75582, n75583, n75584, n75585, n75586, n75587, n75588, n75589,
    n75590, n75591, n75592, n75593, n75595, n75596, n75597, n75598, n75599,
    n75600, n75601, n75602, n75603, n75604, n75605, n75606, n75607, n75608,
    n75609, n75610, n75611, n75612, n75613, n75614, n75615, n75616, n75617,
    n75618, n75619, n75620, n75621, n75622, n75623, n75624, n75625, n75626,
    n75627, n75628, n75629, n75630, n75632, n75633, n75634, n75635, n75636,
    n75637, n75638, n75639, n75640, n75641, n75642, n75643, n75644, n75645,
    n75646, n75647, n75648, n75649, n75650, n75651, n75652, n75653, n75654,
    n75655, n75656, n75657, n75658, n75659, n75660, n75661, n75662, n75663,
    n75664, n75665, n75666, n75667, n75668, n75669, n75670, n75671, n75672,
    n75673, n75674, n75675, n75677, n75678, n75679, n75680, n75681, n75682,
    n75683, n75684, n75685, n75686, n75687, n75688, n75689, n75690, n75691,
    n75692, n75693, n75694, n75695, n75696, n75697, n75698, n75699, n75700,
    n75701, n75702, n75703, n75704, n75705, n75706, n75707, n75708, n75709,
    n75711, n75712, n75713, n75714, n75715, n75716, n75717, n75718, n75719,
    n75720, n75721, n75722, n75723, n75724, n75725, n75726, n75727, n75728,
    n75729, n75730, n75731, n75732, n75733, n75734, n75735, n75736, n75737,
    n75738, n75739, n75740, n75741, n75742, n75743, n75744, n75745, n75746,
    n75747, n75749, n75750, n75751, n75752, n75753, n75754, n75755, n75756,
    n75757, n75758, n75759, n75760, n75761, n75762, n75763, n75764, n75765,
    n75766, n75767, n75768, n75769, n75770, n75771, n75772, n75773, n75774,
    n75775, n75776, n75777, n75779, n75780, n75781, n75782, n75783, n75784,
    n75785, n75786, n75787, n75788, n75789, n75790, n75791, n75792, n75793,
    n75794, n75795, n75796, n75797, n75798, n75799, n75800, n75801, n75802,
    n75803, n75804, n75805, n75806, n75807, n75808, n75809, n75810, n75811,
    n75812, n75813, n75814, n75815, n75816, n75817, n75818, n75819, n75820,
    n75821, n75822, n75823, n75824, n75825, n75826, n75827, n75828, n75829,
    n75830, n75831, n75832, n75833, n75834, n75835, n75836, n75837, n75838,
    n75839, n75840, n75841, n75842, n75843, n75844, n75845, n75846, n75847,
    n75848, n75849, n75850, n75851, n75852, n75853, n75854, n75855, n75856,
    n75857, n75858, n75859, n75860, n75861, n75862, n75863, n75864, n75865,
    n75866, n75867, n75868, n75869, n75871, n75872, n75873, n75874, n75875,
    n75876, n75877, n75878, n75879, n75880, n75881, n75882, n75883, n75884,
    n75885, n75886, n75887, n75888, n75889, n75890, n75891, n75892, n75893,
    n75894, n75895, n75897, n75898, n75899, n75900, n75901, n75902, n75903,
    n75904, n75905, n75906, n75907, n75908, n75909, n75910, n75911, n75912,
    n75913, n75914, n75915, n75916, n75917, n75918, n75919, n75920, n75921,
    n75922, n75923, n75924, n75925, n75926, n75927, n75928, n75929, n75930,
    n75931, n75932, n75933, n75934, n75935, n75936, n75937, n75938, n75939,
    n75940, n75941, n75942, n75943, n75945, n75946, n75947, n75948, n75949,
    n75950, n75951, n75952, n75953, n75954, n75955, n75956, n75957, n75958,
    n75959, n75960, n75961, n75962, n75963, n75964, n75965, n75966, n75967,
    n75968, n75969, n75970, n75971, n75972, n75973, n75974, n75975, n75976,
    n75977, n75978, n75980, n75981, n75982, n75983, n75984, n75985, n75986,
    n75987, n75988, n75989, n75990, n75991, n75992, n75993, n75994, n75995,
    n75996, n75997, n75998, n75999, n76000, n76001, n76002, n76003, n76004,
    n76005, n76006, n76007, n76008, n76009, n76010, n76011, n76012, n76013,
    n76014, n76015, n76016, n76017, n76018, n76019, n76020, n76021, n76022,
    n76023, n76024, n76025, n76026, n76027, n76028, n76029, n76030, n76031,
    n76032, n76033, n76034, n76035, n76036, n76037, n76038, n76039, n76040,
    n76041, n76042, n76043, n76044, n76045, n76046, n76047, n76048, n76049,
    n76050, n76051, n76052, n76053, n76054, n76055, n76056, n76057, n76058,
    n76059, n76060, n76061, n76062, n76063, n76064, n76065, n76066, n76067,
    n76069, n76070, n76071, n76072, n76073, n76074, n76075, n76076, n76077,
    n76078, n76079, n76080, n76081, n76082, n76083, n76084, n76085, n76086,
    n76087, n76088, n76089, n76090, n76091, n76092, n76093, n76094, n76095,
    n76096, n76097, n76098, n76099, n76100, n76101, n76102, n76103, n76104,
    n76105, n76106, n76107, n76108, n76109, n76110, n76111, n76113, n76114,
    n76115, n76116, n76117, n76118, n76119, n76120, n76121, n76122, n76123,
    n76124, n76125, n76126, n76127, n76128, n76129, n76130, n76131, n76132,
    n76133, n76134, n76135, n76136, n76137, n76138, n76139, n76140, n76141,
    n76142, n76143, n76144, n76145, n76146, n76147, n76148, n76149, n76150,
    n76151, n76152, n76153, n76154, n76156, n76157, n76158, n76159, n76160,
    n76161, n76162, n76163, n76164, n76165, n76166, n76167, n76168, n76169,
    n76170, n76171, n76172, n76173, n76174, n76175, n76176, n76177, n76178,
    n76179, n76180, n76181, n76182, n76183, n76184, n76185, n76186, n76187,
    n76188, n76189, n76191, n76192, n76193, n76194, n76195, n76196, n76197,
    n76198, n76199, n76200, n76201, n76202, n76203, n76204, n76205, n76206,
    n76207, n76208, n76209, n76210, n76211, n76212, n76213, n76214, n76215,
    n76216, n76217, n76218, n76219, n76220, n76221, n76222, n76223, n76224,
    n76225, n76226, n76227, n76228, n76229, n76230, n76231, n76232, n76233,
    n76234, n76236, n76237, n76238, n76239, n76240, n76241, n76242, n76243,
    n76244, n76245, n76246, n76247, n76248, n76249, n76250, n76251, n76252,
    n76253, n76254, n76255, n76256, n76257, n76258, n76259, n76260, n76261,
    n76262, n76263, n76264, n76265, n76266, n76267, n76269, n76270, n76271,
    n76272, n76273, n76274, n76275, n76276, n76277, n76278, n76279, n76280,
    n76281, n76282, n76283, n76284, n76285, n76286, n76287, n76288, n76289,
    n76290, n76291, n76292, n76293, n76294, n76295, n76296, n76297, n76298,
    n76299, n76300, n76301, n76302, n76303, n76304, n76305, n76306, n76307,
    n76309, n76310, n76311, n76312, n76313, n76314, n76315, n76316, n76317,
    n76318, n76319, n76320, n76321, n76322, n76323, n76324, n76325, n76326,
    n76327, n76328, n76329, n76330, n76331, n76332, n76333, n76334, n76335,
    n76336, n76337, n76338, n76339, n76340, n76341, n76342, n76343, n76345,
    n76346, n76347, n76348, n76349, n76350, n76351, n76352, n76353, n76354,
    n76355, n76356, n76357, n76358, n76359, n76360, n76361, n76362, n76363,
    n76364, n76365, n76366, n76367, n76368, n76369, n76370, n76371, n76372,
    n76373, n76374, n76375, n76376, n76377, n76378, n76379, n76380, n76381,
    n76382, n76383, n76384, n76385, n76386, n76387, n76388, n76389, n76390,
    n76391, n76392, n76393, n76394, n76395, n76396, n76397, n76398, n76399,
    n76400, n76401, n76402, n76403, n76404, n76405, n76406, n76407, n76408,
    n76409, n76410, n76411, n76412, n76413, n76414, n76415, n76416, n76417,
    n76418, n76419, n76420, n76421, n76422, n76423, n76424, n76425, n76426,
    n76427, n76428, n76429, n76430, n76431, n76432, n76433, n76434, n76435,
    n76436, n76437, n76438, n76439, n76440, n76441, n76442, n76443, n76444,
    n76446, n76447, n76448, n76449, n76450, n76451, n76452, n76453, n76454,
    n76455, n76456, n76457, n76458, n76459, n76460, n76461, n76462, n76463,
    n76464, n76465, n76466, n76467, n76468, n76469, n76470, n76471, n76472,
    n76473, n76474, n76475, n76476, n76477, n76478, n76479, n76480, n76481,
    n76482, n76483, n76484, n76485, n76486, n76487, n76488, n76489, n76490,
    n76491, n76492, n76493, n76494, n76495, n76496, n76497, n76498, n76499,
    n76500, n76501, n76502, n76503, n76504, n76505, n76506, n76507, n76508,
    n76509, n76510, n76511, n76512, n76513, n76514, n76515, n76516, n76517,
    n76518, n76519, n76520, n76521, n76522, n76523, n76524, n76525, n76526,
    n76527, n76528, n76529, n76530, n76531, n76532, n76533, n76534, n76535,
    n76536, n76537, n76538, n76539, n76540, n76541, n76542, n76543, n76544,
    n76545, n76546, n76548, n76549, n76550, n76551, n76552, n76553, n76554,
    n76555, n76556, n76557, n76558, n76559, n76560, n76561, n76562, n76563,
    n76564, n76565, n76566, n76567, n76568, n76569, n76570, n76571, n76572,
    n76573, n76574, n76575, n76576, n76577, n76578, n76579, n76580, n76581,
    n76583, n76584, n76585, n76586, n76587, n76588, n76589, n76590, n76591,
    n76592, n76593, n76594, n76595, n76596, n76597, n76598, n76599, n76600,
    n76601, n76602, n76603, n76604, n76605, n76606, n76607, n76608, n76609,
    n76610, n76611, n76612, n76613, n76614, n76615, n76616, n76617, n76618,
    n76619, n76620, n76621, n76622, n76623, n76624, n76625, n76626, n76627,
    n76628, n76629, n76631, n76632, n76633, n76634, n76635, n76636, n76637,
    n76638, n76639, n76640, n76641, n76642, n76643, n76644, n76645, n76646,
    n76647, n76648, n76649, n76650, n76651, n76652, n76653, n76654, n76655,
    n76656, n76657, n76658, n76659, n76660, n76661, n76662, n76663, n76664,
    n76665, n76666, n76667, n76668, n76669, n76670, n76671, n76672, n76673,
    n76674, n76675, n76676, n76677, n76678, n76679, n76680, n76681, n76682,
    n76683, n76684, n76685, n76686, n76687, n76688, n76689, n76690, n76691,
    n76692, n76693, n76694, n76695, n76696, n76697, n76698, n76699, n76700,
    n76701, n76702, n76703, n76704, n76705, n76706, n76707, n76708, n76709,
    n76710, n76711, n76712, n76713, n76714, n76715, n76716, n76717, n76718,
    n76719, n76720, n76721, n76722, n76723, n76724, n76725, n76726, n76727,
    n76728, n76729, n76730, n76731, n76732, n76733, n76734, n76735, n76736,
    n76737, n76738, n76740, n76741, n76742, n76743, n76744, n76745, n76746,
    n76747, n76748, n76749, n76750, n76751, n76752, n76753, n76754, n76755,
    n76756, n76757, n76758, n76759, n76760, n76761, n76762, n76763, n76764,
    n76765, n76766, n76767, n76768, n76769, n76770, n76771, n76772, n76773,
    n76774, n76775, n76776, n76777, n76778, n76779, n76780, n76781, n76782,
    n76783, n76784, n76785, n76786, n76787, n76788, n76789, n76790, n76791,
    n76792, n76793, n76794, n76795, n76796, n76797, n76798, n76799, n76800,
    n76801, n76802, n76803, n76804, n76805, n76806, n76807, n76808, n76809,
    n76810, n76811, n76812, n76813, n76814, n76815, n76816, n76817, n76818,
    n76819, n76820, n76821, n76822, n76823, n76824, n76825, n76826, n76827,
    n76828, n76829, n76830, n76831, n76832, n76833, n76834, n76835, n76836,
    n76837, n76838, n76839, n76840, n76842, n76843, n76844, n76845, n76846,
    n76847, n76848, n76849, n76850, n76851, n76852, n76853, n76854, n76855,
    n76856, n76857, n76858, n76859, n76860, n76861, n76862, n76863, n76864,
    n76865, n76866, n76867, n76868, n76869, n76870, n76871, n76872, n76873,
    n76874, n76876, n76877, n76878, n76879, n76880, n76881, n76882, n76883,
    n76884, n76885, n76886, n76887, n76888, n76889, n76890, n76891, n76892,
    n76893, n76894, n76895, n76896, n76897, n76898, n76899, n76900, n76901,
    n76902, n76903, n76904, n76905, n76906, n76907, n76908, n76909, n76910,
    n76911, n76912, n76913, n76914, n76915, n76916, n76917, n76918, n76919,
    n76920, n76921, n76922, n76923, n76924, n76925, n76926, n76927, n76928,
    n76929, n76930, n76931, n76932, n76933, n76934, n76935, n76936, n76937,
    n76938, n76939, n76940, n76941, n76942, n76943, n76944, n76945, n76946,
    n76947, n76948, n76949, n76950, n76951, n76952, n76953, n76954, n76955,
    n76956, n76957, n76958, n76959, n76960, n76961, n76962, n76963, n76964,
    n76966, n76967, n76968, n76969, n76970, n76971, n76972, n76973, n76974,
    n76975, n76976, n76977, n76978, n76979, n76980, n76981, n76982, n76983,
    n76984, n76985, n76986, n76987, n76988, n76989, n76990, n76991, n76992,
    n76993, n76994, n76995, n76996, n76997, n76998, n77000, n77001, n77002,
    n77003, n77004, n77005, n77006, n77007, n77008, n77009, n77010, n77011,
    n77012, n77013, n77014, n77015, n77016, n77017, n77018, n77019, n77020,
    n77021, n77022, n77023, n77024, n77025, n77026, n77027, n77028, n77029,
    n77030, n77031, n77032, n77033, n77034, n77035, n77036, n77037, n77038,
    n77040, n77041, n77042, n77043, n77044, n77045, n77046, n77047, n77048,
    n77049, n77050, n77051, n77052, n77053, n77054, n77055, n77056, n77057,
    n77058, n77059, n77060, n77061, n77062, n77063, n77064, n77065, n77066,
    n77067, n77068, n77069, n77070, n77071, n77072, n77073, n77074, n77075,
    n77076, n77077, n77078, n77079, n77080, n77081, n77082, n77083, n77084,
    n77085, n77086, n77087, n77089, n77090, n77091, n77092, n77093, n77094,
    n77095, n77096, n77097, n77098, n77099, n77100, n77101, n77102, n77103,
    n77104, n77105, n77106, n77107, n77108, n77109, n77110, n77111, n77112,
    n77113, n77114, n77115, n77116, n77117, n77118, n77119, n77120, n77121,
    n77122, n77124, n77125, n77126, n77127, n77128, n77129, n77130, n77131,
    n77132, n77133, n77134, n77135, n77136, n77137, n77138, n77139, n77140,
    n77141, n77142, n77143, n77144, n77145, n77146, n77147, n77148, n77149,
    n77150, n77151, n77152, n77153, n77154, n77155, n77156, n77157, n77158,
    n77159, n77160, n77161, n77162, n77163, n77164, n77165, n77166, n77167,
    n77168, n77169, n77170, n77171, n77172, n77173, n77174, n77175, n77176,
    n77177, n77178, n77179, n77180, n77181, n77182, n77183, n77184, n77185,
    n77186, n77187, n77188, n77189, n77190, n77191, n77192, n77193, n77194,
    n77195, n77196, n77197, n77198, n77199, n77200, n77201, n77202, n77203,
    n77204, n77205, n77206, n77207, n77208, n77209, n77210, n77211, n77213,
    n77214, n77215, n77216, n77217, n77218, n77219, n77220, n77221, n77222,
    n77223, n77224, n77225, n77226, n77227, n77228, n77229, n77230, n77231,
    n77232, n77233, n77234, n77235, n77236, n77237, n77238, n77239, n77240,
    n77241, n77242, n77243, n77244, n77245, n77246, n77247, n77248, n77249,
    n77250, n77251, n77252, n77253, n77254, n77255, n77257, n77258, n77259,
    n77260, n77261, n77262, n77263, n77264, n77265, n77266, n77267, n77268,
    n77269, n77270, n77271, n77272, n77273, n77274, n77275, n77276, n77277,
    n77278, n77279, n77280, n77281, n77282, n77283, n77284, n77285, n77286,
    n77287, n77288, n77289, n77290, n77291, n77292, n77293, n77294, n77295,
    n77296, n77297, n77298, n77299, n77300, n77301, n77303, n77304, n77305,
    n77306, n77307, n77308, n77309, n77310, n77311, n77312, n77313, n77314,
    n77315, n77316, n77317, n77318, n77319, n77320, n77321, n77322, n77323,
    n77324, n77325, n77326, n77327, n77328, n77329, n77330, n77331, n77332,
    n77333, n77334, n77335, n77336, n77337, n77338, n77339, n77340, n77341,
    n77342, n77343, n77344, n77345, n77346, n77347, n77348, n77349, n77350,
    n77351, n77352, n77353, n77354, n77355, n77356, n77357, n77358, n77359,
    n77360, n77361, n77362, n77363, n77364, n77365, n77366, n77367, n77368,
    n77369, n77370, n77371, n77372, n77373, n77374, n77375, n77376, n77377,
    n77378, n77379, n77380, n77381, n77382, n77383, n77384, n77385, n77386,
    n77387, n77388, n77389, n77390, n77391, n77392, n77393, n77394, n77395,
    n77396, n77397, n77398, n77399, n77400, n77402, n77403, n77404, n77405,
    n77406, n77407, n77408, n77409, n77410, n77411, n77412, n77413, n77414,
    n77415, n77416, n77417, n77418, n77419, n77420, n77421, n77422, n77423,
    n77424, n77425, n77426, n77427, n77428, n77429, n77430, n77431, n77432,
    n77433, n77434, n77435, n77436, n77437, n77438, n77439, n77440, n77441,
    n77442, n77443, n77444, n77445, n77446, n77447, n77448, n77450, n77451,
    n77452, n77453, n77454, n77455, n77456, n77457, n77458, n77459, n77460,
    n77461, n77462, n77463, n77464, n77465, n77466, n77467, n77468, n77469,
    n77470, n77471, n77472, n77473, n77474, n77475, n77476, n77477, n77478,
    n77479, n77480, n77481, n77482, n77483, n77484, n77485, n77486, n77487,
    n77488, n77489, n77490, n77491, n77492, n77493, n77494, n77495, n77496,
    n77497, n77498, n77499, n77501, n77502, n77503, n77504, n77505, n77506,
    n77507, n77508, n77509, n77510, n77511, n77512, n77513, n77514, n77515,
    n77516, n77517, n77518, n77519, n77520, n77521, n77522, n77523, n77524,
    n77525, n77526, n77527, n77528, n77529, n77530, n77531, n77532, n77533,
    n77534, n77535, n77536, n77537, n77538, n77539, n77540, n77542, n77543,
    n77544, n77545, n77546, n77547, n77548, n77549, n77550, n77551, n77552,
    n77553, n77554, n77555, n77556, n77557, n77558, n77559, n77560, n77561,
    n77562, n77563, n77564, n77565, n77566, n77567, n77568, n77569, n77570,
    n77571, n77572, n77573, n77575, n77576, n77577, n77578, n77579, n77580,
    n77581, n77582, n77583, n77584, n77585, n77586, n77587, n77588, n77589,
    n77590, n77591, n77592, n77593, n77594, n77595, n77596, n77597, n77598,
    n77599, n77600, n77601, n77602, n77603, n77604, n77605, n77606, n77607,
    n77608, n77609, n77610, n77611, n77612, n77613, n77614, n77615, n77616,
    n77618, n77619, n77620, n77621, n77622, n77623, n77624, n77625, n77626,
    n77627, n77628, n77629, n77630, n77631, n77632, n77633, n77634, n77635,
    n77636, n77637, n77638, n77639, n77640, n77641, n77642, n77643, n77644,
    n77645, n77646, n77647, n77648, n77649, n77650, n77651, n77652, n77653,
    n77655, n77656, n77657, n77658, n77659, n77660, n77661, n77662, n77663,
    n77664, n77665, n77666, n77667, n77668, n77669, n77670, n77671, n77672,
    n77673, n77674, n77675, n77676, n77677, n77678, n77679, n77680, n77681,
    n77682, n77683, n77684, n77685, n77686, n77687, n77689, n77690, n77691,
    n77692, n77693, n77694, n77695, n77696, n77697, n77698, n77699, n77700,
    n77701, n77702, n77703, n77704, n77705, n77706, n77707, n77708, n77709,
    n77710, n77711, n77712, n77713, n77714, n77715, n77716, n77717, n77718,
    n77719, n77720, n77721, n77722, n77724, n77725, n77726, n77727, n77728,
    n77729, n77730, n77731, n77732, n77733, n77734, n77735, n77736, n77737,
    n77738, n77739, n77740, n77741, n77742, n77743, n77744, n77745, n77746,
    n77747, n77748, n77749, n77750, n77751, n77752, n77753, n77754, n77755,
    n77756, n77757, n77759, n77760, n77761, n77762, n77763, n77764, n77765,
    n77766, n77767, n77768, n77769, n77770, n77771, n77772, n77773, n77774,
    n77775, n77776, n77777, n77778, n77779, n77780, n77781, n77782, n77783,
    n77784, n77785, n77786, n77787, n77788, n77789, n77790, n77791, n77792,
    n77793, n77794, n77795, n77796, n77797, n77798, n77799, n77800, n77801,
    n77802, n77803, n77804, n77805, n77806, n77807, n77808, n77809, n77810,
    n77811, n77812, n77813, n77814, n77815, n77816, n77817, n77818, n77819,
    n77820, n77821, n77822, n77823, n77824, n77825, n77826, n77827, n77828,
    n77829, n77830, n77831, n77832, n77833, n77834, n77835, n77836, n77837,
    n77838, n77839, n77840, n77841, n77842, n77843, n77844, n77845, n77846,
    n77847, n77848, n77849, n77850, n77851, n77852, n77853, n77854, n77855,
    n77857, n77858, n77859, n77860, n77861, n77862, n77863, n77864, n77865,
    n77866, n77867, n77868, n77869, n77870, n77871, n77872, n77873, n77874,
    n77875, n77876, n77877, n77878, n77879, n77880, n77881, n77882, n77883,
    n77884, n77885, n77887, n77888, n77889, n77890, n77891, n77892, n77893,
    n77894, n77895, n77896, n77897, n77898, n77899, n77900, n77901, n77902,
    n77903, n77904, n77905, n77906, n77907, n77908, n77909, n77910, n77911,
    n77913, n77914, n77915, n77916, n77917, n77918, n77919, n77920, n77921,
    n77922, n77923, n77924, n77925, n77926, n77927, n77928, n77929, n77930,
    n77931, n77932, n77933, n77934, n77935, n77936, n77937, n77938, n77939,
    n77940, n77942, n77943, n77944, n77945, n77946, n77947, n77948, n77949,
    n77950, n77951, n77952, n77953, n77954, n77955, n77956, n77957, n77958,
    n77959, n77960, n77961, n77962, n77963, n77964, n77965, n77966, n77967,
    n77968, n77969, n77970, n77971, n77972, n77973, n77974, n77975, n77976,
    n77977, n77978, n77979, n77980, n77981, n77982, n77983, n77984, n77985,
    n77986, n77987, n77988, n77989, n77990, n77991, n77993, n77994, n77995,
    n77996, n77997, n77998, n77999, n78000, n78001, n78002, n78003, n78004,
    n78005, n78006, n78007, n78008, n78009, n78010, n78011, n78012, n78013,
    n78014, n78015, n78016, n78017, n78018, n78019, n78020, n78021, n78022,
    n78023, n78024, n78025, n78026, n78027, n78029, n78030, n78031, n78032,
    n78033, n78034, n78035, n78036, n78037, n78038, n78039, n78040, n78041,
    n78042, n78043, n78044, n78045, n78046, n78047, n78048, n78049, n78050,
    n78051, n78052, n78053, n78054, n78055, n78056, n78057, n78059, n78060,
    n78061, n78062, n78063, n78064, n78065, n78066, n78067, n78068, n78069,
    n78070, n78071, n78072, n78073, n78074, n78075, n78076, n78077, n78078,
    n78079, n78080, n78081, n78082, n78083, n78084, n78085, n78086, n78087,
    n78088, n78089, n78090, n78091, n78092, n78093, n78094, n78095, n78096,
    n78097, n78098, n78099, n78100, n78101, n78102, n78103, n78104, n78105,
    n78106, n78107, n78108, n78109, n78110, n78111, n78112, n78113, n78114,
    n78115, n78116, n78117, n78118, n78119, n78120, n78121, n78122, n78123,
    n78124, n78125, n78126, n78127, n78128, n78129, n78130, n78131, n78132,
    n78133, n78134, n78135, n78136, n78137, n78138, n78139, n78140, n78141,
    n78142, n78143, n78144, n78145, n78146, n78147, n78148, n78149, n78150,
    n78151, n78152, n78153, n78154, n78155, n78156, n78157, n78158, n78159,
    n78160, n78161, n78163, n78164, n78165, n78166, n78167, n78168, n78169,
    n78170, n78171, n78172, n78173, n78174, n78175, n78176, n78177, n78178,
    n78179, n78180, n78181, n78182, n78183, n78184, n78185, n78186, n78187,
    n78188, n78189, n78190, n78191, n78192, n78193, n78194, n78195, n78196,
    n78197, n78198, n78199, n78200, n78201, n78202, n78203, n78204, n78205,
    n78206, n78207, n78209, n78210, n78211, n78212, n78213, n78214, n78215,
    n78216, n78217, n78218, n78219, n78220, n78221, n78222, n78223, n78224,
    n78225, n78226, n78227, n78228, n78229, n78230, n78231, n78232, n78233,
    n78234, n78235, n78236, n78237, n78238, n78239, n78241, n78242, n78243,
    n78244, n78245, n78246, n78247, n78248, n78249, n78250, n78251, n78252,
    n78253, n78254, n78255, n78256, n78257, n78258, n78259, n78260, n78261,
    n78262, n78263, n78264, n78265, n78266, n78267, n78268, n78269, n78270,
    n78271, n78272, n78273, n78274, n78275, n78277, n78278, n78279, n78280,
    n78281, n78282, n78283, n78284, n78285, n78286, n78287, n78288, n78289,
    n78290, n78291, n78292, n78293, n78294, n78295, n78296, n78297, n78298,
    n78299, n78300, n78301, n78302, n78303, n78304, n78305, n78306, n78307,
    n78308, n78309, n78310, n78311, n78312, n78313, n78314, n78315, n78316,
    n78317, n78318, n78319, n78320, n78321, n78322, n78323, n78324, n78325,
    n78326, n78327, n78328, n78329, n78330, n78331, n78332, n78333, n78334,
    n78335, n78336, n78337, n78338, n78339, n78340, n78341, n78342, n78343,
    n78344, n78345, n78346, n78347, n78348, n78349, n78350, n78351, n78352,
    n78353, n78354, n78355, n78356, n78357, n78358, n78359, n78360, n78361,
    n78362, n78363, n78364, n78365, n78366, n78367, n78368, n78369, n78370,
    n78371, n78372, n78373, n78374, n78375, n78376, n78377, n78378, n78380,
    n78381, n78382, n78383, n78384, n78385, n78386, n78387, n78388, n78389,
    n78390, n78391, n78392, n78393, n78394, n78395, n78396, n78397, n78398,
    n78399, n78400, n78401, n78402, n78403, n78404, n78405, n78406, n78407,
    n78408, n78409, n78410, n78411, n78412, n78413, n78414, n78415, n78416,
    n78417, n78418, n78419, n78420, n78421, n78422, n78423, n78424, n78425,
    n78426, n78427, n78428, n78429, n78430, n78431, n78432, n78433, n78434,
    n78435, n78436, n78437, n78438, n78439, n78440, n78441, n78442, n78443,
    n78444, n78445, n78446, n78447, n78448, n78449, n78450, n78451, n78452,
    n78453, n78454, n78455, n78456, n78457, n78458, n78459, n78460, n78461,
    n78462, n78463, n78464, n78465, n78466, n78467, n78468, n78469, n78470,
    n78471, n78472, n78473, n78474, n78475, n78476, n78477, n78478, n78479,
    n78480, n78481, n78483, n78484, n78485, n78486, n78487, n78488, n78489,
    n78490, n78491, n78492, n78493, n78494, n78495, n78496, n78497, n78498,
    n78499, n78500, n78501, n78502, n78503, n78504, n78505, n78506, n78507,
    n78508, n78509, n78510, n78511, n78512, n78513, n78514, n78515, n78516,
    n78517, n78518, n78519, n78520, n78521, n78522, n78523, n78524, n78525,
    n78526, n78527, n78528, n78529, n78530, n78531, n78532, n78533, n78534,
    n78535, n78536, n78537, n78538, n78539, n78540, n78541, n78542, n78543,
    n78544, n78545, n78546, n78547, n78548, n78549, n78550, n78551, n78552,
    n78553, n78554, n78555, n78556, n78557, n78558, n78559, n78560, n78561,
    n78562, n78563, n78564, n78565, n78566, n78567, n78568, n78569, n78570,
    n78571, n78572, n78573, n78574, n78575, n78576, n78577, n78578, n78579,
    n78580, n78581, n78582, n78584, n78585, n78586, n78587, n78588, n78589,
    n78590, n78591, n78592, n78593, n78594, n78595, n78596, n78597, n78598,
    n78599, n78600, n78601, n78602, n78603, n78604, n78605, n78606, n78607,
    n78608, n78609, n78610, n78611, n78612, n78613, n78614, n78615, n78617,
    n78618, n78619, n78620, n78621, n78622, n78623, n78624, n78625, n78626,
    n78627, n78628, n78629, n78630, n78631, n78632, n78633, n78634, n78635,
    n78636, n78637, n78638, n78639, n78640, n78641, n78642, n78643, n78644,
    n78645, n78646, n78647, n78648, n78649, n78650, n78651, n78652, n78653,
    n78654, n78655, n78656, n78657, n78658, n78659, n78660, n78661, n78662,
    n78663, n78664, n78665, n78666, n78667, n78668, n78669, n78670, n78671,
    n78672, n78673, n78674, n78675, n78676, n78677, n78678, n78679, n78680,
    n78681, n78682, n78683, n78684, n78685, n78686, n78687, n78688, n78689,
    n78690, n78691, n78692, n78693, n78694, n78695, n78696, n78697, n78698,
    n78699, n78700, n78701, n78702, n78703, n78704, n78705, n78706, n78707,
    n78708, n78709, n78710, n78712, n78713, n78714, n78715, n78716, n78717,
    n78718, n78719, n78720, n78721, n78722, n78723, n78724, n78725, n78726,
    n78727, n78728, n78729, n78730, n78731, n78732, n78733, n78734, n78735,
    n78736, n78737, n78738, n78739, n78740, n78741, n78742, n78743, n78744,
    n78745, n78746, n78747, n78748, n78749, n78750, n78752, n78753, n78754,
    n78755, n78756, n78757, n78758, n78759, n78760, n78761, n78762, n78763,
    n78764, n78765, n78766, n78767, n78768, n78769, n78770, n78771, n78772,
    n78773, n78774, n78775, n78776, n78777, n78778, n78779, n78780, n78781,
    n78782, n78783, n78784, n78785, n78786, n78787, n78788, n78789, n78790,
    n78791, n78792, n78793, n78794, n78795, n78796, n78797, n78798, n78799,
    n78801, n78802, n78803, n78804, n78805, n78806, n78807, n78808, n78809,
    n78810, n78811, n78812, n78813, n78814, n78815, n78816, n78817, n78818,
    n78819, n78820, n78821, n78822, n78823, n78824, n78825, n78826, n78827,
    n78828, n78829, n78830, n78831, n78832, n78833, n78834, n78835, n78836,
    n78837, n78838, n78839, n78840, n78841, n78842, n78843, n78844, n78845,
    n78847, n78848, n78849, n78850, n78851, n78852, n78853, n78854, n78855,
    n78856, n78857, n78858, n78859, n78860, n78861, n78862, n78863, n78864,
    n78865, n78866, n78867, n78868, n78869, n78870, n78871, n78872, n78873,
    n78874, n78875, n78876, n78877, n78878, n78879, n78880, n78881, n78882,
    n78883, n78884, n78885, n78886, n78887, n78888, n78889, n78890, n78891,
    n78892, n78894, n78895, n78896, n78897, n78898, n78899, n78900, n78901,
    n78902, n78903, n78904, n78905, n78906, n78907, n78908, n78909, n78910,
    n78911, n78912, n78913, n78914, n78915, n78916, n78917, n78918, n78919,
    n78920, n78921, n78922, n78923, n78924, n78925, n78926, n78927, n78928,
    n78929, n78930, n78931, n78932, n78933, n78934, n78935, n78936, n78937,
    n78938, n78939, n78940, n78941, n78943, n78944, n78945, n78946, n78947,
    n78948, n78949, n78950, n78951, n78952, n78953, n78954, n78955, n78956,
    n78957, n78958, n78959, n78960, n78961, n78962, n78963, n78964, n78965,
    n78966, n78967, n78968, n78969, n78970, n78971, n78972, n78973, n78974,
    n78975, n78976, n78977, n78978, n78979, n78980, n78981, n78982, n78983,
    n78984, n78985, n78986, n78987, n78988, n78989, n78990, n78991, n78992,
    n78993, n78994, n78995, n78996, n78997, n78998, n78999, n79000, n79001,
    n79002, n79003, n79004, n79005, n79006, n79007, n79008, n79009, n79010,
    n79011, n79012, n79013, n79014, n79015, n79016, n79017, n79018, n79019,
    n79020, n79021, n79022, n79023, n79024, n79025, n79026, n79027, n79028,
    n79029, n79030, n79031, n79033, n79034, n79035, n79036, n79037, n79038,
    n79039, n79040, n79041, n79042, n79043, n79044, n79045, n79046, n79047,
    n79048, n79049, n79050, n79051, n79052, n79053, n79054, n79055, n79056,
    n79057, n79058, n79059, n79060, n79061, n79062, n79063, n79064, n79065,
    n79066, n79067, n79068, n79069, n79070, n79071, n79072, n79073, n79074,
    n79075, n79076, n79077, n79078, n79079, n79080, n79081, n79082, n79083,
    n79084, n79085, n79086, n79087, n79088, n79089, n79090, n79091, n79092,
    n79093, n79094, n79095, n79096, n79097, n79098, n79099, n79100, n79101,
    n79102, n79103, n79104, n79105, n79106, n79107, n79108, n79109, n79110,
    n79111, n79112, n79113, n79114, n79115, n79116, n79117, n79118, n79119,
    n79120, n79121, n79122, n79123, n79124, n79125, n79126, n79127, n79128,
    n79129, n79131, n79132, n79133, n79134, n79135, n79136, n79137, n79138,
    n79139, n79140, n79141, n79142, n79143, n79144, n79145, n79146, n79147,
    n79148, n79149, n79150, n79151, n79152, n79153, n79154, n79155, n79156,
    n79157, n79158, n79159, n79160, n79161, n79162, n79163, n79164, n79165,
    n79166, n79168, n79169, n79170, n79171, n79172, n79173, n79174, n79175,
    n79176, n79177, n79178, n79179, n79180, n79181, n79182, n79183, n79184,
    n79185, n79186, n79187, n79188, n79189, n79190, n79191, n79192, n79193,
    n79194, n79195, n79196, n79197, n79198, n79199, n79200, n79202, n79203,
    n79204, n79205, n79206, n79207, n79208, n79209, n79210, n79211, n79212,
    n79213, n79214, n79215, n79216, n79217, n79218, n79219, n79220, n79221,
    n79222, n79223, n79224, n79225, n79226, n79227, n79228, n79229, n79230,
    n79231, n79232, n79233, n79234, n79235, n79236, n79237, n79238, n79239,
    n79240, n79241, n79242, n79243, n79244, n79245, n79246, n79247, n79248,
    n79249, n79250, n79251, n79252, n79253, n79254, n79255, n79256, n79257,
    n79258, n79259, n79260, n79261, n79262, n79263, n79264, n79265, n79266,
    n79267, n79268, n79269, n79270, n79271, n79272, n79273, n79274, n79275,
    n79276, n79277, n79278, n79279, n79280, n79281, n79282, n79283, n79284,
    n79285, n79286, n79287, n79288, n79289, n79290, n79291, n79292, n79294,
    n79295, n79296, n79297, n79298, n79299, n79300, n79301, n79302, n79303,
    n79304, n79305, n79306, n79307, n79308, n79309, n79310, n79311, n79312,
    n79313, n79314, n79315, n79316, n79317, n79318, n79319, n79320, n79321,
    n79322, n79324, n79325, n79326, n79327, n79328, n79329, n79330, n79331,
    n79332, n79333, n79334, n79335, n79336, n79337, n79338, n79339, n79340,
    n79341, n79342, n79343, n79344, n79345, n79346, n79347, n79348, n79349,
    n79350, n79351, n79352, n79353, n79354, n79355, n79356, n79357, n79358,
    n79359, n79360, n79361, n79363, n79364, n79365, n79366, n79367, n79368,
    n79369, n79370, n79371, n79372, n79373, n79374, n79375, n79376, n79377,
    n79378, n79379, n79380, n79381, n79382, n79383, n79384, n79385, n79386,
    n79387, n79388, n79389, n79390, n79391, n79392, n79393, n79394, n79395,
    n79396, n79397, n79398, n79399, n79400, n79401, n79402, n79403, n79404,
    n79405, n79406, n79407, n79408, n79409, n79410, n79411, n79412, n79413,
    n79415, n79416, n79417, n79418, n79419, n79420, n79421, n79422, n79423,
    n79424, n79425, n79426, n79427, n79428, n79429, n79430, n79431, n79432,
    n79433, n79434, n79435, n79436, n79437, n79438, n79439, n79440, n79441,
    n79442, n79443, n79444, n79445, n79446, n79447, n79448, n79449, n79451,
    n79452, n79453, n79454, n79455, n79456, n79457, n79458, n79459, n79460,
    n79461, n79462, n79463, n79464, n79465, n79466, n79467, n79468, n79469,
    n79470, n79471, n79472, n79473, n79474, n79475, n79476, n79477, n79478,
    n79479, n79480, n79481, n79482, n79483, n79484, n79485, n79486, n79487,
    n79489, n79490, n79491, n79492, n79493, n79494, n79495, n79496, n79497,
    n79498, n79499, n79500, n79501, n79502, n79503, n79504, n79505, n79506,
    n79507, n79508, n79509, n79510, n79511, n79512, n79513, n79514, n79515,
    n79516, n79517, n79518, n79519, n79520, n79521, n79522, n79523, n79524,
    n79525, n79526, n79527, n79528, n79529, n79530, n79531, n79532, n79533,
    n79534, n79535, n79536, n79537, n79538, n79539, n79540, n79541, n79542,
    n79543, n79545, n79546, n79547, n79548, n79549, n79550, n79551, n79552,
    n79553, n79554, n79555, n79556, n79557, n79558, n79559, n79560, n79561,
    n79562, n79563, n79564, n79565, n79566, n79567, n79568, n79569, n79570,
    n79571, n79572, n79573, n79575, n79576, n79577, n79578, n79579, n79580,
    n79581, n79582, n79583, n79584, n79585, n79586, n79587, n79588, n79589,
    n79590, n79591, n79592, n79593, n79594, n79595, n79596, n79597, n79598,
    n79599, n79600, n79601, n79602, n79603, n79604, n79605, n79606, n79607,
    n79608, n79609, n79610, n79611, n79612, n79613, n79615, n79616, n79617,
    n79618, n79619, n79620, n79621, n79622, n79623, n79624, n79625, n79626,
    n79627, n79628, n79629, n79630, n79631, n79632, n79633, n79634, n79635,
    n79636, n79637, n79638, n79639, n79640, n79641, n79642, n79643, n79644,
    n79645, n79646, n79647, n79648, n79649, n79651, n79652, n79653, n79654,
    n79655, n79656, n79657, n79658, n79659, n79660, n79661, n79662, n79663,
    n79664, n79665, n79666, n79667, n79668, n79669, n79670, n79671, n79672,
    n79673, n79674, n79675, n79676, n79677, n79678, n79679, n79680, n79681,
    n79682, n79684, n79685, n79686, n79687, n79688, n79689, n79690, n79691,
    n79692, n79693, n79694, n79695, n79696, n79697, n79698, n79699, n79700,
    n79701, n79702, n79703, n79704, n79705, n79706, n79707, n79708, n79709,
    n79710, n79711, n79712, n79713, n79714, n79715, n79716, n79717, n79718,
    n79719, n79720, n79722, n79723, n79724, n79725, n79726, n79727, n79728,
    n79729, n79730, n79731, n79732, n79733, n79734, n79735, n79736, n79737,
    n79738, n79739, n79740, n79741, n79742, n79743, n79744, n79745, n79746,
    n79747, n79748, n79749, n79750, n79751, n79752, n79753, n79754, n79755,
    n79756, n79757, n79758, n79759, n79761, n79762, n79763, n79764, n79765,
    n79766, n79767, n79768, n79769, n79770, n79771, n79772, n79773, n79774,
    n79775, n79776, n79777, n79778, n79779, n79780, n79781, n79782, n79783,
    n79784, n79785, n79787, n79788, n79789, n79790, n79791, n79792, n79793,
    n79794, n79795, n79796, n79797, n79798, n79799, n79800, n79801, n79802,
    n79803, n79804, n79805, n79806, n79807, n79808, n79809, n79810, n79811,
    n79812, n79813, n79814, n79815, n79816, n79817, n79818, n79819, n79820,
    n79821, n79822, n79823, n79824, n79825, n79826, n79827, n79828, n79829,
    n79830, n79831, n79832, n79833, n79834, n79835, n79836, n79837, n79838,
    n79839, n79840, n79841, n79842, n79843, n79844, n79845, n79846, n79847,
    n79848, n79849, n79850, n79851, n79852, n79853, n79854, n79855, n79856,
    n79857, n79858, n79859, n79860, n79861, n79862, n79863, n79864, n79865,
    n79866, n79867, n79868, n79869, n79870, n79871, n79872, n79873, n79874,
    n79875, n79876, n79877, n79878, n79879, n79880, n79881, n79882, n79883,
    n79884, n79885, n79886, n79888, n79889, n79890, n79891, n79892, n79893,
    n79894, n79895, n79896, n79897, n79898, n79899, n79900, n79901, n79902,
    n79903, n79904, n79905, n79906, n79907, n79908, n79909, n79910, n79911,
    n79912, n79913, n79914, n79915, n79916, n79917, n79918, n79919, n79920,
    n79921, n79922, n79923, n79924, n79925, n79926, n79927, n79929, n79930,
    n79931, n79932, n79933, n79934, n79935, n79936, n79937, n79938, n79939,
    n79940, n79941, n79942, n79943, n79944, n79945, n79946, n79947, n79948,
    n79949, n79950, n79951, n79952, n79953, n79954, n79955, n79956, n79957,
    n79958, n79959, n79960, n79961, n79962, n79963, n79964, n79965, n79966,
    n79967, n79968, n79969, n79970, n79971, n79972, n79973, n79974, n79975,
    n79976, n79977, n79978, n79979, n79980, n79981, n79982, n79983, n79984,
    n79985, n79986, n79987, n79988, n79989, n79990, n79991, n79992, n79993,
    n79994, n79995, n79996, n79997, n79998, n79999, n80000, n80001, n80002,
    n80003, n80004, n80005, n80006, n80007, n80008, n80009, n80010, n80011,
    n80012, n80013, n80014, n80015, n80016, n80017, n80018, n80019, n80020,
    n80021, n80022, n80023, n80024, n80025, n80026, n80027, n80028, n80029,
    n80030, n80031, n80032, n80033, n80034, n80036, n80037, n80038, n80039,
    n80040, n80041, n80042, n80043, n80044, n80045, n80046, n80047, n80048,
    n80049, n80050, n80051, n80052, n80053, n80054, n80055, n80056, n80057,
    n80058, n80059, n80060, n80061, n80062, n80063, n80064, n80065, n80066,
    n80067, n80068, n80069, n80070, n80071, n80072, n80073, n80074, n80076,
    n80077, n80078, n80079, n80080, n80081, n80082, n80083, n80084, n80085,
    n80086, n80087, n80088, n80089, n80090, n80091, n80092, n80093, n80094,
    n80095, n80096, n80097, n80098, n80099, n80100, n80101, n80102, n80103,
    n80104, n80105, n80106, n80107, n80108, n80109, n80110, n80111, n80112,
    n80113, n80114, n80115, n80117, n80118, n80119, n80120, n80121, n80122,
    n80123, n80124, n80125, n80126, n80127, n80128, n80129, n80130, n80131,
    n80132, n80133, n80134, n80135, n80136, n80137, n80138, n80139, n80140,
    n80141, n80142, n80143, n80144, n80145, n80146, n80147, n80148, n80149,
    n80150, n80151, n80152, n80153, n80154, n80155, n80156, n80157, n80158,
    n80159, n80160, n80161, n80162, n80163, n80164, n80165, n80166, n80167,
    n80168, n80169, n80170, n80171, n80172, n80173, n80174, n80175, n80176,
    n80177, n80178, n80179, n80180, n80181, n80182, n80183, n80184, n80185,
    n80186, n80187, n80188, n80189, n80190, n80191, n80192, n80193, n80194,
    n80195, n80196, n80197, n80198, n80199, n80200, n80201, n80202, n80203,
    n80204, n80205, n80206, n80207, n80208, n80209, n80210, n80211, n80213,
    n80214, n80215, n80216, n80217, n80218, n80219, n80220, n80221, n80222,
    n80223, n80224, n80225, n80226, n80227, n80228, n80229, n80230, n80231,
    n80232, n80233, n80234, n80235, n80236, n80237, n80238, n80239, n80240,
    n80241, n80242, n80243, n80244, n80245, n80246, n80247, n80248, n80249,
    n80250, n80251, n80252, n80253, n80254, n80255, n80257, n80258, n80259,
    n80260, n80261, n80262, n80263, n80264, n80265, n80266, n80267, n80268,
    n80269, n80270, n80271, n80272, n80273, n80274, n80275, n80276, n80277,
    n80278, n80279, n80280, n80281, n80282, n80283, n80284, n80285, n80286,
    n80287, n80288, n80289, n80290, n80291, n80292, n80293, n80294, n80295,
    n80296, n80297, n80298, n80299, n80300, n80301, n80302, n80303, n80304,
    n80305, n80306, n80307, n80308, n80309, n80310, n80311, n80312, n80313,
    n80314, n80315, n80316, n80317, n80318, n80319, n80320, n80321, n80322,
    n80323, n80324, n80325, n80326, n80327, n80328, n80329, n80330, n80331,
    n80332, n80333, n80334, n80335, n80336, n80337, n80338, n80339, n80340,
    n80341, n80342, n80343, n80344, n80345, n80346, n80347, n80348, n80349,
    n80350, n80351, n80352, n80353, n80354, n80355, n80356, n80357, n80358,
    n80359, n80360, n80361, n80363, n80364, n80365, n80366, n80367, n80368,
    n80369, n80370, n80371, n80372, n80373, n80374, n80375, n80376, n80377,
    n80378, n80379, n80380, n80381, n80382, n80383, n80384, n80385, n80386,
    n80387, n80388, n80389, n80390, n80391, n80392, n80393, n80394, n80395,
    n80396, n80397, n80398, n80399, n80400, n80401, n80402, n80403, n80404,
    n80405, n80406, n80407, n80408, n80409, n80410, n80411, n80412, n80413,
    n80414, n80415, n80416, n80417, n80418, n80419, n80420, n80421, n80422,
    n80423, n80424, n80425, n80426, n80427, n80428, n80429, n80430, n80431,
    n80432, n80433, n80434, n80435, n80436, n80437, n80438, n80439, n80440,
    n80441, n80442, n80443, n80444, n80445, n80446, n80447, n80448, n80449,
    n80450, n80451, n80452, n80453, n80454, n80455, n80456, n80457, n80458,
    n80459, n80460, n80461, n80462, n80463, n80464, n80465, n80466, n80468,
    n80469, n80470, n80471, n80472, n80473, n80474, n80475, n80476, n80477,
    n80478, n80479, n80480, n80481, n80482, n80483, n80484, n80485, n80486,
    n80487, n80488, n80489, n80490, n80491, n80492, n80493, n80494, n80495,
    n80496, n80497, n80498, n80499, n80500, n80501, n80502, n80504, n80505,
    n80506, n80507, n80508, n80509, n80510, n80511, n80512, n80513, n80514,
    n80515, n80516, n80517, n80518, n80519, n80520, n80521, n80522, n80523,
    n80524, n80525, n80526, n80527, n80528, n80529, n80530, n80531, n80532,
    n80533, n80534, n80535, n80536, n80537, n80538, n80539, n80540, n80541,
    n80543, n80544, n80545, n80546, n80547, n80548, n80549, n80550, n80551,
    n80552, n80553, n80554, n80555, n80556, n80557, n80558, n80559, n80560,
    n80561, n80562, n80563, n80564, n80565, n80566, n80567, n80568, n80569,
    n80570, n80571, n80573, n80574, n80575, n80576, n80577, n80578, n80579,
    n80580, n80581, n80582, n80583, n80584, n80585, n80586, n80587, n80588,
    n80589, n80590, n80591, n80592, n80593, n80594, n80595, n80596, n80597,
    n80598, n80599, n80600, n80601, n80602, n80603, n80604, n80605, n80606,
    n80607, n80608, n80609, n80610, n80611, n80612, n80613, n80614, n80615,
    n80616, n80617, n80618, n80619, n80620, n80621, n80622, n80623, n80624,
    n80625, n80626, n80627, n80628, n80629, n80630, n80631, n80632, n80633,
    n80634, n80635, n80636, n80637, n80638, n80639, n80640, n80641, n80642,
    n80643, n80644, n80645, n80646, n80647, n80648, n80649, n80650, n80651,
    n80652, n80653, n80654, n80655, n80656, n80657, n80658, n80659, n80660,
    n80661, n80662, n80663, n80664, n80665, n80666, n80667, n80668, n80669,
    n80670, n80672, n80673, n80674, n80675, n80676, n80677, n80678, n80679,
    n80680, n80681, n80682, n80683, n80684, n80685, n80686, n80687, n80688,
    n80689, n80690, n80691, n80692, n80693, n80694, n80695, n80696, n80697,
    n80698, n80699, n80700, n80701, n80702, n80703, n80704, n80705, n80706,
    n80707, n80708, n80709, n80710, n80711, n80712, n80713, n80714, n80715,
    n80717, n80718, n80719, n80720, n80721, n80722, n80723, n80724, n80725,
    n80726, n80727, n80728, n80729, n80730, n80731, n80732, n80733, n80734,
    n80735, n80736, n80737, n80738, n80739, n80740, n80741, n80742, n80743,
    n80744, n80745, n80746, n80747, n80748, n80749, n80750, n80751, n80752,
    n80753, n80754, n80755, n80756, n80757, n80759, n80760, n80761, n80762,
    n80763, n80764, n80765, n80766, n80767, n80768, n80769, n80770, n80771,
    n80772, n80773, n80774, n80775, n80776, n80777, n80778, n80779, n80780,
    n80781, n80782, n80783, n80784, n80785, n80786, n80787, n80788, n80789,
    n80790, n80791, n80792, n80793, n80794, n80795, n80797, n80798, n80799,
    n80800, n80801, n80802, n80803, n80804, n80805, n80806, n80807, n80808,
    n80809, n80810, n80811, n80812, n80813, n80814, n80815, n80816, n80817,
    n80818, n80819, n80820, n80821, n80822, n80823, n80824, n80825, n80827,
    n80828, n80829, n80830, n80831, n80832, n80833, n80834, n80835, n80836,
    n80837, n80838, n80839, n80840, n80841, n80842, n80843, n80844, n80845,
    n80846, n80847, n80848, n80849, n80850, n80851, n80852, n80853, n80854,
    n80855, n80857, n80858, n80859, n80860, n80861, n80862, n80863, n80864,
    n80865, n80866, n80867, n80868, n80869, n80870, n80871, n80872, n80873,
    n80874, n80875, n80876, n80877, n80878, n80879, n80880, n80881, n80882,
    n80883, n80884, n80885, n80886, n80887, n80888, n80889, n80890, n80891,
    n80893, n80894, n80895, n80896, n80897, n80898, n80899, n80900, n80901,
    n80902, n80903, n80904, n80905, n80906, n80907, n80908, n80909, n80910,
    n80911, n80912, n80913, n80914, n80915, n80916, n80917, n80918, n80919,
    n80920, n80921, n80922, n80923, n80924, n80925, n80926, n80927, n80928,
    n80929, n80930, n80932, n80933, n80934, n80935, n80936, n80937, n80938,
    n80939, n80940, n80941, n80942, n80943, n80944, n80945, n80946, n80947,
    n80948, n80949, n80950, n80951, n80952, n80953, n80954, n80955, n80956,
    n80957, n80959, n80960, n80961, n80962, n80963, n80964, n80965, n80966,
    n80967, n80968, n80969, n80970, n80971, n80972, n80973, n80974, n80975,
    n80976, n80977, n80978, n80979, n80980, n80981, n80982, n80983, n80984,
    n80985, n80986, n80987, n80988, n80989, n80990, n80991, n80992, n80993,
    n80994, n80995, n80996, n80997, n80998, n80999, n81000, n81001, n81002,
    n81003, n81004, n81005, n81006, n81007, n81008, n81009, n81010, n81011,
    n81012, n81013, n81014, n81015, n81016, n81017, n81018, n81019, n81020,
    n81021, n81022, n81023, n81024, n81025, n81026, n81027, n81028, n81029,
    n81030, n81031, n81032, n81033, n81034, n81035, n81036, n81037, n81038,
    n81039, n81040, n81041, n81042, n81043, n81044, n81045, n81046, n81047,
    n81048, n81049, n81050, n81051, n81052, n81053, n81054, n81055, n81056,
    n81057, n81058, n81059, n81061, n81062, n81063, n81064, n81065, n81066,
    n81067, n81068, n81069, n81070, n81071, n81072, n81073, n81074, n81075,
    n81076, n81077, n81078, n81079, n81080, n81081, n81082, n81083, n81084,
    n81085, n81086, n81087, n81088, n81089, n81090, n81091, n81092, n81094,
    n81095, n81096, n81097, n81098, n81099, n81100, n81101, n81102, n81103,
    n81104, n81105, n81106, n81107, n81108, n81109, n81110, n81111, n81112,
    n81113, n81114, n81115, n81116, n81117, n81118, n81119, n81120, n81121,
    n81122, n81123, n81124, n81125, n81126, n81127, n81128, n81129, n81130,
    n81131, n81132, n81134, n81135, n81136, n81137, n81138, n81139, n81140,
    n81141, n81142, n81143, n81144, n81145, n81146, n81147, n81148, n81149,
    n81150, n81151, n81152, n81153, n81154, n81155, n81156, n81157, n81158,
    n81159, n81160, n81161, n81162, n81163, n81164, n81165, n81166, n81167,
    n81168, n81169, n81170, n81171, n81172, n81173, n81175, n81176, n81177,
    n81178, n81179, n81180, n81181, n81182, n81183, n81184, n81185, n81186,
    n81187, n81188, n81189, n81190, n81191, n81192, n81193, n81194, n81195,
    n81196, n81197, n81198, n81199, n81200, n81201, n81202, n81203, n81204,
    n81205, n81206, n81207, n81208, n81209, n81210, n81211, n81212, n81213,
    n81214, n81215, n81216, n81217, n81219, n81220, n81221, n81222, n81223,
    n81224, n81225, n81226, n81227, n81228, n81229, n81230, n81231, n81232,
    n81233, n81234, n81235, n81236, n81237, n81238, n81239, n81240, n81241,
    n81242, n81243, n81244, n81245, n81246, n81247, n81248, n81249, n81250,
    n81251, n81252, n81253, n81254, n81255, n81256, n81257, n81258, n81259,
    n81260, n81261, n81262, n81263, n81264, n81265, n81266, n81267, n81268,
    n81269, n81270, n81271, n81272, n81273, n81274, n81275, n81276, n81277,
    n81278, n81279, n81280, n81281, n81282, n81283, n81284, n81285, n81286,
    n81287, n81288, n81289, n81290, n81291, n81292, n81293, n81294, n81295,
    n81296, n81297, n81298, n81299, n81300, n81301, n81302, n81303, n81304,
    n81305, n81306, n81307, n81308, n81309, n81310, n81311, n81312, n81314,
    n81315, n81316, n81317, n81318, n81319, n81320, n81321, n81322, n81323,
    n81324, n81325, n81326, n81327, n81328, n81329, n81330, n81331, n81332,
    n81333, n81334, n81335, n81336, n81337, n81338, n81339, n81340, n81341,
    n81342, n81343, n81344, n81345, n81346, n81347, n81348, n81349, n81351,
    n81352, n81353, n81354, n81355, n81356, n81357, n81358, n81359, n81360,
    n81361, n81362, n81363, n81364, n81365, n81366, n81367, n81368, n81369,
    n81370, n81371, n81372, n81373, n81374, n81375, n81376, n81377, n81378,
    n81379, n81380, n81381, n81382, n81383, n81384, n81385, n81386, n81387,
    n81388, n81389, n81390, n81391, n81392, n81394, n81395, n81396, n81397,
    n81398, n81399, n81400, n81401, n81402, n81403, n81404, n81405, n81406,
    n81407, n81408, n81409, n81410, n81411, n81412, n81413, n81414, n81415,
    n81416, n81417, n81418, n81419, n81420, n81421, n81422, n81423, n81424,
    n81425, n81426, n81427, n81428, n81429, n81430, n81431, n81433, n81434,
    n81435, n81436, n81437, n81438, n81439, n81440, n81441, n81442, n81443,
    n81444, n81445, n81446, n81447, n81448, n81449, n81450, n81451, n81452,
    n81453, n81454, n81455, n81456, n81457, n81458, n81459, n81460, n81461,
    n81462, n81463, n81464, n81465, n81466, n81467, n81469, n81470, n81471,
    n81472, n81473, n81474, n81475, n81476, n81477, n81478, n81479, n81480,
    n81481, n81482, n81483, n81484, n81485, n81486, n81487, n81488, n81489,
    n81490, n81491, n81492, n81493, n81494, n81495, n81496, n81497, n81498,
    n81499, n81500, n81502, n81503, n81504, n81505, n81506, n81507, n81508,
    n81509, n81510, n81511, n81512, n81513, n81514, n81515, n81516, n81517,
    n81518, n81519, n81520, n81521, n81522, n81523, n81524, n81525, n81526,
    n81527, n81528, n81529, n81530, n81531, n81532, n81533, n81534, n81535,
    n81536, n81537, n81538, n81539, n81540, n81541, n81542, n81543, n81544,
    n81545, n81546, n81547, n81548, n81549, n81550, n81551, n81552, n81553,
    n81554, n81555, n81556, n81557, n81558, n81559, n81560, n81561, n81562,
    n81563, n81564, n81565, n81566, n81567, n81568, n81569, n81570, n81571,
    n81572, n81573, n81574, n81575, n81576, n81577, n81578, n81579, n81580,
    n81581, n81582, n81583, n81584, n81585, n81586, n81587, n81588, n81589,
    n81590, n81591, n81592, n81593, n81594, n81595, n81596, n81597, n81598,
    n81599, n81600, n81601, n81602, n81604, n81605, n81606, n81607, n81608,
    n81609, n81610, n81611, n81612, n81613, n81614, n81615, n81616, n81617,
    n81618, n81619, n81620, n81621, n81622, n81623, n81624, n81625, n81626,
    n81627, n81628, n81629, n81630, n81631, n81632, n81633, n81634, n81635,
    n81636, n81637, n81638, n81639, n81640, n81641, n81642, n81643, n81644,
    n81645, n81646, n81647, n81648, n81649, n81650, n81651, n81652, n81653,
    n81654, n81655, n81656, n81657, n81658, n81659, n81660, n81661, n81662,
    n81663, n81664, n81665, n81666, n81667, n81668, n81669, n81670, n81671,
    n81672, n81673, n81674, n81675, n81676, n81677, n81678, n81679, n81680,
    n81681, n81682, n81683, n81684, n81685, n81686, n81687, n81688, n81689,
    n81690, n81691, n81692, n81693, n81694, n81695, n81696, n81697, n81698,
    n81699, n81700, n81701, n81702, n81703, n81704, n81706, n81707, n81708,
    n81709, n81710, n81711, n81712, n81713, n81714, n81715, n81716, n81717,
    n81718, n81719, n81720, n81721, n81722, n81723, n81724, n81725, n81726,
    n81727, n81728, n81729, n81730, n81731, n81732, n81733, n81734, n81735,
    n81736, n81737, n81738, n81739, n81740, n81741, n81742, n81743, n81744,
    n81745, n81746, n81747, n81749, n81750, n81751, n81752, n81753, n81754,
    n81755, n81756, n81757, n81758, n81759, n81760, n81761, n81762, n81763,
    n81764, n81765, n81766, n81767, n81768, n81769, n81770, n81771, n81772,
    n81773, n81774, n81775, n81776, n81777, n81779, n81780, n81781, n81782,
    n81783, n81784, n81785, n81786, n81787, n81788, n81789, n81790, n81791,
    n81792, n81793, n81794, n81795, n81796, n81797, n81798, n81799, n81800,
    n81801, n81802, n81803, n81804, n81805, n81806, n81807, n81808, n81809,
    n81810, n81811, n81812, n81813, n81814, n81815, n81816, n81817, n81818,
    n81819, n81820, n81821, n81822, n81823, n81824, n81826, n81827, n81828,
    n81829, n81830, n81831, n81832, n81833, n81834, n81835, n81836, n81837,
    n81838, n81839, n81840, n81841, n81842, n81843, n81844, n81845, n81846,
    n81847, n81848, n81849, n81850, n81851, n81852, n81853, n81854, n81855,
    n81856, n81857, n81858, n81859, n81860, n81861, n81862, n81864, n81865,
    n81866, n81867, n81868, n81869, n81870, n81871, n81872, n81873, n81874,
    n81875, n81876, n81877, n81878, n81879, n81880, n81881, n81882, n81883,
    n81884, n81885, n81886, n81887, n81888, n81889, n81890, n81891, n81892,
    n81893, n81894, n81895, n81896, n81897, n81898, n81900, n81901, n81902,
    n81903, n81904, n81905, n81906, n81907, n81908, n81909, n81910, n81911,
    n81912, n81913, n81914, n81915, n81916, n81917, n81918, n81919, n81920,
    n81921, n81922, n81923, n81924, n81925, n81926, n81927, n81928, n81929,
    n81930, n81931, n81932, n81933, n81934, n81935, n81936, n81937, n81938,
    n81939, n81940, n81941, n81942, n81943, n81944, n81945, n81946, n81947,
    n81948, n81949, n81950, n81951, n81952, n81953, n81954, n81955, n81956,
    n81957, n81958, n81959, n81960, n81961, n81962, n81963, n81964, n81965,
    n81966, n81967, n81968, n81969, n81970, n81971, n81972, n81973, n81974,
    n81975, n81976, n81977, n81978, n81979, n81980, n81981, n81982, n81983,
    n81984, n81985, n81986, n81987, n81988, n81989, n81990, n81991, n81992,
    n81993, n81994, n81995, n81996, n81997, n81998, n81999, n82000, n82001,
    n82002, n82003, n82005, n82006, n82007, n82008, n82009, n82010, n82011,
    n82012, n82013, n82014, n82015, n82016, n82017, n82018, n82019, n82020,
    n82021, n82022, n82023, n82024, n82025, n82026, n82027, n82028, n82029,
    n82030, n82031, n82032, n82033, n82034, n82035, n82036, n82037, n82038,
    n82039, n82040, n82041, n82042, n82043, n82044, n82045, n82046, n82047,
    n82048, n82049, n82050, n82051, n82052, n82053, n82054, n82055, n82056,
    n82057, n82058, n82059, n82060, n82061, n82062, n82063, n82064, n82065,
    n82066, n82067, n82068, n82069, n82070, n82071, n82072, n82073, n82074,
    n82075, n82076, n82077, n82078, n82079, n82080, n82081, n82082, n82083,
    n82084, n82085, n82086, n82087, n82088, n82089, n82090, n82091, n82092,
    n82093, n82094, n82096, n82097, n82098, n82099, n82100, n82101, n82102,
    n82103, n82104, n82105, n82106, n82107, n82108, n82109, n82110, n82111,
    n82112, n82113, n82114, n82115, n82116, n82117, n82118, n82119, n82120,
    n82121, n82122, n82123, n82124, n82125, n82126, n82127, n82128, n82129,
    n82130, n82131, n82132, n82133, n82134, n82135, n82136, n82137, n82138,
    n82139, n82140, n82141, n82142, n82143, n82144, n82145, n82146, n82147,
    n82148, n82149, n82150, n82151, n82152, n82153, n82154, n82155, n82156,
    n82157, n82158, n82159, n82160, n82161, n82162, n82163, n82164, n82165,
    n82166, n82167, n82168, n82169, n82170, n82171, n82172, n82173, n82174,
    n82175, n82176, n82177, n82178, n82179, n82180, n82181, n82182, n82183,
    n82184, n82185, n82186, n82187, n82188, n82189, n82190, n82191, n82192,
    n82193, n82194, n82195, n82196, n82197, n82198, n82200, n82201, n82202,
    n82203, n82204, n82205, n82206, n82207, n82208, n82209, n82210, n82211,
    n82212, n82213, n82214, n82215, n82216, n82217, n82218, n82219, n82220,
    n82221, n82222, n82223, n82224, n82225, n82226, n82227, n82228, n82229,
    n82230, n82231, n82232, n82233, n82234, n82235, n82236, n82237, n82238,
    n82239, n82240, n82241, n82242, n82243, n82244, n82245, n82246, n82247,
    n82249, n82250, n82251, n82252, n82253, n82254, n82255, n82256, n82257,
    n82258, n82259, n82260, n82261, n82262, n82263, n82264, n82265, n82266,
    n82267, n82268, n82269, n82270, n82271, n82272, n82273, n82274, n82275,
    n82276, n82277, n82278, n82279, n82280, n82281, n82282, n82283, n82284,
    n82285, n82286, n82287, n82288, n82289, n82290, n82291, n82292, n82293,
    n82294, n82295, n82296, n82298, n82299, n82300, n82301, n82302, n82303,
    n82304, n82305, n82306, n82307, n82308, n82309, n82310, n82311, n82312,
    n82313, n82314, n82315, n82316, n82317, n82318, n82319, n82320, n82321,
    n82322, n82323, n82324, n82325, n82326, n82327, n82328, n82329, n82330,
    n82332, n82333, n82334, n82335, n82336, n82337, n82338, n82339, n82340,
    n82341, n82342, n82343, n82344, n82345, n82346, n82347, n82348, n82349,
    n82350, n82351, n82352, n82353, n82354, n82355, n82356, n82357, n82358,
    n82359, n82360, n82361, n82362, n82363, n82364, n82365, n82366, n82367,
    n82368, n82369, n82370, n82371, n82372, n82373, n82374, n82376, n82377,
    n82378, n82379, n82380, n82381, n82382, n82383, n82384, n82385, n82386,
    n82387, n82388, n82389, n82390, n82391, n82392, n82393, n82394, n82395,
    n82396, n82397, n82398, n82399, n82400, n82401, n82402, n82403, n82404,
    n82406, n82407, n82408, n82409, n82410, n82411, n82412, n82413, n82414,
    n82415, n82416, n82417, n82418, n82419, n82420, n82421, n82422, n82423,
    n82424, n82425, n82426, n82427, n82428, n82429, n82430, n82431, n82432,
    n82433, n82434, n82435, n82436, n82437, n82438, n82440, n82441, n82442,
    n82443, n82444, n82445, n82446, n82447, n82448, n82449, n82450, n82451,
    n82452, n82453, n82454, n82455, n82456, n82457, n82458, n82459, n82460,
    n82461, n82462, n82463, n82464, n82465, n82466, n82467, n82468, n82469,
    n82470, n82471, n82472, n82473, n82474, n82475, n82476, n82477, n82478,
    n82479, n82480, n82481, n82482, n82483, n82484, n82485, n82486, n82487,
    n82488, n82489, n82490, n82491, n82492, n82493, n82494, n82495, n82496,
    n82497, n82498, n82499, n82500, n82501, n82502, n82503, n82504, n82505,
    n82506, n82507, n82508, n82509, n82510, n82511, n82512, n82513, n82514,
    n82515, n82516, n82517, n82518, n82519, n82520, n82521, n82522, n82523,
    n82524, n82525, n82526, n82527, n82528, n82529, n82530, n82531, n82532,
    n82533, n82534, n82535, n82536, n82537, n82538, n82539, n82540, n82541,
    n82542, n82543, n82544, n82545, n82547, n82548, n82549, n82550, n82551,
    n82552, n82553, n82554, n82555, n82556, n82557, n82558, n82559, n82560,
    n82561, n82562, n82563, n82564, n82565, n82566, n82567, n82568, n82569,
    n82570, n82571, n82572, n82573, n82574, n82575, n82576, n82577, n82578,
    n82579, n82580, n82581, n82582, n82583, n82584, n82585, n82586, n82587,
    n82588, n82589, n82590, n82591, n82592, n82593, n82594, n82595, n82596,
    n82597, n82598, n82599, n82600, n82601, n82602, n82603, n82604, n82605,
    n82606, n82607, n82608, n82609, n82610, n82611, n82612, n82613, n82614,
    n82615, n82616, n82617, n82618, n82619, n82620, n82621, n82622, n82623,
    n82624, n82625, n82626, n82627, n82628, n82629, n82630, n82631, n82632,
    n82633, n82634, n82635, n82636, n82637, n82638, n82639, n82640, n82642,
    n82643, n82644, n82645, n82646, n82647, n82648, n82649, n82650, n82651,
    n82652, n82653, n82654, n82655, n82656, n82657, n82658, n82659, n82660,
    n82661, n82662, n82663, n82664, n82665, n82666, n82667, n82668, n82669,
    n82670, n82671, n82672, n82673, n82674, n82675, n82676, n82677, n82678,
    n82679, n82681, n82682, n82683, n82684, n82685, n82686, n82687, n82688,
    n82689, n82690, n82691, n82692, n82693, n82694, n82695, n82696, n82697,
    n82698, n82699, n82700, n82701, n82702, n82703, n82704, n82705, n82706,
    n82707, n82708, n82709, n82710, n82711, n82712, n82713, n82714, n82715,
    n82716, n82717, n82718, n82719, n82720, n82721, n82722, n82723, n82724,
    n82725, n82726, n82727, n82728, n82729, n82730, n82731, n82732, n82733,
    n82734, n82735, n82736, n82737, n82738, n82739, n82740, n82741, n82742,
    n82743, n82744, n82745, n82746, n82747, n82748, n82749, n82750, n82751,
    n82752, n82753, n82754, n82755, n82756, n82757, n82758, n82759, n82760,
    n82761, n82762, n82763, n82764, n82765, n82766, n82767, n82768, n82769,
    n82770, n82771, n82772, n82773, n82774, n82775, n82776, n82778, n82779,
    n82780, n82781, n82782, n82783, n82784, n82785, n82786, n82787, n82788,
    n82789, n82790, n82791, n82792, n82793, n82794, n82795, n82796, n82797,
    n82798, n82799, n82800, n82801, n82802, n82803, n82804, n82805, n82806,
    n82807, n82808, n82809, n82810, n82811, n82812, n82813, n82814, n82815,
    n82816, n82817, n82818, n82819, n82820, n82821, n82822, n82824, n82825,
    n82826, n82827, n82828, n82829, n82830, n82831, n82832, n82833, n82834,
    n82835, n82836, n82837, n82838, n82839, n82840, n82841, n82842, n82843,
    n82844, n82845, n82846, n82847, n82848, n82849, n82850, n82851, n82852,
    n82853, n82854, n82855, n82856, n82857, n82858, n82860, n82861, n82862,
    n82863, n82864, n82865, n82866, n82867, n82868, n82869, n82870, n82871,
    n82872, n82873, n82874, n82875, n82876, n82877, n82878, n82879, n82880,
    n82881, n82882, n82883, n82884, n82885, n82886, n82887, n82888, n82889,
    n82890, n82891, n82892, n82893, n82894, n82895, n82896, n82897, n82898,
    n82899, n82900, n82901, n82902, n82904, n82905, n82906, n82907, n82908,
    n82909, n82910, n82911, n82912, n82913, n82914, n82915, n82916, n82917,
    n82918, n82919, n82920, n82921, n82922, n82923, n82924, n82925, n82926,
    n82927, n82928, n82929, n82930, n82931, n82932, n82933, n82934, n82935,
    n82936, n82937, n82939, n82940, n82941, n82942, n82943, n82944, n82945,
    n82946, n82947, n82948, n82949, n82950, n82951, n82952, n82953, n82954,
    n82955, n82956, n82957, n82958, n82959, n82960, n82961, n82962, n82963,
    n82964, n82965, n82966, n82967, n82968, n82969, n82970, n82971, n82972,
    n82973, n82974, n82975, n82976, n82977, n82978, n82979, n82980, n82981,
    n82982, n82983, n82985, n82986, n82987, n82988, n82989, n82990, n82991,
    n82992, n82993, n82994, n82995, n82996, n82997, n82998, n82999, n83000,
    n83001, n83002, n83003, n83004, n83005, n83006, n83007, n83008, n83009,
    n83010, n83011, n83012, n83013, n83014, n83015, n83016, n83017, n83018,
    n83019, n83020, n83021, n83022, n83023, n83024, n83025, n83026, n83027,
    n83028, n83029, n83030, n83032, n83033, n83034, n83035, n83036, n83037,
    n83038, n83039, n83040, n83041, n83042, n83043, n83044, n83045, n83046,
    n83047, n83048, n83049, n83050, n83051, n83052, n83053, n83054, n83055,
    n83056, n83057, n83058, n83059, n83060, n83061, n83062, n83063, n83064,
    n83065, n83066, n83068, n83069, n83070, n83071, n83072, n83073, n83074,
    n83075, n83076, n83077, n83078, n83079, n83080, n83081, n83082, n83083,
    n83084, n83085, n83086, n83087, n83088, n83089, n83090, n83091, n83092,
    n83094, n83095, n83096, n83097, n83098, n83099, n83100, n83101, n83102,
    n83103, n83104, n83105, n83106, n83107, n83108, n83109, n83110, n83111,
    n83112, n83113, n83114, n83115, n83116, n83117, n83118, n83119, n83120,
    n83121, n83122, n83123, n83124, n83125, n83126, n83127, n83129, n83130,
    n83131, n83132, n83133, n83134, n83135, n83136, n83137, n83138, n83139,
    n83140, n83141, n83142, n83143, n83144, n83145, n83146, n83147, n83148,
    n83149, n83150, n83151, n83152, n83153, n83154, n83155, n83156, n83157,
    n83158, n83159, n83160, n83161, n83163, n83164, n83165, n83166, n83167,
    n83168, n83169, n83170, n83171, n83172, n83173, n83174, n83175, n83176,
    n83177, n83178, n83179, n83180, n83181, n83182, n83183, n83184, n83185,
    n83186, n83187, n83188, n83189, n83190, n83191, n83193, n83194, n83195,
    n83196, n83197, n83198, n83199, n83200, n83201, n83202, n83203, n83204,
    n83205, n83206, n83207, n83208, n83209, n83210, n83211, n83212, n83213,
    n83214, n83215, n83216, n83217, n83218, n83219, n83220, n83221, n83223,
    n83224, n83225, n83226, n83227, n83228, n83229, n83230, n83231, n83232,
    n83233, n83234, n83235, n83236, n83237, n83238, n83239, n83240, n83241,
    n83242, n83243, n83244, n83245, n83246, n83247, n83248, n83249, n83250,
    n83251, n83252, n83253, n83254, n83255, n83256, n83257, n83258, n83259,
    n83260, n83261, n83262, n83263, n83264, n83265, n83266, n83267, n83268,
    n83269, n83270, n83271, n83272, n83273, n83274, n83275, n83276, n83277,
    n83278, n83279, n83280, n83281, n83282, n83283, n83284, n83285, n83286,
    n83287, n83288, n83289, n83290, n83291, n83292, n83293, n83294, n83295,
    n83296, n83297, n83298, n83299, n83300, n83301, n83302, n83303, n83304,
    n83305, n83306, n83307, n83308, n83309, n83310, n83311, n83312, n83313,
    n83314, n83315, n83316, n83317, n83318, n83319, n83320, n83322, n83323,
    n83324, n83325, n83326, n83327, n83328, n83329, n83330, n83331, n83332,
    n83333, n83334, n83335, n83336, n83337, n83338, n83339, n83340, n83341,
    n83342, n83343, n83344, n83345, n83346, n83347, n83348, n83349, n83350,
    n83351, n83352, n83353, n83354, n83355, n83356, n83357, n83358, n83359,
    n83360, n83362, n83363, n83364, n83365, n83366, n83367, n83368, n83369,
    n83370, n83371, n83372, n83373, n83374, n83375, n83376, n83377, n83378,
    n83379, n83380, n83381, n83382, n83383, n83384, n83385, n83386, n83387,
    n83388, n83389, n83390, n83391, n83392, n83393, n83394, n83395, n83396,
    n83397, n83398, n83399, n83400, n83401, n83402, n83403, n83404, n83405,
    n83406, n83407, n83408, n83409, n83410, n83411, n83412, n83413, n83414,
    n83415, n83416, n83417, n83418, n83419, n83420, n83421, n83422, n83423,
    n83424, n83425, n83426, n83427, n83428, n83429, n83430, n83431, n83432,
    n83433, n83434, n83435, n83436, n83437, n83438, n83439, n83440, n83441,
    n83442, n83443, n83444, n83445, n83446, n83447, n83448, n83449, n83450,
    n83451, n83452, n83453, n83454, n83455, n83456, n83457, n83458, n83459,
    n83461, n83462, n83463, n83464, n83465, n83466, n83467, n83468, n83469,
    n83470, n83471, n83472, n83473, n83474, n83475, n83476, n83477, n83478,
    n83479, n83480, n83481, n83482, n83483, n83484, n83485, n83486, n83487,
    n83488, n83489, n83490, n83491, n83492, n83493, n83494, n83495, n83496,
    n83497, n83499, n83500, n83501, n83502, n83503, n83504, n83505, n83506,
    n83507, n83508, n83509, n83510, n83511, n83512, n83513, n83514, n83515,
    n83516, n83517, n83518, n83519, n83520, n83521, n83522, n83523, n83524,
    n83525, n83526, n83527, n83528, n83529, n83530, n83531, n83532, n83533,
    n83534, n83536, n83537, n83538, n83539, n83540, n83541, n83542, n83543,
    n83544, n83545, n83546, n83547, n83548, n83549, n83550, n83551, n83552,
    n83553, n83554, n83555, n83556, n83557, n83558, n83559, n83560, n83561,
    n83562, n83563, n83564, n83565, n83566, n83567, n83568, n83569, n83570,
    n83571, n83572, n83573, n83574, n83575, n83576, n83577, n83578, n83579,
    n83580, n83581, n83582, n83583, n83584, n83585, n83586, n83587, n83588,
    n83589, n83590, n83591, n83592, n83593, n83594, n83595, n83596, n83597,
    n83598, n83599, n83600, n83601, n83602, n83603, n83604, n83605, n83606,
    n83607, n83608, n83609, n83610, n83611, n83612, n83613, n83614, n83615,
    n83616, n83617, n83618, n83619, n83620, n83621, n83622, n83623, n83624,
    n83625, n83626, n83627, n83628, n83629, n83630, n83631, n83632, n83633,
    n83634, n83635, n83636, n83638, n83639, n83640, n83641, n83642, n83643,
    n83644, n83645, n83646, n83647, n83648, n83649, n83650, n83651, n83652,
    n83653, n83654, n83655, n83656, n83657, n83658, n83659, n83660, n83661,
    n83662, n83663, n83664, n83665, n83666, n83667, n83668, n83669, n83670,
    n83671, n83672, n83673, n83674, n83675, n83676, n83677, n83678, n83679,
    n83680, n83681, n83682, n83683, n83684, n83685, n83686, n83687, n83688,
    n83689, n83690, n83691, n83692, n83693, n83694, n83695, n83696, n83697,
    n83698, n83699, n83700, n83701, n83702, n83703, n83704, n83705, n83706,
    n83707, n83708, n83709, n83710, n83711, n83712, n83713, n83714, n83715,
    n83716, n83717, n83718, n83719, n83720, n83721, n83722, n83723, n83724,
    n83725, n83726, n83727, n83728, n83729, n83730, n83731, n83732, n83733,
    n83734, n83735, n83736, n83737, n83739, n83740, n83741, n83742, n83743,
    n83744, n83745, n83746, n83747, n83748, n83749, n83750, n83751, n83752,
    n83753, n83754, n83755, n83756, n83757, n83758, n83759, n83760, n83761,
    n83762, n83763, n83764, n83765, n83766, n83767, n83768, n83769, n83770,
    n83771, n83772, n83773, n83774, n83775, n83776, n83777, n83778, n83779,
    n83780, n83781, n83782, n83783, n83784, n83785, n83786, n83787, n83788,
    n83789, n83790, n83791, n83792, n83793, n83794, n83795, n83796, n83797,
    n83798, n83799, n83800, n83801, n83802, n83803, n83804, n83805, n83806,
    n83807, n83808, n83809, n83810, n83811, n83812, n83813, n83814, n83815,
    n83816, n83817, n83818, n83819, n83820, n83821, n83822, n83823, n83824,
    n83825, n83826, n83827, n83828, n83829, n83830, n83831, n83832, n83833,
    n83834, n83835, n83836, n83837, n83839, n83840, n83841, n83842, n83843,
    n83844, n83845, n83846, n83847, n83848, n83849, n83850, n83851, n83852,
    n83853, n83854, n83855, n83856, n83857, n83858, n83859, n83860, n83861,
    n83862, n83863, n83864, n83865, n83866, n83867, n83868, n83869, n83870,
    n83871, n83872, n83873, n83874, n83875, n83876, n83877, n83878, n83879,
    n83880, n83881, n83882, n83883, n83884, n83885, n83887, n83888, n83889,
    n83890, n83891, n83892, n83893, n83894, n83895, n83896, n83897, n83898,
    n83899, n83900, n83901, n83902, n83903, n83904, n83905, n83906, n83907,
    n83908, n83909, n83910, n83911, n83912, n83913, n83914, n83915, n83916,
    n83917, n83918, n83920, n83921, n83922, n83923, n83924, n83925, n83926,
    n83927, n83928, n83929, n83930, n83931, n83932, n83933, n83934, n83935,
    n83936, n83937, n83938, n83939, n83940, n83941, n83942, n83943, n83944,
    n83945, n83946, n83947, n83948, n83949, n83950, n83951, n83952, n83954,
    n83955, n83956, n83957, n83958, n83959, n83960, n83961, n83962, n83963,
    n83964, n83965, n83966, n83967, n83968, n83969, n83970, n83971, n83972,
    n83973, n83974, n83975, n83976, n83977, n83978, n83979, n83980, n83981,
    n83982, n83983, n83984, n83985, n83986, n83987, n83988, n83989, n83990,
    n83991, n83992, n83994, n83995, n83996, n83997, n83998, n83999, n84000,
    n84001, n84002, n84003, n84004, n84005, n84006, n84007, n84008, n84009,
    n84010, n84011, n84012, n84013, n84014, n84015, n84016, n84017, n84018,
    n84019, n84020, n84021, n84022, n84023, n84024, n84025, n84026, n84027,
    n84028, n84029, n84030, n84031, n84032, n84033, n84034, n84035, n84036,
    n84037, n84038, n84039, n84040, n84041, n84042, n84043, n84044, n84045,
    n84046, n84047, n84048, n84049, n84050, n84051, n84052, n84053, n84054,
    n84055, n84056, n84057, n84058, n84059, n84060, n84061, n84062, n84063,
    n84064, n84065, n84066, n84067, n84068, n84069, n84070, n84071, n84072,
    n84073, n84074, n84075, n84076, n84077, n84078, n84079, n84080, n84081,
    n84082, n84083, n84084, n84085, n84086, n84087, n84088, n84089, n84090,
    n84091, n84092, n84093, n84094, n84095, n84096, n84097, n84098, n84099,
    n84101, n84102, n84103, n84104, n84105, n84106, n84107, n84108, n84109,
    n84110, n84111, n84112, n84113, n84114, n84115, n84116, n84117, n84118,
    n84119, n84120, n84121, n84122, n84123, n84124, n84125, n84126, n84127,
    n84128, n84129, n84130, n84131, n84132, n84133, n84134, n84136, n84137,
    n84138, n84139, n84140, n84141, n84142, n84143, n84144, n84145, n84146,
    n84147, n84148, n84149, n84150, n84151, n84152, n84153, n84154, n84155,
    n84156, n84157, n84158, n84159, n84160, n84161, n84162, n84163, n84164,
    n84165, n84166, n84167, n84168, n84169, n84170, n84171, n84172, n84173,
    n84174, n84175, n84177, n84178, n84179, n84180, n84181, n84182, n84183,
    n84184, n84185, n84186, n84187, n84188, n84189, n84190, n84191, n84192,
    n84193, n84194, n84195, n84196, n84197, n84198, n84199, n84200, n84201,
    n84202, n84203, n84204, n84205, n84206, n84207, n84208, n84209, n84210,
    n84211, n84212, n84213, n84214, n84215, n84216, n84217, n84218, n84219,
    n84221, n84222, n84223, n84224, n84225, n84226, n84227, n84228, n84229,
    n84230, n84231, n84232, n84233, n84234, n84235, n84236, n84237, n84238,
    n84239, n84240, n84241, n84242, n84243, n84244, n84245, n84246, n84247,
    n84248, n84249, n84250, n84251, n84252, n84253, n84254, n84255, n84256,
    n84258, n84259, n84260, n84261, n84262, n84263, n84264, n84265, n84266,
    n84267, n84268, n84269, n84270, n84271, n84272, n84273, n84274, n84275,
    n84276, n84277, n84278, n84279, n84280, n84281, n84282, n84283, n84284,
    n84285, n84286, n84287, n84288, n84289, n84290, n84291, n84292, n84293,
    n84294, n84295, n84296, n84297, n84298, n84299, n84300, n84301, n84302,
    n84303, n84304, n84305, n84306, n84307, n84308, n84309, n84310, n84311,
    n84312, n84313, n84314, n84315, n84316, n84317, n84318, n84319, n84320,
    n84321, n84322, n84323, n84324, n84325, n84326, n84327, n84328, n84329,
    n84330, n84331, n84332, n84333, n84334, n84335, n84336, n84337, n84338,
    n84339, n84340, n84341, n84342, n84343, n84344, n84345, n84346, n84347,
    n84348, n84349, n84350, n84351, n84352, n84353, n84354, n84356, n84357,
    n84358, n84359, n84360, n84361, n84362, n84363, n84364, n84365, n84366,
    n84367, n84368, n84369, n84370, n84371, n84372, n84373, n84374, n84375,
    n84376, n84377, n84378, n84379, n84380, n84381, n84382, n84383, n84384,
    n84385, n84386, n84387, n84388, n84389, n84390, n84391, n84392, n84393,
    n84395, n84396, n84397, n84398, n84399, n84400, n84401, n84402, n84403,
    n84404, n84405, n84406, n84407, n84408, n84409, n84410, n84411, n84412,
    n84413, n84414, n84415, n84416, n84417, n84418, n84419, n84420, n84421,
    n84422, n84423, n84424, n84425, n84426, n84427, n84428, n84429, n84430,
    n84431, n84432, n84433, n84434, n84435, n84436, n84437, n84438, n84439,
    n84440, n84441, n84442, n84443, n84444, n84445, n84446, n84447, n84448,
    n84449, n84450, n84451, n84452, n84453, n84454, n84455, n84456, n84457,
    n84458, n84459, n84460, n84461, n84462, n84463, n84464, n84465, n84466,
    n84467, n84468, n84469, n84470, n84471, n84472, n84473, n84474, n84475,
    n84476, n84477, n84478, n84479, n84480, n84481, n84482, n84483, n84485,
    n84486, n84487, n84488, n84489, n84490, n84491, n84492, n84493, n84494,
    n84495, n84496, n84497, n84498, n84499, n84500, n84501, n84502, n84503,
    n84504, n84505, n84506, n84507, n84508, n84509, n84510, n84511, n84512,
    n84513, n84514, n84515, n84516, n84517, n84518, n84519, n84520, n84521,
    n84522, n84523, n84524, n84525, n84526, n84527, n84528, n84529, n84531,
    n84532, n84533, n84534, n84535, n84536, n84537, n84538, n84539, n84540,
    n84541, n84542, n84543, n84544, n84545, n84546, n84547, n84548, n84549,
    n84550, n84551, n84552, n84553, n84554, n84555, n84556, n84557, n84558,
    n84559, n84560, n84561, n84562, n84563, n84564, n84566, n84567, n84568,
    n84569, n84570, n84571, n84572, n84573, n84574, n84575, n84576, n84577,
    n84578, n84579, n84580, n84581, n84582, n84583, n84584, n84585, n84586,
    n84587, n84588, n84589, n84590, n84591, n84592, n84593, n84594, n84595,
    n84596, n84597, n84598, n84599, n84600, n84601, n84602, n84603, n84604,
    n84605, n84607, n84608, n84609, n84610, n84611, n84612, n84613, n84614,
    n84615, n84616, n84617, n84618, n84619, n84620, n84621, n84622, n84623,
    n84624, n84625, n84626, n84627, n84628, n84629, n84630, n84631, n84632,
    n84633, n84634, n84635, n84636, n84637, n84638, n84639, n84640, n84641,
    n84642, n84643, n84644, n84645, n84646, n84647, n84648, n84649, n84650,
    n84651, n84652, n84653, n84654, n84655, n84656, n84658, n84659, n84660,
    n84661, n84662, n84663, n84664, n84665, n84666, n84667, n84668, n84669,
    n84670, n84671, n84672, n84673, n84674, n84675, n84676, n84677, n84678,
    n84679, n84680, n84681, n84682, n84683, n84684, n84685, n84686, n84687,
    n84688, n84689, n84690, n84691, n84693, n84694, n84695, n84696, n84697,
    n84698, n84699, n84700, n84701, n84702, n84703, n84704, n84705, n84706,
    n84707, n84708, n84709, n84710, n84711, n84712, n84713, n84714, n84715,
    n84716, n84717, n84718, n84719, n84720, n84721, n84722, n84723, n84724,
    n84725, n84726, n84727, n84728, n84729, n84730, n84731, n84733, n84734,
    n84735, n84736, n84737, n84738, n84739, n84740, n84741, n84742, n84743,
    n84744, n84745, n84746, n84747, n84748, n84749, n84750, n84751, n84752,
    n84753, n84754, n84755, n84756, n84757, n84758, n84759, n84760, n84761,
    n84762, n84763, n84764, n84765, n84766, n84767, n84768, n84769, n84770,
    n84771, n84772, n84773, n84774, n84775, n84776, n84777, n84779, n84780,
    n84781, n84782, n84783, n84784, n84785, n84786, n84787, n84788, n84789,
    n84790, n84791, n84792, n84793, n84794, n84795, n84796, n84797, n84798,
    n84799, n84800, n84801, n84802, n84803, n84804, n84805, n84806, n84807,
    n84809, n84810, n84811, n84812, n84813, n84814, n84815, n84816, n84817,
    n84818, n84819, n84820, n84821, n84822, n84823, n84824, n84825, n84826,
    n84827, n84828, n84829, n84830, n84831, n84832, n84833, n84834, n84835,
    n84836, n84837, n84839, n84840, n84841, n84842, n84843, n84844, n84845,
    n84846, n84847, n84848, n84849, n84850, n84851, n84852, n84853, n84854,
    n84855, n84856, n84857, n84858, n84859, n84860, n84861, n84862, n84863,
    n84864, n84865, n84866, n84867, n84868, n84869, n84870, n84871, n84872,
    n84873, n84874, n84875, n84877, n84878, n84879, n84880, n84881, n84882,
    n84883, n84884, n84885, n84886, n84887, n84888, n84889, n84890, n84891,
    n84892, n84893, n84894, n84895, n84896, n84897, n84898, n84899, n84900,
    n84901, n84902, n84903, n84904, n84905, n84906, n84907, n84908, n84909,
    n84911, n84912, n84913, n84914, n84915, n84916, n84917, n84918, n84919,
    n84920, n84921, n84922, n84923, n84924, n84925, n84926, n84927, n84928,
    n84929, n84930, n84931, n84932, n84933, n84934, n84935, n84937, n84938,
    n84939, n84940, n84941, n84942, n84943, n84944, n84945, n84946, n84947,
    n84948, n84949, n84950, n84951, n84952, n84953, n84954, n84955, n84956,
    n84957, n84958, n84959, n84960, n84961, n84962, n84963, n84964, n84965,
    n84966, n84967, n84968, n84969, n84970, n84971, n84972, n84973, n84974,
    n84975, n84976, n84977, n84978, n84979, n84980, n84981, n84982, n84983,
    n84984, n84985, n84986, n84987, n84988, n84989, n84990, n84991, n84992,
    n84993, n84994, n84995, n84996, n84997, n84998, n84999, n85000, n85001,
    n85002, n85003, n85004, n85005, n85006, n85007, n85008, n85009, n85010,
    n85011, n85012, n85013, n85014, n85015, n85016, n85017, n85018, n85019,
    n85020, n85021, n85022, n85023, n85024, n85025, n85026, n85027, n85028,
    n85029, n85030, n85031, n85032, n85033, n85034, n85035, n85036, n85037,
    n85039, n85040, n85041, n85042, n85043, n85044, n85045, n85046, n85047,
    n85048, n85049, n85050, n85051, n85052, n85053, n85054, n85055, n85056,
    n85057, n85058, n85059, n85060, n85061, n85062, n85063, n85064, n85065,
    n85066, n85067, n85068, n85069, n85070, n85071, n85072, n85073, n85074,
    n85075, n85076, n85077, n85078, n85079, n85080, n85081, n85082, n85083,
    n85084, n85086, n85087, n85088, n85089, n85090, n85091, n85092, n85093,
    n85094, n85095, n85096, n85097, n85098, n85099, n85100, n85101, n85102,
    n85103, n85104, n85105, n85106, n85107, n85108, n85109, n85110, n85111,
    n85112, n85113, n85114, n85115, n85116, n85117, n85118, n85120, n85121,
    n85122, n85123, n85124, n85125, n85126, n85127, n85128, n85129, n85130,
    n85131, n85132, n85133, n85134, n85135, n85136, n85137, n85138, n85139,
    n85140, n85141, n85142, n85143, n85144, n85145, n85146, n85147, n85148,
    n85149, n85150, n85151, n85152, n85153, n85154, n85155, n85156, n85157,
    n85158, n85159, n85160, n85161, n85162, n85163, n85164, n85165, n85166,
    n85167, n85168, n85169, n85170, n85171, n85172, n85173, n85174, n85175,
    n85176, n85177, n85178, n85179, n85180, n85181, n85182, n85183, n85184,
    n85185, n85186, n85187, n85188, n85189, n85190, n85191, n85192, n85193,
    n85194, n85195, n85196, n85197, n85198, n85199, n85200, n85201, n85202,
    n85203, n85204, n85205, n85206, n85207, n85208, n85209, n85210, n85211,
    n85212, n85213, n85214, n85215, n85216, n85217, n85218, n85219, n85220,
    n85221, n85222, n85224, n85225, n85226, n85227, n85228, n85229, n85230,
    n85231, n85232, n85233, n85234, n85235, n85236, n85237, n85238, n85239,
    n85240, n85241, n85242, n85243, n85244, n85245, n85246, n85247, n85248,
    n85249, n85250, n85251, n85252, n85253, n85254, n85255, n85256, n85257,
    n85258, n85259, n85260, n85261, n85262, n85263, n85264, n85265, n85266,
    n85267, n85268, n85269, n85270, n85271, n85272, n85273, n85274, n85275,
    n85276, n85277, n85278, n85279, n85280, n85281, n85282, n85283, n85284,
    n85285, n85286, n85287, n85288, n85289, n85290, n85291, n85292, n85293,
    n85294, n85295, n85296, n85297, n85298, n85299, n85300, n85301, n85302,
    n85303, n85304, n85305, n85306, n85307, n85308, n85309, n85310, n85311,
    n85312, n85313, n85314, n85315, n85316, n85317, n85318, n85319, n85320,
    n85321, n85322, n85323, n85325, n85326, n85327, n85328, n85329, n85330,
    n85331, n85332, n85333, n85334, n85335, n85336, n85337, n85338, n85339,
    n85340, n85341, n85342, n85343, n85344, n85345, n85346, n85347, n85348,
    n85349, n85350, n85351, n85352, n85353, n85354, n85355, n85356, n85357,
    n85358, n85359, n85360, n85361, n85362, n85363, n85364, n85365, n85366,
    n85367, n85368, n85369, n85370, n85371, n85372, n85373, n85374, n85375,
    n85376, n85377, n85378, n85379, n85380, n85381, n85382, n85383, n85384,
    n85385, n85386, n85387, n85388, n85389, n85390, n85391, n85392, n85393,
    n85394, n85395, n85396, n85397, n85398, n85399, n85400, n85401, n85402,
    n85403, n85404, n85405, n85406, n85407, n85408, n85409, n85410, n85411,
    n85412, n85413, n85414, n85415, n85417, n85418, n85419, n85420, n85421,
    n85422, n85423, n85424, n85425, n85426, n85427, n85428, n85429, n85430,
    n85431, n85432, n85433, n85434, n85435, n85436, n85437, n85438, n85439,
    n85440, n85441, n85442, n85443, n85444, n85445, n85446, n85447, n85448,
    n85449, n85450, n85451, n85453, n85454, n85455, n85456, n85457, n85458,
    n85459, n85460, n85461, n85462, n85463, n85464, n85465, n85466, n85467,
    n85468, n85469, n85470, n85471, n85472, n85473, n85474, n85475, n85476,
    n85477, n85478, n85479, n85480, n85481, n85482, n85483, n85484, n85485,
    n85486, n85487, n85488, n85489, n85490, n85491, n85492, n85493, n85494,
    n85495, n85496, n85497, n85498, n85499, n85500, n85501, n85502, n85503,
    n85504, n85505, n85506, n85507, n85508, n85509, n85510, n85511, n85512,
    n85513, n85514, n85515, n85516, n85517, n85518, n85519, n85520, n85521,
    n85522, n85523, n85524, n85525, n85526, n85527, n85528, n85529, n85530,
    n85531, n85532, n85533, n85534, n85535, n85536, n85537, n85538, n85539,
    n85540, n85541, n85542, n85543, n85544, n85545, n85546, n85548, n85549,
    n85550, n85551, n85552, n85553, n85554, n85555, n85556, n85557, n85558,
    n85559, n85560, n85561, n85562, n85563, n85564, n85565, n85566, n85567,
    n85568, n85569, n85570, n85571, n85572, n85573, n85574, n85575, n85576,
    n85577, n85578, n85579, n85580, n85581, n85582, n85583, n85584, n85585,
    n85586, n85587, n85588, n85590, n85591, n85592, n85593, n85594, n85595,
    n85596, n85597, n85598, n85599, n85600, n85601, n85602, n85603, n85604,
    n85605, n85606, n85607, n85608, n85609, n85610, n85611, n85612, n85613,
    n85614, n85615, n85616, n85617, n85618, n85619, n85620, n85621, n85622,
    n85623, n85624, n85625, n85626, n85627, n85628, n85629, n85630, n85631,
    n85632, n85633, n85634, n85635, n85636, n85637, n85638, n85639, n85640,
    n85641, n85642, n85643, n85645, n85646, n85647, n85648, n85649, n85650,
    n85651, n85652, n85653, n85654, n85655, n85656, n85657, n85658, n85659,
    n85660, n85661, n85662, n85663, n85664, n85665, n85666, n85667, n85668,
    n85669, n85670, n85671, n85672, n85673, n85674, n85675, n85676, n85677,
    n85678, n85679, n85680, n85681, n85682, n85683, n85684, n85685, n85686,
    n85687, n85688, n85689, n85690, n85691, n85692, n85693, n85694, n85695,
    n85696, n85697, n85698, n85699, n85700, n85701, n85702, n85703, n85704,
    n85705, n85706, n85707, n85708, n85709, n85710, n85711, n85712, n85713,
    n85714, n85715, n85716, n85717, n85718, n85719, n85720, n85721, n85722,
    n85723, n85724, n85725, n85726, n85727, n85728, n85729, n85730, n85731,
    n85732, n85733, n85734, n85735, n85736, n85737, n85738, n85739, n85740,
    n85741, n85742, n85743, n85744, n85745, n85746, n85748, n85749, n85750,
    n85751, n85752, n85753, n85754, n85755, n85756, n85757, n85758, n85759,
    n85760, n85761, n85762, n85763, n85764, n85765, n85766, n85767, n85768,
    n85769, n85770, n85771, n85772, n85773, n85774, n85775, n85776, n85777,
    n85778, n85779, n85780, n85781, n85782, n85783, n85785, n85786, n85787,
    n85788, n85789, n85790, n85791, n85792, n85793, n85794, n85795, n85796,
    n85797, n85798, n85799, n85800, n85801, n85802, n85803, n85804, n85805,
    n85806, n85807, n85808, n85809, n85810, n85811, n85812, n85813, n85814,
    n85815, n85816, n85817, n85818, n85819, n85820, n85821, n85822, n85823,
    n85824, n85825, n85826, n85827, n85828, n85829, n85830, n85831, n85832,
    n85833, n85834, n85835, n85836, n85837, n85838, n85839, n85840, n85841,
    n85842, n85843, n85844, n85845, n85846, n85847, n85848, n85849, n85850,
    n85851, n85852, n85853, n85854, n85855, n85856, n85857, n85858, n85859,
    n85860, n85861, n85862, n85863, n85864, n85865, n85866, n85867, n85868,
    n85869, n85870, n85871, n85872, n85873, n85874, n85875, n85876, n85877,
    n85878, n85879, n85880, n85881, n85882, n85883, n85885, n85886, n85887,
    n85888, n85889, n85890, n85891, n85892, n85893, n85894, n85895, n85896,
    n85897, n85898, n85899, n85900, n85901, n85902, n85903, n85904, n85905,
    n85906, n85907, n85908, n85909, n85910, n85911, n85912, n85914, n85915,
    n85916, n85917, n85918, n85919, n85920, n85921, n85922, n85923, n85924,
    n85925, n85926, n85927, n85928, n85929, n85930, n85931, n85932, n85933,
    n85934, n85935, n85936, n85937, n85938, n85939, n85940, n85941, n85942,
    n85944, n85945, n85946, n85947, n85948, n85949, n85950, n85951, n85952,
    n85953, n85954, n85955, n85956, n85957, n85958, n85959, n85960, n85961,
    n85962, n85963, n85964, n85965, n85966, n85967, n85968, n85969, n85970,
    n85971, n85972, n85973, n85974, n85976, n85977, n85978, n85979, n85980,
    n85981, n85982, n85983, n85984, n85985, n85986, n85987, n85988, n85989,
    n85990, n85991, n85992, n85993, n85994, n85995, n85996, n85997, n85998,
    n85999, n86000, n86001, n86002, n86003, n86004, n86005, n86006, n86007,
    n86008, n86009, n86010, n86011, n86012, n86013, n86014, n86015, n86016,
    n86017, n86018, n86020, n86021, n86022, n86023, n86024, n86025, n86026,
    n86027, n86028, n86029, n86030, n86031, n86032, n86033, n86034, n86035,
    n86036, n86037, n86038, n86039, n86040, n86041, n86042, n86043, n86044,
    n86045, n86046, n86047, n86048, n86049, n86050, n86051, n86052, n86053,
    n86054, n86055, n86056, n86057, n86058, n86059, n86060, n86061, n86062,
    n86063, n86064, n86065, n86067, n86068, n86069, n86070, n86071, n86072,
    n86073, n86074, n86075, n86076, n86077, n86078, n86079, n86080, n86081,
    n86082, n86083, n86084, n86085, n86086, n86087, n86088, n86089, n86090,
    n86091, n86092, n86093, n86094, n86095, n86096, n86097, n86098, n86099,
    n86100, n86101, n86102, n86103, n86105, n86106, n86107, n86108, n86109,
    n86110, n86111, n86112, n86113, n86114, n86115, n86116, n86117, n86118,
    n86119, n86120, n86121, n86122, n86123, n86124, n86125, n86126, n86127,
    n86128, n86129, n86130, n86131, n86132, n86133, n86134, n86135, n86136,
    n86137, n86138, n86139, n86140, n86141, n86142, n86143, n86145, n86146,
    n86147, n86148, n86149, n86150, n86151, n86152, n86153, n86154, n86155,
    n86156, n86157, n86158, n86159, n86160, n86161, n86162, n86163, n86164,
    n86165, n86166, n86167, n86168, n86169, n86170, n86171, n86172, n86173,
    n86174, n86175, n86176, n86177, n86178, n86179, n86180, n86181, n86182,
    n86183, n86184, n86186, n86187, n86188, n86189, n86190, n86191, n86192,
    n86193, n86194, n86195, n86196, n86197, n86198, n86199, n86200, n86201,
    n86202, n86203, n86204, n86205, n86206, n86207, n86208, n86209, n86210,
    n86211, n86212, n86213, n86214, n86215, n86216, n86217, n86218, n86219,
    n86220, n86221, n86222, n86223, n86224, n86225, n86226, n86227, n86228,
    n86229, n86230, n86231, n86233, n86234, n86235, n86236, n86237, n86238,
    n86239, n86240, n86241, n86242, n86243, n86244, n86245, n86246, n86247,
    n86248, n86249, n86250, n86251, n86252, n86253, n86254, n86255, n86256,
    n86257, n86258, n86259, n86260, n86261, n86262, n86263, n86264, n86265,
    n86266, n86267, n86268, n86269, n86270, n86271, n86272, n86273, n86274,
    n86275, n86276, n86277, n86278, n86279, n86281, n86282, n86283, n86284,
    n86285, n86286, n86287, n86288, n86289, n86290, n86291, n86292, n86293,
    n86294, n86295, n86296, n86297, n86298, n86299, n86300, n86301, n86302,
    n86303, n86304, n86305, n86306, n86307, n86308, n86309, n86310, n86311,
    n86312, n86313, n86314, n86315, n86316, n86317, n86318, n86319, n86320,
    n86321, n86322, n86323, n86324, n86325, n86326, n86327, n86328, n86329,
    n86330, n86331, n86332, n86333, n86334, n86335, n86336, n86337, n86338,
    n86339, n86340, n86341, n86342, n86343, n86344, n86345, n86346, n86347,
    n86348, n86349, n86350, n86351, n86352, n86353, n86354, n86355, n86356,
    n86357, n86358, n86359, n86360, n86361, n86362, n86363, n86364, n86365,
    n86366, n86367, n86368, n86369, n86370, n86371, n86372, n86373, n86374,
    n86375, n86376, n86377, n86379, n86380, n86381, n86382, n86383, n86384,
    n86385, n86386, n86387, n86388, n86389, n86390, n86391, n86392, n86393,
    n86394, n86395, n86396, n86397, n86398, n86399, n86400, n86401, n86402,
    n86403, n86404, n86405, n86406, n86407, n86408, n86409, n86410, n86411,
    n86412, n86413, n86414, n86416, n86417, n86418, n86419, n86420, n86421,
    n86422, n86423, n86424, n86425, n86426, n86427, n86428, n86429, n86430,
    n86431, n86432, n86433, n86434, n86435, n86436, n86437, n86438, n86439,
    n86440, n86441, n86442, n86443, n86444, n86446, n86447, n86448, n86449,
    n86450, n86451, n86452, n86453, n86454, n86455, n86456, n86457, n86458,
    n86459, n86460, n86461, n86462, n86463, n86464, n86465, n86466, n86467,
    n86468, n86469, n86470, n86471, n86472, n86473, n86474, n86475, n86476,
    n86477, n86478, n86479, n86480, n86481, n86482, n86483, n86484, n86485,
    n86486, n86487, n86488, n86490, n86491, n86492, n86493, n86494, n86495,
    n86496, n86497, n86498, n86499, n86500, n86501, n86502, n86503, n86504,
    n86505, n86506, n86507, n86508, n86509, n86510, n86511, n86512, n86513,
    n86514, n86515, n86516, n86517, n86518, n86519, n86520, n86521, n86522,
    n86523, n86525, n86526, n86527, n86528, n86529, n86530, n86531, n86532,
    n86533, n86534, n86535, n86536, n86537, n86538, n86539, n86540, n86541,
    n86542, n86543, n86544, n86545, n86546, n86547, n86548, n86549, n86550,
    n86551, n86552, n86553, n86554, n86555, n86556, n86557, n86558, n86560,
    n86561, n86562, n86563, n86564, n86565, n86566, n86567, n86568, n86569,
    n86570, n86571, n86572, n86573, n86574, n86575, n86576, n86577, n86578,
    n86579, n86580, n86581, n86582, n86583, n86584, n86585, n86586, n86587,
    n86588, n86589, n86590, n86591, n86592, n86593, n86594, n86595, n86596,
    n86598, n86599, n86600, n86601, n86602, n86603, n86604, n86605, n86606,
    n86607, n86608, n86609, n86610, n86611, n86612, n86613, n86614, n86615,
    n86616, n86617, n86618, n86619, n86620, n86621, n86622, n86623, n86625,
    n86626, n86627, n86628, n86629, n86630, n86631, n86632, n86633, n86634,
    n86635, n86636, n86637, n86638, n86639, n86640, n86641, n86642, n86643,
    n86644, n86645, n86646, n86647, n86648, n86649, n86650, n86651, n86652,
    n86653, n86654, n86655, n86656, n86658, n86659, n86660, n86661, n86662,
    n86663, n86664, n86665, n86666, n86667, n86668, n86669, n86670, n86671,
    n86672, n86673, n86674, n86675, n86676, n86677, n86678, n86679, n86680,
    n86681, n86682, n86683, n86684, n86685, n86686, n86687, n86688, n86689,
    n86690, n86691, n86692, n86693, n86694, n86695, n86696, n86697, n86698,
    n86699, n86700, n86701, n86702, n86703, n86704, n86705, n86706, n86707,
    n86708, n86709, n86710, n86711, n86712, n86713, n86714, n86715, n86716,
    n86717, n86718, n86719, n86720, n86721, n86722, n86723, n86724, n86725,
    n86726, n86727, n86728, n86729, n86730, n86731, n86732, n86733, n86734,
    n86735, n86736, n86737, n86738, n86739, n86740, n86741, n86742, n86743,
    n86744, n86745, n86746, n86747, n86748, n86749, n86750, n86751, n86752,
    n86753, n86754, n86755, n86756, n86757, n86758, n86760, n86761, n86762,
    n86763, n86764, n86765, n86766, n86767, n86768, n86769, n86770, n86771,
    n86772, n86773, n86774, n86775, n86776, n86777, n86778, n86779, n86780,
    n86781, n86782, n86783, n86784, n86785, n86786, n86787, n86788, n86789,
    n86790, n86791, n86792, n86793, n86794, n86795, n86796, n86797, n86798,
    n86799, n86800, n86801, n86802, n86803, n86804, n86805, n86806, n86807,
    n86808, n86809, n86810, n86811, n86812, n86813, n86814, n86815, n86816,
    n86817, n86818, n86819, n86820, n86821, n86822, n86823, n86824, n86825,
    n86826, n86827, n86828, n86829, n86830, n86831, n86832, n86833, n86834,
    n86835, n86836, n86837, n86838, n86839, n86840, n86841, n86842, n86843,
    n86844, n86845, n86846, n86847, n86848, n86849, n86850, n86851, n86852,
    n86853, n86854, n86855, n86856, n86857, n86858, n86859, n86860, n86861,
    n86863, n86864, n86865, n86866, n86867, n86868, n86869, n86870, n86871,
    n86872, n86873, n86874, n86875, n86876, n86877, n86878, n86879, n86880,
    n86881, n86882, n86883, n86884, n86885, n86886, n86887, n86888, n86889,
    n86890, n86891, n86892, n86893, n86894, n86896, n86897, n86898, n86899,
    n86900, n86901, n86902, n86903, n86904, n86905, n86906, n86907, n86908,
    n86909, n86910, n86911, n86912, n86913, n86914, n86915, n86916, n86917,
    n86918, n86919, n86920, n86921, n86922, n86923, n86924, n86925, n86926,
    n86927, n86928, n86929, n86930, n86931, n86932, n86933, n86934, n86935,
    n86936, n86937, n86938, n86939, n86940, n86941, n86942, n86943, n86944,
    n86945, n86946, n86947, n86948, n86949, n86950, n86951, n86952, n86953,
    n86954, n86955, n86956, n86957, n86958, n86959, n86960, n86961, n86962,
    n86963, n86964, n86965, n86966, n86967, n86968, n86969, n86970, n86971,
    n86972, n86973, n86974, n86975, n86976, n86977, n86978, n86979, n86980,
    n86981, n86982, n86983, n86984, n86985, n86986, n86987, n86988, n86989,
    n86990, n86991, n86992, n86993, n86994, n86995, n86996, n86998, n86999,
    n87000, n87001, n87002, n87003, n87004, n87005, n87006, n87007, n87008,
    n87009, n87010, n87011, n87012, n87013, n87014, n87015, n87016, n87017,
    n87018, n87019, n87020, n87021, n87022, n87023, n87024, n87025, n87026,
    n87027, n87028, n87029, n87030, n87031, n87032, n87033, n87034, n87035,
    n87036, n87038, n87039, n87040, n87041, n87042, n87043, n87044, n87045,
    n87046, n87047, n87048, n87049, n87050, n87051, n87052, n87053, n87054,
    n87055, n87056, n87057, n87058, n87059, n87060, n87061, n87062, n87063,
    n87064, n87065, n87066, n87067, n87068, n87069, n87070, n87071, n87072,
    n87073, n87074, n87075, n87076, n87077, n87078, n87079, n87080, n87081,
    n87082, n87083, n87084, n87085, n87086, n87087, n87088, n87089, n87090,
    n87091, n87092, n87093, n87094, n87095, n87096, n87097, n87098, n87099,
    n87100, n87101, n87102, n87103, n87104, n87105, n87106, n87107, n87108,
    n87109, n87110, n87111, n87112, n87113, n87114, n87115, n87116, n87117,
    n87118, n87119, n87120, n87121, n87122, n87123, n87124, n87125, n87126,
    n87127, n87128, n87129, n87130, n87131, n87132, n87133, n87134, n87135,
    n87136, n87137, n87138, n87139, n87140, n87141, n87142, n87144, n87145,
    n87146, n87147, n87148, n87149, n87150, n87151, n87152, n87153, n87154,
    n87155, n87156, n87157, n87158, n87159, n87160, n87161, n87162, n87163,
    n87164, n87165, n87166, n87167, n87168, n87169, n87170, n87171, n87172,
    n87173, n87174, n87175, n87176, n87177, n87178, n87179, n87180, n87181,
    n87182, n87183, n87184, n87185, n87186, n87187, n87189, n87190, n87191,
    n87192, n87193, n87194, n87195, n87196, n87197, n87198, n87199, n87200,
    n87201, n87202, n87203, n87204, n87205, n87206, n87207, n87208, n87209,
    n87210, n87211, n87212, n87213, n87214, n87215, n87216, n87217, n87218,
    n87219, n87220, n87221, n87222, n87223, n87224, n87225, n87226, n87227,
    n87229, n87230, n87231, n87232, n87233, n87234, n87235, n87236, n87237,
    n87238, n87239, n87240, n87241, n87242, n87243, n87244, n87245, n87246,
    n87247, n87248, n87249, n87250, n87251, n87252, n87253, n87254, n87255,
    n87256, n87257, n87258, n87259, n87260, n87261, n87262, n87263, n87264,
    n87265, n87266, n87267, n87268, n87269, n87270, n87271, n87272, n87273,
    n87274, n87275, n87276, n87277, n87278, n87279, n87280, n87281, n87282,
    n87283, n87284, n87285, n87286, n87287, n87288, n87289, n87290, n87291,
    n87292, n87293, n87294, n87295, n87296, n87297, n87298, n87299, n87300,
    n87301, n87302, n87303, n87304, n87305, n87306, n87307, n87308, n87309,
    n87310, n87311, n87312, n87313, n87314, n87315, n87316, n87317, n87319,
    n87320, n87321, n87322, n87323, n87324, n87325, n87326, n87327, n87328,
    n87329, n87330, n87331, n87332, n87333, n87334, n87335, n87336, n87337,
    n87338, n87339, n87340, n87341, n87342, n87343, n87344, n87345, n87346,
    n87347, n87348, n87349, n87350, n87351, n87352, n87353, n87354, n87355,
    n87356, n87357, n87358, n87360, n87361, n87362, n87363, n87364, n87365,
    n87366, n87367, n87368, n87369, n87370, n87371, n87372, n87373, n87374,
    n87375, n87376, n87377, n87378, n87379, n87380, n87381, n87382, n87383,
    n87384, n87385, n87386, n87387, n87388, n87389, n87390, n87391, n87392,
    n87393, n87394, n87395, n87396, n87397, n87398, n87399, n87400, n87401,
    n87402, n87403, n87404, n87405, n87406, n87407, n87408, n87409, n87410,
    n87411, n87412, n87413, n87414, n87415, n87416, n87417, n87418, n87419,
    n87420, n87421, n87422, n87423, n87424, n87425, n87426, n87427, n87428,
    n87429, n87430, n87431, n87432, n87433, n87434, n87435, n87436, n87437,
    n87438, n87439, n87440, n87441, n87442, n87443, n87444, n87445, n87446,
    n87447, n87448, n87449, n87451, n87452, n87453, n87454, n87455, n87456,
    n87457, n87458, n87459, n87460, n87461, n87462, n87463, n87464, n87465,
    n87466, n87467, n87468, n87469, n87470, n87471, n87472, n87473, n87474,
    n87475, n87476, n87477, n87478, n87479, n87480, n87481, n87482, n87483,
    n87484, n87485, n87486, n87488, n87489, n87490, n87491, n87492, n87493,
    n87494, n87495, n87496, n87497, n87498, n87499, n87500, n87501, n87502,
    n87503, n87504, n87505, n87506, n87507, n87508, n87509, n87510, n87511,
    n87512, n87513, n87514, n87515, n87516, n87517, n87518, n87519, n87520,
    n87521, n87522, n87523, n87524, n87525, n87526, n87527, n87528, n87529,
    n87530, n87531, n87532, n87533, n87534, n87535, n87536, n87537, n87538,
    n87539, n87540, n87541, n87542, n87543, n87544, n87545, n87546, n87547,
    n87548, n87549, n87550, n87551, n87552, n87553, n87554, n87555, n87556,
    n87557, n87558, n87559, n87560, n87561, n87562, n87563, n87564, n87565,
    n87566, n87567, n87568, n87569, n87570, n87571, n87572, n87573, n87574,
    n87575, n87576, n87577, n87578, n87579, n87580, n87581, n87582, n87583,
    n87584, n87585, n87587, n87588, n87589, n87590, n87591, n87592, n87593,
    n87594, n87595, n87596, n87597, n87598, n87599, n87600, n87601, n87602,
    n87603, n87604, n87605, n87606, n87607, n87608, n87609, n87610, n87611,
    n87612, n87613, n87614, n87615, n87616, n87617, n87618, n87619, n87620,
    n87621, n87622, n87623, n87624, n87625, n87626, n87627, n87628, n87629,
    n87630, n87631, n87632, n87633, n87635, n87636, n87637, n87638, n87639,
    n87640, n87641, n87642, n87643, n87644, n87645, n87646, n87647, n87648,
    n87649, n87650, n87651, n87652, n87653, n87654, n87655, n87656, n87657,
    n87658, n87659, n87660, n87661, n87662, n87663, n87664, n87665, n87666,
    n87667, n87668, n87669, n87670, n87671, n87672, n87674, n87675, n87676,
    n87677, n87678, n87679, n87680, n87681, n87682, n87683, n87684, n87685,
    n87686, n87687, n87688, n87689, n87690, n87691, n87692, n87693, n87694,
    n87695, n87696, n87697, n87698, n87699, n87700, n87701, n87702, n87704,
    n87705, n87706, n87707, n87708, n87709, n87710, n87711, n87712, n87713,
    n87714, n87715, n87716, n87717, n87718, n87719, n87720, n87721, n87722,
    n87723, n87724, n87725, n87726, n87727, n87728, n87729, n87730, n87731,
    n87732, n87733, n87734, n87735, n87736, n87737, n87738, n87739, n87740,
    n87741, n87742, n87743, n87744, n87746, n87747, n87748, n87749, n87750,
    n87751, n87752, n87753, n87754, n87755, n87756, n87757, n87758, n87759,
    n87760, n87761, n87762, n87763, n87764, n87765, n87766, n87767, n87768,
    n87769, n87770, n87771, n87772, n87773, n87774, n87775, n87776, n87777,
    n87778, n87779, n87780, n87781, n87782, n87783, n87784, n87785, n87787,
    n87788, n87789, n87790, n87791, n87792, n87793, n87794, n87795, n87796,
    n87797, n87798, n87799, n87800, n87801, n87802, n87803, n87804, n87805,
    n87806, n87807, n87808, n87809, n87810, n87811, n87812, n87813, n87814,
    n87815, n87816, n87817, n87818, n87819, n87820, n87821, n87822, n87823,
    n87824, n87826, n87827, n87828, n87829, n87830, n87831, n87832, n87833,
    n87834, n87835, n87836, n87837, n87838, n87839, n87840, n87841, n87842,
    n87843, n87844, n87845, n87846, n87847, n87848, n87849, n87850, n87851,
    n87852, n87853, n87854, n87855, n87856, n87857, n87858, n87859, n87860,
    n87861, n87862, n87863, n87864, n87865, n87866, n87867, n87868, n87869,
    n87870, n87871, n87872, n87873, n87874, n87876, n87877, n87878, n87879,
    n87880, n87881, n87882, n87883, n87884, n87885, n87886, n87887, n87888,
    n87889, n87890, n87891, n87892, n87893, n87894, n87895, n87896, n87897,
    n87898, n87899, n87900, n87901, n87902, n87903, n87904, n87905, n87906,
    n87907, n87908, n87909, n87911, n87912, n87913, n87914, n87915, n87916,
    n87917, n87918, n87919, n87920, n87921, n87922, n87923, n87924, n87925,
    n87926, n87927, n87928, n87929, n87930, n87931, n87932, n87933, n87934,
    n87935, n87936, n87937, n87938, n87939, n87940, n87941, n87942, n87943,
    n87944, n87945, n87946, n87947, n87948, n87949, n87950, n87951, n87953,
    n87954, n87955, n87956, n87957, n87958, n87959, n87960, n87961, n87962,
    n87963, n87964, n87965, n87966, n87967, n87968, n87969, n87970, n87971,
    n87972, n87973, n87974, n87975, n87976, n87977, n87978, n87979, n87980,
    n87981, n87982, n87983, n87984, n87985, n87986, n87987, n87988, n87989,
    n87990, n87992, n87993, n87994, n87995, n87996, n87997, n87998, n87999,
    n88000, n88001, n88002, n88003, n88004, n88005, n88006, n88007, n88008,
    n88009, n88010, n88011, n88012, n88013, n88014, n88015, n88016, n88017,
    n88018, n88019, n88020, n88021, n88022, n88023, n88024, n88025, n88026,
    n88027, n88028, n88029, n88030, n88031, n88032, n88033, n88034, n88035,
    n88036, n88037, n88039, n88040, n88041, n88042, n88043, n88044, n88045,
    n88046, n88047, n88048, n88049, n88050, n88051, n88052, n88053, n88054,
    n88055, n88056, n88057, n88058, n88059, n88060, n88061, n88062, n88063,
    n88064, n88065, n88066, n88067, n88068, n88069, n88070, n88071, n88072,
    n88073, n88074, n88075, n88076, n88077, n88078, n88079, n88080, n88081,
    n88082, n88083, n88084, n88085, n88086, n88087, n88088, n88089, n88090,
    n88091, n88092, n88093, n88094, n88095, n88096, n88097, n88098, n88099,
    n88100, n88101, n88102, n88103, n88104, n88105, n88106, n88107, n88108,
    n88109, n88110, n88111, n88112, n88113, n88114, n88115, n88116, n88117,
    n88118, n88119, n88120, n88121, n88122, n88123, n88124, n88125, n88126,
    n88127, n88128, n88129, n88130, n88131, n88132, n88133, n88134, n88135,
    n88137, n88138, n88139, n88140, n88141, n88142, n88143, n88144, n88145,
    n88146, n88147, n88148, n88149, n88150, n88151, n88152, n88153, n88154,
    n88155, n88156, n88157, n88158, n88159, n88160, n88161, n88162, n88163,
    n88164, n88165, n88166, n88167, n88168, n88169, n88170, n88171, n88173,
    n88174, n88175, n88176, n88177, n88178, n88179, n88180, n88181, n88182,
    n88183, n88184, n88185, n88186, n88187, n88188, n88189, n88190, n88191,
    n88192, n88193, n88194, n88195, n88196, n88197, n88198, n88199, n88200,
    n88201, n88202, n88203, n88204, n88206, n88207, n88208, n88209, n88210,
    n88211, n88212, n88213, n88214, n88215, n88216, n88217, n88218, n88219,
    n88220, n88221, n88222, n88223, n88224, n88225, n88226, n88227, n88228,
    n88229, n88230, n88231, n88233, n88234, n88235, n88236, n88237, n88238,
    n88239, n88240, n88241, n88242, n88243, n88244, n88245, n88246, n88247,
    n88248, n88249, n88250, n88251, n88252, n88253, n88254, n88255, n88256,
    n88257, n88258, n88259, n88260, n88261, n88262, n88263, n88264, n88265,
    n88266, n88267, n88268, n88269, n88270, n88271, n88272, n88273, n88274,
    n88275, n88276, n88278, n88279, n88280, n88281, n88282, n88283, n88284,
    n88285, n88286, n88287, n88288, n88289, n88290, n88291, n88292, n88293,
    n88294, n88295, n88296, n88297, n88298, n88299, n88300, n88301, n88302,
    n88303, n88304, n88305, n88306, n88307, n88308, n88309, n88310, n88311,
    n88312, n88314, n88315, n88316, n88317, n88318, n88319, n88320, n88321,
    n88322, n88323, n88324, n88325, n88326, n88327, n88328, n88329, n88330,
    n88331, n88332, n88333, n88334, n88335, n88336, n88337, n88338, n88339,
    n88340, n88341, n88342, n88343, n88344, n88345, n88347, n88348, n88349,
    n88350, n88351, n88352, n88353, n88354, n88355, n88356, n88357, n88358,
    n88359, n88360, n88361, n88362, n88363, n88364, n88365, n88366, n88367,
    n88368, n88369, n88370, n88371, n88372, n88373, n88374, n88375, n88377,
    n88378, n88379, n88380, n88381, n88382, n88383, n88384, n88385, n88386,
    n88387, n88388, n88389, n88390, n88391, n88392, n88393, n88394, n88395,
    n88396, n88397, n88398, n88399, n88400, n88401, n88402, n88403, n88404,
    n88405, n88406, n88407, n88408, n88409, n88410, n88411, n88412, n88413,
    n88414, n88415, n88416, n88417, n88418, n88419, n88420, n88421, n88422,
    n88423, n88424, n88425, n88426, n88427, n88428, n88429, n88430, n88431,
    n88432, n88433, n88434, n88435, n88436, n88437, n88438, n88439, n88440,
    n88441, n88442, n88443, n88444, n88445, n88446, n88447, n88448, n88449,
    n88450, n88451, n88452, n88453, n88454, n88455, n88456, n88457, n88458,
    n88459, n88460, n88461, n88462, n88463, n88464, n88465, n88466, n88467,
    n88468, n88469, n88470, n88471, n88472, n88473, n88474, n88476, n88477,
    n88478, n88479, n88480, n88481, n88482, n88483, n88484, n88485, n88486,
    n88487, n88488, n88489, n88490, n88491, n88492, n88493, n88494, n88495,
    n88496, n88497, n88498, n88499, n88500, n88501, n88502, n88503, n88504,
    n88505, n88506, n88507, n88508, n88509, n88510, n88511, n88512, n88513,
    n88514, n88515, n88516, n88517, n88518, n88519, n88520, n88522, n88523,
    n88524, n88525, n88526, n88527, n88528, n88529, n88530, n88531, n88532,
    n88533, n88534, n88535, n88536, n88537, n88538, n88539, n88540, n88541,
    n88542, n88543, n88544, n88545, n88546, n88547, n88548, n88549, n88550,
    n88551, n88552, n88553, n88554, n88555, n88556, n88557, n88558, n88559,
    n88560, n88561, n88562, n88563, n88564, n88565, n88566, n88567, n88568,
    n88569, n88570, n88571, n88572, n88573, n88574, n88575, n88576, n88577,
    n88578, n88579, n88580, n88581, n88582, n88583, n88584, n88585, n88586,
    n88587, n88588, n88589, n88590, n88591, n88592, n88593, n88594, n88595,
    n88596, n88597, n88598, n88599, n88600, n88601, n88602, n88603, n88604,
    n88605, n88606, n88607, n88608, n88609, n88610, n88611, n88612, n88613,
    n88614, n88615, n88616, n88617, n88618, n88619, n88620, n88621, n88623,
    n88624, n88625, n88626, n88627, n88628, n88629, n88630, n88631, n88632,
    n88633, n88634, n88635, n88636, n88637, n88638, n88639, n88640, n88641,
    n88642, n88643, n88644, n88645, n88646, n88647, n88648, n88649, n88650,
    n88651, n88652, n88653, n88655, n88656, n88657, n88658, n88659, n88660,
    n88661, n88662, n88663, n88664, n88665, n88666, n88667, n88668, n88669,
    n88670, n88671, n88672, n88673, n88674, n88675, n88676, n88677, n88678,
    n88679, n88680, n88681, n88682, n88683, n88684, n88685, n88686, n88687,
    n88688, n88689, n88691, n88692, n88693, n88694, n88695, n88696, n88697,
    n88698, n88699, n88700, n88701, n88702, n88703, n88704, n88705, n88706,
    n88707, n88708, n88709, n88710, n88711, n88712, n88713, n88714, n88715,
    n88716, n88717, n88718, n88719, n88720, n88721, n88722, n88723, n88724,
    n88725, n88726, n88727, n88728, n88729, n88730, n88731, n88732, n88733,
    n88734, n88735, n88736, n88737, n88738, n88739, n88740, n88741, n88742,
    n88743, n88744, n88745, n88746, n88747, n88748, n88749, n88750, n88751,
    n88752, n88753, n88754, n88755, n88756, n88757, n88758, n88759, n88760,
    n88761, n88762, n88763, n88764, n88765, n88766, n88767, n88768, n88769,
    n88770, n88771, n88772, n88773, n88774, n88775, n88776, n88777, n88778,
    n88779, n88780, n88781, n88782, n88783, n88784, n88785, n88786, n88787,
    n88788, n88790, n88791, n88792, n88793, n88794, n88795, n88796, n88797,
    n88798, n88799, n88800, n88801, n88802, n88803, n88804, n88805, n88806,
    n88807, n88808, n88809, n88810, n88811, n88812, n88813, n88814, n88815,
    n88816, n88817, n88818, n88819, n88820, n88821, n88822, n88823, n88824,
    n88825, n88826, n88827, n88828, n88829, n88830, n88831, n88832, n88833,
    n88834, n88835, n88836, n88837, n88838, n88839, n88840, n88841, n88842,
    n88843, n88844, n88845, n88846, n88847, n88848, n88849, n88850, n88851,
    n88852, n88853, n88854, n88855, n88856, n88857, n88858, n88859, n88860,
    n88861, n88862, n88863, n88864, n88865, n88866, n88867, n88868, n88869,
    n88870, n88871, n88872, n88873, n88874, n88875, n88876, n88877, n88878,
    n88879, n88880, n88881, n88882, n88883, n88884, n88885, n88886, n88887,
    n88888, n88889, n88890, n88892, n88893, n88894, n88895, n88896, n88897,
    n88898, n88899, n88900, n88901, n88902, n88903, n88904, n88905, n88906,
    n88907, n88908, n88909, n88910, n88911, n88912, n88913, n88914, n88915,
    n88916, n88917, n88918, n88919, n88920, n88921, n88922, n88923, n88925,
    n88926, n88927, n88928, n88929, n88930, n88931, n88932, n88933, n88934,
    n88935, n88936, n88937, n88938, n88939, n88940, n88941, n88942, n88943,
    n88944, n88945, n88946, n88947, n88948, n88949, n88950, n88951, n88952,
    n88953, n88954, n88955, n88956, n88957, n88958, n88959, n88960, n88961,
    n88962, n88963, n88964, n88965, n88966, n88967, n88968, n88969, n88970,
    n88971, n88972, n88973, n88974, n88975, n88976, n88977, n88978, n88979,
    n88980, n88981, n88982, n88983, n88984, n88985, n88986, n88987, n88988,
    n88989, n88990, n88991, n88992, n88993, n88994, n88995, n88996, n88997,
    n88998, n88999, n89000, n89001, n89002, n89003, n89004, n89005, n89006,
    n89007, n89008, n89009, n89010, n89011, n89012, n89013, n89014, n89015,
    n89016, n89017, n89018, n89019, n89020, n89021, n89022, n89023, n89024,
    n89025, n89026, n89027, n89029, n89030, n89031, n89032, n89033, n89034,
    n89035, n89036, n89037, n89038, n89039, n89040, n89041, n89042, n89043,
    n89044, n89045, n89046, n89047, n89048, n89049, n89050, n89051, n89052,
    n89053, n89054, n89055, n89056, n89057, n89058, n89059, n89060, n89061,
    n89062, n89063, n89064, n89065, n89066, n89068, n89069, n89070, n89071,
    n89072, n89073, n89074, n89075, n89076, n89077, n89078, n89079, n89080,
    n89081, n89082, n89083, n89084, n89085, n89086, n89087, n89088, n89089,
    n89090, n89091, n89092, n89093, n89094, n89095, n89096, n89097, n89098,
    n89099, n89100, n89101, n89102, n89103, n89104, n89105, n89106, n89107,
    n89108, n89109, n89110, n89111, n89112, n89113, n89114, n89115, n89116,
    n89117, n89118, n89119, n89120, n89121, n89122, n89123, n89124, n89125,
    n89126, n89127, n89128, n89129, n89130, n89131, n89132, n89133, n89134,
    n89135, n89136, n89137, n89138, n89139, n89140, n89141, n89142, n89143,
    n89144, n89145, n89146, n89147, n89148, n89149, n89150, n89151, n89152,
    n89153, n89154, n89155, n89156, n89157, n89158, n89159, n89160, n89161,
    n89162, n89163, n89164, n89165, n89167, n89168, n89169, n89170, n89171,
    n89172, n89173, n89174, n89175, n89176, n89177, n89178, n89179, n89180,
    n89181, n89182, n89183, n89184, n89185, n89186, n89187, n89188, n89189,
    n89190, n89191, n89192, n89193, n89194, n89195, n89196, n89197, n89198,
    n89199, n89200, n89201, n89202, n89203, n89204, n89205, n89206, n89207,
    n89208, n89209, n89210, n89211, n89212, n89214, n89215, n89216, n89217,
    n89218, n89219, n89220, n89221, n89222, n89223, n89224, n89225, n89226,
    n89227, n89228, n89229, n89230, n89231, n89232, n89233, n89234, n89235,
    n89236, n89237, n89238, n89239, n89240, n89241, n89242, n89243, n89244,
    n89245, n89246, n89247, n89248, n89249, n89250, n89251, n89252, n89253,
    n89254, n89255, n89256, n89257, n89258, n89259, n89260, n89261, n89262,
    n89263, n89264, n89265, n89266, n89267, n89268, n89269, n89270, n89271,
    n89272, n89273, n89274, n89275, n89276, n89277, n89278, n89279, n89280,
    n89281, n89282, n89283, n89284, n89285, n89286, n89287, n89288, n89289,
    n89290, n89291, n89292, n89293, n89294, n89295, n89296, n89297, n89298,
    n89299, n89300, n89301, n89302, n89303, n89304, n89306, n89307, n89308,
    n89309, n89310, n89311, n89312, n89313, n89314, n89315, n89316, n89317,
    n89318, n89319, n89320, n89321, n89322, n89323, n89324, n89325, n89326,
    n89327, n89328, n89329, n89330, n89331, n89332, n89333, n89334, n89335,
    n89336, n89337, n89338, n89339, n89340, n89341, n89342, n89343, n89344,
    n89345, n89346, n89347, n89348, n89349, n89350, n89351, n89352, n89354,
    n89355, n89356, n89357, n89358, n89359, n89360, n89361, n89362, n89363,
    n89364, n89365, n89366, n89367, n89368, n89369, n89370, n89371, n89372,
    n89373, n89374, n89375, n89376, n89377, n89378, n89379, n89380, n89381,
    n89382, n89383, n89384, n89385, n89386, n89387, n89388, n89389, n89390,
    n89391, n89392, n89393, n89394, n89395, n89396, n89397, n89398, n89399,
    n89400, n89401, n89402, n89403, n89404, n89405, n89406, n89407, n89408,
    n89409, n89410, n89411, n89412, n89413, n89414, n89415, n89416, n89417,
    n89418, n89419, n89420, n89421, n89422, n89423, n89424, n89425, n89426,
    n89427, n89428, n89429, n89430, n89431, n89432, n89433, n89434, n89435,
    n89436, n89437, n89438, n89439, n89440, n89441, n89442, n89444, n89445,
    n89446, n89447, n89448, n89449, n89450, n89451, n89452, n89453, n89454,
    n89455, n89456, n89457, n89458, n89459, n89460, n89461, n89462, n89463,
    n89464, n89465, n89466, n89467, n89468, n89469, n89470, n89471, n89472,
    n89473, n89474, n89475, n89476, n89477, n89478, n89479, n89480, n89481,
    n89482, n89483, n89484, n89485, n89486, n89487, n89488, n89489, n89490,
    n89491, n89492, n89493, n89494, n89495, n89496, n89497, n89499, n89500,
    n89501, n89502, n89503, n89504, n89505, n89506, n89507, n89508, n89509,
    n89510, n89511, n89512, n89513, n89514, n89515, n89516, n89517, n89518,
    n89519, n89520, n89521, n89522, n89523, n89524, n89525, n89526, n89527,
    n89528, n89529, n89530, n89531, n89532, n89533, n89534, n89535, n89537,
    n89538, n89539, n89540, n89541, n89542, n89543, n89544, n89545, n89546,
    n89547, n89548, n89549, n89550, n89551, n89552, n89553, n89554, n89555,
    n89556, n89557, n89558, n89559, n89560, n89561, n89562, n89563, n89564,
    n89565, n89566, n89567, n89568, n89569, n89570, n89571, n89572, n89573,
    n89574, n89575, n89577, n89578, n89579, n89580, n89581, n89582, n89583,
    n89584, n89585, n89586, n89587, n89588, n89589, n89590, n89591, n89592,
    n89593, n89594, n89595, n89596, n89597, n89598, n89599, n89600, n89601,
    n89602, n89603, n89604, n89605, n89607, n89608, n89609, n89610, n89611,
    n89612, n89613, n89614, n89615, n89616, n89617, n89618, n89619, n89620,
    n89621, n89622, n89623, n89624, n89625, n89626, n89627, n89628, n89629,
    n89630, n89631, n89632, n89633, n89634, n89635, n89636, n89637, n89638,
    n89639, n89641, n89642, n89643, n89644, n89645, n89646, n89647, n89648,
    n89649, n89650, n89651, n89652, n89653, n89654, n89655, n89656, n89657,
    n89658, n89659, n89660, n89661, n89662, n89663, n89664, n89665, n89666,
    n89667, n89668, n89669, n89670, n89671, n89672, n89673, n89674, n89675,
    n89676, n89677, n89679, n89680, n89681, n89682, n89683, n89684, n89685,
    n89686, n89687, n89688, n89689, n89690, n89691, n89692, n89693, n89694,
    n89695, n89696, n89697, n89698, n89699, n89700, n89701, n89702, n89703,
    n89704, n89705, n89706, n89707, n89708, n89709, n89710, n89711, n89712,
    n89713, n89714, n89715, n89716, n89717, n89718, n89719, n89720, n89722,
    n89723, n89724, n89725, n89726, n89727, n89728, n89729, n89730, n89731,
    n89732, n89733, n89734, n89735, n89736, n89737, n89738, n89739, n89740,
    n89741, n89742, n89743, n89744, n89745, n89746, n89747, n89748, n89749,
    n89750, n89751, n89752, n89753, n89754, n89755, n89756, n89757, n89758,
    n89759, n89760, n89761, n89762, n89763, n89764, n89765, n89766, n89767,
    n89769, n89770, n89771, n89772, n89773, n89774, n89775, n89776, n89777,
    n89778, n89779, n89780, n89781, n89782, n89783, n89784, n89785, n89786,
    n89787, n89788, n89789, n89790, n89791, n89792, n89793, n89794, n89795,
    n89796, n89797, n89798, n89799, n89800, n89801, n89802, n89803, n89804,
    n89805, n89806, n89807, n89808, n89809, n89810, n89811, n89812, n89813,
    n89814, n89815, n89816, n89817, n89818, n89819, n89821, n89822, n89823,
    n89824, n89825, n89826, n89827, n89828, n89829, n89830, n89831, n89832,
    n89833, n89834, n89835, n89836, n89837, n89838, n89839, n89840, n89841,
    n89842, n89843, n89844, n89845, n89846, n89847, n89848, n89849, n89850,
    n89851, n89852, n89853, n89854, n89856, n89857, n89858, n89859, n89860,
    n89861, n89862, n89863, n89864, n89865, n89866, n89867, n89868, n89869,
    n89870, n89871, n89872, n89873, n89874, n89875, n89876, n89877, n89878,
    n89879, n89880, n89881, n89882, n89883, n89884, n89885, n89886, n89887,
    n89888, n89889, n89890, n89892, n89893, n89894, n89895, n89896, n89897,
    n89898, n89899, n89900, n89901, n89902, n89903, n89904, n89905, n89906,
    n89907, n89908, n89909, n89910, n89911, n89912, n89913, n89914, n89915,
    n89916, n89917, n89918, n89919, n89920, n89922, n89923, n89924, n89925,
    n89926, n89927, n89928, n89929, n89930, n89931, n89932, n89933, n89934,
    n89935, n89936, n89937, n89938, n89939, n89940, n89941, n89942, n89943,
    n89944, n89945, n89946, n89947, n89948, n89949, n89950, n89951, n89952,
    n89953, n89954, n89955, n89956, n89957, n89958, n89960, n89961, n89962,
    n89963, n89964, n89965, n89966, n89967, n89968, n89969, n89970, n89971,
    n89972, n89973, n89974, n89975, n89976, n89977, n89978, n89979, n89980,
    n89981, n89982, n89983, n89984, n89985, n89986, n89987, n89988, n89989,
    n89990, n89991, n89992, n89993, n89995, n89996, n89997, n89998, n89999,
    n90000, n90001, n90002, n90003, n90004, n90005, n90006, n90007, n90008,
    n90009, n90010, n90011, n90012, n90013, n90014, n90015, n90016, n90017,
    n90018, n90019, n90020, n90021, n90022, n90023, n90024, n90025, n90026,
    n90027, n90028, n90029, n90030, n90031, n90033, n90034, n90035, n90036,
    n90037, n90038, n90039, n90040, n90041, n90042, n90043, n90044, n90045,
    n90046, n90047, n90048, n90049, n90050, n90051, n90052, n90053, n90054,
    n90055, n90056, n90057, n90058, n90059, n90060, n90061, n90062, n90063,
    n90064, n90065, n90067, n90068, n90069, n90070, n90071, n90072, n90073,
    n90074, n90075, n90076, n90077, n90078, n90079, n90080, n90081, n90082,
    n90083, n90084, n90085, n90086, n90087, n90088, n90089, n90090, n90091,
    n90093, n90094, n90095, n90096, n90097, n90098, n90099, n90100, n90101,
    n90102, n90103, n90104, n90105, n90106, n90107, n90108, n90109, n90110,
    n90111, n90112, n90113, n90114, n90115, n90116, n90117, n90118, n90119,
    n90120, n90121, n90122, n90123, n90124, n90125, n90126, n90127, n90128,
    n90129, n90130, n90131, n90132, n90133, n90134, n90135, n90136, n90137,
    n90138, n90139, n90140, n90141, n90142, n90143, n90144, n90145, n90146,
    n90147, n90148, n90149, n90150, n90151, n90152, n90153, n90154, n90155,
    n90156, n90157, n90158, n90159, n90160, n90161, n90162, n90163, n90164,
    n90165, n90166, n90167, n90168, n90169, n90170, n90171, n90172, n90173,
    n90174, n90175, n90176, n90177, n90178, n90179, n90180, n90181, n90182,
    n90183, n90184, n90185, n90186, n90187, n90188, n90189, n90190, n90192,
    n90193, n90194, n90195, n90196, n90197, n90198, n90199, n90200, n90201,
    n90202, n90203, n90204, n90205, n90206, n90207, n90208, n90209, n90210,
    n90211, n90212, n90213, n90214, n90215, n90216, n90217, n90218, n90219,
    n90220, n90221, n90222, n90223, n90224, n90225, n90226, n90227, n90228,
    n90229, n90230, n90231, n90233, n90234, n90235, n90236, n90237, n90238,
    n90239, n90240, n90241, n90242, n90243, n90244, n90245, n90246, n90247,
    n90248, n90249, n90250, n90251, n90252, n90253, n90254, n90255, n90256,
    n90257, n90258, n90259, n90260, n90261, n90262, n90263, n90264, n90265,
    n90266, n90267, n90268, n90269, n90270, n90271, n90272, n90273, n90274,
    n90275, n90276, n90277, n90278, n90279, n90280, n90281, n90282, n90283,
    n90284, n90285, n90286, n90287, n90288, n90289, n90290, n90291, n90292,
    n90293, n90294, n90295, n90296, n90297, n90298, n90299, n90300, n90301,
    n90302, n90303, n90304, n90305, n90306, n90307, n90308, n90309, n90310,
    n90311, n90312, n90313, n90314, n90315, n90316, n90317, n90318, n90319,
    n90320, n90321, n90323, n90324, n90325, n90326, n90327, n90328, n90329,
    n90330, n90331, n90332, n90333, n90334, n90335, n90336, n90337, n90338,
    n90339, n90340, n90341, n90342, n90343, n90344, n90345, n90346, n90347,
    n90348, n90349, n90350, n90351, n90352, n90353, n90354, n90355, n90356,
    n90357, n90358, n90359, n90360, n90361, n90362, n90363, n90364, n90365,
    n90366, n90367, n90368, n90369, n90370, n90371, n90372, n90373, n90374,
    n90375, n90376, n90377, n90378, n90379, n90380, n90381, n90382, n90383,
    n90384, n90385, n90386, n90387, n90388, n90389, n90390, n90391, n90392,
    n90393, n90394, n90395, n90396, n90397, n90398, n90399, n90400, n90401,
    n90402, n90403, n90404, n90405, n90406, n90407, n90408, n90409, n90410,
    n90411, n90412, n90413, n90414, n90415, n90416, n90417, n90418, n90419,
    n90420, n90421, n90422, n90423, n90425, n90426, n90427, n90428, n90429,
    n90430, n90431, n90432, n90433, n90434, n90435, n90436, n90437, n90438,
    n90439, n90440, n90441, n90442, n90443, n90444, n90445, n90446, n90447,
    n90448, n90449, n90450, n90451, n90452, n90453, n90454, n90455, n90456,
    n90457, n90458, n90459, n90460, n90461, n90462, n90463, n90464, n90465,
    n90466, n90467, n90468, n90469, n90470, n90471, n90472, n90473, n90475,
    n90476, n90477, n90478, n90479, n90480, n90481, n90482, n90483, n90484,
    n90485, n90486, n90487, n90488, n90489, n90490, n90491, n90492, n90493,
    n90494, n90495, n90496, n90497, n90498, n90499, n90500, n90501, n90502,
    n90503, n90504, n90505, n90506, n90507, n90508, n90509, n90510, n90511,
    n90512, n90513, n90514, n90515, n90516, n90517, n90518, n90519, n90520,
    n90521, n90522, n90523, n90524, n90525, n90526, n90527, n90528, n90529,
    n90530, n90531, n90532, n90533, n90534, n90535, n90536, n90537, n90538,
    n90539, n90540, n90541, n90542, n90543, n90544, n90545, n90546, n90547,
    n90548, n90549, n90550, n90551, n90552, n90553, n90554, n90555, n90556,
    n90557, n90558, n90559, n90560, n90561, n90562, n90563, n90564, n90565,
    n90566, n90567, n90568, n90569, n90570, n90571, n90572, n90573, n90574,
    n90575, n90576, n90577, n90578, n90579, n90581, n90582, n90583, n90584,
    n90585, n90586, n90587, n90588, n90589, n90590, n90591, n90592, n90593,
    n90594, n90595, n90596, n90597, n90598, n90599, n90600, n90601, n90602,
    n90603, n90604, n90605, n90606, n90607, n90608, n90609, n90610, n90611,
    n90612, n90613, n90614, n90615, n90616, n90617, n90618, n90619, n90620,
    n90621, n90622, n90623, n90624, n90625, n90626, n90627, n90628, n90629,
    n90630, n90631, n90632, n90633, n90634, n90635, n90636, n90637, n90638,
    n90639, n90640, n90641, n90642, n90643, n90644, n90645, n90646, n90647,
    n90648, n90649, n90650, n90651, n90652, n90653, n90654, n90655, n90656,
    n90657, n90658, n90659, n90660, n90661, n90662, n90663, n90664, n90665,
    n90666, n90667, n90668, n90669, n90670, n90671, n90672, n90673, n90674,
    n90675, n90676, n90677, n90678, n90679, n90680, n90681, n90682, n90683,
    n90685, n90686, n90687, n90688, n90689, n90690, n90691, n90692, n90693,
    n90694, n90695, n90696, n90697, n90698, n90699, n90700, n90701, n90702,
    n90703, n90704, n90705, n90706, n90707, n90708, n90709, n90710, n90711,
    n90712, n90713, n90714, n90715, n90716, n90717, n90718, n90719, n90720,
    n90721, n90722, n90723, n90724, n90725, n90726, n90727, n90728, n90729,
    n90730, n90731, n90732, n90733, n90734, n90735, n90736, n90737, n90738,
    n90739, n90740, n90741, n90742, n90743, n90744, n90745, n90746, n90747,
    n90748, n90749, n90750, n90751, n90752, n90753, n90754, n90755, n90756,
    n90757, n90758, n90759, n90760, n90761, n90762, n90763, n90764, n90765,
    n90766, n90767, n90768, n90769, n90770, n90771, n90772, n90773, n90774,
    n90775, n90776, n90777, n90778, n90779, n90780, n90781, n90782, n90783,
    n90784, n90785, n90786, n90787, n90788, n90789, n90790, n90792, n90793,
    n90794, n90795, n90796, n90797, n90798, n90799, n90800, n90801, n90802,
    n90803, n90804, n90805, n90806, n90807, n90808, n90809, n90810, n90811,
    n90812, n90813, n90814, n90815, n90816, n90817, n90818, n90819, n90820,
    n90821, n90822, n90823, n90824, n90825, n90826, n90827, n90828, n90829,
    n90830, n90831, n90832, n90833, n90834, n90835, n90836, n90837, n90838,
    n90839, n90840, n90841, n90842, n90843, n90844, n90845, n90846, n90847,
    n90848, n90849, n90850, n90851, n90852, n90853, n90854, n90855, n90856,
    n90857, n90858, n90859, n90860, n90861, n90862, n90863, n90864, n90865,
    n90866, n90867, n90868, n90869, n90870, n90871, n90872, n90873, n90874,
    n90875, n90876, n90877, n90878, n90879, n90880, n90881, n90882, n90883,
    n90884, n90885, n90886, n90887, n90888, n90889, n90890, n90892, n90893,
    n90894, n90895, n90896, n90897, n90898, n90899, n90900, n90901, n90902,
    n90903, n90904, n90905, n90906, n90907, n90908, n90909, n90910, n90911,
    n90912, n90913, n90914, n90915, n90916, n90917, n90918, n90919, n90920,
    n90921, n90922, n90923, n90924, n90925, n90926, n90927, n90928, n90929,
    n90930, n90931, n90932, n90933, n90934, n90935, n90936, n90937, n90938,
    n90939, n90940, n90941, n90942, n90944, n90945, n90946, n90947, n90948,
    n90949, n90950, n90951, n90952, n90953, n90954, n90955, n90956, n90957,
    n90958, n90959, n90960, n90961, n90962, n90963, n90964, n90965, n90966,
    n90967, n90968, n90969, n90970, n90971, n90972, n90973, n90974, n90975,
    n90976, n90977, n90978, n90979, n90980, n90981, n90982, n90983, n90985,
    n90986, n90987, n90988, n90989, n90990, n90991, n90992, n90993, n90994,
    n90995, n90996, n90997, n90998, n90999, n91000, n91001, n91002, n91003,
    n91004, n91005, n91006, n91007, n91008, n91009, n91010, n91011, n91012,
    n91013, n91014, n91015, n91016, n91017, n91018, n91019, n91020, n91021,
    n91022, n91023, n91024, n91025, n91026, n91027, n91028, n91029, n91030,
    n91032, n91033, n91034, n91035, n91036, n91037, n91038, n91039, n91040,
    n91041, n91042, n91043, n91044, n91045, n91046, n91047, n91048, n91049,
    n91050, n91051, n91052, n91053, n91054, n91055, n91056, n91057, n91058,
    n91059, n91060, n91061, n91062, n91063, n91064, n91065, n91066, n91067,
    n91068, n91069, n91070, n91071, n91073, n91074, n91075, n91076, n91077,
    n91078, n91079, n91080, n91081, n91082, n91083, n91084, n91085, n91086,
    n91087, n91088, n91089, n91090, n91091, n91092, n91093, n91094, n91095,
    n91096, n91097, n91098, n91099, n91100, n91101, n91102, n91103, n91104,
    n91105, n91106, n91107, n91108, n91109, n91110, n91111, n91112, n91113,
    n91114, n91116, n91117, n91118, n91119, n91120, n91121, n91122, n91123,
    n91124, n91125, n91126, n91127, n91128, n91129, n91130, n91131, n91132,
    n91133, n91134, n91135, n91136, n91137, n91138, n91139, n91140, n91141,
    n91142, n91143, n91144, n91146, n91147, n91148, n91149, n91150, n91151,
    n91152, n91153, n91154, n91155, n91156, n91157, n91158, n91159, n91160,
    n91161, n91162, n91163, n91164, n91165, n91166, n91167, n91168, n91169,
    n91170, n91171, n91172, n91173, n91174, n91175, n91176, n91177, n91178,
    n91179, n91180, n91181, n91183, n91184, n91185, n91186, n91187, n91188,
    n91189, n91190, n91191, n91192, n91193, n91194, n91195, n91196, n91197,
    n91198, n91199, n91200, n91201, n91202, n91203, n91204, n91205, n91206,
    n91207, n91208, n91209, n91210, n91211, n91212, n91213, n91215, n91216,
    n91217, n91218, n91219, n91220, n91221, n91222, n91223, n91224, n91225,
    n91226, n91227, n91228, n91229, n91230, n91231, n91232, n91233, n91234,
    n91235, n91236, n91237, n91238, n91239, n91240, n91241, n91242, n91243,
    n91244, n91246, n91247, n91248, n91249, n91250, n91251, n91252, n91253,
    n91254, n91255, n91256, n91257, n91258, n91259, n91260, n91261, n91262,
    n91263, n91264, n91265, n91266, n91267, n91268, n91269, n91270, n91271,
    n91272, n91273, n91274, n91275, n91276, n91278, n91279, n91280, n91281,
    n91282, n91283, n91284, n91285, n91286, n91287, n91288, n91289, n91290,
    n91291, n91292, n91293, n91294, n91295, n91296, n91297, n91298, n91299,
    n91300, n91301, n91302, n91303, n91304, n91305, n91306, n91307, n91308,
    n91309, n91310, n91311, n91312, n91313, n91315, n91316, n91317, n91318,
    n91319, n91320, n91321, n91322, n91323, n91324, n91325, n91326, n91327,
    n91328, n91329, n91330, n91331, n91332, n91333, n91334, n91335, n91336,
    n91337, n91338, n91339, n91340, n91341, n91342, n91343, n91344, n91345,
    n91346, n91347, n91348, n91349, n91350, n91351, n91353, n91354, n91355,
    n91356, n91357, n91358, n91359, n91360, n91361, n91362, n91363, n91364,
    n91365, n91366, n91367, n91368, n91369, n91370, n91371, n91372, n91373,
    n91374, n91375, n91376, n91377, n91378, n91379, n91380, n91381, n91383,
    n91384, n91385, n91386, n91387, n91388, n91389, n91390, n91391, n91392,
    n91393, n91394, n91395, n91396, n91397, n91398, n91399, n91400, n91401,
    n91402, n91403, n91404, n91405, n91406, n91407, n91408, n91409, n91410,
    n91411, n91412, n91413, n91414, n91415, n91416, n91417, n91418, n91419,
    n91420, n91421, n91422, n91423, n91424, n91425, n91426, n91427, n91428,
    n91429, n91430, n91431, n91432, n91433, n91434, n91435, n91436, n91437,
    n91438, n91439, n91440, n91441, n91442, n91443, n91444, n91445, n91446,
    n91447, n91448, n91449, n91450, n91451, n91452, n91453, n91454, n91455,
    n91456, n91457, n91458, n91459, n91460, n91461, n91462, n91463, n91464,
    n91465, n91466, n91467, n91468, n91469, n91470, n91471, n91472, n91473,
    n91474, n91475, n91476, n91477, n91478, n91479, n91481, n91482, n91483,
    n91484, n91485, n91486, n91487, n91488, n91489, n91490, n91491, n91492,
    n91493, n91494, n91495, n91496, n91497, n91498, n91499, n91500, n91501,
    n91502, n91503, n91504, n91505, n91506, n91507, n91508, n91509, n91510,
    n91511, n91512, n91513, n91514, n91515, n91516, n91517, n91518, n91519,
    n91521, n91522, n91523, n91524, n91525, n91526, n91527, n91528, n91529,
    n91530, n91531, n91532, n91533, n91534, n91535, n91536, n91537, n91538,
    n91539, n91540, n91541, n91542, n91543, n91544, n91545, n91546, n91547,
    n91548, n91549, n91550, n91551, n91552, n91553, n91554, n91555, n91556,
    n91557, n91558, n91559, n91560, n91561, n91562, n91563, n91564, n91565,
    n91567, n91568, n91569, n91570, n91571, n91572, n91573, n91574, n91575,
    n91576, n91577, n91578, n91579, n91580, n91581, n91582, n91583, n91584,
    n91585, n91586, n91587, n91588, n91589, n91590, n91591, n91592, n91593,
    n91594, n91595, n91596, n91597, n91598, n91599, n91600, n91601, n91602,
    n91603, n91604, n91605, n91606, n91608, n91609, n91610, n91611, n91612,
    n91613, n91614, n91615, n91616, n91617, n91618, n91619, n91620, n91621,
    n91622, n91623, n91624, n91625, n91626, n91627, n91628, n91629, n91630,
    n91631, n91632, n91634, n91635, n91636, n91637, n91638, n91639, n91640,
    n91641, n91642, n91643, n91644, n91645, n91646, n91647, n91648, n91649,
    n91650, n91651, n91652, n91653, n91654, n91655, n91656, n91657, n91658,
    n91659, n91660, n91661, n91662, n91663, n91664, n91665, n91666, n91668,
    n91669, n91670, n91671, n91672, n91673, n91674, n91675, n91676, n91677,
    n91678, n91679, n91680, n91681, n91682, n91683, n91684, n91685, n91686,
    n91687, n91688, n91689, n91690, n91691, n91692, n91693, n91694, n91695,
    n91696, n91697, n91698, n91699, n91700, n91701, n91702, n91703, n91704,
    n91705, n91706, n91707, n91708, n91709, n91710, n91711, n91713, n91714,
    n91715, n91716, n91717, n91718, n91719, n91720, n91721, n91722, n91723,
    n91724, n91725, n91726, n91727, n91728, n91729, n91730, n91731, n91732,
    n91733, n91734, n91735, n91736, n91737, n91738, n91739, n91740, n91741,
    n91742, n91743, n91744, n91745, n91746, n91747, n91749, n91750, n91751,
    n91752, n91753, n91754, n91755, n91756, n91757, n91758, n91759, n91760,
    n91761, n91762, n91763, n91764, n91765, n91766, n91767, n91768, n91769,
    n91770, n91771, n91772, n91773, n91774, n91775, n91776, n91777, n91778,
    n91779, n91780, n91781, n91782, n91783, n91784, n91786, n91787, n91788,
    n91789, n91790, n91791, n91792, n91793, n91794, n91795, n91796, n91797,
    n91798, n91799, n91800, n91801, n91802, n91803, n91804, n91805, n91806,
    n91807, n91808, n91809, n91810, n91811, n91812, n91813, n91814, n91815,
    n91816, n91817, n91819, n91820, n91821, n91822, n91823, n91824, n91825,
    n91826, n91827, n91828, n91829, n91830, n91831, n91832, n91833, n91834,
    n91835, n91836, n91837, n91838, n91839, n91840, n91841, n91842, n91843,
    n91844, n91845, n91846, n91847, n91848, n91849, n91850, n91851, n91852,
    n91853, n91854, n91855, n91856, n91857, n91858, n91859, n91860, n91861,
    n91862, n91863, n91864, n91865, n91866, n91867, n91868, n91869, n91870,
    n91871, n91872, n91873, n91874, n91875, n91876, n91877, n91878, n91879,
    n91880, n91881, n91882, n91883, n91884, n91885, n91886, n91887, n91888,
    n91889, n91890, n91891, n91892, n91893, n91894, n91895, n91896, n91897,
    n91898, n91899, n91900, n91901, n91902, n91903, n91904, n91905, n91906,
    n91907, n91908, n91909, n91910, n91911, n91912, n91913, n91914, n91915,
    n91916, n91917, n91918, n91919, n91921, n91922, n91923, n91924, n91925,
    n91926, n91927, n91928, n91929, n91930, n91931, n91932, n91933, n91934,
    n91935, n91936, n91937, n91938, n91939, n91940, n91941, n91942, n91943,
    n91944, n91945, n91946, n91947, n91948, n91949, n91950, n91951, n91952,
    n91953, n91954, n91955, n91956, n91957, n91958, n91959, n91960, n91961,
    n91962, n91963, n91964, n91965, n91966, n91967, n91968, n91969, n91970,
    n91971, n91972, n91973, n91974, n91975, n91976, n91977, n91978, n91979,
    n91980, n91981, n91982, n91983, n91984, n91985, n91986, n91987, n91988,
    n91989, n91990, n91991, n91992, n91993, n91994, n91995, n91996, n91997,
    n91998, n91999, n92000, n92001, n92002, n92003, n92004, n92005, n92006,
    n92007, n92008, n92009, n92010, n92011, n92012, n92013, n92014, n92015,
    n92016, n92017, n92018, n92019, n92020, n92022, n92023, n92024, n92025,
    n92026, n92027, n92028, n92029, n92030, n92031, n92032, n92033, n92034,
    n92035, n92036, n92037, n92038, n92039, n92040, n92041, n92042, n92043,
    n92044, n92045, n92046, n92047, n92048, n92049, n92050, n92051, n92052,
    n92053, n92054, n92055, n92056, n92057, n92058, n92059, n92060, n92061,
    n92062, n92063, n92064, n92065, n92066, n92067, n92068, n92069, n92070,
    n92071, n92072, n92073, n92074, n92075, n92076, n92077, n92078, n92079,
    n92080, n92081, n92082, n92083, n92084, n92085, n92086, n92087, n92088,
    n92089, n92090, n92091, n92092, n92093, n92094, n92095, n92096, n92097,
    n92098, n92099, n92100, n92101, n92102, n92103, n92104, n92105, n92106,
    n92107, n92108, n92109, n92110, n92111, n92112, n92113, n92114, n92115,
    n92116, n92117, n92118, n92119, n92120, n92121, n92122, n92123, n92124,
    n92126, n92127, n92128, n92129, n92130, n92131, n92132, n92133, n92134,
    n92135, n92136, n92137, n92138, n92139, n92140, n92141, n92142, n92143,
    n92144, n92145, n92146, n92147, n92148, n92149, n92150, n92151, n92152,
    n92153, n92154, n92155, n92156, n92157, n92158, n92159, n92160, n92161,
    n92162, n92163, n92164, n92165, n92166, n92167, n92169, n92170, n92171,
    n92172, n92173, n92174, n92175, n92176, n92177, n92178, n92179, n92180,
    n92181, n92182, n92183, n92184, n92185, n92186, n92187, n92188, n92189,
    n92190, n92191, n92192, n92193, n92194, n92195, n92196, n92197, n92198,
    n92199, n92200, n92201, n92202, n92203, n92204, n92205, n92206, n92207,
    n92208, n92209, n92210, n92211, n92212, n92213, n92214, n92215, n92216,
    n92217, n92218, n92219, n92220, n92221, n92222, n92223, n92224, n92225,
    n92226, n92227, n92228, n92229, n92230, n92231, n92232, n92233, n92234,
    n92235, n92236, n92237, n92238, n92239, n92240, n92241, n92242, n92243,
    n92244, n92245, n92246, n92247, n92248, n92249, n92250, n92251, n92252,
    n92253, n92254, n92255, n92256, n92257, n92258, n92259, n92260, n92261,
    n92262, n92263, n92264, n92265, n92266, n92267, n92268, n92270, n92271,
    n92272, n92273, n92274, n92275, n92276, n92277, n92278, n92279, n92280,
    n92281, n92282, n92283, n92284, n92285, n92286, n92287, n92288, n92289,
    n92290, n92291, n92292, n92293, n92294, n92295, n92296, n92297, n92298,
    n92300, n92301, n92302, n92303, n92304, n92305, n92306, n92307, n92308,
    n92309, n92310, n92311, n92312, n92313, n92314, n92315, n92316, n92317,
    n92318, n92319, n92320, n92321, n92322, n92323, n92324, n92325, n92326,
    n92327, n92328, n92329, n92330, n92331, n92332, n92333, n92334, n92335,
    n92336, n92337, n92338, n92339, n92340, n92341, n92342, n92343, n92344,
    n92345, n92346, n92347, n92348, n92349, n92350, n92351, n92352, n92353,
    n92354, n92355, n92356, n92357, n92358, n92359, n92360, n92361, n92362,
    n92363, n92364, n92365, n92366, n92367, n92368, n92369, n92370, n92371,
    n92372, n92373, n92374, n92375, n92376, n92377, n92378, n92379, n92380,
    n92381, n92382, n92383, n92384, n92385, n92386, n92387, n92388, n92389,
    n92391, n92392, n92393, n92394, n92395, n92396, n92397, n92398, n92399,
    n92400, n92401, n92402, n92403, n92404, n92405, n92406, n92407, n92408,
    n92409, n92410, n92411, n92412, n92413, n92414, n92415, n92416, n92417,
    n92418, n92419, n92420, n92421, n92422, n92423, n92424, n92425, n92426,
    n92427, n92428, n92429, n92430, n92431, n92432, n92433, n92434, n92435,
    n92436, n92437, n92438, n92439, n92440, n92441, n92442, n92443, n92444,
    n92446, n92447, n92448, n92449, n92450, n92451, n92452, n92453, n92454,
    n92455, n92456, n92457, n92458, n92459, n92460, n92461, n92462, n92463,
    n92464, n92465, n92466, n92467, n92468, n92469, n92470, n92471, n92472,
    n92473, n92474, n92475, n92476, n92477, n92478, n92479, n92480, n92481,
    n92482, n92483, n92484, n92485, n92486, n92487, n92488, n92489, n92490,
    n92491, n92492, n92493, n92494, n92495, n92496, n92497, n92498, n92499,
    n92500, n92501, n92502, n92503, n92504, n92505, n92506, n92507, n92508,
    n92509, n92510, n92511, n92512, n92513, n92514, n92515, n92516, n92517,
    n92518, n92519, n92520, n92521, n92522, n92523, n92524, n92525, n92526,
    n92527, n92528, n92529, n92530, n92531, n92532, n92533, n92534, n92535,
    n92536, n92537, n92538, n92539, n92540, n92541, n92542, n92543, n92544,
    n92545, n92546, n92547, n92548, n92549, n92551, n92552, n92553, n92554,
    n92555, n92556, n92557, n92558, n92559, n92560, n92561, n92562, n92563,
    n92564, n92565, n92566, n92567, n92568, n92569, n92570, n92571, n92572,
    n92573, n92574, n92575, n92576, n92577, n92578, n92579, n92580, n92581,
    n92582, n92583, n92584, n92585, n92586, n92587, n92588, n92589, n92590,
    n92591, n92592, n92593, n92594, n92595, n92596, n92597, n92598, n92599,
    n92601, n92602, n92603, n92604, n92605, n92606, n92607, n92608, n92609,
    n92610, n92611, n92612, n92613, n92614, n92615, n92616, n92617, n92618,
    n92619, n92620, n92621, n92622, n92623, n92624, n92625, n92626, n92627,
    n92628, n92629, n92630, n92631, n92632, n92633, n92634, n92635, n92636,
    n92637, n92638, n92639, n92640, n92641, n92642, n92644, n92645, n92646,
    n92647, n92648, n92649, n92650, n92651, n92652, n92653, n92654, n92655,
    n92656, n92657, n92658, n92659, n92660, n92661, n92662, n92663, n92664,
    n92665, n92666, n92667, n92668, n92669, n92670, n92671, n92672, n92673,
    n92674, n92675, n92676, n92677, n92678, n92679, n92680, n92681, n92682,
    n92683, n92684, n92685, n92686, n92687, n92688, n92689, n92690, n92691,
    n92692, n92693, n92694, n92695, n92696, n92697, n92698, n92699, n92700,
    n92701, n92702, n92703, n92704, n92705, n92706, n92707, n92708, n92709,
    n92710, n92711, n92712, n92713, n92714, n92715, n92716, n92717, n92718,
    n92719, n92720, n92721, n92722, n92723, n92724, n92725, n92726, n92727,
    n92728, n92729, n92730, n92731, n92732, n92733, n92734, n92735, n92737,
    n92738, n92739, n92740, n92741, n92742, n92743, n92744, n92745, n92746,
    n92747, n92748, n92749, n92750, n92751, n92752, n92753, n92754, n92755,
    n92756, n92757, n92758, n92759, n92760, n92761, n92762, n92763, n92764,
    n92765, n92766, n92767, n92768, n92769, n92770, n92771, n92773, n92774,
    n92775, n92776, n92777, n92778, n92779, n92780, n92781, n92782, n92783,
    n92784, n92785, n92786, n92787, n92788, n92789, n92790, n92791, n92792,
    n92793, n92794, n92795, n92796, n92797, n92798, n92799, n92800, n92801,
    n92802, n92803, n92804, n92805, n92806, n92807, n92808, n92810, n92811,
    n92812, n92813, n92814, n92815, n92816, n92817, n92818, n92819, n92820,
    n92821, n92822, n92823, n92824, n92825, n92826, n92827, n92828, n92829,
    n92830, n92831, n92832, n92833, n92834, n92835, n92836, n92837, n92838,
    n92839, n92840, n92841, n92842, n92843, n92844, n92845, n92846, n92847,
    n92848, n92849, n92850, n92851, n92852, n92853, n92854, n92855, n92856,
    n92857, n92858, n92859, n92861, n92862, n92863, n92864, n92865, n92866,
    n92867, n92868, n92869, n92870, n92871, n92872, n92873, n92874, n92875,
    n92876, n92877, n92878, n92879, n92880, n92881, n92882, n92883, n92884,
    n92885, n92886, n92887, n92888, n92889, n92890, n92891, n92892, n92893,
    n92894, n92895, n92896, n92897, n92898, n92900, n92901, n92902, n92903,
    n92904, n92905, n92906, n92907, n92908, n92909, n92910, n92911, n92912,
    n92913, n92914, n92915, n92916, n92917, n92918, n92919, n92920, n92921,
    n92922, n92923, n92924, n92925, n92926, n92927, n92928, n92930, n92931,
    n92932, n92933, n92934, n92935, n92936, n92937, n92938, n92939, n92940,
    n92941, n92942, n92943, n92944, n92945, n92946, n92947, n92948, n92949,
    n92950, n92951, n92952, n92953, n92954, n92955, n92956, n92957, n92958,
    n92960, n92961, n92962, n92963, n92964, n92965, n92966, n92967, n92968,
    n92969, n92970, n92971, n92972, n92973, n92974, n92975, n92976, n92977,
    n92978, n92979, n92980, n92981, n92982, n92983, n92984, n92985, n92986,
    n92987, n92988, n92989, n92990, n92991, n92992, n92993, n92994, n92995,
    n92996, n92997, n92999, n93000, n93001, n93002, n93003, n93004, n93005,
    n93006, n93007, n93008, n93009, n93010, n93011, n93012, n93013, n93014,
    n93015, n93016, n93017, n93018, n93019, n93020, n93021, n93022, n93023,
    n93024, n93025, n93026, n93027, n93028, n93029, n93030, n93031, n93032,
    n93033, n93034, n93035, n93036, n93037, n93038, n93040, n93041, n93042,
    n93043, n93044, n93045, n93046, n93047, n93048, n93049, n93050, n93051,
    n93052, n93053, n93054, n93055, n93056, n93057, n93058, n93059, n93060,
    n93061, n93062, n93063, n93064, n93065, n93066, n93067, n93069, n93070,
    n93071, n93072, n93073, n93074, n93075, n93076, n93077, n93078, n93079,
    n93080, n93081, n93082, n93083, n93084, n93085, n93086, n93087, n93088,
    n93089, n93090, n93091, n93092, n93093, n93094, n93095, n93096, n93097,
    n93098, n93099, n93100, n93101, n93102, n93103, n93104, n93105, n93106,
    n93107, n93108, n93109, n93110, n93111, n93112, n93113, n93114, n93115,
    n93116, n93118, n93119, n93120, n93121, n93122, n93123, n93124, n93125,
    n93126, n93127, n93128, n93129, n93130, n93131, n93132, n93133, n93134,
    n93135, n93136, n93137, n93138, n93139, n93140, n93141, n93142, n93143,
    n93144, n93145, n93146, n93147, n93148, n93149, n93150, n93151, n93152,
    n93153, n93154, n93155, n93156, n93157, n93158, n93160, n93161, n93162,
    n93163, n93164, n93165, n93166, n93167, n93168, n93169, n93170, n93171,
    n93172, n93173, n93174, n93175, n93176, n93177, n93178, n93179, n93180,
    n93181, n93182, n93183, n93184, n93185, n93186, n93187, n93188, n93189,
    n93190, n93191, n93192, n93193, n93194, n93195, n93196, n93197, n93198,
    n93199, n93200, n93201, n93202, n93203, n93204, n93205, n93206, n93207,
    n93208, n93209, n93210, n93211, n93212, n93213, n93214, n93215, n93216,
    n93217, n93218, n93219, n93220, n93221, n93222, n93223, n93224, n93225,
    n93226, n93227, n93228, n93229, n93230, n93231, n93232, n93233, n93234,
    n93235, n93236, n93237, n93238, n93239, n93240, n93241, n93242, n93243,
    n93244, n93245, n93246, n93247, n93248, n93249, n93250, n93251, n93252,
    n93253, n93254, n93256, n93257, n93258, n93259, n93260, n93261, n93262,
    n93263, n93264, n93265, n93266, n93267, n93268, n93269, n93270, n93271,
    n93272, n93273, n93274, n93275, n93276, n93277, n93278, n93279, n93280,
    n93281, n93282, n93283, n93284, n93285, n93286, n93287, n93288, n93289,
    n93290, n93291, n93292, n93293, n93294, n93295, n93296, n93297, n93298,
    n93299, n93301, n93302, n93303, n93304, n93305, n93306, n93307, n93308,
    n93309, n93310, n93311, n93312, n93313, n93314, n93315, n93316, n93317,
    n93318, n93319, n93320, n93321, n93322, n93323, n93324, n93325, n93326,
    n93327, n93328, n93329, n93330, n93331, n93332, n93333, n93334, n93335,
    n93336, n93337, n93338, n93339, n93340, n93341, n93342, n93344, n93345,
    n93346, n93347, n93348, n93349, n93350, n93351, n93352, n93353, n93354,
    n93355, n93356, n93357, n93358, n93359, n93360, n93361, n93362, n93363,
    n93364, n93365, n93366, n93367, n93368, n93369, n93370, n93371, n93372,
    n93373, n93374, n93375, n93376, n93378, n93379, n93380, n93381, n93382,
    n93383, n93384, n93385, n93386, n93387, n93388, n93389, n93390, n93391,
    n93392, n93393, n93394, n93395, n93396, n93397, n93398, n93399, n93400,
    n93401, n93402, n93403, n93404, n93405, n93406, n93407, n93408, n93409,
    n93410, n93411, n93413, n93414, n93415, n93416, n93417, n93418, n93419,
    n93420, n93421, n93422, n93423, n93424, n93425, n93426, n93427, n93428,
    n93429, n93430, n93431, n93432, n93433, n93434, n93435, n93436, n93437,
    n93438, n93439, n93440, n93441, n93442, n93443, n93444, n93445, n93446,
    n93447, n93449, n93450, n93451, n93452, n93453, n93454, n93455, n93456,
    n93457, n93458, n93459, n93460, n93461, n93462, n93463, n93464, n93465,
    n93466, n93467, n93468, n93469, n93470, n93471, n93472, n93473, n93474,
    n93475, n93476, n93477, n93478, n93479, n93480, n93482, n93483, n93484,
    n93485, n93486, n93487, n93488, n93489, n93490, n93491, n93492, n93493,
    n93494, n93495, n93496, n93497, n93498, n93499, n93500, n93501, n93502,
    n93503, n93504, n93505, n93506, n93507, n93508, n93509, n93510, n93511,
    n93512, n93513, n93514, n93516, n93517, n93518, n93519, n93520, n93521,
    n93522, n93523, n93524, n93525, n93526, n93527, n93528, n93529, n93530,
    n93531, n93532, n93533, n93534, n93535, n93536, n93537, n93538, n93539,
    n93540, n93541, n93543, n93544, n93545, n93546, n93547, n93548, n93549,
    n93550, n93551, n93552, n93553, n93554, n93555, n93556, n93557, n93558,
    n93559, n93560, n93561, n93562, n93563, n93564, n93565, n93566, n93567,
    n93568, n93569, n93570, n93571, n93572, n93573, n93574, n93575, n93576,
    n93577, n93578, n93579, n93580, n93581, n93582, n93583, n93584, n93585,
    n93586, n93587, n93588, n93589, n93590, n93591, n93592, n93593, n93594,
    n93595, n93596, n93597, n93598, n93599, n93600, n93601, n93602, n93603,
    n93604, n93605, n93606, n93607, n93608, n93609, n93610, n93611, n93612,
    n93613, n93614, n93615, n93616, n93617, n93618, n93619, n93620, n93621,
    n93622, n93623, n93624, n93625, n93626, n93627, n93628, n93629, n93630,
    n93631, n93632, n93633, n93634, n93635, n93636, n93637, n93638, n93639,
    n93640, n93641, n93643, n93644, n93645, n93646, n93647, n93648, n93649,
    n93650, n93651, n93652, n93653, n93654, n93655, n93656, n93657, n93658,
    n93659, n93660, n93661, n93662, n93663, n93664, n93665, n93666, n93667,
    n93668, n93669, n93670, n93671, n93672, n93673, n93674, n93675, n93676,
    n93677, n93678, n93679, n93680, n93681, n93682, n93683, n93684, n93685,
    n93686, n93687, n93688, n93689, n93690, n93691, n93692, n93693, n93694,
    n93695, n93696, n93697, n93698, n93699, n93700, n93701, n93702, n93703,
    n93704, n93705, n93706, n93707, n93708, n93709, n93710, n93711, n93712,
    n93713, n93714, n93715, n93716, n93717, n93718, n93719, n93720, n93721,
    n93722, n93723, n93724, n93725, n93726, n93727, n93728, n93729, n93730,
    n93731, n93732, n93733, n93734, n93735, n93736, n93737, n93738, n93739,
    n93740, n93741, n93743, n93744, n93745, n93746, n93747, n93748, n93749,
    n93750, n93751, n93752, n93753, n93754, n93755, n93756, n93757, n93758,
    n93759, n93760, n93761, n93762, n93763, n93764, n93765, n93766, n93767,
    n93768, n93769, n93770, n93771, n93772, n93773, n93774, n93775, n93776,
    n93777, n93778, n93779, n93780, n93781, n93782, n93783, n93784, n93785,
    n93786, n93787, n93788, n93789, n93790, n93792, n93793, n93794, n93795,
    n93796, n93797, n93798, n93799, n93800, n93801, n93802, n93803, n93804,
    n93805, n93806, n93807, n93808, n93809, n93810, n93811, n93812, n93813,
    n93814, n93815, n93816, n93817, n93818, n93819, n93820, n93821, n93822,
    n93823, n93824, n93825, n93826, n93827, n93828, n93829, n93830, n93831,
    n93832, n93833, n93834, n93835, n93836, n93837, n93838, n93839, n93840,
    n93841, n93842, n93843, n93844, n93845, n93846, n93847, n93848, n93849,
    n93850, n93851, n93852, n93853, n93854, n93855, n93856, n93857, n93858,
    n93859, n93860, n93861, n93862, n93863, n93864, n93865, n93866, n93867,
    n93868, n93869, n93870, n93871, n93872, n93873, n93874, n93875, n93876,
    n93877, n93878, n93879, n93880, n93881, n93882, n93883, n93884, n93885,
    n93886, n93887, n93888, n93889, n93890, n93891, n93892, n93894, n93895,
    n93896, n93897, n93898, n93899, n93900, n93901, n93902, n93903, n93904,
    n93905, n93906, n93907, n93908, n93909, n93910, n93911, n93912, n93913,
    n93914, n93915, n93916, n93917, n93918, n93919, n93920, n93921, n93922,
    n93924, n93925, n93926, n93927, n93928, n93929, n93930, n93931, n93932,
    n93933, n93934, n93935, n93936, n93937, n93938, n93939, n93940, n93941,
    n93942, n93943, n93944, n93945, n93946, n93947, n93948, n93949, n93950,
    n93951, n93952, n93953, n93954, n93955, n93957, n93958, n93959, n93960,
    n93961, n93962, n93963, n93964, n93965, n93966, n93967, n93968, n93969,
    n93970, n93971, n93972, n93973, n93974, n93975, n93976, n93977, n93978,
    n93979, n93980, n93981, n93982, n93983, n93984, n93985, n93986, n93987,
    n93988, n93989, n93990, n93991, n93992, n93993, n93994, n93995, n93996,
    n93997, n93998, n93999, n94000, n94001, n94002, n94003, n94004, n94005,
    n94006, n94007, n94008, n94009, n94010, n94011, n94012, n94013, n94014,
    n94015, n94016, n94017, n94018, n94019, n94020, n94021, n94022, n94023,
    n94024, n94025, n94026, n94027, n94028, n94029, n94030, n94031, n94032,
    n94033, n94034, n94035, n94036, n94037, n94038, n94039, n94040, n94041,
    n94042, n94043, n94044, n94045, n94046, n94047, n94048, n94049, n94050,
    n94051, n94052, n94053, n94054, n94055, n94056, n94057, n94058, n94059,
    n94060, n94061, n94063, n94064, n94065, n94066, n94067, n94068, n94069,
    n94070, n94071, n94072, n94073, n94074, n94075, n94076, n94077, n94078,
    n94079, n94080, n94081, n94082, n94083, n94084, n94085, n94086, n94087,
    n94088, n94089, n94090, n94091, n94092, n94093, n94094, n94095, n94096,
    n94097, n94099, n94100, n94101, n94102, n94103, n94104, n94105, n94106,
    n94107, n94108, n94109, n94110, n94111, n94112, n94113, n94114, n94115,
    n94116, n94117, n94118, n94119, n94120, n94121, n94122, n94123, n94124,
    n94125, n94126, n94127, n94128, n94129, n94130, n94131, n94132, n94133,
    n94134, n94135, n94136, n94137, n94138, n94140, n94141, n94142, n94143,
    n94144, n94145, n94146, n94147, n94148, n94149, n94150, n94151, n94152,
    n94153, n94154, n94155, n94156, n94157, n94158, n94159, n94160, n94161,
    n94162, n94163, n94164, n94165, n94166, n94167, n94168, n94169, n94170,
    n94171, n94172, n94173, n94174, n94175, n94176, n94177, n94178, n94179,
    n94181, n94182, n94183, n94184, n94185, n94186, n94187, n94188, n94189,
    n94190, n94191, n94192, n94193, n94194, n94195, n94196, n94197, n94198,
    n94199, n94200, n94201, n94202, n94203, n94204, n94205, n94206, n94207,
    n94208, n94209, n94210, n94211, n94212, n94213, n94214, n94215, n94216,
    n94217, n94218, n94219, n94220, n94221, n94222, n94223, n94224, n94225,
    n94226, n94227, n94228, n94229, n94230, n94231, n94232, n94233, n94234,
    n94235, n94236, n94237, n94238, n94239, n94240, n94241, n94242, n94243,
    n94244, n94245, n94246, n94247, n94248, n94249, n94250, n94251, n94252,
    n94253, n94254, n94255, n94256, n94257, n94258, n94259, n94260, n94261,
    n94262, n94263, n94264, n94265, n94266, n94267, n94268, n94269, n94270,
    n94271, n94272, n94273, n94274, n94276, n94277, n94278, n94279, n94280,
    n94281, n94282, n94283, n94284, n94285, n94286, n94287, n94288, n94289,
    n94290, n94291, n94292, n94293, n94294, n94295, n94296, n94297, n94298,
    n94299, n94300, n94301, n94302, n94303, n94304, n94305, n94306, n94307,
    n94308, n94309, n94310, n94311, n94312, n94313, n94314, n94315, n94316,
    n94317, n94318, n94320, n94321, n94322, n94323, n94324, n94325, n94326,
    n94327, n94328, n94329, n94330, n94331, n94332, n94333, n94334, n94335,
    n94336, n94337, n94338, n94339, n94340, n94341, n94342, n94343, n94344,
    n94345, n94346, n94347, n94348, n94349, n94350, n94351, n94352, n94353,
    n94354, n94355, n94356, n94357, n94358, n94359, n94360, n94361, n94362,
    n94363, n94365, n94366, n94367, n94368, n94369, n94370, n94371, n94372,
    n94373, n94374, n94375, n94376, n94377, n94378, n94379, n94380, n94381,
    n94382, n94383, n94384, n94385, n94386, n94387, n94388, n94389, n94390,
    n94391, n94392, n94393, n94394, n94395, n94396, n94397, n94398, n94399,
    n94400, n94401, n94402, n94403, n94404, n94405, n94406, n94407, n94408,
    n94409, n94410, n94411, n94412, n94413, n94414, n94415, n94416, n94417,
    n94418, n94419, n94420, n94421, n94422, n94423, n94424, n94425, n94426,
    n94427, n94428, n94429, n94430, n94431, n94432, n94433, n94434, n94435,
    n94436, n94437, n94438, n94439, n94440, n94441, n94442, n94443, n94444,
    n94445, n94446, n94447, n94448, n94449, n94450, n94451, n94452, n94453,
    n94454, n94455, n94456, n94457, n94458, n94459, n94460, n94461, n94462,
    n94463, n94464, n94465, n94466, n94467, n94468, n94470, n94471, n94472,
    n94473, n94474, n94475, n94476, n94477, n94478, n94479, n94480, n94481,
    n94482, n94483, n94484, n94485, n94486, n94487, n94488, n94489, n94490,
    n94491, n94492, n94493, n94494, n94495, n94496, n94497, n94498, n94499,
    n94500, n94501, n94502, n94503, n94504, n94505, n94506, n94508, n94509,
    n94510, n94511, n94512, n94513, n94514, n94515, n94516, n94517, n94518,
    n94519, n94520, n94521, n94522, n94523, n94524, n94525, n94526, n94527,
    n94528, n94529, n94530, n94531, n94532, n94533, n94534, n94535, n94536,
    n94537, n94538, n94539, n94540, n94541, n94542, n94543, n94544, n94545,
    n94546, n94548, n94549, n94550, n94551, n94552, n94553, n94554, n94555,
    n94556, n94557, n94558, n94559, n94560, n94561, n94562, n94563, n94564,
    n94565, n94566, n94567, n94568, n94569, n94570, n94571, n94572, n94573,
    n94574, n94575, n94576, n94578, n94579, n94580, n94581, n94582, n94583,
    n94584, n94585, n94586, n94587, n94588, n94589, n94590, n94591, n94592,
    n94593, n94594, n94595, n94596, n94597, n94598, n94599, n94600, n94601,
    n94602, n94603, n94604, n94605, n94606, n94607, n94608, n94609, n94610,
    n94611, n94612, n94613, n94614, n94615, n94616, n94617, n94618, n94619,
    n94620, n94621, n94622, n94623, n94624, n94625, n94626, n94627, n94628,
    n94629, n94630, n94631, n94632, n94633, n94634, n94635, n94636, n94637,
    n94638, n94639, n94640, n94641, n94642, n94643, n94644, n94645, n94646,
    n94647, n94648, n94649, n94650, n94651, n94652, n94653, n94654, n94655,
    n94656, n94657, n94658, n94659, n94660, n94661, n94662, n94663, n94664,
    n94665, n94666, n94668, n94669, n94670, n94671, n94672, n94673, n94674,
    n94675, n94676, n94677, n94678, n94679, n94680, n94681, n94682, n94683,
    n94684, n94685, n94686, n94687, n94688, n94689, n94690, n94691, n94692,
    n94693, n94694, n94695, n94696, n94697, n94698, n94699, n94700, n94701,
    n94702, n94703, n94704, n94705, n94706, n94707, n94708, n94709, n94710,
    n94711, n94712, n94713, n94714, n94715, n94717, n94718, n94719, n94720,
    n94721, n94722, n94723, n94724, n94725, n94726, n94727, n94728, n94729,
    n94730, n94731, n94732, n94733, n94734, n94735, n94736, n94737, n94738,
    n94739, n94740, n94741, n94742, n94743, n94744, n94745, n94746, n94747,
    n94748, n94750, n94751, n94752, n94753, n94754, n94755, n94756, n94757,
    n94758, n94759, n94760, n94761, n94762, n94763, n94764, n94765, n94766,
    n94767, n94768, n94769, n94770, n94771, n94772, n94773, n94774, n94775,
    n94776, n94777, n94778, n94779, n94780, n94781, n94782, n94783, n94784,
    n94785, n94786, n94787, n94788, n94789, n94790, n94791, n94792, n94793,
    n94794, n94796, n94797, n94798, n94799, n94800, n94801, n94802, n94803,
    n94804, n94805, n94806, n94807, n94808, n94809, n94810, n94811, n94812,
    n94813, n94814, n94815, n94816, n94817, n94818, n94819, n94820, n94821,
    n94822, n94823, n94824, n94825, n94826, n94827, n94828, n94830, n94831,
    n94832, n94833, n94834, n94835, n94836, n94837, n94838, n94839, n94840,
    n94841, n94842, n94843, n94844, n94845, n94846, n94847, n94848, n94849,
    n94850, n94851, n94852, n94853, n94854, n94855, n94856, n94857, n94858,
    n94859, n94860, n94861, n94862, n94863, n94864, n94865, n94866, n94867,
    n94868, n94869, n94870, n94871, n94872, n94873, n94874, n94875, n94876,
    n94877, n94878, n94879, n94880, n94881, n94882, n94883, n94884, n94885,
    n94886, n94887, n94888, n94889, n94890, n94891, n94892, n94893, n94894,
    n94895, n94896, n94897, n94898, n94899, n94900, n94901, n94902, n94903,
    n94904, n94905, n94906, n94907, n94908, n94909, n94910, n94911, n94912,
    n94913, n94914, n94915, n94916, n94917, n94919, n94920, n94921, n94922,
    n94923, n94924, n94925, n94926, n94927, n94928, n94929, n94930, n94931,
    n94932, n94933, n94934, n94935, n94936, n94937, n94938, n94939, n94940,
    n94941, n94942, n94943, n94944, n94945, n94946, n94947, n94948, n94949,
    n94950, n94951, n94952, n94953, n94954, n94956, n94957, n94958, n94959,
    n94960, n94961, n94962, n94963, n94964, n94965, n94966, n94967, n94968,
    n94969, n94970, n94971, n94972, n94973, n94974, n94975, n94976, n94977,
    n94978, n94979, n94980, n94981, n94982, n94983, n94984, n94985, n94986,
    n94987, n94988, n94989, n94990, n94991, n94992, n94993, n94994, n94995,
    n94996, n94997, n94998, n94999, n95000, n95001, n95002, n95003, n95004,
    n95006, n95007, n95008, n95009, n95010, n95011, n95012, n95013, n95014,
    n95015, n95016, n95017, n95018, n95019, n95020, n95021, n95022, n95023,
    n95024, n95025, n95026, n95027, n95028, n95029, n95030, n95031, n95032,
    n95033, n95034, n95035, n95036, n95037, n95038, n95039, n95040, n95041,
    n95042, n95043, n95044, n95045, n95046, n95047, n95048, n95049, n95051,
    n95052, n95053, n95054, n95055, n95056, n95057, n95058, n95059, n95060,
    n95061, n95062, n95063, n95064, n95065, n95066, n95067, n95068, n95069,
    n95070, n95071, n95072, n95073, n95074, n95075, n95076, n95077, n95078,
    n95079, n95080, n95081, n95082, n95083, n95084, n95085, n95086, n95087,
    n95088, n95089, n95090, n95091, n95093, n95094, n95095, n95096, n95097,
    n95098, n95099, n95100, n95101, n95102, n95103, n95104, n95105, n95106,
    n95107, n95108, n95109, n95110, n95111, n95112, n95113, n95114, n95115,
    n95116, n95117, n95118, n95119, n95120, n95121, n95122, n95123, n95124,
    n95125, n95126, n95128, n95129, n95130, n95131, n95132, n95133, n95134,
    n95135, n95136, n95137, n95138, n95139, n95140, n95141, n95142, n95143,
    n95144, n95145, n95146, n95147, n95148, n95149, n95150, n95151, n95152,
    n95153, n95154, n95155, n95156, n95157, n95158, n95159, n95160, n95161,
    n95162, n95164, n95165, n95166, n95167, n95168, n95169, n95170, n95171,
    n95172, n95173, n95174, n95175, n95176, n95177, n95178, n95179, n95180,
    n95181, n95182, n95183, n95184, n95185, n95186, n95187, n95188, n95189,
    n95190, n95191, n95192, n95193, n95194, n95195, n95196, n95197, n95198,
    n95199, n95200, n95201, n95202, n95204, n95205, n95206, n95207, n95208,
    n95209, n95210, n95211, n95212, n95213, n95214, n95215, n95216, n95217,
    n95218, n95219, n95220, n95221, n95222, n95223, n95224, n95225, n95226,
    n95227, n95228, n95229, n95230, n95231, n95232, n95234, n95235, n95236,
    n95237, n95238, n95239, n95240, n95241, n95242, n95243, n95244, n95245,
    n95246, n95247, n95248, n95249, n95250, n95251, n95252, n95253, n95254,
    n95255, n95256, n95257, n95258, n95260, n95261, n95262, n95263, n95264,
    n95265, n95266, n95267, n95268, n95269, n95270, n95271, n95272, n95273,
    n95274, n95275, n95276, n95277, n95278, n95279, n95280, n95281, n95282,
    n95283, n95284, n95285, n95286, n95287, n95288, n95289, n95290, n95291,
    n95292, n95293, n95294, n95295, n95296, n95297, n95298, n95299, n95300,
    n95301, n95302, n95303, n95304, n95305, n95306, n95307, n95308, n95309,
    n95310, n95311, n95312, n95313, n95314, n95315, n95316, n95317, n95318,
    n95319, n95320, n95321, n95322, n95323, n95324, n95325, n95326, n95327,
    n95328, n95329, n95330, n95331, n95332, n95333, n95334, n95335, n95336,
    n95337, n95338, n95339, n95340, n95341, n95342, n95343, n95344, n95345,
    n95346, n95347, n95348, n95349, n95350, n95351, n95352, n95353, n95354,
    n95355, n95356, n95357, n95358, n95359, n95360, n95361, n95362, n95364,
    n95365, n95366, n95367, n95368, n95369, n95370, n95371, n95372, n95373,
    n95374, n95375, n95376, n95377, n95378, n95379, n95380, n95381, n95382,
    n95383, n95384, n95385, n95386, n95387, n95388, n95389, n95390, n95391,
    n95392, n95393, n95394, n95395, n95396, n95397, n95398, n95399, n95400,
    n95401, n95402, n95403, n95404, n95405, n95406, n95407, n95408, n95409,
    n95410, n95411, n95412, n95413, n95414, n95415, n95416, n95417, n95418,
    n95419, n95420, n95421, n95422, n95423, n95424, n95425, n95426, n95427,
    n95428, n95429, n95430, n95431, n95432, n95433, n95434, n95435, n95436,
    n95437, n95438, n95439, n95440, n95441, n95442, n95443, n95444, n95445,
    n95446, n95447, n95448, n95449, n95450, n95451, n95452, n95453, n95454,
    n95455, n95456, n95457, n95458, n95459, n95460, n95461, n95462, n95463,
    n95464, n95466, n95467, n95468, n95469, n95470, n95471, n95472, n95473,
    n95474, n95475, n95476, n95477, n95478, n95479, n95480, n95481, n95482,
    n95483, n95484, n95485, n95486, n95487, n95488, n95489, n95490, n95491,
    n95492, n95493, n95494, n95495, n95496, n95497, n95498, n95499, n95500,
    n95501, n95502, n95503, n95504, n95505, n95506, n95507, n95508, n95509,
    n95510, n95511, n95512, n95513, n95514, n95515, n95516, n95517, n95518,
    n95519, n95520, n95521, n95522, n95523, n95524, n95525, n95526, n95527,
    n95528, n95529, n95530, n95531, n95532, n95533, n95534, n95535, n95536,
    n95537, n95538, n95539, n95540, n95541, n95542, n95543, n95544, n95545,
    n95546, n95547, n95548, n95549, n95550, n95551, n95552, n95553, n95554,
    n95555, n95557, n95558, n95559, n95560, n95561, n95562, n95563, n95564,
    n95565, n95566, n95567, n95568, n95569, n95570, n95571, n95572, n95573,
    n95574, n95575, n95576, n95577, n95578, n95579, n95580, n95581, n95582,
    n95583, n95584, n95585, n95586, n95587, n95588, n95589, n95590, n95591,
    n95592, n95593, n95594, n95595, n95596, n95597, n95598, n95599, n95600,
    n95601, n95602, n95603, n95604, n95605, n95606, n95607, n95608, n95609,
    n95610, n95611, n95612, n95613, n95614, n95615, n95616, n95617, n95618,
    n95619, n95620, n95621, n95622, n95623, n95624, n95625, n95626, n95627,
    n95628, n95629, n95630, n95631, n95632, n95633, n95634, n95635, n95636,
    n95637, n95638, n95639, n95640, n95641, n95642, n95643, n95644, n95645,
    n95646, n95647, n95648, n95649, n95650, n95651, n95652, n95653, n95654,
    n95655, n95656, n95657, n95658, n95659, n95660, n95662, n95663, n95664,
    n95665, n95666, n95667, n95668, n95669, n95670, n95671, n95672, n95673,
    n95674, n95675, n95676, n95677, n95678, n95679, n95680, n95681, n95682,
    n95683, n95684, n95685, n95686, n95687, n95688, n95689, n95690, n95691,
    n95692, n95693, n95694, n95695, n95696, n95697, n95698, n95699, n95700,
    n95701, n95702, n95703, n95704, n95705, n95706, n95707, n95708, n95709,
    n95710, n95711, n95712, n95713, n95714, n95715, n95716, n95717, n95718,
    n95719, n95720, n95721, n95722, n95723, n95724, n95725, n95726, n95727,
    n95728, n95729, n95730, n95731, n95732, n95733, n95734, n95735, n95736,
    n95737, n95738, n95739, n95740, n95741, n95742, n95743, n95744, n95745,
    n95746, n95747, n95748, n95749, n95750, n95751, n95752, n95753, n95754,
    n95755, n95756, n95757, n95758, n95759, n95760, n95761, n95762, n95763,
    n95764, n95765, n95766, n95767, n95768, n95770, n95771, n95772, n95773,
    n95774, n95775, n95776, n95777, n95778, n95779, n95780, n95781, n95782,
    n95783, n95784, n95785, n95786, n95787, n95788, n95789, n95790, n95791,
    n95792, n95793, n95794, n95795, n95796, n95797, n95798, n95799, n95800,
    n95801, n95802, n95803, n95804, n95805, n95806, n95807, n95808, n95809,
    n95810, n95811, n95812, n95813, n95814, n95815, n95816, n95817, n95818,
    n95819, n95820, n95821, n95822, n95823, n95824, n95825, n95826, n95827,
    n95828, n95829, n95830, n95831, n95832, n95833, n95834, n95835, n95836,
    n95837, n95838, n95839, n95840, n95841, n95842, n95843, n95844, n95845,
    n95846, n95847, n95848, n95849, n95850, n95851, n95852, n95853, n95854,
    n95855, n95856, n95857, n95858, n95859, n95860, n95861, n95862, n95863,
    n95864, n95865, n95866, n95867, n95868, n95870, n95871, n95872, n95873,
    n95874, n95875, n95876, n95877, n95878, n95879, n95880, n95881, n95882,
    n95883, n95884, n95885, n95886, n95887, n95888, n95889, n95890, n95891,
    n95892, n95893, n95894, n95895, n95896, n95897, n95898, n95899, n95900,
    n95901, n95902, n95903, n95904, n95905, n95906, n95907, n95908, n95909,
    n95910, n95911, n95913, n95914, n95915, n95916, n95917, n95918, n95919,
    n95920, n95921, n95922, n95923, n95924, n95925, n95926, n95927, n95928,
    n95929, n95930, n95931, n95932, n95933, n95934, n95935, n95936, n95937,
    n95938, n95939, n95940, n95941, n95942, n95943, n95944, n95945, n95946,
    n95947, n95948, n95949, n95950, n95951, n95952, n95953, n95954, n95955,
    n95956, n95957, n95958, n95959, n95960, n95961, n95963, n95964, n95965,
    n95966, n95967, n95968, n95969, n95970, n95971, n95972, n95973, n95974,
    n95975, n95976, n95977, n95978, n95979, n95980, n95981, n95982, n95983,
    n95984, n95985, n95986, n95987, n95988, n95989, n95990, n95991, n95992,
    n95993, n95994, n95995, n95996, n95997, n95998, n95999, n96000, n96001,
    n96002, n96003, n96004, n96005, n96006, n96007, n96008, n96009, n96010,
    n96011, n96012, n96013, n96014, n96015, n96016, n96017, n96018, n96019,
    n96020, n96021, n96022, n96023, n96024, n96025, n96026, n96027, n96028,
    n96029, n96030, n96031, n96032, n96033, n96034, n96035, n96036, n96037,
    n96038, n96039, n96040, n96041, n96042, n96043, n96044, n96045, n96046,
    n96047, n96048, n96049, n96050, n96051, n96052, n96053, n96054, n96055,
    n96056, n96057, n96058, n96059, n96060, n96061, n96062, n96064, n96065,
    n96066, n96067, n96068, n96069, n96070, n96071, n96072, n96073, n96074,
    n96075, n96076, n96077, n96078, n96079, n96080, n96081, n96082, n96083,
    n96084, n96085, n96086, n96087, n96088, n96089, n96090, n96091, n96092,
    n96093, n96094, n96096, n96097, n96098, n96099, n96100, n96101, n96102,
    n96103, n96104, n96105, n96106, n96107, n96108, n96109, n96110, n96111,
    n96112, n96113, n96114, n96115, n96116, n96117, n96118, n96119, n96120,
    n96121, n96122, n96123, n96124, n96125, n96126, n96128, n96129, n96130,
    n96131, n96132, n96133, n96134, n96135, n96136, n96137, n96138, n96139,
    n96140, n96141, n96142, n96143, n96144, n96145, n96146, n96147, n96148,
    n96149, n96150, n96151, n96152, n96153, n96154, n96155, n96156, n96157,
    n96158, n96159, n96160, n96161, n96162, n96164, n96165, n96166, n96167,
    n96168, n96169, n96170, n96171, n96172, n96173, n96174, n96175, n96176,
    n96177, n96178, n96179, n96180, n96181, n96182, n96183, n96184, n96185,
    n96186, n96187, n96188, n96189, n96190, n96191, n96192, n96193, n96194,
    n96195, n96196, n96197, n96198, n96199, n96200, n96202, n96203, n96204,
    n96205, n96206, n96207, n96208, n96209, n96210, n96211, n96212, n96213,
    n96214, n96215, n96216, n96217, n96218, n96219, n96220, n96221, n96222,
    n96223, n96224, n96225, n96226, n96227, n96228, n96229, n96230, n96231,
    n96232, n96233, n96234, n96235, n96236, n96237, n96238, n96239, n96240,
    n96242, n96243, n96244, n96245, n96246, n96247, n96248, n96249, n96250,
    n96251, n96252, n96253, n96254, n96255, n96256, n96257, n96258, n96259,
    n96260, n96261, n96262, n96263, n96264, n96265, n96266, n96267, n96268,
    n96269, n96270, n96271, n96272, n96273, n96274, n96275, n96276, n96277,
    n96278, n96279, n96280, n96282, n96283, n96284, n96285, n96286, n96287,
    n96288, n96289, n96290, n96291, n96292, n96293, n96294, n96295, n96296,
    n96297, n96298, n96299, n96300, n96301, n96302, n96303, n96304, n96305,
    n96306, n96307, n96308, n96309, n96310, n96311, n96312, n96314, n96315,
    n96316, n96317, n96318, n96319, n96320, n96321, n96322, n96323, n96324,
    n96325, n96326, n96327, n96328, n96329, n96330, n96331, n96332, n96333,
    n96334, n96335, n96336, n96337, n96338, n96339, n96340, n96341, n96342,
    n96343, n96344, n96345, n96346, n96347, n96348, n96349, n96350, n96351,
    n96352, n96353, n96354, n96355, n96356, n96357, n96358, n96359, n96360,
    n96361, n96363, n96364, n96365, n96366, n96367, n96368, n96369, n96370,
    n96371, n96372, n96373, n96374, n96375, n96376, n96377, n96378, n96379,
    n96380, n96381, n96382, n96383, n96384, n96385, n96386, n96387, n96388,
    n96389, n96390, n96391, n96392, n96393, n96394, n96395, n96396, n96397,
    n96398, n96399, n96400, n96402, n96403, n96404, n96405, n96406, n96407,
    n96408, n96409, n96410, n96411, n96412, n96413, n96414, n96415, n96416,
    n96417, n96418, n96419, n96420, n96421, n96422, n96423, n96424, n96425,
    n96426, n96427, n96428, n96429, n96430, n96431, n96432, n96433, n96434,
    n96435, n96436, n96438, n96439, n96440, n96441, n96442, n96443, n96444,
    n96445, n96446, n96447, n96448, n96449, n96450, n96451, n96452, n96453,
    n96454, n96455, n96456, n96457, n96458, n96459, n96460, n96461, n96462,
    n96463, n96464, n96465, n96466, n96467, n96468, n96469, n96470, n96471,
    n96472, n96473, n96474, n96475, n96477, n96478, n96479, n96480, n96481,
    n96482, n96483, n96484, n96485, n96486, n96487, n96488, n96489, n96490,
    n96491, n96492, n96493, n96494, n96495, n96496, n96497, n96498, n96499,
    n96500, n96501, n96502, n96503, n96504, n96505, n96506, n96507, n96508,
    n96509, n96510, n96511, n96512, n96513, n96514, n96515, n96516, n96518,
    n96519, n96520, n96521, n96522, n96523, n96524, n96525, n96526, n96527,
    n96528, n96529, n96530, n96531, n96532, n96533, n96534, n96535, n96536,
    n96537, n96538, n96539, n96540, n96541, n96542, n96543, n96544, n96545,
    n96546, n96547, n96548, n96549, n96550, n96551, n96552, n96553, n96554,
    n96555, n96556, n96557, n96558, n96559, n96560, n96561, n96562, n96563,
    n96565, n96566, n96567, n96568, n96569, n96570, n96571, n96572, n96573,
    n96574, n96575, n96576, n96577, n96578, n96579, n96580, n96581, n96582,
    n96583, n96584, n96585, n96586, n96587, n96588, n96589, n96590, n96591,
    n96592, n96593, n96595, n96596, n96597, n96598, n96599, n96600, n96601,
    n96602, n96603, n96604, n96605, n96606, n96607, n96608, n96609, n96610,
    n96611, n96612, n96613, n96614, n96615, n96616, n96617, n96618, n96619,
    n96620, n96621, n96622, n96623, n96624, n96625, n96626, n96627, n96628,
    n96629, n96630, n96631, n96632, n96633, n96634, n96635, n96636, n96637,
    n96638, n96640, n96641, n96642, n96643, n96644, n96645, n96646, n96647,
    n96648, n96649, n96650, n96651, n96652, n96653, n96654, n96655, n96656,
    n96657, n96658, n96659, n96660, n96661, n96662, n96663, n96664, n96665,
    n96666, n96667, n96668, n96669, n96670, n96671, n96672, n96673, n96674,
    n96675, n96676, n96677, n96679, n96680, n96681, n96682, n96683, n96684,
    n96685, n96686, n96687, n96688, n96689, n96690, n96691, n96692, n96693,
    n96694, n96695, n96696, n96697, n96698, n96699, n96700, n96701, n96702,
    n96703, n96704, n96705, n96706, n96707, n96708, n96709, n96710, n96711,
    n96712, n96713, n96714, n96715, n96716, n96717, n96718, n96719, n96720,
    n96721, n96722, n96723, n96724, n96725, n96726, n96727, n96728, n96729,
    n96730, n96731, n96732, n96733, n96734, n96735, n96736, n96737, n96738,
    n96739, n96740, n96741, n96742, n96743, n96744, n96745, n96746, n96747,
    n96748, n96749, n96750, n96751, n96752, n96753, n96754, n96755, n96756,
    n96757, n96758, n96759, n96760, n96761, n96762, n96763, n96764, n96765,
    n96766, n96767, n96768, n96769, n96770, n96771, n96772, n96773, n96774,
    n96775, n96777, n96778, n96779, n96780, n96781, n96782, n96783, n96784,
    n96785, n96786, n96787, n96788, n96789, n96790, n96791, n96792, n96793,
    n96794, n96795, n96796, n96797, n96798, n96799, n96800, n96801, n96803,
    n96804, n96805, n96806, n96807, n96808, n96809, n96810, n96811, n96812,
    n96813, n96814, n96815, n96816, n96817, n96818, n96819, n96820, n96821,
    n96822, n96823, n96824, n96825, n96826, n96827, n96828, n96829, n96830,
    n96831, n96832, n96833, n96835, n96836, n96837, n96838, n96839, n96840,
    n96841, n96842, n96843, n96844, n96845, n96846, n96847, n96848, n96849,
    n96850, n96851, n96852, n96853, n96854, n96855, n96856, n96857, n96858,
    n96859, n96860, n96861, n96862, n96863, n96864, n96865, n96866, n96867,
    n96868, n96869, n96870, n96871, n96872, n96873, n96874, n96876, n96877,
    n96878, n96879, n96880, n96881, n96882, n96883, n96884, n96885, n96886,
    n96887, n96888, n96889, n96890, n96891, n96892, n96893, n96894, n96895,
    n96896, n96897, n96898, n96899, n96900, n96901, n96902, n96903, n96904,
    n96905, n96906, n96907, n96908, n96909, n96910, n96911, n96912, n96914,
    n96915, n96916, n96917, n96918, n96919, n96920, n96921, n96922, n96923,
    n96924, n96925, n96926, n96927, n96928, n96929, n96930, n96931, n96932,
    n96933, n96934, n96935, n96936, n96937, n96938, n96939, n96940, n96941,
    n96942, n96944, n96945, n96946, n96947, n96948, n96949, n96950, n96951,
    n96952, n96953, n96954, n96955, n96956, n96957, n96958, n96959, n96960,
    n96961, n96962, n96963, n96964, n96965, n96966, n96967, n96968, n96969,
    n96970, n96971, n96972, n96973, n96974, n96975, n96976, n96977, n96979,
    n96980, n96981, n96982, n96983, n96984, n96985, n96986, n96987, n96988,
    n96989, n96990, n96991, n96992, n96993, n96994, n96995, n96996, n96997,
    n96998, n96999, n97000, n97001, n97002, n97003, n97004, n97005, n97006,
    n97007, n97008, n97009, n97010, n97011, n97012, n97013, n97014, n97015,
    n97016, n97017, n97018, n97019, n97020, n97021, n97022, n97023, n97024,
    n97025, n97026, n97027, n97028, n97029, n97030, n97031, n97032, n97033,
    n97034, n97035, n97036, n97037, n97038, n97039, n97040, n97041, n97042,
    n97043, n97044, n97045, n97046, n97047, n97048, n97049, n97050, n97051,
    n97052, n97053, n97054, n97055, n97056, n97057, n97058, n97059, n97060,
    n97061, n97062, n97063, n97064, n97065, n97066, n97067, n97068, n97069,
    n97070, n97071, n97072, n97073, n97074, n97075, n97076, n97077, n97078,
    n97079, n97080, n97082, n97083, n97084, n97085, n97086, n97087, n97088,
    n97089, n97090, n97091, n97092, n97093, n97094, n97095, n97096, n97097,
    n97098, n97099, n97100, n97101, n97102, n97103, n97104, n97105, n97106,
    n97107, n97108, n97109, n97110, n97111, n97112, n97113, n97114, n97115,
    n97116, n97117, n97118, n97119, n97120, n97121, n97122, n97123, n97124,
    n97125, n97126, n97127, n97128, n97129, n97130, n97131, n97132, n97133,
    n97134, n97135, n97136, n97137, n97138, n97139, n97140, n97141, n97142,
    n97143, n97144, n97145, n97146, n97147, n97148, n97149, n97150, n97151,
    n97152, n97153, n97154, n97155, n97156, n97157, n97158, n97159, n97160,
    n97161, n97162, n97163, n97164, n97165, n97166, n97167, n97168, n97169,
    n97170, n97171, n97172, n97173, n97174, n97175, n97176, n97177, n97178,
    n97179, n97180, n97181, n97182, n97183, n97184, n97185, n97186, n97187,
    n97188, n97190, n97191, n97192, n97193, n97194, n97195, n97196, n97197,
    n97198, n97199, n97200, n97201, n97202, n97203, n97204, n97205, n97206,
    n97207, n97208, n97209, n97210, n97211, n97212, n97213, n97214, n97215,
    n97216, n97217, n97218, n97219, n97221, n97222, n97223, n97224, n97225,
    n97226, n97227, n97228, n97229, n97230, n97231, n97232, n97233, n97234,
    n97235, n97236, n97237, n97238, n97239, n97240, n97241, n97242, n97243,
    n97244, n97245, n97246, n97247, n97248, n97249, n97250, n97251, n97252,
    n97253, n97254, n97255, n97256, n97257, n97258, n97259, n97260, n97261,
    n97262, n97263, n97264, n97265, n97266, n97267, n97268, n97269, n97270,
    n97271, n97272, n97273, n97274, n97275, n97276, n97277, n97278, n97279,
    n97280, n97281, n97282, n97283, n97284, n97285, n97286, n97287, n97288,
    n97289, n97290, n97291, n97292, n97293, n97294, n97295, n97296, n97297,
    n97298, n97299, n97300, n97301, n97302, n97303, n97304, n97305, n97306,
    n97307, n97308, n97309, n97310, n97311, n97312, n97313, n97314, n97315,
    n97316, n97317, n97318, n97319, n97320, n97321, n97322, n97324, n97325,
    n97326, n97327, n97328, n97329, n97330, n97331, n97332, n97333, n97334,
    n97335, n97336, n97337, n97338, n97339, n97340, n97341, n97342, n97343,
    n97344, n97345, n97346, n97347, n97348, n97349, n97350, n97351, n97352,
    n97353, n97354, n97355, n97356, n97357, n97358, n97359, n97360, n97361,
    n97362, n97363, n97364, n97365, n97366, n97367, n97368, n97369, n97370,
    n97371, n97372, n97373, n97374, n97375, n97376, n97377, n97378, n97379,
    n97380, n97381, n97382, n97383, n97384, n97385, n97386, n97387, n97388,
    n97389, n97390, n97391, n97392, n97393, n97394, n97395, n97396, n97397,
    n97398, n97399, n97400, n97401, n97402, n97403, n97404, n97405, n97406,
    n97407, n97408, n97409, n97410, n97411, n97412, n97413, n97414, n97415,
    n97416, n97417, n97418, n97419, n97420, n97421, n97423, n97424, n97425,
    n97426, n97427, n97428, n97429, n97430, n97431, n97432, n97433, n97434,
    n97435, n97436, n97437, n97438, n97439, n97440, n97441, n97442, n97443,
    n97444, n97445, n97446, n97447, n97448, n97449, n97450, n97451, n97452,
    n97453, n97454, n97455, n97456, n97457, n97458, n97459, n97460, n97461,
    n97462, n97463, n97464, n97465, n97466, n97467, n97468, n97469, n97471,
    n97472, n97473, n97474, n97475, n97476, n97477, n97478, n97479, n97480,
    n97481, n97482, n97483, n97484, n97485, n97486, n97487, n97488, n97489,
    n97490, n97491, n97492, n97493, n97494, n97495, n97496, n97497, n97498,
    n97499, n97500, n97501, n97502, n97503, n97504, n97505, n97506, n97507,
    n97508, n97509, n97511, n97512, n97513, n97514, n97515, n97516, n97517,
    n97518, n97519, n97520, n97521, n97522, n97523, n97524, n97525, n97526,
    n97527, n97528, n97529, n97530, n97531, n97532, n97533, n97534, n97535,
    n97536, n97537, n97538, n97539, n97540, n97541, n97542, n97543, n97544,
    n97545, n97546, n97547, n97548, n97549, n97550, n97551, n97552, n97553,
    n97554, n97555, n97556, n97557, n97558, n97559, n97560, n97561, n97562,
    n97563, n97564, n97565, n97566, n97567, n97568, n97569, n97570, n97571,
    n97572, n97573, n97574, n97575, n97576, n97577, n97578, n97579, n97580,
    n97581, n97582, n97583, n97584, n97585, n97586, n97587, n97588, n97589,
    n97590, n97591, n97592, n97593, n97594, n97595, n97596, n97597, n97598,
    n97599, n97600, n97601, n97602, n97603, n97604, n97605, n97606, n97608,
    n97609, n97610, n97611, n97612, n97613, n97614, n97615, n97616, n97617,
    n97618, n97619, n97620, n97621, n97622, n97623, n97624, n97625, n97626,
    n97627, n97628, n97629, n97630, n97631, n97632, n97633, n97634, n97635,
    n97636, n97637, n97638, n97639, n97640, n97641, n97642, n97643, n97644,
    n97645, n97646, n97647, n97648, n97649, n97650, n97651, n97652, n97654,
    n97655, n97656, n97657, n97658, n97659, n97660, n97661, n97662, n97663,
    n97664, n97665, n97666, n97667, n97668, n97669, n97670, n97671, n97672,
    n97673, n97674, n97675, n97676, n97677, n97678, n97679, n97680, n97681,
    n97682, n97683, n97684, n97686, n97687, n97688, n97689, n97690, n97691,
    n97692, n97693, n97694, n97695, n97696, n97697, n97698, n97699, n97700,
    n97701, n97702, n97703, n97704, n97705, n97706, n97707, n97708, n97709,
    n97710, n97711, n97712, n97713, n97714, n97715, n97716, n97717, n97718,
    n97719, n97720, n97721, n97722, n97723, n97724, n97725, n97726, n97727,
    n97728, n97729, n97730, n97731, n97732, n97733, n97734, n97735, n97736,
    n97737, n97738, n97739, n97740, n97741, n97742, n97743, n97744, n97745,
    n97746, n97747, n97748, n97749, n97750, n97751, n97752, n97753, n97754,
    n97755, n97756, n97757, n97758, n97759, n97760, n97761, n97762, n97763,
    n97764, n97765, n97766, n97767, n97768, n97769, n97770, n97771, n97772,
    n97773, n97774, n97775, n97777, n97778, n97779, n97780, n97781, n97782,
    n97783, n97784, n97785, n97786, n97787, n97788, n97789, n97790, n97791,
    n97792, n97793, n97794, n97795, n97796, n97797, n97798, n97799, n97800,
    n97801, n97802, n97803, n97804, n97805, n97806, n97807, n97808, n97809,
    n97810, n97811, n97813, n97814, n97815, n97816, n97817, n97818, n97819,
    n97820, n97821, n97822, n97823, n97824, n97825, n97826, n97827, n97828,
    n97829, n97830, n97831, n97832, n97833, n97834, n97835, n97836, n97837,
    n97838, n97839, n97840, n97841, n97842, n97843, n97844, n97845, n97846,
    n97847, n97849, n97850, n97851, n97852, n97853, n97854, n97855, n97856,
    n97857, n97858, n97859, n97860, n97861, n97862, n97863, n97864, n97865,
    n97866, n97867, n97868, n97869, n97870, n97871, n97872, n97873, n97874,
    n97875, n97876, n97877, n97878, n97879, n97880, n97881, n97882, n97883,
    n97884, n97885, n97886, n97887, n97888, n97889, n97890, n97891, n97893,
    n97894, n97895, n97896, n97897, n97898, n97899, n97900, n97901, n97902,
    n97903, n97904, n97905, n97906, n97907, n97908, n97909, n97910, n97911,
    n97912, n97913, n97914, n97915, n97916, n97917, n97918, n97919, n97920,
    n97921, n97922, n97923, n97924, n97925, n97926, n97927, n97928, n97929,
    n97930, n97931, n97932, n97933, n97934, n97936, n97937, n97938, n97939,
    n97940, n97941, n97942, n97943, n97944, n97945, n97946, n97947, n97948,
    n97949, n97950, n97951, n97952, n97953, n97954, n97955, n97956, n97957,
    n97958, n97959, n97960, n97961, n97962, n97963, n97964, n97965, n97966,
    n97967, n97968, n97969, n97970, n97971, n97972, n97973, n97974, n97975,
    n97977, n97978, n97979, n97980, n97981, n97982, n97983, n97984, n97985,
    n97986, n97987, n97988, n97989, n97990, n97991, n97992, n97993, n97994,
    n97995, n97996, n97997, n97998, n97999, n98000, n98001, n98002, n98003,
    n98004, n98005, n98006, n98007, n98008, n98009, n98010, n98011, n98012,
    n98013, n98014, n98015, n98016, n98017, n98018, n98019, n98020, n98021,
    n98022, n98023, n98024, n98025, n98026, n98027, n98028, n98029, n98030,
    n98031, n98032, n98033, n98034, n98035, n98036, n98037, n98038, n98039,
    n98040, n98041, n98042, n98043, n98044, n98045, n98046, n98047, n98048,
    n98049, n98050, n98051, n98052, n98053, n98054, n98055, n98056, n98057,
    n98058, n98059, n98060, n98061, n98062, n98063, n98064, n98065, n98066,
    n98067, n98068, n98069, n98071, n98072, n98073, n98074, n98075, n98076,
    n98077, n98078, n98079, n98080, n98081, n98082, n98083, n98084, n98085,
    n98086, n98087, n98088, n98089, n98090, n98091, n98092, n98093, n98094,
    n98095, n98096, n98097, n98098, n98099, n98100, n98101, n98102, n98103,
    n98104, n98105, n98106, n98107, n98108, n98109, n98110, n98111, n98113,
    n98114, n98115, n98116, n98117, n98118, n98119, n98120, n98121, n98122,
    n98123, n98124, n98125, n98126, n98127, n98128, n98129, n98130, n98131,
    n98132, n98133, n98134, n98135, n98136, n98137, n98138, n98139, n98140,
    n98141, n98142, n98143, n98144, n98145, n98146, n98147, n98148, n98149,
    n98150, n98151, n98152, n98153, n98154, n98155, n98156, n98157, n98159,
    n98160, n98161, n98162, n98163, n98164, n98165, n98166, n98167, n98168,
    n98169, n98170, n98171, n98172, n98173, n98174, n98175, n98176, n98177,
    n98178, n98179, n98180, n98181, n98182, n98183, n98184, n98185, n98186,
    n98187, n98188, n98189, n98190, n98191, n98193, n98194, n98195, n98196,
    n98197, n98198, n98199, n98200, n98201, n98202, n98203, n98204, n98205,
    n98206, n98207, n98208, n98209, n98210, n98211, n98212, n98213, n98214,
    n98215, n98216, n98217, n98218, n98219, n98220, n98221, n98222, n98223,
    n98224, n98225, n98226, n98227, n98228, n98229, n98230, n98231, n98232,
    n98233, n98234, n98235, n98236, n98237, n98238, n98239, n98240, n98241,
    n98242, n98243, n98244, n98245, n98246, n98247, n98248, n98249, n98250,
    n98251, n98252, n98253, n98254, n98255, n98256, n98257, n98258, n98259,
    n98260, n98261, n98262, n98263, n98264, n98265, n98266, n98267, n98268,
    n98269, n98270, n98271, n98272, n98273, n98274, n98275, n98276, n98277,
    n98278, n98279, n98280, n98281, n98282, n98283, n98284, n98285, n98286,
    n98287, n98288, n98289, n98290, n98292, n98293, n98294, n98295, n98296,
    n98297, n98298, n98299, n98300, n98301, n98302, n98303, n98304, n98305,
    n98306, n98307, n98308, n98309, n98310, n98311, n98312, n98313, n98314,
    n98315, n98316, n98317, n98318, n98319, n98320, n98322, n98323, n98324,
    n98325, n98326, n98327, n98328, n98329, n98330, n98331, n98332, n98333,
    n98334, n98335, n98336, n98337, n98338, n98339, n98340, n98341, n98342,
    n98343, n98344, n98345, n98346, n98347, n98348, n98349, n98350, n98351,
    n98352, n98353, n98354, n98355, n98357, n98358, n98359, n98360, n98361,
    n98362, n98363, n98364, n98365, n98366, n98367, n98368, n98369, n98370,
    n98371, n98372, n98373, n98374, n98375, n98376, n98377, n98378, n98379,
    n98380, n98381, n98382, n98383, n98384, n98385, n98386, n98387, n98388,
    n98389, n98390, n98391, n98392, n98393, n98394, n98395, n98396, n98397,
    n98398, n98399, n98400, n98401, n98402, n98403, n98405, n98406, n98407,
    n98408, n98409, n98410, n98411, n98412, n98413, n98414, n98415, n98416,
    n98417, n98418, n98419, n98420, n98421, n98422, n98423, n98424, n98425,
    n98426, n98427, n98428, n98429, n98430, n98431, n98432, n98433, n98434,
    n98435, n98436, n98437, n98438, n98439, n98440, n98441, n98442, n98443,
    n98444, n98445, n98446, n98448, n98449, n98450, n98451, n98452, n98453,
    n98454, n98455, n98456, n98457, n98458, n98459, n98460, n98461, n98462,
    n98463, n98464, n98465, n98466, n98467, n98468, n98469, n98470, n98471,
    n98472, n98473, n98474, n98475, n98476, n98477, n98478, n98480, n98481,
    n98482, n98483, n98484, n98485, n98486, n98487, n98488, n98489, n98490,
    n98491, n98492, n98493, n98494, n98495, n98496, n98497, n98498, n98499,
    n98500, n98501, n98502, n98503, n98504, n98505, n98506, n98507, n98508,
    n98509, n98510, n98511, n98512, n98513, n98514, n98515, n98516, n98518,
    n98519, n98520, n98521, n98522, n98523, n98524, n98525, n98526, n98527,
    n98528, n98529, n98530, n98531, n98532, n98533, n98534, n98535, n98536,
    n98537, n98538, n98539, n98540, n98541, n98542, n98543, n98544, n98545,
    n98546, n98547, n98548, n98549, n98550, n98551, n98552, n98553, n98554,
    n98555, n98556, n98557, n98559, n98560, n98561, n98562, n98563, n98564,
    n98565, n98566, n98567, n98568, n98569, n98570, n98571, n98572, n98573,
    n98574, n98575, n98576, n98577, n98578, n98579, n98580, n98581, n98582,
    n98583, n98584, n98585, n98586, n98587, n98588, n98589, n98590, n98591,
    n98592, n98594, n98595, n98596, n98597, n98598, n98599, n98600, n98601,
    n98602, n98603, n98604, n98605, n98606, n98607, n98608, n98609, n98610,
    n98611, n98612, n98613, n98614, n98615, n98616, n98617, n98618, n98619,
    n98620, n98621, n98622, n98623, n98624, n98625, n98626, n98627, n98628,
    n98629, n98630, n98631, n98632, n98633, n98634, n98635, n98636, n98637,
    n98638, n98639, n98641, n98642, n98643, n98644, n98645, n98646, n98647,
    n98648, n98649, n98650, n98651, n98652, n98653, n98654, n98655, n98656,
    n98657, n98658, n98659, n98660, n98661, n98662, n98663, n98664, n98665,
    n98667, n98668, n98669, n98670, n98671, n98672, n98673, n98674, n98675,
    n98676, n98677, n98678, n98679, n98680, n98681, n98682, n98683, n98684,
    n98685, n98686, n98687, n98688, n98689, n98690, n98691, n98692, n98693,
    n98694, n98695, n98697, n98698, n98699, n98700, n98701, n98702, n98703,
    n98704, n98705, n98706, n98707, n98708, n98709, n98710, n98711, n98712,
    n98713, n98714, n98715, n98716, n98717, n98718, n98719, n98720, n98721,
    n98722, n98723, n98724, n98725, n98726, n98727, n98728, n98729, n98730,
    n98731, n98732, n98733, n98734, n98735, n98736, n98737, n98738, n98739,
    n98740, n98741, n98742, n98743, n98744, n98745, n98746, n98747, n98748,
    n98749, n98750, n98751, n98752, n98753, n98754, n98755, n98756, n98757,
    n98758, n98759, n98760, n98761, n98762, n98763, n98764, n98765, n98766,
    n98767, n98768, n98769, n98770, n98771, n98772, n98773, n98774, n98775,
    n98776, n98777, n98778, n98779, n98780, n98781, n98782, n98783, n98784,
    n98785, n98786, n98787, n98788, n98789, n98790, n98791, n98792, n98793,
    n98794, n98795, n98797, n98798, n98799, n98800, n98801, n98802, n98803,
    n98804, n98805, n98806, n98807, n98808, n98809, n98810, n98811, n98812,
    n98813, n98814, n98815, n98816, n98817, n98818, n98819, n98820, n98821,
    n98822, n98823, n98824, n98825, n98826, n98827, n98828, n98829, n98830,
    n98831, n98832, n98833, n98834, n98835, n98836, n98837, n98838, n98839,
    n98840, n98841, n98842, n98843, n98845, n98846, n98847, n98848, n98849,
    n98850, n98851, n98852, n98853, n98854, n98855, n98856, n98857, n98858,
    n98859, n98860, n98861, n98862, n98863, n98864, n98865, n98866, n98867,
    n98868, n98869, n98870, n98871, n98872, n98873, n98874, n98875, n98876,
    n98877, n98878, n98879, n98880, n98881, n98882, n98883, n98884, n98885,
    n98886, n98887, n98888, n98889, n98890, n98891, n98892, n98893, n98894,
    n98895, n98896, n98897, n98898, n98899, n98900, n98901, n98902, n98903,
    n98904, n98905, n98906, n98907, n98908, n98909, n98910, n98911, n98912,
    n98913, n98914, n98915, n98916, n98917, n98918, n98919, n98920, n98921,
    n98922, n98923, n98924, n98925, n98926, n98927, n98928, n98929, n98930,
    n98931, n98932, n98933, n98934, n98935, n98936, n98937, n98938, n98939,
    n98940, n98941, n98942, n98943, n98944, n98945, n98946, n98947, n98948,
    n98949, n98950, n98951, n98953, n98954, n98955, n98956, n98957, n98958,
    n98959, n98960, n98961, n98962, n98963, n98964, n98965, n98966, n98967,
    n98968, n98969, n98970, n98971, n98972, n98973, n98974, n98975, n98976,
    n98977, n98978, n98979, n98980, n98981, n98982, n98983, n98984, n98985,
    n98986, n98987, n98988, n98989, n98990, n98991, n98992, n98993, n98994,
    n98995, n98996, n98997, n98998, n98999, n99000, n99001, n99002, n99003,
    n99004, n99005, n99006, n99007, n99008, n99009, n99010, n99011, n99012,
    n99013, n99014, n99015, n99016, n99017, n99018, n99019, n99020, n99021,
    n99022, n99023, n99024, n99025, n99026, n99027, n99028, n99029, n99030,
    n99031, n99032, n99033, n99034, n99035, n99036, n99037, n99038, n99039,
    n99040, n99041, n99042, n99043, n99044, n99045, n99046, n99047, n99048,
    n99049, n99050, n99051, n99052, n99053, n99054, n99056, n99057, n99058,
    n99059, n99060, n99061, n99062, n99063, n99064, n99065, n99066, n99067,
    n99068, n99069, n99070, n99071, n99072, n99073, n99074, n99075, n99076,
    n99077, n99078, n99079, n99080, n99081, n99082, n99083, n99084, n99085,
    n99086, n99087, n99088, n99089, n99090, n99091, n99092, n99093, n99094,
    n99095, n99096, n99097, n99098, n99099, n99100, n99101, n99102, n99103,
    n99104, n99105, n99106, n99107, n99108, n99109, n99110, n99111, n99112,
    n99113, n99114, n99115, n99116, n99117, n99118, n99119, n99120, n99121,
    n99122, n99123, n99124, n99125, n99126, n99127, n99128, n99129, n99130,
    n99131, n99132, n99133, n99134, n99135, n99136, n99137, n99138, n99139,
    n99140, n99141, n99142, n99143, n99144, n99145, n99146, n99147, n99148,
    n99149, n99150, n99151, n99152, n99153, n99154, n99155, n99157, n99158,
    n99159, n99160, n99161, n99162, n99163, n99164, n99165, n99166, n99167,
    n99168, n99169, n99170, n99171, n99172, n99173, n99174, n99175, n99176,
    n99177, n99178, n99179, n99180, n99181, n99182, n99183, n99184, n99185,
    n99186, n99187, n99188, n99189, n99190, n99191, n99192, n99193, n99194,
    n99195, n99196, n99197, n99198, n99199, n99200, n99201, n99202, n99203,
    n99204, n99205, n99206, n99207, n99208, n99209, n99210, n99211, n99212,
    n99213, n99214, n99215, n99216, n99217, n99218, n99219, n99220, n99221,
    n99222, n99223, n99224, n99225, n99226, n99227, n99228, n99229, n99230,
    n99231, n99232, n99233, n99234, n99235, n99236, n99237, n99238, n99239,
    n99240, n99241, n99242, n99243, n99244, n99246, n99247, n99248, n99249,
    n99250, n99251, n99252, n99253, n99254, n99255, n99256, n99257, n99258,
    n99259, n99260, n99261, n99262, n99263, n99264, n99265, n99266, n99267,
    n99268, n99269, n99270, n99271, n99272, n99273, n99274, n99275, n99276,
    n99277, n99278, n99279, n99280, n99281, n99282, n99283, n99284, n99285,
    n99286, n99287, n99288, n99289, n99290, n99291, n99293, n99294, n99295,
    n99296, n99297, n99298, n99299, n99300, n99301, n99302, n99303, n99304,
    n99305, n99306, n99307, n99308, n99309, n99310, n99311, n99312, n99313,
    n99314, n99315, n99316, n99317, n99318, n99319, n99320, n99321, n99322,
    n99323, n99324, n99325, n99326, n99327, n99328, n99329, n99330, n99331,
    n99332, n99333, n99334, n99335, n99336, n99337, n99338, n99339, n99340,
    n99341, n99342, n99343, n99344, n99345, n99346, n99347, n99348, n99349,
    n99350, n99351, n99352, n99353, n99354, n99355, n99356, n99357, n99358,
    n99359, n99360, n99361, n99362, n99363, n99364, n99365, n99366, n99367,
    n99368, n99369, n99370, n99371, n99372, n99373, n99374, n99375, n99376,
    n99377, n99378, n99379, n99380, n99381, n99382, n99383, n99384, n99385,
    n99386, n99387, n99388, n99389, n99390, n99391, n99393, n99394, n99395,
    n99396, n99397, n99398, n99399, n99400, n99401, n99402, n99403, n99404,
    n99405, n99406, n99407, n99408, n99409, n99410, n99411, n99412, n99413,
    n99414, n99415, n99416, n99417, n99418, n99419, n99420, n99421, n99422,
    n99423, n99424, n99425, n99426, n99427, n99428, n99429, n99430, n99431,
    n99432, n99433, n99434, n99435, n99436, n99437, n99438, n99439, n99440,
    n99441, n99443, n99444, n99445, n99446, n99447, n99448, n99449, n99450,
    n99451, n99452, n99453, n99454, n99455, n99456, n99457, n99458, n99459,
    n99460, n99461, n99462, n99463, n99464, n99465, n99466, n99467, n99468,
    n99469, n99470, n99471, n99472, n99473, n99474, n99475, n99477, n99478,
    n99479, n99480, n99481, n99482, n99483, n99484, n99485, n99486, n99487,
    n99488, n99489, n99490, n99491, n99492, n99493, n99494, n99495, n99496,
    n99497, n99498, n99499, n99500, n99501, n99502, n99503, n99504, n99505,
    n99506, n99507, n99508, n99509, n99510, n99511, n99512, n99513, n99514,
    n99515, n99517, n99518, n99519, n99520, n99521, n99522, n99523, n99524,
    n99525, n99526, n99527, n99528, n99529, n99530, n99531, n99532, n99533,
    n99534, n99535, n99536, n99537, n99538, n99539, n99540, n99541, n99542,
    n99543, n99544, n99545, n99546, n99547, n99548, n99549, n99550, n99551,
    n99552, n99553, n99554, n99555, n99556, n99557, n99558, n99559, n99560,
    n99561, n99562, n99563, n99564, n99565, n99566, n99567, n99568, n99569,
    n99570, n99571, n99572, n99573, n99574, n99575, n99576, n99577, n99578,
    n99579, n99580, n99581, n99582, n99583, n99584, n99585, n99586, n99587,
    n99588, n99589, n99590, n99591, n99592, n99593, n99594, n99595, n99596,
    n99597, n99598, n99599, n99600, n99601, n99602, n99603, n99604, n99605,
    n99606, n99607, n99609, n99610, n99611, n99612, n99613, n99614, n99615,
    n99616, n99617, n99618, n99619, n99620, n99621, n99622, n99623, n99624,
    n99625, n99626, n99627, n99628, n99629, n99630, n99631, n99632, n99633,
    n99634, n99635, n99636, n99637, n99638, n99639, n99640, n99641, n99642,
    n99643, n99644, n99645, n99646, n99647, n99649, n99650, n99651, n99652,
    n99653, n99654, n99655, n99656, n99657, n99658, n99659, n99660, n99661,
    n99662, n99663, n99664, n99665, n99666, n99667, n99668, n99669, n99670,
    n99671, n99672, n99673, n99674, n99675, n99676, n99677, n99678, n99679,
    n99680, n99681, n99682, n99683, n99684, n99685, n99686, n99687, n99688,
    n99689, n99690, n99692, n99693, n99694, n99695, n99696, n99697, n99698,
    n99699, n99700, n99701, n99702, n99703, n99704, n99705, n99706, n99707,
    n99708, n99709, n99710, n99711, n99712, n99713, n99714, n99715, n99716,
    n99717, n99718, n99719, n99720, n99721, n99722, n99723, n99724, n99725,
    n99726, n99727, n99728, n99730, n99731, n99732, n99733, n99734, n99735,
    n99736, n99737, n99738, n99739, n99740, n99741, n99742, n99743, n99744,
    n99745, n99746, n99747, n99748, n99749, n99750, n99751, n99752, n99753,
    n99754, n99755, n99756, n99757, n99758, n99759, n99760, n99761, n99762,
    n99763, n99764, n99765, n99766, n99767, n99768, n99769, n99771, n99772,
    n99773, n99774, n99775, n99776, n99777, n99778, n99779, n99780, n99781,
    n99782, n99783, n99784, n99785, n99786, n99787, n99788, n99789, n99790,
    n99791, n99792, n99793, n99794, n99795, n99796, n99797, n99798, n99799,
    n99800, n99801, n99802, n99803, n99804, n99805, n99806, n99807, n99808,
    n99809, n99810, n99811, n99812, n99813, n99814, n99815, n99816, n99817,
    n99818, n99819, n99820, n99821, n99822, n99823, n99824, n99825, n99826,
    n99827, n99828, n99829, n99830, n99831, n99832, n99833, n99834, n99835,
    n99836, n99837, n99838, n99839, n99840, n99841, n99842, n99843, n99844,
    n99845, n99846, n99847, n99848, n99849, n99850, n99851, n99852, n99853,
    n99854, n99855, n99856, n99857, n99858, n99859, n99860, n99861, n99862,
    n99863, n99864, n99865, n99866, n99868, n99869, n99870, n99871, n99872,
    n99873, n99874, n99875, n99876, n99877, n99878, n99879, n99880, n99881,
    n99882, n99883, n99884, n99885, n99886, n99887, n99888, n99889, n99890,
    n99891, n99892, n99893, n99895, n99896, n99897, n99898, n99899, n99900,
    n99901, n99902, n99903, n99904, n99905, n99906, n99907, n99908, n99909,
    n99910, n99911, n99912, n99913, n99914, n99915, n99916, n99917, n99918,
    n99919, n99920, n99921, n99922, n99923, n99924, n99925, n99926, n99927,
    n99928, n99929, n99930, n99931, n99932, n99933, n99934, n99935, n99936,
    n99937, n99938, n99939, n99940, n99942, n99943, n99944, n99945, n99946,
    n99947, n99948, n99949, n99950, n99951, n99952, n99953, n99954, n99955,
    n99956, n99957, n99958, n99959, n99960, n99961, n99962, n99963, n99964,
    n99965, n99966, n99967, n99968, n99969, n99970, n99971, n99972, n99973,
    n99974, n99975, n99977, n99978, n99979, n99980, n99981, n99982, n99983,
    n99984, n99985, n99986, n99987, n99988, n99989, n99990, n99991, n99992,
    n99993, n99994, n99995, n99996, n99997, n99998, n99999, n100000,
    n100001, n100002, n100003, n100004, n100005, n100006, n100007, n100008,
    n100009, n100010, n100011, n100013, n100014, n100015, n100016, n100017,
    n100018, n100019, n100020, n100021, n100022, n100023, n100024, n100025,
    n100026, n100027, n100028, n100029, n100030, n100031, n100032, n100033,
    n100034, n100035, n100036, n100037, n100038, n100039, n100040, n100041,
    n100042, n100043, n100044, n100045, n100046, n100047, n100048, n100049,
    n100050, n100052, n100053, n100054, n100055, n100056, n100057, n100058,
    n100059, n100060, n100061, n100062, n100063, n100064, n100065, n100066,
    n100067, n100068, n100069, n100070, n100071, n100072, n100073, n100074,
    n100075, n100076, n100077, n100078, n100079, n100080, n100081, n100082,
    n100083, n100084, n100086, n100087, n100088, n100089, n100090, n100091,
    n100092, n100093, n100094, n100095, n100096, n100097, n100098, n100099,
    n100100, n100101, n100102, n100103, n100104, n100105, n100106, n100107,
    n100108, n100109, n100110, n100111, n100112, n100113, n100114, n100115,
    n100116, n100117, n100118, n100119, n100120, n100121, n100122, n100123,
    n100124, n100125, n100126, n100127, n100129, n100130, n100131, n100132,
    n100133, n100134, n100135, n100136, n100137, n100138, n100139, n100140,
    n100141, n100142, n100143, n100144, n100145, n100146, n100147, n100148,
    n100149, n100150, n100151, n100152, n100153, n100154, n100155, n100156,
    n100157, n100158, n100159, n100161, n100162, n100163, n100164, n100165,
    n100166, n100167, n100168, n100169, n100170, n100171, n100172, n100173,
    n100174, n100175, n100176, n100177, n100178, n100179, n100180, n100181,
    n100182, n100183, n100184, n100185, n100186, n100187, n100189, n100190,
    n100191, n100192, n100193, n100194, n100195, n100196, n100197, n100198,
    n100199, n100200, n100201, n100202, n100203, n100204, n100205, n100206,
    n100207, n100208, n100209, n100210, n100211, n100212, n100213, n100214,
    n100215, n100216, n100217, n100218, n100219, n100220, n100221, n100222,
    n100223, n100224, n100225, n100226, n100227, n100228, n100230, n100231,
    n100232, n100233, n100234, n100235, n100236, n100237, n100238, n100239,
    n100240, n100241, n100242, n100243, n100244, n100245, n100246, n100247,
    n100248, n100249, n100250, n100251, n100252, n100253, n100254, n100255,
    n100256, n100257, n100258, n100259, n100260, n100261, n100262, n100263,
    n100264, n100266, n100267, n100268, n100269, n100270, n100271, n100272,
    n100273, n100274, n100275, n100276, n100277, n100278, n100279, n100280,
    n100281, n100282, n100283, n100284, n100285, n100286, n100287, n100288,
    n100289, n100290, n100291, n100292, n100294, n100295, n100296, n100297,
    n100298, n100299, n100300, n100301, n100302, n100303, n100304, n100305,
    n100306, n100307, n100308, n100309, n100310, n100311, n100312, n100313,
    n100314, n100315, n100316, n100317, n100318, n100319, n100320, n100321,
    n100322, n100323, n100324, n100325, n100326, n100327, n100328, n100329,
    n100330, n100331, n100332, n100333, n100334, n100336, n100337, n100338,
    n100339, n100340, n100341, n100342, n100343, n100344, n100345, n100346,
    n100347, n100348, n100349, n100350, n100351, n100352, n100353, n100354,
    n100355, n100356, n100357, n100358, n100359, n100360, n100362, n100363,
    n100364, n100365, n100366, n100367, n100368, n100369, n100370, n100371,
    n100372, n100373, n100374, n100375, n100376, n100377, n100378, n100379,
    n100380, n100381, n100382, n100383, n100384, n100385, n100386, n100387,
    n100388, n100389, n100390, n100391, n100392, n100393, n100394, n100396,
    n100397, n100399, n100400, n100402, n100403, n100405, n100406, n100408,
    n100409, n100411, n100412, n100414, n100415, n100417, n100418, n100420,
    n100421, n100423, n100424, n100426, n100427, n100429, n100430, n100432,
    n100433, n100435, n100436, n100438, n100439, n100441, n100442, n100444,
    n100445, n100447, n100448, n100450, n100451, n100453, n100454, n100456,
    n100457, n100459, n100460, n100462, n100463, n100465, n100466, n100468,
    n100469, n100471, n100472, n100474, n100475, n100477, n100478, n100480,
    n100481, n100483, n100484, n100486, n100487, n100489, n100490, n100492,
    n100493, n100495, n100496, n100498, n100499, n100501, n100502, n100504,
    n100505, n100507, n100508, n100510, n100511, n100513, n100514, n100516,
    n100517, n100519, n100520, n100522, n100523, n100525, n100526, n100528,
    n100529, n100531, n100532, n100534, n100535, n100537, n100538, n100540,
    n100541, n100543, n100544, n100546, n100547, n100549, n100550, n100552,
    n100553, n100555, n100556, n100558, n100559, n100561, n100562, n100564,
    n100565, n100567, n100568, n100570, n100571, n100573, n100574, n100576,
    n100577, n100579, n100580, n100582, n100583, n100585, n100586, n100588,
    n100589, n100591, n100592, n100594, n100595, n100597, n100598, n100600,
    n100601, n100603, n100604, n100606, n100607, n100609, n100610, n100612,
    n100613, n100615, n100616, n100618, n100619, n100621, n100622, n100624,
    n100625, n100627, n100628, n100630, n100631, n100633, n100634, n100636,
    n100637, n100639, n100640, n100642, n100643, n100645, n100646, n100648,
    n100649, n100651, n100652, n100654, n100655, n100657, n100658, n100660,
    n100661, n100663, n100664, n100666, n100667, n100669, n100670, n100672,
    n100673, n100675, n100676, n100678, n100679, n100681, n100682, n100684,
    n100685, n100687, n100688, n100690, n100691, n100693, n100694, n100696,
    n100697, n100699, n100700, n100702, n100703, n100705, n100706, n100708,
    n100709, n100711, n100712, n100714, n100715, n100717, n100718, n100720,
    n100721, n100723, n100724, n100726, n100727, n100729, n100730;
  assign n18082 = pi3105 & pi9040;
  assign n18083 = pi3001 & ~pi9040;
  assign n18084 = ~n18082 & ~n18083;
  assign n18085 = ~pi0077 & ~n18084;
  assign n18086 = pi0077 & n18084;
  assign n18087 = ~n18085 & ~n18086;
  assign n18088 = pi2986 & ~pi9040;
  assign n18089 = pi2984 & pi9040;
  assign n18090 = ~n18088 & ~n18089;
  assign n18091 = pi0070 & n18090;
  assign n18092 = ~pi0070 & ~n18090;
  assign n18093 = ~n18091 & ~n18092;
  assign n18094 = pi3008 & ~pi9040;
  assign n18095 = pi2998 & pi9040;
  assign n18096 = ~n18094 & ~n18095;
  assign n18097 = ~pi0066 & n18096;
  assign n18098 = pi0066 & ~n18096;
  assign n18099 = ~n18097 & ~n18098;
  assign n18100 = pi2992 & ~pi9040;
  assign n18101 = pi3003 & pi9040;
  assign n18102 = ~n18100 & ~n18101;
  assign n18103 = ~pi0036 & ~n18102;
  assign n18104 = pi0036 & n18102;
  assign n18105 = ~n18103 & ~n18104;
  assign n18106 = n18099 & ~n18105;
  assign n18107 = n18093 & n18106;
  assign n18108 = pi3010 & pi9040;
  assign n18109 = pi2991 & ~pi9040;
  assign n18110 = ~n18108 & ~n18109;
  assign n18111 = ~pi0067 & ~n18110;
  assign n18112 = pi0067 & n18110;
  assign n18113 = ~n18111 & ~n18112;
  assign n18114 = pi3103 & ~pi9040;
  assign n18115 = pi2982 & pi9040;
  assign n18116 = ~n18114 & ~n18115;
  assign n18117 = ~pi0095 & n18116;
  assign n18118 = pi0095 & ~n18116;
  assign n18119 = ~n18117 & ~n18118;
  assign n18120 = n18113 & n18119;
  assign n18121 = n18107 & n18120;
  assign n18122 = ~n18099 & ~n18113;
  assign n18123 = ~n18093 & n18122;
  assign n18124 = ~n18093 & ~n18113;
  assign n18125 = ~n18105 & n18124;
  assign n18126 = ~n18123 & ~n18125;
  assign n18127 = n18119 & ~n18126;
  assign n18128 = ~n18121 & ~n18127;
  assign n18129 = ~n18087 & ~n18128;
  assign n18130 = ~n18093 & n18105;
  assign n18131 = n18113 & ~n18119;
  assign n18132 = n18130 & n18131;
  assign n18133 = ~n18099 & n18132;
  assign n18134 = ~n18113 & ~n18119;
  assign n18135 = n18093 & n18105;
  assign n18136 = n18134 & n18135;
  assign n18137 = ~n18105 & n18122;
  assign n18138 = ~n18093 & n18137;
  assign n18139 = n18093 & ~n18105;
  assign n18140 = ~n18099 & n18139;
  assign n18141 = ~n18119 & n18140;
  assign n18142 = n18113 & n18141;
  assign n18143 = ~n18138 & ~n18142;
  assign n18144 = ~n18136 & n18143;
  assign n18145 = ~n18133 & n18144;
  assign n18146 = n18099 & ~n18113;
  assign n18147 = n18105 & n18146;
  assign n18148 = n18093 & n18147;
  assign n18149 = n18145 & ~n18148;
  assign n18150 = ~n18087 & ~n18149;
  assign n18151 = ~n18093 & ~n18105;
  assign n18152 = n18099 & n18113;
  assign n18153 = ~n18119 & n18152;
  assign n18154 = n18151 & n18153;
  assign n18155 = n18093 & ~n18099;
  assign n18156 = n18105 & n18155;
  assign n18157 = n18113 & n18156;
  assign n18158 = ~n18137 & ~n18157;
  assign n18159 = n18099 & n18130;
  assign n18160 = n18113 & n18159;
  assign n18161 = n18158 & ~n18160;
  assign n18162 = n18119 & ~n18161;
  assign n18163 = ~n18154 & ~n18162;
  assign n18164 = ~n18150 & n18163;
  assign n18165 = ~n18129 & n18164;
  assign n18166 = n18093 & n18099;
  assign n18167 = n18134 & n18166;
  assign n18168 = ~n18093 & n18113;
  assign n18169 = n18099 & n18168;
  assign n18170 = ~n18099 & n18119;
  assign n18171 = n18093 & n18170;
  assign n18172 = ~n18169 & ~n18171;
  assign n18173 = ~n18159 & n18172;
  assign n18174 = n18107 & ~n18113;
  assign n18175 = n18173 & ~n18174;
  assign n18176 = ~n18119 & n18130;
  assign n18177 = ~n18113 & n18176;
  assign n18178 = n18099 & n18105;
  assign n18179 = n18113 & n18151;
  assign n18180 = ~n18178 & ~n18179;
  assign n18181 = ~n18119 & ~n18180;
  assign n18182 = ~n18177 & ~n18181;
  assign n18183 = n18175 & n18182;
  assign n18184 = n18087 & ~n18183;
  assign n18185 = ~n18167 & ~n18184;
  assign po0068 = n18165 & n18185;
  assign n18187 = ~n18099 & n18151;
  assign n18188 = n18113 & n18187;
  assign n18189 = ~n18099 & n18130;
  assign n18190 = ~n18113 & n18189;
  assign n18191 = ~n18188 & ~n18190;
  assign n18192 = ~n18119 & ~n18191;
  assign n18193 = ~n18099 & n18113;
  assign n18194 = n18105 & n18193;
  assign n18195 = ~n18113 & n18140;
  assign n18196 = ~n18194 & ~n18195;
  assign n18197 = n18093 & n18120;
  assign n18198 = ~n18093 & n18099;
  assign n18199 = n18119 & n18198;
  assign n18200 = ~n18113 & n18199;
  assign n18201 = ~n18093 & ~n18099;
  assign n18202 = ~n18168 & ~n18201;
  assign n18203 = ~n18148 & n18202;
  assign n18204 = ~n18119 & ~n18203;
  assign n18205 = ~n18200 & ~n18204;
  assign n18206 = ~n18197 & n18205;
  assign n18207 = n18196 & n18206;
  assign n18208 = n18087 & ~n18207;
  assign n18209 = ~n18192 & ~n18208;
  assign n18210 = ~n18107 & ~n18156;
  assign n18211 = ~n18119 & ~n18210;
  assign n18212 = ~n18160 & ~n18211;
  assign n18213 = n18113 & n18140;
  assign n18214 = n18212 & ~n18213;
  assign n18215 = ~n18135 & ~n18151;
  assign n18216 = n18099 & ~n18215;
  assign n18217 = ~n18125 & ~n18216;
  assign n18218 = n18119 & ~n18217;
  assign n18219 = n18214 & ~n18218;
  assign n18220 = ~n18087 & ~n18219;
  assign po0070 = n18209 & ~n18220;
  assign n18222 = pi3046 & ~pi9040;
  assign n18223 = pi3001 & pi9040;
  assign n18224 = ~n18222 & ~n18223;
  assign n18225 = pi0036 & n18224;
  assign n18226 = ~pi0036 & ~n18224;
  assign n18227 = ~n18225 & ~n18226;
  assign n18228 = pi2983 & ~pi9040;
  assign n18229 = pi3045 & pi9040;
  assign n18230 = ~n18228 & ~n18229;
  assign n18231 = ~pi0077 & n18230;
  assign n18232 = pi0077 & ~n18230;
  assign n18233 = ~n18231 & ~n18232;
  assign n18234 = pi2991 & pi9040;
  assign n18235 = pi2999 & ~pi9040;
  assign n18236 = ~n18234 & ~n18235;
  assign n18237 = ~pi0088 & n18236;
  assign n18238 = pi0088 & ~n18236;
  assign n18239 = ~n18237 & ~n18238;
  assign n18240 = n18233 & n18239;
  assign n18241 = n18227 & n18240;
  assign n18242 = pi2987 & pi9040;
  assign n18243 = pi2984 & ~pi9040;
  assign n18244 = ~n18242 & ~n18243;
  assign n18245 = pi0091 & n18244;
  assign n18246 = ~pi0091 & ~n18244;
  assign n18247 = ~n18245 & ~n18246;
  assign n18248 = n18233 & ~n18239;
  assign n18249 = ~n18227 & n18248;
  assign n18250 = n18247 & n18249;
  assign n18251 = ~n18227 & ~n18233;
  assign n18252 = n18239 & n18251;
  assign n18253 = ~n18247 & n18252;
  assign n18254 = ~n18250 & ~n18253;
  assign n18255 = ~n18241 & n18254;
  assign n18256 = pi2995 & pi9040;
  assign n18257 = pi3003 & ~pi9040;
  assign n18258 = ~n18256 & ~n18257;
  assign n18259 = ~pi0071 & n18258;
  assign n18260 = pi0071 & ~n18258;
  assign n18261 = ~n18259 & ~n18260;
  assign n18262 = pi3064 & pi9040;
  assign n18263 = pi3000 & ~pi9040;
  assign n18264 = ~n18262 & ~n18263;
  assign n18265 = ~pi0086 & n18264;
  assign n18266 = pi0086 & ~n18264;
  assign n18267 = ~n18265 & ~n18266;
  assign n18268 = n18261 & n18267;
  assign n18269 = ~n18255 & n18268;
  assign n18270 = ~n18227 & n18247;
  assign n18271 = ~n18233 & n18270;
  assign n18272 = ~n18233 & ~n18239;
  assign n18273 = n18247 & n18272;
  assign n18274 = ~n18271 & ~n18273;
  assign n18275 = ~n18261 & ~n18274;
  assign n18276 = n18227 & n18248;
  assign n18277 = ~n18247 & n18276;
  assign n18278 = ~n18275 & ~n18277;
  assign n18279 = ~n18247 & ~n18261;
  assign n18280 = n18248 & n18279;
  assign n18281 = ~n18227 & n18240;
  assign n18282 = ~n18227 & n18272;
  assign n18283 = ~n18281 & ~n18282;
  assign n18284 = ~n18261 & ~n18283;
  assign n18285 = ~n18233 & n18239;
  assign n18286 = ~n18261 & n18285;
  assign n18287 = ~n18247 & n18286;
  assign n18288 = n18227 & n18287;
  assign n18289 = ~n18284 & ~n18288;
  assign n18290 = ~n18280 & n18289;
  assign n18291 = n18278 & n18290;
  assign n18292 = n18267 & ~n18291;
  assign n18293 = ~n18269 & ~n18292;
  assign n18294 = n18247 & n18285;
  assign n18295 = n18227 & n18294;
  assign n18296 = n18227 & n18272;
  assign n18297 = ~n18247 & n18296;
  assign n18298 = ~n18295 & ~n18297;
  assign n18299 = n18261 & ~n18298;
  assign n18300 = n18247 & n18248;
  assign n18301 = ~n18227 & ~n18247;
  assign n18302 = n18239 & n18301;
  assign n18303 = ~n18300 & ~n18302;
  assign n18304 = ~n18261 & ~n18303;
  assign n18305 = n18239 & n18270;
  assign n18306 = ~n18282 & ~n18305;
  assign n18307 = n18261 & ~n18306;
  assign n18308 = ~n18304 & ~n18307;
  assign n18309 = ~n18239 & ~n18247;
  assign n18310 = n18261 & n18309;
  assign n18311 = ~n18227 & n18310;
  assign n18312 = n18241 & ~n18247;
  assign n18313 = ~n18311 & ~n18312;
  assign n18314 = n18247 & n18276;
  assign n18315 = n18298 & ~n18314;
  assign n18316 = n18313 & n18315;
  assign n18317 = n18308 & n18316;
  assign n18318 = ~n18267 & ~n18317;
  assign n18319 = ~n18299 & ~n18318;
  assign po0073 = n18293 & n18319;
  assign n18321 = ~n18106 & ~n18189;
  assign n18322 = n18134 & ~n18321;
  assign n18323 = ~n18107 & ~n18159;
  assign n18324 = ~n18156 & ~n18187;
  assign n18325 = n18323 & n18324;
  assign n18326 = n18113 & ~n18325;
  assign n18327 = ~n18322 & ~n18326;
  assign n18328 = ~n18195 & n18327;
  assign n18329 = n18087 & ~n18328;
  assign n18330 = n18113 & n18189;
  assign n18331 = ~n18113 & n18156;
  assign n18332 = ~n18330 & ~n18331;
  assign n18333 = n18119 & ~n18332;
  assign n18334 = n18113 & n18216;
  assign n18335 = n18119 & ~n18321;
  assign n18336 = ~n18334 & ~n18335;
  assign n18337 = ~n18105 & n18193;
  assign n18338 = ~n18178 & ~n18337;
  assign n18339 = ~n18187 & n18338;
  assign n18340 = ~n18119 & ~n18339;
  assign n18341 = n18336 & ~n18340;
  assign n18342 = ~n18331 & n18341;
  assign n18343 = ~n18087 & ~n18342;
  assign n18344 = ~n18333 & ~n18343;
  assign po0076 = n18329 | ~n18344;
  assign n18346 = pi3042 & pi9040;
  assign n18347 = pi2981 & ~pi9040;
  assign n18348 = ~n18346 & ~n18347;
  assign n18349 = ~pi0087 & n18348;
  assign n18350 = pi0087 & ~n18348;
  assign n18351 = ~n18349 & ~n18350;
  assign n18352 = pi3044 & ~pi9040;
  assign n18353 = pi3004 & pi9040;
  assign n18354 = ~n18352 & ~n18353;
  assign n18355 = ~pi0068 & ~n18354;
  assign n18356 = pi0068 & ~n18352;
  assign n18357 = ~n18353 & n18356;
  assign n18358 = ~n18355 & ~n18357;
  assign n18359 = pi3063 & pi9040;
  assign n18360 = pi3068 & ~pi9040;
  assign n18361 = ~n18359 & ~n18360;
  assign n18362 = ~pi0076 & n18361;
  assign n18363 = pi0076 & ~n18361;
  assign n18364 = ~n18362 & ~n18363;
  assign n18365 = pi2985 & pi9040;
  assign n18366 = pi3006 & ~pi9040;
  assign n18367 = ~n18365 & ~n18366;
  assign n18368 = ~pi0050 & ~n18367;
  assign n18369 = pi0050 & n18367;
  assign n18370 = ~n18368 & ~n18369;
  assign n18371 = n18364 & n18370;
  assign n18372 = n18358 & n18371;
  assign n18373 = n18351 & n18372;
  assign n18374 = ~n18351 & ~n18358;
  assign n18375 = n18364 & n18374;
  assign n18376 = n18351 & ~n18358;
  assign n18377 = ~n18364 & n18376;
  assign n18378 = n18370 & n18377;
  assign n18379 = ~n18375 & ~n18378;
  assign n18380 = ~n18373 & n18379;
  assign n18381 = pi3043 & pi9040;
  assign n18382 = pi3016 & ~pi9040;
  assign n18383 = ~n18381 & ~n18382;
  assign n18384 = pi0069 & n18383;
  assign n18385 = ~pi0069 & ~n18383;
  assign n18386 = ~n18384 & ~n18385;
  assign n18387 = ~n18380 & ~n18386;
  assign n18388 = ~n18351 & ~n18364;
  assign n18389 = n18370 & n18388;
  assign n18390 = n18351 & ~n18364;
  assign n18391 = ~n18370 & n18390;
  assign n18392 = ~n18389 & ~n18391;
  assign n18393 = n18386 & ~n18392;
  assign n18394 = ~n18387 & ~n18393;
  assign n18395 = pi3011 & pi9040;
  assign n18396 = ~pi3033 & ~pi9040;
  assign n18397 = ~n18395 & ~n18396;
  assign n18398 = ~pi0061 & ~n18397;
  assign n18399 = pi0061 & n18397;
  assign n18400 = ~n18398 & ~n18399;
  assign n18401 = n18351 & n18358;
  assign n18402 = ~n18364 & n18401;
  assign n18403 = n18364 & ~n18370;
  assign n18404 = n18358 & n18403;
  assign n18405 = ~n18351 & n18404;
  assign n18406 = ~n18402 & ~n18405;
  assign n18407 = n18386 & ~n18406;
  assign n18408 = n18364 & n18376;
  assign n18409 = ~n18370 & n18408;
  assign n18410 = ~n18373 & ~n18409;
  assign n18411 = ~n18351 & n18364;
  assign n18412 = n18370 & n18411;
  assign n18413 = ~n18351 & n18358;
  assign n18414 = ~n18364 & n18413;
  assign n18415 = ~n18370 & n18414;
  assign n18416 = ~n18412 & ~n18415;
  assign n18417 = ~n18386 & ~n18416;
  assign n18418 = n18410 & ~n18417;
  assign n18419 = ~n18407 & n18418;
  assign n18420 = n18400 & ~n18419;
  assign n18421 = ~n18358 & n18364;
  assign n18422 = ~n18386 & n18421;
  assign n18423 = ~n18370 & n18422;
  assign n18424 = n18386 & n18401;
  assign n18425 = ~n18370 & n18424;
  assign n18426 = n18370 & n18408;
  assign n18427 = ~n18364 & n18374;
  assign n18428 = ~n18426 & ~n18427;
  assign n18429 = n18370 & n18413;
  assign n18430 = n18428 & ~n18429;
  assign n18431 = n18386 & ~n18430;
  assign n18432 = ~n18370 & n18375;
  assign n18433 = ~n18370 & ~n18386;
  assign n18434 = n18411 & n18433;
  assign n18435 = ~n18432 & ~n18434;
  assign n18436 = ~n18431 & n18435;
  assign n18437 = ~n18425 & n18436;
  assign n18438 = ~n18370 & n18402;
  assign n18439 = n18370 & n18414;
  assign n18440 = ~n18438 & ~n18439;
  assign n18441 = n18437 & n18440;
  assign n18442 = ~n18400 & ~n18441;
  assign n18443 = ~n18423 & ~n18442;
  assign n18444 = ~n18420 & n18443;
  assign po0079 = n18394 & n18444;
  assign n18446 = ~n18247 & n18282;
  assign n18447 = n18240 & ~n18247;
  assign n18448 = ~n18276 & ~n18447;
  assign n18449 = n18261 & ~n18448;
  assign n18450 = ~n18446 & ~n18449;
  assign n18451 = ~n18250 & n18450;
  assign n18452 = ~n18233 & n18279;
  assign n18453 = n18241 & n18247;
  assign n18454 = ~n18296 & ~n18453;
  assign n18455 = ~n18252 & n18454;
  assign n18456 = ~n18261 & ~n18455;
  assign n18457 = ~n18452 & ~n18456;
  assign n18458 = n18451 & n18457;
  assign n18459 = ~n18267 & ~n18458;
  assign n18460 = n18233 & n18270;
  assign n18461 = ~n18295 & ~n18460;
  assign n18462 = n18261 & ~n18461;
  assign n18463 = n18247 & ~n18283;
  assign n18464 = ~n18295 & ~n18463;
  assign n18465 = n18267 & ~n18464;
  assign n18466 = ~n18261 & n18267;
  assign n18467 = ~n18448 & n18466;
  assign n18468 = ~n18465 & ~n18467;
  assign n18469 = n18227 & ~n18233;
  assign n18470 = ~n18247 & n18285;
  assign n18471 = ~n18469 & ~n18470;
  assign n18472 = ~n18249 & n18471;
  assign n18473 = n18268 & ~n18472;
  assign n18474 = n18468 & ~n18473;
  assign n18475 = ~n18462 & n18474;
  assign po0082 = n18459 | ~n18475;
  assign n18477 = n18106 & ~n18113;
  assign n18478 = n18113 & n18135;
  assign n18479 = ~n18155 & ~n18478;
  assign n18480 = n18119 & ~n18479;
  assign n18481 = ~n18119 & n18187;
  assign n18482 = n18113 & n18176;
  assign n18483 = ~n18194 & ~n18482;
  assign n18484 = ~n18481 & n18483;
  assign n18485 = ~n18480 & n18484;
  assign n18486 = ~n18477 & n18485;
  assign n18487 = ~n18087 & ~n18486;
  assign n18488 = n18087 & n18119;
  assign n18489 = n18107 & n18113;
  assign n18490 = ~n18159 & ~n18489;
  assign n18491 = ~n18187 & n18490;
  assign n18492 = n18488 & ~n18491;
  assign n18493 = ~n18119 & n18189;
  assign n18494 = ~n18154 & ~n18493;
  assign n18495 = ~n18148 & n18494;
  assign n18496 = ~n18142 & n18495;
  assign n18497 = n18087 & ~n18496;
  assign n18498 = ~n18492 & ~n18497;
  assign n18499 = n18120 & n18156;
  assign n18500 = ~n18113 & n18159;
  assign n18501 = ~n18195 & ~n18500;
  assign n18502 = n18119 & ~n18501;
  assign n18503 = ~n18499 & ~n18502;
  assign n18504 = ~n18167 & n18503;
  assign n18505 = ~n18113 & n18481;
  assign n18506 = n18504 & ~n18505;
  assign n18507 = n18498 & n18506;
  assign po0085 = n18487 | ~n18507;
  assign n18509 = pi2980 & pi9040;
  assign n18510 = pi3066 & ~pi9040;
  assign n18511 = ~n18509 & ~n18510;
  assign n18512 = ~pi0058 & n18511;
  assign n18513 = pi0058 & ~n18511;
  assign n18514 = ~n18512 & ~n18513;
  assign n18515 = pi3106 & ~pi9040;
  assign n18516 = pi3068 & pi9040;
  assign n18517 = ~n18515 & ~n18516;
  assign n18518 = ~pi0076 & ~n18517;
  assign n18519 = pi0076 & n18517;
  assign n18520 = ~n18518 & ~n18519;
  assign n18521 = ~n18514 & n18520;
  assign n18522 = pi2997 & pi9040;
  assign n18523 = pi3047 & ~pi9040;
  assign n18524 = ~n18522 & ~n18523;
  assign n18525 = pi0064 & n18524;
  assign n18526 = ~pi0064 & ~n18524;
  assign n18527 = ~n18525 & ~n18526;
  assign n18528 = ~pi3042 & ~pi9040;
  assign n18529 = ~pi3009 & pi9040;
  assign n18530 = ~n18528 & ~n18529;
  assign n18531 = ~pi0090 & n18530;
  assign n18532 = pi0090 & ~n18530;
  assign n18533 = ~n18531 & ~n18532;
  assign n18534 = ~n18527 & ~n18533;
  assign n18535 = n18521 & n18534;
  assign n18536 = pi2990 & pi9040;
  assign n18537 = pi2985 & ~pi9040;
  assign n18538 = ~n18536 & ~n18537;
  assign n18539 = ~pi0060 & n18538;
  assign n18540 = pi0060 & ~n18538;
  assign n18541 = ~n18539 & ~n18540;
  assign n18542 = ~n18514 & n18541;
  assign n18543 = n18520 & n18542;
  assign n18544 = n18527 & n18543;
  assign n18545 = ~n18514 & ~n18520;
  assign n18546 = ~n18541 & n18545;
  assign n18547 = ~n18544 & ~n18546;
  assign n18548 = n18514 & n18520;
  assign n18549 = ~n18527 & n18548;
  assign n18550 = n18547 & ~n18549;
  assign n18551 = n18533 & ~n18550;
  assign n18552 = n18541 & n18548;
  assign n18553 = n18527 & n18552;
  assign n18554 = n18514 & ~n18520;
  assign n18555 = ~n18541 & n18554;
  assign n18556 = ~n18553 & ~n18555;
  assign n18557 = ~n18533 & ~n18556;
  assign n18558 = ~n18527 & n18541;
  assign n18559 = ~n18520 & n18558;
  assign n18560 = ~n18514 & n18559;
  assign n18561 = ~n18557 & ~n18560;
  assign n18562 = ~n18551 & n18561;
  assign n18563 = ~n18535 & n18562;
  assign n18564 = ~pi3033 & pi9040;
  assign n18565 = pi2979 & ~pi9040;
  assign n18566 = ~n18564 & ~n18565;
  assign n18567 = ~pi0087 & n18566;
  assign n18568 = pi0087 & ~n18566;
  assign n18569 = ~n18567 & ~n18568;
  assign n18570 = ~n18563 & n18569;
  assign n18571 = n18520 & n18527;
  assign n18572 = ~n18541 & n18571;
  assign n18573 = n18514 & ~n18527;
  assign n18574 = ~n18527 & ~n18541;
  assign n18575 = ~n18520 & n18574;
  assign n18576 = ~n18573 & ~n18575;
  assign n18577 = ~n18533 & ~n18576;
  assign n18578 = ~n18527 & n18533;
  assign n18579 = n18521 & n18578;
  assign n18580 = ~n18527 & n18555;
  assign n18581 = ~n18579 & ~n18580;
  assign n18582 = ~n18577 & n18581;
  assign n18583 = ~n18572 & n18582;
  assign n18584 = ~n18569 & ~n18583;
  assign n18585 = ~n18570 & ~n18584;
  assign n18586 = n18541 & n18545;
  assign n18587 = n18521 & ~n18541;
  assign n18588 = ~n18586 & ~n18587;
  assign n18589 = n18527 & n18588;
  assign n18590 = ~n18527 & ~n18554;
  assign n18591 = ~n18589 & ~n18590;
  assign n18592 = ~n18533 & n18591;
  assign n18593 = n18527 & n18533;
  assign n18594 = ~n18541 & n18548;
  assign n18595 = n18541 & n18554;
  assign n18596 = ~n18546 & ~n18595;
  assign n18597 = ~n18594 & n18596;
  assign n18598 = n18593 & ~n18597;
  assign n18599 = ~n18592 & ~n18598;
  assign po0088 = n18585 & n18599;
  assign n18601 = pi3000 & pi9040;
  assign n18602 = pi3038 & ~pi9040;
  assign n18603 = ~n18601 & ~n18602;
  assign n18604 = pi0059 & n18603;
  assign n18605 = ~pi0059 & ~n18603;
  assign n18606 = ~n18604 & ~n18605;
  assign n18607 = pi3046 & pi9040;
  assign n18608 = pi2996 & ~pi9040;
  assign n18609 = ~n18607 & ~n18608;
  assign n18610 = pi0089 & n18609;
  assign n18611 = ~pi0089 & ~n18609;
  assign n18612 = ~n18610 & ~n18611;
  assign n18613 = pi3040 & pi9040;
  assign n18614 = pi2995 & ~pi9040;
  assign n18615 = ~n18613 & ~n18614;
  assign n18616 = pi0084 & n18615;
  assign n18617 = ~pi0084 & ~n18615;
  assign n18618 = ~n18616 & ~n18617;
  assign n18619 = pi2987 & ~pi9040;
  assign n18620 = pi3008 & pi9040;
  assign n18621 = ~n18619 & ~n18620;
  assign n18622 = ~pi0049 & n18621;
  assign n18623 = pi0049 & ~n18621;
  assign n18624 = ~n18622 & ~n18623;
  assign n18625 = pi2983 & pi9040;
  assign n18626 = pi3105 & ~pi9040;
  assign n18627 = ~n18625 & ~n18626;
  assign n18628 = pi0083 & n18627;
  assign n18629 = ~pi0083 & ~n18627;
  assign n18630 = ~n18628 & ~n18629;
  assign n18631 = n18624 & ~n18630;
  assign n18632 = ~n18618 & n18631;
  assign n18633 = ~n18612 & n18632;
  assign n18634 = n18612 & ~n18618;
  assign n18635 = ~n18630 & n18634;
  assign n18636 = ~n18624 & n18635;
  assign n18637 = ~n18633 & ~n18636;
  assign n18638 = n18606 & ~n18637;
  assign n18639 = pi2978 & ~pi9040;
  assign n18640 = pi2986 & pi9040;
  assign n18641 = ~n18639 & ~n18640;
  assign n18642 = ~pi0092 & ~n18641;
  assign n18643 = pi0092 & n18641;
  assign n18644 = ~n18642 & ~n18643;
  assign n18645 = n18624 & n18630;
  assign n18646 = n18618 & n18645;
  assign n18647 = ~n18612 & n18646;
  assign n18648 = ~n18624 & ~n18630;
  assign n18649 = n18618 & n18648;
  assign n18650 = n18606 & n18649;
  assign n18651 = ~n18647 & ~n18650;
  assign n18652 = n18612 & n18618;
  assign n18653 = n18630 & n18652;
  assign n18654 = ~n18624 & n18653;
  assign n18655 = ~n18606 & n18612;
  assign n18656 = n18631 & n18655;
  assign n18657 = ~n18618 & n18656;
  assign n18658 = ~n18612 & ~n18618;
  assign n18659 = ~n18624 & n18658;
  assign n18660 = ~n18612 & n18618;
  assign n18661 = n18624 & n18660;
  assign n18662 = ~n18659 & ~n18661;
  assign n18663 = ~n18606 & ~n18662;
  assign n18664 = n18606 & ~n18618;
  assign n18665 = n18630 & n18664;
  assign n18666 = n18624 & n18665;
  assign n18667 = ~n18663 & ~n18666;
  assign n18668 = ~n18657 & n18667;
  assign n18669 = ~n18654 & n18668;
  assign n18670 = n18651 & n18669;
  assign n18671 = n18644 & ~n18670;
  assign n18672 = ~n18606 & n18647;
  assign n18673 = ~n18612 & n18650;
  assign n18674 = ~n18672 & ~n18673;
  assign n18675 = ~n18671 & n18674;
  assign n18676 = ~n18638 & n18675;
  assign n18677 = n18618 & n18631;
  assign n18678 = n18612 & n18677;
  assign n18679 = ~n18633 & ~n18678;
  assign n18680 = n18606 & n18612;
  assign n18681 = n18618 & n18624;
  assign n18682 = n18680 & n18681;
  assign n18683 = n18606 & n18632;
  assign n18684 = n18612 & n18648;
  assign n18685 = ~n18618 & n18630;
  assign n18686 = ~n18684 & ~n18685;
  assign n18687 = ~n18606 & ~n18686;
  assign n18688 = ~n18624 & n18630;
  assign n18689 = ~n18618 & n18688;
  assign n18690 = ~n18612 & n18689;
  assign n18691 = n18618 & n18688;
  assign n18692 = n18606 & n18691;
  assign n18693 = ~n18690 & ~n18692;
  assign n18694 = ~n18687 & n18693;
  assign n18695 = ~n18683 & n18694;
  assign n18696 = ~n18682 & n18695;
  assign n18697 = n18679 & n18696;
  assign n18698 = ~n18644 & ~n18697;
  assign po0091 = n18676 & ~n18698;
  assign n18700 = pi2980 & ~pi9040;
  assign n18701 = pi2988 & pi9040;
  assign n18702 = ~n18700 & ~n18701;
  assign n18703 = pi0094 & n18702;
  assign n18704 = ~pi0094 & ~n18702;
  assign n18705 = ~n18703 & ~n18704;
  assign n18706 = pi3028 & ~pi9040;
  assign n18707 = pi2976 & pi9040;
  assign n18708 = ~n18706 & ~n18707;
  assign n18709 = ~pi0085 & ~n18708;
  assign n18710 = pi0085 & n18708;
  assign n18711 = ~n18709 & ~n18710;
  assign n18712 = pi3044 & pi9040;
  assign n18713 = pi2997 & ~pi9040;
  assign n18714 = ~n18712 & ~n18713;
  assign n18715 = ~pi0083 & ~n18714;
  assign n18716 = pi0083 & n18714;
  assign n18717 = ~n18715 & ~n18716;
  assign n18718 = pi2993 & pi9040;
  assign n18719 = pi2990 & ~pi9040;
  assign n18720 = ~n18718 & ~n18719;
  assign n18721 = ~pi0092 & n18720;
  assign n18722 = pi0092 & ~n18720;
  assign n18723 = ~n18721 & ~n18722;
  assign n18724 = pi3016 & pi9040;
  assign n18725 = pi3058 & ~pi9040;
  assign n18726 = ~n18724 & ~n18725;
  assign n18727 = ~pi0060 & ~n18726;
  assign n18728 = pi0060 & n18726;
  assign n18729 = ~n18727 & ~n18728;
  assign n18730 = n18723 & ~n18729;
  assign n18731 = ~n18717 & n18730;
  assign n18732 = ~n18711 & n18731;
  assign n18733 = n18723 & n18729;
  assign n18734 = n18717 & n18733;
  assign n18735 = ~n18711 & n18734;
  assign n18736 = ~n18732 & ~n18735;
  assign n18737 = ~n18705 & ~n18736;
  assign n18738 = ~n18723 & n18729;
  assign n18739 = n18717 & n18738;
  assign n18740 = ~n18711 & n18739;
  assign n18741 = n18705 & n18740;
  assign n18742 = ~n18737 & ~n18741;
  assign n18743 = ~n18717 & n18733;
  assign n18744 = n18705 & n18733;
  assign n18745 = ~n18705 & n18738;
  assign n18746 = ~n18744 & ~n18745;
  assign n18747 = n18717 & ~n18729;
  assign n18748 = ~n18723 & n18747;
  assign n18749 = n18746 & ~n18748;
  assign n18750 = ~n18743 & n18749;
  assign n18751 = n18711 & ~n18750;
  assign n18752 = ~n18717 & n18738;
  assign n18753 = ~n18705 & n18752;
  assign n18754 = ~n18751 & ~n18753;
  assign n18755 = ~n18705 & n18748;
  assign n18756 = ~n18723 & ~n18729;
  assign n18757 = ~n18717 & n18756;
  assign n18758 = n18705 & n18757;
  assign n18759 = ~n18755 & ~n18758;
  assign n18760 = n18754 & n18759;
  assign n18761 = n18742 & n18760;
  assign n18762 = pi2994 & ~pi9040;
  assign n18763 = pi3106 & pi9040;
  assign n18764 = ~n18762 & ~n18763;
  assign n18765 = ~pi0058 & ~n18764;
  assign n18766 = pi0058 & n18764;
  assign n18767 = ~n18765 & ~n18766;
  assign n18768 = ~n18761 & n18767;
  assign n18769 = n18717 & n18730;
  assign n18770 = n18705 & n18769;
  assign n18771 = n18705 & n18743;
  assign n18772 = ~n18770 & ~n18771;
  assign n18773 = ~n18711 & ~n18772;
  assign n18774 = ~n18768 & ~n18773;
  assign n18775 = ~n18705 & n18769;
  assign n18776 = n18705 & n18747;
  assign n18777 = ~n18705 & n18757;
  assign n18778 = ~n18776 & ~n18777;
  assign n18779 = ~n18705 & n18717;
  assign n18780 = n18729 & n18779;
  assign n18781 = ~n18723 & n18780;
  assign n18782 = n18778 & ~n18781;
  assign n18783 = ~n18743 & n18782;
  assign n18784 = ~n18711 & ~n18783;
  assign n18785 = n18723 & n18779;
  assign n18786 = n18705 & n18738;
  assign n18787 = ~n18785 & ~n18786;
  assign n18788 = ~n18731 & n18787;
  assign n18789 = n18711 & ~n18788;
  assign n18790 = n18705 & n18752;
  assign n18791 = ~n18789 & ~n18790;
  assign n18792 = ~n18784 & n18791;
  assign n18793 = ~n18775 & n18792;
  assign n18794 = ~n18767 & ~n18793;
  assign n18795 = n18705 & n18731;
  assign n18796 = ~n18755 & ~n18795;
  assign n18797 = n18711 & ~n18796;
  assign n18798 = ~n18794 & ~n18797;
  assign po0094 = n18774 & n18798;
  assign n18800 = n18520 & ~n18541;
  assign n18801 = n18578 & n18800;
  assign n18802 = ~n18521 & ~n18554;
  assign n18803 = n18527 & ~n18802;
  assign n18804 = ~n18595 & ~n18803;
  assign n18805 = ~n18533 & ~n18804;
  assign n18806 = n18514 & ~n18541;
  assign n18807 = ~n18527 & n18806;
  assign n18808 = ~n18594 & ~n18807;
  assign n18809 = n18527 & n18546;
  assign n18810 = n18808 & ~n18809;
  assign n18811 = n18533 & ~n18810;
  assign n18812 = ~n18805 & ~n18811;
  assign n18813 = ~n18533 & n18545;
  assign n18814 = ~n18527 & n18813;
  assign n18815 = n18527 & n18595;
  assign n18816 = ~n18544 & ~n18815;
  assign n18817 = ~n18527 & n18552;
  assign n18818 = n18816 & ~n18817;
  assign n18819 = ~n18814 & n18818;
  assign n18820 = n18812 & n18819;
  assign n18821 = ~n18569 & ~n18820;
  assign n18822 = ~n18520 & ~n18527;
  assign n18823 = n18541 & n18822;
  assign n18824 = n18527 & n18555;
  assign n18825 = ~n18823 & ~n18824;
  assign n18826 = n18588 & n18825;
  assign n18827 = n18533 & ~n18826;
  assign n18828 = ~n18553 & ~n18827;
  assign n18829 = n18569 & ~n18828;
  assign n18830 = ~n18533 & n18569;
  assign n18831 = n18521 & ~n18527;
  assign n18832 = ~n18809 & ~n18831;
  assign n18833 = ~n18807 & n18832;
  assign n18834 = n18830 & ~n18833;
  assign n18835 = ~n18829 & ~n18834;
  assign n18836 = ~n18821 & n18835;
  assign n18837 = ~n18560 & n18836;
  assign po0097 = n18801 | ~n18837;
  assign n18839 = n18527 & n18587;
  assign n18840 = ~n18533 & n18594;
  assign n18841 = ~n18839 & ~n18840;
  assign n18842 = ~n18514 & n18527;
  assign n18843 = ~n18542 & ~n18842;
  assign n18844 = ~n18555 & n18843;
  assign n18845 = n18533 & ~n18844;
  assign n18846 = n18841 & ~n18845;
  assign n18847 = ~n18533 & n18595;
  assign n18848 = n18846 & ~n18847;
  assign n18849 = n18569 & ~n18848;
  assign n18850 = n18533 & n18552;
  assign n18851 = ~n18575 & ~n18817;
  assign n18852 = ~n18514 & n18574;
  assign n18853 = n18533 & n18852;
  assign n18854 = n18527 & n18800;
  assign n18855 = n18514 & n18854;
  assign n18856 = ~n18533 & n18542;
  assign n18857 = ~n18815 & ~n18856;
  assign n18858 = ~n18855 & n18857;
  assign n18859 = ~n18853 & n18858;
  assign n18860 = n18851 & n18859;
  assign n18861 = ~n18850 & n18860;
  assign n18862 = ~n18569 & ~n18861;
  assign n18863 = n18533 & n18817;
  assign n18864 = ~n18527 & n18546;
  assign n18865 = ~n18533 & n18864;
  assign n18866 = ~n18863 & ~n18865;
  assign n18867 = ~n18527 & n18543;
  assign n18868 = ~n18533 & n18867;
  assign n18869 = n18866 & ~n18868;
  assign n18870 = ~n18862 & n18869;
  assign po0100 = n18849 | ~n18870;
  assign n18872 = n18705 & ~n18717;
  assign n18873 = ~n18711 & n18872;
  assign n18874 = ~n18723 & n18873;
  assign n18875 = n18711 & n18747;
  assign n18876 = ~n18705 & n18875;
  assign n18877 = n18705 & n18734;
  assign n18878 = ~n18876 & ~n18877;
  assign n18879 = n18717 & n18723;
  assign n18880 = n18705 & n18879;
  assign n18881 = ~n18757 & ~n18880;
  assign n18882 = ~n18711 & ~n18881;
  assign n18883 = ~n18717 & n18723;
  assign n18884 = ~n18711 & n18883;
  assign n18885 = ~n18705 & n18884;
  assign n18886 = ~n18882 & ~n18885;
  assign n18887 = n18878 & n18886;
  assign n18888 = ~n18767 & ~n18887;
  assign n18889 = ~n18705 & n18743;
  assign n18890 = n18705 & ~n18723;
  assign n18891 = n18717 & n18890;
  assign n18892 = ~n18729 & n18891;
  assign n18893 = ~n18795 & ~n18892;
  assign n18894 = ~n18889 & n18893;
  assign n18895 = n18711 & ~n18894;
  assign n18896 = ~n18752 & ~n18785;
  assign n18897 = ~n18711 & ~n18896;
  assign n18898 = ~n18780 & ~n18897;
  assign n18899 = ~n18705 & ~n18717;
  assign n18900 = ~n18729 & n18899;
  assign n18901 = n18705 & n18730;
  assign n18902 = ~n18900 & ~n18901;
  assign n18903 = ~n18883 & n18902;
  assign n18904 = ~n18739 & n18903;
  assign n18905 = n18711 & ~n18904;
  assign n18906 = n18898 & ~n18905;
  assign n18907 = ~n18892 & n18906;
  assign n18908 = n18767 & ~n18907;
  assign n18909 = ~n18895 & ~n18908;
  assign n18910 = ~n18888 & n18909;
  assign n18911 = ~n18781 & n18910;
  assign po0103 = n18874 | ~n18911;
  assign n18913 = ~n18261 & n18469;
  assign n18914 = ~n18247 & n18913;
  assign n18915 = n18247 & n18281;
  assign n18916 = ~n18261 & n18915;
  assign n18917 = n18247 & n18469;
  assign n18918 = ~n18294 & ~n18917;
  assign n18919 = ~n18249 & n18918;
  assign n18920 = n18261 & ~n18919;
  assign n18921 = n18227 & n18239;
  assign n18922 = ~n18249 & ~n18921;
  assign n18923 = ~n18247 & ~n18922;
  assign n18924 = n18247 & ~n18261;
  assign n18925 = n18282 & n18924;
  assign n18926 = ~n18923 & ~n18925;
  assign n18927 = ~n18311 & n18926;
  assign n18928 = ~n18920 & n18927;
  assign n18929 = ~n18314 & n18928;
  assign n18930 = n18267 & ~n18929;
  assign n18931 = ~n18247 & n18249;
  assign n18932 = ~n18314 & ~n18931;
  assign n18933 = n18261 & ~n18932;
  assign n18934 = n18247 & n18261;
  assign n18935 = ~n18240 & ~n18282;
  assign n18936 = n18934 & ~n18935;
  assign n18937 = n18240 & n18261;
  assign n18938 = ~n18227 & n18937;
  assign n18939 = ~n18936 & ~n18938;
  assign n18940 = n18227 & n18279;
  assign n18941 = ~n18913 & ~n18940;
  assign n18942 = n18939 & n18941;
  assign n18943 = ~n18253 & n18942;
  assign n18944 = ~n18297 & n18943;
  assign n18945 = ~n18267 & ~n18944;
  assign n18946 = ~n18933 & ~n18945;
  assign n18947 = ~n18930 & n18946;
  assign n18948 = ~n18916 & n18947;
  assign po0106 = n18914 | ~n18948;
  assign n18950 = ~n18618 & n18645;
  assign n18951 = n18612 & n18950;
  assign n18952 = ~n18678 & ~n18951;
  assign n18953 = ~n18654 & n18952;
  assign n18954 = n18606 & ~n18953;
  assign n18955 = ~n18612 & n18649;
  assign n18956 = ~n18612 & n18631;
  assign n18957 = ~n18636 & ~n18956;
  assign n18958 = n18606 & ~n18957;
  assign n18959 = ~n18647 & ~n18654;
  assign n18960 = ~n18612 & n18648;
  assign n18961 = ~n18689 & ~n18960;
  assign n18962 = ~n18606 & ~n18961;
  assign n18963 = n18959 & ~n18962;
  assign n18964 = ~n18958 & n18963;
  assign n18965 = ~n18955 & n18964;
  assign n18966 = ~n18644 & ~n18965;
  assign n18967 = n18624 & n18634;
  assign n18968 = n18612 & n18649;
  assign n18969 = ~n18967 & ~n18968;
  assign n18970 = n18644 & ~n18969;
  assign n18971 = n18630 & n18660;
  assign n18972 = ~n18661 & ~n18971;
  assign n18973 = ~n18646 & n18972;
  assign n18974 = ~n18606 & ~n18973;
  assign n18975 = n18644 & n18974;
  assign n18976 = ~n18970 & ~n18975;
  assign n18977 = n18649 & n18655;
  assign n18978 = ~n18657 & ~n18977;
  assign n18979 = ~n18659 & ~n18685;
  assign n18980 = n18606 & ~n18979;
  assign n18981 = n18644 & n18980;
  assign n18982 = n18978 & ~n18981;
  assign n18983 = n18976 & n18982;
  assign n18984 = ~n18966 & n18983;
  assign po0109 = n18954 | ~n18984;
  assign n18986 = ~n18527 & n18847;
  assign n18987 = n18521 & n18527;
  assign n18988 = ~n18580 & ~n18987;
  assign n18989 = n18533 & ~n18988;
  assign n18990 = ~n18863 & ~n18989;
  assign n18991 = n18527 & n18806;
  assign n18992 = ~n18587 & ~n18991;
  assign n18993 = ~n18560 & n18992;
  assign n18994 = n18533 & ~n18993;
  assign n18995 = ~n18527 & n18594;
  assign n18996 = n18514 & n18541;
  assign n18997 = ~n18545 & ~n18996;
  assign n18998 = n18527 & ~n18997;
  assign n18999 = ~n18995 & ~n18998;
  assign n19000 = ~n18867 & n18999;
  assign n19001 = ~n18533 & ~n19000;
  assign n19002 = ~n18994 & ~n19001;
  assign n19003 = ~n18569 & ~n19002;
  assign n19004 = ~n18865 & ~n19003;
  assign n19005 = n18514 & n18578;
  assign n19006 = ~n18852 & ~n18991;
  assign n19007 = ~n18533 & ~n19006;
  assign n19008 = ~n18814 & ~n19007;
  assign n19009 = ~n18544 & ~n18864;
  assign n19010 = n18542 & n18593;
  assign n19011 = ~n18850 & ~n19010;
  assign n19012 = n19009 & n19011;
  assign n19013 = n19008 & n19012;
  assign n19014 = ~n19005 & n19013;
  assign n19015 = n18569 & ~n19014;
  assign n19016 = n19004 & ~n19015;
  assign n19017 = n18990 & n19016;
  assign po0112 = n18986 | ~n19017;
  assign n19019 = ~n18370 & n18377;
  assign n19020 = ~n18432 & ~n19019;
  assign n19021 = ~n18351 & n18372;
  assign n19022 = n18370 & n18402;
  assign n19023 = n18364 & n18401;
  assign n19024 = ~n18386 & n19023;
  assign n19025 = ~n19022 & ~n19024;
  assign n19026 = ~n18426 & n19025;
  assign n19027 = ~n19021 & n19026;
  assign n19028 = n18358 & ~n18364;
  assign n19029 = ~n18351 & n18370;
  assign n19030 = ~n18421 & ~n19029;
  assign n19031 = ~n19028 & n19030;
  assign n19032 = n18386 & ~n19031;
  assign n19033 = n19027 & ~n19032;
  assign n19034 = n19020 & n19033;
  assign n19035 = ~n18400 & ~n19034;
  assign n19036 = n18370 & n18375;
  assign n19037 = ~n18388 & ~n18409;
  assign n19038 = ~n18386 & ~n19037;
  assign n19039 = ~n19036 & ~n19038;
  assign n19040 = ~n18405 & n19039;
  assign n19041 = n18373 & n18386;
  assign n19042 = ~n18438 & ~n19041;
  assign n19043 = ~n18378 & n19042;
  assign n19044 = n19040 & n19043;
  assign n19045 = n18400 & ~n19044;
  assign po0115 = ~n19035 & ~n19045;
  assign n19047 = ~n18711 & n18758;
  assign n19048 = n18711 & n18739;
  assign n19049 = ~n18705 & n18733;
  assign n19050 = ~n18734 & ~n19049;
  assign n19051 = ~n18752 & n19050;
  assign n19052 = ~n18711 & ~n19051;
  assign n19053 = ~n18705 & n18711;
  assign n19054 = n18757 & n19053;
  assign n19055 = ~n18785 & ~n19054;
  assign n19056 = n18893 & n19055;
  assign n19057 = ~n19052 & n19056;
  assign n19058 = ~n19048 & n19057;
  assign n19059 = ~n18767 & ~n19058;
  assign n19060 = ~n18705 & ~n18723;
  assign n19061 = ~n18711 & n19060;
  assign n19062 = ~n18705 & n18731;
  assign n19063 = ~n18752 & ~n19062;
  assign n19064 = n18711 & ~n19063;
  assign n19065 = ~n19061 & ~n19064;
  assign n19066 = n18772 & n19065;
  assign n19067 = n18767 & ~n19066;
  assign n19068 = n18734 & n19053;
  assign n19069 = n18705 & n18875;
  assign n19070 = ~n19068 & ~n19069;
  assign n19071 = n18711 & n18771;
  assign n19072 = n19070 & ~n19071;
  assign n19073 = ~n19067 & n19072;
  assign n19074 = ~n19059 & n19073;
  assign po0118 = n19047 | ~n19074;
  assign n19076 = ~n18673 & ~n18682;
  assign n19077 = ~n18618 & n18648;
  assign n19078 = ~n18647 & ~n19077;
  assign n19079 = ~n18684 & n19078;
  assign n19080 = ~n18606 & ~n19079;
  assign n19081 = ~n18654 & ~n18951;
  assign n19082 = n18606 & ~n18612;
  assign n19083 = n18689 & n19082;
  assign n19084 = n19081 & ~n19083;
  assign n19085 = n18606 & n18677;
  assign n19086 = n19084 & ~n19085;
  assign n19087 = ~n19080 & n19086;
  assign n19088 = n18644 & ~n19087;
  assign n19089 = n18606 & n18645;
  assign n19090 = ~n18612 & n19089;
  assign n19091 = ~n18624 & n18634;
  assign n19092 = ~n19077 & ~n19091;
  assign n19093 = n18606 & ~n19092;
  assign n19094 = ~n19090 & ~n19093;
  assign n19095 = ~n18606 & ~n18612;
  assign n19096 = n18688 & n19095;
  assign n19097 = ~n18606 & n18632;
  assign n19098 = ~n19096 & ~n19097;
  assign n19099 = n19094 & n19098;
  assign n19100 = ~n18624 & n18660;
  assign n19101 = ~n18633 & ~n19100;
  assign n19102 = ~n18678 & n19101;
  assign n19103 = n19099 & n19102;
  assign n19104 = ~n18644 & ~n19103;
  assign n19105 = ~n18633 & n19081;
  assign n19106 = ~n18606 & ~n19105;
  assign n19107 = ~n19104 & ~n19106;
  assign n19108 = ~n19088 & n19107;
  assign po0121 = ~n19076 | ~n19108;
  assign n19110 = pi3043 & ~pi9040;
  assign n19111 = pi3066 & pi9040;
  assign n19112 = ~n19110 & ~n19111;
  assign n19113 = ~pi0070 & ~n19112;
  assign n19114 = pi0070 & n19112;
  assign n19115 = ~n19113 & ~n19114;
  assign n19116 = pi3028 & pi9040;
  assign n19117 = ~pi2977 & ~pi9040;
  assign n19118 = ~n19116 & ~n19117;
  assign n19119 = pi0074 & n19118;
  assign n19120 = ~pi0074 & ~n19118;
  assign n19121 = ~n19119 & ~n19120;
  assign n19122 = pi2994 & pi9040;
  assign n19123 = pi3009 & ~pi9040;
  assign n19124 = ~n19122 & ~n19123;
  assign n19125 = ~pi0061 & n19124;
  assign n19126 = pi0061 & ~n19124;
  assign n19127 = ~n19125 & ~n19126;
  assign n19128 = pi3063 & ~pi9040;
  assign n19129 = pi3047 & pi9040;
  assign n19130 = ~n19128 & ~n19129;
  assign n19131 = pi0093 & n19130;
  assign n19132 = ~pi0093 & ~n19130;
  assign n19133 = ~n19131 & ~n19132;
  assign n19134 = pi2993 & ~pi9040;
  assign n19135 = pi3002 & pi9040;
  assign n19136 = ~n19134 & ~n19135;
  assign n19137 = ~pi0068 & n19136;
  assign n19138 = pi0068 & ~n19136;
  assign n19139 = ~n19137 & ~n19138;
  assign n19140 = ~n19133 & n19139;
  assign n19141 = n19127 & n19140;
  assign n19142 = ~n19121 & ~n19141;
  assign n19143 = pi2988 & ~pi9040;
  assign n19144 = pi2979 & pi9040;
  assign n19145 = ~n19143 & ~n19144;
  assign n19146 = ~pi0066 & n19145;
  assign n19147 = pi0066 & ~n19145;
  assign n19148 = ~n19146 & ~n19147;
  assign n19149 = n19133 & ~n19139;
  assign n19150 = n19148 & n19149;
  assign n19151 = ~n19127 & ~n19148;
  assign n19152 = ~n19127 & n19139;
  assign n19153 = ~n19151 & ~n19152;
  assign n19154 = ~n19133 & ~n19153;
  assign n19155 = n19127 & n19148;
  assign n19156 = ~n19139 & n19155;
  assign n19157 = n19121 & ~n19156;
  assign n19158 = ~n19154 & n19157;
  assign n19159 = ~n19150 & n19158;
  assign n19160 = ~n19142 & ~n19159;
  assign n19161 = n19127 & n19149;
  assign n19162 = ~n19148 & n19161;
  assign n19163 = ~n19160 & ~n19162;
  assign n19164 = n19115 & ~n19163;
  assign n19165 = ~n19121 & n19133;
  assign n19166 = n19152 & n19165;
  assign n19167 = n19115 & n19166;
  assign n19168 = ~n19164 & ~n19167;
  assign n19169 = ~n19127 & n19148;
  assign n19170 = ~n19139 & n19169;
  assign n19171 = ~n19133 & n19170;
  assign n19172 = ~n19121 & n19171;
  assign n19173 = ~n19121 & ~n19127;
  assign n19174 = ~n19133 & n19173;
  assign n19175 = ~n19139 & ~n19148;
  assign n19176 = n19133 & n19155;
  assign n19177 = ~n19175 & ~n19176;
  assign n19178 = ~n19121 & ~n19177;
  assign n19179 = ~n19174 & ~n19178;
  assign n19180 = n19139 & n19169;
  assign n19181 = n19133 & n19180;
  assign n19182 = n19127 & ~n19148;
  assign n19183 = n19139 & n19182;
  assign n19184 = ~n19181 & ~n19183;
  assign n19185 = n19121 & ~n19184;
  assign n19186 = ~n19139 & n19151;
  assign n19187 = n19133 & n19186;
  assign n19188 = ~n19185 & ~n19187;
  assign n19189 = n19179 & n19188;
  assign n19190 = ~n19171 & n19189;
  assign n19191 = ~n19115 & ~n19190;
  assign n19192 = n19133 & n19183;
  assign n19193 = n19133 & n19156;
  assign n19194 = n19139 & n19155;
  assign n19195 = ~n19133 & n19194;
  assign n19196 = ~n19193 & ~n19195;
  assign n19197 = ~n19192 & n19196;
  assign n19198 = n19139 & n19151;
  assign n19199 = ~n19133 & n19198;
  assign n19200 = n19197 & ~n19199;
  assign n19201 = n19121 & ~n19200;
  assign n19202 = ~n19191 & ~n19201;
  assign n19203 = ~n19172 & n19202;
  assign po0124 = ~n19168 | ~n19203;
  assign n19205 = ~n18612 & n18677;
  assign n19206 = ~n18612 & n18691;
  assign n19207 = ~n19205 & ~n19206;
  assign n19208 = ~n18606 & ~n19207;
  assign n19209 = ~n18606 & n19077;
  assign n19210 = ~n18612 & n19209;
  assign n19211 = ~n19208 & ~n19210;
  assign n19212 = ~n18647 & ~n18659;
  assign n19213 = n18618 & n18680;
  assign n19214 = ~n18645 & n19213;
  assign n19215 = ~n18650 & ~n19214;
  assign n19216 = n19212 & n19215;
  assign n19217 = ~n18644 & ~n19216;
  assign n19218 = ~n18618 & ~n18630;
  assign n19219 = ~n18967 & ~n19218;
  assign n19220 = ~n18606 & ~n19219;
  assign n19221 = ~n18644 & n19220;
  assign n19222 = n18606 & n18647;
  assign n19223 = ~n19221 & ~n19222;
  assign n19224 = ~n19217 & n19223;
  assign n19225 = n19211 & n19224;
  assign n19226 = n18612 & n19089;
  assign n19227 = ~n18968 & ~n19205;
  assign n19228 = ~n18612 & n18950;
  assign n19229 = n18612 & n18688;
  assign n19230 = ~n19228 & ~n19229;
  assign n19231 = ~n18606 & ~n19230;
  assign n19232 = n18612 & n18646;
  assign n19233 = ~n19231 & ~n19232;
  assign n19234 = ~n18683 & n19233;
  assign n19235 = n19227 & n19234;
  assign n19236 = ~n19226 & n19235;
  assign n19237 = n18644 & ~n19236;
  assign n19238 = n19225 & ~n19237;
  assign po0127 = ~n19083 & n19238;
  assign n19240 = n18373 & ~n18386;
  assign n19241 = ~n18370 & n18374;
  assign n19242 = n18364 & n18413;
  assign n19243 = ~n19241 & ~n19242;
  assign n19244 = ~n18386 & ~n19243;
  assign n19245 = ~n18378 & ~n19244;
  assign n19246 = ~n18373 & ~n18439;
  assign n19247 = n18370 & n18421;
  assign n19248 = ~n19028 & ~n19247;
  assign n19249 = ~n18408 & n19248;
  assign n19250 = n18386 & ~n19249;
  assign n19251 = ~n18370 & n18427;
  assign n19252 = ~n19250 & ~n19251;
  assign n19253 = n19246 & n19252;
  assign n19254 = n19245 & n19253;
  assign n19255 = ~n18400 & ~n19254;
  assign n19256 = n18370 & n18390;
  assign n19257 = ~n18415 & ~n19256;
  assign n19258 = n18386 & ~n19257;
  assign n19259 = ~n18374 & ~n18401;
  assign n19260 = n18403 & ~n19259;
  assign n19261 = ~n19021 & ~n19260;
  assign n19262 = ~n18377 & n19261;
  assign n19263 = n18386 & ~n19262;
  assign n19264 = n18370 & n18427;
  assign n19265 = ~n19263 & ~n19264;
  assign n19266 = ~n18370 & n19028;
  assign n19267 = n18370 & n18374;
  assign n19268 = ~n19266 & ~n19267;
  assign n19269 = ~n18408 & n19268;
  assign n19270 = ~n18386 & ~n19269;
  assign n19271 = n19265 & ~n19270;
  assign n19272 = n18400 & ~n19271;
  assign n19273 = ~n19258 & ~n19272;
  assign n19274 = ~n19255 & n19273;
  assign po0130 = n19240 | ~n19274;
  assign n19276 = ~n18755 & ~n18790;
  assign n19277 = ~n19062 & n19276;
  assign n19278 = ~n18711 & ~n19277;
  assign n19279 = ~n19054 & ~n19071;
  assign n19280 = ~n18758 & ~n18781;
  assign n19281 = ~n18745 & ~n18769;
  assign n19282 = n18711 & ~n19281;
  assign n19283 = ~n18735 & ~n19282;
  assign n19284 = n19280 & n19283;
  assign n19285 = n18767 & ~n19284;
  assign n19286 = ~n18717 & n18729;
  assign n19287 = ~n18883 & ~n19286;
  assign n19288 = n18705 & ~n19287;
  assign n19289 = ~n18748 & ~n19049;
  assign n19290 = n18711 & ~n19289;
  assign n19291 = n18705 & n18729;
  assign n19292 = ~n18752 & ~n19291;
  assign n19293 = ~n18730 & n19292;
  assign n19294 = ~n18711 & ~n19293;
  assign n19295 = ~n19290 & ~n19294;
  assign n19296 = ~n19288 & n19295;
  assign n19297 = ~n18767 & ~n19296;
  assign n19298 = ~n19285 & ~n19297;
  assign n19299 = n19279 & n19298;
  assign po0133 = n19278 | ~n19299;
  assign n19301 = ~n18261 & n18922;
  assign n19302 = ~n18247 & n18272;
  assign n19303 = ~n18252 & ~n19302;
  assign n19304 = n18261 & n19303;
  assign n19305 = ~n19301 & ~n19304;
  assign n19306 = ~n18915 & ~n19305;
  assign n19307 = ~n18267 & ~n19306;
  assign n19308 = n18261 & n18276;
  assign n19309 = ~n19307 & ~n19308;
  assign n19310 = ~n18273 & ~n18312;
  assign n19311 = ~n18261 & ~n19310;
  assign n19312 = n18227 & n18934;
  assign n19313 = ~n18301 & ~n19312;
  assign n19314 = n18233 & ~n19313;
  assign n19315 = n18247 & n18282;
  assign n19316 = ~n18261 & n18296;
  assign n19317 = ~n19315 & ~n19316;
  assign n19318 = ~n18295 & n19317;
  assign n19319 = ~n18302 & n19318;
  assign n19320 = ~n19314 & n19319;
  assign n19321 = n18267 & ~n19320;
  assign n19322 = ~n19311 & ~n19321;
  assign po0136 = ~n19309 | ~n19322;
  assign n19324 = ~n19133 & n19186;
  assign n19325 = n19133 & n19152;
  assign n19326 = ~n19170 & ~n19325;
  assign n19327 = n19121 & ~n19326;
  assign n19328 = ~n19324 & ~n19327;
  assign n19329 = ~n19121 & n19151;
  assign n19330 = ~n19133 & n19329;
  assign n19331 = n19165 & n19182;
  assign n19332 = ~n19330 & ~n19331;
  assign n19333 = ~n19121 & n19156;
  assign n19334 = n19332 & ~n19333;
  assign n19335 = ~n19181 & ~n19195;
  assign n19336 = ~n19161 & n19335;
  assign n19337 = n19334 & n19336;
  assign n19338 = n19328 & n19337;
  assign n19339 = ~n19115 & ~n19338;
  assign n19340 = ~n19170 & ~n19194;
  assign n19341 = n19133 & ~n19340;
  assign n19342 = n19140 & ~n19148;
  assign n19343 = ~n19139 & n19182;
  assign n19344 = ~n19342 & ~n19343;
  assign n19345 = ~n19127 & ~n19139;
  assign n19346 = n19133 & n19345;
  assign n19347 = n19344 & ~n19346;
  assign n19348 = n19121 & ~n19347;
  assign n19349 = ~n19133 & n19169;
  assign n19350 = n19133 & n19198;
  assign n19351 = ~n19349 & ~n19350;
  assign n19352 = ~n19121 & ~n19351;
  assign n19353 = ~n19133 & n19183;
  assign n19354 = ~n19352 & ~n19353;
  assign n19355 = ~n19348 & n19354;
  assign n19356 = ~n19341 & n19355;
  assign n19357 = n19115 & ~n19356;
  assign n19358 = n19121 & n19141;
  assign n19359 = ~n19357 & ~n19358;
  assign n19360 = ~n19121 & n19324;
  assign n19361 = n19359 & ~n19360;
  assign po0138 = ~n19339 & n19361;
  assign n19363 = ~n18370 & n18413;
  assign n19364 = ~n19019 & ~n19363;
  assign n19365 = n18386 & ~n19364;
  assign n19366 = ~n18426 & ~n19365;
  assign n19367 = ~n18400 & ~n19366;
  assign n19368 = ~n18386 & ~n18426;
  assign n19369 = ~n18364 & ~n19259;
  assign n19370 = n18370 & n19369;
  assign n19371 = ~n19021 & ~n19370;
  assign n19372 = n18386 & n19371;
  assign n19373 = ~n19368 & ~n19372;
  assign n19374 = ~n18386 & n19364;
  assign n19375 = n18351 & n18364;
  assign n19376 = ~n18370 & n19375;
  assign n19377 = ~n19369 & ~n19376;
  assign n19378 = ~n19256 & ~n19267;
  assign n19379 = n18386 & n19378;
  assign n19380 = n19377 & n19379;
  assign n19381 = ~n19374 & ~n19380;
  assign n19382 = n19371 & ~n19381;
  assign n19383 = n18400 & ~n19382;
  assign n19384 = n18370 & n18376;
  assign n19385 = ~n18439 & ~n19384;
  assign n19386 = ~n18386 & ~n19385;
  assign n19387 = ~n18386 & ~n19259;
  assign n19388 = n18364 & n19387;
  assign n19389 = ~n19386 & ~n19388;
  assign n19390 = ~n18370 & n19387;
  assign n19391 = n19389 & ~n19390;
  assign n19392 = ~n18400 & ~n19391;
  assign n19393 = ~n19383 & ~n19392;
  assign n19394 = ~n19373 & n19393;
  assign po0142 = n19367 | ~n19394;
  assign n19396 = ~n19193 & ~n19199;
  assign n19397 = ~n19121 & ~n19396;
  assign n19398 = n19139 & n19148;
  assign n19399 = n19133 & n19169;
  assign n19400 = ~n19398 & ~n19399;
  assign n19401 = ~n19133 & ~n19139;
  assign n19402 = ~n19148 & n19401;
  assign n19403 = n19400 & ~n19402;
  assign n19404 = n19121 & ~n19403;
  assign n19405 = ~n19192 & ~n19404;
  assign n19406 = n19133 & n19329;
  assign n19407 = ~n19333 & ~n19406;
  assign n19408 = n19405 & n19407;
  assign n19409 = ~n19115 & ~n19408;
  assign n19410 = n19121 & n19398;
  assign n19411 = n19133 & n19410;
  assign n19412 = ~n19409 & ~n19411;
  assign n19413 = ~n19133 & n19156;
  assign n19414 = ~n19186 & ~n19413;
  assign n19415 = n19121 & ~n19414;
  assign n19416 = ~n19170 & ~n19343;
  assign n19417 = ~n19141 & n19416;
  assign n19418 = ~n19121 & ~n19417;
  assign n19419 = ~n19162 & ~n19181;
  assign n19420 = ~n19342 & n19419;
  assign n19421 = ~n19418 & n19420;
  assign n19422 = ~n19415 & n19421;
  assign n19423 = n19115 & ~n19422;
  assign n19424 = n19412 & ~n19423;
  assign n19425 = ~n19172 & n19424;
  assign po0145 = n19397 | ~n19425;
  assign n19427 = ~pi3053 & ~pi9040;
  assign n19428 = pi2996 & pi9040;
  assign n19429 = ~n19427 & ~n19428;
  assign n19430 = ~pi0049 & ~n19429;
  assign n19431 = pi0049 & n19429;
  assign n19432 = ~n19430 & ~n19431;
  assign n19433 = pi2992 & pi9040;
  assign n19434 = pi3045 & ~pi9040;
  assign n19435 = ~n19433 & ~n19434;
  assign n19436 = pi0075 & n19435;
  assign n19437 = ~pi0075 & ~n19435;
  assign n19438 = ~n19436 & ~n19437;
  assign n19439 = pi3038 & pi9040;
  assign n19440 = pi2989 & ~pi9040;
  assign n19441 = ~n19439 & ~n19440;
  assign n19442 = ~pi0088 & ~n19441;
  assign n19443 = pi0088 & n19441;
  assign n19444 = ~n19442 & ~n19443;
  assign n19445 = pi3040 & ~pi9040;
  assign n19446 = pi3007 & pi9040;
  assign n19447 = ~n19445 & ~n19446;
  assign n19448 = ~pi0084 & n19447;
  assign n19449 = pi0084 & ~n19447;
  assign n19450 = ~n19448 & ~n19449;
  assign n19451 = pi3103 & pi9040;
  assign n19452 = pi3005 & ~pi9040;
  assign n19453 = ~n19451 & ~n19452;
  assign n19454 = ~pi0086 & n19453;
  assign n19455 = pi0086 & ~n19453;
  assign n19456 = ~n19454 & ~n19455;
  assign n19457 = n19450 & ~n19456;
  assign n19458 = n19444 & n19457;
  assign n19459 = pi2978 & pi9040;
  assign n19460 = pi3010 & ~pi9040;
  assign n19461 = ~n19459 & ~n19460;
  assign n19462 = pi0065 & n19461;
  assign n19463 = ~pi0065 & ~n19461;
  assign n19464 = ~n19462 & ~n19463;
  assign n19465 = ~n19450 & n19464;
  assign n19466 = n19456 & n19465;
  assign n19467 = ~n19444 & ~n19464;
  assign n19468 = ~n19450 & ~n19456;
  assign n19469 = n19450 & n19456;
  assign n19470 = ~n19468 & ~n19469;
  assign n19471 = n19467 & ~n19470;
  assign n19472 = ~n19466 & ~n19471;
  assign n19473 = ~n19458 & n19472;
  assign n19474 = ~n19438 & ~n19473;
  assign n19475 = ~n19432 & n19474;
  assign n19476 = n19464 & n19469;
  assign n19477 = ~n19450 & n19456;
  assign n19478 = ~n19464 & n19477;
  assign n19479 = ~n19456 & n19464;
  assign n19480 = ~n19444 & n19479;
  assign n19481 = ~n19478 & ~n19480;
  assign n19482 = n19444 & n19469;
  assign n19483 = n19481 & ~n19482;
  assign n19484 = ~n19476 & n19483;
  assign n19485 = n19438 & ~n19484;
  assign n19486 = ~n19444 & n19457;
  assign n19487 = n19464 & n19486;
  assign n19488 = ~n19485 & ~n19487;
  assign n19489 = ~n19432 & ~n19488;
  assign n19490 = n19438 & ~n19464;
  assign n19491 = n19444 & ~n19450;
  assign n19492 = n19456 & n19491;
  assign n19493 = n19490 & n19492;
  assign n19494 = ~n19456 & n19467;
  assign n19495 = n19450 & n19494;
  assign n19496 = n19438 & n19495;
  assign n19497 = ~n19493 & ~n19496;
  assign n19498 = ~n19438 & ~n19467;
  assign n19499 = ~n19470 & n19498;
  assign n19500 = ~n19444 & n19477;
  assign n19501 = ~n19438 & ~n19464;
  assign n19502 = n19500 & n19501;
  assign n19503 = ~n19477 & n19490;
  assign n19504 = ~n19444 & n19503;
  assign n19505 = n19444 & ~n19456;
  assign n19506 = n19464 & n19505;
  assign n19507 = ~n19466 & ~n19506;
  assign n19508 = n19438 & ~n19507;
  assign n19509 = ~n19504 & ~n19508;
  assign n19510 = ~n19495 & n19509;
  assign n19511 = ~n19502 & n19510;
  assign n19512 = ~n19499 & n19511;
  assign n19513 = n19432 & ~n19512;
  assign n19514 = n19497 & ~n19513;
  assign n19515 = n19444 & n19468;
  assign n19516 = ~n19438 & n19464;
  assign n19517 = n19515 & n19516;
  assign n19518 = n19514 & ~n19517;
  assign n19519 = ~n19489 & n19518;
  assign po0148 = n19475 | ~n19519;
  assign n19521 = ~n19162 & ~n19353;
  assign n19522 = n19121 & ~n19521;
  assign n19523 = ~n19115 & ~n19121;
  assign n19524 = n19152 & n19523;
  assign n19525 = n19148 & n19401;
  assign n19526 = ~n19345 & ~n19525;
  assign n19527 = ~n19183 & n19526;
  assign n19528 = n19121 & ~n19527;
  assign n19529 = ~n19133 & n19180;
  assign n19530 = ~n19528 & ~n19529;
  assign n19531 = ~n19115 & ~n19530;
  assign n19532 = ~n19524 & ~n19531;
  assign n19533 = ~n19133 & n19343;
  assign n19534 = n19196 & ~n19533;
  assign n19535 = ~n19325 & n19534;
  assign n19536 = ~n19121 & ~n19535;
  assign n19537 = n19139 & ~n19148;
  assign n19538 = n19165 & n19537;
  assign n19539 = ~n19133 & n19345;
  assign n19540 = ~n19193 & ~n19539;
  assign n19541 = ~n19350 & n19540;
  assign n19542 = ~n19538 & n19541;
  assign n19543 = n19121 & n19194;
  assign n19544 = n19542 & ~n19543;
  assign n19545 = n19115 & ~n19544;
  assign n19546 = ~n19536 & ~n19545;
  assign n19547 = n19532 & n19546;
  assign po0151 = n19522 | ~n19547;
  assign n19549 = n19438 & n19458;
  assign n19550 = ~n19444 & ~n19450;
  assign n19551 = ~n19466 & ~n19550;
  assign n19552 = n19438 & ~n19551;
  assign n19553 = ~n19549 & ~n19552;
  assign n19554 = n19432 & ~n19553;
  assign n19555 = n19432 & n19482;
  assign n19556 = n19464 & n19555;
  assign n19557 = ~n19554 & ~n19556;
  assign n19558 = ~n19444 & n19464;
  assign n19559 = ~n19450 & n19558;
  assign n19560 = ~n19464 & n19469;
  assign n19561 = ~n19444 & n19560;
  assign n19562 = ~n19559 & ~n19561;
  assign n19563 = n19438 & ~n19562;
  assign n19564 = n19464 & n19492;
  assign n19565 = ~n19438 & n19564;
  assign n19566 = n19444 & ~n19464;
  assign n19567 = ~n19470 & n19566;
  assign n19568 = ~n19495 & ~n19567;
  assign n19569 = n19458 & n19464;
  assign n19570 = ~n19444 & ~n19470;
  assign n19571 = n19464 & n19570;
  assign n19572 = ~n19569 & ~n19571;
  assign n19573 = ~n19502 & n19572;
  assign n19574 = n19568 & n19573;
  assign n19575 = ~n19565 & n19574;
  assign n19576 = n19444 & n19490;
  assign n19577 = n19456 & n19576;
  assign n19578 = n19575 & ~n19577;
  assign n19579 = ~n19432 & ~n19578;
  assign n19580 = ~n19486 & ~n19515;
  assign n19581 = ~n19450 & n19566;
  assign n19582 = n19580 & ~n19581;
  assign n19583 = n19432 & ~n19438;
  assign n19584 = ~n19582 & n19583;
  assign n19585 = ~n19579 & ~n19584;
  assign n19586 = ~n19563 & n19585;
  assign po0154 = ~n19557 | ~n19586;
  assign n19588 = ~n19476 & ~n19478;
  assign n19589 = n19438 & ~n19588;
  assign n19590 = ~n19496 & ~n19589;
  assign n19591 = n19432 & ~n19590;
  assign n19592 = ~n19444 & ~n19456;
  assign n19593 = ~n19468 & ~n19592;
  assign n19594 = ~n19464 & ~n19593;
  assign n19595 = ~n19492 & ~n19594;
  assign n19596 = ~n19438 & ~n19595;
  assign n19597 = ~n19471 & ~n19596;
  assign n19598 = n19464 & n19500;
  assign n19599 = n19450 & n19566;
  assign n19600 = n19464 & ~n19593;
  assign n19601 = ~n19599 & ~n19600;
  assign n19602 = n19438 & ~n19601;
  assign n19603 = ~n19598 & ~n19602;
  assign n19604 = n19597 & n19603;
  assign n19605 = ~n19432 & ~n19604;
  assign n19606 = n19438 & n19558;
  assign n19607 = n19468 & n19606;
  assign n19608 = n19444 & n19450;
  assign n19609 = n19516 & n19608;
  assign n19610 = ~n19607 & ~n19609;
  assign n19611 = n19444 & n19464;
  assign n19612 = n19432 & ~n19468;
  assign n19613 = n19611 & n19612;
  assign n19614 = n19610 & ~n19613;
  assign n19615 = ~n19479 & ~n19482;
  assign n19616 = n19583 & ~n19615;
  assign n19617 = n19614 & ~n19616;
  assign n19618 = ~n19605 & n19617;
  assign po0157 = n19591 | ~n19618;
  assign n19620 = ~n19444 & n19476;
  assign n19621 = ~n19569 & ~n19620;
  assign n19622 = n19438 & ~n19621;
  assign n19623 = n19457 & ~n19464;
  assign n19624 = ~n19476 & ~n19623;
  assign n19625 = ~n19438 & ~n19624;
  assign n19626 = ~n19564 & ~n19625;
  assign n19627 = n19438 & n19482;
  assign n19628 = ~n19500 & ~n19627;
  assign n19629 = n19580 & n19628;
  assign n19630 = ~n19464 & ~n19629;
  assign n19631 = n19626 & ~n19630;
  assign n19632 = n19432 & ~n19631;
  assign n19633 = ~n19500 & ~n19560;
  assign n19634 = ~n19515 & n19633;
  assign n19635 = ~n19438 & ~n19634;
  assign n19636 = ~n19444 & n19468;
  assign n19637 = ~n19492 & ~n19636;
  assign n19638 = n19438 & ~n19637;
  assign n19639 = ~n19635 & ~n19638;
  assign n19640 = ~n19549 & n19639;
  assign n19641 = ~n19561 & n19640;
  assign n19642 = ~n19432 & ~n19641;
  assign n19643 = n19516 & n19592;
  assign n19644 = ~n19642 & ~n19643;
  assign n19645 = ~n19632 & n19644;
  assign po0160 = n19622 | ~n19645;
  assign n19647 = pi3035 & pi9040;
  assign n19648 = pi3067 & ~pi9040;
  assign n19649 = ~n19647 & ~n19648;
  assign n19650 = ~pi0129 & n19649;
  assign n19651 = pi0129 & ~n19649;
  assign n19652 = ~n19650 & ~n19651;
  assign n19653 = pi3062 & pi9040;
  assign n19654 = pi3029 & ~pi9040;
  assign n19655 = ~n19653 & ~n19654;
  assign n19656 = ~pi0146 & n19655;
  assign n19657 = pi0146 & ~n19655;
  assign n19658 = ~n19656 & ~n19657;
  assign n19659 = pi3165 & pi9040;
  assign n19660 = pi3097 & ~pi9040;
  assign n19661 = ~n19659 & ~n19660;
  assign n19662 = ~pi0127 & n19661;
  assign n19663 = pi0127 & ~n19661;
  assign n19664 = ~n19662 & ~n19663;
  assign n19665 = n19658 & n19664;
  assign n19666 = pi3054 & pi9040;
  assign n19667 = pi3127 & ~pi9040;
  assign n19668 = ~n19666 & ~n19667;
  assign n19669 = pi0156 & n19668;
  assign n19670 = ~pi0156 & ~n19668;
  assign n19671 = ~n19669 & ~n19670;
  assign n19672 = pi3031 & pi9040;
  assign n19673 = pi3013 & ~pi9040;
  assign n19674 = ~n19672 & ~n19673;
  assign n19675 = ~pi0107 & ~n19674;
  assign n19676 = pi0107 & n19674;
  assign n19677 = ~n19675 & ~n19676;
  assign n19678 = n19671 & n19677;
  assign n19679 = n19665 & n19678;
  assign n19680 = ~n19658 & n19664;
  assign n19681 = ~n19677 & n19680;
  assign n19682 = n19671 & n19681;
  assign n19683 = ~n19679 & ~n19682;
  assign n19684 = ~n19658 & ~n19664;
  assign n19685 = ~n19677 & n19684;
  assign n19686 = ~n19671 & n19685;
  assign n19687 = n19665 & ~n19677;
  assign n19688 = ~n19671 & n19687;
  assign n19689 = ~n19686 & ~n19688;
  assign n19690 = n19683 & n19689;
  assign n19691 = ~n19652 & ~n19690;
  assign n19692 = n19671 & ~n19677;
  assign n19693 = ~n19664 & n19692;
  assign n19694 = n19658 & n19693;
  assign n19695 = ~n19681 & ~n19694;
  assign n19696 = ~n19652 & ~n19695;
  assign n19697 = ~n19664 & ~n19671;
  assign n19698 = n19652 & n19697;
  assign n19699 = ~n19658 & n19677;
  assign n19700 = n19665 & n19671;
  assign n19701 = ~n19699 & ~n19700;
  assign n19702 = n19652 & ~n19701;
  assign n19703 = ~n19698 & ~n19702;
  assign n19704 = n19658 & ~n19664;
  assign n19705 = n19677 & n19704;
  assign n19706 = ~n19671 & n19705;
  assign n19707 = n19703 & ~n19706;
  assign n19708 = ~n19664 & n19699;
  assign n19709 = n19671 & n19708;
  assign n19710 = n19707 & ~n19709;
  assign n19711 = ~n19696 & n19710;
  assign n19712 = pi3029 & pi9040;
  assign n19713 = pi3065 & ~pi9040;
  assign n19714 = ~n19712 & ~n19713;
  assign n19715 = pi0150 & n19714;
  assign n19716 = ~pi0150 & ~n19714;
  assign n19717 = ~n19715 & ~n19716;
  assign n19718 = ~n19711 & ~n19717;
  assign n19719 = ~n19664 & ~n19677;
  assign n19720 = n19652 & n19671;
  assign n19721 = n19717 & n19720;
  assign n19722 = n19719 & n19721;
  assign n19723 = ~n19671 & ~n19677;
  assign n19724 = n19664 & n19723;
  assign n19725 = n19652 & ~n19724;
  assign n19726 = n19658 & n19678;
  assign n19727 = ~n19684 & ~n19719;
  assign n19728 = ~n19671 & ~n19727;
  assign n19729 = n19665 & n19677;
  assign n19730 = ~n19728 & ~n19729;
  assign n19731 = ~n19652 & n19730;
  assign n19732 = ~n19726 & n19731;
  assign n19733 = ~n19725 & ~n19732;
  assign n19734 = n19677 & n19680;
  assign n19735 = n19671 & n19734;
  assign n19736 = ~n19733 & ~n19735;
  assign n19737 = n19717 & ~n19736;
  assign n19738 = ~n19722 & ~n19737;
  assign n19739 = ~n19718 & n19738;
  assign n19740 = ~n19691 & n19739;
  assign n19741 = n19652 & n19706;
  assign n19742 = n19740 & ~n19741;
  assign n19743 = pi0162 & ~n19742;
  assign n19744 = ~pi0162 & ~n19741;
  assign n19745 = n19739 & n19744;
  assign n19746 = ~n19691 & n19745;
  assign po0166 = n19743 | n19746;
  assign n19748 = pi3057 & pi9040;
  assign n19749 = pi3027 & ~pi9040;
  assign n19750 = ~n19748 & ~n19749;
  assign n19751 = pi0155 & n19750;
  assign n19752 = ~pi0155 & ~n19750;
  assign n19753 = ~n19751 & ~n19752;
  assign n19754 = pi3114 & pi9040;
  assign n19755 = pi3054 & ~pi9040;
  assign n19756 = ~n19754 & ~n19755;
  assign n19757 = pi0107 & n19756;
  assign n19758 = ~pi0107 & ~n19756;
  assign n19759 = ~n19757 & ~n19758;
  assign n19760 = pi3013 & pi9040;
  assign n19761 = pi3035 & ~pi9040;
  assign n19762 = ~n19760 & ~n19761;
  assign n19763 = pi0143 & n19762;
  assign n19764 = ~pi0143 & ~n19762;
  assign n19765 = ~n19763 & ~n19764;
  assign n19766 = pi3099 & pi9040;
  assign n19767 = pi3165 & ~pi9040;
  assign n19768 = ~n19766 & ~n19767;
  assign n19769 = pi0142 & n19768;
  assign n19770 = ~pi0142 & ~n19768;
  assign n19771 = ~n19769 & ~n19770;
  assign n19772 = ~n19765 & ~n19771;
  assign n19773 = n19759 & n19772;
  assign n19774 = n19753 & n19773;
  assign n19775 = n19765 & ~n19771;
  assign n19776 = ~n19759 & n19775;
  assign n19777 = n19753 & n19776;
  assign n19778 = pi3126 & pi9040;
  assign n19779 = pi3114 & ~pi9040;
  assign n19780 = ~n19778 & ~n19779;
  assign n19781 = ~pi0149 & n19780;
  assign n19782 = pi0149 & ~n19780;
  assign n19783 = ~n19781 & ~n19782;
  assign n19784 = ~n19759 & n19772;
  assign n19785 = ~n19753 & n19784;
  assign n19786 = n19753 & n19771;
  assign n19787 = ~n19785 & ~n19786;
  assign n19788 = ~n19783 & ~n19787;
  assign n19789 = ~n19777 & ~n19788;
  assign n19790 = ~n19774 & n19789;
  assign n19791 = n19765 & n19771;
  assign n19792 = ~n19759 & n19791;
  assign n19793 = ~n19753 & n19792;
  assign n19794 = ~n19753 & n19759;
  assign n19795 = n19771 & n19794;
  assign n19796 = ~n19765 & n19795;
  assign n19797 = ~n19771 & n19794;
  assign n19798 = n19765 & n19783;
  assign n19799 = n19797 & n19798;
  assign n19800 = ~n19796 & ~n19799;
  assign n19801 = ~n19793 & n19800;
  assign n19802 = n19790 & n19801;
  assign n19803 = pi3022 & pi9040;
  assign n19804 = pi3048 & ~pi9040;
  assign n19805 = ~n19803 & ~n19804;
  assign n19806 = pi0127 & n19805;
  assign n19807 = ~pi0127 & ~n19805;
  assign n19808 = ~n19806 & ~n19807;
  assign n19809 = ~n19802 & n19808;
  assign n19810 = n19753 & n19759;
  assign n19811 = ~n19771 & n19810;
  assign n19812 = n19765 & n19811;
  assign n19813 = ~n19753 & n19776;
  assign n19814 = ~n19812 & ~n19813;
  assign n19815 = ~n19783 & n19797;
  assign n19816 = n19765 & n19795;
  assign n19817 = ~n19815 & ~n19816;
  assign n19818 = n19753 & ~n19759;
  assign n19819 = ~n19771 & n19818;
  assign n19820 = ~n19765 & n19819;
  assign n19821 = ~n19753 & ~n19759;
  assign n19822 = n19771 & n19821;
  assign n19823 = ~n19765 & n19822;
  assign n19824 = ~n19820 & ~n19823;
  assign n19825 = n19759 & n19771;
  assign n19826 = n19753 & n19765;
  assign n19827 = ~n19825 & ~n19826;
  assign n19828 = ~n19759 & ~n19771;
  assign n19829 = n19827 & ~n19828;
  assign n19830 = n19783 & ~n19829;
  assign n19831 = n19824 & ~n19830;
  assign n19832 = n19817 & n19831;
  assign n19833 = n19814 & n19832;
  assign n19834 = ~n19808 & ~n19833;
  assign n19835 = ~n19809 & ~n19834;
  assign n19836 = pi0166 & ~n19835;
  assign n19837 = ~pi0166 & ~n19809;
  assign n19838 = ~n19834 & n19837;
  assign po0179 = n19836 | n19838;
  assign n19840 = pi3123 & pi9040;
  assign n19841 = pi3032 & ~pi9040;
  assign n19842 = ~n19840 & ~n19841;
  assign n19843 = ~pi0145 & n19842;
  assign n19844 = pi0145 & ~n19842;
  assign n19845 = ~n19843 & ~n19844;
  assign n19846 = pi3056 & pi9040;
  assign n19847 = pi3102 & ~pi9040;
  assign n19848 = ~n19846 & ~n19847;
  assign n19849 = ~pi0157 & n19848;
  assign n19850 = pi0157 & ~n19848;
  assign n19851 = ~n19849 & ~n19850;
  assign n19852 = pi3019 & pi9040;
  assign n19853 = pi3024 & ~pi9040;
  assign n19854 = ~n19852 & ~n19853;
  assign n19855 = ~pi0140 & ~n19854;
  assign n19856 = pi0140 & ~n19852;
  assign n19857 = ~n19853 & n19856;
  assign n19858 = ~n19855 & ~n19857;
  assign n19859 = pi3098 & pi9040;
  assign n19860 = pi3056 & ~pi9040;
  assign n19861 = ~n19859 & ~n19860;
  assign n19862 = ~pi0131 & n19861;
  assign n19863 = pi0131 & ~n19861;
  assign n19864 = ~n19862 & ~n19863;
  assign n19865 = pi3037 & pi9040;
  assign n19866 = pi3041 & ~pi9040;
  assign n19867 = ~n19865 & ~n19866;
  assign n19868 = ~pi0122 & ~n19867;
  assign n19869 = pi0122 & n19867;
  assign n19870 = ~n19868 & ~n19869;
  assign n19871 = ~n19864 & ~n19870;
  assign n19872 = n19858 & n19871;
  assign n19873 = n19851 & n19872;
  assign n19874 = ~n19845 & n19873;
  assign n19875 = ~n19864 & n19870;
  assign n19876 = ~n19858 & n19875;
  assign n19877 = ~n19845 & n19876;
  assign n19878 = n19851 & n19877;
  assign n19879 = pi3041 & pi9040;
  assign n19880 = pi3061 & ~pi9040;
  assign n19881 = ~n19879 & ~n19880;
  assign n19882 = pi0153 & n19881;
  assign n19883 = ~pi0153 & ~n19881;
  assign n19884 = ~n19882 & ~n19883;
  assign n19885 = n19845 & ~n19884;
  assign n19886 = ~n19851 & ~n19858;
  assign n19887 = ~n19870 & n19886;
  assign n19888 = ~n19858 & n19864;
  assign n19889 = ~n19887 & ~n19888;
  assign n19890 = n19885 & ~n19889;
  assign n19891 = ~n19878 & ~n19890;
  assign n19892 = ~n19845 & n19871;
  assign n19893 = ~n19851 & n19892;
  assign n19894 = n19864 & ~n19870;
  assign n19895 = ~n19858 & n19894;
  assign n19896 = ~n19845 & n19895;
  assign n19897 = n19864 & n19870;
  assign n19898 = n19858 & n19897;
  assign n19899 = ~n19851 & n19898;
  assign n19900 = n19858 & n19894;
  assign n19901 = n19851 & n19900;
  assign n19902 = ~n19899 & ~n19901;
  assign n19903 = ~n19851 & n19872;
  assign n19904 = ~n19858 & ~n19870;
  assign n19905 = ~n19864 & n19904;
  assign n19906 = n19851 & n19905;
  assign n19907 = ~n19851 & n19875;
  assign n19908 = ~n19906 & ~n19907;
  assign n19909 = n19845 & ~n19908;
  assign n19910 = ~n19903 & ~n19909;
  assign n19911 = n19902 & n19910;
  assign n19912 = ~n19896 & n19911;
  assign n19913 = ~n19893 & n19912;
  assign n19914 = n19884 & ~n19913;
  assign n19915 = n19858 & n19875;
  assign n19916 = n19851 & n19915;
  assign n19917 = ~n19901 & ~n19916;
  assign n19918 = n19845 & ~n19917;
  assign n19919 = ~n19858 & n19897;
  assign n19920 = n19845 & n19919;
  assign n19921 = n19851 & n19920;
  assign n19922 = ~n19918 & ~n19921;
  assign n19923 = n19851 & n19870;
  assign n19924 = ~n19858 & n19923;
  assign n19925 = ~n19873 & ~n19924;
  assign n19926 = ~n19845 & ~n19851;
  assign n19927 = n19858 & n19926;
  assign n19928 = ~n19871 & n19927;
  assign n19929 = ~n19845 & n19898;
  assign n19930 = ~n19928 & ~n19929;
  assign n19931 = n19925 & n19930;
  assign n19932 = ~n19884 & ~n19931;
  assign n19933 = n19922 & ~n19932;
  assign n19934 = ~n19914 & n19933;
  assign n19935 = n19891 & n19934;
  assign n19936 = ~n19874 & n19935;
  assign n19937 = pi0168 & n19936;
  assign n19938 = ~pi0168 & ~n19936;
  assign po0180 = n19937 | n19938;
  assign n19940 = n19851 & ~n19858;
  assign n19941 = n19864 & n19940;
  assign n19942 = ~n19870 & n19941;
  assign n19943 = ~n19851 & n19919;
  assign n19944 = ~n19942 & ~n19943;
  assign n19945 = ~n19845 & ~n19944;
  assign n19946 = ~n19873 & ~n19929;
  assign n19947 = n19851 & n19858;
  assign n19948 = ~n19870 & n19947;
  assign n19949 = ~n19924 & ~n19948;
  assign n19950 = n19845 & ~n19949;
  assign n19951 = n19845 & ~n19851;
  assign n19952 = n19894 & n19951;
  assign n19953 = ~n19858 & n19952;
  assign n19954 = ~n19851 & n19915;
  assign n19955 = ~n19845 & ~n19858;
  assign n19956 = ~n19864 & n19955;
  assign n19957 = ~n19870 & n19956;
  assign n19958 = ~n19954 & ~n19957;
  assign n19959 = ~n19953 & n19958;
  assign n19960 = ~n19950 & n19959;
  assign n19961 = n19946 & n19960;
  assign n19962 = n19884 & ~n19961;
  assign n19963 = n19845 & n19851;
  assign n19964 = n19872 & n19963;
  assign n19965 = ~n19845 & n19851;
  assign n19966 = n19897 & n19965;
  assign n19967 = n19858 & n19966;
  assign n19968 = ~n19964 & ~n19967;
  assign n19969 = ~n19962 & n19968;
  assign n19970 = ~n19945 & n19969;
  assign n19971 = n19858 & ~n19870;
  assign n19972 = n19926 & n19971;
  assign n19973 = ~n19896 & ~n19972;
  assign n19974 = n19851 & n19876;
  assign n19975 = ~n19845 & n19915;
  assign n19976 = ~n19974 & ~n19975;
  assign n19977 = ~n19851 & n19858;
  assign n19978 = n19864 & n19977;
  assign n19979 = ~n19870 & n19978;
  assign n19980 = ~n19942 & ~n19979;
  assign n19981 = ~n19851 & n19897;
  assign n19982 = ~n19858 & ~n19864;
  assign n19983 = ~n19981 & ~n19982;
  assign n19984 = n19845 & ~n19983;
  assign n19985 = n19980 & ~n19984;
  assign n19986 = n19976 & n19985;
  assign n19987 = n19973 & n19986;
  assign n19988 = ~n19884 & ~n19987;
  assign n19989 = n19970 & ~n19988;
  assign n19990 = ~pi0160 & ~n19989;
  assign n19991 = pi0160 & n19989;
  assign po0188 = n19990 | n19991;
  assign n19993 = ~n19671 & n19681;
  assign n19994 = ~n19735 & ~n19993;
  assign n19995 = ~n19652 & ~n19994;
  assign n19996 = ~n19664 & n19677;
  assign n19997 = ~n19671 & n19677;
  assign n19998 = n19658 & n19997;
  assign n19999 = ~n19996 & ~n19998;
  assign n20000 = ~n19681 & n19999;
  assign n20001 = ~n19652 & ~n20000;
  assign n20002 = ~n19677 & n19704;
  assign n20003 = ~n19671 & n20002;
  assign n20004 = ~n20001 & ~n20003;
  assign n20005 = ~n19717 & ~n20004;
  assign n20006 = ~n19717 & n19719;
  assign n20007 = n19652 & n20006;
  assign n20008 = ~n20005 & ~n20007;
  assign n20009 = ~n19995 & n20008;
  assign n20010 = ~n19658 & ~n19677;
  assign n20011 = n19652 & n20010;
  assign n20012 = n19671 & n20011;
  assign n20013 = ~n19658 & n19693;
  assign n20014 = ~n19671 & n19996;
  assign n20015 = ~n19679 & ~n20014;
  assign n20016 = ~n20013 & n20015;
  assign n20017 = ~n20012 & n20016;
  assign n20018 = ~n19652 & ~n19677;
  assign n20019 = n19665 & n20018;
  assign n20020 = n20017 & ~n20019;
  assign n20021 = n19717 & ~n20020;
  assign n20022 = ~n19679 & ~n19688;
  assign n20023 = ~n19671 & n19734;
  assign n20024 = ~n19664 & n19671;
  assign n20025 = ~n19677 & n20024;
  assign n20026 = ~n20023 & ~n20025;
  assign n20027 = n20022 & n20026;
  assign n20028 = n19652 & ~n20027;
  assign n20029 = ~n20021 & ~n20028;
  assign n20030 = n20009 & n20029;
  assign n20031 = pi0190 & n20030;
  assign n20032 = ~pi0190 & ~n20030;
  assign po0189 = n20031 | n20032;
  assign n20034 = ~n19688 & ~n19694;
  assign n20035 = n19652 & ~n19671;
  assign n20036 = ~n19664 & n20035;
  assign n20037 = ~n19658 & n20036;
  assign n20038 = n19680 & n19720;
  assign n20039 = ~n20037 & ~n20038;
  assign n20040 = n19652 & n19677;
  assign n20041 = n19665 & n20040;
  assign n20042 = n20039 & ~n20041;
  assign n20043 = ~n19671 & n19708;
  assign n20044 = ~n19705 & ~n20025;
  assign n20045 = ~n19652 & ~n20044;
  assign n20046 = ~n20043 & ~n20045;
  assign n20047 = n19664 & n19678;
  assign n20048 = n20046 & ~n20047;
  assign n20049 = n20042 & n20048;
  assign n20050 = n20034 & n20049;
  assign n20051 = ~n19717 & ~n20050;
  assign n20052 = ~n19687 & ~n19705;
  assign n20053 = n19671 & ~n20052;
  assign n20054 = ~n19671 & n19704;
  assign n20055 = ~n20013 & ~n20054;
  assign n20056 = n19652 & ~n20055;
  assign n20057 = ~n19658 & n19723;
  assign n20058 = ~n19734 & ~n20057;
  assign n20059 = n19671 & n19996;
  assign n20060 = n20058 & ~n20059;
  assign n20061 = ~n19652 & ~n20060;
  assign n20062 = ~n19993 & ~n20061;
  assign n20063 = ~n20056 & n20062;
  assign n20064 = ~n20053 & n20063;
  assign n20065 = n19717 & ~n20064;
  assign n20066 = ~n19652 & n19724;
  assign n20067 = ~n20065 & ~n20066;
  assign n20068 = n19699 & n20035;
  assign n20069 = ~n19664 & n20068;
  assign n20070 = n20067 & ~n20069;
  assign n20071 = ~n20051 & n20070;
  assign n20072 = ~pi0191 & ~n20071;
  assign n20073 = pi0191 & n20067;
  assign n20074 = ~n20051 & n20073;
  assign n20075 = ~n20069 & n20074;
  assign po0190 = n20072 | n20075;
  assign n20077 = pi3095 & pi9040;
  assign n20078 = pi3012 & ~pi9040;
  assign n20079 = ~n20077 & ~n20078;
  assign n20080 = ~pi0144 & ~n20079;
  assign n20081 = pi0144 & ~n20077;
  assign n20082 = ~n20078 & n20081;
  assign n20083 = ~n20080 & ~n20082;
  assign n20084 = pi3012 & pi9040;
  assign n20085 = pi3164 & ~pi9040;
  assign n20086 = ~n20084 & ~n20085;
  assign n20087 = pi0119 & n20086;
  assign n20088 = ~pi0119 & ~n20086;
  assign n20089 = ~n20087 & ~n20088;
  assign n20090 = pi3061 & pi9040;
  assign n20091 = pi3019 & ~pi9040;
  assign n20092 = ~n20090 & ~n20091;
  assign n20093 = pi0152 & n20092;
  assign n20094 = ~pi0152 & ~n20092;
  assign n20095 = ~n20093 & ~n20094;
  assign n20096 = n20089 & ~n20095;
  assign n20097 = pi3052 & pi9040;
  assign n20098 = pi3020 & ~pi9040;
  assign n20099 = ~n20097 & ~n20098;
  assign n20100 = ~pi0151 & n20099;
  assign n20101 = pi0151 & ~n20099;
  assign n20102 = ~n20100 & ~n20101;
  assign n20103 = pi3164 & pi9040;
  assign n20104 = pi3026 & ~pi9040;
  assign n20105 = ~n20103 & ~n20104;
  assign n20106 = ~pi0120 & n20105;
  assign n20107 = pi0120 & ~n20105;
  assign n20108 = ~n20106 & ~n20107;
  assign n20109 = ~n20102 & ~n20108;
  assign n20110 = n20096 & n20109;
  assign n20111 = ~n20102 & n20108;
  assign n20112 = ~n20089 & n20111;
  assign n20113 = ~n20110 & ~n20112;
  assign n20114 = ~n20083 & ~n20113;
  assign n20115 = pi3051 & pi9040;
  assign n20116 = pi3059 & ~pi9040;
  assign n20117 = ~n20115 & ~n20116;
  assign n20118 = pi0148 & n20117;
  assign n20119 = ~pi0148 & ~n20117;
  assign n20120 = ~n20118 & ~n20119;
  assign n20121 = n20089 & n20102;
  assign n20122 = n20083 & n20121;
  assign n20123 = n20096 & n20108;
  assign n20124 = n20089 & n20095;
  assign n20125 = ~n20108 & n20124;
  assign n20126 = ~n20123 & ~n20125;
  assign n20127 = ~n20089 & ~n20095;
  assign n20128 = ~n20108 & n20127;
  assign n20129 = ~n20102 & n20128;
  assign n20130 = n20126 & ~n20129;
  assign n20131 = n20083 & ~n20130;
  assign n20132 = ~n20122 & ~n20131;
  assign n20133 = ~n20089 & n20095;
  assign n20134 = n20108 & n20133;
  assign n20135 = ~n20102 & n20134;
  assign n20136 = n20132 & ~n20135;
  assign n20137 = n20102 & n20127;
  assign n20138 = ~n20089 & ~n20108;
  assign n20139 = n20095 & n20138;
  assign n20140 = ~n20137 & ~n20139;
  assign n20141 = ~n20083 & ~n20140;
  assign n20142 = n20108 & n20124;
  assign n20143 = n20102 & n20142;
  assign n20144 = ~n20141 & ~n20143;
  assign n20145 = n20136 & n20144;
  assign n20146 = n20120 & ~n20145;
  assign n20147 = ~n20114 & ~n20146;
  assign n20148 = n20083 & ~n20120;
  assign n20149 = ~n20140 & n20148;
  assign n20150 = n20108 & n20127;
  assign n20151 = ~n20142 & ~n20150;
  assign n20152 = ~n20102 & ~n20151;
  assign n20153 = ~n20110 & ~n20152;
  assign n20154 = ~n20120 & ~n20153;
  assign n20155 = ~n20149 & ~n20154;
  assign n20156 = ~n20083 & ~n20120;
  assign n20157 = n20096 & n20102;
  assign n20158 = ~n20134 & ~n20157;
  assign n20159 = n20089 & ~n20108;
  assign n20160 = n20158 & ~n20159;
  assign n20161 = n20156 & ~n20160;
  assign n20162 = n20155 & ~n20161;
  assign n20163 = n20147 & n20162;
  assign n20164 = ~pi0174 & ~n20163;
  assign n20165 = pi0174 & n20155;
  assign n20166 = n20147 & n20165;
  assign n20167 = ~n20161 & n20166;
  assign po0191 = n20164 | n20167;
  assign n20169 = ~n19765 & n19783;
  assign n20170 = n19794 & n20169;
  assign n20171 = n19771 & n19818;
  assign n20172 = ~n19813 & ~n20171;
  assign n20173 = n19765 & n19810;
  assign n20174 = n20172 & ~n20173;
  assign n20175 = n19783 & ~n20174;
  assign n20176 = n19753 & ~n19771;
  assign n20177 = ~n19765 & ~n19783;
  assign n20178 = n20176 & n20177;
  assign n20179 = ~n19820 & ~n20178;
  assign n20180 = ~n20175 & n20179;
  assign n20181 = ~n20170 & n20180;
  assign n20182 = n19771 & n19810;
  assign n20183 = n19765 & n20182;
  assign n20184 = ~n19796 & ~n20183;
  assign n20185 = n20181 & n20184;
  assign n20186 = ~n19808 & ~n20185;
  assign n20187 = n19765 & n19797;
  assign n20188 = ~n19793 & ~n19819;
  assign n20189 = ~n20187 & n20188;
  assign n20190 = ~n19783 & ~n20189;
  assign n20191 = ~n19753 & n19771;
  assign n20192 = ~n19765 & n20191;
  assign n20193 = n19765 & n19786;
  assign n20194 = ~n20192 & ~n20193;
  assign n20195 = n19783 & ~n20194;
  assign n20196 = ~n20190 & ~n20195;
  assign n20197 = ~n19774 & ~n19795;
  assign n20198 = n19783 & ~n20197;
  assign n20199 = ~n19785 & ~n20187;
  assign n20200 = n19753 & n19775;
  assign n20201 = ~n19765 & n20182;
  assign n20202 = ~n20200 & ~n20201;
  assign n20203 = ~n19783 & ~n20202;
  assign n20204 = n20199 & ~n20203;
  assign n20205 = ~n20198 & n20204;
  assign n20206 = n19808 & ~n20205;
  assign n20207 = ~n19783 & n19828;
  assign n20208 = ~n19765 & n20207;
  assign n20209 = ~n20206 & ~n20208;
  assign n20210 = n20196 & n20209;
  assign n20211 = ~n20186 & n20210;
  assign n20212 = pi0171 & n20211;
  assign n20213 = ~pi0171 & ~n20211;
  assign po0194 = n20212 | n20213;
  assign n20215 = n19851 & n19892;
  assign n20216 = n19870 & n19886;
  assign n20217 = ~n19919 & ~n20216;
  assign n20218 = ~n19845 & ~n20217;
  assign n20219 = ~n20215 & ~n20218;
  assign n20220 = n19875 & n19963;
  assign n20221 = n19845 & n19895;
  assign n20222 = ~n20220 & ~n20221;
  assign n20223 = n20219 & n20222;
  assign n20224 = n19870 & n19947;
  assign n20225 = ~n19942 & ~n20224;
  assign n20226 = ~n19979 & n20225;
  assign n20227 = n20223 & n20226;
  assign n20228 = ~n19884 & ~n20227;
  assign n20229 = ~n19873 & ~n19919;
  assign n20230 = ~n19981 & n20229;
  assign n20231 = n19845 & ~n20230;
  assign n20232 = ~n19851 & n19905;
  assign n20233 = ~n19954 & ~n20232;
  assign n20234 = ~n19878 & n20233;
  assign n20235 = ~n19845 & n19900;
  assign n20236 = n20234 & ~n20235;
  assign n20237 = ~n20231 & n20236;
  assign n20238 = n19884 & ~n20237;
  assign n20239 = ~n19942 & n20233;
  assign n20240 = n19845 & ~n20239;
  assign n20241 = ~n19967 & ~n19972;
  assign n20242 = ~n20240 & n20241;
  assign n20243 = ~n20238 & n20242;
  assign n20244 = ~n20228 & n20243;
  assign n20245 = pi0163 & n20244;
  assign n20246 = ~pi0163 & ~n20244;
  assign po0195 = n20245 | n20246;
  assign n20248 = ~n19887 & ~n19899;
  assign n20249 = n19884 & ~n20248;
  assign n20250 = n19845 & n19872;
  assign n20251 = ~n19864 & n19947;
  assign n20252 = ~n19948 & ~n20251;
  assign n20253 = n19845 & ~n20252;
  assign n20254 = ~n20250 & ~n20253;
  assign n20255 = n19884 & ~n20254;
  assign n20256 = ~n20249 & ~n20255;
  assign n20257 = n19898 & n19951;
  assign n20258 = ~n19924 & ~n19982;
  assign n20259 = ~n19845 & ~n20258;
  assign n20260 = n19884 & n20259;
  assign n20261 = ~n20257 & ~n20260;
  assign n20262 = ~n19953 & n20261;
  assign n20263 = n19851 & n19898;
  assign n20264 = n19851 & n19894;
  assign n20265 = ~n19943 & ~n20264;
  assign n20266 = ~n19845 & ~n20265;
  assign n20267 = ~n19873 & ~n19954;
  assign n20268 = n19851 & n19897;
  assign n20269 = ~n19876 & ~n20268;
  assign n20270 = n19845 & ~n20269;
  assign n20271 = n20267 & ~n20270;
  assign n20272 = ~n20266 & n20271;
  assign n20273 = ~n20263 & n20272;
  assign n20274 = ~n19884 & ~n20273;
  assign n20275 = ~n19979 & n20233;
  assign n20276 = ~n19845 & ~n20275;
  assign n20277 = ~n20274 & ~n20276;
  assign n20278 = n20262 & n20277;
  assign n20279 = n20256 & n20278;
  assign n20280 = ~pi0167 & ~n20279;
  assign n20281 = pi0167 & n20262;
  assign n20282 = n20256 & n20281;
  assign n20283 = n20277 & n20282;
  assign po0196 = n20280 | n20283;
  assign n20285 = ~n20083 & ~n20102;
  assign n20286 = ~n20127 & ~n20142;
  assign n20287 = n20285 & ~n20286;
  assign n20288 = ~n20083 & n20108;
  assign n20289 = n20127 & n20288;
  assign n20290 = ~n20287 & ~n20289;
  assign n20291 = n20120 & ~n20290;
  assign n20292 = n20102 & ~n20108;
  assign n20293 = n20095 & n20292;
  assign n20294 = n20089 & n20293;
  assign n20295 = ~n20159 & ~n20292;
  assign n20296 = n20083 & ~n20295;
  assign n20297 = n20102 & n20108;
  assign n20298 = ~n20095 & n20297;
  assign n20299 = n20089 & n20298;
  assign n20300 = ~n20296 & ~n20299;
  assign n20301 = ~n20294 & n20300;
  assign n20302 = n20120 & ~n20301;
  assign n20303 = ~n20291 & ~n20302;
  assign n20304 = n20095 & n20109;
  assign n20305 = ~n20089 & n20304;
  assign n20306 = n20102 & n20134;
  assign n20307 = ~n20305 & ~n20306;
  assign n20308 = ~n20083 & ~n20307;
  assign n20309 = ~n20095 & ~n20108;
  assign n20310 = ~n20134 & ~n20309;
  assign n20311 = n20102 & ~n20310;
  assign n20312 = n20095 & n20102;
  assign n20313 = n20288 & n20312;
  assign n20314 = ~n20096 & ~n20159;
  assign n20315 = ~n20102 & ~n20314;
  assign n20316 = ~n20134 & ~n20315;
  assign n20317 = ~n20083 & ~n20316;
  assign n20318 = n20083 & ~n20102;
  assign n20319 = n20124 & n20318;
  assign n20320 = n20108 & n20319;
  assign n20321 = ~n20317 & ~n20320;
  assign n20322 = ~n20313 & n20321;
  assign n20323 = ~n20311 & n20322;
  assign n20324 = ~n20305 & n20323;
  assign n20325 = ~n20120 & ~n20324;
  assign n20326 = n20102 & n20159;
  assign n20327 = ~n20102 & n20150;
  assign n20328 = ~n20326 & ~n20327;
  assign n20329 = n20083 & ~n20328;
  assign n20330 = ~n20325 & ~n20329;
  assign n20331 = ~n20308 & n20330;
  assign n20332 = n20303 & n20331;
  assign n20333 = pi0179 & n20332;
  assign n20334 = ~pi0179 & ~n20332;
  assign po0197 = n20333 | n20334;
  assign n20336 = pi3015 & pi9040;
  assign n20337 = pi3031 & ~pi9040;
  assign n20338 = ~n20336 & ~n20337;
  assign n20339 = ~pi0141 & n20338;
  assign n20340 = pi0141 & ~n20338;
  assign n20341 = ~n20339 & ~n20340;
  assign n20342 = pi3017 & ~pi9040;
  assign n20343 = pi3067 & pi9040;
  assign n20344 = ~n20342 & ~n20343;
  assign n20345 = ~pi0155 & ~n20344;
  assign n20346 = pi0155 & n20344;
  assign n20347 = ~n20345 & ~n20346;
  assign n20348 = n20341 & ~n20347;
  assign n20349 = pi3100 & pi9040;
  assign n20350 = pi3124 & ~pi9040;
  assign n20351 = ~n20349 & ~n20350;
  assign n20352 = ~pi0114 & n20351;
  assign n20353 = pi0114 & ~n20351;
  assign n20354 = ~n20352 & ~n20353;
  assign n20355 = pi3055 & pi9040;
  assign n20356 = pi3039 & ~pi9040;
  assign n20357 = ~n20355 & ~n20356;
  assign n20358 = ~pi0147 & ~n20357;
  assign n20359 = pi0147 & n20357;
  assign n20360 = ~n20358 & ~n20359;
  assign n20361 = pi3017 & pi9040;
  assign n20362 = pi3101 & ~pi9040;
  assign n20363 = ~n20361 & ~n20362;
  assign n20364 = ~pi0132 & ~n20363;
  assign n20365 = pi0132 & ~n20361;
  assign n20366 = ~n20362 & n20365;
  assign n20367 = ~n20364 & ~n20366;
  assign n20368 = n20360 & ~n20367;
  assign n20369 = n20354 & n20368;
  assign n20370 = pi3124 & pi9040;
  assign n20371 = pi3015 & ~pi9040;
  assign n20372 = ~n20370 & ~n20371;
  assign n20373 = ~pi0142 & n20372;
  assign n20374 = pi0142 & ~n20372;
  assign n20375 = ~n20373 & ~n20374;
  assign n20376 = n20367 & n20375;
  assign n20377 = n20360 & n20376;
  assign n20378 = ~n20354 & n20377;
  assign n20379 = n20367 & ~n20375;
  assign n20380 = n20354 & n20379;
  assign n20381 = ~n20378 & ~n20380;
  assign n20382 = ~n20369 & n20381;
  assign n20383 = n20348 & ~n20382;
  assign n20384 = n20354 & n20375;
  assign n20385 = ~n20360 & n20384;
  assign n20386 = ~n20367 & n20375;
  assign n20387 = n20360 & n20386;
  assign n20388 = ~n20354 & n20387;
  assign n20389 = ~n20385 & ~n20388;
  assign n20390 = ~n20360 & n20376;
  assign n20391 = n20360 & n20379;
  assign n20392 = ~n20390 & ~n20391;
  assign n20393 = n20389 & n20392;
  assign n20394 = ~n20341 & ~n20393;
  assign n20395 = ~n20367 & ~n20375;
  assign n20396 = ~n20360 & n20395;
  assign n20397 = ~n20354 & n20396;
  assign n20398 = ~n20394 & ~n20397;
  assign n20399 = ~n20347 & ~n20398;
  assign n20400 = ~n20383 & ~n20399;
  assign n20401 = ~n20341 & n20354;
  assign n20402 = n20360 & n20401;
  assign n20403 = ~n20375 & n20402;
  assign n20404 = n20354 & n20390;
  assign n20405 = ~n20403 & ~n20404;
  assign n20406 = ~n20379 & ~n20386;
  assign n20407 = ~n20354 & ~n20406;
  assign n20408 = ~n20360 & n20386;
  assign n20409 = ~n20407 & ~n20408;
  assign n20410 = n20341 & ~n20409;
  assign n20411 = n20360 & n20395;
  assign n20412 = ~n20369 & ~n20411;
  assign n20413 = ~n20378 & n20412;
  assign n20414 = ~n20341 & ~n20413;
  assign n20415 = ~n20410 & ~n20414;
  assign n20416 = n20341 & n20354;
  assign n20417 = n20376 & n20416;
  assign n20418 = ~n20354 & ~n20360;
  assign n20419 = n20375 & n20418;
  assign n20420 = ~n20367 & n20419;
  assign n20421 = ~n20360 & n20367;
  assign n20422 = ~n20375 & n20421;
  assign n20423 = ~n20354 & n20422;
  assign n20424 = ~n20420 & ~n20423;
  assign n20425 = n20354 & ~n20360;
  assign n20426 = ~n20375 & n20425;
  assign n20427 = ~n20367 & n20426;
  assign n20428 = n20424 & ~n20427;
  assign n20429 = ~n20417 & n20428;
  assign n20430 = n20415 & n20429;
  assign n20431 = n20347 & ~n20430;
  assign n20432 = n20405 & ~n20431;
  assign n20433 = n20400 & n20432;
  assign n20434 = pi0164 & ~n20433;
  assign n20435 = ~pi0164 & n20405;
  assign n20436 = n20400 & n20435;
  assign n20437 = ~n20431 & n20436;
  assign po0198 = n20434 | n20437;
  assign n20439 = n19658 & ~n19677;
  assign n20440 = ~n19652 & n20439;
  assign n20441 = n19671 & n20440;
  assign n20442 = n19671 & n19704;
  assign n20443 = ~n20439 & ~n20442;
  assign n20444 = ~n19658 & n19997;
  assign n20445 = n20443 & ~n20444;
  assign n20446 = ~n19652 & ~n20445;
  assign n20447 = ~n19682 & ~n20446;
  assign n20448 = ~n19717 & ~n20447;
  assign n20449 = n19652 & n19684;
  assign n20450 = n19671 & n20449;
  assign n20451 = ~n20041 & ~n20450;
  assign n20452 = ~n19717 & ~n20451;
  assign n20453 = ~n20448 & ~n20452;
  assign n20454 = ~n19705 & ~n19724;
  assign n20455 = ~n19734 & n20454;
  assign n20456 = n19652 & ~n20455;
  assign n20457 = ~n19671 & n19729;
  assign n20458 = ~n19708 & ~n20457;
  assign n20459 = ~n19652 & ~n20458;
  assign n20460 = ~n20057 & ~n20459;
  assign n20461 = ~n20456 & n20460;
  assign n20462 = ~n19694 & ~n19735;
  assign n20463 = n20461 & n20462;
  assign n20464 = n19717 & ~n20463;
  assign n20465 = ~n19679 & ~n19686;
  assign n20466 = n19652 & ~n20465;
  assign n20467 = ~n19741 & ~n20466;
  assign n20468 = ~n20464 & n20467;
  assign n20469 = n20453 & n20468;
  assign n20470 = ~n20441 & n20469;
  assign n20471 = pi0195 & n20470;
  assign n20472 = ~pi0195 & ~n20470;
  assign po0199 = n20471 | n20472;
  assign n20474 = ~n19783 & n20187;
  assign n20475 = ~n19794 & ~n19818;
  assign n20476 = n19772 & ~n20475;
  assign n20477 = ~n19822 & ~n20476;
  assign n20478 = ~n19812 & n20477;
  assign n20479 = n19783 & ~n20478;
  assign n20480 = n19765 & n20171;
  assign n20481 = ~n20479 & ~n20480;
  assign n20482 = n19765 & n19818;
  assign n20483 = ~n19771 & n19821;
  assign n20484 = ~n19765 & n19825;
  assign n20485 = ~n20483 & ~n20484;
  assign n20486 = ~n20482 & n20485;
  assign n20487 = ~n19783 & ~n20486;
  assign n20488 = n20481 & ~n20487;
  assign n20489 = n19808 & ~n20488;
  assign n20490 = ~n20474 & ~n20489;
  assign n20491 = ~n19765 & n19818;
  assign n20492 = ~n19811 & ~n20491;
  assign n20493 = ~n19783 & ~n20492;
  assign n20494 = ~n19793 & ~n20493;
  assign n20495 = ~n20183 & ~n20187;
  assign n20496 = n19765 & n19828;
  assign n20497 = ~n19825 & ~n20496;
  assign n20498 = ~n20483 & n20497;
  assign n20499 = n19783 & ~n20498;
  assign n20500 = ~n19765 & n20171;
  assign n20501 = ~n20499 & ~n20500;
  assign n20502 = n20495 & n20501;
  assign n20503 = n20494 & n20502;
  assign n20504 = ~n19808 & ~n20503;
  assign n20505 = n19765 & n20191;
  assign n20506 = ~n20201 & ~n20505;
  assign n20507 = n19783 & ~n20506;
  assign n20508 = ~n20504 & ~n20507;
  assign n20509 = n20490 & n20508;
  assign n20510 = pi0197 & n20509;
  assign n20511 = ~pi0197 & ~n20509;
  assign po0200 = n20510 | n20511;
  assign n20513 = ~n19783 & ~n20475;
  assign n20514 = ~n19765 & n20513;
  assign n20515 = n19765 & n19821;
  assign n20516 = ~n20183 & ~n20515;
  assign n20517 = ~n19783 & ~n20516;
  assign n20518 = ~n19771 & n20513;
  assign n20519 = ~n20517 & ~n20518;
  assign n20520 = ~n20514 & n20519;
  assign n20521 = ~n19808 & ~n20520;
  assign n20522 = n19771 & ~n20475;
  assign n20523 = n19765 & n20522;
  assign n20524 = ~n19812 & ~n20523;
  assign n20525 = ~n19765 & n19810;
  assign n20526 = ~n19823 & ~n20525;
  assign n20527 = ~n19783 & n20526;
  assign n20528 = ~n19753 & n19772;
  assign n20529 = ~n20482 & ~n20528;
  assign n20530 = n19783 & n20529;
  assign n20531 = ~n20522 & n20530;
  assign n20532 = ~n20505 & n20531;
  assign n20533 = ~n20527 & ~n20532;
  assign n20534 = n20524 & ~n20533;
  assign n20535 = n19808 & ~n20534;
  assign n20536 = ~n20521 & ~n20535;
  assign n20537 = n19783 & ~n20526;
  assign n20538 = ~n19813 & ~n20537;
  assign n20539 = ~n19808 & ~n20538;
  assign n20540 = ~n19783 & n19813;
  assign n20541 = n19783 & ~n20524;
  assign n20542 = ~n20540 & ~n20541;
  assign n20543 = ~n20539 & n20542;
  assign n20544 = n20536 & n20543;
  assign n20545 = pi0200 & n20544;
  assign n20546 = ~pi0200 & ~n20544;
  assign po0201 = n20545 | n20546;
  assign n20548 = pi3096 & ~pi9040;
  assign n20549 = pi3021 & pi9040;
  assign n20550 = ~n20548 & ~n20549;
  assign n20551 = ~pi0119 & ~n20550;
  assign n20552 = pi0119 & n20550;
  assign n20553 = ~n20551 & ~n20552;
  assign n20554 = pi3032 & pi9040;
  assign n20555 = pi3014 & ~pi9040;
  assign n20556 = ~n20554 & ~n20555;
  assign n20557 = ~pi0146 & n20556;
  assign n20558 = pi0146 & ~n20556;
  assign n20559 = ~n20557 & ~n20558;
  assign n20560 = pi3014 & pi9040;
  assign n20561 = pi3023 & ~pi9040;
  assign n20562 = ~n20560 & ~n20561;
  assign n20563 = ~pi0150 & n20562;
  assign n20564 = pi0150 & ~n20562;
  assign n20565 = ~n20563 & ~n20564;
  assign n20566 = pi3034 & pi9040;
  assign n20567 = pi3098 & ~pi9040;
  assign n20568 = ~n20566 & ~n20567;
  assign n20569 = ~pi0120 & ~n20568;
  assign n20570 = pi0120 & n20568;
  assign n20571 = ~n20569 & ~n20570;
  assign n20572 = n20565 & n20571;
  assign n20573 = pi3036 & ~pi9040;
  assign n20574 = pi3023 & pi9040;
  assign n20575 = ~n20573 & ~n20574;
  assign n20576 = ~pi0133 & n20575;
  assign n20577 = pi0133 & ~n20575;
  assign n20578 = ~n20576 & ~n20577;
  assign n20579 = pi3102 & pi9040;
  assign n20580 = pi3051 & ~pi9040;
  assign n20581 = ~n20579 & ~n20580;
  assign n20582 = ~pi0159 & n20581;
  assign n20583 = pi0159 & ~n20581;
  assign n20584 = ~n20582 & ~n20583;
  assign n20585 = ~n20578 & ~n20584;
  assign n20586 = n20572 & n20585;
  assign n20587 = ~n20559 & n20586;
  assign n20588 = n20578 & ~n20584;
  assign n20589 = ~n20565 & n20571;
  assign n20590 = n20588 & n20589;
  assign n20591 = ~n20559 & n20578;
  assign n20592 = ~n20571 & n20591;
  assign n20593 = n20565 & n20592;
  assign n20594 = ~n20565 & ~n20571;
  assign n20595 = ~n20559 & n20594;
  assign n20596 = ~n20584 & n20595;
  assign n20597 = ~n20578 & n20596;
  assign n20598 = ~n20593 & ~n20597;
  assign n20599 = ~n20590 & n20598;
  assign n20600 = ~n20587 & n20599;
  assign n20601 = n20559 & n20578;
  assign n20602 = n20571 & n20601;
  assign n20603 = ~n20565 & n20602;
  assign n20604 = n20600 & ~n20603;
  assign n20605 = ~n20553 & ~n20604;
  assign n20606 = ~n20559 & ~n20565;
  assign n20607 = n20571 & n20606;
  assign n20608 = ~n20578 & n20607;
  assign n20609 = ~n20592 & ~n20608;
  assign n20610 = n20559 & n20572;
  assign n20611 = ~n20578 & n20610;
  assign n20612 = n20609 & ~n20611;
  assign n20613 = n20584 & ~n20612;
  assign n20614 = n20559 & ~n20571;
  assign n20615 = ~n20565 & n20614;
  assign n20616 = ~n20578 & n20584;
  assign n20617 = n20615 & n20616;
  assign n20618 = n20565 & n20591;
  assign n20619 = n20565 & ~n20571;
  assign n20620 = n20578 & n20619;
  assign n20621 = ~n20618 & ~n20620;
  assign n20622 = n20584 & ~n20621;
  assign n20623 = ~n20617 & ~n20622;
  assign n20624 = ~n20553 & ~n20623;
  assign n20625 = ~n20613 & ~n20624;
  assign n20626 = ~n20605 & n20625;
  assign n20627 = n20559 & ~n20578;
  assign n20628 = ~n20584 & n20627;
  assign n20629 = n20619 & n20628;
  assign n20630 = n20559 & n20588;
  assign n20631 = ~n20565 & n20630;
  assign n20632 = n20584 & n20606;
  assign n20633 = n20565 & ~n20578;
  assign n20634 = n20559 & n20633;
  assign n20635 = ~n20610 & ~n20634;
  assign n20636 = ~n20632 & n20635;
  assign n20637 = n20578 & n20615;
  assign n20638 = n20636 & ~n20637;
  assign n20639 = n20572 & ~n20584;
  assign n20640 = n20578 & n20639;
  assign n20641 = n20559 & n20571;
  assign n20642 = ~n20578 & n20619;
  assign n20643 = ~n20641 & ~n20642;
  assign n20644 = ~n20584 & ~n20643;
  assign n20645 = ~n20640 & ~n20644;
  assign n20646 = n20638 & n20645;
  assign n20647 = n20553 & ~n20646;
  assign n20648 = ~n20631 & ~n20647;
  assign n20649 = ~n20629 & n20648;
  assign n20650 = n20626 & n20649;
  assign n20651 = pi0172 & n20650;
  assign n20652 = ~pi0172 & ~n20650;
  assign po0204 = n20651 | n20652;
  assign n20654 = ~n20354 & n20368;
  assign n20655 = ~n20391 & ~n20654;
  assign n20656 = ~n20404 & n20655;
  assign n20657 = ~n20341 & ~n20656;
  assign n20658 = n20354 & ~n20375;
  assign n20659 = n20421 & n20658;
  assign n20660 = n20354 & n20411;
  assign n20661 = ~n20360 & ~n20367;
  assign n20662 = ~n20376 & ~n20661;
  assign n20663 = ~n20354 & ~n20662;
  assign n20664 = ~n20660 & ~n20663;
  assign n20665 = ~n20659 & n20664;
  assign n20666 = n20341 & ~n20665;
  assign n20667 = ~n20657 & ~n20666;
  assign n20668 = n20347 & ~n20667;
  assign n20669 = ~n20367 & n20401;
  assign n20670 = n20354 & n20360;
  assign n20671 = n20367 & n20670;
  assign n20672 = ~n20654 & ~n20671;
  assign n20673 = n20341 & ~n20672;
  assign n20674 = ~n20417 & ~n20673;
  assign n20675 = ~n20341 & ~n20354;
  assign n20676 = n20421 & n20675;
  assign n20677 = ~n20341 & n20396;
  assign n20678 = ~n20676 & ~n20677;
  assign n20679 = n20354 & n20377;
  assign n20680 = ~n20423 & ~n20679;
  assign n20681 = n20678 & n20680;
  assign n20682 = n20674 & n20681;
  assign n20683 = ~n20669 & n20682;
  assign n20684 = ~n20347 & ~n20683;
  assign n20685 = n20408 & n20416;
  assign n20686 = n20360 & n20417;
  assign n20687 = ~n20685 & ~n20686;
  assign n20688 = ~n20341 & n20427;
  assign n20689 = n20687 & ~n20688;
  assign n20690 = n20354 & n20387;
  assign n20691 = ~n20354 & n20379;
  assign n20692 = ~n20690 & ~n20691;
  assign n20693 = ~n20341 & ~n20692;
  assign n20694 = n20689 & ~n20693;
  assign n20695 = ~n20684 & n20694;
  assign n20696 = ~n20668 & n20695;
  assign n20697 = ~pi0161 & n20696;
  assign n20698 = pi0161 & ~n20696;
  assign po0205 = n20697 | n20698;
  assign n20700 = pi3127 & pi9040;
  assign n20701 = pi3057 & ~pi9040;
  assign n20702 = ~n20700 & ~n20701;
  assign n20703 = ~pi0132 & ~n20702;
  assign n20704 = pi0132 & n20702;
  assign n20705 = ~n20703 & ~n20704;
  assign n20706 = pi3048 & pi9040;
  assign n20707 = pi3126 & ~pi9040;
  assign n20708 = ~n20706 & ~n20707;
  assign n20709 = pi0154 & n20708;
  assign n20710 = ~pi0154 & ~n20708;
  assign n20711 = ~n20709 & ~n20710;
  assign n20712 = pi3027 & pi9040;
  assign n20713 = pi3030 & ~pi9040;
  assign n20714 = ~n20712 & ~n20713;
  assign n20715 = ~pi0153 & ~n20714;
  assign n20716 = pi0153 & ~n20712;
  assign n20717 = ~n20713 & n20716;
  assign n20718 = ~n20715 & ~n20717;
  assign n20719 = pi3018 & pi9040;
  assign n20720 = pi3099 & ~pi9040;
  assign n20721 = ~n20719 & ~n20720;
  assign n20722 = ~pi0131 & n20721;
  assign n20723 = pi0131 & ~n20721;
  assign n20724 = ~n20722 & ~n20723;
  assign n20725 = pi3101 & pi9040;
  assign n20726 = pi3018 & ~pi9040;
  assign n20727 = ~n20725 & ~n20726;
  assign n20728 = ~pi0147 & ~n20727;
  assign n20729 = pi0147 & n20727;
  assign n20730 = ~n20728 & ~n20729;
  assign n20731 = ~n20724 & ~n20730;
  assign n20732 = n20718 & n20731;
  assign n20733 = n20711 & n20732;
  assign n20734 = ~n20711 & ~n20724;
  assign n20735 = n20730 & n20734;
  assign n20736 = pi3039 & pi9040;
  assign n20737 = pi3022 & ~pi9040;
  assign n20738 = ~n20736 & ~n20737;
  assign n20739 = ~pi0112 & n20738;
  assign n20740 = pi0112 & ~n20738;
  assign n20741 = ~n20739 & ~n20740;
  assign n20742 = ~n20718 & n20734;
  assign n20743 = n20718 & n20730;
  assign n20744 = n20724 & n20743;
  assign n20745 = ~n20742 & ~n20744;
  assign n20746 = n20741 & ~n20745;
  assign n20747 = ~n20735 & ~n20746;
  assign n20748 = ~n20724 & n20743;
  assign n20749 = ~n20718 & n20724;
  assign n20750 = n20724 & ~n20730;
  assign n20751 = ~n20711 & n20750;
  assign n20752 = ~n20718 & ~n20730;
  assign n20753 = n20711 & n20752;
  assign n20754 = ~n20751 & ~n20753;
  assign n20755 = ~n20749 & n20754;
  assign n20756 = ~n20748 & n20755;
  assign n20757 = ~n20741 & ~n20756;
  assign n20758 = n20747 & ~n20757;
  assign n20759 = ~n20733 & n20758;
  assign n20760 = n20705 & ~n20759;
  assign n20761 = ~n20718 & n20730;
  assign n20762 = n20724 & n20761;
  assign n20763 = ~n20711 & n20762;
  assign n20764 = n20724 & n20752;
  assign n20765 = n20711 & n20764;
  assign n20766 = ~n20733 & ~n20765;
  assign n20767 = ~n20763 & n20766;
  assign n20768 = ~n20741 & ~n20767;
  assign n20769 = ~n20760 & ~n20768;
  assign n20770 = n20718 & n20735;
  assign n20771 = n20711 & n20724;
  assign n20772 = n20741 & n20771;
  assign n20773 = n20718 & n20772;
  assign n20774 = ~n20711 & ~n20741;
  assign n20775 = n20731 & n20774;
  assign n20776 = ~n20724 & n20761;
  assign n20777 = n20711 & n20776;
  assign n20778 = ~n20775 & ~n20777;
  assign n20779 = ~n20718 & ~n20724;
  assign n20780 = n20711 & n20779;
  assign n20781 = n20718 & ~n20730;
  assign n20782 = n20724 & n20781;
  assign n20783 = ~n20780 & ~n20782;
  assign n20784 = n20741 & ~n20783;
  assign n20785 = n20741 & n20749;
  assign n20786 = ~n20711 & n20785;
  assign n20787 = ~n20784 & ~n20786;
  assign n20788 = n20778 & n20787;
  assign n20789 = ~n20705 & ~n20788;
  assign n20790 = ~n20773 & ~n20789;
  assign n20791 = ~n20770 & n20790;
  assign n20792 = n20769 & n20791;
  assign n20793 = ~pi0169 & ~n20792;
  assign n20794 = ~n20760 & ~n20770;
  assign n20795 = ~n20768 & n20794;
  assign n20796 = n20790 & n20795;
  assign n20797 = pi0169 & n20796;
  assign po0206 = n20793 | n20797;
  assign n20799 = ~n20341 & n20379;
  assign n20800 = n20354 & n20799;
  assign n20801 = ~n20690 & ~n20800;
  assign n20802 = n20354 & ~n20367;
  assign n20803 = n20375 & n20670;
  assign n20804 = ~n20802 & ~n20803;
  assign n20805 = n20341 & ~n20804;
  assign n20806 = ~n20354 & n20360;
  assign n20807 = ~n20375 & n20806;
  assign n20808 = ~n20805 & ~n20807;
  assign n20809 = n20801 & n20808;
  assign n20810 = n20347 & ~n20809;
  assign n20811 = ~n20377 & ~n20423;
  assign n20812 = n20354 & n20395;
  assign n20813 = n20811 & ~n20812;
  assign n20814 = ~n20341 & ~n20813;
  assign n20815 = n20379 & n20416;
  assign n20816 = ~n20404 & ~n20815;
  assign n20817 = ~n20814 & n20816;
  assign n20818 = ~n20387 & ~n20397;
  assign n20819 = n20341 & ~n20818;
  assign n20820 = n20817 & ~n20819;
  assign n20821 = ~n20347 & ~n20820;
  assign n20822 = ~n20810 & ~n20821;
  assign n20823 = ~n20408 & ~n20411;
  assign n20824 = ~n20377 & n20823;
  assign n20825 = ~n20354 & ~n20824;
  assign n20826 = ~n20341 & n20825;
  assign n20827 = n20354 & ~n20386;
  assign n20828 = ~n20354 & n20392;
  assign n20829 = ~n20827 & ~n20828;
  assign n20830 = n20341 & n20829;
  assign n20831 = ~n20826 & ~n20830;
  assign n20832 = n20822 & n20831;
  assign n20833 = ~pi0165 & ~n20832;
  assign n20834 = ~n20821 & n20831;
  assign n20835 = pi0165 & n20834;
  assign n20836 = ~n20810 & n20835;
  assign po0207 = n20833 | n20836;
  assign n20838 = ~n20559 & n20565;
  assign n20839 = ~n20603 & ~n20838;
  assign n20840 = ~n20633 & n20839;
  assign n20841 = ~n20584 & ~n20840;
  assign n20842 = ~n20565 & n20616;
  assign n20843 = ~n20559 & ~n20578;
  assign n20844 = n20571 & n20843;
  assign n20845 = n20578 & n20595;
  assign n20846 = ~n20844 & ~n20845;
  assign n20847 = n20559 & n20565;
  assign n20848 = n20578 & n20584;
  assign n20849 = n20847 & n20848;
  assign n20850 = n20846 & ~n20849;
  assign n20851 = ~n20842 & n20850;
  assign n20852 = ~n20841 & n20851;
  assign n20853 = n20553 & ~n20852;
  assign n20854 = ~n20559 & n20572;
  assign n20855 = n20578 & n20854;
  assign n20856 = ~n20571 & n20838;
  assign n20857 = ~n20578 & n20856;
  assign n20858 = ~n20855 & ~n20857;
  assign n20859 = ~n20584 & ~n20858;
  assign n20860 = ~n20853 & ~n20859;
  assign n20861 = ~n20578 & n20595;
  assign n20862 = ~n20607 & ~n20615;
  assign n20863 = ~n20584 & ~n20862;
  assign n20864 = ~n20861 & ~n20863;
  assign n20865 = ~n20611 & n20864;
  assign n20866 = ~n20553 & ~n20865;
  assign n20867 = ~n20589 & ~n20619;
  assign n20868 = n20559 & ~n20867;
  assign n20869 = ~n20620 & ~n20868;
  assign n20870 = n20584 & ~n20869;
  assign n20871 = ~n20553 & n20870;
  assign n20872 = ~n20866 & ~n20871;
  assign n20873 = n20860 & n20872;
  assign n20874 = pi0173 & ~n20873;
  assign n20875 = ~pi0173 & n20860;
  assign n20876 = n20872 & n20875;
  assign po0213 = n20874 | n20876;
  assign n20878 = ~n20095 & n20111;
  assign n20879 = ~n20142 & ~n20878;
  assign n20880 = ~n20083 & ~n20879;
  assign n20881 = ~n20102 & n20133;
  assign n20882 = ~n20298 & ~n20881;
  assign n20883 = n20083 & ~n20882;
  assign n20884 = n20102 & n20128;
  assign n20885 = ~n20313 & ~n20884;
  assign n20886 = ~n20110 & n20885;
  assign n20887 = ~n20883 & n20886;
  assign n20888 = ~n20880 & n20887;
  assign n20889 = ~n20294 & ~n20305;
  assign n20890 = n20888 & n20889;
  assign n20891 = n20120 & ~n20890;
  assign n20892 = n20096 & n20292;
  assign n20893 = n20151 & ~n20892;
  assign n20894 = n20083 & ~n20893;
  assign n20895 = n20102 & n20139;
  assign n20896 = ~n20894 & ~n20895;
  assign n20897 = n20089 & n20111;
  assign n20898 = ~n20102 & n20124;
  assign n20899 = ~n20897 & ~n20898;
  assign n20900 = n20083 & ~n20899;
  assign n20901 = n20083 & n20133;
  assign n20902 = n20102 & n20901;
  assign n20903 = ~n20900 & ~n20902;
  assign n20904 = n20896 & n20903;
  assign n20905 = ~n20120 & ~n20904;
  assign n20906 = ~n20128 & ~n20135;
  assign n20907 = ~n20299 & n20906;
  assign n20908 = n20156 & ~n20907;
  assign n20909 = ~n20905 & ~n20908;
  assign n20910 = ~n20110 & ~n20294;
  assign n20911 = ~n20083 & ~n20910;
  assign n20912 = n20909 & ~n20911;
  assign n20913 = ~n20891 & n20912;
  assign n20914 = ~pi0192 & n20913;
  assign n20915 = pi0192 & ~n20913;
  assign po0214 = n20914 | n20915;
  assign n20917 = n20354 & n20422;
  assign n20918 = n20341 & n20917;
  assign n20919 = ~n20686 & ~n20918;
  assign n20920 = ~n20427 & ~n20803;
  assign n20921 = ~n20341 & n20367;
  assign n20922 = n20670 & n20921;
  assign n20923 = ~n20354 & n20411;
  assign n20924 = n20341 & n20421;
  assign n20925 = ~n20923 & ~n20924;
  assign n20926 = ~n20420 & n20925;
  assign n20927 = ~n20922 & n20926;
  assign n20928 = n20920 & n20927;
  assign n20929 = ~n20677 & n20928;
  assign n20930 = n20347 & ~n20929;
  assign n20931 = ~n20354 & n20367;
  assign n20932 = ~n20421 & ~n20931;
  assign n20933 = ~n20387 & n20932;
  assign n20934 = ~n20341 & ~n20933;
  assign n20935 = n20341 & ~n20823;
  assign n20936 = ~n20354 & n20391;
  assign n20937 = ~n20935 & ~n20936;
  assign n20938 = ~n20934 & n20937;
  assign n20939 = ~n20347 & ~n20938;
  assign n20940 = ~n20930 & ~n20939;
  assign n20941 = ~n20688 & n20940;
  assign n20942 = n20919 & n20941;
  assign n20943 = pi0175 & n20942;
  assign n20944 = ~pi0175 & ~n20942;
  assign po0215 = n20943 | n20944;
  assign n20946 = ~n20711 & n20741;
  assign n20947 = n20718 & n20946;
  assign n20948 = ~n20724 & n20752;
  assign n20949 = n20711 & n20948;
  assign n20950 = n20711 & n20762;
  assign n20951 = ~n20949 & ~n20950;
  assign n20952 = ~n20711 & n20764;
  assign n20953 = ~n20744 & ~n20952;
  assign n20954 = ~n20741 & ~n20953;
  assign n20955 = n20951 & ~n20954;
  assign n20956 = ~n20947 & n20955;
  assign n20957 = n20705 & ~n20956;
  assign n20958 = n20711 & n20718;
  assign n20959 = n20724 & n20958;
  assign n20960 = ~n20730 & n20959;
  assign n20961 = n20741 & n20960;
  assign n20962 = n20774 & n20782;
  assign n20963 = ~n20742 & ~n20962;
  assign n20964 = ~n20744 & ~n20776;
  assign n20965 = ~n20711 & n20761;
  assign n20966 = n20964 & ~n20965;
  assign n20967 = n20741 & ~n20966;
  assign n20968 = ~n20741 & n20748;
  assign n20969 = n20766 & ~n20968;
  assign n20970 = ~n20967 & n20969;
  assign n20971 = n20963 & n20970;
  assign n20972 = ~n20705 & ~n20971;
  assign n20973 = ~n20961 & ~n20972;
  assign n20974 = ~n20957 & n20973;
  assign n20975 = n20774 & n20776;
  assign n20976 = n20731 & ~n20741;
  assign n20977 = n20711 & n20976;
  assign n20978 = ~n20975 & ~n20977;
  assign n20979 = ~n20741 & n20950;
  assign n20980 = n20978 & ~n20979;
  assign n20981 = n20974 & n20980;
  assign n20982 = ~pi0170 & ~n20981;
  assign n20983 = pi0170 & n20980;
  assign n20984 = n20973 & n20983;
  assign n20985 = ~n20957 & n20984;
  assign po0216 = n20982 | n20985;
  assign n20987 = pi3049 & pi9040;
  assign n20988 = pi3037 & ~pi9040;
  assign n20989 = ~n20987 & ~n20988;
  assign n20990 = ~pi0152 & ~n20989;
  assign n20991 = pi0152 & n20989;
  assign n20992 = ~n20990 & ~n20991;
  assign n20993 = pi3050 & pi9040;
  assign n20994 = pi3123 & ~pi9040;
  assign n20995 = ~n20993 & ~n20994;
  assign n20996 = ~pi0148 & n20995;
  assign n20997 = pi0148 & ~n20995;
  assign n20998 = ~n20996 & ~n20997;
  assign n20999 = pi3036 & pi9040;
  assign n21000 = pi3034 & ~pi9040;
  assign n21001 = ~n20999 & ~n21000;
  assign n21002 = ~pi0140 & n21001;
  assign n21003 = pi0140 & ~n21001;
  assign n21004 = ~n21002 & ~n21003;
  assign n21005 = n20998 & ~n21004;
  assign n21006 = n20992 & n21005;
  assign n21007 = pi3024 & pi9040;
  assign n21008 = pi3021 & ~pi9040;
  assign n21009 = ~n21007 & ~n21008;
  assign n21010 = pi0106 & n21009;
  assign n21011 = ~pi0106 & ~n21009;
  assign n21012 = ~n21010 & ~n21011;
  assign n21013 = pi3020 & pi9040;
  assign n21014 = pi3025 & ~pi9040;
  assign n21015 = ~n21013 & ~n21014;
  assign n21016 = pi0134 & n21015;
  assign n21017 = ~pi0134 & ~n21015;
  assign n21018 = ~n21016 & ~n21017;
  assign n21019 = n21012 & ~n21018;
  assign n21020 = n21006 & n21019;
  assign n21021 = ~n20998 & n21004;
  assign n21022 = n21019 & n21021;
  assign n21023 = ~n20992 & n21022;
  assign n21024 = ~n21020 & ~n21023;
  assign n21025 = ~n20992 & n21005;
  assign n21026 = ~n21012 & n21025;
  assign n21027 = ~n21018 & n21026;
  assign n21028 = ~n20992 & n21021;
  assign n21029 = ~n21018 & n21028;
  assign n21030 = ~n21027 & ~n21029;
  assign n21031 = ~n20998 & n21018;
  assign n21032 = n20992 & n21031;
  assign n21033 = n21005 & n21018;
  assign n21034 = ~n21032 & ~n21033;
  assign n21035 = n21012 & ~n21034;
  assign n21036 = ~n20998 & ~n21004;
  assign n21037 = n20998 & n21004;
  assign n21038 = ~n21036 & ~n21037;
  assign n21039 = ~n20992 & ~n21018;
  assign n21040 = ~n21012 & ~n21039;
  assign n21041 = ~n21038 & n21040;
  assign n21042 = ~n20992 & ~n21005;
  assign n21043 = n21012 & n21042;
  assign n21044 = ~n21018 & n21043;
  assign n21045 = ~n21041 & ~n21044;
  assign n21046 = ~n21035 & n21045;
  assign n21047 = n21030 & n21046;
  assign n21048 = pi3096 & pi9040;
  assign n21049 = pi3050 & ~pi9040;
  assign n21050 = ~n21048 & ~n21049;
  assign n21051 = ~pi0122 & n21050;
  assign n21052 = pi0122 & ~n21050;
  assign n21053 = ~n21051 & ~n21052;
  assign n21054 = ~n21047 & ~n21053;
  assign n21055 = n21024 & ~n21054;
  assign n21056 = n20992 & n21036;
  assign n21057 = ~n21012 & n21056;
  assign n21058 = n21018 & n21057;
  assign n21059 = ~n21012 & n21053;
  assign n21060 = n20992 & n21021;
  assign n21061 = ~n21038 & n21039;
  assign n21062 = ~n21033 & ~n21061;
  assign n21063 = ~n21060 & n21062;
  assign n21064 = n21059 & ~n21063;
  assign n21065 = n21018 & n21028;
  assign n21066 = ~n20992 & n21031;
  assign n21067 = n21018 & n21037;
  assign n21068 = ~n21066 & ~n21067;
  assign n21069 = n21005 & ~n21018;
  assign n21070 = n20992 & n21037;
  assign n21071 = ~n21069 & ~n21070;
  assign n21072 = n21068 & n21071;
  assign n21073 = n21012 & ~n21072;
  assign n21074 = ~n21065 & ~n21073;
  assign n21075 = n21053 & ~n21074;
  assign n21076 = ~n21064 & ~n21075;
  assign n21077 = ~n21058 & n21076;
  assign n21078 = n21055 & n21077;
  assign n21079 = pi0186 & ~n21078;
  assign n21080 = ~pi0186 & n21055;
  assign n21081 = n21077 & n21080;
  assign po0217 = n21079 | n21081;
  assign n21083 = ~n20578 & ~n20867;
  assign n21084 = n20559 & n21083;
  assign n21085 = ~n20571 & n20843;
  assign n21086 = ~n20641 & ~n21085;
  assign n21087 = ~n20856 & n21086;
  assign n21088 = ~n20584 & ~n21087;
  assign n21089 = ~n20614 & ~n20854;
  assign n21090 = n20584 & ~n21089;
  assign n21091 = ~n21088 & ~n21090;
  assign n21092 = ~n21084 & n21091;
  assign n21093 = n20578 & n20607;
  assign n21094 = n21092 & ~n21093;
  assign n21095 = ~n20553 & ~n21094;
  assign n21096 = n20588 & ~n21089;
  assign n21097 = ~n20610 & ~n20615;
  assign n21098 = ~n20607 & ~n20856;
  assign n21099 = n21097 & n21098;
  assign n21100 = ~n20578 & ~n21099;
  assign n21101 = ~n21096 & ~n21100;
  assign n21102 = ~n20845 & n21101;
  assign n21103 = n20553 & ~n21102;
  assign n21104 = ~n21095 & ~n21103;
  assign n21105 = ~n20578 & n20854;
  assign n21106 = ~n21093 & ~n21105;
  assign n21107 = n20584 & ~n21106;
  assign n21108 = n21104 & ~n21107;
  assign n21109 = pi0189 & ~n21108;
  assign n21110 = ~pi0189 & ~n21107;
  assign n21111 = ~n21103 & n21110;
  assign n21112 = ~n21095 & n21111;
  assign po0218 = n21109 | n21112;
  assign n21114 = ~n20730 & n20734;
  assign n21115 = ~n20718 & n21114;
  assign n21116 = ~n20762 & ~n20770;
  assign n21117 = n20711 & n20731;
  assign n21118 = ~n20711 & n20782;
  assign n21119 = ~n21117 & ~n21118;
  assign n21120 = n21116 & n21119;
  assign n21121 = n20741 & ~n21120;
  assign n21122 = n20711 & n20743;
  assign n21123 = ~n20742 & ~n21122;
  assign n21124 = ~n20764 & n21123;
  assign n21125 = ~n20741 & ~n21124;
  assign n21126 = n20730 & n20771;
  assign n21127 = n20718 & n21126;
  assign n21128 = ~n21125 & ~n21127;
  assign n21129 = ~n21121 & n21128;
  assign n21130 = ~n21115 & n21129;
  assign n21131 = ~n20705 & ~n21130;
  assign n21132 = n20711 & n20741;
  assign n21133 = n20748 & n21132;
  assign n21134 = n20741 & n20764;
  assign n21135 = n20741 & n20776;
  assign n21136 = ~n21134 & ~n21135;
  assign n21137 = ~n20711 & ~n21136;
  assign n21138 = ~n21133 & ~n21137;
  assign n21139 = n20711 & n20761;
  assign n21140 = ~n20711 & n20743;
  assign n21141 = ~n21139 & ~n21140;
  assign n21142 = ~n20732 & n21141;
  assign n21143 = ~n20762 & n21142;
  assign n21144 = ~n20741 & ~n21143;
  assign n21145 = ~n20711 & n20744;
  assign n21146 = ~n21144 & ~n21145;
  assign n21147 = ~n20711 & n20732;
  assign n21148 = ~n20960 & ~n21147;
  assign n21149 = n21146 & n21148;
  assign n21150 = n21138 & n21149;
  assign n21151 = n20705 & ~n21150;
  assign n21152 = n20741 & ~n20951;
  assign n21153 = ~n21151 & ~n21152;
  assign n21154 = ~n20765 & ~n21147;
  assign n21155 = ~n20741 & ~n21154;
  assign n21156 = n21153 & ~n21155;
  assign n21157 = ~n21131 & n21156;
  assign n21158 = pi0178 & ~n21157;
  assign n21159 = ~pi0178 & n21157;
  assign po0219 = n21158 | n21159;
  assign n21161 = ~n20584 & n20856;
  assign n21162 = ~n20578 & n20639;
  assign n21163 = ~n21161 & ~n21162;
  assign n21164 = ~n20844 & n21163;
  assign n21165 = n20578 & n20614;
  assign n21166 = ~n20578 & n20589;
  assign n21167 = ~n20606 & ~n21166;
  assign n21168 = n20584 & ~n21167;
  assign n21169 = ~n21165 & ~n21168;
  assign n21170 = n21164 & n21169;
  assign n21171 = ~n20553 & ~n21170;
  assign n21172 = ~n20584 & n20854;
  assign n21173 = ~n20603 & ~n20629;
  assign n21174 = ~n20597 & n21173;
  assign n21175 = ~n21172 & n21174;
  assign n21176 = n20553 & ~n21175;
  assign n21177 = n20553 & n20584;
  assign n21178 = ~n20565 & ~n20578;
  assign n21179 = n20559 & n21178;
  assign n21180 = ~n20571 & n21179;
  assign n21181 = ~n20856 & ~n21180;
  assign n21182 = ~n20610 & n21181;
  assign n21183 = n21177 & ~n21182;
  assign n21184 = ~n21176 & ~n21183;
  assign n21185 = n20607 & n20616;
  assign n21186 = n20578 & n20610;
  assign n21187 = ~n20845 & ~n21186;
  assign n21188 = n20584 & ~n21187;
  assign n21189 = ~n21185 & ~n21188;
  assign n21190 = ~n20631 & n21189;
  assign n21191 = n20578 & n21161;
  assign n21192 = n21190 & ~n21191;
  assign n21193 = n21184 & n21192;
  assign n21194 = ~n21171 & n21193;
  assign n21195 = ~pi0194 & n21194;
  assign n21196 = pi0194 & ~n21194;
  assign po0220 = n21195 | n21196;
  assign n21198 = n20992 & ~n21018;
  assign n21199 = ~n21004 & n21198;
  assign n21200 = ~n21028 & ~n21056;
  assign n21201 = ~n21199 & n21200;
  assign n21202 = ~n21012 & ~n21053;
  assign n21203 = ~n21201 & n21202;
  assign n21204 = n21018 & ~n21053;
  assign n21205 = n21070 & n21204;
  assign n21206 = ~n20992 & ~n21004;
  assign n21207 = ~n21033 & ~n21206;
  assign n21208 = n21012 & ~n21207;
  assign n21209 = n21012 & n21060;
  assign n21210 = ~n21208 & ~n21209;
  assign n21211 = ~n21053 & ~n21210;
  assign n21212 = ~n21205 & ~n21211;
  assign n21213 = ~n20992 & n21018;
  assign n21214 = ~n21004 & n21213;
  assign n21215 = ~n21018 & n21037;
  assign n21216 = ~n20992 & n21215;
  assign n21217 = ~n21214 & ~n21216;
  assign n21218 = n21012 & ~n21217;
  assign n21219 = n21212 & ~n21218;
  assign n21220 = n20992 & n21018;
  assign n21221 = n21004 & n21220;
  assign n21222 = ~n20998 & n21221;
  assign n21223 = ~n21012 & n21018;
  assign n21224 = n21005 & n21223;
  assign n21225 = n20992 & n21224;
  assign n21226 = ~n21038 & n21213;
  assign n21227 = ~n21225 & ~n21226;
  assign n21228 = ~n21222 & n21227;
  assign n21229 = ~n21038 & n21198;
  assign n21230 = ~n21029 & ~n21229;
  assign n21231 = n20992 & n20998;
  assign n21232 = n21019 & n21231;
  assign n21233 = ~n21027 & ~n21232;
  assign n21234 = n21230 & n21233;
  assign n21235 = n21228 & n21234;
  assign n21236 = n21053 & ~n21235;
  assign n21237 = n21219 & ~n21236;
  assign n21238 = ~n21203 & n21237;
  assign n21239 = ~pi0199 & ~n21238;
  assign n21240 = pi0199 & n21219;
  assign n21241 = ~n21203 & n21240;
  assign n21242 = ~n21236 & n21241;
  assign po0221 = n21239 | n21242;
  assign n21244 = ~n20992 & ~n20998;
  assign n21245 = ~n21012 & n21244;
  assign n21246 = n21018 & n21245;
  assign n21247 = ~n21025 & ~n21215;
  assign n21248 = ~n21056 & n21247;
  assign n21249 = ~n21012 & ~n21248;
  assign n21250 = ~n20992 & n21036;
  assign n21251 = ~n21006 & ~n21250;
  assign n21252 = n21012 & ~n21251;
  assign n21253 = ~n21249 & ~n21252;
  assign n21254 = ~n21209 & ~n21216;
  assign n21255 = n21253 & n21254;
  assign n21256 = n21053 & ~n21255;
  assign n21257 = n21006 & n21018;
  assign n21258 = ~n21018 & n21021;
  assign n21259 = ~n21067 & ~n21258;
  assign n21260 = ~n21012 & ~n21259;
  assign n21261 = ~n21257 & ~n21260;
  assign n21262 = n21012 & n21070;
  assign n21263 = n21200 & ~n21262;
  assign n21264 = ~n21025 & n21263;
  assign n21265 = ~n21018 & ~n21264;
  assign n21266 = n21261 & ~n21265;
  assign n21267 = ~n21053 & ~n21266;
  assign n21268 = ~n21256 & ~n21267;
  assign n21269 = ~n21246 & n21268;
  assign n21270 = ~n20992 & n21067;
  assign n21271 = ~n21222 & ~n21270;
  assign n21272 = n21012 & ~n21271;
  assign n21273 = n21269 & ~n21272;
  assign n21274 = ~pi0183 & ~n21273;
  assign n21275 = n21268 & ~n21272;
  assign n21276 = pi0183 & n21275;
  assign n21277 = ~n21246 & n21276;
  assign po0222 = n21274 | n21277;
  assign n21279 = ~n21067 & ~n21069;
  assign n21280 = n21012 & ~n21279;
  assign n21281 = ~n21023 & ~n21280;
  assign n21282 = ~n21053 & ~n21281;
  assign n21283 = ~n21036 & n21220;
  assign n21284 = ~n21053 & n21283;
  assign n21285 = n21012 & n21213;
  assign n21286 = n21036 & n21285;
  assign n21287 = n20992 & n21223;
  assign n21288 = n21004 & n21287;
  assign n21289 = ~n21286 & ~n21288;
  assign n21290 = ~n21284 & n21289;
  assign n21291 = ~n21036 & ~n21244;
  assign n21292 = ~n21018 & ~n21291;
  assign n21293 = ~n21006 & ~n21292;
  assign n21294 = ~n21012 & ~n21293;
  assign n21295 = ~n21061 & ~n21294;
  assign n21296 = n21018 & n21025;
  assign n21297 = n21004 & n21198;
  assign n21298 = n21018 & ~n21291;
  assign n21299 = ~n21297 & ~n21298;
  assign n21300 = n21012 & ~n21299;
  assign n21301 = ~n21296 & ~n21300;
  assign n21302 = n21295 & n21301;
  assign n21303 = n21053 & ~n21302;
  assign n21304 = ~n21031 & ~n21070;
  assign n21305 = n21202 & ~n21304;
  assign n21306 = ~n21303 & ~n21305;
  assign n21307 = n21290 & n21306;
  assign n21308 = ~n21282 & n21307;
  assign n21309 = pi0187 & ~n21308;
  assign n21310 = ~pi0187 & n21308;
  assign po0223 = n21309 | n21310;
  assign n21312 = ~n20083 & n20139;
  assign n21313 = n20102 & n20124;
  assign n21314 = ~n20123 & ~n21313;
  assign n21315 = ~n20083 & ~n21314;
  assign n21316 = n20083 & ~n20310;
  assign n21317 = ~n21315 & ~n21316;
  assign n21318 = ~n20327 & n21317;
  assign n21319 = n20120 & ~n21318;
  assign n21320 = ~n21312 & ~n21319;
  assign n21321 = ~n20108 & n20285;
  assign n21322 = ~n20297 & ~n21321;
  assign n21323 = ~n20089 & ~n21322;
  assign n21324 = ~n20110 & ~n21323;
  assign n21325 = ~n20298 & n21324;
  assign n21326 = ~n20102 & n20142;
  assign n21327 = n20083 & n20125;
  assign n21328 = ~n21326 & ~n21327;
  assign n21329 = n21325 & n21328;
  assign n21330 = ~n20120 & ~n21329;
  assign n21331 = ~n20884 & ~n20898;
  assign n21332 = n20083 & ~n21331;
  assign n21333 = ~n21330 & ~n21332;
  assign n21334 = n21320 & n21333;
  assign n21335 = ~pi0210 & ~n21334;
  assign n21336 = pi0210 & n21320;
  assign n21337 = n21333 & n21336;
  assign po0224 = n21335 | n21337;
  assign n21339 = ~n20952 & ~n21147;
  assign n21340 = ~n21127 & n21339;
  assign n21341 = n20741 & ~n21340;
  assign n21342 = ~n20962 & ~n20979;
  assign n21343 = ~n20960 & ~n21135;
  assign n21344 = ~n20948 & ~n21140;
  assign n21345 = ~n20741 & ~n21344;
  assign n21346 = ~n20770 & ~n21345;
  assign n21347 = n21343 & n21346;
  assign n21348 = n20705 & ~n21347;
  assign n21349 = n20724 & n20730;
  assign n21350 = ~n20749 & ~n21349;
  assign n21351 = n20711 & ~n21350;
  assign n21352 = ~n20732 & ~n20965;
  assign n21353 = ~n20741 & ~n21352;
  assign n21354 = n20711 & n20730;
  assign n21355 = ~n20744 & ~n21354;
  assign n21356 = ~n20752 & n21355;
  assign n21357 = n20741 & ~n21356;
  assign n21358 = ~n21353 & ~n21357;
  assign n21359 = ~n21351 & n21358;
  assign n21360 = ~n20705 & ~n21359;
  assign n21361 = ~n21348 & ~n21360;
  assign n21362 = n21342 & n21361;
  assign n21363 = ~n21341 & n21362;
  assign n21364 = ~pi0188 & ~n21363;
  assign n21365 = pi0188 & n21342;
  assign n21366 = ~n21341 & n21365;
  assign n21367 = n21361 & n21366;
  assign po0225 = n21364 | n21367;
  assign n21369 = pi3153 & ~pi9040;
  assign n21370 = pi3115 & pi9040;
  assign n21371 = ~n21369 & ~n21370;
  assign n21372 = ~pi0211 & ~n21371;
  assign n21373 = pi0211 & n21371;
  assign n21374 = ~n21372 & ~n21373;
  assign n21375 = pi3188 & pi9040;
  assign n21376 = pi3110 & ~pi9040;
  assign n21377 = ~n21375 & ~n21376;
  assign n21378 = ~pi0209 & n21377;
  assign n21379 = pi0209 & ~n21377;
  assign n21380 = ~n21378 & ~n21379;
  assign n21381 = pi3172 & pi9040;
  assign n21382 = pi3228 & ~pi9040;
  assign n21383 = ~n21381 & ~n21382;
  assign n21384 = pi0201 & n21383;
  assign n21385 = ~pi0201 & ~n21383;
  assign n21386 = ~n21384 & ~n21385;
  assign n21387 = pi3104 & pi9040;
  assign n21388 = pi3115 & ~pi9040;
  assign n21389 = ~n21387 & ~n21388;
  assign n21390 = ~pi0216 & n21389;
  assign n21391 = pi0216 & ~n21389;
  assign n21392 = ~n21390 & ~n21391;
  assign n21393 = pi3116 & pi9040;
  assign n21394 = pi3172 & ~pi9040;
  assign n21395 = ~n21393 & ~n21394;
  assign n21396 = ~pi0177 & ~n21395;
  assign n21397 = pi0177 & ~n21393;
  assign n21398 = ~n21394 & n21397;
  assign n21399 = ~n21396 & ~n21398;
  assign n21400 = ~n21392 & ~n21399;
  assign n21401 = n21386 & n21400;
  assign n21402 = pi3089 & pi9040;
  assign n21403 = pi3169 & ~pi9040;
  assign n21404 = ~n21402 & ~n21403;
  assign n21405 = ~pi0196 & n21404;
  assign n21406 = pi0196 & ~n21404;
  assign n21407 = ~n21405 & ~n21406;
  assign n21408 = n21399 & ~n21407;
  assign n21409 = ~n21392 & n21408;
  assign n21410 = ~n21401 & ~n21409;
  assign n21411 = n21399 & n21407;
  assign n21412 = n21392 & n21411;
  assign n21413 = ~n21386 & n21412;
  assign n21414 = n21410 & ~n21413;
  assign n21415 = ~n21380 & ~n21414;
  assign n21416 = n21392 & n21399;
  assign n21417 = ~n21386 & n21416;
  assign n21418 = ~n21407 & n21417;
  assign n21419 = ~n21399 & ~n21407;
  assign n21420 = ~n21392 & n21419;
  assign n21421 = ~n21386 & n21420;
  assign n21422 = n21392 & ~n21399;
  assign n21423 = ~n21411 & ~n21422;
  assign n21424 = n21386 & ~n21423;
  assign n21425 = ~n21421 & ~n21424;
  assign n21426 = ~n21418 & n21425;
  assign n21427 = n21380 & ~n21426;
  assign n21428 = ~n21415 & ~n21427;
  assign n21429 = n21374 & ~n21428;
  assign n21430 = ~n21380 & ~n21386;
  assign n21431 = ~n21399 & n21430;
  assign n21432 = n21380 & ~n21386;
  assign n21433 = n21411 & n21432;
  assign n21434 = ~n21386 & ~n21392;
  assign n21435 = n21399 & n21434;
  assign n21436 = ~n21401 & ~n21435;
  assign n21437 = n21380 & ~n21436;
  assign n21438 = ~n21433 & ~n21437;
  assign n21439 = ~n21392 & n21411;
  assign n21440 = ~n21386 & n21439;
  assign n21441 = ~n21407 & n21416;
  assign n21442 = n21386 & n21441;
  assign n21443 = ~n21440 & ~n21442;
  assign n21444 = ~n21380 & n21386;
  assign n21445 = n21416 & n21444;
  assign n21446 = n21392 & n21419;
  assign n21447 = ~n21380 & n21446;
  assign n21448 = ~n21445 & ~n21447;
  assign n21449 = n21443 & n21448;
  assign n21450 = n21438 & n21449;
  assign n21451 = ~n21431 & n21450;
  assign n21452 = ~n21374 & ~n21451;
  assign n21453 = ~n21399 & n21407;
  assign n21454 = n21392 & n21453;
  assign n21455 = n21432 & n21454;
  assign n21456 = ~n21392 & n21433;
  assign n21457 = ~n21455 & ~n21456;
  assign n21458 = ~n21386 & n21392;
  assign n21459 = ~n21407 & n21458;
  assign n21460 = ~n21399 & n21459;
  assign n21461 = ~n21380 & n21460;
  assign n21462 = n21457 & ~n21461;
  assign n21463 = n21386 & n21408;
  assign n21464 = ~n21392 & n21453;
  assign n21465 = ~n21386 & n21464;
  assign n21466 = ~n21463 & ~n21465;
  assign n21467 = ~n21380 & ~n21466;
  assign n21468 = n21462 & ~n21467;
  assign n21469 = ~n21452 & n21468;
  assign n21470 = ~n21429 & n21469;
  assign n21471 = ~pi0233 & ~n21470;
  assign n21472 = pi0233 & n21470;
  assign po0236 = n21471 | n21472;
  assign n21474 = ~n21374 & n21380;
  assign n21475 = ~n21386 & n21400;
  assign n21476 = n21386 & n21439;
  assign n21477 = ~n21386 & n21408;
  assign n21478 = ~n21476 & ~n21477;
  assign n21479 = ~n21475 & n21478;
  assign n21480 = n21474 & ~n21479;
  assign n21481 = n21407 & n21458;
  assign n21482 = n21386 & n21464;
  assign n21483 = ~n21481 & ~n21482;
  assign n21484 = ~n21409 & ~n21412;
  assign n21485 = n21483 & n21484;
  assign n21486 = ~n21380 & ~n21485;
  assign n21487 = n21386 & n21446;
  assign n21488 = ~n21486 & ~n21487;
  assign n21489 = ~n21374 & ~n21488;
  assign n21490 = ~n21480 & ~n21489;
  assign n21491 = ~n21392 & n21430;
  assign n21492 = ~n21407 & n21491;
  assign n21493 = ~n21413 & ~n21492;
  assign n21494 = ~n21408 & ~n21453;
  assign n21495 = n21386 & ~n21494;
  assign n21496 = ~n21454 & ~n21495;
  assign n21497 = n21380 & ~n21496;
  assign n21498 = ~n21420 & ~n21475;
  assign n21499 = ~n21476 & n21498;
  assign n21500 = ~n21380 & ~n21499;
  assign n21501 = ~n21497 & ~n21500;
  assign n21502 = n21386 & n21392;
  assign n21503 = n21407 & n21502;
  assign n21504 = ~n21399 & n21503;
  assign n21505 = ~n21442 & ~n21504;
  assign n21506 = ~n21460 & n21505;
  assign n21507 = ~n21433 & n21506;
  assign n21508 = n21501 & n21507;
  assign n21509 = n21374 & ~n21508;
  assign n21510 = n21493 & ~n21509;
  assign n21511 = n21490 & n21510;
  assign n21512 = pi0234 & ~n21511;
  assign n21513 = ~pi0234 & n21493;
  assign n21514 = n21490 & n21513;
  assign n21515 = ~n21509 & n21514;
  assign po0237 = n21512 | n21515;
  assign n21517 = ~n21420 & ~n21454;
  assign n21518 = n21380 & ~n21517;
  assign n21519 = n21386 & n21409;
  assign n21520 = ~n21518 & ~n21519;
  assign n21521 = n21386 & n21399;
  assign n21522 = ~n21416 & ~n21521;
  assign n21523 = ~n21464 & n21522;
  assign n21524 = ~n21380 & ~n21523;
  assign n21525 = n21520 & ~n21524;
  assign n21526 = ~n21374 & ~n21525;
  assign n21527 = ~n21386 & n21441;
  assign n21528 = n21380 & n21527;
  assign n21529 = ~n21456 & ~n21528;
  assign n21530 = ~n21461 & n21529;
  assign n21531 = ~n21380 & n21399;
  assign n21532 = n21434 & n21531;
  assign n21533 = n21386 & n21420;
  assign n21534 = n21380 & n21416;
  assign n21535 = ~n21533 & ~n21534;
  assign n21536 = ~n21504 & n21535;
  assign n21537 = ~n21532 & n21536;
  assign n21538 = n21407 & n21434;
  assign n21539 = ~n21460 & ~n21538;
  assign n21540 = n21537 & n21539;
  assign n21541 = ~n21447 & n21540;
  assign n21542 = n21374 & ~n21541;
  assign n21543 = n21530 & ~n21542;
  assign n21544 = ~n21526 & n21543;
  assign n21545 = ~pi0241 & ~n21544;
  assign n21546 = pi0241 & n21530;
  assign n21547 = ~n21526 & n21546;
  assign n21548 = ~n21542 & n21547;
  assign po0242 = n21545 | n21548;
  assign n21550 = pi3078 & pi9040;
  assign n21551 = pi3160 & ~pi9040;
  assign n21552 = ~n21550 & ~n21551;
  assign n21553 = ~pi0218 & n21552;
  assign n21554 = pi0218 & ~n21552;
  assign n21555 = ~n21553 & ~n21554;
  assign n21556 = pi3088 & pi9040;
  assign n21557 = pi3108 & ~pi9040;
  assign n21558 = ~n21556 & ~n21557;
  assign n21559 = pi0184 & n21558;
  assign n21560 = ~pi0184 & ~n21558;
  assign n21561 = ~n21559 & ~n21560;
  assign n21562 = pi3160 & pi9040;
  assign n21563 = pi3113 & ~pi9040;
  assign n21564 = ~n21562 & ~n21563;
  assign n21565 = pi0196 & n21564;
  assign n21566 = ~pi0196 & ~n21564;
  assign n21567 = ~n21565 & ~n21566;
  assign n21568 = pi3228 & pi9040;
  assign n21569 = pi3077 & ~pi9040;
  assign n21570 = ~n21568 & ~n21569;
  assign n21571 = ~pi0211 & n21570;
  assign n21572 = pi0211 & ~n21570;
  assign n21573 = ~n21571 & ~n21572;
  assign n21574 = n21567 & n21573;
  assign n21575 = ~n21561 & n21574;
  assign n21576 = n21567 & ~n21573;
  assign n21577 = n21561 & n21576;
  assign n21578 = ~n21575 & ~n21577;
  assign n21579 = n21555 & ~n21578;
  assign n21580 = pi3074 & pi9040;
  assign n21581 = pi3084 & ~pi9040;
  assign n21582 = ~n21580 & ~n21581;
  assign n21583 = pi0207 & n21582;
  assign n21584 = ~pi0207 & ~n21582;
  assign n21585 = ~n21583 & ~n21584;
  assign n21586 = pi3137 & pi9040;
  assign n21587 = pi3180 & ~pi9040;
  assign n21588 = ~n21586 & ~n21587;
  assign n21589 = ~pi0182 & ~n21588;
  assign n21590 = pi0182 & n21588;
  assign n21591 = ~n21589 & ~n21590;
  assign n21592 = n21573 & n21591;
  assign n21593 = n21555 & ~n21561;
  assign n21594 = n21592 & n21593;
  assign n21595 = ~n21567 & ~n21573;
  assign n21596 = ~n21555 & ~n21561;
  assign n21597 = n21595 & n21596;
  assign n21598 = ~n21573 & ~n21591;
  assign n21599 = n21567 & n21598;
  assign n21600 = n21561 & ~n21567;
  assign n21601 = ~n21591 & n21600;
  assign n21602 = n21573 & n21601;
  assign n21603 = ~n21599 & ~n21602;
  assign n21604 = ~n21573 & n21591;
  assign n21605 = n21561 & n21604;
  assign n21606 = n21603 & ~n21605;
  assign n21607 = n21555 & ~n21606;
  assign n21608 = ~n21597 & ~n21607;
  assign n21609 = ~n21594 & n21608;
  assign n21610 = n21567 & n21604;
  assign n21611 = n21561 & n21610;
  assign n21612 = ~n21567 & n21598;
  assign n21613 = ~n21561 & n21612;
  assign n21614 = n21567 & n21592;
  assign n21615 = ~n21561 & n21614;
  assign n21616 = ~n21613 & ~n21615;
  assign n21617 = ~n21611 & n21616;
  assign n21618 = n21609 & n21617;
  assign n21619 = ~n21585 & ~n21618;
  assign n21620 = ~n21561 & ~n21567;
  assign n21621 = n21591 & n21620;
  assign n21622 = ~n21573 & n21621;
  assign n21623 = ~n21614 & ~n21622;
  assign n21624 = n21555 & ~n21623;
  assign n21625 = ~n21591 & n21620;
  assign n21626 = n21573 & n21625;
  assign n21627 = ~n21567 & n21592;
  assign n21628 = n21561 & n21627;
  assign n21629 = ~n21626 & ~n21628;
  assign n21630 = ~n21573 & n21600;
  assign n21631 = ~n21561 & n21610;
  assign n21632 = ~n21630 & ~n21631;
  assign n21633 = ~n21555 & ~n21632;
  assign n21634 = n21629 & ~n21633;
  assign n21635 = ~n21624 & n21634;
  assign n21636 = n21585 & ~n21635;
  assign n21637 = ~n21567 & ~n21591;
  assign n21638 = ~n21555 & n21637;
  assign n21639 = ~n21561 & n21638;
  assign n21640 = n21573 & ~n21591;
  assign n21641 = n21567 & n21640;
  assign n21642 = n21561 & n21641;
  assign n21643 = ~n21612 & ~n21642;
  assign n21644 = ~n21628 & n21643;
  assign n21645 = ~n21555 & ~n21644;
  assign n21646 = ~n21639 & ~n21645;
  assign n21647 = ~n21636 & n21646;
  assign n21648 = ~n21619 & n21647;
  assign n21649 = ~n21579 & n21648;
  assign n21650 = ~pi0225 & ~n21649;
  assign n21651 = pi0225 & n21649;
  assign po0244 = n21650 | n21651;
  assign n21653 = ~n21386 & ~n21399;
  assign n21654 = ~n21538 & ~n21653;
  assign n21655 = n21380 & ~n21654;
  assign n21656 = n21386 & ~n21392;
  assign n21657 = ~n21407 & n21656;
  assign n21658 = ~n21655 & ~n21657;
  assign n21659 = ~n21380 & n21408;
  assign n21660 = ~n21386 & n21659;
  assign n21661 = ~n21465 & ~n21660;
  assign n21662 = n21658 & n21661;
  assign n21663 = n21374 & ~n21662;
  assign n21664 = ~n21439 & ~n21442;
  assign n21665 = ~n21386 & n21419;
  assign n21666 = n21664 & ~n21665;
  assign n21667 = ~n21380 & ~n21666;
  assign n21668 = n21408 & n21432;
  assign n21669 = ~n21413 & ~n21668;
  assign n21670 = ~n21667 & n21669;
  assign n21671 = ~n21464 & ~n21487;
  assign n21672 = n21380 & ~n21671;
  assign n21673 = n21670 & ~n21672;
  assign n21674 = ~n21374 & ~n21673;
  assign n21675 = ~n21663 & ~n21674;
  assign n21676 = ~n21386 & n21453;
  assign n21677 = n21386 & ~n21484;
  assign n21678 = ~n21676 & ~n21677;
  assign n21679 = n21380 & ~n21678;
  assign n21680 = ~n21439 & n21517;
  assign n21681 = n21444 & ~n21680;
  assign n21682 = ~n21679 & ~n21681;
  assign n21683 = n21675 & n21682;
  assign n21684 = ~pi0236 & ~n21683;
  assign n21685 = ~n21674 & n21682;
  assign n21686 = pi0236 & n21685;
  assign n21687 = ~n21663 & n21686;
  assign po0249 = n21684 | n21687;
  assign n21689 = pi3069 & pi9040;
  assign n21690 = pi3107 & ~pi9040;
  assign n21691 = ~n21689 & ~n21690;
  assign n21692 = pi0202 & n21691;
  assign n21693 = ~pi0202 & ~n21691;
  assign n21694 = ~n21692 & ~n21693;
  assign n21695 = pi3113 & pi9040;
  assign n21696 = pi3076 & ~pi9040;
  assign n21697 = ~n21695 & ~n21696;
  assign n21698 = ~pi0182 & n21697;
  assign n21699 = pi0182 & ~n21697;
  assign n21700 = ~n21698 & ~n21699;
  assign n21701 = pi3108 & pi9040;
  assign n21702 = pi3137 & ~pi9040;
  assign n21703 = ~n21701 & ~n21702;
  assign n21704 = ~pi0193 & n21703;
  assign n21705 = pi0193 & ~n21703;
  assign n21706 = ~n21704 & ~n21705;
  assign n21707 = pi3180 & pi9040;
  assign n21708 = pi3088 & ~pi9040;
  assign n21709 = ~n21707 & ~n21708;
  assign n21710 = ~pi0207 & n21709;
  assign n21711 = pi0207 & ~n21709;
  assign n21712 = ~n21710 & ~n21711;
  assign n21713 = ~n21706 & ~n21712;
  assign n21714 = n21700 & n21713;
  assign n21715 = pi3070 & pi9040;
  assign n21716 = pi3080 & ~pi9040;
  assign n21717 = ~n21715 & ~n21716;
  assign n21718 = pi0212 & n21717;
  assign n21719 = ~pi0212 & ~n21717;
  assign n21720 = ~n21718 & ~n21719;
  assign n21721 = n21714 & ~n21720;
  assign n21722 = n21706 & n21712;
  assign n21723 = n21700 & n21722;
  assign n21724 = ~n21720 & n21723;
  assign n21725 = ~n21721 & ~n21724;
  assign n21726 = ~n21700 & n21720;
  assign n21727 = n21722 & n21726;
  assign n21728 = ~n21706 & n21712;
  assign n21729 = n21700 & n21728;
  assign n21730 = n21720 & n21729;
  assign n21731 = ~n21727 & ~n21730;
  assign n21732 = n21725 & n21731;
  assign n21733 = n21694 & ~n21732;
  assign n21734 = n21706 & ~n21712;
  assign n21735 = n21700 & n21734;
  assign n21736 = n21720 & n21735;
  assign n21737 = ~n21729 & ~n21736;
  assign n21738 = n21694 & ~n21737;
  assign n21739 = ~n21712 & ~n21720;
  assign n21740 = ~n21694 & n21739;
  assign n21741 = ~n21700 & ~n21706;
  assign n21742 = n21720 & n21722;
  assign n21743 = ~n21741 & ~n21742;
  assign n21744 = ~n21694 & ~n21743;
  assign n21745 = ~n21740 & ~n21744;
  assign n21746 = ~n21700 & n21734;
  assign n21747 = ~n21720 & n21746;
  assign n21748 = n21745 & ~n21747;
  assign n21749 = ~n21712 & n21741;
  assign n21750 = n21720 & n21749;
  assign n21751 = n21748 & ~n21750;
  assign n21752 = ~n21738 & n21751;
  assign n21753 = pi3107 & pi9040;
  assign n21754 = pi3070 & ~pi9040;
  assign n21755 = ~n21753 & ~n21754;
  assign n21756 = ~pi0223 & ~n21755;
  assign n21757 = pi0223 & n21755;
  assign n21758 = ~n21756 & ~n21757;
  assign n21759 = ~n21752 & ~n21758;
  assign n21760 = n21700 & ~n21712;
  assign n21761 = ~n21694 & n21720;
  assign n21762 = n21758 & n21761;
  assign n21763 = n21760 & n21762;
  assign n21764 = n21700 & ~n21720;
  assign n21765 = n21712 & n21764;
  assign n21766 = ~n21694 & ~n21765;
  assign n21767 = n21706 & n21726;
  assign n21768 = ~n21713 & ~n21760;
  assign n21769 = ~n21720 & ~n21768;
  assign n21770 = ~n21700 & n21722;
  assign n21771 = n21694 & ~n21770;
  assign n21772 = ~n21769 & n21771;
  assign n21773 = ~n21767 & n21772;
  assign n21774 = ~n21766 & ~n21773;
  assign n21775 = ~n21700 & n21728;
  assign n21776 = n21720 & n21775;
  assign n21777 = ~n21774 & ~n21776;
  assign n21778 = n21758 & ~n21777;
  assign n21779 = ~n21763 & ~n21778;
  assign n21780 = ~n21759 & n21779;
  assign n21781 = ~n21733 & n21780;
  assign n21782 = ~n21694 & ~n21720;
  assign n21783 = n21734 & n21782;
  assign n21784 = ~n21700 & n21783;
  assign n21785 = n21781 & ~n21784;
  assign n21786 = pi0227 & ~n21785;
  assign n21787 = n21780 & ~n21784;
  assign n21788 = ~pi0227 & n21787;
  assign n21789 = ~n21733 & n21788;
  assign po0250 = n21786 | n21789;
  assign n21791 = ~n21573 & n21601;
  assign n21792 = ~n21576 & ~n21626;
  assign n21793 = ~n21555 & ~n21792;
  assign n21794 = ~n21791 & ~n21793;
  assign n21795 = ~n21622 & n21794;
  assign n21796 = n21555 & n21561;
  assign n21797 = n21627 & n21796;
  assign n21798 = ~n21615 & ~n21797;
  assign n21799 = ~n21642 & n21798;
  assign n21800 = n21795 & n21799;
  assign n21801 = n21585 & ~n21800;
  assign n21802 = ~n21567 & n21604;
  assign n21803 = n21561 & n21802;
  assign n21804 = ~n21602 & ~n21803;
  assign n21805 = ~n21561 & n21641;
  assign n21806 = ~n21613 & ~n21805;
  assign n21807 = ~n21555 & n21627;
  assign n21808 = n21561 & n21614;
  assign n21809 = ~n21807 & ~n21808;
  assign n21810 = n21567 & n21591;
  assign n21811 = n21561 & ~n21573;
  assign n21812 = ~n21810 & ~n21811;
  assign n21813 = ~n21637 & n21812;
  assign n21814 = n21555 & ~n21813;
  assign n21815 = n21809 & ~n21814;
  assign n21816 = n21806 & n21815;
  assign n21817 = n21804 & n21816;
  assign n21818 = ~n21585 & ~n21817;
  assign n21819 = ~n21801 & ~n21818;
  assign n21820 = pi0224 & ~n21819;
  assign n21821 = ~pi0224 & ~n21801;
  assign n21822 = ~n21818 & n21821;
  assign po0252 = n21820 | n21822;
  assign n21824 = pi3075 & pi9040;
  assign n21825 = pi3091 & ~pi9040;
  assign n21826 = ~n21824 & ~n21825;
  assign n21827 = ~pi0220 & n21826;
  assign n21828 = pi0220 & ~n21826;
  assign n21829 = ~n21827 & ~n21828;
  assign n21830 = pi3109 & pi9040;
  assign n21831 = pi3157 & ~pi9040;
  assign n21832 = ~n21830 & ~n21831;
  assign n21833 = pi0198 & n21832;
  assign n21834 = ~pi0198 & ~n21832;
  assign n21835 = ~n21833 & ~n21834;
  assign n21836 = pi3111 & pi9040;
  assign n21837 = pi3109 & ~pi9040;
  assign n21838 = ~n21836 & ~n21837;
  assign n21839 = ~pi0214 & n21838;
  assign n21840 = pi0214 & ~n21838;
  assign n21841 = ~n21839 & ~n21840;
  assign n21842 = n21835 & n21841;
  assign n21843 = pi3083 & pi9040;
  assign n21844 = pi3118 & ~pi9040;
  assign n21845 = ~n21843 & ~n21844;
  assign n21846 = pi0219 & n21845;
  assign n21847 = ~pi0219 & ~n21845;
  assign n21848 = ~n21846 & ~n21847;
  assign n21849 = pi3163 & pi9040;
  assign n21850 = pi3085 & ~pi9040;
  assign n21851 = ~n21849 & ~n21850;
  assign n21852 = ~pi0180 & ~n21851;
  assign n21853 = pi0180 & n21851;
  assign n21854 = ~n21852 & ~n21853;
  assign n21855 = n21848 & n21854;
  assign n21856 = n21842 & n21855;
  assign n21857 = n21848 & ~n21854;
  assign n21858 = ~n21835 & n21857;
  assign n21859 = ~n21856 & ~n21858;
  assign n21860 = n21829 & ~n21859;
  assign n21861 = pi3085 & pi9040;
  assign n21862 = pi3081 & ~pi9040;
  assign n21863 = ~n21861 & ~n21862;
  assign n21864 = ~pi0205 & ~n21863;
  assign n21865 = pi0205 & n21863;
  assign n21866 = ~n21864 & ~n21865;
  assign n21867 = ~n21829 & ~n21848;
  assign n21868 = n21835 & n21867;
  assign n21869 = n21842 & ~n21854;
  assign n21870 = n21835 & ~n21841;
  assign n21871 = n21854 & n21870;
  assign n21872 = ~n21869 & ~n21871;
  assign n21873 = ~n21835 & n21841;
  assign n21874 = n21854 & n21873;
  assign n21875 = n21848 & n21874;
  assign n21876 = n21872 & ~n21875;
  assign n21877 = ~n21829 & ~n21876;
  assign n21878 = ~n21868 & ~n21877;
  assign n21879 = ~n21835 & ~n21841;
  assign n21880 = ~n21854 & n21879;
  assign n21881 = n21848 & n21880;
  assign n21882 = n21878 & ~n21881;
  assign n21883 = ~n21848 & n21873;
  assign n21884 = ~n21835 & n21854;
  assign n21885 = ~n21841 & n21884;
  assign n21886 = ~n21883 & ~n21885;
  assign n21887 = n21829 & ~n21886;
  assign n21888 = ~n21854 & n21870;
  assign n21889 = ~n21848 & n21888;
  assign n21890 = ~n21887 & ~n21889;
  assign n21891 = n21882 & n21890;
  assign n21892 = n21866 & ~n21891;
  assign n21893 = ~n21860 & ~n21892;
  assign n21894 = ~n21829 & ~n21866;
  assign n21895 = ~n21886 & n21894;
  assign n21896 = ~n21854 & n21873;
  assign n21897 = ~n21888 & ~n21896;
  assign n21898 = n21848 & ~n21897;
  assign n21899 = ~n21856 & ~n21898;
  assign n21900 = ~n21866 & ~n21899;
  assign n21901 = ~n21895 & ~n21900;
  assign n21902 = n21829 & ~n21866;
  assign n21903 = n21842 & ~n21848;
  assign n21904 = ~n21880 & ~n21903;
  assign n21905 = n21835 & n21854;
  assign n21906 = n21904 & ~n21905;
  assign n21907 = n21902 & ~n21906;
  assign n21908 = n21901 & ~n21907;
  assign n21909 = n21893 & n21908;
  assign n21910 = ~pi0231 & ~n21909;
  assign n21911 = pi0231 & n21901;
  assign n21912 = n21893 & n21911;
  assign n21913 = ~n21907 & n21912;
  assign po0257 = n21910 | n21913;
  assign n21915 = pi3086 & pi9040;
  assign n21916 = pi3121 & ~pi9040;
  assign n21917 = ~n21915 & ~n21916;
  assign n21918 = ~pi0198 & ~n21917;
  assign n21919 = pi0198 & n21917;
  assign n21920 = ~n21918 & ~n21919;
  assign n21921 = pi3112 & pi9040;
  assign n21922 = pi3111 & ~pi9040;
  assign n21923 = ~n21921 & ~n21922;
  assign n21924 = ~pi0193 & n21923;
  assign n21925 = pi0193 & ~n21923;
  assign n21926 = ~n21924 & ~n21925;
  assign n21927 = pi3081 & pi9040;
  assign n21928 = pi3073 & ~pi9040;
  assign n21929 = ~n21927 & ~n21928;
  assign n21930 = ~pi0223 & n21929;
  assign n21931 = pi0223 & ~n21929;
  assign n21932 = ~n21930 & ~n21931;
  assign n21933 = pi3093 & pi9040;
  assign n21934 = pi3225 & ~pi9040;
  assign n21935 = ~n21933 & ~n21934;
  assign n21936 = ~pi0180 & n21935;
  assign n21937 = pi0180 & ~n21935;
  assign n21938 = ~n21936 & ~n21937;
  assign n21939 = n21932 & ~n21938;
  assign n21940 = pi3072 & pi9040;
  assign n21941 = pi3168 & ~pi9040;
  assign n21942 = ~n21940 & ~n21941;
  assign n21943 = pi0208 & n21942;
  assign n21944 = ~pi0208 & ~n21942;
  assign n21945 = ~n21943 & ~n21944;
  assign n21946 = pi3157 & pi9040;
  assign n21947 = pi3112 & ~pi9040;
  assign n21948 = ~n21946 & ~n21947;
  assign n21949 = ~pi0213 & n21948;
  assign n21950 = pi0213 & ~n21948;
  assign n21951 = ~n21949 & ~n21950;
  assign n21952 = n21945 & ~n21951;
  assign n21953 = n21939 & n21952;
  assign n21954 = ~n21926 & n21953;
  assign n21955 = ~n21945 & ~n21951;
  assign n21956 = ~n21932 & ~n21938;
  assign n21957 = n21955 & n21956;
  assign n21958 = n21932 & n21938;
  assign n21959 = ~n21926 & n21958;
  assign n21960 = ~n21945 & n21959;
  assign n21961 = ~n21932 & n21938;
  assign n21962 = ~n21926 & n21961;
  assign n21963 = ~n21951 & n21962;
  assign n21964 = n21945 & n21963;
  assign n21965 = ~n21960 & ~n21964;
  assign n21966 = ~n21957 & n21965;
  assign n21967 = ~n21954 & n21966;
  assign n21968 = n21926 & ~n21945;
  assign n21969 = ~n21938 & n21968;
  assign n21970 = ~n21932 & n21969;
  assign n21971 = n21967 & ~n21970;
  assign n21972 = ~n21920 & ~n21971;
  assign n21973 = n21926 & n21938;
  assign n21974 = ~n21932 & n21973;
  assign n21975 = n21945 & n21951;
  assign n21976 = n21974 & n21975;
  assign n21977 = ~n21926 & ~n21945;
  assign n21978 = n21932 & n21977;
  assign n21979 = ~n21945 & n21958;
  assign n21980 = ~n21978 & ~n21979;
  assign n21981 = n21951 & ~n21980;
  assign n21982 = ~n21976 & ~n21981;
  assign n21983 = ~n21920 & ~n21982;
  assign n21984 = n21938 & n21977;
  assign n21985 = ~n21926 & ~n21932;
  assign n21986 = ~n21938 & n21985;
  assign n21987 = n21945 & n21986;
  assign n21988 = ~n21984 & ~n21987;
  assign n21989 = n21926 & n21939;
  assign n21990 = n21945 & n21989;
  assign n21991 = n21988 & ~n21990;
  assign n21992 = n21951 & ~n21991;
  assign n21993 = ~n21983 & ~n21992;
  assign n21994 = ~n21972 & n21993;
  assign n21995 = n21926 & n21945;
  assign n21996 = ~n21951 & n21995;
  assign n21997 = n21958 & n21996;
  assign n21998 = n21926 & ~n21932;
  assign n21999 = n21955 & n21998;
  assign n22000 = n21951 & n21985;
  assign n22001 = n21932 & n21945;
  assign n22002 = n21926 & n22001;
  assign n22003 = ~n21989 & ~n22002;
  assign n22004 = ~n22000 & n22003;
  assign n22005 = ~n21945 & n21974;
  assign n22006 = n22004 & ~n22005;
  assign n22007 = n21939 & ~n21951;
  assign n22008 = ~n21945 & n22007;
  assign n22009 = n21926 & ~n21938;
  assign n22010 = n21945 & n21958;
  assign n22011 = ~n22009 & ~n22010;
  assign n22012 = ~n21951 & ~n22011;
  assign n22013 = ~n22008 & ~n22012;
  assign n22014 = n22006 & n22013;
  assign n22015 = n21920 & ~n22014;
  assign n22016 = ~n21999 & ~n22015;
  assign n22017 = ~n21997 & n22016;
  assign n22018 = n21994 & n22017;
  assign n22019 = pi0228 & n22018;
  assign n22020 = ~pi0228 & ~n22018;
  assign po0259 = n22019 | n22020;
  assign n22022 = ~n21926 & n21932;
  assign n22023 = ~n21970 & ~n22022;
  assign n22024 = ~n22001 & n22023;
  assign n22025 = ~n21951 & ~n22024;
  assign n22026 = ~n21932 & n21975;
  assign n22027 = ~n21926 & n21945;
  assign n22028 = ~n21938 & n22027;
  assign n22029 = ~n21945 & n21962;
  assign n22030 = ~n22028 & ~n22029;
  assign n22031 = n21926 & n21932;
  assign n22032 = ~n21945 & n21951;
  assign n22033 = n22031 & n22032;
  assign n22034 = n22030 & ~n22033;
  assign n22035 = ~n22026 & n22034;
  assign n22036 = ~n22025 & n22035;
  assign n22037 = n21920 & ~n22036;
  assign n22038 = ~n21926 & n21939;
  assign n22039 = ~n21945 & n22038;
  assign n22040 = n21945 & n21959;
  assign n22041 = ~n22039 & ~n22040;
  assign n22042 = ~n21951 & ~n22041;
  assign n22043 = ~n22037 & ~n22042;
  assign n22044 = n21945 & n21962;
  assign n22045 = ~n21974 & ~n21986;
  assign n22046 = ~n21951 & ~n22045;
  assign n22047 = ~n22044 & ~n22046;
  assign n22048 = ~n21990 & n22047;
  assign n22049 = ~n21920 & ~n22048;
  assign n22050 = ~n21956 & ~n21958;
  assign n22051 = n21926 & ~n22050;
  assign n22052 = ~n21979 & ~n22051;
  assign n22053 = n21951 & ~n22052;
  assign n22054 = ~n21920 & n22053;
  assign n22055 = ~n22049 & ~n22054;
  assign n22056 = n22043 & n22055;
  assign n22057 = pi0229 & ~n22056;
  assign n22058 = ~pi0229 & n22043;
  assign n22059 = n22055 & n22058;
  assign po0261 = n22057 | n22059;
  assign n22061 = pi3184 & pi9040;
  assign n22062 = pi3087 & ~pi9040;
  assign n22063 = ~n22061 & ~n22062;
  assign n22064 = ~pi0215 & n22063;
  assign n22065 = pi0215 & ~n22063;
  assign n22066 = ~n22064 & ~n22065;
  assign n22067 = pi3091 & pi9040;
  assign n22068 = pi3184 & ~pi9040;
  assign n22069 = ~n22067 & ~n22068;
  assign n22070 = ~pi0206 & n22069;
  assign n22071 = pi0206 & ~n22069;
  assign n22072 = ~n22070 & ~n22071;
  assign n22073 = pi3073 & pi9040;
  assign n22074 = pi3163 & ~pi9040;
  assign n22075 = ~n22073 & ~n22074;
  assign n22076 = ~pi0217 & ~n22075;
  assign n22077 = pi0217 & n22075;
  assign n22078 = ~n22076 & ~n22077;
  assign n22079 = pi3122 & pi9040;
  assign n22080 = pi3079 & ~pi9040;
  assign n22081 = ~n22079 & ~n22080;
  assign n22082 = ~pi0203 & ~n22081;
  assign n22083 = pi0203 & n22081;
  assign n22084 = ~n22082 & ~n22083;
  assign n22085 = pi3071 & pi9040;
  assign n22086 = pi3082 & ~pi9040;
  assign n22087 = ~n22085 & ~n22086;
  assign n22088 = ~pi0204 & n22087;
  assign n22089 = pi0204 & ~n22087;
  assign n22090 = ~n22088 & ~n22089;
  assign n22091 = ~n22084 & n22090;
  assign n22092 = ~n22078 & n22091;
  assign n22093 = n22072 & n22092;
  assign n22094 = ~n22072 & ~n22078;
  assign n22095 = n22090 & n22094;
  assign n22096 = n22084 & n22095;
  assign n22097 = ~n22093 & ~n22096;
  assign n22098 = ~n22066 & ~n22097;
  assign n22099 = ~n22084 & ~n22090;
  assign n22100 = n22078 & n22099;
  assign n22101 = n22072 & n22100;
  assign n22102 = n22066 & n22101;
  assign n22103 = pi3087 & pi9040;
  assign n22104 = pi3075 & ~pi9040;
  assign n22105 = ~n22103 & ~n22104;
  assign n22106 = ~pi0221 & ~n22105;
  assign n22107 = pi0221 & ~n22103;
  assign n22108 = ~n22104 & n22107;
  assign n22109 = ~n22106 & ~n22108;
  assign n22110 = n22084 & n22090;
  assign n22111 = n22078 & n22110;
  assign n22112 = ~n22066 & n22111;
  assign n22113 = ~n22101 & ~n22112;
  assign n22114 = n22072 & n22084;
  assign n22115 = ~n22078 & n22114;
  assign n22116 = n22072 & n22078;
  assign n22117 = ~n22084 & n22116;
  assign n22118 = ~n22115 & ~n22117;
  assign n22119 = n22066 & ~n22118;
  assign n22120 = n22066 & ~n22072;
  assign n22121 = n22091 & n22120;
  assign n22122 = ~n22078 & n22121;
  assign n22123 = ~n22072 & n22078;
  assign n22124 = ~n22090 & n22123;
  assign n22125 = n22084 & n22124;
  assign n22126 = ~n22078 & n22099;
  assign n22127 = ~n22066 & n22126;
  assign n22128 = ~n22125 & ~n22127;
  assign n22129 = ~n22122 & n22128;
  assign n22130 = ~n22119 & n22129;
  assign n22131 = n22113 & n22130;
  assign n22132 = n22109 & ~n22131;
  assign n22133 = n22072 & n22112;
  assign n22134 = ~n22132 & ~n22133;
  assign n22135 = ~n22102 & n22134;
  assign n22136 = ~n22098 & n22135;
  assign n22137 = ~n22066 & ~n22072;
  assign n22138 = n22078 & ~n22084;
  assign n22139 = n22137 & n22138;
  assign n22140 = ~n22066 & n22092;
  assign n22141 = ~n22139 & ~n22140;
  assign n22142 = n22084 & ~n22090;
  assign n22143 = n22078 & n22142;
  assign n22144 = ~n22066 & n22143;
  assign n22145 = ~n22078 & n22142;
  assign n22146 = n22072 & n22145;
  assign n22147 = ~n22144 & ~n22146;
  assign n22148 = n22078 & n22091;
  assign n22149 = ~n22072 & n22148;
  assign n22150 = ~n22093 & ~n22149;
  assign n22151 = ~n22072 & n22110;
  assign n22152 = ~n22078 & ~n22090;
  assign n22153 = ~n22151 & ~n22152;
  assign n22154 = n22066 & ~n22153;
  assign n22155 = n22150 & ~n22154;
  assign n22156 = n22147 & n22155;
  assign n22157 = n22141 & n22156;
  assign n22158 = ~n22109 & ~n22157;
  assign n22159 = n22136 & ~n22158;
  assign n22160 = ~pi0226 & ~n22159;
  assign n22161 = pi0226 & n22136;
  assign n22162 = ~n22158 & n22161;
  assign po0262 = n22160 | n22162;
  assign n22164 = n21829 & n21848;
  assign n22165 = ~n21873 & ~n21888;
  assign n22166 = n22164 & ~n22165;
  assign n22167 = n21829 & ~n21854;
  assign n22168 = n21873 & n22167;
  assign n22169 = ~n22166 & ~n22168;
  assign n22170 = n21866 & ~n22169;
  assign n22171 = ~n21848 & n21854;
  assign n22172 = ~n21841 & n22171;
  assign n22173 = n21835 & n22172;
  assign n22174 = ~n21905 & ~n22171;
  assign n22175 = ~n21829 & ~n22174;
  assign n22176 = ~n21848 & ~n21854;
  assign n22177 = n21841 & n22176;
  assign n22178 = n21835 & n22177;
  assign n22179 = ~n22175 & ~n22178;
  assign n22180 = ~n22173 & n22179;
  assign n22181 = n21866 & ~n22180;
  assign n22182 = ~n22170 & ~n22181;
  assign n22183 = ~n21841 & n21855;
  assign n22184 = ~n21835 & n22183;
  assign n22185 = ~n21848 & n21880;
  assign n22186 = ~n22184 & ~n22185;
  assign n22187 = n21829 & ~n22186;
  assign n22188 = ~n21842 & ~n21905;
  assign n22189 = n21848 & ~n22188;
  assign n22190 = ~n21880 & ~n22189;
  assign n22191 = n21829 & ~n22190;
  assign n22192 = ~n21841 & ~n21848;
  assign n22193 = n21829 & n22192;
  assign n22194 = ~n21854 & n22193;
  assign n22195 = n21841 & n21854;
  assign n22196 = ~n21880 & ~n22195;
  assign n22197 = ~n21848 & ~n22196;
  assign n22198 = ~n21829 & n21848;
  assign n22199 = n21870 & n22198;
  assign n22200 = ~n21854 & n22199;
  assign n22201 = ~n22197 & ~n22200;
  assign n22202 = ~n22194 & n22201;
  assign n22203 = ~n22191 & n22202;
  assign n22204 = ~n22184 & n22203;
  assign n22205 = ~n21866 & ~n22204;
  assign n22206 = ~n21848 & n21905;
  assign n22207 = n21848 & n21896;
  assign n22208 = ~n22206 & ~n22207;
  assign n22209 = ~n21829 & ~n22208;
  assign n22210 = ~n22205 & ~n22209;
  assign n22211 = ~n22187 & n22210;
  assign n22212 = n22182 & n22211;
  assign n22213 = pi0235 & n22212;
  assign n22214 = ~pi0235 & ~n22212;
  assign po0263 = n22213 | n22214;
  assign n22216 = ~n22066 & n22099;
  assign n22217 = n22072 & n22216;
  assign n22218 = ~n22078 & n22110;
  assign n22219 = n22084 & n22094;
  assign n22220 = ~n22218 & ~n22219;
  assign n22221 = ~n22066 & ~n22220;
  assign n22222 = ~n22217 & ~n22221;
  assign n22223 = n22066 & n22072;
  assign n22224 = n22142 & n22223;
  assign n22225 = n22066 & n22092;
  assign n22226 = ~n22224 & ~n22225;
  assign n22227 = n22222 & n22226;
  assign n22228 = n22084 & n22116;
  assign n22229 = ~n22093 & ~n22228;
  assign n22230 = ~n22149 & n22229;
  assign n22231 = n22227 & n22230;
  assign n22232 = ~n22109 & ~n22231;
  assign n22233 = ~n22133 & ~n22139;
  assign n22234 = ~n22101 & ~n22218;
  assign n22235 = ~n22151 & n22234;
  assign n22236 = n22066 & ~n22235;
  assign n22237 = ~n22090 & n22094;
  assign n22238 = ~n22084 & n22237;
  assign n22239 = ~n22125 & ~n22238;
  assign n22240 = ~n22066 & n22072;
  assign n22241 = n22145 & n22240;
  assign n22242 = n22239 & ~n22241;
  assign n22243 = ~n22066 & n22148;
  assign n22244 = n22242 & ~n22243;
  assign n22245 = ~n22236 & n22244;
  assign n22246 = n22109 & ~n22245;
  assign n22247 = ~n22093 & n22239;
  assign n22248 = n22066 & ~n22247;
  assign n22249 = ~n22246 & ~n22248;
  assign n22250 = n22233 & n22249;
  assign n22251 = ~n22232 & n22250;
  assign n22252 = pi0230 & ~n22251;
  assign n22253 = ~pi0230 & n22251;
  assign po0264 = n22252 | n22253;
  assign n22255 = n21841 & n21857;
  assign n22256 = ~n21888 & ~n22255;
  assign n22257 = n21829 & ~n22256;
  assign n22258 = n21848 & n21879;
  assign n22259 = ~n22177 & ~n22258;
  assign n22260 = ~n21829 & ~n22259;
  assign n22261 = ~n21848 & n21874;
  assign n22262 = ~n22194 & ~n22261;
  assign n22263 = ~n22260 & n22262;
  assign n22264 = ~n21856 & n22263;
  assign n22265 = ~n22257 & n22264;
  assign n22266 = ~n22173 & ~n22184;
  assign n22267 = n22265 & n22266;
  assign n22268 = n21866 & ~n22267;
  assign n22269 = n21835 & n21857;
  assign n22270 = n21848 & n21870;
  assign n22271 = ~n22269 & ~n22270;
  assign n22272 = ~n21829 & ~n22271;
  assign n22273 = ~n21829 & n21879;
  assign n22274 = ~n21848 & n22273;
  assign n22275 = ~n22272 & ~n22274;
  assign n22276 = n21842 & n22171;
  assign n22277 = n21897 & ~n22276;
  assign n22278 = ~n21829 & ~n22277;
  assign n22279 = ~n21848 & n21885;
  assign n22280 = ~n22278 & ~n22279;
  assign n22281 = n22275 & n22280;
  assign n22282 = ~n21866 & ~n22281;
  assign n22283 = ~n21874 & ~n21881;
  assign n22284 = ~n22178 & n22283;
  assign n22285 = n21902 & ~n22284;
  assign n22286 = ~n22282 & ~n22285;
  assign n22287 = ~n21856 & ~n22173;
  assign n22288 = n21829 & ~n22287;
  assign n22289 = n22286 & ~n22288;
  assign n22290 = ~n22268 & n22289;
  assign n22291 = ~pi0248 & n22290;
  assign n22292 = pi0248 & ~n22290;
  assign po0270 = n22291 | n22292;
  assign n22294 = ~n21945 & n21989;
  assign n22295 = ~n22029 & ~n22294;
  assign n22296 = n21951 & ~n22295;
  assign n22297 = n21975 & n21986;
  assign n22298 = ~n22296 & ~n22297;
  assign n22299 = ~n21999 & n22298;
  assign n22300 = ~n21932 & n21945;
  assign n22301 = n21926 & n22300;
  assign n22302 = n21938 & n22301;
  assign n22303 = ~n21959 & ~n22302;
  assign n22304 = ~n21989 & n22303;
  assign n22305 = n21951 & ~n22304;
  assign n22306 = n21920 & n22305;
  assign n22307 = ~n21926 & ~n21951;
  assign n22308 = n21938 & n22307;
  assign n22309 = n21932 & n22308;
  assign n22310 = ~n21945 & n22309;
  assign n22311 = ~n21951 & n22038;
  assign n22312 = ~n21970 & ~n21997;
  assign n22313 = ~n21964 & n22312;
  assign n22314 = ~n22311 & n22313;
  assign n22315 = n21920 & ~n22314;
  assign n22316 = n21945 & n22007;
  assign n22317 = ~n22309 & ~n22316;
  assign n22318 = ~n22028 & n22317;
  assign n22319 = n21938 & n21968;
  assign n22320 = n21945 & n21956;
  assign n22321 = ~n21985 & ~n22320;
  assign n22322 = n21951 & ~n22321;
  assign n22323 = ~n22319 & ~n22322;
  assign n22324 = n22318 & n22323;
  assign n22325 = ~n21920 & ~n22324;
  assign n22326 = ~n22315 & ~n22325;
  assign n22327 = ~n22310 & n22326;
  assign n22328 = ~n22306 & n22327;
  assign n22329 = n22299 & n22328;
  assign n22330 = pi0238 & ~n22329;
  assign n22331 = ~pi0238 & n22299;
  assign n22332 = n22328 & n22331;
  assign po0271 = n22330 | n22332;
  assign n22334 = pi3117 & pi9040;
  assign n22335 = pi3104 & ~pi9040;
  assign n22336 = ~n22334 & ~n22335;
  assign n22337 = pi0177 & n22336;
  assign n22338 = ~pi0177 & ~n22336;
  assign n22339 = ~n22337 & ~n22338;
  assign n22340 = pi3119 & pi9040;
  assign n22341 = pi3120 & ~pi9040;
  assign n22342 = ~n22340 & ~n22341;
  assign n22343 = pi0222 & n22342;
  assign n22344 = ~pi0222 & ~n22342;
  assign n22345 = ~n22343 & ~n22344;
  assign n22346 = pi3169 & pi9040;
  assign n22347 = pi3074 & ~pi9040;
  assign n22348 = ~n22346 & ~n22347;
  assign n22349 = ~pi0221 & ~n22348;
  assign n22350 = pi0221 & ~n22346;
  assign n22351 = ~n22347 & n22350;
  assign n22352 = ~n22349 & ~n22351;
  assign n22353 = pi3120 & pi9040;
  assign n22354 = pi3188 & ~pi9040;
  assign n22355 = ~n22353 & ~n22354;
  assign n22356 = ~pi0204 & n22355;
  assign n22357 = pi0204 & ~n22355;
  assign n22358 = ~n22356 & ~n22357;
  assign n22359 = pi3084 & pi9040;
  assign n22360 = pi3089 & ~pi9040;
  assign n22361 = ~n22359 & ~n22360;
  assign n22362 = ~pi0216 & ~n22361;
  assign n22363 = pi0216 & n22361;
  assign n22364 = ~n22362 & ~n22363;
  assign n22365 = ~n22358 & ~n22364;
  assign n22366 = n22352 & n22365;
  assign n22367 = n22345 & n22366;
  assign n22368 = pi3077 & pi9040;
  assign n22369 = pi3116 & ~pi9040;
  assign n22370 = ~n22368 & ~n22369;
  assign n22371 = ~pi0185 & n22370;
  assign n22372 = pi0185 & ~n22370;
  assign n22373 = ~n22371 & ~n22372;
  assign n22374 = n22352 & n22364;
  assign n22375 = ~n22358 & n22374;
  assign n22376 = ~n22352 & n22358;
  assign n22377 = n22358 & ~n22364;
  assign n22378 = ~n22345 & n22377;
  assign n22379 = ~n22352 & ~n22364;
  assign n22380 = n22345 & n22379;
  assign n22381 = ~n22378 & ~n22380;
  assign n22382 = ~n22376 & n22381;
  assign n22383 = ~n22375 & n22382;
  assign n22384 = ~n22373 & ~n22383;
  assign n22385 = ~n22345 & ~n22358;
  assign n22386 = n22364 & n22385;
  assign n22387 = ~n22352 & n22385;
  assign n22388 = n22358 & n22374;
  assign n22389 = ~n22387 & ~n22388;
  assign n22390 = n22373 & ~n22389;
  assign n22391 = ~n22386 & ~n22390;
  assign n22392 = ~n22384 & n22391;
  assign n22393 = ~n22367 & n22392;
  assign n22394 = n22339 & ~n22393;
  assign n22395 = ~n22352 & n22364;
  assign n22396 = n22358 & n22395;
  assign n22397 = ~n22345 & n22396;
  assign n22398 = n22358 & n22379;
  assign n22399 = n22345 & n22398;
  assign n22400 = ~n22367 & ~n22399;
  assign n22401 = ~n22397 & n22400;
  assign n22402 = ~n22373 & ~n22401;
  assign n22403 = ~n22394 & ~n22402;
  assign n22404 = ~n22345 & n22375;
  assign n22405 = n22345 & n22358;
  assign n22406 = n22373 & n22405;
  assign n22407 = n22352 & n22406;
  assign n22408 = ~n22358 & n22395;
  assign n22409 = n22345 & n22408;
  assign n22410 = ~n22364 & ~n22373;
  assign n22411 = ~n22358 & n22410;
  assign n22412 = ~n22345 & n22411;
  assign n22413 = ~n22409 & ~n22412;
  assign n22414 = ~n22352 & ~n22358;
  assign n22415 = n22345 & n22414;
  assign n22416 = n22352 & ~n22364;
  assign n22417 = n22358 & n22416;
  assign n22418 = ~n22415 & ~n22417;
  assign n22419 = n22373 & ~n22418;
  assign n22420 = n22373 & n22376;
  assign n22421 = ~n22345 & n22420;
  assign n22422 = ~n22419 & ~n22421;
  assign n22423 = n22413 & n22422;
  assign n22424 = ~n22339 & ~n22423;
  assign n22425 = ~n22407 & ~n22424;
  assign n22426 = ~n22404 & n22425;
  assign n22427 = n22403 & n22426;
  assign n22428 = ~pi0242 & ~n22427;
  assign n22429 = ~n22394 & ~n22404;
  assign n22430 = ~n22402 & n22429;
  assign n22431 = n22425 & n22430;
  assign n22432 = pi0242 & n22431;
  assign po0272 = n22428 | n22432;
  assign n22434 = ~n22072 & n22100;
  assign n22435 = ~n22072 & n22142;
  assign n22436 = n22072 & n22126;
  assign n22437 = ~n22435 & ~n22436;
  assign n22438 = n22066 & ~n22437;
  assign n22439 = ~n22434 & ~n22438;
  assign n22440 = ~n22072 & n22216;
  assign n22441 = ~n22140 & ~n22440;
  assign n22442 = n22439 & n22441;
  assign n22443 = ~n22072 & n22111;
  assign n22444 = n22072 & n22148;
  assign n22445 = ~n22443 & ~n22444;
  assign n22446 = n22442 & n22445;
  assign n22447 = n22109 & ~n22446;
  assign n22448 = n22218 & n22223;
  assign n22449 = n22078 & n22137;
  assign n22450 = ~n22099 & n22449;
  assign n22451 = ~n22112 & ~n22450;
  assign n22452 = ~n22101 & ~n22115;
  assign n22453 = n22451 & n22452;
  assign n22454 = ~n22109 & ~n22453;
  assign n22455 = ~n22084 & n22094;
  assign n22456 = ~n22078 & n22090;
  assign n22457 = ~n22455 & ~n22456;
  assign n22458 = n22066 & ~n22109;
  assign n22459 = ~n22457 & n22458;
  assign n22460 = ~n22454 & ~n22459;
  assign n22461 = n22072 & n22143;
  assign n22462 = ~n22444 & ~n22461;
  assign n22463 = n22066 & ~n22462;
  assign n22464 = ~n22066 & n22101;
  assign n22465 = ~n22463 & ~n22464;
  assign n22466 = n22460 & n22465;
  assign n22467 = ~n22448 & n22466;
  assign n22468 = ~n22447 & n22467;
  assign n22469 = ~n22241 & n22468;
  assign n22470 = ~pi0239 & ~n22469;
  assign n22471 = pi0239 & ~n22241;
  assign n22472 = n22467 & n22471;
  assign n22473 = ~n22447 & n22472;
  assign po0273 = n22470 | n22473;
  assign n22475 = ~n21561 & n21604;
  assign n22476 = ~n21805 & ~n22475;
  assign n22477 = ~n21555 & n22476;
  assign n22478 = n21561 & n21574;
  assign n22479 = ~n21592 & ~n21598;
  assign n22480 = n21567 & ~n22479;
  assign n22481 = n21573 & n21620;
  assign n22482 = n21561 & n21598;
  assign n22483 = ~n22481 & ~n22482;
  assign n22484 = n21555 & n22483;
  assign n22485 = ~n22480 & n22484;
  assign n22486 = ~n22478 & n22485;
  assign n22487 = ~n22477 & ~n22486;
  assign n22488 = n21561 & n22480;
  assign n22489 = ~n21803 & ~n22488;
  assign n22490 = ~n22487 & n22489;
  assign n22491 = n21585 & ~n22490;
  assign n22492 = ~n21555 & ~n22479;
  assign n22493 = ~n21561 & n22492;
  assign n22494 = n21561 & n21640;
  assign n22495 = ~n21611 & ~n22494;
  assign n22496 = ~n21555 & ~n22495;
  assign n22497 = ~n21567 & n22492;
  assign n22498 = ~n22496 & ~n22497;
  assign n22499 = ~n22493 & n22498;
  assign n22500 = ~n21585 & ~n22499;
  assign n22501 = ~n22491 & ~n22500;
  assign n22502 = n21555 & ~n22476;
  assign n22503 = ~n21602 & ~n22502;
  assign n22504 = ~n21585 & ~n22503;
  assign n22505 = ~n21555 & n21602;
  assign n22506 = n21555 & ~n22489;
  assign n22507 = ~n22505 & ~n22506;
  assign n22508 = ~n22504 & n22507;
  assign n22509 = n22501 & n22508;
  assign n22510 = pi0240 & ~n22509;
  assign n22511 = ~pi0240 & n22508;
  assign n22512 = ~n22500 & n22511;
  assign n22513 = ~n22491 & n22512;
  assign po0274 = n22510 | n22513;
  assign n22515 = n21700 & ~n21706;
  assign n22516 = ~n21694 & n22515;
  assign n22517 = n21720 & n22516;
  assign n22518 = n21700 & n21720;
  assign n22519 = ~n21712 & n22518;
  assign n22520 = ~n21706 & n22519;
  assign n22521 = ~n21700 & ~n21712;
  assign n22522 = ~n21720 & n22521;
  assign n22523 = ~n21727 & ~n22522;
  assign n22524 = ~n22520 & n22523;
  assign n22525 = ~n22517 & n22524;
  assign n22526 = n21694 & n21723;
  assign n22527 = n22525 & ~n22526;
  assign n22528 = n21758 & ~n22527;
  assign n22529 = ~n21724 & ~n21727;
  assign n22530 = ~n21720 & n21775;
  assign n22531 = n21720 & n21760;
  assign n22532 = ~n22530 & ~n22531;
  assign n22533 = n22529 & n22532;
  assign n22534 = ~n21694 & ~n22533;
  assign n22535 = ~n22528 & ~n22534;
  assign n22536 = ~n21706 & n21765;
  assign n22537 = ~n21776 & ~n22536;
  assign n22538 = n21694 & ~n22537;
  assign n22539 = ~n21700 & ~n21720;
  assign n22540 = n21706 & n22539;
  assign n22541 = ~n22521 & ~n22540;
  assign n22542 = ~n21729 & n22541;
  assign n22543 = n21694 & ~n22542;
  assign n22544 = ~n21720 & n21735;
  assign n22545 = ~n22543 & ~n22544;
  assign n22546 = ~n21758 & ~n22545;
  assign n22547 = ~n21758 & n21760;
  assign n22548 = ~n21694 & n22547;
  assign n22549 = ~n22546 & ~n22548;
  assign n22550 = ~n22538 & n22549;
  assign n22551 = n22535 & n22550;
  assign n22552 = ~pi0247 & ~n22551;
  assign n22553 = pi0247 & n22535;
  assign n22554 = n22550 & n22553;
  assign po0275 = n22552 | n22554;
  assign n22556 = ~n22443 & ~n22455;
  assign n22557 = n22109 & ~n22556;
  assign n22558 = n22066 & n22100;
  assign n22559 = ~n22090 & n22116;
  assign n22560 = ~n22117 & ~n22559;
  assign n22561 = n22066 & ~n22560;
  assign n22562 = ~n22558 & ~n22561;
  assign n22563 = n22109 & ~n22562;
  assign n22564 = ~n22557 & ~n22563;
  assign n22565 = n22111 & n22120;
  assign n22566 = ~n22122 & ~n22565;
  assign n22567 = ~n22115 & ~n22152;
  assign n22568 = ~n22066 & ~n22567;
  assign n22569 = n22109 & n22568;
  assign n22570 = n22566 & ~n22569;
  assign n22571 = n22090 & n22116;
  assign n22572 = n22084 & n22571;
  assign n22573 = n22072 & n22091;
  assign n22574 = ~n22096 & ~n22573;
  assign n22575 = ~n22066 & ~n22574;
  assign n22576 = ~n22101 & ~n22125;
  assign n22577 = n22072 & n22110;
  assign n22578 = ~n22145 & ~n22577;
  assign n22579 = n22066 & ~n22578;
  assign n22580 = n22576 & ~n22579;
  assign n22581 = ~n22575 & n22580;
  assign n22582 = ~n22572 & n22581;
  assign n22583 = ~n22109 & ~n22582;
  assign n22584 = ~n22149 & n22239;
  assign n22585 = ~n22066 & ~n22584;
  assign n22586 = ~n22583 & ~n22585;
  assign n22587 = n22570 & n22586;
  assign n22588 = n22564 & n22587;
  assign n22589 = ~pi0237 & ~n22588;
  assign n22590 = pi0237 & n22570;
  assign n22591 = n22564 & n22590;
  assign n22592 = n22586 & n22591;
  assign po0276 = n22589 | n22592;
  assign n22594 = ~n21720 & n21749;
  assign n22595 = ~n21746 & ~n22531;
  assign n22596 = n21694 & ~n22595;
  assign n22597 = ~n22594 & ~n22596;
  assign n22598 = ~n21712 & n21782;
  assign n22599 = ~n21706 & n22598;
  assign n22600 = n21728 & n21761;
  assign n22601 = ~n22599 & ~n22600;
  assign n22602 = ~n21694 & n21770;
  assign n22603 = n22601 & ~n22602;
  assign n22604 = ~n21724 & ~n21736;
  assign n22605 = n21712 & n21726;
  assign n22606 = n22604 & ~n22605;
  assign n22607 = n22603 & n22606;
  assign n22608 = n22597 & n22607;
  assign n22609 = ~n21758 & ~n22608;
  assign n22610 = ~n21723 & ~n21746;
  assign n22611 = n21720 & ~n22610;
  assign n22612 = ~n21706 & n21764;
  assign n22613 = ~n21775 & ~n22612;
  assign n22614 = n21720 & n22521;
  assign n22615 = n22613 & ~n22614;
  assign n22616 = n21694 & ~n22615;
  assign n22617 = ~n21720 & n21734;
  assign n22618 = ~n22520 & ~n22617;
  assign n22619 = ~n21694 & ~n22618;
  assign n22620 = ~n22536 & ~n22619;
  assign n22621 = ~n22616 & n22620;
  assign n22622 = ~n22611 & n22621;
  assign n22623 = n21758 & ~n22622;
  assign n22624 = n21694 & n21765;
  assign n22625 = ~n22623 & ~n22624;
  assign n22626 = n21741 & n21782;
  assign n22627 = ~n21712 & n22626;
  assign n22628 = n22625 & ~n22627;
  assign n22629 = ~n22609 & n22628;
  assign n22630 = ~pi0249 & ~n22629;
  assign n22631 = pi0249 & n22625;
  assign n22632 = ~n22609 & n22631;
  assign n22633 = ~n22627 & n22632;
  assign po0277 = n22630 | n22633;
  assign n22635 = ~n22358 & n22379;
  assign n22636 = n22345 & n22635;
  assign n22637 = n22345 & n22396;
  assign n22638 = ~n22636 & ~n22637;
  assign n22639 = ~n22345 & n22398;
  assign n22640 = ~n22388 & ~n22639;
  assign n22641 = ~n22373 & ~n22640;
  assign n22642 = n22638 & ~n22641;
  assign n22643 = ~n22345 & n22373;
  assign n22644 = n22352 & n22643;
  assign n22645 = n22642 & ~n22644;
  assign n22646 = n22339 & ~n22645;
  assign n22647 = n22345 & n22352;
  assign n22648 = n22358 & n22647;
  assign n22649 = ~n22364 & n22648;
  assign n22650 = n22373 & n22649;
  assign n22651 = ~n22345 & ~n22373;
  assign n22652 = n22417 & n22651;
  assign n22653 = ~n22387 & ~n22652;
  assign n22654 = ~n22388 & ~n22408;
  assign n22655 = ~n22345 & n22395;
  assign n22656 = n22654 & ~n22655;
  assign n22657 = n22373 & ~n22656;
  assign n22658 = ~n22373 & n22375;
  assign n22659 = n22400 & ~n22658;
  assign n22660 = ~n22657 & n22659;
  assign n22661 = n22653 & n22660;
  assign n22662 = ~n22339 & ~n22661;
  assign n22663 = ~n22650 & ~n22662;
  assign n22664 = ~n22646 & n22663;
  assign n22665 = n22408 & n22651;
  assign n22666 = n22345 & n22411;
  assign n22667 = ~n22665 & ~n22666;
  assign n22668 = ~n22373 & n22637;
  assign n22669 = n22667 & ~n22668;
  assign n22670 = n22664 & n22669;
  assign n22671 = ~pi0243 & ~n22670;
  assign n22672 = ~n22646 & n22669;
  assign n22673 = n22663 & n22672;
  assign n22674 = pi0243 & n22673;
  assign po0278 = n22671 | n22674;
  assign n22676 = n21700 & n21706;
  assign n22677 = n21694 & n22676;
  assign n22678 = n21720 & n22677;
  assign n22679 = ~n21694 & n21713;
  assign n22680 = n21720 & n22679;
  assign n22681 = ~n22602 & ~n22680;
  assign n22682 = n21720 & n21734;
  assign n22683 = ~n22676 & ~n22682;
  assign n22684 = ~n21706 & n22539;
  assign n22685 = n22683 & ~n22684;
  assign n22686 = n21694 & ~n22685;
  assign n22687 = ~n21730 & ~n22686;
  assign n22688 = n22681 & n22687;
  assign n22689 = ~n21758 & ~n22688;
  assign n22690 = ~n21746 & ~n21765;
  assign n22691 = ~n21775 & n22690;
  assign n22692 = ~n21694 & ~n22691;
  assign n22693 = ~n21720 & n21770;
  assign n22694 = ~n21749 & ~n22693;
  assign n22695 = n21694 & ~n22694;
  assign n22696 = ~n22612 & ~n22695;
  assign n22697 = ~n22692 & n22696;
  assign n22698 = ~n21736 & ~n21776;
  assign n22699 = n22697 & n22698;
  assign n22700 = n21758 & ~n22699;
  assign n22701 = ~n21721 & ~n21727;
  assign n22702 = ~n21694 & ~n22701;
  assign n22703 = ~n21784 & ~n22702;
  assign n22704 = ~n22700 & n22703;
  assign n22705 = ~n22689 & n22704;
  assign n22706 = ~n22678 & n22705;
  assign n22707 = pi0252 & n22706;
  assign n22708 = ~pi0252 & ~n22706;
  assign po0279 = n22707 | n22708;
  assign n22710 = ~n21555 & n21628;
  assign n22711 = n21620 & ~n22479;
  assign n22712 = ~n21641 & ~n22711;
  assign n22713 = ~n21803 & n22712;
  assign n22714 = n21555 & ~n22713;
  assign n22715 = n21561 & n21599;
  assign n22716 = ~n22714 & ~n22715;
  assign n22717 = ~n21567 & n21640;
  assign n22718 = ~n21561 & n21810;
  assign n22719 = ~n22717 & ~n22718;
  assign n22720 = ~n22482 & n22719;
  assign n22721 = ~n21555 & ~n22720;
  assign n22722 = n22716 & ~n22721;
  assign n22723 = n21585 & ~n22722;
  assign n22724 = ~n22710 & ~n22723;
  assign n22725 = ~n21561 & n21598;
  assign n22726 = ~n21802 & ~n22725;
  assign n22727 = ~n21555 & ~n22726;
  assign n22728 = ~n21642 & ~n22727;
  assign n22729 = ~n21611 & ~n21628;
  assign n22730 = n21561 & n21637;
  assign n22731 = ~n21810 & ~n22730;
  assign n22732 = ~n22717 & n22731;
  assign n22733 = n21555 & ~n22732;
  assign n22734 = ~n21561 & n21599;
  assign n22735 = ~n22733 & ~n22734;
  assign n22736 = n22729 & n22735;
  assign n22737 = n22728 & n22736;
  assign n22738 = ~n21585 & ~n22737;
  assign n22739 = ~n21631 & ~n22478;
  assign n22740 = n21555 & ~n22739;
  assign n22741 = ~n22738 & ~n22740;
  assign n22742 = n22724 & n22741;
  assign n22743 = pi0244 & n22742;
  assign n22744 = ~pi0244 & ~n22742;
  assign po0280 = n22743 | n22744;
  assign n22746 = pi3090 & pi9040;
  assign n22747 = pi3094 & ~pi9040;
  assign n22748 = ~n22746 & ~n22747;
  assign n22749 = pi0214 & n22748;
  assign n22750 = ~pi0214 & ~n22748;
  assign n22751 = ~n22749 & ~n22750;
  assign n22752 = pi3118 & pi9040;
  assign n22753 = pi3086 & ~pi9040;
  assign n22754 = ~n22752 & ~n22753;
  assign n22755 = pi0217 & n22754;
  assign n22756 = ~pi0217 & ~n22754;
  assign n22757 = ~n22755 & ~n22756;
  assign n22758 = pi3082 & pi9040;
  assign n22759 = pi3122 & ~pi9040;
  assign n22760 = ~n22758 & ~n22759;
  assign n22761 = ~pi0205 & n22760;
  assign n22762 = pi0205 & ~n22760;
  assign n22763 = ~n22761 & ~n22762;
  assign n22764 = ~n22757 & ~n22763;
  assign n22765 = ~n22751 & n22764;
  assign n22766 = n22757 & ~n22763;
  assign n22767 = n22751 & n22766;
  assign n22768 = ~n22765 & ~n22767;
  assign n22769 = pi3094 & pi9040;
  assign n22770 = pi3093 & ~pi9040;
  assign n22771 = ~n22769 & ~n22770;
  assign n22772 = pi0181 & n22771;
  assign n22773 = ~pi0181 & ~n22771;
  assign n22774 = ~n22772 & ~n22773;
  assign n22775 = n22751 & ~n22774;
  assign n22776 = n22757 & n22775;
  assign n22777 = n22768 & ~n22776;
  assign n22778 = pi3168 & pi9040;
  assign n22779 = pi3092 & ~pi9040;
  assign n22780 = ~n22778 & ~n22779;
  assign n22781 = ~pi0176 & n22780;
  assign n22782 = pi0176 & ~n22780;
  assign n22783 = ~n22781 & ~n22782;
  assign n22784 = pi3225 & pi9040;
  assign n22785 = pi3090 & ~pi9040;
  assign n22786 = ~n22784 & ~n22785;
  assign n22787 = ~pi0203 & n22786;
  assign n22788 = pi0203 & ~n22786;
  assign n22789 = ~n22787 & ~n22788;
  assign n22790 = n22783 & ~n22789;
  assign n22791 = ~n22777 & n22790;
  assign n22792 = ~n22757 & n22763;
  assign n22793 = n22751 & n22792;
  assign n22794 = ~n22789 & n22793;
  assign n22795 = n22774 & n22794;
  assign n22796 = n22751 & n22764;
  assign n22797 = ~n22783 & n22796;
  assign n22798 = ~n22751 & n22757;
  assign n22799 = n22757 & n22763;
  assign n22800 = n22774 & n22799;
  assign n22801 = ~n22798 & ~n22800;
  assign n22802 = ~n22783 & ~n22801;
  assign n22803 = ~n22797 & ~n22802;
  assign n22804 = ~n22789 & ~n22803;
  assign n22805 = ~n22795 & ~n22804;
  assign n22806 = ~n22751 & n22774;
  assign n22807 = n22757 & n22806;
  assign n22808 = ~n22751 & ~n22774;
  assign n22809 = ~n22757 & n22808;
  assign n22810 = n22763 & n22809;
  assign n22811 = ~n22807 & ~n22810;
  assign n22812 = ~n22783 & ~n22811;
  assign n22813 = n22805 & ~n22812;
  assign n22814 = n22774 & n22783;
  assign n22815 = n22799 & n22814;
  assign n22816 = n22751 & n22815;
  assign n22817 = ~n22766 & ~n22792;
  assign n22818 = n22775 & ~n22817;
  assign n22819 = n22765 & ~n22774;
  assign n22820 = ~n22818 & ~n22819;
  assign n22821 = ~n22751 & n22799;
  assign n22822 = n22783 & n22821;
  assign n22823 = ~n22774 & n22822;
  assign n22824 = n22806 & ~n22817;
  assign n22825 = n22774 & n22796;
  assign n22826 = ~n22824 & ~n22825;
  assign n22827 = ~n22823 & n22826;
  assign n22828 = n22820 & n22827;
  assign n22829 = ~n22816 & n22828;
  assign n22830 = ~n22774 & ~n22783;
  assign n22831 = n22751 & n22830;
  assign n22832 = n22763 & n22831;
  assign n22833 = n22829 & ~n22832;
  assign n22834 = n22789 & ~n22833;
  assign n22835 = n22813 & ~n22834;
  assign n22836 = ~n22791 & n22835;
  assign n22837 = ~pi0259 & ~n22836;
  assign n22838 = pi0259 & n22813;
  assign n22839 = ~n22791 & n22838;
  assign n22840 = ~n22834 & n22839;
  assign po0281 = n22837 | n22840;
  assign n22842 = n21945 & ~n22050;
  assign n22843 = n21926 & n22842;
  assign n22844 = n21938 & n22027;
  assign n22845 = ~n22009 & ~n22844;
  assign n22846 = ~n21959 & n22845;
  assign n22847 = ~n21951 & ~n22846;
  assign n22848 = ~n21973 & ~n22038;
  assign n22849 = n21951 & ~n22848;
  assign n22850 = ~n22847 & ~n22849;
  assign n22851 = ~n22843 & n22850;
  assign n22852 = ~n21945 & n21986;
  assign n22853 = n22851 & ~n22852;
  assign n22854 = ~n21920 & ~n22853;
  assign n22855 = n21955 & ~n22848;
  assign n22856 = ~n21974 & ~n21989;
  assign n22857 = ~n21959 & ~n21986;
  assign n22858 = n22856 & n22857;
  assign n22859 = n21945 & ~n22858;
  assign n22860 = ~n22855 & ~n22859;
  assign n22861 = ~n22029 & n22860;
  assign n22862 = n21920 & ~n22861;
  assign n22863 = ~n22854 & ~n22862;
  assign n22864 = n21945 & n22038;
  assign n22865 = ~n22852 & ~n22864;
  assign n22866 = n21951 & ~n22865;
  assign n22867 = n22863 & ~n22866;
  assign n22868 = pi0232 & ~n22867;
  assign n22869 = ~pi0232 & ~n22866;
  assign n22870 = ~n22862 & n22869;
  assign n22871 = ~n22854 & n22870;
  assign po0282 = n22868 | n22871;
  assign n22873 = n22774 & n22792;
  assign n22874 = ~n22751 & n22873;
  assign n22875 = ~n22825 & ~n22874;
  assign n22876 = ~n22783 & ~n22875;
  assign n22877 = ~n22751 & n22766;
  assign n22878 = n22751 & n22799;
  assign n22879 = ~n22877 & ~n22878;
  assign n22880 = ~n22783 & ~n22879;
  assign n22881 = ~n22774 & n22792;
  assign n22882 = ~n22767 & ~n22881;
  assign n22883 = ~n22821 & n22882;
  assign n22884 = n22783 & ~n22883;
  assign n22885 = ~n22880 & ~n22884;
  assign n22886 = ~n22797 & ~n22810;
  assign n22887 = n22885 & n22886;
  assign n22888 = n22789 & ~n22887;
  assign n22889 = n22774 & n22878;
  assign n22890 = n22764 & ~n22774;
  assign n22891 = ~n22873 & ~n22890;
  assign n22892 = n22783 & ~n22891;
  assign n22893 = ~n22889 & ~n22892;
  assign n22894 = n22751 & ~n22783;
  assign n22895 = ~n22757 & n22894;
  assign n22896 = n22763 & n22895;
  assign n22897 = n22768 & ~n22896;
  assign n22898 = ~n22821 & n22897;
  assign n22899 = ~n22774 & ~n22898;
  assign n22900 = n22893 & ~n22899;
  assign n22901 = ~n22789 & ~n22900;
  assign n22902 = ~n22888 & ~n22901;
  assign n22903 = ~n22751 & ~n22763;
  assign n22904 = n22814 & n22903;
  assign n22905 = n22902 & ~n22904;
  assign n22906 = ~n22876 & n22905;
  assign n22907 = ~pi0253 & ~n22906;
  assign n22908 = pi0253 & ~n22876;
  assign n22909 = n22902 & n22908;
  assign n22910 = ~n22904 & n22909;
  assign po0283 = n22907 | n22910;
  assign n22912 = n21829 & n21885;
  assign n22913 = ~n21848 & n21870;
  assign n22914 = ~n21869 & ~n22913;
  assign n22915 = n21829 & ~n22914;
  assign n22916 = ~n21829 & ~n22196;
  assign n22917 = ~n22915 & ~n22916;
  assign n22918 = ~n22207 & n22917;
  assign n22919 = n21866 & ~n22918;
  assign n22920 = ~n22912 & ~n22919;
  assign n22921 = n21854 & n22164;
  assign n22922 = ~n22176 & ~n22921;
  assign n22923 = ~n21835 & ~n22922;
  assign n22924 = ~n21856 & ~n22923;
  assign n22925 = ~n22177 & n22924;
  assign n22926 = ~n21829 & n21871;
  assign n22927 = n21848 & n21888;
  assign n22928 = ~n22926 & ~n22927;
  assign n22929 = n22925 & n22928;
  assign n22930 = ~n21866 & ~n22929;
  assign n22931 = ~n22261 & ~n22270;
  assign n22932 = ~n21829 & ~n22931;
  assign n22933 = ~n22930 & ~n22932;
  assign n22934 = n22920 & n22933;
  assign n22935 = ~pi0267 & ~n22934;
  assign n22936 = pi0267 & n22933;
  assign n22937 = ~n22919 & n22936;
  assign n22938 = ~n22912 & n22937;
  assign po0284 = n22935 | n22938;
  assign n22940 = ~n22783 & n22878;
  assign n22941 = ~n22774 & n22940;
  assign n22942 = n22764 & n22830;
  assign n22943 = ~n22751 & n22942;
  assign n22944 = ~n22941 & ~n22943;
  assign n22945 = ~n22819 & ~n22823;
  assign n22946 = ~n22763 & n22774;
  assign n22947 = n22751 & n22946;
  assign n22948 = ~n22800 & ~n22947;
  assign n22949 = ~n22783 & ~n22948;
  assign n22950 = n22783 & ~n22808;
  assign n22951 = ~n22817 & n22950;
  assign n22952 = ~n22751 & ~n22799;
  assign n22953 = ~n22783 & n22952;
  assign n22954 = ~n22774 & n22953;
  assign n22955 = ~n22951 & ~n22954;
  assign n22956 = ~n22949 & n22955;
  assign n22957 = n22945 & n22956;
  assign n22958 = ~n22789 & ~n22957;
  assign n22959 = n22944 & ~n22958;
  assign n22960 = n22767 & n22783;
  assign n22961 = n22774 & n22960;
  assign n22962 = n22783 & n22789;
  assign n22963 = n22808 & ~n22817;
  assign n22964 = ~n22800 & ~n22963;
  assign n22965 = ~n22796 & n22964;
  assign n22966 = n22962 & ~n22965;
  assign n22967 = n22765 & n22774;
  assign n22968 = ~n22751 & n22946;
  assign n22969 = ~n22873 & ~n22968;
  assign n22970 = ~n22774 & n22799;
  assign n22971 = ~n22793 & ~n22970;
  assign n22972 = n22969 & n22971;
  assign n22973 = ~n22783 & ~n22972;
  assign n22974 = ~n22967 & ~n22973;
  assign n22975 = n22789 & ~n22974;
  assign n22976 = ~n22966 & ~n22975;
  assign n22977 = ~n22961 & n22976;
  assign n22978 = n22959 & n22977;
  assign n22979 = pi0260 & ~n22978;
  assign n22980 = ~pi0260 & n22959;
  assign n22981 = n22977 & n22980;
  assign po0285 = n22979 | n22981;
  assign n22983 = ~n22793 & ~n22946;
  assign n22984 = n22790 & ~n22983;
  assign n22985 = n22751 & n22774;
  assign n22986 = ~n22766 & n22985;
  assign n22987 = ~n22789 & n22986;
  assign n22988 = ~n22783 & n22806;
  assign n22989 = n22766 & n22988;
  assign n22990 = n22751 & n22814;
  assign n22991 = ~n22757 & n22990;
  assign n22992 = ~n22989 & ~n22991;
  assign n22993 = ~n22987 & n22992;
  assign n22994 = ~n22873 & ~n22970;
  assign n22995 = ~n22783 & ~n22994;
  assign n22996 = ~n22943 & ~n22995;
  assign n22997 = ~n22789 & ~n22996;
  assign n22998 = ~n22766 & ~n22903;
  assign n22999 = ~n22774 & ~n22998;
  assign n23000 = ~n22878 & ~n22999;
  assign n23001 = n22783 & ~n23000;
  assign n23002 = ~n22963 & ~n23001;
  assign n23003 = n22774 & n22821;
  assign n23004 = ~n22757 & n22775;
  assign n23005 = n22774 & ~n22998;
  assign n23006 = ~n23004 & ~n23005;
  assign n23007 = ~n22783 & ~n23006;
  assign n23008 = ~n23003 & ~n23007;
  assign n23009 = n23002 & n23008;
  assign n23010 = n22789 & ~n23009;
  assign n23011 = ~n22997 & ~n23010;
  assign n23012 = n22993 & n23011;
  assign n23013 = ~n22984 & n23012;
  assign n23014 = pi0268 & ~n23013;
  assign n23015 = ~pi0268 & n22993;
  assign n23016 = ~n22984 & n23015;
  assign n23017 = n23011 & n23016;
  assign po0286 = n23014 | n23017;
  assign n23019 = ~n22364 & n22385;
  assign n23020 = ~n22352 & n23019;
  assign n23021 = ~n22396 & ~n22404;
  assign n23022 = n22345 & n22365;
  assign n23023 = ~n22345 & n22417;
  assign n23024 = ~n23022 & ~n23023;
  assign n23025 = n23021 & n23024;
  assign n23026 = n22373 & ~n23025;
  assign n23027 = n22345 & n22374;
  assign n23028 = ~n22387 & ~n23027;
  assign n23029 = ~n22398 & n23028;
  assign n23030 = ~n22373 & ~n23029;
  assign n23031 = n22364 & n22405;
  assign n23032 = n22352 & n23031;
  assign n23033 = ~n23030 & ~n23032;
  assign n23034 = ~n23026 & n23033;
  assign n23035 = ~n23020 & n23034;
  assign n23036 = ~n22339 & ~n23035;
  assign n23037 = n22345 & n22373;
  assign n23038 = n22375 & n23037;
  assign n23039 = n22373 & n22398;
  assign n23040 = n22373 & n22408;
  assign n23041 = ~n23039 & ~n23040;
  assign n23042 = ~n22345 & ~n23041;
  assign n23043 = ~n23038 & ~n23042;
  assign n23044 = ~n22345 & n22366;
  assign n23045 = ~n22649 & ~n23044;
  assign n23046 = n22345 & n22395;
  assign n23047 = ~n22345 & n22374;
  assign n23048 = ~n23046 & ~n23047;
  assign n23049 = ~n22366 & n23048;
  assign n23050 = ~n22396 & n23049;
  assign n23051 = ~n22373 & ~n23050;
  assign n23052 = ~n22345 & n22388;
  assign n23053 = ~n23051 & ~n23052;
  assign n23054 = n23045 & n23053;
  assign n23055 = n23043 & n23054;
  assign n23056 = n22339 & ~n23055;
  assign n23057 = n22373 & ~n22638;
  assign n23058 = ~n23056 & ~n23057;
  assign n23059 = ~n22399 & ~n23044;
  assign n23060 = ~n22373 & ~n23059;
  assign n23061 = n23058 & ~n23060;
  assign n23062 = ~n23036 & n23061;
  assign n23063 = pi0246 & ~n23062;
  assign n23064 = ~pi0246 & n23062;
  assign po0287 = n23063 | n23064;
  assign n23066 = ~n22639 & ~n23044;
  assign n23067 = ~n23032 & n23066;
  assign n23068 = n22373 & ~n23067;
  assign n23069 = ~n22652 & ~n22668;
  assign n23070 = ~n22649 & ~n23040;
  assign n23071 = ~n22635 & ~n23047;
  assign n23072 = ~n22373 & ~n23071;
  assign n23073 = ~n22404 & ~n23072;
  assign n23074 = n23070 & n23073;
  assign n23075 = n22339 & ~n23074;
  assign n23076 = n22358 & n22364;
  assign n23077 = ~n22376 & ~n23076;
  assign n23078 = n22345 & ~n23077;
  assign n23079 = ~n22366 & ~n22655;
  assign n23080 = ~n22373 & ~n23079;
  assign n23081 = n22345 & n22364;
  assign n23082 = ~n22388 & ~n23081;
  assign n23083 = ~n22379 & n23082;
  assign n23084 = n22373 & ~n23083;
  assign n23085 = ~n23080 & ~n23084;
  assign n23086 = ~n23078 & n23085;
  assign n23087 = ~n22339 & ~n23086;
  assign n23088 = ~n23075 & ~n23087;
  assign n23089 = n23069 & n23088;
  assign n23090 = ~n23068 & n23089;
  assign n23091 = ~pi0258 & ~n23090;
  assign n23092 = pi0258 & n23069;
  assign n23093 = ~n23068 & n23092;
  assign n23094 = n23088 & n23093;
  assign po0289 = n23091 | n23094;
  assign n23096 = pi3183 & ~pi9040;
  assign n23097 = pi3136 & pi9040;
  assign n23098 = ~n23096 & ~n23097;
  assign n23099 = ~pi0285 & ~n23098;
  assign n23100 = pi0285 & n23098;
  assign n23101 = ~n23099 & ~n23100;
  assign n23102 = pi3182 & pi9040;
  assign n23103 = pi3152 & ~pi9040;
  assign n23104 = ~n23102 & ~n23103;
  assign n23105 = ~pi0264 & n23104;
  assign n23106 = pi0264 & ~n23104;
  assign n23107 = ~n23105 & ~n23106;
  assign n23108 = pi3196 & pi9040;
  assign n23109 = pi3171 & ~pi9040;
  assign n23110 = ~n23108 & ~n23109;
  assign n23111 = pi0245 & n23110;
  assign n23112 = ~pi0245 & ~n23110;
  assign n23113 = ~n23111 & ~n23112;
  assign n23114 = pi3171 & pi9040;
  assign n23115 = pi3181 & ~pi9040;
  assign n23116 = ~n23114 & ~n23115;
  assign n23117 = ~pi0279 & n23116;
  assign n23118 = pi0279 & ~n23116;
  assign n23119 = ~n23117 & ~n23118;
  assign n23120 = pi3151 & pi9040;
  assign n23121 = pi3235 & ~pi9040;
  assign n23122 = ~n23120 & ~n23121;
  assign n23123 = ~pi0256 & ~n23122;
  assign n23124 = pi0256 & ~n23120;
  assign n23125 = ~n23121 & n23124;
  assign n23126 = ~n23123 & ~n23125;
  assign n23127 = ~n23119 & ~n23126;
  assign n23128 = n23113 & n23127;
  assign n23129 = pi3158 & pi9040;
  assign n23130 = pi3128 & ~pi9040;
  assign n23131 = ~n23129 & ~n23130;
  assign n23132 = ~pi0272 & n23131;
  assign n23133 = pi0272 & ~n23131;
  assign n23134 = ~n23132 & ~n23133;
  assign n23135 = n23126 & ~n23134;
  assign n23136 = ~n23119 & n23135;
  assign n23137 = ~n23128 & ~n23136;
  assign n23138 = n23126 & n23134;
  assign n23139 = n23119 & n23138;
  assign n23140 = ~n23113 & n23139;
  assign n23141 = n23137 & ~n23140;
  assign n23142 = ~n23107 & ~n23141;
  assign n23143 = n23119 & n23126;
  assign n23144 = ~n23113 & ~n23134;
  assign n23145 = n23143 & n23144;
  assign n23146 = ~n23126 & ~n23134;
  assign n23147 = ~n23119 & n23146;
  assign n23148 = ~n23113 & n23147;
  assign n23149 = n23119 & ~n23126;
  assign n23150 = ~n23138 & ~n23149;
  assign n23151 = n23113 & ~n23150;
  assign n23152 = ~n23148 & ~n23151;
  assign n23153 = ~n23145 & n23152;
  assign n23154 = n23107 & ~n23153;
  assign n23155 = ~n23142 & ~n23154;
  assign n23156 = n23101 & ~n23155;
  assign n23157 = ~n23107 & ~n23113;
  assign n23158 = ~n23126 & n23157;
  assign n23159 = n23107 & n23138;
  assign n23160 = ~n23113 & n23159;
  assign n23161 = ~n23113 & ~n23119;
  assign n23162 = n23126 & n23161;
  assign n23163 = ~n23128 & ~n23162;
  assign n23164 = n23107 & ~n23163;
  assign n23165 = ~n23160 & ~n23164;
  assign n23166 = ~n23119 & n23138;
  assign n23167 = ~n23113 & n23166;
  assign n23168 = ~n23134 & n23143;
  assign n23169 = n23113 & n23168;
  assign n23170 = ~n23167 & ~n23169;
  assign n23171 = ~n23107 & n23113;
  assign n23172 = n23143 & n23171;
  assign n23173 = n23119 & n23146;
  assign n23174 = ~n23107 & n23173;
  assign n23175 = ~n23172 & ~n23174;
  assign n23176 = n23170 & n23175;
  assign n23177 = n23165 & n23176;
  assign n23178 = ~n23158 & n23177;
  assign n23179 = ~n23101 & ~n23178;
  assign n23180 = ~n23126 & n23134;
  assign n23181 = n23119 & n23180;
  assign n23182 = n23107 & ~n23113;
  assign n23183 = n23181 & n23182;
  assign n23184 = n23138 & n23182;
  assign n23185 = ~n23119 & n23184;
  assign n23186 = ~n23183 & ~n23185;
  assign n23187 = ~n23134 & n23149;
  assign n23188 = ~n23113 & n23187;
  assign n23189 = ~n23107 & n23188;
  assign n23190 = n23186 & ~n23189;
  assign n23191 = n23113 & n23135;
  assign n23192 = ~n23119 & n23180;
  assign n23193 = ~n23113 & n23192;
  assign n23194 = ~n23191 & ~n23193;
  assign n23195 = ~n23107 & ~n23194;
  assign n23196 = n23190 & ~n23195;
  assign n23197 = ~n23179 & n23196;
  assign n23198 = ~n23156 & n23197;
  assign n23199 = ~pi0291 & ~n23198;
  assign n23200 = pi0291 & n23198;
  assign po0306 = n23199 | n23200;
  assign n23202 = pi3175 & pi9040;
  assign n23203 = pi3154 & ~pi9040;
  assign n23204 = ~n23202 & ~n23203;
  assign n23205 = ~pi0278 & n23204;
  assign n23206 = pi0278 & ~n23204;
  assign n23207 = ~n23205 & ~n23206;
  assign n23208 = pi3156 & pi9040;
  assign n23209 = pi3224 & ~pi9040;
  assign n23210 = ~n23208 & ~n23209;
  assign n23211 = ~pi0277 & n23210;
  assign n23212 = pi0277 & ~n23210;
  assign n23213 = ~n23211 & ~n23212;
  assign n23214 = pi3147 & pi9040;
  assign n23215 = pi3308 & ~pi9040;
  assign n23216 = ~n23214 & ~n23215;
  assign n23217 = ~pi0276 & ~n23216;
  assign n23218 = pi0276 & n23216;
  assign n23219 = ~n23217 & ~n23218;
  assign n23220 = pi3224 & pi9040;
  assign n23221 = pi3167 & ~pi9040;
  assign n23222 = ~n23220 & ~n23221;
  assign n23223 = ~pi0251 & ~n23222;
  assign n23224 = pi0251 & n23222;
  assign n23225 = ~n23223 & ~n23224;
  assign n23226 = pi3198 & pi9040;
  assign n23227 = pi3159 & ~pi9040;
  assign n23228 = ~n23226 & ~n23227;
  assign n23229 = ~pi0255 & n23228;
  assign n23230 = pi0255 & ~n23228;
  assign n23231 = ~n23229 & ~n23230;
  assign n23232 = ~n23225 & n23231;
  assign n23233 = ~n23219 & n23232;
  assign n23234 = n23213 & n23233;
  assign n23235 = ~n23213 & ~n23219;
  assign n23236 = n23231 & n23235;
  assign n23237 = n23225 & n23236;
  assign n23238 = ~n23234 & ~n23237;
  assign n23239 = ~n23207 & ~n23238;
  assign n23240 = ~n23225 & ~n23231;
  assign n23241 = n23219 & n23240;
  assign n23242 = n23213 & n23241;
  assign n23243 = n23207 & n23242;
  assign n23244 = pi3155 & pi9040;
  assign n23245 = pi3198 & ~pi9040;
  assign n23246 = ~n23244 & ~n23245;
  assign n23247 = ~pi0286 & ~n23246;
  assign n23248 = pi0286 & ~n23244;
  assign n23249 = ~n23245 & n23248;
  assign n23250 = ~n23247 & ~n23249;
  assign n23251 = n23225 & n23231;
  assign n23252 = n23219 & n23251;
  assign n23253 = ~n23207 & n23252;
  assign n23254 = ~n23242 & ~n23253;
  assign n23255 = n23213 & n23225;
  assign n23256 = ~n23219 & n23255;
  assign n23257 = n23213 & n23219;
  assign n23258 = ~n23225 & n23257;
  assign n23259 = ~n23256 & ~n23258;
  assign n23260 = n23207 & ~n23259;
  assign n23261 = n23207 & ~n23213;
  assign n23262 = n23232 & n23261;
  assign n23263 = ~n23219 & n23262;
  assign n23264 = ~n23213 & n23219;
  assign n23265 = ~n23231 & n23264;
  assign n23266 = n23225 & n23265;
  assign n23267 = ~n23219 & n23240;
  assign n23268 = ~n23207 & n23267;
  assign n23269 = ~n23266 & ~n23268;
  assign n23270 = ~n23263 & n23269;
  assign n23271 = ~n23260 & n23270;
  assign n23272 = n23254 & n23271;
  assign n23273 = n23250 & ~n23272;
  assign n23274 = n23213 & n23253;
  assign n23275 = ~n23273 & ~n23274;
  assign n23276 = ~n23243 & n23275;
  assign n23277 = ~n23239 & n23276;
  assign n23278 = ~n23207 & ~n23213;
  assign n23279 = n23219 & ~n23225;
  assign n23280 = n23278 & n23279;
  assign n23281 = ~n23207 & n23233;
  assign n23282 = ~n23280 & ~n23281;
  assign n23283 = n23219 & n23232;
  assign n23284 = ~n23213 & n23283;
  assign n23285 = ~n23234 & ~n23284;
  assign n23286 = n23225 & ~n23231;
  assign n23287 = n23219 & n23286;
  assign n23288 = ~n23207 & n23287;
  assign n23289 = ~n23219 & n23286;
  assign n23290 = n23213 & n23289;
  assign n23291 = ~n23288 & ~n23290;
  assign n23292 = ~n23213 & n23251;
  assign n23293 = ~n23219 & ~n23231;
  assign n23294 = ~n23292 & ~n23293;
  assign n23295 = n23207 & ~n23294;
  assign n23296 = n23291 & ~n23295;
  assign n23297 = n23285 & n23296;
  assign n23298 = n23282 & n23297;
  assign n23299 = ~n23250 & ~n23298;
  assign n23300 = n23277 & ~n23299;
  assign n23301 = ~pi0293 & ~n23300;
  assign n23302 = pi0293 & n23277;
  assign n23303 = ~n23299 & n23302;
  assign po0307 = n23301 | n23303;
  assign n23305 = pi3145 & pi9040;
  assign n23306 = pi3134 & ~pi9040;
  assign n23307 = ~n23305 & ~n23306;
  assign n23308 = pi0254 & n23307;
  assign n23309 = ~pi0254 & ~n23307;
  assign n23310 = ~n23308 & ~n23309;
  assign n23311 = pi3296 & pi9040;
  assign n23312 = pi3176 & ~pi9040;
  assign n23313 = ~n23311 & ~n23312;
  assign n23314 = ~pi0262 & ~n23313;
  assign n23315 = pi0262 & ~n23311;
  assign n23316 = ~n23312 & n23315;
  assign n23317 = ~n23314 & ~n23316;
  assign n23318 = pi3148 & pi9040;
  assign n23319 = pi3240 & ~pi9040;
  assign n23320 = ~n23318 & ~n23319;
  assign n23321 = pi0271 & n23320;
  assign n23322 = ~pi0271 & ~n23320;
  assign n23323 = ~n23321 & ~n23322;
  assign n23324 = pi3132 & pi9040;
  assign n23325 = pi3129 & ~pi9040;
  assign n23326 = ~n23324 & ~n23325;
  assign n23327 = ~pi0266 & n23326;
  assign n23328 = pi0266 & ~n23326;
  assign n23329 = ~n23327 & ~n23328;
  assign n23330 = n23323 & ~n23329;
  assign n23331 = ~n23317 & n23330;
  assign n23332 = pi3183 & pi9040;
  assign n23333 = pi3194 & ~pi9040;
  assign n23334 = ~n23332 & ~n23333;
  assign n23335 = ~pi0287 & n23334;
  assign n23336 = pi0287 & ~n23334;
  assign n23337 = ~n23335 & ~n23336;
  assign n23338 = n23331 & n23337;
  assign n23339 = ~n23323 & n23329;
  assign n23340 = ~n23317 & n23339;
  assign n23341 = n23337 & n23340;
  assign n23342 = ~n23338 & ~n23341;
  assign n23343 = n23317 & ~n23337;
  assign n23344 = n23339 & n23343;
  assign n23345 = n23323 & n23329;
  assign n23346 = ~n23317 & n23345;
  assign n23347 = ~n23337 & n23346;
  assign n23348 = ~n23344 & ~n23347;
  assign n23349 = n23342 & n23348;
  assign n23350 = n23310 & ~n23349;
  assign n23351 = ~n23317 & ~n23337;
  assign n23352 = ~n23329 & n23351;
  assign n23353 = ~n23323 & n23352;
  assign n23354 = ~n23346 & ~n23353;
  assign n23355 = n23310 & ~n23354;
  assign n23356 = ~n23329 & n23337;
  assign n23357 = ~n23310 & n23356;
  assign n23358 = n23317 & n23323;
  assign n23359 = ~n23337 & n23339;
  assign n23360 = ~n23358 & ~n23359;
  assign n23361 = ~n23310 & ~n23360;
  assign n23362 = ~n23357 & ~n23361;
  assign n23363 = ~n23323 & ~n23329;
  assign n23364 = n23317 & n23363;
  assign n23365 = n23337 & n23364;
  assign n23366 = n23362 & ~n23365;
  assign n23367 = ~n23329 & n23358;
  assign n23368 = ~n23337 & n23367;
  assign n23369 = n23366 & ~n23368;
  assign n23370 = ~n23355 & n23369;
  assign n23371 = ~pi3132 & ~pi9040;
  assign n23372 = ~pi3181 & pi9040;
  assign n23373 = ~n23371 & ~n23372;
  assign n23374 = ~pi0273 & n23373;
  assign n23375 = pi0273 & ~n23373;
  assign n23376 = ~n23374 & ~n23375;
  assign n23377 = ~n23370 & ~n23376;
  assign n23378 = ~n23317 & ~n23329;
  assign n23379 = ~n23310 & ~n23337;
  assign n23380 = n23376 & n23379;
  assign n23381 = n23378 & n23380;
  assign n23382 = ~n23317 & n23337;
  assign n23383 = n23329 & n23382;
  assign n23384 = ~n23310 & ~n23383;
  assign n23385 = ~n23323 & n23343;
  assign n23386 = ~n23330 & ~n23378;
  assign n23387 = n23337 & ~n23386;
  assign n23388 = n23317 & n23339;
  assign n23389 = ~n23387 & ~n23388;
  assign n23390 = ~n23385 & n23389;
  assign n23391 = n23310 & n23390;
  assign n23392 = ~n23384 & ~n23391;
  assign n23393 = n23317 & n23345;
  assign n23394 = ~n23337 & n23393;
  assign n23395 = ~n23392 & ~n23394;
  assign n23396 = n23376 & ~n23395;
  assign n23397 = ~n23381 & ~n23396;
  assign n23398 = ~n23377 & n23397;
  assign n23399 = ~n23350 & n23398;
  assign n23400 = ~n23310 & n23365;
  assign n23401 = n23399 & ~n23400;
  assign n23402 = pi0288 & ~n23401;
  assign n23403 = ~pi0288 & ~n23400;
  assign n23404 = n23398 & n23403;
  assign n23405 = ~n23350 & n23404;
  assign po0310 = n23402 | n23405;
  assign n23407 = ~n23207 & n23240;
  assign n23408 = n23213 & n23407;
  assign n23409 = ~n23219 & n23251;
  assign n23410 = n23225 & n23235;
  assign n23411 = ~n23409 & ~n23410;
  assign n23412 = ~n23207 & ~n23411;
  assign n23413 = ~n23408 & ~n23412;
  assign n23414 = n23207 & n23213;
  assign n23415 = n23286 & n23414;
  assign n23416 = n23207 & n23233;
  assign n23417 = ~n23415 & ~n23416;
  assign n23418 = n23413 & n23417;
  assign n23419 = n23225 & n23257;
  assign n23420 = ~n23234 & ~n23419;
  assign n23421 = ~n23284 & n23420;
  assign n23422 = n23418 & n23421;
  assign n23423 = ~n23250 & ~n23422;
  assign n23424 = ~n23274 & ~n23280;
  assign n23425 = ~n23242 & ~n23409;
  assign n23426 = ~n23292 & n23425;
  assign n23427 = n23207 & ~n23426;
  assign n23428 = ~n23231 & n23235;
  assign n23429 = ~n23225 & n23428;
  assign n23430 = ~n23266 & ~n23429;
  assign n23431 = ~n23207 & n23213;
  assign n23432 = n23289 & n23431;
  assign n23433 = n23430 & ~n23432;
  assign n23434 = ~n23207 & n23283;
  assign n23435 = n23433 & ~n23434;
  assign n23436 = ~n23427 & n23435;
  assign n23437 = n23250 & ~n23436;
  assign n23438 = ~n23234 & n23430;
  assign n23439 = n23207 & ~n23438;
  assign n23440 = ~n23437 & ~n23439;
  assign n23441 = n23424 & n23440;
  assign n23442 = ~n23423 & n23441;
  assign n23443 = pi0300 & ~n23442;
  assign n23444 = ~pi0300 & n23442;
  assign po0311 = n23443 | n23444;
  assign n23446 = ~n23101 & n23107;
  assign n23447 = ~n23113 & n23135;
  assign n23448 = ~n23113 & n23127;
  assign n23449 = n23113 & n23166;
  assign n23450 = ~n23448 & ~n23449;
  assign n23451 = ~n23447 & n23450;
  assign n23452 = n23446 & ~n23451;
  assign n23453 = ~n23113 & n23119;
  assign n23454 = n23134 & n23453;
  assign n23455 = n23113 & n23192;
  assign n23456 = ~n23454 & ~n23455;
  assign n23457 = ~n23136 & ~n23139;
  assign n23458 = n23456 & n23457;
  assign n23459 = ~n23107 & ~n23458;
  assign n23460 = n23113 & n23173;
  assign n23461 = ~n23459 & ~n23460;
  assign n23462 = ~n23101 & ~n23461;
  assign n23463 = ~n23452 & ~n23462;
  assign n23464 = ~n23119 & n23157;
  assign n23465 = ~n23134 & n23464;
  assign n23466 = ~n23140 & ~n23465;
  assign n23467 = ~n23135 & ~n23180;
  assign n23468 = n23113 & ~n23467;
  assign n23469 = ~n23181 & ~n23468;
  assign n23470 = n23107 & ~n23469;
  assign n23471 = ~n23147 & ~n23448;
  assign n23472 = ~n23449 & n23471;
  assign n23473 = ~n23107 & ~n23472;
  assign n23474 = ~n23470 & ~n23473;
  assign n23475 = n23113 & n23119;
  assign n23476 = n23134 & n23475;
  assign n23477 = ~n23126 & n23476;
  assign n23478 = ~n23169 & ~n23477;
  assign n23479 = ~n23188 & n23478;
  assign n23480 = ~n23160 & n23479;
  assign n23481 = n23474 & n23480;
  assign n23482 = n23101 & ~n23481;
  assign n23483 = n23466 & ~n23482;
  assign n23484 = n23463 & n23483;
  assign n23485 = pi0290 & ~n23484;
  assign n23486 = ~pi0290 & n23484;
  assign po0312 = n23485 | n23486;
  assign n23488 = ~n23213 & n23252;
  assign n23489 = n23213 & n23283;
  assign n23490 = ~n23488 & ~n23489;
  assign n23491 = ~n23213 & n23241;
  assign n23492 = ~n23213 & n23286;
  assign n23493 = n23213 & n23267;
  assign n23494 = ~n23492 & ~n23493;
  assign n23495 = n23207 & ~n23494;
  assign n23496 = ~n23491 & ~n23495;
  assign n23497 = ~n23213 & n23407;
  assign n23498 = ~n23281 & ~n23497;
  assign n23499 = n23496 & n23498;
  assign n23500 = n23490 & n23499;
  assign n23501 = n23250 & ~n23500;
  assign n23502 = n23207 & ~n23250;
  assign n23503 = ~n23225 & n23235;
  assign n23504 = ~n23219 & n23231;
  assign n23505 = ~n23503 & ~n23504;
  assign n23506 = n23502 & ~n23505;
  assign n23507 = n23213 & n23409;
  assign n23508 = n23207 & n23507;
  assign n23509 = n23213 & n23287;
  assign n23510 = ~n23489 & ~n23509;
  assign n23511 = n23207 & ~n23510;
  assign n23512 = ~n23508 & ~n23511;
  assign n23513 = ~n23242 & ~n23256;
  assign n23514 = n23219 & n23278;
  assign n23515 = ~n23240 & n23514;
  assign n23516 = ~n23253 & ~n23515;
  assign n23517 = n23513 & n23516;
  assign n23518 = ~n23250 & ~n23517;
  assign n23519 = n23241 & n23431;
  assign n23520 = ~n23518 & ~n23519;
  assign n23521 = n23512 & n23520;
  assign n23522 = ~n23506 & n23521;
  assign n23523 = ~n23501 & n23522;
  assign n23524 = ~n23432 & n23523;
  assign n23525 = ~pi0310 & ~n23524;
  assign n23526 = ~n23432 & n23522;
  assign n23527 = pi0310 & n23526;
  assign n23528 = ~n23501 & n23527;
  assign po0314 = n23525 | n23528;
  assign n23530 = ~n23147 & ~n23181;
  assign n23531 = n23107 & ~n23530;
  assign n23532 = n23113 & n23136;
  assign n23533 = ~n23531 & ~n23532;
  assign n23534 = n23113 & n23126;
  assign n23535 = ~n23143 & ~n23534;
  assign n23536 = ~n23192 & n23535;
  assign n23537 = ~n23107 & ~n23536;
  assign n23538 = n23533 & ~n23537;
  assign n23539 = ~n23101 & ~n23538;
  assign n23540 = ~n23113 & n23168;
  assign n23541 = n23107 & n23540;
  assign n23542 = ~n23185 & ~n23541;
  assign n23543 = ~n23189 & n23542;
  assign n23544 = ~n23107 & n23126;
  assign n23545 = n23161 & n23544;
  assign n23546 = n23113 & n23147;
  assign n23547 = n23107 & n23143;
  assign n23548 = ~n23546 & ~n23547;
  assign n23549 = ~n23477 & n23548;
  assign n23550 = ~n23545 & n23549;
  assign n23551 = n23134 & n23161;
  assign n23552 = ~n23188 & ~n23551;
  assign n23553 = n23550 & n23552;
  assign n23554 = ~n23174 & n23553;
  assign n23555 = n23101 & ~n23554;
  assign n23556 = n23543 & ~n23555;
  assign n23557 = ~n23539 & n23556;
  assign n23558 = ~pi0296 & ~n23557;
  assign n23559 = pi0296 & n23543;
  assign n23560 = ~n23539 & n23559;
  assign n23561 = ~n23555 & n23560;
  assign po0315 = n23558 | n23561;
  assign n23563 = ~n23488 & ~n23503;
  assign n23564 = n23250 & ~n23563;
  assign n23565 = n23207 & n23241;
  assign n23566 = ~n23231 & n23257;
  assign n23567 = ~n23258 & ~n23566;
  assign n23568 = n23207 & ~n23567;
  assign n23569 = ~n23565 & ~n23568;
  assign n23570 = n23250 & ~n23569;
  assign n23571 = ~n23564 & ~n23570;
  assign n23572 = n23252 & n23261;
  assign n23573 = ~n23263 & ~n23572;
  assign n23574 = ~n23256 & ~n23293;
  assign n23575 = ~n23207 & ~n23574;
  assign n23576 = n23250 & n23575;
  assign n23577 = n23573 & ~n23576;
  assign n23578 = n23231 & n23257;
  assign n23579 = n23225 & n23578;
  assign n23580 = n23213 & n23232;
  assign n23581 = ~n23237 & ~n23580;
  assign n23582 = ~n23207 & ~n23581;
  assign n23583 = ~n23242 & ~n23266;
  assign n23584 = n23213 & n23251;
  assign n23585 = ~n23289 & ~n23584;
  assign n23586 = n23207 & ~n23585;
  assign n23587 = n23583 & ~n23586;
  assign n23588 = ~n23582 & n23587;
  assign n23589 = ~n23579 & n23588;
  assign n23590 = ~n23250 & ~n23589;
  assign n23591 = ~n23284 & n23430;
  assign n23592 = ~n23207 & ~n23591;
  assign n23593 = ~n23590 & ~n23592;
  assign n23594 = n23577 & n23593;
  assign n23595 = n23571 & n23594;
  assign n23596 = ~pi0306 & ~n23595;
  assign n23597 = pi0306 & n23577;
  assign n23598 = n23571 & n23597;
  assign n23599 = n23593 & n23598;
  assign po0323 = n23596 | n23599;
  assign n23601 = pi3235 & pi9040;
  assign n23602 = pi3145 & ~pi9040;
  assign n23603 = ~n23601 & ~n23602;
  assign n23604 = pi0256 & n23603;
  assign n23605 = ~pi0256 & ~n23603;
  assign n23606 = ~n23604 & ~n23605;
  assign n23607 = pi3176 & pi9040;
  assign n23608 = pi3158 & ~pi9040;
  assign n23609 = ~n23607 & ~n23608;
  assign n23610 = ~pi0282 & n23609;
  assign n23611 = pi0282 & ~n23609;
  assign n23612 = ~n23610 & ~n23611;
  assign n23613 = pi3139 & pi9040;
  assign n23614 = pi3151 & ~pi9040;
  assign n23615 = ~n23613 & ~n23614;
  assign n23616 = ~pi0286 & ~n23615;
  assign n23617 = pi0286 & ~n23613;
  assign n23618 = ~n23614 & n23617;
  assign n23619 = ~n23616 & ~n23618;
  assign n23620 = pi3174 & pi9040;
  assign n23621 = pi3139 & ~pi9040;
  assign n23622 = ~n23620 & ~n23621;
  assign n23623 = ~pi0255 & n23622;
  assign n23624 = pi0255 & ~n23622;
  assign n23625 = ~n23623 & ~n23624;
  assign n23626 = pi3150 & pi9040;
  assign n23627 = pi3251 & ~pi9040;
  assign n23628 = ~n23626 & ~n23627;
  assign n23629 = pi0279 & n23628;
  assign n23630 = ~pi0279 & ~n23628;
  assign n23631 = ~n23629 & ~n23630;
  assign n23632 = ~n23625 & ~n23631;
  assign n23633 = n23619 & n23632;
  assign n23634 = ~n23612 & n23633;
  assign n23635 = n23612 & ~n23625;
  assign n23636 = n23631 & n23635;
  assign n23637 = pi3128 & pi9040;
  assign n23638 = pi3142 & ~pi9040;
  assign n23639 = ~n23637 & ~n23638;
  assign n23640 = ~pi0270 & n23639;
  assign n23641 = pi0270 & ~n23639;
  assign n23642 = ~n23640 & ~n23641;
  assign n23643 = ~n23619 & n23635;
  assign n23644 = n23619 & n23631;
  assign n23645 = n23625 & n23644;
  assign n23646 = ~n23643 & ~n23645;
  assign n23647 = n23642 & ~n23646;
  assign n23648 = ~n23636 & ~n23647;
  assign n23649 = ~n23625 & n23644;
  assign n23650 = ~n23619 & n23625;
  assign n23651 = n23625 & ~n23631;
  assign n23652 = n23612 & n23651;
  assign n23653 = ~n23619 & ~n23631;
  assign n23654 = ~n23612 & n23653;
  assign n23655 = ~n23652 & ~n23654;
  assign n23656 = ~n23650 & n23655;
  assign n23657 = ~n23649 & n23656;
  assign n23658 = ~n23642 & ~n23657;
  assign n23659 = n23648 & ~n23658;
  assign n23660 = ~n23634 & n23659;
  assign n23661 = n23606 & ~n23660;
  assign n23662 = ~n23619 & n23631;
  assign n23663 = n23625 & n23662;
  assign n23664 = n23612 & n23663;
  assign n23665 = n23625 & n23653;
  assign n23666 = ~n23612 & n23665;
  assign n23667 = ~n23634 & ~n23666;
  assign n23668 = ~n23664 & n23667;
  assign n23669 = ~n23642 & ~n23668;
  assign n23670 = ~n23661 & ~n23669;
  assign n23671 = n23612 & n23649;
  assign n23672 = n23625 & n23642;
  assign n23673 = n23619 & n23672;
  assign n23674 = ~n23612 & n23673;
  assign n23675 = n23612 & ~n23642;
  assign n23676 = n23632 & n23675;
  assign n23677 = ~n23625 & n23662;
  assign n23678 = ~n23612 & n23677;
  assign n23679 = ~n23676 & ~n23678;
  assign n23680 = ~n23619 & ~n23625;
  assign n23681 = ~n23612 & n23680;
  assign n23682 = n23619 & ~n23631;
  assign n23683 = n23625 & n23682;
  assign n23684 = ~n23681 & ~n23683;
  assign n23685 = n23642 & ~n23684;
  assign n23686 = n23642 & n23650;
  assign n23687 = n23612 & n23686;
  assign n23688 = ~n23685 & ~n23687;
  assign n23689 = n23679 & n23688;
  assign n23690 = ~n23606 & ~n23689;
  assign n23691 = ~n23674 & ~n23690;
  assign n23692 = ~n23671 & n23691;
  assign n23693 = n23670 & n23692;
  assign n23694 = ~pi0309 & ~n23693;
  assign n23695 = ~n23661 & ~n23671;
  assign n23696 = ~n23669 & n23695;
  assign n23697 = n23691 & n23696;
  assign n23698 = pi0309 & n23697;
  assign po0326 = n23694 | n23698;
  assign n23700 = ~n23113 & ~n23126;
  assign n23701 = ~n23551 & ~n23700;
  assign n23702 = n23107 & ~n23701;
  assign n23703 = n23113 & ~n23119;
  assign n23704 = ~n23134 & n23703;
  assign n23705 = ~n23702 & ~n23704;
  assign n23706 = ~n23107 & n23135;
  assign n23707 = ~n23113 & n23706;
  assign n23708 = ~n23193 & ~n23707;
  assign n23709 = n23705 & n23708;
  assign n23710 = n23101 & ~n23709;
  assign n23711 = ~n23166 & ~n23169;
  assign n23712 = ~n23113 & n23146;
  assign n23713 = n23711 & ~n23712;
  assign n23714 = ~n23107 & ~n23713;
  assign n23715 = n23135 & n23182;
  assign n23716 = ~n23140 & ~n23715;
  assign n23717 = ~n23714 & n23716;
  assign n23718 = ~n23192 & ~n23460;
  assign n23719 = n23107 & ~n23718;
  assign n23720 = n23717 & ~n23719;
  assign n23721 = ~n23101 & ~n23720;
  assign n23722 = ~n23710 & ~n23721;
  assign n23723 = ~n23113 & n23180;
  assign n23724 = n23113 & ~n23457;
  assign n23725 = ~n23723 & ~n23724;
  assign n23726 = n23107 & ~n23725;
  assign n23727 = ~n23166 & n23530;
  assign n23728 = n23171 & ~n23727;
  assign n23729 = ~n23726 & ~n23728;
  assign n23730 = n23722 & n23729;
  assign n23731 = ~pi0295 & ~n23730;
  assign n23732 = ~n23721 & n23729;
  assign n23733 = pi0295 & n23732;
  assign n23734 = ~n23710 & n23733;
  assign po0328 = n23731 | n23734;
  assign n23736 = pi3152 & pi9040;
  assign n23737 = pi3196 & ~pi9040;
  assign n23738 = ~n23736 & ~n23737;
  assign n23739 = ~pi0266 & ~n23738;
  assign n23740 = pi0266 & n23738;
  assign n23741 = ~n23739 & ~n23740;
  assign n23742 = pi3251 & pi9040;
  assign n23743 = pi3136 & ~pi9040;
  assign n23744 = ~n23742 & ~n23743;
  assign n23745 = ~pi0285 & ~n23744;
  assign n23746 = pi0285 & n23744;
  assign n23747 = ~n23745 & ~n23746;
  assign n23748 = pi3134 & pi9040;
  assign n23749 = pi3296 & ~pi9040;
  assign n23750 = ~n23748 & ~n23749;
  assign n23751 = ~pi0262 & n23750;
  assign n23752 = pi0262 & ~n23750;
  assign n23753 = ~n23751 & ~n23752;
  assign n23754 = ~n23747 & ~n23753;
  assign n23755 = pi3194 & pi9040;
  assign n23756 = pi3179 & ~pi9040;
  assign n23757 = ~n23755 & ~n23756;
  assign n23758 = pi0265 & n23757;
  assign n23759 = ~pi0265 & ~n23757;
  assign n23760 = ~n23758 & ~n23759;
  assign n23761 = pi3179 & pi9040;
  assign n23762 = pi3182 & ~pi9040;
  assign n23763 = ~n23761 & ~n23762;
  assign n23764 = ~pi0281 & n23763;
  assign n23765 = pi0281 & ~n23763;
  assign n23766 = ~n23764 & ~n23765;
  assign n23767 = ~n23760 & n23766;
  assign n23768 = n23754 & n23767;
  assign n23769 = pi3240 & pi9040;
  assign n23770 = pi3130 & ~pi9040;
  assign n23771 = ~n23769 & ~n23770;
  assign n23772 = ~pi0272 & ~n23771;
  assign n23773 = pi0272 & n23771;
  assign n23774 = ~n23772 & ~n23773;
  assign n23775 = n23747 & n23753;
  assign n23776 = n23774 & n23775;
  assign n23777 = n23753 & ~n23774;
  assign n23778 = ~n23747 & n23777;
  assign n23779 = n23760 & n23778;
  assign n23780 = ~n23776 & ~n23779;
  assign n23781 = n23747 & ~n23753;
  assign n23782 = n23760 & n23781;
  assign n23783 = n23780 & ~n23782;
  assign n23784 = n23766 & ~n23783;
  assign n23785 = n23747 & ~n23774;
  assign n23786 = ~n23760 & ~n23766;
  assign n23787 = n23785 & n23786;
  assign n23788 = ~n23774 & n23775;
  assign n23789 = ~n23760 & n23788;
  assign n23790 = ~n23787 & ~n23789;
  assign n23791 = ~n23784 & n23790;
  assign n23792 = ~n23768 & n23791;
  assign n23793 = n23754 & n23774;
  assign n23794 = ~n23760 & n23793;
  assign n23795 = n23774 & n23781;
  assign n23796 = n23760 & n23795;
  assign n23797 = ~n23794 & ~n23796;
  assign n23798 = n23792 & n23797;
  assign n23799 = ~n23741 & ~n23798;
  assign n23800 = ~n23760 & ~n23774;
  assign n23801 = ~n23753 & n23800;
  assign n23802 = n23747 & n23801;
  assign n23803 = ~n23793 & ~n23802;
  assign n23804 = n23766 & ~n23803;
  assign n23805 = n23754 & ~n23774;
  assign n23806 = n23760 & n23805;
  assign n23807 = ~n23760 & n23777;
  assign n23808 = ~n23747 & n23807;
  assign n23809 = ~n23806 & ~n23808;
  assign n23810 = n23760 & ~n23774;
  assign n23811 = n23747 & n23810;
  assign n23812 = ~n23760 & n23795;
  assign n23813 = ~n23811 & ~n23812;
  assign n23814 = ~n23766 & ~n23813;
  assign n23815 = n23809 & ~n23814;
  assign n23816 = ~n23804 & n23815;
  assign n23817 = n23741 & ~n23816;
  assign n23818 = ~n23747 & n23753;
  assign n23819 = n23774 & n23818;
  assign n23820 = n23760 & n23819;
  assign n23821 = ~n23788 & ~n23820;
  assign n23822 = ~n23806 & n23821;
  assign n23823 = ~n23766 & ~n23822;
  assign n23824 = ~n23747 & n23774;
  assign n23825 = ~n23760 & n23824;
  assign n23826 = n23747 & n23774;
  assign n23827 = n23760 & n23826;
  assign n23828 = ~n23825 & ~n23827;
  assign n23829 = n23766 & ~n23828;
  assign n23830 = ~n23823 & ~n23829;
  assign n23831 = ~n23766 & n23777;
  assign n23832 = ~n23760 & n23831;
  assign n23833 = n23830 & ~n23832;
  assign n23834 = ~n23817 & n23833;
  assign n23835 = ~n23799 & n23834;
  assign n23836 = ~pi0292 & ~n23835;
  assign n23837 = pi0292 & n23835;
  assign po0331 = n23836 | n23837;
  assign n23839 = pi3143 & pi9040;
  assign n23840 = pi3195 & ~pi9040;
  assign n23841 = ~n23839 & ~n23840;
  assign n23842 = pi0275 & n23841;
  assign n23843 = ~pi0275 & ~n23841;
  assign n23844 = ~n23842 & ~n23843;
  assign n23845 = pi3166 & pi9040;
  assign n23846 = pi3177 & ~pi9040;
  assign n23847 = ~n23845 & ~n23846;
  assign n23848 = ~pi0271 & n23847;
  assign n23849 = pi0271 & ~n23847;
  assign n23850 = ~n23848 & ~n23849;
  assign n23851 = pi3178 & pi9040;
  assign n23852 = pi3140 & ~pi9040;
  assign n23853 = ~n23851 & ~n23852;
  assign n23854 = ~pi0273 & n23853;
  assign n23855 = pi0273 & ~n23853;
  assign n23856 = ~n23854 & ~n23855;
  assign n23857 = pi3167 & pi9040;
  assign n23858 = pi3227 & ~pi9040;
  assign n23859 = ~n23857 & ~n23858;
  assign n23860 = ~pi0250 & n23859;
  assign n23861 = pi0250 & ~n23859;
  assign n23862 = ~n23860 & ~n23861;
  assign n23863 = n23856 & ~n23862;
  assign n23864 = pi3133 & pi9040;
  assign n23865 = pi3141 & ~pi9040;
  assign n23866 = ~n23864 & ~n23865;
  assign n23867 = pi0263 & n23866;
  assign n23868 = ~pi0263 & ~n23866;
  assign n23869 = ~n23867 & ~n23868;
  assign n23870 = pi3308 & pi9040;
  assign n23871 = pi3155 & ~pi9040;
  assign n23872 = ~n23870 & ~n23871;
  assign n23873 = ~pi0283 & n23872;
  assign n23874 = pi0283 & ~n23872;
  assign n23875 = ~n23873 & ~n23874;
  assign n23876 = n23869 & ~n23875;
  assign n23877 = n23863 & n23876;
  assign n23878 = ~n23850 & n23877;
  assign n23879 = ~n23869 & ~n23875;
  assign n23880 = ~n23856 & ~n23862;
  assign n23881 = n23879 & n23880;
  assign n23882 = n23856 & n23862;
  assign n23883 = ~n23850 & n23882;
  assign n23884 = ~n23869 & n23883;
  assign n23885 = ~n23856 & n23862;
  assign n23886 = ~n23850 & n23885;
  assign n23887 = ~n23875 & n23886;
  assign n23888 = n23869 & n23887;
  assign n23889 = ~n23884 & ~n23888;
  assign n23890 = ~n23881 & n23889;
  assign n23891 = ~n23878 & n23890;
  assign n23892 = n23850 & ~n23869;
  assign n23893 = ~n23862 & n23892;
  assign n23894 = ~n23856 & n23893;
  assign n23895 = n23891 & ~n23894;
  assign n23896 = ~n23844 & ~n23895;
  assign n23897 = n23850 & n23862;
  assign n23898 = ~n23856 & n23897;
  assign n23899 = n23869 & n23875;
  assign n23900 = n23898 & n23899;
  assign n23901 = ~n23850 & ~n23869;
  assign n23902 = n23856 & n23901;
  assign n23903 = ~n23869 & n23882;
  assign n23904 = ~n23902 & ~n23903;
  assign n23905 = n23875 & ~n23904;
  assign n23906 = ~n23900 & ~n23905;
  assign n23907 = ~n23844 & ~n23906;
  assign n23908 = n23862 & n23901;
  assign n23909 = ~n23850 & ~n23856;
  assign n23910 = ~n23862 & n23909;
  assign n23911 = n23869 & n23910;
  assign n23912 = ~n23908 & ~n23911;
  assign n23913 = n23850 & n23863;
  assign n23914 = n23869 & n23913;
  assign n23915 = n23912 & ~n23914;
  assign n23916 = n23875 & ~n23915;
  assign n23917 = ~n23907 & ~n23916;
  assign n23918 = ~n23896 & n23917;
  assign n23919 = n23850 & n23869;
  assign n23920 = ~n23875 & n23919;
  assign n23921 = n23882 & n23920;
  assign n23922 = n23850 & ~n23856;
  assign n23923 = n23879 & n23922;
  assign n23924 = n23875 & n23909;
  assign n23925 = n23856 & n23869;
  assign n23926 = n23850 & n23925;
  assign n23927 = ~n23913 & ~n23926;
  assign n23928 = ~n23924 & n23927;
  assign n23929 = ~n23869 & n23898;
  assign n23930 = n23928 & ~n23929;
  assign n23931 = n23863 & ~n23875;
  assign n23932 = ~n23869 & n23931;
  assign n23933 = n23850 & ~n23862;
  assign n23934 = n23869 & n23882;
  assign n23935 = ~n23933 & ~n23934;
  assign n23936 = ~n23875 & ~n23935;
  assign n23937 = ~n23932 & ~n23936;
  assign n23938 = n23930 & n23937;
  assign n23939 = n23844 & ~n23938;
  assign n23940 = ~n23923 & ~n23939;
  assign n23941 = ~n23921 & n23940;
  assign n23942 = n23918 & n23941;
  assign n23943 = pi0299 & n23942;
  assign n23944 = ~pi0299 & ~n23942;
  assign po0332 = n23943 | n23944;
  assign n23946 = n23753 & n23810;
  assign n23947 = n23747 & n23946;
  assign n23948 = ~n23808 & ~n23826;
  assign n23949 = ~n23766 & ~n23948;
  assign n23950 = ~n23947 & ~n23949;
  assign n23951 = ~n23802 & n23950;
  assign n23952 = n23760 & n23766;
  assign n23953 = n23805 & n23952;
  assign n23954 = ~n23794 & ~n23953;
  assign n23955 = ~n23820 & n23954;
  assign n23956 = n23951 & n23955;
  assign n23957 = n23741 & ~n23956;
  assign n23958 = ~n23774 & n23781;
  assign n23959 = n23760 & n23958;
  assign n23960 = ~n23779 & ~n23959;
  assign n23961 = ~n23760 & n23819;
  assign n23962 = ~n23789 & ~n23961;
  assign n23963 = ~n23766 & n23805;
  assign n23964 = n23760 & n23793;
  assign n23965 = ~n23963 & ~n23964;
  assign n23966 = ~n23753 & n23774;
  assign n23967 = n23747 & n23760;
  assign n23968 = ~n23966 & ~n23967;
  assign n23969 = ~n23777 & n23968;
  assign n23970 = n23766 & ~n23969;
  assign n23971 = n23965 & ~n23970;
  assign n23972 = n23962 & n23971;
  assign n23973 = n23960 & n23972;
  assign n23974 = ~n23741 & ~n23973;
  assign n23975 = ~n23957 & ~n23974;
  assign n23976 = pi0289 & ~n23975;
  assign n23977 = ~pi0289 & ~n23957;
  assign n23978 = ~n23974 & n23977;
  assign po0333 = n23976 | n23978;
  assign n23980 = ~n23850 & n23856;
  assign n23981 = ~n23894 & ~n23980;
  assign n23982 = ~n23925 & n23981;
  assign n23983 = ~n23875 & ~n23982;
  assign n23984 = ~n23856 & n23899;
  assign n23985 = ~n23850 & n23869;
  assign n23986 = ~n23862 & n23985;
  assign n23987 = ~n23869 & n23886;
  assign n23988 = ~n23986 & ~n23987;
  assign n23989 = n23850 & n23856;
  assign n23990 = ~n23869 & n23875;
  assign n23991 = n23989 & n23990;
  assign n23992 = n23988 & ~n23991;
  assign n23993 = ~n23984 & n23992;
  assign n23994 = ~n23983 & n23993;
  assign n23995 = n23844 & ~n23994;
  assign n23996 = ~n23850 & n23863;
  assign n23997 = ~n23869 & n23996;
  assign n23998 = n23869 & n23883;
  assign n23999 = ~n23997 & ~n23998;
  assign n24000 = ~n23875 & ~n23999;
  assign n24001 = ~n23995 & ~n24000;
  assign n24002 = n23869 & n23886;
  assign n24003 = ~n23898 & ~n23910;
  assign n24004 = ~n23875 & ~n24003;
  assign n24005 = ~n24002 & ~n24004;
  assign n24006 = ~n23914 & n24005;
  assign n24007 = ~n23844 & ~n24006;
  assign n24008 = ~n23880 & ~n23882;
  assign n24009 = n23850 & ~n24008;
  assign n24010 = ~n23903 & ~n24009;
  assign n24011 = n23875 & ~n24010;
  assign n24012 = ~n23844 & n24011;
  assign n24013 = ~n24007 & ~n24012;
  assign n24014 = n24001 & n24013;
  assign n24015 = pi0301 & ~n24014;
  assign n24016 = ~pi0301 & n24001;
  assign n24017 = n24013 & n24016;
  assign po0334 = n24015 | n24017;
  assign n24019 = n23612 & n23642;
  assign n24020 = n23619 & n24019;
  assign n24021 = ~n23625 & n23653;
  assign n24022 = ~n23612 & n24021;
  assign n24023 = ~n23612 & n23663;
  assign n24024 = ~n24022 & ~n24023;
  assign n24025 = n23612 & n23665;
  assign n24026 = ~n23645 & ~n24025;
  assign n24027 = ~n23642 & ~n24026;
  assign n24028 = n24024 & ~n24027;
  assign n24029 = ~n24020 & n24028;
  assign n24030 = n23606 & ~n24029;
  assign n24031 = ~n23612 & n23619;
  assign n24032 = n23625 & n24031;
  assign n24033 = ~n23631 & n24032;
  assign n24034 = n23642 & n24033;
  assign n24035 = n23675 & n23683;
  assign n24036 = ~n23643 & ~n24035;
  assign n24037 = ~n23645 & ~n23677;
  assign n24038 = n23612 & n23662;
  assign n24039 = n24037 & ~n24038;
  assign n24040 = n23642 & ~n24039;
  assign n24041 = ~n23642 & n23649;
  assign n24042 = n23667 & ~n24041;
  assign n24043 = ~n24040 & n24042;
  assign n24044 = n24036 & n24043;
  assign n24045 = ~n23606 & ~n24044;
  assign n24046 = ~n24034 & ~n24045;
  assign n24047 = ~n24030 & n24046;
  assign n24048 = n23675 & n23677;
  assign n24049 = n23632 & ~n23642;
  assign n24050 = ~n23612 & n24049;
  assign n24051 = ~n24048 & ~n24050;
  assign n24052 = ~n23642 & n24023;
  assign n24053 = n24051 & ~n24052;
  assign n24054 = n24047 & n24053;
  assign n24055 = ~pi0297 & ~n24054;
  assign n24056 = pi0297 & n24053;
  assign n24057 = n24046 & n24056;
  assign n24058 = ~n24030 & n24057;
  assign po0335 = n24055 | n24058;
  assign n24060 = ~n23631 & n23635;
  assign n24061 = ~n23619 & n24060;
  assign n24062 = ~n23663 & ~n23671;
  assign n24063 = ~n23612 & n23632;
  assign n24064 = n23612 & n23683;
  assign n24065 = ~n24063 & ~n24064;
  assign n24066 = n24062 & n24065;
  assign n24067 = n23642 & ~n24066;
  assign n24068 = ~n23612 & n23644;
  assign n24069 = ~n23643 & ~n24068;
  assign n24070 = ~n23665 & n24069;
  assign n24071 = ~n23642 & ~n24070;
  assign n24072 = ~n23612 & n23625;
  assign n24073 = n23631 & n24072;
  assign n24074 = n23619 & n24073;
  assign n24075 = ~n24071 & ~n24074;
  assign n24076 = ~n24067 & n24075;
  assign n24077 = ~n24061 & n24076;
  assign n24078 = ~n23606 & ~n24077;
  assign n24079 = ~n23612 & n23642;
  assign n24080 = n23649 & n24079;
  assign n24081 = n23642 & n23665;
  assign n24082 = n23642 & n23677;
  assign n24083 = ~n24081 & ~n24082;
  assign n24084 = n23612 & ~n24083;
  assign n24085 = ~n24080 & ~n24084;
  assign n24086 = n23612 & n23633;
  assign n24087 = ~n24033 & ~n24086;
  assign n24088 = ~n23612 & n23662;
  assign n24089 = n23612 & n23644;
  assign n24090 = ~n24088 & ~n24089;
  assign n24091 = ~n23633 & n24090;
  assign n24092 = ~n23663 & n24091;
  assign n24093 = ~n23642 & ~n24092;
  assign n24094 = n23612 & n23645;
  assign n24095 = ~n24093 & ~n24094;
  assign n24096 = n24087 & n24095;
  assign n24097 = n24085 & n24096;
  assign n24098 = n23606 & ~n24097;
  assign n24099 = n23642 & ~n24024;
  assign n24100 = ~n24098 & ~n24099;
  assign n24101 = ~n23666 & ~n24086;
  assign n24102 = ~n23642 & ~n24101;
  assign n24103 = n24100 & ~n24102;
  assign n24104 = ~n24078 & n24103;
  assign n24105 = pi0307 & ~n24104;
  assign n24106 = ~pi0307 & n24104;
  assign po0336 = n24105 | n24106;
  assign n24108 = pi3177 & pi9040;
  assign n24109 = pi3161 & ~pi9040;
  assign n24110 = ~n24108 & ~n24109;
  assign n24111 = pi0269 & n24110;
  assign n24112 = ~pi0269 & ~n24110;
  assign n24113 = ~n24111 & ~n24112;
  assign n24114 = pi3140 & pi9040;
  assign n24115 = pi3175 & ~pi9040;
  assign n24116 = ~n24114 & ~n24115;
  assign n24117 = pi0275 & n24116;
  assign n24118 = ~pi0275 & ~n24116;
  assign n24119 = ~n24117 & ~n24118;
  assign n24120 = pi3149 & pi9040;
  assign n24121 = pi3156 & ~pi9040;
  assign n24122 = ~n24120 & ~n24121;
  assign n24123 = pi0274 & n24122;
  assign n24124 = ~pi0274 & ~n24122;
  assign n24125 = ~n24123 & ~n24124;
  assign n24126 = n24119 & ~n24125;
  assign n24127 = pi3138 & pi9040;
  assign n24128 = pi3146 & ~pi9040;
  assign n24129 = ~n24127 & ~n24128;
  assign n24130 = ~pi0284 & n24129;
  assign n24131 = pi0284 & ~n24129;
  assign n24132 = ~n24130 & ~n24131;
  assign n24133 = pi3141 & pi9040;
  assign n24134 = pi3166 & ~pi9040;
  assign n24135 = ~n24133 & ~n24134;
  assign n24136 = ~pi0250 & n24135;
  assign n24137 = pi0250 & ~n24135;
  assign n24138 = ~n24136 & ~n24137;
  assign n24139 = ~n24132 & ~n24138;
  assign n24140 = n24126 & n24139;
  assign n24141 = ~n24132 & n24138;
  assign n24142 = ~n24119 & n24141;
  assign n24143 = ~n24140 & ~n24142;
  assign n24144 = ~n24113 & ~n24143;
  assign n24145 = pi3135 & pi9040;
  assign n24146 = pi3149 & ~pi9040;
  assign n24147 = ~n24145 & ~n24146;
  assign n24148 = ~pi0280 & ~n24147;
  assign n24149 = pi0280 & n24147;
  assign n24150 = ~n24148 & ~n24149;
  assign n24151 = n24113 & n24132;
  assign n24152 = n24119 & n24151;
  assign n24153 = n24126 & n24138;
  assign n24154 = n24119 & n24125;
  assign n24155 = ~n24138 & n24154;
  assign n24156 = ~n24153 & ~n24155;
  assign n24157 = ~n24119 & ~n24125;
  assign n24158 = ~n24138 & n24157;
  assign n24159 = ~n24132 & n24158;
  assign n24160 = n24156 & ~n24159;
  assign n24161 = n24113 & ~n24160;
  assign n24162 = ~n24152 & ~n24161;
  assign n24163 = ~n24119 & n24125;
  assign n24164 = n24138 & n24163;
  assign n24165 = ~n24132 & n24164;
  assign n24166 = n24162 & ~n24165;
  assign n24167 = n24132 & n24157;
  assign n24168 = ~n24119 & ~n24138;
  assign n24169 = n24125 & n24168;
  assign n24170 = ~n24167 & ~n24169;
  assign n24171 = ~n24113 & ~n24170;
  assign n24172 = n24138 & n24154;
  assign n24173 = n24132 & n24172;
  assign n24174 = ~n24171 & ~n24173;
  assign n24175 = n24166 & n24174;
  assign n24176 = n24150 & ~n24175;
  assign n24177 = ~n24144 & ~n24176;
  assign n24178 = n24113 & ~n24150;
  assign n24179 = ~n24170 & n24178;
  assign n24180 = n24138 & n24157;
  assign n24181 = ~n24172 & ~n24180;
  assign n24182 = ~n24132 & ~n24181;
  assign n24183 = ~n24140 & ~n24182;
  assign n24184 = ~n24150 & ~n24183;
  assign n24185 = ~n24179 & ~n24184;
  assign n24186 = ~n24113 & ~n24150;
  assign n24187 = n24126 & n24132;
  assign n24188 = ~n24164 & ~n24187;
  assign n24189 = n24119 & ~n24138;
  assign n24190 = n24188 & ~n24189;
  assign n24191 = n24186 & ~n24190;
  assign n24192 = n24185 & ~n24191;
  assign n24193 = n24177 & n24192;
  assign n24194 = ~pi0294 & ~n24193;
  assign n24195 = pi0294 & n24185;
  assign n24196 = n24177 & n24195;
  assign n24197 = ~n24191 & n24196;
  assign po0337 = n24194 | n24197;
  assign n24199 = ~n24113 & ~n24132;
  assign n24200 = ~n24157 & ~n24172;
  assign n24201 = n24199 & ~n24200;
  assign n24202 = ~n24113 & n24138;
  assign n24203 = n24157 & n24202;
  assign n24204 = ~n24201 & ~n24203;
  assign n24205 = n24150 & ~n24204;
  assign n24206 = n24132 & ~n24138;
  assign n24207 = n24125 & n24206;
  assign n24208 = n24119 & n24207;
  assign n24209 = ~n24189 & ~n24206;
  assign n24210 = n24113 & ~n24209;
  assign n24211 = n24132 & n24138;
  assign n24212 = ~n24125 & n24211;
  assign n24213 = n24119 & n24212;
  assign n24214 = ~n24210 & ~n24213;
  assign n24215 = ~n24208 & n24214;
  assign n24216 = n24150 & ~n24215;
  assign n24217 = ~n24205 & ~n24216;
  assign n24218 = n24125 & n24139;
  assign n24219 = ~n24119 & n24218;
  assign n24220 = n24132 & n24164;
  assign n24221 = ~n24219 & ~n24220;
  assign n24222 = ~n24113 & ~n24221;
  assign n24223 = ~n24125 & ~n24138;
  assign n24224 = ~n24164 & ~n24223;
  assign n24225 = n24132 & ~n24224;
  assign n24226 = n24125 & n24132;
  assign n24227 = ~n24113 & n24226;
  assign n24228 = n24138 & n24227;
  assign n24229 = ~n24126 & ~n24189;
  assign n24230 = ~n24132 & ~n24229;
  assign n24231 = ~n24164 & ~n24230;
  assign n24232 = ~n24113 & ~n24231;
  assign n24233 = n24113 & ~n24132;
  assign n24234 = n24154 & n24233;
  assign n24235 = n24138 & n24234;
  assign n24236 = ~n24232 & ~n24235;
  assign n24237 = ~n24228 & n24236;
  assign n24238 = ~n24225 & n24237;
  assign n24239 = ~n24219 & n24238;
  assign n24240 = ~n24150 & ~n24239;
  assign n24241 = n24132 & n24189;
  assign n24242 = ~n24132 & n24180;
  assign n24243 = ~n24241 & ~n24242;
  assign n24244 = n24113 & ~n24243;
  assign n24245 = ~n24240 & ~n24244;
  assign n24246 = ~n24222 & n24245;
  assign n24247 = n24217 & n24246;
  assign n24248 = pi0316 & n24247;
  assign n24249 = ~pi0316 & ~n24247;
  assign po0338 = n24248 | n24249;
  assign n24251 = ~n23869 & n23913;
  assign n24252 = ~n23987 & ~n24251;
  assign n24253 = n23875 & ~n24252;
  assign n24254 = n23899 & n23910;
  assign n24255 = ~n24253 & ~n24254;
  assign n24256 = ~n23923 & n24255;
  assign n24257 = ~n23850 & ~n23875;
  assign n24258 = n23862 & n24257;
  assign n24259 = n23856 & n24258;
  assign n24260 = ~n23869 & n24259;
  assign n24261 = ~n23856 & n23869;
  assign n24262 = n23850 & n24261;
  assign n24263 = n23862 & n24262;
  assign n24264 = ~n23883 & ~n24263;
  assign n24265 = ~n23913 & n24264;
  assign n24266 = n23875 & ~n24265;
  assign n24267 = n23844 & n24266;
  assign n24268 = ~n23875 & n23996;
  assign n24269 = ~n23894 & ~n23921;
  assign n24270 = ~n23888 & n24269;
  assign n24271 = ~n24268 & n24270;
  assign n24272 = n23844 & ~n24271;
  assign n24273 = n23869 & n23931;
  assign n24274 = ~n24259 & ~n24273;
  assign n24275 = ~n23986 & n24274;
  assign n24276 = n23862 & n23892;
  assign n24277 = n23869 & n23880;
  assign n24278 = ~n23909 & ~n24277;
  assign n24279 = n23875 & ~n24278;
  assign n24280 = ~n24276 & ~n24279;
  assign n24281 = n24275 & n24280;
  assign n24282 = ~n23844 & ~n24281;
  assign n24283 = ~n24272 & ~n24282;
  assign n24284 = ~n24267 & n24283;
  assign n24285 = ~n24260 & n24284;
  assign n24286 = n24256 & n24285;
  assign n24287 = pi0311 & ~n24286;
  assign n24288 = ~pi0311 & n24256;
  assign n24289 = n24285 & n24288;
  assign po0339 = n24287 | n24289;
  assign n24291 = pi3131 & pi9040;
  assign n24292 = pi3143 & ~pi9040;
  assign n24293 = ~n24291 & ~n24292;
  assign n24294 = pi0257 & n24293;
  assign n24295 = ~pi0257 & ~n24293;
  assign n24296 = ~n24294 & ~n24295;
  assign n24297 = pi3146 & pi9040;
  assign n24298 = pi3135 & ~pi9040;
  assign n24299 = ~n24297 & ~n24298;
  assign n24300 = ~pi0261 & n24299;
  assign n24301 = pi0261 & ~n24299;
  assign n24302 = ~n24300 & ~n24301;
  assign n24303 = pi3159 & pi9040;
  assign n24304 = pi3144 & ~pi9040;
  assign n24305 = ~n24303 & ~n24304;
  assign n24306 = pi0274 & n24305;
  assign n24307 = ~pi0274 & ~n24305;
  assign n24308 = ~n24306 & ~n24307;
  assign n24309 = pi3161 & pi9040;
  assign n24310 = pi3131 & ~pi9040;
  assign n24311 = ~n24309 & ~n24310;
  assign n24312 = ~pi0280 & n24311;
  assign n24313 = pi0280 & ~n24311;
  assign n24314 = ~n24312 & ~n24313;
  assign n24315 = pi3144 & pi9040;
  assign n24316 = pi3170 & ~pi9040;
  assign n24317 = ~n24315 & ~n24316;
  assign n24318 = pi0276 & n24317;
  assign n24319 = ~pi0276 & ~n24317;
  assign n24320 = ~n24318 & ~n24319;
  assign n24321 = n24314 & n24320;
  assign n24322 = n24308 & n24321;
  assign n24323 = ~n24302 & n24322;
  assign n24324 = ~n24296 & n24323;
  assign n24325 = ~n24314 & ~n24320;
  assign n24326 = ~n24296 & ~n24302;
  assign n24327 = n24325 & n24326;
  assign n24328 = ~n24308 & n24327;
  assign n24329 = ~n24324 & ~n24328;
  assign n24330 = ~n24308 & n24321;
  assign n24331 = n24302 & n24330;
  assign n24332 = ~n24296 & n24331;
  assign n24333 = ~n24308 & n24325;
  assign n24334 = ~n24296 & n24333;
  assign n24335 = ~n24332 & ~n24334;
  assign n24336 = n24296 & ~n24314;
  assign n24337 = n24308 & n24336;
  assign n24338 = n24296 & n24321;
  assign n24339 = ~n24337 & ~n24338;
  assign n24340 = ~n24302 & ~n24339;
  assign n24341 = ~n24314 & n24320;
  assign n24342 = n24314 & ~n24320;
  assign n24343 = ~n24341 & ~n24342;
  assign n24344 = ~n24296 & ~n24308;
  assign n24345 = n24302 & ~n24344;
  assign n24346 = ~n24343 & n24345;
  assign n24347 = ~n24308 & ~n24321;
  assign n24348 = ~n24302 & n24347;
  assign n24349 = ~n24296 & n24348;
  assign n24350 = ~n24346 & ~n24349;
  assign n24351 = ~n24340 & n24350;
  assign n24352 = n24335 & n24351;
  assign n24353 = pi3217 & pi9040;
  assign n24354 = pi3138 & ~pi9040;
  assign n24355 = ~n24353 & ~n24354;
  assign n24356 = ~pi0251 & n24355;
  assign n24357 = pi0251 & ~n24355;
  assign n24358 = ~n24356 & ~n24357;
  assign n24359 = ~n24352 & ~n24358;
  assign n24360 = n24329 & ~n24359;
  assign n24361 = n24308 & n24341;
  assign n24362 = n24302 & n24361;
  assign n24363 = n24296 & n24362;
  assign n24364 = n24302 & n24358;
  assign n24365 = n24308 & n24325;
  assign n24366 = ~n24343 & n24344;
  assign n24367 = ~n24338 & ~n24366;
  assign n24368 = ~n24365 & n24367;
  assign n24369 = n24364 & ~n24368;
  assign n24370 = n24296 & n24333;
  assign n24371 = ~n24308 & n24336;
  assign n24372 = n24296 & n24342;
  assign n24373 = ~n24371 & ~n24372;
  assign n24374 = ~n24296 & n24321;
  assign n24375 = n24308 & n24342;
  assign n24376 = ~n24374 & ~n24375;
  assign n24377 = n24373 & n24376;
  assign n24378 = ~n24302 & ~n24377;
  assign n24379 = ~n24370 & ~n24378;
  assign n24380 = n24358 & ~n24379;
  assign n24381 = ~n24369 & ~n24380;
  assign n24382 = ~n24363 & n24381;
  assign n24383 = n24360 & n24382;
  assign n24384 = pi0298 & ~n24383;
  assign n24385 = ~pi0298 & n24360;
  assign n24386 = n24382 & n24385;
  assign po0341 = n24384 | n24386;
  assign n24388 = ~n24336 & ~n24375;
  assign n24389 = n24302 & ~n24358;
  assign n24390 = ~n24388 & n24389;
  assign n24391 = n24296 & n24308;
  assign n24392 = ~n24341 & n24391;
  assign n24393 = ~n24358 & n24392;
  assign n24394 = n24296 & ~n24308;
  assign n24395 = ~n24302 & n24394;
  assign n24396 = n24341 & n24395;
  assign n24397 = n24296 & n24302;
  assign n24398 = n24308 & n24397;
  assign n24399 = ~n24320 & n24398;
  assign n24400 = ~n24396 & ~n24399;
  assign n24401 = ~n24393 & n24400;
  assign n24402 = ~n24372 & ~n24374;
  assign n24403 = ~n24302 & ~n24402;
  assign n24404 = ~n24328 & ~n24403;
  assign n24405 = ~n24358 & ~n24404;
  assign n24406 = ~n24308 & ~n24314;
  assign n24407 = ~n24341 & ~n24406;
  assign n24408 = ~n24296 & ~n24407;
  assign n24409 = ~n24322 & ~n24408;
  assign n24410 = n24302 & ~n24409;
  assign n24411 = ~n24366 & ~n24410;
  assign n24412 = n24296 & n24330;
  assign n24413 = ~n24296 & n24308;
  assign n24414 = ~n24320 & n24413;
  assign n24415 = n24296 & ~n24407;
  assign n24416 = ~n24414 & ~n24415;
  assign n24417 = ~n24302 & ~n24416;
  assign n24418 = ~n24412 & ~n24417;
  assign n24419 = n24411 & n24418;
  assign n24420 = n24358 & ~n24419;
  assign n24421 = ~n24405 & ~n24420;
  assign n24422 = n24401 & n24421;
  assign n24423 = ~n24390 & n24422;
  assign n24424 = pi0319 & ~n24423;
  assign n24425 = ~pi0319 & n24401;
  assign n24426 = ~n24390 & n24425;
  assign n24427 = n24421 & n24426;
  assign po0342 = n24424 | n24427;
  assign n24429 = ~n24025 & ~n24086;
  assign n24430 = ~n24074 & n24429;
  assign n24431 = n23642 & ~n24430;
  assign n24432 = ~n24035 & ~n24052;
  assign n24433 = ~n24033 & ~n24082;
  assign n24434 = ~n24021 & ~n24089;
  assign n24435 = ~n23642 & ~n24434;
  assign n24436 = ~n23671 & ~n24435;
  assign n24437 = n24433 & n24436;
  assign n24438 = n23606 & ~n24437;
  assign n24439 = n23625 & n23631;
  assign n24440 = ~n23650 & ~n24439;
  assign n24441 = ~n23612 & ~n24440;
  assign n24442 = ~n23633 & ~n24038;
  assign n24443 = ~n23642 & ~n24442;
  assign n24444 = ~n23612 & n23631;
  assign n24445 = ~n23645 & ~n24444;
  assign n24446 = ~n23653 & n24445;
  assign n24447 = n23642 & ~n24446;
  assign n24448 = ~n24443 & ~n24447;
  assign n24449 = ~n24441 & n24448;
  assign n24450 = ~n23606 & ~n24449;
  assign n24451 = ~n24438 & ~n24450;
  assign n24452 = n24432 & n24451;
  assign n24453 = ~n24431 & n24452;
  assign n24454 = ~pi0320 & ~n24453;
  assign n24455 = pi0320 & n24432;
  assign n24456 = ~n24431 & n24455;
  assign n24457 = n24451 & n24456;
  assign po0343 = n24454 | n24457;
  assign n24459 = n23869 & ~n24008;
  assign n24460 = n23850 & n24459;
  assign n24461 = n23862 & n23985;
  assign n24462 = ~n23933 & ~n24461;
  assign n24463 = ~n23883 & n24462;
  assign n24464 = ~n23875 & ~n24463;
  assign n24465 = ~n23897 & ~n23996;
  assign n24466 = n23875 & ~n24465;
  assign n24467 = ~n24464 & ~n24466;
  assign n24468 = ~n24460 & n24467;
  assign n24469 = ~n23869 & n23910;
  assign n24470 = n24468 & ~n24469;
  assign n24471 = ~n23844 & ~n24470;
  assign n24472 = n23879 & ~n24465;
  assign n24473 = ~n23898 & ~n23913;
  assign n24474 = ~n23883 & ~n23910;
  assign n24475 = n24473 & n24474;
  assign n24476 = n23869 & ~n24475;
  assign n24477 = ~n24472 & ~n24476;
  assign n24478 = ~n23987 & n24477;
  assign n24479 = n23844 & ~n24478;
  assign n24480 = ~n24471 & ~n24479;
  assign n24481 = n23869 & n23996;
  assign n24482 = ~n24469 & ~n24481;
  assign n24483 = n23875 & ~n24482;
  assign n24484 = n24480 & ~n24483;
  assign n24485 = pi0321 & ~n24484;
  assign n24486 = ~pi0321 & ~n24483;
  assign n24487 = ~n24479 & n24486;
  assign n24488 = ~n24471 & n24487;
  assign po0344 = n24485 | n24488;
  assign n24490 = ~n23317 & n23323;
  assign n24491 = ~n23310 & n24490;
  assign n24492 = ~n23337 & n24491;
  assign n24493 = n23323 & n23352;
  assign n24494 = n23317 & ~n23329;
  assign n24495 = n23337 & n24494;
  assign n24496 = ~n23344 & ~n24495;
  assign n24497 = ~n24493 & n24496;
  assign n24498 = ~n24492 & n24497;
  assign n24499 = n23310 & n23340;
  assign n24500 = n24498 & ~n24499;
  assign n24501 = n23376 & ~n24500;
  assign n24502 = ~n23341 & ~n23344;
  assign n24503 = n23337 & n23393;
  assign n24504 = ~n23329 & ~n23337;
  assign n24505 = ~n23317 & n24504;
  assign n24506 = ~n24503 & ~n24505;
  assign n24507 = n24502 & n24506;
  assign n24508 = ~n23310 & ~n24507;
  assign n24509 = ~n24501 & ~n24508;
  assign n24510 = n23337 & n23346;
  assign n24511 = ~n23394 & ~n24510;
  assign n24512 = n23310 & ~n24511;
  assign n24513 = n23317 & n23337;
  assign n24514 = ~n23323 & n24513;
  assign n24515 = ~n24494 & ~n24514;
  assign n24516 = ~n23346 & n24515;
  assign n24517 = n23310 & ~n24516;
  assign n24518 = ~n23317 & n23363;
  assign n24519 = n23337 & n24518;
  assign n24520 = ~n24517 & ~n24519;
  assign n24521 = ~n23376 & ~n24520;
  assign n24522 = ~n23376 & n23378;
  assign n24523 = ~n23310 & n24522;
  assign n24524 = ~n24521 & ~n24523;
  assign n24525 = ~n24512 & n24524;
  assign n24526 = n24509 & n24525;
  assign n24527 = ~pi0305 & ~n24526;
  assign n24528 = pi0305 & n24509;
  assign n24529 = n24525 & n24528;
  assign po0345 = n24527 | n24529;
  assign n24531 = n23337 & n23367;
  assign n24532 = ~n23364 & ~n24505;
  assign n24533 = n23310 & ~n24532;
  assign n24534 = ~n24531 & ~n24533;
  assign n24535 = ~n23310 & n23337;
  assign n24536 = ~n23329 & n24535;
  assign n24537 = n23323 & n24536;
  assign n24538 = n23345 & n23379;
  assign n24539 = ~n24537 & ~n24538;
  assign n24540 = ~n23310 & n23317;
  assign n24541 = n23339 & n24540;
  assign n24542 = n24539 & ~n24541;
  assign n24543 = ~n23341 & ~n23353;
  assign n24544 = n23329 & n23343;
  assign n24545 = n24543 & ~n24544;
  assign n24546 = n24542 & n24545;
  assign n24547 = n24534 & n24546;
  assign n24548 = ~n23376 & ~n24547;
  assign n24549 = n23337 & n23363;
  assign n24550 = ~n24493 & ~n24549;
  assign n24551 = ~n23310 & ~n24550;
  assign n24552 = n23323 & n23382;
  assign n24553 = ~n23393 & ~n24552;
  assign n24554 = ~n23337 & n24494;
  assign n24555 = n24553 & ~n24554;
  assign n24556 = n23310 & ~n24555;
  assign n24557 = ~n23340 & ~n23364;
  assign n24558 = ~n23337 & ~n24557;
  assign n24559 = ~n24510 & ~n24558;
  assign n24560 = ~n24556 & n24559;
  assign n24561 = ~n24551 & n24560;
  assign n24562 = n23376 & ~n24561;
  assign n24563 = n23310 & n23383;
  assign n24564 = ~n24562 & ~n24563;
  assign n24565 = n23358 & n24535;
  assign n24566 = ~n23329 & n24565;
  assign n24567 = n24564 & ~n24566;
  assign n24568 = ~n24548 & n24567;
  assign n24569 = ~pi0308 & ~n24568;
  assign n24570 = pi0308 & n24564;
  assign n24571 = ~n24548 & n24570;
  assign n24572 = ~n24566 & n24571;
  assign po0346 = n24569 | n24572;
  assign n24574 = ~n24125 & n24141;
  assign n24575 = ~n24172 & ~n24574;
  assign n24576 = ~n24113 & ~n24575;
  assign n24577 = ~n24132 & n24163;
  assign n24578 = ~n24212 & ~n24577;
  assign n24579 = n24113 & ~n24578;
  assign n24580 = n24132 & n24158;
  assign n24581 = ~n24228 & ~n24580;
  assign n24582 = ~n24140 & n24581;
  assign n24583 = ~n24579 & n24582;
  assign n24584 = ~n24576 & n24583;
  assign n24585 = ~n24208 & ~n24219;
  assign n24586 = n24584 & n24585;
  assign n24587 = n24150 & ~n24586;
  assign n24588 = n24126 & n24206;
  assign n24589 = n24181 & ~n24588;
  assign n24590 = n24113 & ~n24589;
  assign n24591 = n24132 & n24169;
  assign n24592 = ~n24590 & ~n24591;
  assign n24593 = n24119 & n24141;
  assign n24594 = ~n24132 & n24154;
  assign n24595 = ~n24593 & ~n24594;
  assign n24596 = n24113 & ~n24595;
  assign n24597 = n24113 & n24163;
  assign n24598 = n24132 & n24597;
  assign n24599 = ~n24596 & ~n24598;
  assign n24600 = n24592 & n24599;
  assign n24601 = ~n24150 & ~n24600;
  assign n24602 = ~n24158 & ~n24165;
  assign n24603 = ~n24213 & n24602;
  assign n24604 = n24186 & ~n24603;
  assign n24605 = ~n24601 & ~n24604;
  assign n24606 = ~n24140 & ~n24208;
  assign n24607 = ~n24113 & ~n24606;
  assign n24608 = n24605 & ~n24607;
  assign n24609 = ~n24587 & n24608;
  assign n24610 = ~pi0303 & n24609;
  assign n24611 = pi0303 & ~n24609;
  assign po0347 = n24610 | n24611;
  assign n24613 = ~n23338 & ~n23344;
  assign n24614 = ~n23310 & ~n24613;
  assign n24615 = ~n23400 & ~n24614;
  assign n24616 = ~n23317 & ~n23323;
  assign n24617 = n23310 & n24616;
  assign n24618 = ~n23337 & n24617;
  assign n24619 = ~n23310 & n23330;
  assign n24620 = ~n23337 & n24619;
  assign n24621 = ~n24541 & ~n24620;
  assign n24622 = n23323 & n24513;
  assign n24623 = ~n23337 & n23363;
  assign n24624 = ~n24622 & ~n24623;
  assign n24625 = ~n24616 & n24624;
  assign n24626 = n23310 & ~n24625;
  assign n24627 = ~n23347 & ~n24626;
  assign n24628 = n24621 & n24627;
  assign n24629 = ~n23376 & ~n24628;
  assign n24630 = ~n24618 & ~n24629;
  assign n24631 = ~n23364 & ~n23383;
  assign n24632 = ~n23393 & n24631;
  assign n24633 = ~n23310 & ~n24632;
  assign n24634 = n23337 & n23388;
  assign n24635 = ~n23367 & ~n24634;
  assign n24636 = n23310 & ~n24635;
  assign n24637 = ~n24552 & ~n24636;
  assign n24638 = ~n24633 & n24637;
  assign n24639 = ~n23353 & ~n23394;
  assign n24640 = n24638 & n24639;
  assign n24641 = n23376 & ~n24640;
  assign n24642 = n24630 & ~n24641;
  assign n24643 = n24615 & n24642;
  assign n24644 = ~pi0317 & ~n24643;
  assign n24645 = pi0317 & n24630;
  assign n24646 = n24615 & n24645;
  assign n24647 = ~n24641 & n24646;
  assign po0348 = n24644 | n24647;
  assign n24649 = ~n24333 & ~n24361;
  assign n24650 = n24320 & n24413;
  assign n24651 = n24649 & ~n24650;
  assign n24652 = n24389 & ~n24651;
  assign n24653 = ~n24358 & n24375;
  assign n24654 = n24296 & n24653;
  assign n24655 = ~n24302 & n24365;
  assign n24656 = ~n24308 & n24320;
  assign n24657 = ~n24338 & ~n24656;
  assign n24658 = ~n24302 & ~n24657;
  assign n24659 = ~n24655 & ~n24658;
  assign n24660 = ~n24358 & ~n24659;
  assign n24661 = ~n24654 & ~n24660;
  assign n24662 = n24320 & n24394;
  assign n24663 = ~n24320 & n24344;
  assign n24664 = n24314 & n24663;
  assign n24665 = ~n24662 & ~n24664;
  assign n24666 = ~n24302 & ~n24665;
  assign n24667 = n24661 & ~n24666;
  assign n24668 = n24321 & n24397;
  assign n24669 = n24308 & n24668;
  assign n24670 = ~n24343 & n24413;
  assign n24671 = ~n24334 & ~n24670;
  assign n24672 = ~n24343 & n24394;
  assign n24673 = n24296 & n24365;
  assign n24674 = ~n24672 & ~n24673;
  assign n24675 = ~n24332 & n24674;
  assign n24676 = n24671 & n24675;
  assign n24677 = ~n24669 & n24676;
  assign n24678 = n24308 & n24326;
  assign n24679 = n24314 & n24678;
  assign n24680 = n24677 & ~n24679;
  assign n24681 = n24358 & ~n24680;
  assign n24682 = n24667 & ~n24681;
  assign n24683 = ~n24652 & n24682;
  assign n24684 = ~pi0313 & ~n24683;
  assign n24685 = pi0313 & n24667;
  assign n24686 = ~n24652 & n24685;
  assign n24687 = ~n24681 & n24686;
  assign po0349 = n24684 | n24687;
  assign n24689 = ~n23760 & n23781;
  assign n24690 = ~n23961 & ~n24689;
  assign n24691 = ~n23766 & n24690;
  assign n24692 = n23760 & n23824;
  assign n24693 = ~n23754 & ~n23775;
  assign n24694 = n23774 & ~n24693;
  assign n24695 = ~n23747 & n23800;
  assign n24696 = n23760 & n23775;
  assign n24697 = ~n24695 & ~n24696;
  assign n24698 = n23766 & n24697;
  assign n24699 = ~n24694 & n24698;
  assign n24700 = ~n24692 & n24699;
  assign n24701 = ~n24691 & ~n24700;
  assign n24702 = n23760 & n24694;
  assign n24703 = ~n23959 & ~n24702;
  assign n24704 = ~n24701 & n24703;
  assign n24705 = n23741 & ~n24704;
  assign n24706 = ~n23766 & ~n24693;
  assign n24707 = ~n23760 & n24706;
  assign n24708 = n23760 & n23818;
  assign n24709 = ~n23796 & ~n24708;
  assign n24710 = ~n23766 & ~n24709;
  assign n24711 = ~n23774 & n24706;
  assign n24712 = ~n24710 & ~n24711;
  assign n24713 = ~n24707 & n24712;
  assign n24714 = ~n23741 & ~n24713;
  assign n24715 = ~n24705 & ~n24714;
  assign n24716 = n23766 & ~n24690;
  assign n24717 = ~n23779 & ~n24716;
  assign n24718 = ~n23741 & ~n24717;
  assign n24719 = ~n23766 & n23779;
  assign n24720 = n23766 & ~n24703;
  assign n24721 = ~n24719 & ~n24720;
  assign n24722 = ~n24718 & n24721;
  assign n24723 = n24715 & n24722;
  assign n24724 = pi0314 & ~n24723;
  assign n24725 = ~pi0314 & n24722;
  assign n24726 = ~n24714 & n24725;
  assign n24727 = ~n24705 & n24726;
  assign po0350 = n24724 | n24727;
  assign n24729 = ~n24308 & n24372;
  assign n24730 = ~n24673 & ~n24729;
  assign n24731 = ~n24302 & ~n24730;
  assign n24732 = ~n24308 & n24341;
  assign n24733 = ~n24322 & ~n24732;
  assign n24734 = ~n24302 & ~n24733;
  assign n24735 = ~n24296 & n24342;
  assign n24736 = ~n24361 & ~n24735;
  assign n24737 = ~n24330 & n24736;
  assign n24738 = n24302 & ~n24737;
  assign n24739 = ~n24734 & ~n24738;
  assign n24740 = ~n24655 & ~n24664;
  assign n24741 = n24739 & n24740;
  assign n24742 = n24358 & ~n24741;
  assign n24743 = n24296 & n24322;
  assign n24744 = ~n24296 & n24325;
  assign n24745 = ~n24372 & ~n24744;
  assign n24746 = n24302 & ~n24745;
  assign n24747 = ~n24743 & ~n24746;
  assign n24748 = ~n24302 & n24308;
  assign n24749 = ~n24320 & n24748;
  assign n24750 = n24314 & n24749;
  assign n24751 = n24649 & ~n24750;
  assign n24752 = ~n24330 & n24751;
  assign n24753 = ~n24296 & ~n24752;
  assign n24754 = n24747 & ~n24753;
  assign n24755 = ~n24358 & ~n24754;
  assign n24756 = ~n24742 & ~n24755;
  assign n24757 = n24397 & n24406;
  assign n24758 = n24756 & ~n24757;
  assign n24759 = ~n24731 & n24758;
  assign n24760 = ~pi0304 & ~n24759;
  assign n24761 = pi0304 & ~n24731;
  assign n24762 = n24756 & n24761;
  assign n24763 = ~n24757 & n24762;
  assign po0351 = n24760 | n24763;
  assign n24765 = ~n24113 & n24169;
  assign n24766 = n24132 & n24154;
  assign n24767 = ~n24153 & ~n24766;
  assign n24768 = ~n24113 & ~n24767;
  assign n24769 = n24113 & ~n24224;
  assign n24770 = ~n24768 & ~n24769;
  assign n24771 = ~n24242 & n24770;
  assign n24772 = n24150 & ~n24771;
  assign n24773 = ~n24765 & ~n24772;
  assign n24774 = ~n24138 & n24199;
  assign n24775 = ~n24211 & ~n24774;
  assign n24776 = ~n24119 & ~n24775;
  assign n24777 = ~n24140 & ~n24776;
  assign n24778 = ~n24212 & n24777;
  assign n24779 = ~n24132 & n24172;
  assign n24780 = n24113 & n24155;
  assign n24781 = ~n24779 & ~n24780;
  assign n24782 = n24778 & n24781;
  assign n24783 = ~n24150 & ~n24782;
  assign n24784 = ~n24580 & ~n24594;
  assign n24785 = n24113 & ~n24784;
  assign n24786 = ~n24783 & ~n24785;
  assign n24787 = n24773 & n24786;
  assign n24788 = ~pi0340 & ~n24787;
  assign n24789 = ~n24772 & n24786;
  assign n24790 = pi0340 & n24789;
  assign n24791 = ~n24765 & n24790;
  assign po0352 = n24788 | n24791;
  assign n24793 = ~n23766 & n23806;
  assign n24794 = n23800 & ~n24693;
  assign n24795 = ~n23819 & ~n24794;
  assign n24796 = ~n23959 & n24795;
  assign n24797 = n23766 & ~n24796;
  assign n24798 = n23760 & n23776;
  assign n24799 = ~n24797 & ~n24798;
  assign n24800 = ~n23774 & n23818;
  assign n24801 = ~n23760 & n23966;
  assign n24802 = ~n24800 & ~n24801;
  assign n24803 = ~n24696 & n24802;
  assign n24804 = ~n23766 & ~n24803;
  assign n24805 = n24799 & ~n24804;
  assign n24806 = n23741 & ~n24805;
  assign n24807 = ~n24793 & ~n24806;
  assign n24808 = ~n23760 & n23775;
  assign n24809 = ~n23958 & ~n24808;
  assign n24810 = ~n23766 & ~n24809;
  assign n24811 = ~n23820 & ~n24810;
  assign n24812 = ~n23796 & ~n23806;
  assign n24813 = n23760 & n23777;
  assign n24814 = ~n23966 & ~n24813;
  assign n24815 = ~n24800 & n24814;
  assign n24816 = n23766 & ~n24815;
  assign n24817 = ~n23760 & n23776;
  assign n24818 = ~n24816 & ~n24817;
  assign n24819 = n24812 & n24818;
  assign n24820 = n24811 & n24819;
  assign n24821 = ~n23741 & ~n24820;
  assign n24822 = ~n23812 & ~n24692;
  assign n24823 = n23766 & ~n24822;
  assign n24824 = ~n24821 & ~n24823;
  assign n24825 = n24807 & n24824;
  assign n24826 = pi0318 & n24825;
  assign n24827 = ~pi0318 & ~n24825;
  assign po0353 = n24826 | n24827;
  assign n24829 = pi3232 & pi9040;
  assign n24830 = pi3322 & ~pi9040;
  assign n24831 = ~n24829 & ~n24830;
  assign n24832 = pi0335 & n24831;
  assign n24833 = ~pi0335 & ~n24831;
  assign n24834 = ~n24832 & ~n24833;
  assign n24835 = pi3199 & pi9040;
  assign n24836 = pi3255 & ~pi9040;
  assign n24837 = ~n24835 & ~n24836;
  assign n24838 = pi0341 & n24837;
  assign n24839 = ~pi0341 & ~n24837;
  assign n24840 = ~n24838 & ~n24839;
  assign n24841 = pi3230 & pi9040;
  assign n24842 = pi3250 & ~pi9040;
  assign n24843 = ~n24841 & ~n24842;
  assign n24844 = ~pi0312 & n24843;
  assign n24845 = pi0312 & ~n24843;
  assign n24846 = ~n24844 & ~n24845;
  assign n24847 = pi3208 & pi9040;
  assign n24848 = pi3201 & ~pi9040;
  assign n24849 = ~n24847 & ~n24848;
  assign n24850 = pi0334 & n24849;
  assign n24851 = ~pi0334 & ~n24849;
  assign n24852 = ~n24850 & ~n24851;
  assign n24853 = pi3211 & pi9040;
  assign n24854 = pi3333 & ~pi9040;
  assign n24855 = ~n24853 & ~n24854;
  assign n24856 = pi0345 & n24855;
  assign n24857 = ~pi0345 & ~n24855;
  assign n24858 = ~n24856 & ~n24857;
  assign n24859 = ~n24852 & ~n24858;
  assign n24860 = ~n24846 & n24859;
  assign n24861 = ~n24840 & n24860;
  assign n24862 = pi3295 & pi9040;
  assign n24863 = pi3232 & ~pi9040;
  assign n24864 = ~n24862 & ~n24863;
  assign n24865 = ~pi0336 & ~n24864;
  assign n24866 = pi0336 & n24864;
  assign n24867 = ~n24865 & ~n24866;
  assign n24868 = n24840 & n24846;
  assign n24869 = n24867 & n24868;
  assign n24870 = n24852 & ~n24867;
  assign n24871 = n24846 & n24870;
  assign n24872 = ~n24840 & n24871;
  assign n24873 = ~n24869 & ~n24872;
  assign n24874 = n24840 & ~n24846;
  assign n24875 = n24852 & n24874;
  assign n24876 = n24873 & ~n24875;
  assign n24877 = ~n24858 & ~n24876;
  assign n24878 = n24840 & ~n24867;
  assign n24879 = ~n24852 & n24858;
  assign n24880 = n24878 & n24879;
  assign n24881 = ~n24867 & n24868;
  assign n24882 = ~n24852 & n24881;
  assign n24883 = ~n24880 & ~n24882;
  assign n24884 = ~n24877 & n24883;
  assign n24885 = ~n24861 & n24884;
  assign n24886 = ~n24840 & ~n24846;
  assign n24887 = n24867 & n24886;
  assign n24888 = ~n24852 & n24887;
  assign n24889 = n24852 & n24867;
  assign n24890 = ~n24846 & n24889;
  assign n24891 = n24840 & n24890;
  assign n24892 = ~n24888 & ~n24891;
  assign n24893 = n24885 & n24892;
  assign n24894 = ~n24834 & ~n24893;
  assign n24895 = ~n24867 & n24874;
  assign n24896 = ~n24852 & n24895;
  assign n24897 = ~n24887 & ~n24896;
  assign n24898 = ~n24858 & ~n24897;
  assign n24899 = ~n24867 & n24886;
  assign n24900 = n24852 & n24899;
  assign n24901 = ~n24852 & ~n24867;
  assign n24902 = n24846 & n24901;
  assign n24903 = ~n24840 & n24902;
  assign n24904 = ~n24900 & ~n24903;
  assign n24905 = n24840 & n24870;
  assign n24906 = ~n24852 & n24867;
  assign n24907 = ~n24846 & n24906;
  assign n24908 = n24840 & n24907;
  assign n24909 = ~n24905 & ~n24908;
  assign n24910 = n24858 & ~n24909;
  assign n24911 = n24904 & ~n24910;
  assign n24912 = ~n24898 & n24911;
  assign n24913 = n24834 & ~n24912;
  assign n24914 = ~n24840 & n24846;
  assign n24915 = n24867 & n24914;
  assign n24916 = n24852 & n24915;
  assign n24917 = ~n24881 & ~n24916;
  assign n24918 = ~n24900 & n24917;
  assign n24919 = n24858 & ~n24918;
  assign n24920 = ~n24840 & n24867;
  assign n24921 = ~n24852 & n24920;
  assign n24922 = n24840 & n24867;
  assign n24923 = n24852 & n24922;
  assign n24924 = ~n24921 & ~n24923;
  assign n24925 = ~n24858 & ~n24924;
  assign n24926 = ~n24919 & ~n24925;
  assign n24927 = n24846 & ~n24867;
  assign n24928 = n24858 & n24927;
  assign n24929 = ~n24852 & n24928;
  assign n24930 = n24926 & ~n24929;
  assign n24931 = ~n24913 & n24930;
  assign n24932 = ~n24894 & n24931;
  assign n24933 = ~pi0359 & ~n24932;
  assign n24934 = pi0359 & n24932;
  assign po0375 = n24933 | n24934;
  assign n24936 = pi3213 & pi9040;
  assign n24937 = pi3295 & ~pi9040;
  assign n24938 = ~n24936 & ~n24937;
  assign n24939 = pi0325 & n24938;
  assign n24940 = ~pi0325 & ~n24938;
  assign n24941 = ~n24939 & ~n24940;
  assign n24942 = pi3345 & pi9040;
  assign n24943 = pi3252 & ~pi9040;
  assign n24944 = ~n24942 & ~n24943;
  assign n24945 = ~pi0312 & n24944;
  assign n24946 = pi0312 & ~n24944;
  assign n24947 = ~n24945 & ~n24946;
  assign n24948 = pi3218 & pi9040;
  assign n24949 = pi3282 & ~pi9040;
  assign n24950 = ~n24948 & ~n24949;
  assign n24951 = pi0342 & n24950;
  assign n24952 = ~pi0342 & ~n24950;
  assign n24953 = ~n24951 & ~n24952;
  assign n24954 = pi3215 & pi9040;
  assign n24955 = pi3214 & ~pi9040;
  assign n24956 = ~n24954 & ~n24955;
  assign n24957 = ~pi0335 & n24956;
  assign n24958 = pi0335 & ~n24956;
  assign n24959 = ~n24957 & ~n24958;
  assign n24960 = n24953 & ~n24959;
  assign n24961 = n24947 & n24960;
  assign n24962 = pi3258 & pi9040;
  assign n24963 = pi3219 & ~pi9040;
  assign n24964 = ~n24962 & ~n24963;
  assign n24965 = pi0347 & n24964;
  assign n24966 = ~pi0347 & ~n24964;
  assign n24967 = ~n24965 & ~n24966;
  assign n24968 = n24961 & ~n24967;
  assign n24969 = pi0335 & n24956;
  assign n24970 = ~pi0335 & ~n24956;
  assign n24971 = ~n24969 & ~n24970;
  assign n24972 = ~n24953 & ~n24971;
  assign n24973 = n24947 & n24972;
  assign n24974 = ~n24967 & n24973;
  assign n24975 = ~n24968 & ~n24974;
  assign n24976 = ~n24947 & n24967;
  assign n24977 = n24972 & n24976;
  assign n24978 = n24953 & ~n24971;
  assign n24979 = n24947 & n24978;
  assign n24980 = n24967 & n24979;
  assign n24981 = ~n24977 & ~n24980;
  assign n24982 = n24975 & n24981;
  assign n24983 = n24941 & ~n24982;
  assign n24984 = n24947 & n24967;
  assign n24985 = ~n24959 & n24984;
  assign n24986 = ~n24953 & n24985;
  assign n24987 = ~n24979 & ~n24986;
  assign n24988 = n24941 & ~n24987;
  assign n24989 = ~n24959 & ~n24967;
  assign n24990 = ~n24941 & n24989;
  assign n24991 = ~n24947 & n24953;
  assign n24992 = n24967 & n24972;
  assign n24993 = ~n24991 & ~n24992;
  assign n24994 = ~n24941 & ~n24993;
  assign n24995 = ~n24990 & ~n24994;
  assign n24996 = ~n24953 & ~n24959;
  assign n24997 = ~n24947 & n24996;
  assign n24998 = ~n24967 & n24997;
  assign n24999 = n24995 & ~n24998;
  assign n25000 = ~n24959 & n24991;
  assign n25001 = n24967 & n25000;
  assign n25002 = n24999 & ~n25001;
  assign n25003 = ~n24988 & n25002;
  assign n25004 = pi3255 & pi9040;
  assign n25005 = pi3345 & ~pi9040;
  assign n25006 = ~n25004 & ~n25005;
  assign n25007 = ~pi0350 & ~n25006;
  assign n25008 = pi0350 & n25006;
  assign n25009 = ~n25007 & ~n25008;
  assign n25010 = ~n25003 & ~n25009;
  assign n25011 = n24947 & ~n24959;
  assign n25012 = ~n24941 & n24967;
  assign n25013 = n25009 & n25012;
  assign n25014 = n25011 & n25013;
  assign n25015 = n24947 & ~n24967;
  assign n25016 = ~n24971 & n25015;
  assign n25017 = ~n24941 & ~n25016;
  assign n25018 = ~n24960 & ~n25011;
  assign n25019 = ~n24967 & ~n25018;
  assign n25020 = ~n24953 & n24976;
  assign n25021 = ~n24947 & n24972;
  assign n25022 = ~n25020 & ~n25021;
  assign n25023 = ~n25019 & n25022;
  assign n25024 = n24941 & n25023;
  assign n25025 = ~n25017 & ~n25024;
  assign n25026 = ~n24947 & n24978;
  assign n25027 = n24967 & n25026;
  assign n25028 = ~n25025 & ~n25027;
  assign n25029 = n25009 & ~n25028;
  assign n25030 = ~n25014 & ~n25029;
  assign n25031 = ~n25010 & n25030;
  assign n25032 = ~n24983 & n25031;
  assign n25033 = ~n24941 & n24998;
  assign n25034 = n25032 & ~n25033;
  assign n25035 = pi0352 & ~n25034;
  assign n25036 = ~pi0352 & ~n25033;
  assign n25037 = n25031 & n25036;
  assign n25038 = ~n24983 & n25037;
  assign po0380 = n25035 | n25038;
  assign n25040 = n24852 & n24881;
  assign n25041 = ~n24896 & ~n25040;
  assign n25042 = ~n24903 & ~n24922;
  assign n25043 = n24858 & ~n25042;
  assign n25044 = n25041 & ~n25043;
  assign n25045 = n24852 & ~n24858;
  assign n25046 = n24899 & n25045;
  assign n25047 = ~n24888 & ~n25046;
  assign n25048 = ~n24916 & n25047;
  assign n25049 = n25044 & n25048;
  assign n25050 = n24834 & ~n25049;
  assign n25051 = n24852 & n24895;
  assign n25052 = ~n24872 & ~n25051;
  assign n25053 = ~n24852 & n24915;
  assign n25054 = ~n24882 & ~n25053;
  assign n25055 = n24858 & n24899;
  assign n25056 = n24852 & n24887;
  assign n25057 = ~n25055 & ~n25056;
  assign n25058 = ~n24846 & n24867;
  assign n25059 = n24840 & n24852;
  assign n25060 = ~n25058 & ~n25059;
  assign n25061 = ~n24927 & n25060;
  assign n25062 = ~n24858 & ~n25061;
  assign n25063 = n25057 & ~n25062;
  assign n25064 = n25054 & n25063;
  assign n25065 = n25052 & n25064;
  assign n25066 = ~n24834 & ~n25065;
  assign n25067 = ~n25050 & ~n25066;
  assign n25068 = pi0355 & ~n25067;
  assign n25069 = ~pi0355 & ~n25050;
  assign n25070 = ~n25066 & n25069;
  assign po0381 = n25068 | n25070;
  assign n25072 = pi3307 & ~pi9040;
  assign n25073 = pi3229 & pi9040;
  assign n25074 = ~n25072 & ~n25073;
  assign n25075 = ~pi0329 & ~n25074;
  assign n25076 = pi0329 & n25074;
  assign n25077 = ~n25075 & ~n25076;
  assign n25078 = pi3222 & pi9040;
  assign n25079 = pi3207 & ~pi9040;
  assign n25080 = ~n25078 & ~n25079;
  assign n25081 = ~pi0342 & n25080;
  assign n25082 = pi0342 & ~n25080;
  assign n25083 = ~n25081 & ~n25082;
  assign n25084 = pi3307 & pi9040;
  assign n25085 = pi3234 & ~pi9040;
  assign n25086 = ~n25084 & ~n25085;
  assign n25087 = ~pi0350 & n25086;
  assign n25088 = pi0350 & ~n25086;
  assign n25089 = ~n25087 & ~n25088;
  assign n25090 = pi3226 & pi9040;
  assign n25091 = pi3257 & ~pi9040;
  assign n25092 = ~n25090 & ~n25091;
  assign n25093 = ~pi0302 & n25092;
  assign n25094 = pi0302 & ~n25092;
  assign n25095 = ~n25093 & ~n25094;
  assign n25096 = n25089 & ~n25095;
  assign n25097 = pi3212 & pi9040;
  assign n25098 = pi3298 & ~pi9040;
  assign n25099 = ~n25097 & ~n25098;
  assign n25100 = pi0343 & n25099;
  assign n25101 = ~pi0343 & ~n25099;
  assign n25102 = ~n25100 & ~n25101;
  assign n25103 = pi3298 & pi9040;
  assign n25104 = pi3239 & ~pi9040;
  assign n25105 = ~n25103 & ~n25104;
  assign n25106 = ~pi0348 & n25105;
  assign n25107 = pi0348 & ~n25105;
  assign n25108 = ~n25106 & ~n25107;
  assign n25109 = n25102 & ~n25108;
  assign n25110 = n25096 & n25109;
  assign n25111 = ~n25083 & n25110;
  assign n25112 = ~n25102 & ~n25108;
  assign n25113 = ~n25089 & ~n25095;
  assign n25114 = n25112 & n25113;
  assign n25115 = n25089 & n25095;
  assign n25116 = ~n25083 & n25115;
  assign n25117 = ~n25102 & n25116;
  assign n25118 = ~n25089 & n25095;
  assign n25119 = ~n25083 & n25118;
  assign n25120 = ~n25108 & n25119;
  assign n25121 = n25102 & n25120;
  assign n25122 = ~n25117 & ~n25121;
  assign n25123 = ~n25114 & n25122;
  assign n25124 = ~n25111 & n25123;
  assign n25125 = n25083 & ~n25102;
  assign n25126 = ~n25095 & n25125;
  assign n25127 = ~n25089 & n25126;
  assign n25128 = n25124 & ~n25127;
  assign n25129 = ~n25077 & ~n25128;
  assign n25130 = n25083 & n25095;
  assign n25131 = ~n25089 & n25130;
  assign n25132 = n25102 & n25108;
  assign n25133 = n25131 & n25132;
  assign n25134 = ~n25083 & ~n25102;
  assign n25135 = n25089 & n25134;
  assign n25136 = ~n25102 & n25115;
  assign n25137 = ~n25135 & ~n25136;
  assign n25138 = n25108 & ~n25137;
  assign n25139 = ~n25133 & ~n25138;
  assign n25140 = ~n25077 & ~n25139;
  assign n25141 = n25095 & n25134;
  assign n25142 = ~n25083 & ~n25089;
  assign n25143 = ~n25095 & n25142;
  assign n25144 = n25102 & n25143;
  assign n25145 = ~n25141 & ~n25144;
  assign n25146 = n25083 & n25096;
  assign n25147 = n25102 & n25146;
  assign n25148 = n25145 & ~n25147;
  assign n25149 = n25108 & ~n25148;
  assign n25150 = ~n25140 & ~n25149;
  assign n25151 = ~n25129 & n25150;
  assign n25152 = n25083 & n25102;
  assign n25153 = ~n25108 & n25152;
  assign n25154 = n25115 & n25153;
  assign n25155 = n25083 & ~n25089;
  assign n25156 = n25112 & n25155;
  assign n25157 = n25108 & n25142;
  assign n25158 = n25089 & n25102;
  assign n25159 = n25083 & n25158;
  assign n25160 = ~n25146 & ~n25159;
  assign n25161 = ~n25157 & n25160;
  assign n25162 = ~n25102 & n25131;
  assign n25163 = n25161 & ~n25162;
  assign n25164 = n25096 & ~n25108;
  assign n25165 = ~n25102 & n25164;
  assign n25166 = n25083 & ~n25095;
  assign n25167 = n25102 & n25115;
  assign n25168 = ~n25166 & ~n25167;
  assign n25169 = ~n25108 & ~n25168;
  assign n25170 = ~n25165 & ~n25169;
  assign n25171 = n25163 & n25170;
  assign n25172 = n25077 & ~n25171;
  assign n25173 = ~n25156 & ~n25172;
  assign n25174 = ~n25154 & n25173;
  assign n25175 = n25151 & n25174;
  assign n25176 = pi0373 & n25175;
  assign n25177 = ~pi0373 & ~n25175;
  assign po0384 = n25176 | n25177;
  assign n25179 = ~n25083 & n25089;
  assign n25180 = ~n25127 & ~n25179;
  assign n25181 = ~n25158 & n25180;
  assign n25182 = ~n25108 & ~n25181;
  assign n25183 = ~n25089 & n25132;
  assign n25184 = ~n25083 & n25102;
  assign n25185 = ~n25095 & n25184;
  assign n25186 = ~n25102 & n25119;
  assign n25187 = ~n25185 & ~n25186;
  assign n25188 = n25083 & n25089;
  assign n25189 = ~n25102 & n25108;
  assign n25190 = n25188 & n25189;
  assign n25191 = n25187 & ~n25190;
  assign n25192 = ~n25183 & n25191;
  assign n25193 = ~n25182 & n25192;
  assign n25194 = n25077 & ~n25193;
  assign n25195 = ~n25083 & n25096;
  assign n25196 = ~n25102 & n25195;
  assign n25197 = n25102 & n25116;
  assign n25198 = ~n25196 & ~n25197;
  assign n25199 = ~n25108 & ~n25198;
  assign n25200 = ~n25194 & ~n25199;
  assign n25201 = n25102 & n25119;
  assign n25202 = ~n25131 & ~n25143;
  assign n25203 = ~n25108 & ~n25202;
  assign n25204 = ~n25201 & ~n25203;
  assign n25205 = ~n25147 & n25204;
  assign n25206 = ~n25077 & ~n25205;
  assign n25207 = ~n25113 & ~n25115;
  assign n25208 = n25083 & ~n25207;
  assign n25209 = ~n25136 & ~n25208;
  assign n25210 = n25108 & ~n25209;
  assign n25211 = ~n25077 & n25210;
  assign n25212 = ~n25206 & ~n25211;
  assign n25213 = n25200 & n25212;
  assign n25214 = pi0374 & ~n25213;
  assign n25215 = ~pi0374 & n25200;
  assign n25216 = n25212 & n25215;
  assign po0385 = n25214 | n25216;
  assign n25218 = pi3292 & pi9040;
  assign n25219 = pi3226 & ~pi9040;
  assign n25220 = ~n25218 & ~n25219;
  assign n25221 = ~pi0332 & n25220;
  assign n25222 = pi0332 & ~n25220;
  assign n25223 = ~n25221 & ~n25222;
  assign n25224 = pi3234 & pi9040;
  assign n25225 = pi3263 & ~pi9040;
  assign n25226 = ~n25224 & ~n25225;
  assign n25227 = pi0331 & n25226;
  assign n25228 = ~pi0331 & ~n25226;
  assign n25229 = ~n25227 & ~n25228;
  assign n25230 = pi3200 & pi9040;
  assign n25231 = pi3292 & ~pi9040;
  assign n25232 = ~n25230 & ~n25231;
  assign n25233 = ~pi0344 & n25232;
  assign n25234 = pi0344 & ~n25232;
  assign n25235 = ~n25233 & ~n25234;
  assign n25236 = pi3294 & pi9040;
  assign n25237 = pi3229 & ~pi9040;
  assign n25238 = ~n25236 & ~n25237;
  assign n25239 = ~pi0323 & ~n25238;
  assign n25240 = pi0323 & n25238;
  assign n25241 = ~n25239 & ~n25240;
  assign n25242 = pi3207 & pi9040;
  assign n25243 = pi3206 & ~pi9040;
  assign n25244 = ~n25242 & ~n25243;
  assign n25245 = ~pi0328 & n25244;
  assign n25246 = pi0328 & ~n25244;
  assign n25247 = ~n25245 & ~n25246;
  assign n25248 = ~n25241 & n25247;
  assign n25249 = n25235 & n25248;
  assign n25250 = ~n25229 & n25249;
  assign n25251 = n25229 & n25235;
  assign n25252 = n25247 & n25251;
  assign n25253 = n25241 & n25252;
  assign n25254 = ~n25250 & ~n25253;
  assign n25255 = ~n25223 & ~n25254;
  assign n25256 = ~n25241 & ~n25247;
  assign n25257 = ~n25235 & n25256;
  assign n25258 = ~n25229 & n25257;
  assign n25259 = n25223 & n25258;
  assign n25260 = pi3202 & pi9040;
  assign n25261 = pi3210 & ~pi9040;
  assign n25262 = ~n25260 & ~n25261;
  assign n25263 = ~pi0346 & ~n25262;
  assign n25264 = pi0346 & ~n25260;
  assign n25265 = ~n25261 & n25264;
  assign n25266 = ~n25263 & ~n25265;
  assign n25267 = n25241 & n25247;
  assign n25268 = ~n25235 & n25267;
  assign n25269 = ~n25223 & n25268;
  assign n25270 = ~n25258 & ~n25269;
  assign n25271 = ~n25229 & n25241;
  assign n25272 = n25235 & n25271;
  assign n25273 = ~n25229 & ~n25235;
  assign n25274 = ~n25241 & n25273;
  assign n25275 = ~n25272 & ~n25274;
  assign n25276 = n25223 & ~n25275;
  assign n25277 = n25223 & n25229;
  assign n25278 = n25248 & n25277;
  assign n25279 = n25235 & n25278;
  assign n25280 = n25229 & ~n25235;
  assign n25281 = ~n25247 & n25280;
  assign n25282 = n25241 & n25281;
  assign n25283 = ~n25223 & n25235;
  assign n25284 = ~n25247 & n25283;
  assign n25285 = ~n25241 & n25284;
  assign n25286 = ~n25282 & ~n25285;
  assign n25287 = ~n25279 & n25286;
  assign n25288 = ~n25276 & n25287;
  assign n25289 = n25270 & n25288;
  assign n25290 = n25266 & ~n25289;
  assign n25291 = ~n25229 & n25269;
  assign n25292 = ~n25290 & ~n25291;
  assign n25293 = ~n25259 & n25292;
  assign n25294 = ~n25255 & n25293;
  assign n25295 = ~n25223 & n25229;
  assign n25296 = ~n25235 & ~n25241;
  assign n25297 = n25295 & n25296;
  assign n25298 = ~n25223 & n25249;
  assign n25299 = ~n25297 & ~n25298;
  assign n25300 = n25241 & ~n25247;
  assign n25301 = ~n25235 & n25300;
  assign n25302 = ~n25223 & n25301;
  assign n25303 = n25235 & n25300;
  assign n25304 = ~n25229 & n25303;
  assign n25305 = ~n25302 & ~n25304;
  assign n25306 = ~n25235 & n25248;
  assign n25307 = n25229 & n25306;
  assign n25308 = ~n25250 & ~n25307;
  assign n25309 = n25229 & n25267;
  assign n25310 = n25235 & ~n25247;
  assign n25311 = ~n25309 & ~n25310;
  assign n25312 = n25223 & ~n25311;
  assign n25313 = n25308 & ~n25312;
  assign n25314 = n25305 & n25313;
  assign n25315 = n25299 & n25314;
  assign n25316 = ~n25266 & ~n25315;
  assign n25317 = n25294 & ~n25316;
  assign n25318 = ~pi0361 & ~n25317;
  assign n25319 = pi0361 & n25294;
  assign n25320 = ~n25316 & n25319;
  assign po0386 = n25318 | n25320;
  assign n25322 = ~n25291 & ~n25297;
  assign n25323 = n25235 & n25267;
  assign n25324 = ~n25258 & ~n25323;
  assign n25325 = ~n25309 & n25324;
  assign n25326 = n25223 & ~n25325;
  assign n25327 = n25235 & n25256;
  assign n25328 = n25229 & n25327;
  assign n25329 = ~n25282 & ~n25328;
  assign n25330 = ~n25223 & ~n25229;
  assign n25331 = n25303 & n25330;
  assign n25332 = n25329 & ~n25331;
  assign n25333 = ~n25223 & n25306;
  assign n25334 = n25332 & ~n25333;
  assign n25335 = ~n25326 & n25334;
  assign n25336 = n25266 & ~n25335;
  assign n25337 = ~n25223 & n25256;
  assign n25338 = ~n25229 & n25337;
  assign n25339 = n25241 & n25251;
  assign n25340 = ~n25323 & ~n25339;
  assign n25341 = ~n25223 & ~n25340;
  assign n25342 = ~n25338 & ~n25341;
  assign n25343 = n25223 & ~n25229;
  assign n25344 = n25300 & n25343;
  assign n25345 = n25223 & n25249;
  assign n25346 = ~n25344 & ~n25345;
  assign n25347 = n25342 & n25346;
  assign n25348 = n25241 & n25273;
  assign n25349 = ~n25250 & ~n25348;
  assign n25350 = ~n25307 & n25349;
  assign n25351 = n25347 & n25350;
  assign n25352 = ~n25266 & ~n25351;
  assign n25353 = ~n25250 & n25329;
  assign n25354 = n25223 & ~n25353;
  assign n25355 = ~n25352 & ~n25354;
  assign n25356 = ~n25336 & n25355;
  assign n25357 = n25322 & n25356;
  assign n25358 = pi0367 & ~n25357;
  assign n25359 = ~pi0367 & n25357;
  assign po0387 = n25358 | n25359;
  assign n25361 = pi3385 & pi9040;
  assign n25362 = pi3230 & ~pi9040;
  assign n25363 = ~n25361 & ~n25362;
  assign n25364 = ~pi0333 & ~n25363;
  assign n25365 = pi0333 & n25363;
  assign n25366 = ~n25364 & ~n25365;
  assign n25367 = pi3254 & pi9040;
  assign n25368 = pi3205 & ~pi9040;
  assign n25369 = ~n25367 & ~n25368;
  assign n25370 = ~pi0336 & n25369;
  assign n25371 = pi0336 & ~n25369;
  assign n25372 = ~n25370 & ~n25371;
  assign n25373 = pi3209 & pi9040;
  assign n25374 = pi3256 & ~pi9040;
  assign n25375 = ~n25373 & ~n25374;
  assign n25376 = pi0326 & n25375;
  assign n25377 = ~pi0326 & ~n25375;
  assign n25378 = ~n25376 & ~n25377;
  assign n25379 = n25372 & ~n25378;
  assign n25380 = ~n25366 & n25379;
  assign n25381 = pi3197 & pi9040;
  assign n25382 = pi3213 & ~pi9040;
  assign n25383 = ~n25381 & ~n25382;
  assign n25384 = pi0322 & n25383;
  assign n25385 = ~pi0322 & ~n25383;
  assign n25386 = ~n25384 & ~n25385;
  assign n25387 = pi3282 & pi9040;
  assign n25388 = pi3209 & ~pi9040;
  assign n25389 = ~n25387 & ~n25388;
  assign n25390 = ~pi0337 & n25389;
  assign n25391 = pi0337 & ~n25389;
  assign n25392 = ~n25390 & ~n25391;
  assign n25393 = ~n25386 & n25392;
  assign n25394 = n25380 & n25393;
  assign n25395 = n25372 & n25378;
  assign n25396 = n25393 & n25395;
  assign n25397 = n25366 & n25396;
  assign n25398 = ~n25394 & ~n25397;
  assign n25399 = ~n25366 & ~n25386;
  assign n25400 = ~n25372 & n25399;
  assign n25401 = ~n25378 & n25400;
  assign n25402 = ~n25392 & n25401;
  assign n25403 = n25398 & ~n25402;
  assign n25404 = pi3215 & ~pi9040;
  assign n25405 = pi3205 & pi9040;
  assign n25406 = ~n25404 & ~n25405;
  assign n25407 = ~pi0341 & ~n25406;
  assign n25408 = pi0341 & n25406;
  assign n25409 = ~n25407 & ~n25408;
  assign n25410 = ~n25386 & ~n25392;
  assign n25411 = ~n25378 & n25410;
  assign n25412 = n25392 & n25395;
  assign n25413 = ~n25386 & n25412;
  assign n25414 = n25366 & ~n25378;
  assign n25415 = n25386 & n25414;
  assign n25416 = n25366 & ~n25386;
  assign n25417 = n25378 & n25416;
  assign n25418 = ~n25415 & ~n25417;
  assign n25419 = n25392 & ~n25418;
  assign n25420 = ~n25413 & ~n25419;
  assign n25421 = n25366 & n25395;
  assign n25422 = ~n25386 & n25421;
  assign n25423 = ~n25366 & n25378;
  assign n25424 = ~n25372 & n25423;
  assign n25425 = n25386 & n25424;
  assign n25426 = ~n25422 & ~n25425;
  assign n25427 = n25386 & ~n25392;
  assign n25428 = n25423 & n25427;
  assign n25429 = ~n25372 & ~n25378;
  assign n25430 = ~n25366 & n25429;
  assign n25431 = ~n25392 & n25430;
  assign n25432 = ~n25428 & ~n25431;
  assign n25433 = n25426 & n25432;
  assign n25434 = n25420 & n25433;
  assign n25435 = ~n25411 & n25434;
  assign n25436 = ~n25409 & ~n25435;
  assign n25437 = ~n25372 & n25378;
  assign n25438 = n25366 & n25437;
  assign n25439 = ~n25415 & ~n25438;
  assign n25440 = ~n25366 & n25395;
  assign n25441 = ~n25386 & n25440;
  assign n25442 = n25439 & ~n25441;
  assign n25443 = ~n25392 & ~n25442;
  assign n25444 = ~n25386 & n25424;
  assign n25445 = n25366 & n25429;
  assign n25446 = ~n25386 & n25445;
  assign n25447 = ~n25366 & ~n25378;
  assign n25448 = ~n25395 & ~n25447;
  assign n25449 = n25386 & ~n25448;
  assign n25450 = ~n25446 & ~n25449;
  assign n25451 = ~n25444 & n25450;
  assign n25452 = n25392 & ~n25451;
  assign n25453 = ~n25443 & ~n25452;
  assign n25454 = n25409 & ~n25453;
  assign n25455 = n25386 & n25437;
  assign n25456 = n25366 & n25379;
  assign n25457 = ~n25386 & n25456;
  assign n25458 = ~n25455 & ~n25457;
  assign n25459 = ~n25392 & ~n25458;
  assign n25460 = ~n25454 & ~n25459;
  assign n25461 = ~n25436 & n25460;
  assign n25462 = n25403 & n25461;
  assign n25463 = ~pi0360 & ~n25462;
  assign n25464 = pi0360 & n25462;
  assign po0391 = n25463 | n25464;
  assign n25466 = n25392 & ~n25409;
  assign n25467 = ~n25386 & n25414;
  assign n25468 = n25386 & n25421;
  assign n25469 = ~n25386 & n25437;
  assign n25470 = ~n25468 & ~n25469;
  assign n25471 = ~n25467 & n25470;
  assign n25472 = n25466 & ~n25471;
  assign n25473 = n25372 & n25399;
  assign n25474 = n25386 & n25456;
  assign n25475 = ~n25473 & ~n25474;
  assign n25476 = ~n25438 & ~n25440;
  assign n25477 = n25475 & n25476;
  assign n25478 = ~n25392 & ~n25477;
  assign n25479 = n25386 & n25430;
  assign n25480 = ~n25478 & ~n25479;
  assign n25481 = ~n25409 & ~n25480;
  assign n25482 = ~n25472 & ~n25481;
  assign n25483 = n25366 & n25410;
  assign n25484 = ~n25372 & n25483;
  assign n25485 = ~n25441 & ~n25484;
  assign n25486 = ~n25379 & ~n25437;
  assign n25487 = n25386 & ~n25486;
  assign n25488 = ~n25380 & ~n25487;
  assign n25489 = n25392 & ~n25488;
  assign n25490 = ~n25445 & ~n25467;
  assign n25491 = ~n25468 & n25490;
  assign n25492 = ~n25392 & ~n25491;
  assign n25493 = ~n25489 & ~n25492;
  assign n25494 = ~n25366 & n25386;
  assign n25495 = n25372 & n25494;
  assign n25496 = ~n25378 & n25495;
  assign n25497 = ~n25425 & ~n25496;
  assign n25498 = ~n25401 & n25497;
  assign n25499 = ~n25413 & n25498;
  assign n25500 = n25493 & n25499;
  assign n25501 = n25409 & ~n25500;
  assign n25502 = n25485 & ~n25501;
  assign n25503 = n25482 & n25502;
  assign n25504 = pi0354 & ~n25503;
  assign n25505 = ~pi0354 & n25485;
  assign n25506 = n25482 & n25505;
  assign n25507 = ~n25501 & n25506;
  assign po0392 = n25504 | n25507;
  assign n25509 = pi3216 & pi9040;
  assign n25510 = pi3204 & ~pi9040;
  assign n25511 = ~n25509 & ~n25510;
  assign n25512 = ~pi0330 & ~n25511;
  assign n25513 = pi0330 & n25511;
  assign n25514 = ~n25512 & ~n25513;
  assign n25515 = pi3206 & pi9040;
  assign n25516 = pi3290 & ~pi9040;
  assign n25517 = ~n25515 & ~n25516;
  assign n25518 = pi0338 & n25517;
  assign n25519 = ~pi0338 & ~n25517;
  assign n25520 = ~n25518 & ~n25519;
  assign n25521 = pi3204 & pi9040;
  assign n25522 = pi3223 & ~pi9040;
  assign n25523 = ~n25521 & ~n25522;
  assign n25524 = ~pi0339 & n25523;
  assign n25525 = pi0339 & ~n25523;
  assign n25526 = ~n25524 & ~n25525;
  assign n25527 = n25520 & n25526;
  assign n25528 = pi3290 & pi9040;
  assign n25529 = pi3202 & ~pi9040;
  assign n25530 = ~n25528 & ~n25529;
  assign n25531 = ~pi0302 & n25530;
  assign n25532 = pi0302 & ~n25530;
  assign n25533 = ~n25531 & ~n25532;
  assign n25534 = pi3238 & pi9040;
  assign n25535 = pi3294 & ~pi9040;
  assign n25536 = ~n25534 & ~n25535;
  assign n25537 = ~pi0329 & ~n25536;
  assign n25538 = pi0329 & n25536;
  assign n25539 = ~n25537 & ~n25538;
  assign n25540 = pi3221 & pi9040;
  assign n25541 = pi3203 & ~pi9040;
  assign n25542 = ~n25540 & ~n25541;
  assign n25543 = ~pi0349 & n25542;
  assign n25544 = pi0349 & ~n25542;
  assign n25545 = ~n25543 & ~n25544;
  assign n25546 = n25539 & ~n25545;
  assign n25547 = n25533 & n25546;
  assign n25548 = ~n25539 & n25545;
  assign n25549 = ~n25547 & ~n25548;
  assign n25550 = n25527 & ~n25549;
  assign n25551 = n25526 & n25533;
  assign n25552 = n25548 & n25551;
  assign n25553 = ~n25550 & ~n25552;
  assign n25554 = n25514 & ~n25553;
  assign n25555 = ~n25533 & n25546;
  assign n25556 = ~n25520 & n25555;
  assign n25557 = ~n25533 & n25539;
  assign n25558 = ~n25520 & ~n25533;
  assign n25559 = ~n25557 & ~n25558;
  assign n25560 = ~n25526 & ~n25559;
  assign n25561 = ~n25520 & n25533;
  assign n25562 = n25545 & n25561;
  assign n25563 = n25539 & n25562;
  assign n25564 = ~n25560 & ~n25563;
  assign n25565 = ~n25556 & n25564;
  assign n25566 = n25514 & ~n25565;
  assign n25567 = ~n25554 & ~n25566;
  assign n25568 = n25520 & ~n25533;
  assign n25569 = ~n25545 & n25568;
  assign n25570 = ~n25539 & n25569;
  assign n25571 = ~n25539 & ~n25545;
  assign n25572 = n25533 & n25571;
  assign n25573 = ~n25520 & n25572;
  assign n25574 = ~n25570 & ~n25573;
  assign n25575 = n25526 & ~n25574;
  assign n25576 = ~n25533 & n25545;
  assign n25577 = ~n25572 & ~n25576;
  assign n25578 = ~n25520 & ~n25577;
  assign n25579 = ~n25520 & ~n25545;
  assign n25580 = n25526 & n25579;
  assign n25581 = n25533 & n25580;
  assign n25582 = n25539 & n25545;
  assign n25583 = ~n25557 & ~n25582;
  assign n25584 = n25520 & ~n25583;
  assign n25585 = ~n25572 & ~n25584;
  assign n25586 = n25526 & ~n25585;
  assign n25587 = n25520 & ~n25526;
  assign n25588 = n25546 & n25587;
  assign n25589 = n25533 & n25588;
  assign n25590 = ~n25586 & ~n25589;
  assign n25591 = ~n25581 & n25590;
  assign n25592 = ~n25578 & n25591;
  assign n25593 = ~n25570 & n25592;
  assign n25594 = ~n25514 & ~n25593;
  assign n25595 = ~n25520 & n25557;
  assign n25596 = n25520 & n25533;
  assign n25597 = n25545 & n25596;
  assign n25598 = ~n25539 & n25597;
  assign n25599 = ~n25595 & ~n25598;
  assign n25600 = ~n25526 & ~n25599;
  assign n25601 = ~n25594 & ~n25600;
  assign n25602 = ~n25575 & n25601;
  assign n25603 = n25567 & n25602;
  assign n25604 = pi0364 & n25603;
  assign n25605 = ~pi0364 & ~n25603;
  assign po0393 = n25604 | n25605;
  assign n25607 = ~n25102 & n25146;
  assign n25608 = ~n25186 & ~n25607;
  assign n25609 = n25108 & ~n25608;
  assign n25610 = n25132 & n25143;
  assign n25611 = ~n25609 & ~n25610;
  assign n25612 = ~n25156 & n25611;
  assign n25613 = ~n25089 & n25102;
  assign n25614 = n25083 & n25613;
  assign n25615 = n25095 & n25614;
  assign n25616 = ~n25116 & ~n25615;
  assign n25617 = ~n25146 & n25616;
  assign n25618 = n25108 & ~n25617;
  assign n25619 = n25077 & n25618;
  assign n25620 = ~n25083 & ~n25108;
  assign n25621 = n25095 & n25620;
  assign n25622 = n25089 & n25621;
  assign n25623 = ~n25102 & n25622;
  assign n25624 = ~n25108 & n25195;
  assign n25625 = ~n25127 & ~n25154;
  assign n25626 = ~n25121 & n25625;
  assign n25627 = ~n25624 & n25626;
  assign n25628 = n25077 & ~n25627;
  assign n25629 = n25102 & n25164;
  assign n25630 = ~n25622 & ~n25629;
  assign n25631 = ~n25185 & n25630;
  assign n25632 = n25095 & n25125;
  assign n25633 = n25102 & n25113;
  assign n25634 = ~n25142 & ~n25633;
  assign n25635 = n25108 & ~n25634;
  assign n25636 = ~n25632 & ~n25635;
  assign n25637 = n25631 & n25636;
  assign n25638 = ~n25077 & ~n25637;
  assign n25639 = ~n25628 & ~n25638;
  assign n25640 = ~n25623 & n25639;
  assign n25641 = ~n25619 & n25640;
  assign n25642 = n25612 & n25641;
  assign n25643 = pi0381 & ~n25642;
  assign n25644 = ~pi0381 & n25612;
  assign n25645 = n25641 & n25644;
  assign po0394 = n25643 | n25645;
  assign n25647 = n25229 & n25268;
  assign n25648 = ~n25229 & n25306;
  assign n25649 = ~n25647 & ~n25648;
  assign n25650 = n25229 & n25257;
  assign n25651 = n25229 & n25300;
  assign n25652 = ~n25229 & n25327;
  assign n25653 = ~n25651 & ~n25652;
  assign n25654 = n25223 & ~n25653;
  assign n25655 = ~n25650 & ~n25654;
  assign n25656 = n25229 & n25337;
  assign n25657 = ~n25298 & ~n25656;
  assign n25658 = n25655 & n25657;
  assign n25659 = n25649 & n25658;
  assign n25660 = n25266 & ~n25659;
  assign n25661 = n25223 & ~n25266;
  assign n25662 = ~n25241 & n25251;
  assign n25663 = n25235 & n25247;
  assign n25664 = ~n25662 & ~n25663;
  assign n25665 = n25661 & ~n25664;
  assign n25666 = ~n25258 & ~n25272;
  assign n25667 = ~n25235 & n25295;
  assign n25668 = ~n25256 & n25667;
  assign n25669 = ~n25269 & ~n25668;
  assign n25670 = n25666 & n25669;
  assign n25671 = ~n25266 & ~n25670;
  assign n25672 = n25323 & n25343;
  assign n25673 = ~n25229 & n25301;
  assign n25674 = ~n25648 & ~n25673;
  assign n25675 = n25223 & ~n25674;
  assign n25676 = ~n25672 & ~n25675;
  assign n25677 = n25257 & n25330;
  assign n25678 = n25676 & ~n25677;
  assign n25679 = ~n25671 & n25678;
  assign n25680 = ~n25665 & n25679;
  assign n25681 = ~n25660 & n25680;
  assign n25682 = ~n25331 & n25681;
  assign n25683 = ~pi0357 & ~n25682;
  assign n25684 = pi0357 & ~n25331;
  assign n25685 = n25680 & n25684;
  assign n25686 = ~n25660 & n25685;
  assign po0395 = n25683 | n25686;
  assign n25688 = ~n25520 & n25548;
  assign n25689 = ~n25533 & ~n25539;
  assign n25690 = ~n25545 & n25689;
  assign n25691 = ~n25688 & ~n25690;
  assign n25692 = ~n25514 & ~n25526;
  assign n25693 = ~n25691 & n25692;
  assign n25694 = n25568 & n25582;
  assign n25695 = n25533 & n25548;
  assign n25696 = ~n25547 & ~n25695;
  assign n25697 = n25520 & ~n25696;
  assign n25698 = ~n25694 & ~n25697;
  assign n25699 = ~n25514 & ~n25698;
  assign n25700 = ~n25693 & ~n25699;
  assign n25701 = ~n25539 & n25596;
  assign n25702 = ~n25694 & ~n25701;
  assign n25703 = n25526 & ~n25702;
  assign n25704 = ~n25520 & ~n25526;
  assign n25705 = n25539 & n25704;
  assign n25706 = n25533 & n25582;
  assign n25707 = ~n25555 & ~n25706;
  assign n25708 = ~n25533 & n25548;
  assign n25709 = n25520 & n25708;
  assign n25710 = n25707 & ~n25709;
  assign n25711 = ~n25526 & ~n25710;
  assign n25712 = ~n25705 & ~n25711;
  assign n25713 = n25520 & n25572;
  assign n25714 = n25712 & ~n25713;
  assign n25715 = n25526 & ~n25691;
  assign n25716 = ~n25520 & n25547;
  assign n25717 = ~n25715 & ~n25716;
  assign n25718 = n25714 & n25717;
  assign n25719 = n25514 & ~n25718;
  assign n25720 = ~n25703 & ~n25719;
  assign n25721 = ~n25514 & n25526;
  assign n25722 = ~n25520 & n25582;
  assign n25723 = ~n25572 & ~n25722;
  assign n25724 = ~n25557 & n25723;
  assign n25725 = n25721 & ~n25724;
  assign n25726 = n25720 & ~n25725;
  assign n25727 = n25700 & n25726;
  assign n25728 = ~pi0358 & ~n25727;
  assign n25729 = pi0358 & n25700;
  assign n25730 = n25720 & n25729;
  assign n25731 = ~n25725 & n25730;
  assign po0396 = n25728 | n25731;
  assign n25733 = ~n24852 & n24874;
  assign n25734 = ~n25053 & ~n25733;
  assign n25735 = n24858 & n25734;
  assign n25736 = n24852 & n24920;
  assign n25737 = ~n24868 & ~n24886;
  assign n25738 = n24867 & ~n25737;
  assign n25739 = ~n24840 & n24901;
  assign n25740 = n24852 & n24868;
  assign n25741 = ~n25739 & ~n25740;
  assign n25742 = ~n24858 & n25741;
  assign n25743 = ~n25738 & n25742;
  assign n25744 = ~n25736 & n25743;
  assign n25745 = ~n25735 & ~n25744;
  assign n25746 = n24852 & n25738;
  assign n25747 = ~n25051 & ~n25746;
  assign n25748 = ~n25745 & n25747;
  assign n25749 = n24834 & ~n25748;
  assign n25750 = n24858 & ~n25737;
  assign n25751 = ~n24852 & n25750;
  assign n25752 = n24852 & n24914;
  assign n25753 = ~n24891 & ~n25752;
  assign n25754 = n24858 & ~n25753;
  assign n25755 = ~n24867 & n25750;
  assign n25756 = ~n25754 & ~n25755;
  assign n25757 = ~n25751 & n25756;
  assign n25758 = ~n24834 & ~n25757;
  assign n25759 = ~n25749 & ~n25758;
  assign n25760 = n24858 & n24872;
  assign n25761 = ~n24858 & ~n25747;
  assign n25762 = ~n25760 & ~n25761;
  assign n25763 = ~n24858 & ~n25734;
  assign n25764 = ~n24872 & ~n25763;
  assign n25765 = ~n24834 & ~n25764;
  assign n25766 = n25762 & ~n25765;
  assign n25767 = n25759 & n25766;
  assign n25768 = pi0385 & ~n25767;
  assign n25769 = ~pi0385 & n25766;
  assign n25770 = ~n25758 & n25769;
  assign n25771 = ~n25749 & n25770;
  assign po0399 = n25768 | n25771;
  assign n25773 = ~n25380 & ~n25445;
  assign n25774 = n25392 & ~n25773;
  assign n25775 = n25386 & n25438;
  assign n25776 = ~n25774 & ~n25775;
  assign n25777 = n25378 & n25386;
  assign n25778 = ~n25423 & ~n25777;
  assign n25779 = ~n25456 & n25778;
  assign n25780 = ~n25392 & ~n25779;
  assign n25781 = n25776 & ~n25780;
  assign n25782 = ~n25409 & ~n25781;
  assign n25783 = n25392 & n25444;
  assign n25784 = ~n25397 & ~n25783;
  assign n25785 = ~n25402 & n25784;
  assign n25786 = n25378 & ~n25392;
  assign n25787 = n25416 & n25786;
  assign n25788 = n25386 & n25445;
  assign n25789 = n25392 & n25423;
  assign n25790 = ~n25788 & ~n25789;
  assign n25791 = ~n25496 & n25790;
  assign n25792 = ~n25787 & n25791;
  assign n25793 = n25372 & n25416;
  assign n25794 = ~n25401 & ~n25793;
  assign n25795 = n25792 & n25794;
  assign n25796 = ~n25431 & n25795;
  assign n25797 = n25409 & ~n25796;
  assign n25798 = n25785 & ~n25797;
  assign n25799 = ~n25782 & n25798;
  assign n25800 = ~pi0366 & ~n25799;
  assign n25801 = pi0366 & n25785;
  assign n25802 = ~n25782 & n25801;
  assign n25803 = ~n25797 & n25802;
  assign po0400 = n25800 | n25803;
  assign n25805 = ~n25647 & ~n25662;
  assign n25806 = n25266 & ~n25805;
  assign n25807 = n25223 & n25257;
  assign n25808 = ~n25247 & n25273;
  assign n25809 = ~n25274 & ~n25808;
  assign n25810 = n25223 & ~n25809;
  assign n25811 = ~n25807 & ~n25810;
  assign n25812 = n25266 & ~n25811;
  assign n25813 = ~n25806 & ~n25812;
  assign n25814 = n25268 & n25277;
  assign n25815 = ~n25279 & ~n25814;
  assign n25816 = ~n25272 & ~n25310;
  assign n25817 = ~n25223 & ~n25816;
  assign n25818 = n25266 & n25817;
  assign n25819 = n25815 & ~n25818;
  assign n25820 = n25247 & n25273;
  assign n25821 = n25241 & n25820;
  assign n25822 = ~n25229 & n25248;
  assign n25823 = ~n25253 & ~n25822;
  assign n25824 = ~n25223 & ~n25823;
  assign n25825 = ~n25258 & ~n25282;
  assign n25826 = ~n25229 & n25267;
  assign n25827 = ~n25303 & ~n25826;
  assign n25828 = n25223 & ~n25827;
  assign n25829 = n25825 & ~n25828;
  assign n25830 = ~n25824 & n25829;
  assign n25831 = ~n25821 & n25830;
  assign n25832 = ~n25266 & ~n25831;
  assign n25833 = ~n25307 & n25329;
  assign n25834 = ~n25223 & ~n25833;
  assign n25835 = ~n25832 & ~n25834;
  assign n25836 = n25819 & n25835;
  assign n25837 = n25813 & n25836;
  assign n25838 = ~pi0375 & ~n25837;
  assign n25839 = pi0375 & n25819;
  assign n25840 = n25813 & n25839;
  assign n25841 = n25835 & n25840;
  assign po0401 = n25838 | n25841;
  assign n25843 = pi3322 & pi9040;
  assign n25844 = pi3218 & ~pi9040;
  assign n25845 = ~n25843 & ~n25844;
  assign n25846 = pi0326 & n25845;
  assign n25847 = ~pi0326 & ~n25845;
  assign n25848 = ~n25846 & ~n25847;
  assign n25849 = pi3214 & pi9040;
  assign n25850 = pi3199 & ~pi9040;
  assign n25851 = ~n25849 & ~n25850;
  assign n25852 = pi0351 & n25851;
  assign n25853 = ~pi0351 & ~n25851;
  assign n25854 = ~n25852 & ~n25853;
  assign n25855 = pi3333 & pi9040;
  assign n25856 = pi3253 & ~pi9040;
  assign n25857 = ~n25855 & ~n25856;
  assign n25858 = pi0346 & n25857;
  assign n25859 = ~pi0346 & ~n25857;
  assign n25860 = ~n25858 & ~n25859;
  assign n25861 = pi3201 & pi9040;
  assign n25862 = pi3302 & ~pi9040;
  assign n25863 = ~n25861 & ~n25862;
  assign n25864 = ~pi0328 & n25863;
  assign n25865 = pi0328 & ~n25863;
  assign n25866 = ~n25864 & ~n25865;
  assign n25867 = pi3252 & pi9040;
  assign n25868 = pi3385 & ~pi9040;
  assign n25869 = ~n25867 & ~n25868;
  assign n25870 = pi0333 & n25869;
  assign n25871 = ~pi0333 & ~n25869;
  assign n25872 = ~n25870 & ~n25871;
  assign n25873 = ~n25866 & ~n25872;
  assign n25874 = n25860 & n25873;
  assign n25875 = n25854 & n25874;
  assign n25876 = ~n25854 & ~n25866;
  assign n25877 = n25872 & n25876;
  assign n25878 = pi3302 & pi9040;
  assign n25879 = pi3258 & ~pi9040;
  assign n25880 = ~n25878 & ~n25879;
  assign n25881 = ~pi0324 & n25880;
  assign n25882 = pi0324 & ~n25880;
  assign n25883 = ~n25881 & ~n25882;
  assign n25884 = ~n25860 & n25876;
  assign n25885 = ~pi0346 & n25857;
  assign n25886 = pi0346 & ~n25857;
  assign n25887 = ~n25885 & ~n25886;
  assign n25888 = n25872 & ~n25887;
  assign n25889 = n25866 & n25888;
  assign n25890 = ~n25884 & ~n25889;
  assign n25891 = n25883 & ~n25890;
  assign n25892 = ~n25877 & ~n25891;
  assign n25893 = ~n25866 & n25888;
  assign n25894 = n25866 & n25887;
  assign n25895 = n25866 & ~n25872;
  assign n25896 = ~n25854 & n25895;
  assign n25897 = ~n25860 & ~n25872;
  assign n25898 = n25854 & n25897;
  assign n25899 = ~n25896 & ~n25898;
  assign n25900 = ~n25894 & n25899;
  assign n25901 = ~n25893 & n25900;
  assign n25902 = ~n25883 & ~n25901;
  assign n25903 = n25892 & ~n25902;
  assign n25904 = ~n25875 & n25903;
  assign n25905 = n25848 & ~n25904;
  assign n25906 = ~n25860 & n25872;
  assign n25907 = n25866 & n25906;
  assign n25908 = ~n25854 & n25907;
  assign n25909 = n25866 & n25897;
  assign n25910 = n25854 & n25909;
  assign n25911 = ~n25875 & ~n25910;
  assign n25912 = ~n25908 & n25911;
  assign n25913 = ~n25883 & ~n25912;
  assign n25914 = ~n25905 & ~n25913;
  assign n25915 = ~n25854 & n25893;
  assign n25916 = n25866 & ~n25887;
  assign n25917 = n25883 & n25916;
  assign n25918 = n25854 & n25917;
  assign n25919 = n25854 & ~n25866;
  assign n25920 = n25872 & n25919;
  assign n25921 = ~n25860 & n25920;
  assign n25922 = ~n25872 & ~n25883;
  assign n25923 = ~n25866 & n25922;
  assign n25924 = ~n25854 & n25923;
  assign n25925 = ~n25921 & ~n25924;
  assign n25926 = ~n25860 & ~n25866;
  assign n25927 = n25854 & n25926;
  assign n25928 = ~n25872 & ~n25887;
  assign n25929 = n25866 & n25928;
  assign n25930 = ~n25927 & ~n25929;
  assign n25931 = n25883 & ~n25930;
  assign n25932 = n25883 & n25894;
  assign n25933 = ~n25854 & n25932;
  assign n25934 = ~n25931 & ~n25933;
  assign n25935 = n25925 & n25934;
  assign n25936 = ~n25848 & ~n25935;
  assign n25937 = ~n25918 & ~n25936;
  assign n25938 = ~n25915 & n25937;
  assign n25939 = n25914 & n25938;
  assign n25940 = ~pi0356 & ~n25939;
  assign n25941 = ~n25905 & ~n25915;
  assign n25942 = ~n25913 & n25941;
  assign n25943 = n25937 & n25942;
  assign n25944 = pi0356 & n25943;
  assign po0402 = n25940 | n25944;
  assign n25946 = n24858 & n24900;
  assign n25947 = n24901 & ~n25737;
  assign n25948 = ~n24915 & ~n25947;
  assign n25949 = ~n25051 & n25948;
  assign n25950 = ~n24858 & ~n25949;
  assign n25951 = n24852 & n24869;
  assign n25952 = ~n25950 & ~n25951;
  assign n25953 = ~n24867 & n24914;
  assign n25954 = ~n24852 & n25058;
  assign n25955 = ~n25953 & ~n25954;
  assign n25956 = ~n25740 & n25955;
  assign n25957 = n24858 & ~n25956;
  assign n25958 = n25952 & ~n25957;
  assign n25959 = n24834 & ~n25958;
  assign n25960 = ~n25946 & ~n25959;
  assign n25961 = ~n24852 & n24868;
  assign n25962 = ~n24895 & ~n25961;
  assign n25963 = n24858 & ~n25962;
  assign n25964 = ~n24916 & ~n25963;
  assign n25965 = ~n24891 & ~n24900;
  assign n25966 = n24852 & n24927;
  assign n25967 = ~n25058 & ~n25966;
  assign n25968 = ~n25953 & n25967;
  assign n25969 = ~n24858 & ~n25968;
  assign n25970 = ~n24852 & n24869;
  assign n25971 = ~n25969 & ~n25970;
  assign n25972 = n25965 & n25971;
  assign n25973 = n25964 & n25972;
  assign n25974 = ~n24834 & ~n25973;
  assign n25975 = ~n24908 & ~n25736;
  assign n25976 = ~n24858 & ~n25975;
  assign n25977 = ~n25974 & ~n25976;
  assign n25978 = n25960 & n25977;
  assign n25979 = pi0390 & n25978;
  assign n25980 = ~pi0390 & ~n25978;
  assign po0403 = n25979 | n25980;
  assign n25982 = n25102 & ~n25207;
  assign n25983 = n25083 & n25982;
  assign n25984 = n25095 & n25184;
  assign n25985 = ~n25166 & ~n25984;
  assign n25986 = ~n25116 & n25985;
  assign n25987 = ~n25108 & ~n25986;
  assign n25988 = ~n25130 & ~n25195;
  assign n25989 = n25108 & ~n25988;
  assign n25990 = ~n25987 & ~n25989;
  assign n25991 = ~n25983 & n25990;
  assign n25992 = ~n25102 & n25143;
  assign n25993 = n25991 & ~n25992;
  assign n25994 = ~n25077 & ~n25993;
  assign n25995 = n25112 & ~n25988;
  assign n25996 = ~n25131 & ~n25146;
  assign n25997 = ~n25116 & ~n25143;
  assign n25998 = n25996 & n25997;
  assign n25999 = n25102 & ~n25998;
  assign n26000 = ~n25995 & ~n25999;
  assign n26001 = ~n25186 & n26000;
  assign n26002 = n25077 & ~n26001;
  assign n26003 = ~n25994 & ~n26002;
  assign n26004 = n25102 & n25195;
  assign n26005 = ~n25992 & ~n26004;
  assign n26006 = n25108 & ~n26005;
  assign n26007 = n26003 & ~n26006;
  assign n26008 = pi0370 & ~n26007;
  assign n26009 = ~pi0370 & ~n26006;
  assign n26010 = ~n26002 & n26009;
  assign n26011 = ~n25994 & n26010;
  assign po0404 = n26008 | n26011;
  assign n26013 = ~n25378 & ~n25386;
  assign n26014 = ~n25793 & ~n26013;
  assign n26015 = n25392 & ~n26014;
  assign n26016 = n25366 & n25386;
  assign n26017 = ~n25372 & n26016;
  assign n26018 = ~n26015 & ~n26017;
  assign n26019 = ~n25392 & n25437;
  assign n26020 = ~n25386 & n26019;
  assign n26021 = ~n25457 & ~n26020;
  assign n26022 = n26018 & n26021;
  assign n26023 = n25409 & ~n26022;
  assign n26024 = ~n25421 & ~n25425;
  assign n26025 = ~n25386 & n25429;
  assign n26026 = n26024 & ~n26025;
  assign n26027 = ~n25392 & ~n26026;
  assign n26028 = n25393 & n25437;
  assign n26029 = ~n25441 & ~n26028;
  assign n26030 = ~n26027 & n26029;
  assign n26031 = ~n25456 & ~n25479;
  assign n26032 = n25392 & ~n26031;
  assign n26033 = n26030 & ~n26032;
  assign n26034 = ~n25409 & ~n26033;
  assign n26035 = ~n26023 & ~n26034;
  assign n26036 = n25379 & ~n25386;
  assign n26037 = n25386 & ~n25476;
  assign n26038 = ~n26036 & ~n26037;
  assign n26039 = n25392 & ~n26038;
  assign n26040 = ~n25421 & n25773;
  assign n26041 = n25427 & ~n26040;
  assign n26042 = ~n26039 & ~n26041;
  assign n26043 = n26035 & n26042;
  assign n26044 = ~pi0362 & ~n26043;
  assign n26045 = ~n26034 & n26042;
  assign n26046 = pi0362 & n26045;
  assign n26047 = ~n26023 & n26046;
  assign po0405 = n26044 | n26047;
  assign n26049 = ~n25547 & ~n25597;
  assign n26050 = n25526 & ~n26049;
  assign n26051 = n25520 & n25571;
  assign n26052 = ~n25562 & ~n26051;
  assign n26053 = ~n25526 & ~n26052;
  assign n26054 = ~n25520 & n25708;
  assign n26055 = ~n25581 & ~n26054;
  assign n26056 = ~n25694 & n26055;
  assign n26057 = ~n26053 & n26056;
  assign n26058 = ~n26050 & n26057;
  assign n26059 = ~n25556 & ~n25570;
  assign n26060 = n26058 & n26059;
  assign n26061 = n25514 & ~n26060;
  assign n26062 = n25558 & n25582;
  assign n26063 = n25696 & ~n26062;
  assign n26064 = ~n25526 & ~n26063;
  assign n26065 = ~n25520 & n25690;
  assign n26066 = ~n26064 & ~n26065;
  assign n26067 = n25539 & n25596;
  assign n26068 = n25520 & n25546;
  assign n26069 = ~n26067 & ~n26068;
  assign n26070 = ~n25526 & ~n26069;
  assign n26071 = ~n25526 & n25571;
  assign n26072 = ~n25520 & n26071;
  assign n26073 = ~n26070 & ~n26072;
  assign n26074 = n26066 & n26073;
  assign n26075 = ~n25514 & ~n26074;
  assign n26076 = ~n25708 & ~n25713;
  assign n26077 = ~n25563 & n26076;
  assign n26078 = n25721 & ~n26077;
  assign n26079 = ~n26075 & ~n26078;
  assign n26080 = ~n25556 & ~n25694;
  assign n26081 = n25526 & ~n26080;
  assign n26082 = n26079 & ~n26081;
  assign n26083 = ~n26061 & n26082;
  assign n26084 = ~pi0380 & n26083;
  assign n26085 = pi0380 & ~n26083;
  assign po0406 = n26084 | n26085;
  assign n26087 = ~n25854 & n25874;
  assign n26088 = ~n25910 & ~n26087;
  assign n26089 = ~n25883 & ~n26088;
  assign n26090 = ~n25866 & n25897;
  assign n26091 = n25854 & n26090;
  assign n26092 = n25854 & n25907;
  assign n26093 = ~n26091 & ~n26092;
  assign n26094 = n25883 & ~n26093;
  assign n26095 = ~n26089 & ~n26094;
  assign n26096 = n25854 & n25883;
  assign n26097 = n25893 & n26096;
  assign n26098 = n25883 & n25909;
  assign n26099 = ~n25866 & n25906;
  assign n26100 = n25883 & n26099;
  assign n26101 = ~n26098 & ~n26100;
  assign n26102 = ~n25854 & ~n26101;
  assign n26103 = ~n26097 & ~n26102;
  assign n26104 = n25854 & n25906;
  assign n26105 = ~n25854 & n25888;
  assign n26106 = ~n26104 & ~n26105;
  assign n26107 = ~n25874 & n26106;
  assign n26108 = ~n25907 & n26107;
  assign n26109 = ~n25883 & ~n26108;
  assign n26110 = ~n25854 & n25889;
  assign n26111 = ~n26109 & ~n26110;
  assign n26112 = n25854 & ~n25887;
  assign n26113 = n25866 & n26112;
  assign n26114 = ~n25872 & n26113;
  assign n26115 = ~n26087 & ~n26114;
  assign n26116 = n26111 & n26115;
  assign n26117 = n26103 & n26116;
  assign n26118 = n25848 & ~n26117;
  assign n26119 = n25854 & n25888;
  assign n26120 = ~n25884 & ~n26119;
  assign n26121 = ~n25909 & n26120;
  assign n26122 = ~n25883 & ~n26121;
  assign n26123 = ~n25907 & ~n25915;
  assign n26124 = n25854 & n25873;
  assign n26125 = ~n25854 & n25929;
  assign n26126 = ~n26124 & ~n26125;
  assign n26127 = n26123 & n26126;
  assign n26128 = n25883 & ~n26127;
  assign n26129 = ~n26122 & ~n26128;
  assign n26130 = ~n25854 & n26090;
  assign n26131 = n25854 & n25889;
  assign n26132 = ~n26130 & ~n26131;
  assign n26133 = n26129 & n26132;
  assign n26134 = ~n25848 & ~n26133;
  assign n26135 = ~n26118 & ~n26134;
  assign n26136 = n26095 & n26135;
  assign n26137 = pi0365 & ~n26136;
  assign n26138 = ~pi0365 & n26136;
  assign po0407 = n26137 | n26138;
  assign n26140 = n24947 & n24953;
  assign n26141 = ~n24941 & n26140;
  assign n26142 = n24967 & n26141;
  assign n26143 = n24953 & n24985;
  assign n26144 = ~n24947 & ~n24959;
  assign n26145 = ~n24967 & n26144;
  assign n26146 = ~n24977 & ~n26145;
  assign n26147 = ~n26143 & n26146;
  assign n26148 = ~n26142 & n26147;
  assign n26149 = n24941 & n24973;
  assign n26150 = n26148 & ~n26149;
  assign n26151 = n25009 & ~n26150;
  assign n26152 = ~n24974 & ~n24977;
  assign n26153 = ~n24967 & n25026;
  assign n26154 = n24967 & n25011;
  assign n26155 = ~n26153 & ~n26154;
  assign n26156 = n26152 & n26155;
  assign n26157 = ~n24941 & ~n26156;
  assign n26158 = ~n26151 & ~n26157;
  assign n26159 = ~n24967 & n24979;
  assign n26160 = ~n25027 & ~n26159;
  assign n26161 = n24941 & ~n26160;
  assign n26162 = ~n24947 & ~n24967;
  assign n26163 = ~n24953 & n26162;
  assign n26164 = ~n26144 & ~n26163;
  assign n26165 = ~n24979 & n26164;
  assign n26166 = n24941 & ~n26165;
  assign n26167 = n24947 & n24996;
  assign n26168 = ~n24967 & n26167;
  assign n26169 = ~n26166 & ~n26168;
  assign n26170 = ~n25009 & ~n26169;
  assign n26171 = ~n25009 & n25011;
  assign n26172 = ~n24941 & n26171;
  assign n26173 = ~n26170 & ~n26172;
  assign n26174 = ~n26161 & n26173;
  assign n26175 = n26158 & n26174;
  assign n26176 = ~pi0379 & ~n26175;
  assign n26177 = pi0379 & n26158;
  assign n26178 = n26174 & n26177;
  assign po0408 = n26176 | n26178;
  assign n26180 = ~n24967 & n25000;
  assign n26181 = ~n24997 & ~n26154;
  assign n26182 = n24941 & ~n26181;
  assign n26183 = ~n26180 & ~n26182;
  assign n26184 = ~n24941 & ~n24967;
  assign n26185 = ~n24959 & n26184;
  assign n26186 = n24953 & n26185;
  assign n26187 = n24978 & n25012;
  assign n26188 = ~n26186 & ~n26187;
  assign n26189 = ~n24941 & ~n24947;
  assign n26190 = n24972 & n26189;
  assign n26191 = n26188 & ~n26190;
  assign n26192 = ~n24974 & ~n24986;
  assign n26193 = n24959 & n24976;
  assign n26194 = n26192 & ~n26193;
  assign n26195 = n26191 & n26194;
  assign n26196 = n26183 & n26195;
  assign n26197 = ~n25009 & ~n26196;
  assign n26198 = ~n24967 & n24996;
  assign n26199 = ~n26143 & ~n26198;
  assign n26200 = ~n24941 & ~n26199;
  assign n26201 = n24953 & n25015;
  assign n26202 = ~n25026 & ~n26201;
  assign n26203 = n24967 & n26144;
  assign n26204 = n26202 & ~n26203;
  assign n26205 = n24941 & ~n26204;
  assign n26206 = ~n24973 & ~n24997;
  assign n26207 = n24967 & ~n26206;
  assign n26208 = ~n26159 & ~n26207;
  assign n26209 = ~n26205 & n26208;
  assign n26210 = ~n26200 & n26209;
  assign n26211 = n25009 & ~n26210;
  assign n26212 = n24941 & n25016;
  assign n26213 = ~n26211 & ~n26212;
  assign n26214 = n24991 & n26184;
  assign n26215 = ~n24959 & n26214;
  assign n26216 = n26213 & ~n26215;
  assign n26217 = ~n26197 & n26216;
  assign n26218 = ~pi0368 & ~n26217;
  assign n26219 = pi0368 & n26213;
  assign n26220 = ~n26197 & n26219;
  assign n26221 = ~n26215 & n26220;
  assign po0409 = n26218 | n26221;
  assign n26223 = ~n25854 & n25866;
  assign n26224 = ~n25872 & n26223;
  assign n26225 = ~n25860 & n26224;
  assign n26226 = ~n25889 & ~n26225;
  assign n26227 = ~n25883 & ~n26226;
  assign n26228 = n26093 & ~n26227;
  assign n26229 = ~n25854 & n25883;
  assign n26230 = n25860 & n26229;
  assign n26231 = n26228 & ~n26230;
  assign n26232 = n25848 & ~n26231;
  assign n26233 = n25883 & n26114;
  assign n26234 = ~n25854 & ~n25883;
  assign n26235 = n25929 & n26234;
  assign n26236 = ~n25884 & ~n26235;
  assign n26237 = ~n25889 & ~n26099;
  assign n26238 = ~n25854 & n25906;
  assign n26239 = n26237 & ~n26238;
  assign n26240 = n25883 & ~n26239;
  assign n26241 = ~n25883 & n25893;
  assign n26242 = n25911 & ~n26241;
  assign n26243 = ~n26240 & n26242;
  assign n26244 = n26236 & n26243;
  assign n26245 = ~n25848 & ~n26244;
  assign n26246 = ~n26233 & ~n26245;
  assign n26247 = ~n26232 & n26246;
  assign n26248 = n26099 & n26234;
  assign n26249 = n25854 & n25923;
  assign n26250 = ~n26248 & ~n26249;
  assign n26251 = ~n25883 & n26092;
  assign n26252 = n26250 & ~n26251;
  assign n26253 = n26247 & n26252;
  assign n26254 = ~pi0353 & ~n26253;
  assign n26255 = pi0353 & n26252;
  assign n26256 = n26246 & n26255;
  assign n26257 = ~n26232 & n26256;
  assign po0410 = n26254 | n26257;
  assign n26259 = ~n24968 & ~n24977;
  assign n26260 = ~n24941 & ~n26259;
  assign n26261 = ~n25033 & ~n26260;
  assign n26262 = n24947 & ~n24953;
  assign n26263 = n24941 & n26262;
  assign n26264 = n24967 & n26263;
  assign n26265 = ~n24941 & n24960;
  assign n26266 = n24967 & n26265;
  assign n26267 = ~n26190 & ~n26266;
  assign n26268 = n24953 & n26162;
  assign n26269 = n24967 & n24996;
  assign n26270 = ~n26268 & ~n26269;
  assign n26271 = ~n26262 & n26270;
  assign n26272 = n24941 & ~n26271;
  assign n26273 = ~n24980 & ~n26272;
  assign n26274 = n26267 & n26273;
  assign n26275 = ~n25009 & ~n26274;
  assign n26276 = ~n26264 & ~n26275;
  assign n26277 = ~n24997 & ~n25016;
  assign n26278 = ~n25026 & n26277;
  assign n26279 = ~n24941 & ~n26278;
  assign n26280 = ~n24967 & n25021;
  assign n26281 = ~n25000 & ~n26280;
  assign n26282 = n24941 & ~n26281;
  assign n26283 = ~n26201 & ~n26282;
  assign n26284 = ~n26279 & n26283;
  assign n26285 = ~n24986 & ~n25027;
  assign n26286 = n26284 & n26285;
  assign n26287 = n25009 & ~n26286;
  assign n26288 = n26276 & ~n26287;
  assign n26289 = n26261 & n26288;
  assign n26290 = ~pi0377 & ~n26289;
  assign n26291 = pi0377 & n26276;
  assign n26292 = n26261 & n26291;
  assign n26293 = ~n26287 & n26292;
  assign po0411 = n26290 | n26293;
  assign n26295 = n25526 & n25690;
  assign n26296 = ~n25520 & n25546;
  assign n26297 = ~n25706 & ~n26296;
  assign n26298 = n25526 & ~n26297;
  assign n26299 = ~n25526 & ~n25577;
  assign n26300 = ~n26298 & ~n26299;
  assign n26301 = ~n25598 & n26300;
  assign n26302 = n25514 & ~n26301;
  assign n26303 = ~n26295 & ~n26302;
  assign n26304 = n25527 & ~n25533;
  assign n26305 = ~n25561 & ~n26304;
  assign n26306 = ~n25539 & ~n26305;
  assign n26307 = ~n25694 & ~n26306;
  assign n26308 = ~n25562 & n26307;
  assign n26309 = ~n25526 & n25555;
  assign n26310 = n25520 & n25547;
  assign n26311 = ~n26309 & ~n26310;
  assign n26312 = n26308 & n26311;
  assign n26313 = ~n25514 & ~n26312;
  assign n26314 = ~n26054 & ~n26068;
  assign n26315 = ~n25526 & ~n26314;
  assign n26316 = ~n26313 & ~n26315;
  assign n26317 = n26303 & n26316;
  assign n26318 = ~pi0398 & ~n26317;
  assign n26319 = pi0398 & n26316;
  assign n26320 = ~n26302 & n26319;
  assign n26321 = ~n26295 & n26320;
  assign po0412 = n26318 | n26321;
  assign n26323 = ~n26087 & ~n26225;
  assign n26324 = ~n26131 & n26323;
  assign n26325 = n25883 & ~n26324;
  assign n26326 = ~n26100 & ~n26114;
  assign n26327 = ~n26090 & ~n26105;
  assign n26328 = ~n25883 & ~n26327;
  assign n26329 = ~n25915 & ~n26328;
  assign n26330 = n26326 & n26329;
  assign n26331 = n25848 & ~n26330;
  assign n26332 = n25866 & n25872;
  assign n26333 = ~n25894 & ~n26332;
  assign n26334 = n25854 & ~n26333;
  assign n26335 = ~n25874 & ~n26238;
  assign n26336 = ~n25883 & ~n26335;
  assign n26337 = n25854 & n25872;
  assign n26338 = ~n25889 & ~n26337;
  assign n26339 = ~n25897 & n26338;
  assign n26340 = n25883 & ~n26339;
  assign n26341 = ~n26336 & ~n26340;
  assign n26342 = ~n26334 & n26341;
  assign n26343 = ~n25848 & ~n26342;
  assign n26344 = ~n26331 & ~n26343;
  assign n26345 = ~n26235 & ~n26251;
  assign n26346 = n26344 & n26345;
  assign n26347 = ~n26325 & n26346;
  assign n26348 = ~pi0378 & ~n26347;
  assign n26349 = pi0378 & n26345;
  assign n26350 = ~n26325 & n26349;
  assign n26351 = n26344 & n26350;
  assign po0413 = n26348 | n26351;
  assign n26353 = pi3223 & pi9040;
  assign n26354 = pi3259 & ~pi9040;
  assign n26355 = ~n26353 & ~n26354;
  assign n26356 = pi0349 & n26355;
  assign n26357 = ~pi0349 & ~n26355;
  assign n26358 = ~n26356 & ~n26357;
  assign n26359 = pi3203 & pi9040;
  assign n26360 = pi3220 & ~pi9040;
  assign n26361 = ~n26359 & ~n26360;
  assign n26362 = ~pi0330 & n26361;
  assign n26363 = pi0330 & ~n26361;
  assign n26364 = ~n26362 & ~n26363;
  assign n26365 = pi3220 & pi9040;
  assign n26366 = pi3216 & ~pi9040;
  assign n26367 = ~n26365 & ~n26366;
  assign n26368 = ~pi0344 & n26367;
  assign n26369 = pi0344 & ~n26367;
  assign n26370 = ~n26368 & ~n26369;
  assign n26371 = ~n26364 & ~n26370;
  assign n26372 = n26358 & n26371;
  assign n26373 = ~pi0344 & ~n26367;
  assign n26374 = pi0344 & n26367;
  assign n26375 = ~n26373 & ~n26374;
  assign n26376 = ~n26364 & ~n26375;
  assign n26377 = ~n26358 & n26376;
  assign n26378 = ~n26372 & ~n26377;
  assign n26379 = pi3263 & pi9040;
  assign n26380 = pi3233 & ~pi9040;
  assign n26381 = ~n26379 & ~n26380;
  assign n26382 = pi0327 & n26381;
  assign n26383 = ~pi0327 & ~n26381;
  assign n26384 = ~n26382 & ~n26383;
  assign n26385 = n26358 & ~n26384;
  assign n26386 = n26375 & n26385;
  assign n26387 = n26378 & ~n26386;
  assign n26388 = pi3259 & pi9040;
  assign n26389 = pi3222 & ~pi9040;
  assign n26390 = ~n26388 & ~n26389;
  assign n26391 = pi0315 & n26390;
  assign n26392 = ~pi0315 & ~n26390;
  assign n26393 = ~n26391 & ~n26392;
  assign n26394 = pi3210 & pi9040;
  assign n26395 = pi3212 & ~pi9040;
  assign n26396 = ~n26394 & ~n26395;
  assign n26397 = ~pi0323 & n26396;
  assign n26398 = pi0323 & ~n26396;
  assign n26399 = ~n26397 & ~n26398;
  assign n26400 = ~n26393 & ~n26399;
  assign n26401 = ~n26387 & n26400;
  assign n26402 = n26364 & ~n26375;
  assign n26403 = n26358 & n26402;
  assign n26404 = ~n26399 & n26403;
  assign n26405 = n26384 & n26404;
  assign n26406 = n26358 & n26376;
  assign n26407 = n26393 & n26406;
  assign n26408 = ~n26358 & n26375;
  assign n26409 = n26364 & ~n26370;
  assign n26410 = n26384 & n26409;
  assign n26411 = ~n26408 & ~n26410;
  assign n26412 = n26393 & ~n26411;
  assign n26413 = ~n26407 & ~n26412;
  assign n26414 = ~n26399 & ~n26413;
  assign n26415 = ~n26405 & ~n26414;
  assign n26416 = ~n26358 & n26384;
  assign n26417 = n26375 & n26416;
  assign n26418 = ~n26358 & ~n26384;
  assign n26419 = ~n26375 & n26418;
  assign n26420 = n26364 & n26419;
  assign n26421 = ~n26417 & ~n26420;
  assign n26422 = n26393 & ~n26421;
  assign n26423 = n26415 & ~n26422;
  assign n26424 = n26384 & ~n26393;
  assign n26425 = n26409 & n26424;
  assign n26426 = n26358 & n26425;
  assign n26427 = ~n26371 & ~n26402;
  assign n26428 = n26385 & ~n26427;
  assign n26429 = ~n26364 & n26419;
  assign n26430 = ~n26428 & ~n26429;
  assign n26431 = ~n26358 & n26409;
  assign n26432 = ~n26384 & ~n26393;
  assign n26433 = n26431 & n26432;
  assign n26434 = n26416 & ~n26427;
  assign n26435 = n26384 & n26406;
  assign n26436 = ~n26434 & ~n26435;
  assign n26437 = ~n26433 & n26436;
  assign n26438 = n26430 & n26437;
  assign n26439 = ~n26426 & n26438;
  assign n26440 = ~n26384 & n26393;
  assign n26441 = n26358 & n26440;
  assign n26442 = n26364 & n26441;
  assign n26443 = n26439 & ~n26442;
  assign n26444 = n26399 & ~n26443;
  assign n26445 = n26423 & ~n26444;
  assign n26446 = ~n26401 & n26445;
  assign n26447 = ~pi0369 & ~n26446;
  assign n26448 = pi0369 & n26423;
  assign n26449 = ~n26401 & n26448;
  assign n26450 = ~n26444 & n26449;
  assign po0414 = n26447 | n26450;
  assign n26452 = n26358 & n26409;
  assign n26453 = n26393 & n26452;
  assign n26454 = ~n26384 & n26453;
  assign n26455 = n26376 & n26440;
  assign n26456 = ~n26358 & n26455;
  assign n26457 = ~n26454 & ~n26456;
  assign n26458 = ~n26429 & ~n26433;
  assign n26459 = ~n26364 & n26384;
  assign n26460 = n26358 & n26459;
  assign n26461 = ~n26410 & ~n26460;
  assign n26462 = n26393 & ~n26461;
  assign n26463 = ~n26393 & ~n26418;
  assign n26464 = ~n26427 & n26463;
  assign n26465 = ~n26358 & ~n26409;
  assign n26466 = n26393 & n26465;
  assign n26467 = ~n26384 & n26466;
  assign n26468 = ~n26464 & ~n26467;
  assign n26469 = ~n26462 & n26468;
  assign n26470 = n26458 & n26469;
  assign n26471 = ~n26399 & ~n26470;
  assign n26472 = n26457 & ~n26471;
  assign n26473 = n26372 & ~n26393;
  assign n26474 = n26384 & n26473;
  assign n26475 = ~n26393 & n26399;
  assign n26476 = n26418 & ~n26427;
  assign n26477 = ~n26410 & ~n26476;
  assign n26478 = ~n26406 & n26477;
  assign n26479 = n26475 & ~n26478;
  assign n26480 = n26377 & n26384;
  assign n26481 = ~n26358 & n26459;
  assign n26482 = n26384 & n26402;
  assign n26483 = ~n26481 & ~n26482;
  assign n26484 = ~n26384 & n26409;
  assign n26485 = ~n26403 & ~n26484;
  assign n26486 = n26483 & n26485;
  assign n26487 = n26393 & ~n26486;
  assign n26488 = ~n26480 & ~n26487;
  assign n26489 = n26399 & ~n26488;
  assign n26490 = ~n26479 & ~n26489;
  assign n26491 = ~n26474 & n26490;
  assign n26492 = n26472 & n26491;
  assign n26493 = pi0371 & ~n26492;
  assign n26494 = ~pi0371 & n26472;
  assign n26495 = n26491 & n26494;
  assign po0415 = n26493 | n26495;
  assign n26497 = ~n26358 & n26371;
  assign n26498 = ~n26452 & ~n26497;
  assign n26499 = n26393 & ~n26498;
  assign n26500 = ~n26384 & n26402;
  assign n26501 = ~n26372 & ~n26500;
  assign n26502 = ~n26431 & n26501;
  assign n26503 = ~n26393 & ~n26502;
  assign n26504 = ~n26499 & ~n26503;
  assign n26505 = ~n26407 & ~n26420;
  assign n26506 = n26504 & n26505;
  assign n26507 = n26399 & ~n26506;
  assign n26508 = n26384 & n26452;
  assign n26509 = n26376 & ~n26384;
  assign n26510 = ~n26482 & ~n26509;
  assign n26511 = ~n26393 & ~n26510;
  assign n26512 = ~n26508 & ~n26511;
  assign n26513 = n26393 & n26403;
  assign n26514 = n26378 & ~n26513;
  assign n26515 = ~n26431 & n26514;
  assign n26516 = ~n26384 & ~n26515;
  assign n26517 = n26512 & ~n26516;
  assign n26518 = ~n26399 & ~n26517;
  assign n26519 = ~n26507 & ~n26518;
  assign n26520 = ~n26358 & n26482;
  assign n26521 = ~n26435 & ~n26520;
  assign n26522 = n26393 & ~n26521;
  assign n26523 = ~n26358 & ~n26364;
  assign n26524 = n26424 & n26523;
  assign n26525 = ~n26522 & ~n26524;
  assign n26526 = n26519 & n26525;
  assign n26527 = ~pi0363 & ~n26526;
  assign n26528 = pi0363 & ~n26522;
  assign n26529 = n26519 & n26528;
  assign n26530 = ~n26524 & n26529;
  assign po0416 = n26527 | n26530;
  assign n26532 = ~n26403 & ~n26459;
  assign n26533 = n26400 & ~n26532;
  assign n26534 = ~n26482 & ~n26484;
  assign n26535 = n26393 & ~n26534;
  assign n26536 = ~n26456 & ~n26535;
  assign n26537 = ~n26399 & ~n26536;
  assign n26538 = ~n26371 & ~n26523;
  assign n26539 = ~n26384 & ~n26538;
  assign n26540 = ~n26452 & ~n26539;
  assign n26541 = ~n26393 & ~n26540;
  assign n26542 = ~n26476 & ~n26541;
  assign n26543 = n26384 & n26431;
  assign n26544 = ~n26375 & n26385;
  assign n26545 = n26384 & ~n26538;
  assign n26546 = ~n26544 & ~n26545;
  assign n26547 = n26393 & ~n26546;
  assign n26548 = ~n26543 & ~n26547;
  assign n26549 = n26542 & n26548;
  assign n26550 = n26399 & ~n26549;
  assign n26551 = ~n26537 & ~n26550;
  assign n26552 = n26358 & n26384;
  assign n26553 = ~n26371 & n26552;
  assign n26554 = ~n26399 & n26553;
  assign n26555 = n26393 & n26416;
  assign n26556 = n26371 & n26555;
  assign n26557 = n26358 & n26424;
  assign n26558 = ~n26375 & n26557;
  assign n26559 = ~n26556 & ~n26558;
  assign n26560 = ~n26554 & n26559;
  assign n26561 = n26551 & n26560;
  assign n26562 = ~n26533 & n26561;
  assign n26563 = pi0372 & ~n26562;
  assign n26564 = ~pi0372 & n26560;
  assign n26565 = ~n26533 & n26564;
  assign n26566 = n26551 & n26565;
  assign po0417 = n26563 | n26566;
  assign n26568 = pi3321 & pi9040;
  assign n26569 = pi3402 & ~pi9040;
  assign n26570 = ~n26568 & ~n26569;
  assign n26571 = pi0402 & n26570;
  assign n26572 = ~pi0402 & ~n26570;
  assign n26573 = ~n26571 & ~n26572;
  assign n26574 = pi3287 & pi9040;
  assign n26575 = pi3315 & ~pi9040;
  assign n26576 = ~n26574 & ~n26575;
  assign n26577 = ~pi0382 & ~n26576;
  assign n26578 = pi0382 & ~n26574;
  assign n26579 = ~n26575 & n26578;
  assign n26580 = ~n26577 & ~n26579;
  assign n26581 = pi3283 & pi9040;
  assign n26582 = pi3335 & ~pi9040;
  assign n26583 = ~n26581 & ~n26582;
  assign n26584 = ~pi0405 & ~n26583;
  assign n26585 = pi0405 & ~n26581;
  assign n26586 = ~n26582 & n26585;
  assign n26587 = ~n26584 & ~n26586;
  assign n26588 = pi3334 & pi9040;
  assign n26589 = pi3352 & ~pi9040;
  assign n26590 = ~n26588 & ~n26589;
  assign n26591 = ~pi0389 & n26590;
  assign n26592 = pi0389 & ~n26590;
  assign n26593 = ~n26591 & ~n26592;
  assign n26594 = n26587 & ~n26593;
  assign n26595 = ~n26580 & n26594;
  assign n26596 = pi3289 & pi9040;
  assign n26597 = pi3280 & ~pi9040;
  assign n26598 = ~n26596 & ~n26597;
  assign n26599 = ~pi0401 & n26598;
  assign n26600 = pi0401 & ~n26598;
  assign n26601 = ~n26599 & ~n26600;
  assign n26602 = n26595 & n26601;
  assign n26603 = ~n26587 & n26593;
  assign n26604 = ~n26580 & n26603;
  assign n26605 = n26601 & n26604;
  assign n26606 = ~n26602 & ~n26605;
  assign n26607 = n26580 & ~n26601;
  assign n26608 = n26603 & n26607;
  assign n26609 = n26587 & n26593;
  assign n26610 = ~n26580 & n26609;
  assign n26611 = ~n26601 & n26610;
  assign n26612 = ~n26608 & ~n26611;
  assign n26613 = n26606 & n26612;
  assign n26614 = n26573 & ~n26613;
  assign n26615 = ~n26580 & ~n26601;
  assign n26616 = ~n26593 & n26615;
  assign n26617 = ~n26587 & n26616;
  assign n26618 = ~n26610 & ~n26617;
  assign n26619 = n26573 & ~n26618;
  assign n26620 = ~n26593 & n26601;
  assign n26621 = ~n26573 & n26620;
  assign n26622 = n26580 & n26587;
  assign n26623 = ~n26601 & n26603;
  assign n26624 = ~n26622 & ~n26623;
  assign n26625 = ~n26573 & ~n26624;
  assign n26626 = ~n26621 & ~n26625;
  assign n26627 = ~n26587 & ~n26593;
  assign n26628 = n26580 & n26627;
  assign n26629 = n26601 & n26628;
  assign n26630 = n26626 & ~n26629;
  assign n26631 = ~n26593 & n26622;
  assign n26632 = ~n26601 & n26631;
  assign n26633 = n26630 & ~n26632;
  assign n26634 = ~n26619 & n26633;
  assign n26635 = ~pi3421 & ~pi9040;
  assign n26636 = ~pi3285 & pi9040;
  assign n26637 = ~n26635 & ~n26636;
  assign n26638 = ~pi0415 & n26637;
  assign n26639 = pi0415 & ~n26637;
  assign n26640 = ~n26638 & ~n26639;
  assign n26641 = ~n26634 & ~n26640;
  assign n26642 = ~n26580 & ~n26593;
  assign n26643 = ~n26573 & ~n26601;
  assign n26644 = n26640 & n26643;
  assign n26645 = n26642 & n26644;
  assign n26646 = ~n26580 & n26601;
  assign n26647 = n26593 & n26646;
  assign n26648 = ~n26573 & ~n26647;
  assign n26649 = ~n26587 & n26607;
  assign n26650 = ~n26594 & ~n26642;
  assign n26651 = n26601 & ~n26650;
  assign n26652 = n26580 & n26603;
  assign n26653 = n26573 & ~n26652;
  assign n26654 = ~n26651 & n26653;
  assign n26655 = ~n26649 & n26654;
  assign n26656 = ~n26648 & ~n26655;
  assign n26657 = n26580 & n26609;
  assign n26658 = ~n26601 & n26657;
  assign n26659 = ~n26656 & ~n26658;
  assign n26660 = n26640 & ~n26659;
  assign n26661 = ~n26645 & ~n26660;
  assign n26662 = ~n26641 & n26661;
  assign n26663 = ~n26614 & n26662;
  assign n26664 = ~n26573 & n26629;
  assign n26665 = n26663 & ~n26664;
  assign n26666 = pi0421 & ~n26665;
  assign n26667 = n26662 & ~n26664;
  assign n26668 = ~pi0421 & n26667;
  assign n26669 = ~n26614 & n26668;
  assign po0432 = n26666 | n26669;
  assign n26671 = pi3402 & pi9040;
  assign n26672 = pi3277 & ~pi9040;
  assign n26673 = ~n26671 & ~n26672;
  assign n26674 = ~pi0411 & n26673;
  assign n26675 = pi0411 & ~n26673;
  assign n26676 = ~n26674 & ~n26675;
  assign n26677 = pi3287 & ~pi9040;
  assign n26678 = pi3286 & pi9040;
  assign n26679 = ~n26677 & ~n26678;
  assign n26680 = ~pi0400 & ~n26679;
  assign n26681 = pi0400 & n26679;
  assign n26682 = ~n26680 & ~n26681;
  assign n26683 = n26676 & ~n26682;
  assign n26684 = pi3315 & pi9040;
  assign n26685 = pi3283 & ~pi9040;
  assign n26686 = ~n26684 & ~n26685;
  assign n26687 = ~pi0387 & ~n26686;
  assign n26688 = pi0387 & ~n26684;
  assign n26689 = ~n26685 & n26688;
  assign n26690 = ~n26687 & ~n26689;
  assign n26691 = pi3417 & pi9040;
  assign n26692 = pi3313 & ~pi9040;
  assign n26693 = ~n26691 & ~n26692;
  assign n26694 = ~pi0397 & ~n26693;
  assign n26695 = pi0397 & n26693;
  assign n26696 = ~n26694 & ~n26695;
  assign n26697 = pi3284 & pi9040;
  assign n26698 = pi3401 & ~pi9040;
  assign n26699 = ~n26697 & ~n26698;
  assign n26700 = ~pi0391 & ~n26699;
  assign n26701 = pi0391 & n26699;
  assign n26702 = ~n26700 & ~n26701;
  assign n26703 = n26696 & ~n26702;
  assign n26704 = ~n26690 & n26703;
  assign n26705 = pi3339 & pi9040;
  assign n26706 = pi3285 & ~pi9040;
  assign n26707 = ~n26705 & ~n26706;
  assign n26708 = ~pi0383 & ~n26707;
  assign n26709 = pi0383 & ~n26705;
  assign n26710 = ~n26706 & n26709;
  assign n26711 = ~n26708 & ~n26710;
  assign n26712 = n26702 & ~n26711;
  assign n26713 = n26696 & n26712;
  assign n26714 = n26690 & n26713;
  assign n26715 = n26702 & n26711;
  assign n26716 = ~n26690 & n26715;
  assign n26717 = ~n26714 & ~n26716;
  assign n26718 = ~n26704 & n26717;
  assign n26719 = n26683 & ~n26718;
  assign n26720 = ~n26690 & ~n26696;
  assign n26721 = ~n26711 & n26720;
  assign n26722 = ~n26702 & ~n26711;
  assign n26723 = n26696 & n26722;
  assign n26724 = n26690 & n26723;
  assign n26725 = ~n26721 & ~n26724;
  assign n26726 = ~n26696 & n26712;
  assign n26727 = n26696 & n26715;
  assign n26728 = ~n26726 & ~n26727;
  assign n26729 = n26725 & n26728;
  assign n26730 = ~n26676 & ~n26729;
  assign n26731 = ~n26702 & n26711;
  assign n26732 = ~n26696 & n26731;
  assign n26733 = n26690 & n26732;
  assign n26734 = ~n26730 & ~n26733;
  assign n26735 = ~n26682 & ~n26734;
  assign n26736 = ~n26719 & ~n26735;
  assign n26737 = ~n26676 & ~n26690;
  assign n26738 = n26696 & n26737;
  assign n26739 = n26711 & n26738;
  assign n26740 = ~n26690 & n26726;
  assign n26741 = ~n26739 & ~n26740;
  assign n26742 = ~n26696 & n26722;
  assign n26743 = ~n26715 & ~n26722;
  assign n26744 = n26690 & ~n26743;
  assign n26745 = ~n26742 & ~n26744;
  assign n26746 = n26676 & ~n26745;
  assign n26747 = n26696 & n26731;
  assign n26748 = ~n26704 & ~n26747;
  assign n26749 = ~n26714 & n26748;
  assign n26750 = ~n26676 & ~n26749;
  assign n26751 = ~n26746 & ~n26750;
  assign n26752 = n26676 & ~n26690;
  assign n26753 = n26712 & n26752;
  assign n26754 = n26690 & n26742;
  assign n26755 = ~n26696 & n26702;
  assign n26756 = n26711 & n26755;
  assign n26757 = n26690 & n26756;
  assign n26758 = ~n26754 & ~n26757;
  assign n26759 = n26711 & n26720;
  assign n26760 = ~n26702 & n26759;
  assign n26761 = n26758 & ~n26760;
  assign n26762 = ~n26753 & n26761;
  assign n26763 = n26751 & n26762;
  assign n26764 = n26682 & ~n26763;
  assign n26765 = n26741 & ~n26764;
  assign n26766 = n26736 & n26765;
  assign n26767 = pi0422 & ~n26766;
  assign n26768 = ~pi0422 & n26741;
  assign n26769 = n26736 & n26768;
  assign n26770 = ~n26764 & n26769;
  assign po0442 = n26767 | n26770;
  assign n26772 = n26690 & n26703;
  assign n26773 = ~n26727 & ~n26772;
  assign n26774 = ~n26740 & n26773;
  assign n26775 = ~n26676 & ~n26774;
  assign n26776 = ~n26690 & n26711;
  assign n26777 = n26755 & n26776;
  assign n26778 = ~n26690 & n26747;
  assign n26779 = ~n26696 & ~n26702;
  assign n26780 = ~n26712 & ~n26779;
  assign n26781 = n26690 & ~n26780;
  assign n26782 = ~n26778 & ~n26781;
  assign n26783 = ~n26777 & n26782;
  assign n26784 = n26676 & ~n26783;
  assign n26785 = ~n26775 & ~n26784;
  assign n26786 = n26682 & ~n26785;
  assign n26787 = ~n26702 & n26737;
  assign n26788 = ~n26690 & n26696;
  assign n26789 = n26702 & n26788;
  assign n26790 = ~n26772 & ~n26789;
  assign n26791 = n26676 & ~n26790;
  assign n26792 = ~n26753 & ~n26791;
  assign n26793 = ~n26690 & n26713;
  assign n26794 = ~n26757 & ~n26793;
  assign n26795 = ~n26676 & n26690;
  assign n26796 = n26755 & n26795;
  assign n26797 = ~n26676 & n26732;
  assign n26798 = ~n26796 & ~n26797;
  assign n26799 = n26794 & n26798;
  assign n26800 = n26792 & n26799;
  assign n26801 = ~n26787 & n26800;
  assign n26802 = ~n26682 & ~n26801;
  assign n26803 = n26742 & n26752;
  assign n26804 = n26696 & n26753;
  assign n26805 = ~n26803 & ~n26804;
  assign n26806 = ~n26676 & n26760;
  assign n26807 = n26805 & ~n26806;
  assign n26808 = n26690 & n26715;
  assign n26809 = ~n26690 & n26723;
  assign n26810 = ~n26808 & ~n26809;
  assign n26811 = ~n26676 & ~n26810;
  assign n26812 = n26807 & ~n26811;
  assign n26813 = ~n26802 & n26812;
  assign n26814 = ~n26786 & n26813;
  assign n26815 = ~pi0420 & ~n26814;
  assign n26816 = pi0420 & n26814;
  assign po0445 = n26815 | n26816;
  assign n26818 = pi3293 & pi9040;
  assign n26819 = pi3342 & ~pi9040;
  assign n26820 = ~n26818 & ~n26819;
  assign n26821 = ~pi0389 & ~n26820;
  assign n26822 = pi0389 & n26820;
  assign n26823 = ~n26821 & ~n26822;
  assign n26824 = pi3340 & pi9040;
  assign n26825 = pi3293 & ~pi9040;
  assign n26826 = ~n26824 & ~n26825;
  assign n26827 = ~pi0382 & n26826;
  assign n26828 = pi0382 & ~n26826;
  assign n26829 = ~n26827 & ~n26828;
  assign n26830 = pi3303 & pi9040;
  assign n26831 = pi3340 & ~pi9040;
  assign n26832 = ~n26830 & ~n26831;
  assign n26833 = ~pi0400 & n26832;
  assign n26834 = pi0400 & ~n26832;
  assign n26835 = ~n26833 & ~n26834;
  assign n26836 = ~n26829 & n26835;
  assign n26837 = pi3401 & pi9040;
  assign n26838 = pi3339 & ~pi9040;
  assign n26839 = ~n26837 & ~n26838;
  assign n26840 = pi0384 & n26839;
  assign n26841 = ~pi0384 & ~n26839;
  assign n26842 = ~n26840 & ~n26841;
  assign n26843 = pi3288 & pi9040;
  assign n26844 = pi3291 & ~pi9040;
  assign n26845 = ~n26843 & ~n26844;
  assign n26846 = ~pi0406 & n26845;
  assign n26847 = pi0406 & ~n26845;
  assign n26848 = ~n26846 & ~n26847;
  assign n26849 = ~n26842 & n26848;
  assign n26850 = n26836 & n26849;
  assign n26851 = pi3313 & pi9040;
  assign n26852 = pi3284 & ~pi9040;
  assign n26853 = ~n26851 & ~n26852;
  assign n26854 = pi0383 & n26853;
  assign n26855 = ~pi0383 & ~n26853;
  assign n26856 = ~n26854 & ~n26855;
  assign n26857 = ~n26835 & ~n26856;
  assign n26858 = ~n26842 & ~n26848;
  assign n26859 = n26857 & n26858;
  assign n26860 = n26829 & ~n26835;
  assign n26861 = n26856 & n26860;
  assign n26862 = n26842 & ~n26856;
  assign n26863 = n26829 & n26862;
  assign n26864 = n26835 & n26863;
  assign n26865 = ~n26861 & ~n26864;
  assign n26866 = ~n26829 & ~n26835;
  assign n26867 = n26842 & n26866;
  assign n26868 = n26865 & ~n26867;
  assign n26869 = n26848 & ~n26868;
  assign n26870 = ~n26856 & n26860;
  assign n26871 = ~n26842 & n26870;
  assign n26872 = ~n26869 & ~n26871;
  assign n26873 = ~n26859 & n26872;
  assign n26874 = ~n26850 & n26873;
  assign n26875 = n26836 & n26856;
  assign n26876 = ~n26842 & n26875;
  assign n26877 = n26856 & n26866;
  assign n26878 = n26842 & n26877;
  assign n26879 = ~n26876 & ~n26878;
  assign n26880 = n26874 & n26879;
  assign n26881 = ~n26823 & ~n26880;
  assign n26882 = n26836 & ~n26856;
  assign n26883 = n26842 & n26882;
  assign n26884 = n26829 & n26835;
  assign n26885 = n26856 & n26884;
  assign n26886 = n26842 & n26885;
  assign n26887 = ~n26870 & ~n26886;
  assign n26888 = ~n26883 & n26887;
  assign n26889 = ~n26848 & ~n26888;
  assign n26890 = n26835 & n26856;
  assign n26891 = ~n26842 & n26890;
  assign n26892 = ~n26835 & n26856;
  assign n26893 = n26842 & n26892;
  assign n26894 = ~n26891 & ~n26893;
  assign n26895 = n26848 & ~n26894;
  assign n26896 = ~n26889 & ~n26895;
  assign n26897 = ~n26842 & ~n26856;
  assign n26898 = ~n26829 & n26897;
  assign n26899 = ~n26835 & n26898;
  assign n26900 = ~n26875 & ~n26899;
  assign n26901 = n26848 & ~n26900;
  assign n26902 = n26829 & ~n26856;
  assign n26903 = ~n26842 & n26902;
  assign n26904 = n26835 & n26903;
  assign n26905 = ~n26883 & ~n26904;
  assign n26906 = ~n26835 & n26862;
  assign n26907 = ~n26842 & n26877;
  assign n26908 = ~n26906 & ~n26907;
  assign n26909 = ~n26848 & ~n26908;
  assign n26910 = n26905 & ~n26909;
  assign n26911 = ~n26901 & n26910;
  assign n26912 = n26823 & ~n26911;
  assign n26913 = ~n26848 & n26902;
  assign n26914 = ~n26842 & n26913;
  assign n26915 = ~n26912 & ~n26914;
  assign n26916 = n26896 & n26915;
  assign n26917 = ~n26881 & n26916;
  assign n26918 = ~pi0435 & ~n26917;
  assign n26919 = pi0435 & n26917;
  assign po0452 = n26918 | n26919;
  assign n26921 = ~n26835 & n26863;
  assign n26922 = ~n26892 & ~n26904;
  assign n26923 = ~n26848 & ~n26922;
  assign n26924 = ~n26921 & ~n26923;
  assign n26925 = ~n26899 & n26924;
  assign n26926 = n26842 & n26848;
  assign n26927 = n26882 & n26926;
  assign n26928 = ~n26876 & ~n26927;
  assign n26929 = ~n26886 & n26928;
  assign n26930 = n26925 & n26929;
  assign n26931 = n26823 & ~n26930;
  assign n26932 = ~n26856 & n26866;
  assign n26933 = n26842 & n26932;
  assign n26934 = ~n26864 & ~n26933;
  assign n26935 = ~n26842 & n26885;
  assign n26936 = ~n26871 & ~n26935;
  assign n26937 = ~n26848 & n26882;
  assign n26938 = n26842 & n26875;
  assign n26939 = ~n26937 & ~n26938;
  assign n26940 = ~n26829 & n26856;
  assign n26941 = ~n26835 & n26842;
  assign n26942 = ~n26940 & ~n26941;
  assign n26943 = ~n26902 & n26942;
  assign n26944 = n26848 & ~n26943;
  assign n26945 = n26939 & ~n26944;
  assign n26946 = n26936 & n26945;
  assign n26947 = n26934 & n26946;
  assign n26948 = ~n26823 & ~n26947;
  assign n26949 = ~n26931 & ~n26948;
  assign n26950 = pi0430 & ~n26949;
  assign n26951 = ~pi0430 & ~n26931;
  assign n26952 = ~n26948 & n26951;
  assign po0453 = n26950 | n26952;
  assign n26954 = ~n26742 & ~n26747;
  assign n26955 = n26676 & ~n26954;
  assign n26956 = n26690 & n26727;
  assign n26957 = ~n26955 & ~n26956;
  assign n26958 = n26690 & n26702;
  assign n26959 = ~n26755 & ~n26958;
  assign n26960 = ~n26723 & n26959;
  assign n26961 = ~n26676 & ~n26960;
  assign n26962 = n26957 & ~n26961;
  assign n26963 = ~n26682 & ~n26962;
  assign n26964 = ~n26690 & n26756;
  assign n26965 = n26676 & n26964;
  assign n26966 = ~n26804 & ~n26965;
  assign n26967 = ~n26806 & n26966;
  assign n26968 = ~n26676 & n26702;
  assign n26969 = n26788 & n26968;
  assign n26970 = n26690 & n26747;
  assign n26971 = n26676 & n26755;
  assign n26972 = ~n26970 & ~n26971;
  assign n26973 = ~n26754 & n26972;
  assign n26974 = ~n26969 & n26973;
  assign n26975 = ~n26711 & n26788;
  assign n26976 = ~n26760 & ~n26975;
  assign n26977 = n26974 & n26976;
  assign n26978 = ~n26797 & n26977;
  assign n26979 = n26682 & ~n26978;
  assign n26980 = n26967 & ~n26979;
  assign n26981 = ~n26963 & n26980;
  assign n26982 = ~pi0433 & ~n26981;
  assign n26983 = pi0433 & n26967;
  assign n26984 = ~n26963 & n26983;
  assign n26985 = ~n26979 & n26984;
  assign po0454 = n26982 | n26985;
  assign n26987 = pi3320 & pi9040;
  assign n26988 = pi3341 & ~pi9040;
  assign n26989 = ~n26987 & ~n26988;
  assign n26990 = pi0404 & n26989;
  assign n26991 = ~pi0404 & ~n26989;
  assign n26992 = ~n26990 & ~n26991;
  assign n26993 = pi3276 & pi9040;
  assign n26994 = pi3380 & ~pi9040;
  assign n26995 = ~n26993 & ~n26994;
  assign n26996 = ~pi0405 & n26995;
  assign n26997 = pi0405 & ~n26995;
  assign n26998 = ~n26996 & ~n26997;
  assign n26999 = pi3364 & pi9040;
  assign n27000 = pi3278 & ~pi9040;
  assign n27001 = ~n26999 & ~n27000;
  assign n27002 = ~pi0415 & n27001;
  assign n27003 = pi0415 & ~n27001;
  assign n27004 = ~n27002 & ~n27003;
  assign n27005 = pi3317 & pi9040;
  assign n27006 = pi3364 & ~pi9040;
  assign n27007 = ~n27005 & ~n27006;
  assign n27008 = ~pi0376 & n27007;
  assign n27009 = pi0376 & ~n27007;
  assign n27010 = ~n27008 & ~n27009;
  assign n27011 = n27004 & ~n27010;
  assign n27012 = pi3318 & pi9040;
  assign n27013 = pi3414 & ~pi9040;
  assign n27014 = ~n27012 & ~n27013;
  assign n27015 = pi0392 & n27014;
  assign n27016 = ~pi0392 & ~n27014;
  assign n27017 = ~n27015 & ~n27016;
  assign n27018 = pi3319 & pi9040;
  assign n27019 = pi3317 & ~pi9040;
  assign n27020 = ~n27018 & ~n27019;
  assign n27021 = ~pi0407 & n27020;
  assign n27022 = pi0407 & ~n27020;
  assign n27023 = ~n27021 & ~n27022;
  assign n27024 = n27017 & ~n27023;
  assign n27025 = n27011 & n27024;
  assign n27026 = ~n26998 & n27025;
  assign n27027 = ~n27017 & ~n27023;
  assign n27028 = ~n27004 & ~n27010;
  assign n27029 = n27027 & n27028;
  assign n27030 = n27004 & n27010;
  assign n27031 = ~n26998 & n27030;
  assign n27032 = ~n27017 & n27031;
  assign n27033 = ~n27004 & n27010;
  assign n27034 = ~n26998 & n27033;
  assign n27035 = ~n27023 & n27034;
  assign n27036 = n27017 & n27035;
  assign n27037 = ~n27032 & ~n27036;
  assign n27038 = ~n27029 & n27037;
  assign n27039 = ~n27026 & n27038;
  assign n27040 = n26998 & ~n27017;
  assign n27041 = ~n27010 & n27040;
  assign n27042 = ~n27004 & n27041;
  assign n27043 = n27039 & ~n27042;
  assign n27044 = ~n26992 & ~n27043;
  assign n27045 = n26998 & n27010;
  assign n27046 = ~n27004 & n27045;
  assign n27047 = n27017 & n27023;
  assign n27048 = n27046 & n27047;
  assign n27049 = ~n26998 & ~n27017;
  assign n27050 = n27004 & n27049;
  assign n27051 = ~n27017 & n27030;
  assign n27052 = ~n27050 & ~n27051;
  assign n27053 = n27023 & ~n27052;
  assign n27054 = ~n27048 & ~n27053;
  assign n27055 = ~n26992 & ~n27054;
  assign n27056 = n27010 & n27049;
  assign n27057 = ~n26998 & ~n27004;
  assign n27058 = ~n27010 & n27057;
  assign n27059 = n27017 & n27058;
  assign n27060 = ~n27056 & ~n27059;
  assign n27061 = n26998 & n27011;
  assign n27062 = n27017 & n27061;
  assign n27063 = n27060 & ~n27062;
  assign n27064 = n27023 & ~n27063;
  assign n27065 = ~n27055 & ~n27064;
  assign n27066 = ~n27044 & n27065;
  assign n27067 = n26998 & n27017;
  assign n27068 = ~n27023 & n27067;
  assign n27069 = n27030 & n27068;
  assign n27070 = n26998 & ~n27004;
  assign n27071 = n27027 & n27070;
  assign n27072 = n27023 & n27057;
  assign n27073 = n27004 & n27017;
  assign n27074 = n26998 & n27073;
  assign n27075 = ~n27061 & ~n27074;
  assign n27076 = ~n27072 & n27075;
  assign n27077 = ~n27017 & n27046;
  assign n27078 = n27076 & ~n27077;
  assign n27079 = n27011 & ~n27023;
  assign n27080 = ~n27017 & n27079;
  assign n27081 = n26998 & ~n27010;
  assign n27082 = n27017 & n27030;
  assign n27083 = ~n27081 & ~n27082;
  assign n27084 = ~n27023 & ~n27083;
  assign n27085 = ~n27080 & ~n27084;
  assign n27086 = n27078 & n27085;
  assign n27087 = n26992 & ~n27086;
  assign n27088 = ~n27071 & ~n27087;
  assign n27089 = ~n27069 & n27088;
  assign n27090 = n27066 & n27089;
  assign n27091 = pi0418 & n27090;
  assign n27092 = ~pi0418 & ~n27090;
  assign po0455 = n27091 | n27092;
  assign n27094 = pi3414 & pi9040;
  assign n27095 = pi3320 & ~pi9040;
  assign n27096 = ~n27094 & ~n27095;
  assign n27097 = ~pi0410 & ~n27096;
  assign n27098 = pi0410 & n27096;
  assign n27099 = ~n27097 & ~n27098;
  assign n27100 = pi3300 & pi9040;
  assign n27101 = pi3299 & ~pi9040;
  assign n27102 = ~n27100 & ~n27101;
  assign n27103 = ~pi0394 & n27102;
  assign n27104 = pi0394 & ~n27102;
  assign n27105 = ~n27103 & ~n27104;
  assign n27106 = pi3301 & pi9040;
  assign n27107 = pi3354 & ~pi9040;
  assign n27108 = ~n27106 & ~n27107;
  assign n27109 = ~pi0409 & ~n27108;
  assign n27110 = pi0409 & n27108;
  assign n27111 = ~n27109 & ~n27110;
  assign n27112 = pi3354 & pi9040;
  assign n27113 = pi3305 & ~pi9040;
  assign n27114 = ~n27112 & ~n27113;
  assign n27115 = ~pi0395 & ~n27114;
  assign n27116 = pi0395 & n27114;
  assign n27117 = ~n27115 & ~n27116;
  assign n27118 = pi3338 & pi9040;
  assign n27119 = pi3318 & ~pi9040;
  assign n27120 = ~n27118 & ~n27119;
  assign n27121 = ~pi0403 & n27120;
  assign n27122 = pi0403 & ~n27120;
  assign n27123 = ~n27121 & ~n27122;
  assign n27124 = ~n27117 & n27123;
  assign n27125 = ~n27111 & n27124;
  assign n27126 = n27105 & n27125;
  assign n27127 = ~n27105 & ~n27111;
  assign n27128 = n27123 & n27127;
  assign n27129 = n27117 & n27128;
  assign n27130 = ~n27126 & ~n27129;
  assign n27131 = n27099 & ~n27130;
  assign n27132 = ~n27117 & ~n27123;
  assign n27133 = n27111 & n27132;
  assign n27134 = n27105 & n27133;
  assign n27135 = ~n27099 & n27134;
  assign n27136 = pi3274 & pi9040;
  assign n27137 = pi3400 & ~pi9040;
  assign n27138 = ~n27136 & ~n27137;
  assign n27139 = ~pi0408 & ~n27138;
  assign n27140 = pi0408 & ~n27136;
  assign n27141 = ~n27137 & n27140;
  assign n27142 = ~n27139 & ~n27141;
  assign n27143 = n27117 & n27123;
  assign n27144 = n27111 & n27143;
  assign n27145 = n27099 & n27144;
  assign n27146 = ~n27134 & ~n27145;
  assign n27147 = n27105 & n27117;
  assign n27148 = ~n27111 & n27147;
  assign n27149 = n27105 & n27111;
  assign n27150 = ~n27117 & n27149;
  assign n27151 = ~n27148 & ~n27150;
  assign n27152 = ~n27099 & ~n27151;
  assign n27153 = ~n27099 & ~n27105;
  assign n27154 = n27124 & n27153;
  assign n27155 = ~n27111 & n27154;
  assign n27156 = ~n27105 & n27111;
  assign n27157 = ~n27123 & n27156;
  assign n27158 = n27117 & n27157;
  assign n27159 = ~n27111 & n27132;
  assign n27160 = n27099 & n27159;
  assign n27161 = ~n27158 & ~n27160;
  assign n27162 = ~n27155 & n27161;
  assign n27163 = ~n27152 & n27162;
  assign n27164 = n27146 & n27163;
  assign n27165 = n27142 & ~n27164;
  assign n27166 = n27105 & n27145;
  assign n27167 = ~n27165 & ~n27166;
  assign n27168 = ~n27135 & n27167;
  assign n27169 = ~n27131 & n27168;
  assign n27170 = n27099 & ~n27105;
  assign n27171 = n27111 & ~n27117;
  assign n27172 = n27170 & n27171;
  assign n27173 = n27099 & n27125;
  assign n27174 = ~n27172 & ~n27173;
  assign n27175 = n27117 & ~n27123;
  assign n27176 = n27111 & n27175;
  assign n27177 = n27099 & n27176;
  assign n27178 = ~n27111 & n27175;
  assign n27179 = n27105 & n27178;
  assign n27180 = ~n27177 & ~n27179;
  assign n27181 = n27111 & n27124;
  assign n27182 = ~n27105 & n27181;
  assign n27183 = ~n27126 & ~n27182;
  assign n27184 = ~n27105 & n27143;
  assign n27185 = ~n27111 & ~n27123;
  assign n27186 = ~n27184 & ~n27185;
  assign n27187 = ~n27099 & ~n27186;
  assign n27188 = n27183 & ~n27187;
  assign n27189 = n27180 & n27188;
  assign n27190 = n27174 & n27189;
  assign n27191 = ~n27142 & ~n27190;
  assign n27192 = n27169 & ~n27191;
  assign n27193 = ~pi0429 & ~n27192;
  assign n27194 = pi0429 & n27169;
  assign n27195 = ~n27191 & n27194;
  assign po0456 = n27193 | n27195;
  assign n27197 = n27099 & n27132;
  assign n27198 = n27105 & n27197;
  assign n27199 = ~n27111 & n27143;
  assign n27200 = n27117 & n27127;
  assign n27201 = ~n27199 & ~n27200;
  assign n27202 = n27099 & ~n27201;
  assign n27203 = ~n27198 & ~n27202;
  assign n27204 = ~n27099 & n27105;
  assign n27205 = n27175 & n27204;
  assign n27206 = ~n27099 & n27125;
  assign n27207 = ~n27205 & ~n27206;
  assign n27208 = n27203 & n27207;
  assign n27209 = n27117 & n27149;
  assign n27210 = ~n27126 & ~n27209;
  assign n27211 = ~n27182 & n27210;
  assign n27212 = n27208 & n27211;
  assign n27213 = ~n27142 & ~n27212;
  assign n27214 = ~n27166 & ~n27172;
  assign n27215 = ~n27134 & ~n27199;
  assign n27216 = ~n27184 & n27215;
  assign n27217 = ~n27099 & ~n27216;
  assign n27218 = ~n27123 & n27127;
  assign n27219 = ~n27117 & n27218;
  assign n27220 = ~n27158 & ~n27219;
  assign n27221 = n27099 & n27105;
  assign n27222 = n27178 & n27221;
  assign n27223 = n27220 & ~n27222;
  assign n27224 = n27099 & n27181;
  assign n27225 = n27223 & ~n27224;
  assign n27226 = ~n27217 & n27225;
  assign n27227 = n27142 & ~n27226;
  assign n27228 = ~n27126 & n27220;
  assign n27229 = ~n27099 & ~n27228;
  assign n27230 = ~n27227 & ~n27229;
  assign n27231 = n27214 & n27230;
  assign n27232 = ~n27213 & n27231;
  assign n27233 = pi0436 & ~n27232;
  assign n27234 = ~pi0436 & n27232;
  assign po0457 = n27233 | n27234;
  assign n27236 = ~n26998 & n27004;
  assign n27237 = ~n27042 & ~n27236;
  assign n27238 = ~n27073 & n27237;
  assign n27239 = ~n27023 & ~n27238;
  assign n27240 = ~n27004 & n27047;
  assign n27241 = ~n26998 & n27017;
  assign n27242 = ~n27010 & n27241;
  assign n27243 = ~n27017 & n27034;
  assign n27244 = ~n27242 & ~n27243;
  assign n27245 = n26998 & n27004;
  assign n27246 = ~n27017 & n27023;
  assign n27247 = n27245 & n27246;
  assign n27248 = n27244 & ~n27247;
  assign n27249 = ~n27240 & n27248;
  assign n27250 = ~n27239 & n27249;
  assign n27251 = n26992 & ~n27250;
  assign n27252 = ~n26998 & n27011;
  assign n27253 = ~n27017 & n27252;
  assign n27254 = n27017 & n27031;
  assign n27255 = ~n27253 & ~n27254;
  assign n27256 = ~n27023 & ~n27255;
  assign n27257 = ~n27251 & ~n27256;
  assign n27258 = n27017 & n27034;
  assign n27259 = ~n27046 & ~n27058;
  assign n27260 = ~n27023 & ~n27259;
  assign n27261 = ~n27258 & ~n27260;
  assign n27262 = ~n27062 & n27261;
  assign n27263 = ~n26992 & ~n27262;
  assign n27264 = ~n27028 & ~n27030;
  assign n27265 = n26998 & ~n27264;
  assign n27266 = ~n27051 & ~n27265;
  assign n27267 = n27023 & ~n27266;
  assign n27268 = ~n26992 & n27267;
  assign n27269 = ~n27263 & ~n27268;
  assign n27270 = n27257 & n27269;
  assign n27271 = pi0419 & ~n27270;
  assign n27272 = ~pi0419 & n27257;
  assign n27273 = n27269 & n27272;
  assign po0458 = n27271 | n27273;
  assign n27275 = ~n26690 & ~n26702;
  assign n27276 = ~n26975 & ~n27275;
  assign n27277 = n26676 & ~n27276;
  assign n27278 = n26690 & n26696;
  assign n27279 = n26711 & n27278;
  assign n27280 = ~n27277 & ~n27279;
  assign n27281 = ~n26676 & n26715;
  assign n27282 = ~n26690 & n27281;
  assign n27283 = ~n26809 & ~n27282;
  assign n27284 = n27280 & n27283;
  assign n27285 = n26682 & ~n27284;
  assign n27286 = ~n26713 & ~n26757;
  assign n27287 = ~n26690 & n26731;
  assign n27288 = n27286 & ~n27287;
  assign n27289 = ~n26676 & ~n27288;
  assign n27290 = n26715 & n26752;
  assign n27291 = ~n26740 & ~n27290;
  assign n27292 = ~n27289 & n27291;
  assign n27293 = ~n26723 & ~n26733;
  assign n27294 = n26676 & ~n27293;
  assign n27295 = n27292 & ~n27294;
  assign n27296 = ~n26682 & ~n27295;
  assign n27297 = ~n27285 & ~n27296;
  assign n27298 = ~n26690 & n26722;
  assign n27299 = n26690 & ~n26728;
  assign n27300 = ~n27298 & ~n27299;
  assign n27301 = n26676 & ~n27300;
  assign n27302 = ~n26713 & n26954;
  assign n27303 = n26795 & ~n27302;
  assign n27304 = ~n27301 & ~n27303;
  assign n27305 = n27297 & n27304;
  assign n27306 = ~pi0424 & ~n27305;
  assign n27307 = pi0424 & n27304;
  assign n27308 = ~n27296 & n27307;
  assign n27309 = ~n27285 & n27308;
  assign po0459 = n27306 | n27309;
  assign n27311 = pi3337 & pi9040;
  assign n27312 = pi3288 & ~pi9040;
  assign n27313 = ~n27311 & ~n27312;
  assign n27314 = pi0391 & n27313;
  assign n27315 = ~pi0391 & ~n27313;
  assign n27316 = ~n27314 & ~n27315;
  assign n27317 = pi3280 & pi9040;
  assign n27318 = pi3417 & ~pi9040;
  assign n27319 = ~n27317 & ~n27318;
  assign n27320 = ~pi0414 & n27319;
  assign n27321 = pi0414 & ~n27319;
  assign n27322 = ~n27320 & ~n27321;
  assign n27323 = pi3355 & pi9040;
  assign n27324 = pi3286 & ~pi9040;
  assign n27325 = ~n27323 & ~n27324;
  assign n27326 = ~pi0403 & n27325;
  assign n27327 = pi0403 & ~n27325;
  assign n27328 = ~n27326 & ~n27327;
  assign n27329 = pi3335 & pi9040;
  assign n27330 = pi3289 & ~pi9040;
  assign n27331 = ~n27329 & ~n27330;
  assign n27332 = ~pi0408 & ~n27331;
  assign n27333 = pi0408 & ~n27329;
  assign n27334 = ~n27330 & n27333;
  assign n27335 = ~n27332 & ~n27334;
  assign n27336 = pi3352 & pi9040;
  assign n27337 = pi3321 & ~pi9040;
  assign n27338 = ~n27336 & ~n27337;
  assign n27339 = pi0397 & n27338;
  assign n27340 = ~pi0397 & ~n27338;
  assign n27341 = ~n27339 & ~n27340;
  assign n27342 = ~n27335 & ~n27341;
  assign n27343 = ~n27328 & n27342;
  assign n27344 = ~n27322 & n27343;
  assign n27345 = ~n27335 & n27341;
  assign n27346 = n27328 & n27345;
  assign n27347 = ~n27322 & n27346;
  assign n27348 = ~n27344 & ~n27347;
  assign n27349 = n27335 & n27341;
  assign n27350 = n27328 & n27349;
  assign n27351 = n27328 & n27342;
  assign n27352 = n27322 & n27351;
  assign n27353 = ~n27350 & ~n27352;
  assign n27354 = pi3291 & pi9040;
  assign n27355 = pi3334 & ~pi9040;
  assign n27356 = ~n27354 & ~n27355;
  assign n27357 = ~pi0396 & n27356;
  assign n27358 = pi0396 & ~n27356;
  assign n27359 = ~n27357 & ~n27358;
  assign n27360 = ~n27353 & ~n27359;
  assign n27361 = n27348 & ~n27360;
  assign n27362 = n27322 & n27359;
  assign n27363 = n27335 & n27362;
  assign n27364 = n27361 & ~n27363;
  assign n27365 = n27316 & ~n27364;
  assign n27366 = ~n27322 & n27335;
  assign n27367 = n27328 & n27366;
  assign n27368 = ~n27341 & n27367;
  assign n27369 = n27359 & n27368;
  assign n27370 = n27322 & ~n27359;
  assign n27371 = n27335 & ~n27341;
  assign n27372 = n27328 & n27371;
  assign n27373 = n27370 & n27372;
  assign n27374 = n27322 & ~n27328;
  assign n27375 = ~n27335 & n27374;
  assign n27376 = ~n27373 & ~n27375;
  assign n27377 = ~n27328 & n27345;
  assign n27378 = ~n27350 & ~n27377;
  assign n27379 = n27322 & n27345;
  assign n27380 = n27378 & ~n27379;
  assign n27381 = n27359 & ~n27380;
  assign n27382 = ~n27328 & ~n27341;
  assign n27383 = n27335 & n27382;
  assign n27384 = ~n27322 & n27383;
  assign n27385 = ~n27322 & n27351;
  assign n27386 = ~n27384 & ~n27385;
  assign n27387 = ~n27328 & n27349;
  assign n27388 = ~n27359 & n27387;
  assign n27389 = n27386 & ~n27388;
  assign n27390 = ~n27381 & n27389;
  assign n27391 = n27376 & n27390;
  assign n27392 = ~n27316 & ~n27391;
  assign n27393 = ~n27369 & ~n27392;
  assign n27394 = ~n27365 & n27393;
  assign n27395 = n27370 & n27377;
  assign n27396 = ~n27359 & n27382;
  assign n27397 = ~n27322 & n27396;
  assign n27398 = ~n27395 & ~n27397;
  assign n27399 = n27347 & ~n27359;
  assign n27400 = n27398 & ~n27399;
  assign n27401 = n27394 & n27400;
  assign n27402 = ~pi0427 & ~n27401;
  assign n27403 = pi0427 & n27400;
  assign n27404 = n27393 & n27403;
  assign n27405 = ~n27365 & n27404;
  assign po0460 = n27402 | n27405;
  assign n27407 = ~n27328 & ~n27335;
  assign n27408 = ~n27341 & n27407;
  assign n27409 = n27322 & n27408;
  assign n27410 = n27322 & n27387;
  assign n27411 = ~n27346 & ~n27410;
  assign n27412 = ~n27322 & n27382;
  assign n27413 = n27322 & n27372;
  assign n27414 = ~n27412 & ~n27413;
  assign n27415 = n27411 & n27414;
  assign n27416 = n27359 & ~n27415;
  assign n27417 = ~n27322 & n27349;
  assign n27418 = ~n27375 & ~n27417;
  assign n27419 = ~n27351 & n27418;
  assign n27420 = ~n27359 & ~n27419;
  assign n27421 = ~n27322 & n27328;
  assign n27422 = n27341 & n27421;
  assign n27423 = n27335 & n27422;
  assign n27424 = ~n27420 & ~n27423;
  assign n27425 = ~n27416 & n27424;
  assign n27426 = ~n27409 & n27425;
  assign n27427 = ~n27316 & ~n27426;
  assign n27428 = ~n27322 & n27359;
  assign n27429 = n27387 & n27428;
  assign n27430 = n27351 & n27359;
  assign n27431 = n27359 & n27377;
  assign n27432 = ~n27430 & ~n27431;
  assign n27433 = n27322 & ~n27432;
  assign n27434 = ~n27429 & ~n27433;
  assign n27435 = n27322 & n27383;
  assign n27436 = ~n27368 & ~n27435;
  assign n27437 = ~n27322 & n27345;
  assign n27438 = n27322 & n27349;
  assign n27439 = ~n27437 & ~n27438;
  assign n27440 = ~n27383 & n27439;
  assign n27441 = ~n27346 & n27440;
  assign n27442 = ~n27359 & ~n27441;
  assign n27443 = n27322 & n27350;
  assign n27444 = ~n27442 & ~n27443;
  assign n27445 = n27436 & n27444;
  assign n27446 = n27434 & n27445;
  assign n27447 = n27316 & ~n27446;
  assign n27448 = ~n27348 & n27359;
  assign n27449 = ~n27447 & ~n27448;
  assign n27450 = ~n27385 & ~n27435;
  assign n27451 = ~n27359 & ~n27450;
  assign n27452 = n27449 & ~n27451;
  assign n27453 = ~n27427 & n27452;
  assign n27454 = pi0437 & ~n27453;
  assign n27455 = ~pi0437 & n27453;
  assign po0461 = n27454 | n27455;
  assign n27457 = ~n26580 & n26587;
  assign n27458 = ~n26573 & n27457;
  assign n27459 = ~n26601 & n27458;
  assign n27460 = n26587 & n26616;
  assign n27461 = n26580 & ~n26593;
  assign n27462 = n26601 & n27461;
  assign n27463 = ~n26608 & ~n27462;
  assign n27464 = ~n27460 & n27463;
  assign n27465 = ~n27459 & n27464;
  assign n27466 = n26573 & n26604;
  assign n27467 = n27465 & ~n27466;
  assign n27468 = n26640 & ~n27467;
  assign n27469 = n26601 & n26610;
  assign n27470 = ~n26658 & ~n27469;
  assign n27471 = n26573 & ~n27470;
  assign n27472 = ~n26640 & n26642;
  assign n27473 = ~n26573 & n27472;
  assign n27474 = n26580 & n26601;
  assign n27475 = ~n26587 & n27474;
  assign n27476 = ~n27461 & ~n27475;
  assign n27477 = ~n26610 & n27476;
  assign n27478 = n26573 & ~n27477;
  assign n27479 = ~n26580 & n26627;
  assign n27480 = n26601 & n27479;
  assign n27481 = ~n27478 & ~n27480;
  assign n27482 = ~n26640 & ~n27481;
  assign n27483 = ~n27473 & ~n27482;
  assign n27484 = ~n27471 & n27483;
  assign n27485 = ~n26605 & ~n26608;
  assign n27486 = ~n26593 & ~n26601;
  assign n27487 = ~n26580 & n27486;
  assign n27488 = n26601 & n26657;
  assign n27489 = ~n27487 & ~n27488;
  assign n27490 = n27485 & n27489;
  assign n27491 = ~n26573 & ~n27490;
  assign n27492 = n27484 & ~n27491;
  assign n27493 = ~n27468 & n27492;
  assign n27494 = ~pi0445 & ~n27493;
  assign n27495 = pi0445 & n27484;
  assign n27496 = ~n27468 & n27495;
  assign n27497 = ~n27491 & n27496;
  assign po0462 = n27494 | n27497;
  assign n27499 = ~n26628 & ~n27487;
  assign n27500 = n26573 & ~n27499;
  assign n27501 = ~n26573 & n26601;
  assign n27502 = ~n26593 & n27501;
  assign n27503 = n26587 & n27502;
  assign n27504 = n26609 & n26643;
  assign n27505 = ~n27503 & ~n27504;
  assign n27506 = ~n27500 & n27505;
  assign n27507 = n26593 & n26607;
  assign n27508 = n26601 & n26631;
  assign n27509 = ~n27507 & ~n27508;
  assign n27510 = ~n26605 & n27509;
  assign n27511 = ~n26573 & n26580;
  assign n27512 = n26603 & n27511;
  assign n27513 = ~n26617 & ~n27512;
  assign n27514 = n27510 & n27513;
  assign n27515 = n27506 & n27514;
  assign n27516 = ~n26640 & ~n27515;
  assign n27517 = ~n26604 & ~n26628;
  assign n27518 = ~n26601 & ~n27517;
  assign n27519 = n26587 & n26646;
  assign n27520 = ~n26657 & ~n27519;
  assign n27521 = ~n26601 & n27461;
  assign n27522 = n27520 & ~n27521;
  assign n27523 = n26573 & ~n27522;
  assign n27524 = n26601 & n26627;
  assign n27525 = ~n27460 & ~n27524;
  assign n27526 = ~n26573 & ~n27525;
  assign n27527 = ~n27469 & ~n27526;
  assign n27528 = ~n27523 & n27527;
  assign n27529 = ~n27518 & n27528;
  assign n27530 = n26640 & ~n27529;
  assign n27531 = n26573 & n26647;
  assign n27532 = ~n27530 & ~n27531;
  assign n27533 = n26622 & n27501;
  assign n27534 = ~n26593 & n27533;
  assign n27535 = n27532 & ~n27534;
  assign n27536 = ~n27516 & n27535;
  assign n27537 = ~pi0447 & ~n27536;
  assign n27538 = pi0447 & n27532;
  assign n27539 = ~n27516 & n27538;
  assign n27540 = ~n27534 & n27539;
  assign po0463 = n27537 | n27540;
  assign n27542 = ~n27105 & n27133;
  assign n27543 = ~n27105 & n27175;
  assign n27544 = n27105 & n27159;
  assign n27545 = ~n27543 & ~n27544;
  assign n27546 = ~n27099 & ~n27545;
  assign n27547 = ~n27542 & ~n27546;
  assign n27548 = ~n27105 & n27197;
  assign n27549 = ~n27173 & ~n27548;
  assign n27550 = n27547 & n27549;
  assign n27551 = ~n27105 & n27144;
  assign n27552 = n27105 & n27181;
  assign n27553 = ~n27551 & ~n27552;
  assign n27554 = n27550 & n27553;
  assign n27555 = n27142 & ~n27554;
  assign n27556 = ~n27099 & ~n27142;
  assign n27557 = ~n27117 & n27127;
  assign n27558 = ~n27111 & n27123;
  assign n27559 = ~n27557 & ~n27558;
  assign n27560 = n27556 & ~n27559;
  assign n27561 = ~n27134 & ~n27148;
  assign n27562 = n27111 & n27170;
  assign n27563 = ~n27132 & n27562;
  assign n27564 = ~n27145 & ~n27563;
  assign n27565 = n27561 & n27564;
  assign n27566 = ~n27142 & ~n27565;
  assign n27567 = n27199 & n27204;
  assign n27568 = n27105 & n27176;
  assign n27569 = ~n27552 & ~n27568;
  assign n27570 = ~n27099 & ~n27569;
  assign n27571 = ~n27567 & ~n27570;
  assign n27572 = n27133 & n27221;
  assign n27573 = n27571 & ~n27572;
  assign n27574 = ~n27566 & n27573;
  assign n27575 = ~n27560 & n27574;
  assign n27576 = ~n27555 & n27575;
  assign n27577 = ~n27222 & n27576;
  assign n27578 = ~pi0432 & ~n27577;
  assign n27579 = pi0432 & ~n27222;
  assign n27580 = n27575 & n27579;
  assign n27581 = ~n27555 & n27580;
  assign po0464 = n27578 | n27581;
  assign n27583 = pi3281 & pi9040;
  assign n27584 = pi3275 & ~pi9040;
  assign n27585 = ~n27583 & ~n27584;
  assign n27586 = pi0412 & n27585;
  assign n27587 = ~pi0412 & ~n27585;
  assign n27588 = ~n27586 & ~n27587;
  assign n27589 = pi3297 & pi9040;
  assign n27590 = pi3386 & ~pi9040;
  assign n27591 = ~n27589 & ~n27590;
  assign n27592 = pi0404 & n27591;
  assign n27593 = ~pi0404 & ~n27591;
  assign n27594 = ~n27592 & ~n27593;
  assign n27595 = pi3341 & pi9040;
  assign n27596 = pi3312 & ~pi9040;
  assign n27597 = ~n27595 & ~n27596;
  assign n27598 = pi0413 & n27597;
  assign n27599 = ~pi0413 & ~n27597;
  assign n27600 = ~n27598 & ~n27599;
  assign n27601 = n27594 & ~n27600;
  assign n27602 = pi3275 & pi9040;
  assign n27603 = pi3319 & ~pi9040;
  assign n27604 = ~n27602 & ~n27603;
  assign n27605 = pi0399 & n27604;
  assign n27606 = ~pi0399 & ~n27604;
  assign n27607 = ~n27605 & ~n27606;
  assign n27608 = pi3304 & pi9040;
  assign n27609 = pi3306 & ~pi9040;
  assign n27610 = ~n27608 & ~n27609;
  assign n27611 = pi0376 & n27610;
  assign n27612 = ~pi0376 & ~n27610;
  assign n27613 = ~n27611 & ~n27612;
  assign n27614 = n27607 & n27613;
  assign n27615 = n27601 & n27614;
  assign n27616 = n27607 & ~n27613;
  assign n27617 = ~n27594 & n27616;
  assign n27618 = ~n27615 & ~n27617;
  assign n27619 = ~n27588 & ~n27618;
  assign n27620 = pi3316 & pi9040;
  assign n27621 = pi3338 & ~pi9040;
  assign n27622 = ~n27620 & ~n27621;
  assign n27623 = ~pi0386 & ~n27622;
  assign n27624 = pi0386 & n27622;
  assign n27625 = ~n27623 & ~n27624;
  assign n27626 = n27588 & ~n27607;
  assign n27627 = n27594 & n27626;
  assign n27628 = n27601 & ~n27613;
  assign n27629 = n27594 & n27600;
  assign n27630 = n27613 & n27629;
  assign n27631 = ~n27628 & ~n27630;
  assign n27632 = ~n27594 & ~n27600;
  assign n27633 = n27613 & n27632;
  assign n27634 = n27607 & n27633;
  assign n27635 = n27631 & ~n27634;
  assign n27636 = n27588 & ~n27635;
  assign n27637 = ~n27627 & ~n27636;
  assign n27638 = ~n27594 & n27600;
  assign n27639 = ~n27613 & n27638;
  assign n27640 = n27607 & n27639;
  assign n27641 = n27637 & ~n27640;
  assign n27642 = ~n27607 & n27632;
  assign n27643 = ~n27594 & n27613;
  assign n27644 = n27600 & n27643;
  assign n27645 = ~n27642 & ~n27644;
  assign n27646 = ~n27588 & ~n27645;
  assign n27647 = ~n27613 & n27629;
  assign n27648 = ~n27607 & n27647;
  assign n27649 = ~n27646 & ~n27648;
  assign n27650 = n27641 & n27649;
  assign n27651 = n27625 & ~n27650;
  assign n27652 = ~n27619 & ~n27651;
  assign n27653 = n27588 & ~n27625;
  assign n27654 = ~n27645 & n27653;
  assign n27655 = ~n27613 & n27632;
  assign n27656 = ~n27647 & ~n27655;
  assign n27657 = n27607 & ~n27656;
  assign n27658 = ~n27615 & ~n27657;
  assign n27659 = ~n27625 & ~n27658;
  assign n27660 = ~n27654 & ~n27659;
  assign n27661 = ~n27588 & ~n27625;
  assign n27662 = n27601 & ~n27607;
  assign n27663 = ~n27639 & ~n27662;
  assign n27664 = n27594 & n27613;
  assign n27665 = n27663 & ~n27664;
  assign n27666 = n27661 & ~n27665;
  assign n27667 = n27660 & ~n27666;
  assign n27668 = n27652 & n27667;
  assign n27669 = ~pi0416 & ~n27668;
  assign n27670 = pi0416 & n27660;
  assign n27671 = n27652 & n27670;
  assign n27672 = ~n27666 & n27671;
  assign po0465 = n27669 | n27672;
  assign n27674 = n27341 & n27374;
  assign n27675 = ~n27350 & ~n27375;
  assign n27676 = n27359 & ~n27675;
  assign n27677 = ~n27674 & ~n27676;
  assign n27678 = n27328 & ~n27335;
  assign n27679 = n27328 & ~n27341;
  assign n27680 = n27322 & n27679;
  assign n27681 = ~n27322 & n27342;
  assign n27682 = ~n27680 & ~n27681;
  assign n27683 = ~n27678 & n27682;
  assign n27684 = ~n27387 & n27683;
  assign n27685 = ~n27359 & ~n27684;
  assign n27686 = n27677 & ~n27685;
  assign n27687 = ~n27384 & n27686;
  assign n27688 = n27316 & ~n27687;
  assign n27689 = n27322 & n27346;
  assign n27690 = n27386 & ~n27689;
  assign n27691 = ~n27359 & ~n27690;
  assign n27692 = ~n27688 & ~n27691;
  assign n27693 = n27328 & n27335;
  assign n27694 = n27359 & n27693;
  assign n27695 = ~n27322 & n27694;
  assign n27696 = n27370 & n27382;
  assign n27697 = ~n27322 & n27377;
  assign n27698 = ~n27696 & ~n27697;
  assign n27699 = ~n27322 & n27407;
  assign n27700 = ~n27372 & ~n27699;
  assign n27701 = n27359 & ~n27700;
  assign n27702 = n27359 & n27678;
  assign n27703 = n27322 & n27702;
  assign n27704 = ~n27701 & ~n27703;
  assign n27705 = n27698 & n27704;
  assign n27706 = ~n27316 & ~n27705;
  assign n27707 = ~n27695 & ~n27706;
  assign n27708 = ~n27410 & n27707;
  assign n27709 = n27692 & n27708;
  assign n27710 = ~pi0431 & ~n27709;
  assign n27711 = ~n27410 & ~n27688;
  assign n27712 = ~n27691 & n27711;
  assign n27713 = n27707 & n27712;
  assign n27714 = pi0431 & n27713;
  assign po0466 = n27710 | n27714;
  assign n27716 = ~n27017 & n27061;
  assign n27717 = ~n27243 & ~n27716;
  assign n27718 = n27023 & ~n27717;
  assign n27719 = n27047 & n27058;
  assign n27720 = ~n27718 & ~n27719;
  assign n27721 = ~n27071 & n27720;
  assign n27722 = ~n26998 & ~n27023;
  assign n27723 = n27010 & n27722;
  assign n27724 = n27004 & n27723;
  assign n27725 = ~n27017 & n27724;
  assign n27726 = ~n27023 & n27252;
  assign n27727 = ~n27042 & ~n27069;
  assign n27728 = ~n27036 & n27727;
  assign n27729 = ~n27726 & n27728;
  assign n27730 = n26992 & ~n27729;
  assign n27731 = ~n27004 & n27017;
  assign n27732 = n26998 & n27731;
  assign n27733 = n27010 & n27732;
  assign n27734 = ~n27031 & ~n27733;
  assign n27735 = ~n27061 & n27734;
  assign n27736 = n27023 & ~n27735;
  assign n27737 = n26992 & n27736;
  assign n27738 = n27017 & n27079;
  assign n27739 = ~n27724 & ~n27738;
  assign n27740 = ~n27242 & n27739;
  assign n27741 = n27010 & n27040;
  assign n27742 = n27017 & n27028;
  assign n27743 = ~n27057 & ~n27742;
  assign n27744 = n27023 & ~n27743;
  assign n27745 = ~n27741 & ~n27744;
  assign n27746 = n27740 & n27745;
  assign n27747 = ~n26992 & ~n27746;
  assign n27748 = ~n27737 & ~n27747;
  assign n27749 = ~n27730 & n27748;
  assign n27750 = ~n27725 & n27749;
  assign n27751 = n27721 & n27750;
  assign n27752 = pi0426 & ~n27751;
  assign n27753 = ~pi0426 & n27721;
  assign n27754 = n27750 & n27753;
  assign po0467 = n27752 | n27754;
  assign n27756 = pi3312 & pi9040;
  assign n27757 = pi3304 & ~pi9040;
  assign n27758 = ~n27756 & ~n27757;
  assign n27759 = pi0413 & n27758;
  assign n27760 = ~pi0413 & ~n27758;
  assign n27761 = ~n27759 & ~n27760;
  assign n27762 = pi3299 & pi9040;
  assign n27763 = pi3276 & ~pi9040;
  assign n27764 = ~n27762 & ~n27763;
  assign n27765 = pi0409 & n27764;
  assign n27766 = ~pi0409 & ~n27764;
  assign n27767 = ~n27765 & ~n27766;
  assign n27768 = pi3278 & pi9040;
  assign n27769 = pi3279 & ~pi9040;
  assign n27770 = ~n27768 & ~n27769;
  assign n27771 = ~pi0386 & n27770;
  assign n27772 = pi0386 & ~n27770;
  assign n27773 = ~n27771 & ~n27772;
  assign n27774 = ~n27767 & ~n27773;
  assign n27775 = ~n27761 & n27774;
  assign n27776 = n27767 & ~n27773;
  assign n27777 = n27761 & n27776;
  assign n27778 = ~n27775 & ~n27777;
  assign n27779 = pi3386 & pi9040;
  assign n27780 = pi3316 & ~pi9040;
  assign n27781 = ~n27779 & ~n27780;
  assign n27782 = pi0393 & n27781;
  assign n27783 = ~pi0393 & ~n27781;
  assign n27784 = ~n27782 & ~n27783;
  assign n27785 = n27761 & ~n27784;
  assign n27786 = n27767 & n27785;
  assign n27787 = n27778 & ~n27786;
  assign n27788 = pi3279 & pi9040;
  assign n27789 = pi3274 & ~pi9040;
  assign n27790 = ~n27788 & ~n27789;
  assign n27791 = ~pi0388 & n27790;
  assign n27792 = pi0388 & ~n27790;
  assign n27793 = ~n27791 & ~n27792;
  assign n27794 = pi3380 & pi9040;
  assign n27795 = pi3301 & ~pi9040;
  assign n27796 = ~n27794 & ~n27795;
  assign n27797 = ~pi0395 & n27796;
  assign n27798 = pi0395 & ~n27796;
  assign n27799 = ~n27797 & ~n27798;
  assign n27800 = n27793 & ~n27799;
  assign n27801 = ~n27787 & n27800;
  assign n27802 = ~n27767 & n27773;
  assign n27803 = n27761 & n27802;
  assign n27804 = ~n27799 & n27803;
  assign n27805 = n27784 & n27804;
  assign n27806 = n27761 & n27774;
  assign n27807 = ~n27793 & n27806;
  assign n27808 = ~n27761 & n27767;
  assign n27809 = n27767 & n27773;
  assign n27810 = n27784 & n27809;
  assign n27811 = ~n27808 & ~n27810;
  assign n27812 = ~n27793 & ~n27811;
  assign n27813 = ~n27807 & ~n27812;
  assign n27814 = ~n27799 & ~n27813;
  assign n27815 = ~n27805 & ~n27814;
  assign n27816 = ~n27761 & n27784;
  assign n27817 = n27767 & n27816;
  assign n27818 = ~n27761 & ~n27784;
  assign n27819 = ~n27767 & n27818;
  assign n27820 = n27773 & n27819;
  assign n27821 = ~n27817 & ~n27820;
  assign n27822 = ~n27793 & ~n27821;
  assign n27823 = n27815 & ~n27822;
  assign n27824 = n27784 & n27793;
  assign n27825 = n27809 & n27824;
  assign n27826 = n27761 & n27825;
  assign n27827 = ~n27776 & ~n27802;
  assign n27828 = n27785 & ~n27827;
  assign n27829 = n27775 & ~n27784;
  assign n27830 = ~n27828 & ~n27829;
  assign n27831 = n27816 & ~n27827;
  assign n27832 = n27784 & n27806;
  assign n27833 = ~n27831 & ~n27832;
  assign n27834 = ~n27761 & n27809;
  assign n27835 = n27793 & n27834;
  assign n27836 = ~n27784 & n27835;
  assign n27837 = n27833 & ~n27836;
  assign n27838 = n27830 & n27837;
  assign n27839 = ~n27826 & n27838;
  assign n27840 = ~n27784 & ~n27793;
  assign n27841 = n27761 & n27840;
  assign n27842 = n27773 & n27841;
  assign n27843 = n27839 & ~n27842;
  assign n27844 = n27799 & ~n27843;
  assign n27845 = n27823 & ~n27844;
  assign n27846 = ~n27801 & n27845;
  assign n27847 = ~pi0444 & ~n27846;
  assign n27848 = pi0444 & n27823;
  assign n27849 = ~n27801 & n27848;
  assign n27850 = ~n27844 & n27849;
  assign po0468 = n27847 | n27850;
  assign n27852 = ~n26842 & n26866;
  assign n27853 = ~n26935 & ~n27852;
  assign n27854 = ~n26848 & n27853;
  assign n27855 = n26842 & n26890;
  assign n27856 = ~n26836 & ~n26860;
  assign n27857 = n26856 & ~n27856;
  assign n27858 = n26835 & n26897;
  assign n27859 = n26842 & n26860;
  assign n27860 = ~n27858 & ~n27859;
  assign n27861 = ~n27857 & n27860;
  assign n27862 = n26848 & n27861;
  assign n27863 = ~n27855 & n27862;
  assign n27864 = ~n27854 & ~n27863;
  assign n27865 = n26842 & n27857;
  assign n27866 = ~n26933 & ~n27865;
  assign n27867 = ~n27864 & n27866;
  assign n27868 = n26823 & ~n27867;
  assign n27869 = ~n26848 & ~n27856;
  assign n27870 = ~n26842 & n27869;
  assign n27871 = n26842 & n26884;
  assign n27872 = ~n26878 & ~n27871;
  assign n27873 = ~n26848 & ~n27872;
  assign n27874 = ~n26856 & n27869;
  assign n27875 = ~n27873 & ~n27874;
  assign n27876 = ~n27870 & n27875;
  assign n27877 = ~n26823 & ~n27876;
  assign n27878 = ~n27868 & ~n27877;
  assign n27879 = ~n26848 & n26864;
  assign n27880 = n26848 & ~n27866;
  assign n27881 = ~n27879 & ~n27880;
  assign n27882 = n26848 & ~n27853;
  assign n27883 = ~n26864 & ~n27882;
  assign n27884 = ~n26823 & ~n27883;
  assign n27885 = n27881 & ~n27884;
  assign n27886 = n27878 & n27885;
  assign n27887 = pi0452 & ~n27886;
  assign n27888 = ~pi0452 & n27885;
  assign n27889 = ~n27877 & n27888;
  assign n27890 = ~n27868 & n27889;
  assign po0469 = n27887 | n27890;
  assign n27892 = n27761 & n27809;
  assign n27893 = ~n27793 & n27892;
  assign n27894 = ~n27784 & n27893;
  assign n27895 = n27774 & n27840;
  assign n27896 = ~n27761 & n27895;
  assign n27897 = ~n27894 & ~n27896;
  assign n27898 = ~n27829 & ~n27836;
  assign n27899 = ~n27773 & n27784;
  assign n27900 = n27761 & n27899;
  assign n27901 = ~n27810 & ~n27900;
  assign n27902 = ~n27793 & ~n27901;
  assign n27903 = n27793 & ~n27818;
  assign n27904 = ~n27827 & n27903;
  assign n27905 = ~n27761 & ~n27809;
  assign n27906 = ~n27793 & n27905;
  assign n27907 = ~n27784 & n27906;
  assign n27908 = ~n27904 & ~n27907;
  assign n27909 = ~n27902 & n27908;
  assign n27910 = n27898 & n27909;
  assign n27911 = ~n27799 & ~n27910;
  assign n27912 = n27897 & ~n27911;
  assign n27913 = n27777 & n27793;
  assign n27914 = n27784 & n27913;
  assign n27915 = n27793 & n27799;
  assign n27916 = n27818 & ~n27827;
  assign n27917 = ~n27810 & ~n27916;
  assign n27918 = ~n27806 & n27917;
  assign n27919 = n27915 & ~n27918;
  assign n27920 = n27775 & n27784;
  assign n27921 = ~n27761 & n27899;
  assign n27922 = n27784 & n27802;
  assign n27923 = ~n27921 & ~n27922;
  assign n27924 = ~n27784 & n27809;
  assign n27925 = ~n27803 & ~n27924;
  assign n27926 = n27923 & n27925;
  assign n27927 = ~n27793 & ~n27926;
  assign n27928 = ~n27920 & ~n27927;
  assign n27929 = n27799 & ~n27928;
  assign n27930 = ~n27919 & ~n27929;
  assign n27931 = ~n27914 & n27930;
  assign n27932 = n27912 & n27931;
  assign n27933 = pi0434 & ~n27932;
  assign n27934 = ~pi0434 & n27912;
  assign n27935 = n27931 & n27934;
  assign po0471 = n27933 | n27935;
  assign n27937 = ~n27551 & ~n27557;
  assign n27938 = n27142 & ~n27937;
  assign n27939 = ~n27099 & n27133;
  assign n27940 = ~n27123 & n27149;
  assign n27941 = ~n27150 & ~n27940;
  assign n27942 = ~n27099 & ~n27941;
  assign n27943 = ~n27939 & ~n27942;
  assign n27944 = n27142 & ~n27943;
  assign n27945 = ~n27938 & ~n27944;
  assign n27946 = n27144 & n27153;
  assign n27947 = ~n27155 & ~n27946;
  assign n27948 = ~n27148 & ~n27185;
  assign n27949 = n27099 & ~n27948;
  assign n27950 = n27142 & n27949;
  assign n27951 = n27947 & ~n27950;
  assign n27952 = n27123 & n27149;
  assign n27953 = n27117 & n27952;
  assign n27954 = n27105 & n27124;
  assign n27955 = ~n27129 & ~n27954;
  assign n27956 = n27099 & ~n27955;
  assign n27957 = ~n27134 & ~n27158;
  assign n27958 = n27105 & n27143;
  assign n27959 = ~n27178 & ~n27958;
  assign n27960 = ~n27099 & ~n27959;
  assign n27961 = n27957 & ~n27960;
  assign n27962 = ~n27956 & n27961;
  assign n27963 = ~n27953 & n27962;
  assign n27964 = ~n27142 & ~n27963;
  assign n27965 = ~n27182 & n27220;
  assign n27966 = n27099 & ~n27965;
  assign n27967 = ~n27964 & ~n27966;
  assign n27968 = n27951 & n27967;
  assign n27969 = n27945 & n27968;
  assign n27970 = ~pi0441 & ~n27969;
  assign n27971 = pi0441 & n27951;
  assign n27972 = n27945 & n27971;
  assign n27973 = n27967 & n27972;
  assign po0472 = n27970 | n27973;
  assign n27975 = ~n27588 & n27607;
  assign n27976 = ~n27632 & ~n27647;
  assign n27977 = n27975 & ~n27976;
  assign n27978 = ~n27588 & ~n27613;
  assign n27979 = n27632 & n27978;
  assign n27980 = ~n27977 & ~n27979;
  assign n27981 = n27625 & ~n27980;
  assign n27982 = ~n27607 & n27613;
  assign n27983 = n27600 & n27982;
  assign n27984 = n27594 & n27983;
  assign n27985 = ~n27664 & ~n27982;
  assign n27986 = n27588 & ~n27985;
  assign n27987 = ~n27607 & ~n27613;
  assign n27988 = ~n27600 & n27987;
  assign n27989 = n27594 & n27988;
  assign n27990 = ~n27986 & ~n27989;
  assign n27991 = ~n27984 & n27990;
  assign n27992 = n27625 & ~n27991;
  assign n27993 = ~n27981 & ~n27992;
  assign n27994 = n27600 & n27614;
  assign n27995 = ~n27594 & n27994;
  assign n27996 = ~n27607 & n27639;
  assign n27997 = ~n27995 & ~n27996;
  assign n27998 = ~n27588 & ~n27997;
  assign n27999 = ~n27601 & ~n27664;
  assign n28000 = n27607 & ~n27999;
  assign n28001 = ~n27639 & ~n28000;
  assign n28002 = ~n27588 & ~n28001;
  assign n28003 = n27600 & ~n27607;
  assign n28004 = ~n27588 & n28003;
  assign n28005 = ~n27613 & n28004;
  assign n28006 = ~n27600 & n27613;
  assign n28007 = ~n27639 & ~n28006;
  assign n28008 = ~n27607 & ~n28007;
  assign n28009 = n27588 & n27607;
  assign n28010 = n27629 & n28009;
  assign n28011 = ~n27613 & n28010;
  assign n28012 = ~n28008 & ~n28011;
  assign n28013 = ~n28005 & n28012;
  assign n28014 = ~n28002 & n28013;
  assign n28015 = ~n27995 & n28014;
  assign n28016 = ~n27625 & ~n28015;
  assign n28017 = ~n27607 & n27664;
  assign n28018 = n27607 & n27655;
  assign n28019 = ~n28017 & ~n28018;
  assign n28020 = n27588 & ~n28019;
  assign n28021 = ~n28016 & ~n28020;
  assign n28022 = ~n27998 & n28021;
  assign n28023 = n27993 & n28022;
  assign n28024 = pi0423 & n28023;
  assign n28025 = ~pi0423 & ~n28023;
  assign po0473 = n28024 | n28025;
  assign n28027 = ~n27600 & n27616;
  assign n28028 = ~n27647 & ~n28027;
  assign n28029 = ~n27588 & ~n28028;
  assign n28030 = n27607 & n27638;
  assign n28031 = ~n27988 & ~n28030;
  assign n28032 = n27588 & ~n28031;
  assign n28033 = ~n27607 & n27633;
  assign n28034 = ~n28005 & ~n28033;
  assign n28035 = ~n27615 & n28034;
  assign n28036 = ~n28032 & n28035;
  assign n28037 = ~n28029 & n28036;
  assign n28038 = ~n27984 & ~n27995;
  assign n28039 = n28037 & n28038;
  assign n28040 = n27625 & ~n28039;
  assign n28041 = n27601 & n27982;
  assign n28042 = n27656 & ~n28041;
  assign n28043 = n27588 & ~n28042;
  assign n28044 = ~n27607 & n27644;
  assign n28045 = ~n28043 & ~n28044;
  assign n28046 = n27594 & n27616;
  assign n28047 = n27607 & n27629;
  assign n28048 = ~n28046 & ~n28047;
  assign n28049 = n27588 & ~n28048;
  assign n28050 = n27588 & n27638;
  assign n28051 = ~n27607 & n28050;
  assign n28052 = ~n28049 & ~n28051;
  assign n28053 = n28045 & n28052;
  assign n28054 = ~n27625 & ~n28053;
  assign n28055 = ~n27633 & ~n27640;
  assign n28056 = ~n27989 & n28055;
  assign n28057 = n27661 & ~n28056;
  assign n28058 = ~n28054 & ~n28057;
  assign n28059 = ~n27615 & ~n27984;
  assign n28060 = ~n27588 & ~n28059;
  assign n28061 = n28058 & ~n28060;
  assign n28062 = ~n28040 & n28061;
  assign n28063 = ~pi0425 & n28062;
  assign n28064 = pi0425 & ~n28062;
  assign po0474 = n28063 | n28064;
  assign n28066 = ~n26602 & ~n26608;
  assign n28067 = ~n26573 & ~n28066;
  assign n28068 = ~n26664 & ~n28067;
  assign n28069 = ~n26580 & ~n26587;
  assign n28070 = n26573 & n28069;
  assign n28071 = ~n26601 & n28070;
  assign n28072 = ~n26573 & n26594;
  assign n28073 = ~n26601 & n28072;
  assign n28074 = ~n27512 & ~n28073;
  assign n28075 = n26587 & n27474;
  assign n28076 = ~n26601 & n26627;
  assign n28077 = ~n28075 & ~n28076;
  assign n28078 = ~n28069 & n28077;
  assign n28079 = n26573 & ~n28078;
  assign n28080 = ~n26611 & ~n28079;
  assign n28081 = n28074 & n28080;
  assign n28082 = ~n26640 & ~n28081;
  assign n28083 = ~n28071 & ~n28082;
  assign n28084 = ~n26628 & ~n26647;
  assign n28085 = ~n26657 & n28084;
  assign n28086 = ~n26573 & ~n28085;
  assign n28087 = n26601 & n26652;
  assign n28088 = ~n26631 & ~n28087;
  assign n28089 = n26573 & ~n28088;
  assign n28090 = ~n27519 & ~n28089;
  assign n28091 = ~n28086 & n28090;
  assign n28092 = ~n26617 & ~n26658;
  assign n28093 = n28091 & n28092;
  assign n28094 = n26640 & ~n28093;
  assign n28095 = n28083 & ~n28094;
  assign n28096 = n28068 & n28095;
  assign n28097 = ~pi0449 & ~n28096;
  assign n28098 = pi0449 & n28083;
  assign n28099 = n28068 & n28098;
  assign n28100 = ~n28094 & n28099;
  assign po0475 = n28097 | n28100;
  assign n28102 = ~n27761 & n27922;
  assign n28103 = ~n27832 & ~n28102;
  assign n28104 = ~n27793 & ~n28103;
  assign n28105 = ~n27761 & n27776;
  assign n28106 = ~n27892 & ~n28105;
  assign n28107 = ~n27793 & ~n28106;
  assign n28108 = ~n27784 & n27802;
  assign n28109 = ~n27777 & ~n28108;
  assign n28110 = ~n27834 & n28109;
  assign n28111 = n27793 & ~n28110;
  assign n28112 = ~n28107 & ~n28111;
  assign n28113 = ~n27807 & ~n27820;
  assign n28114 = n28112 & n28113;
  assign n28115 = n27799 & ~n28114;
  assign n28116 = n27784 & n27892;
  assign n28117 = n27774 & ~n27784;
  assign n28118 = ~n27922 & ~n28117;
  assign n28119 = n27793 & ~n28118;
  assign n28120 = ~n28116 & ~n28119;
  assign n28121 = n27761 & ~n27793;
  assign n28122 = ~n27767 & n28121;
  assign n28123 = n27773 & n28122;
  assign n28124 = n27778 & ~n28123;
  assign n28125 = ~n27834 & n28124;
  assign n28126 = ~n27784 & ~n28125;
  assign n28127 = n28120 & ~n28126;
  assign n28128 = ~n27799 & ~n28127;
  assign n28129 = ~n28115 & ~n28128;
  assign n28130 = ~n27761 & ~n27773;
  assign n28131 = n27824 & n28130;
  assign n28132 = n28129 & ~n28131;
  assign n28133 = ~n28104 & n28132;
  assign n28134 = ~pi0428 & ~n28133;
  assign n28135 = pi0428 & ~n28104;
  assign n28136 = n28129 & n28135;
  assign n28137 = ~n28131 & n28136;
  assign po0476 = n28134 | n28137;
  assign n28139 = ~n27803 & ~n27899;
  assign n28140 = n27800 & ~n28139;
  assign n28141 = n27761 & n27784;
  assign n28142 = ~n27776 & n28141;
  assign n28143 = ~n27799 & n28142;
  assign n28144 = ~n27793 & n27816;
  assign n28145 = n27776 & n28144;
  assign n28146 = n27761 & n27824;
  assign n28147 = ~n27767 & n28146;
  assign n28148 = ~n28145 & ~n28147;
  assign n28149 = ~n28143 & n28148;
  assign n28150 = ~n27922 & ~n27924;
  assign n28151 = ~n27793 & ~n28150;
  assign n28152 = ~n27896 & ~n28151;
  assign n28153 = ~n27799 & ~n28152;
  assign n28154 = ~n27776 & ~n28130;
  assign n28155 = ~n27784 & ~n28154;
  assign n28156 = ~n27892 & ~n28155;
  assign n28157 = n27793 & ~n28156;
  assign n28158 = ~n27916 & ~n28157;
  assign n28159 = n27784 & n27834;
  assign n28160 = ~n27767 & n27785;
  assign n28161 = n27784 & ~n28154;
  assign n28162 = ~n28160 & ~n28161;
  assign n28163 = ~n27793 & ~n28162;
  assign n28164 = ~n28159 & ~n28163;
  assign n28165 = n28158 & n28164;
  assign n28166 = n27799 & ~n28165;
  assign n28167 = ~n28153 & ~n28166;
  assign n28168 = n28149 & n28167;
  assign n28169 = ~n28140 & n28168;
  assign n28170 = pi0438 & ~n28169;
  assign n28171 = ~pi0438 & n28149;
  assign n28172 = ~n28140 & n28171;
  assign n28173 = n28167 & n28172;
  assign po0477 = n28170 | n28173;
  assign n28175 = ~n27352 & ~n27435;
  assign n28176 = ~n27423 & n28175;
  assign n28177 = n27359 & ~n28176;
  assign n28178 = ~n27373 & ~n27399;
  assign n28179 = ~n27368 & ~n27431;
  assign n28180 = ~n27343 & ~n27438;
  assign n28181 = ~n27359 & ~n28180;
  assign n28182 = ~n27410 & ~n28181;
  assign n28183 = n28179 & n28182;
  assign n28184 = n27316 & ~n28183;
  assign n28185 = n27328 & n27341;
  assign n28186 = ~n27678 & ~n28185;
  assign n28187 = ~n27322 & ~n28186;
  assign n28188 = ~n27379 & ~n27383;
  assign n28189 = ~n27359 & ~n28188;
  assign n28190 = ~n27322 & n27341;
  assign n28191 = ~n27350 & ~n28190;
  assign n28192 = ~n27342 & n28191;
  assign n28193 = n27359 & ~n28192;
  assign n28194 = ~n28189 & ~n28193;
  assign n28195 = ~n28187 & n28194;
  assign n28196 = ~n27316 & ~n28195;
  assign n28197 = ~n28184 & ~n28196;
  assign n28198 = n28178 & n28197;
  assign n28199 = ~n28177 & n28198;
  assign n28200 = ~pi0439 & ~n28199;
  assign n28201 = pi0439 & n28178;
  assign n28202 = ~n28177 & n28201;
  assign n28203 = n28197 & n28202;
  assign po0478 = n28200 | n28203;
  assign n28205 = n27017 & ~n27264;
  assign n28206 = n26998 & n28205;
  assign n28207 = n27010 & n27241;
  assign n28208 = ~n27081 & ~n28207;
  assign n28209 = ~n27031 & n28208;
  assign n28210 = ~n27023 & ~n28209;
  assign n28211 = ~n27045 & ~n27252;
  assign n28212 = n27023 & ~n28211;
  assign n28213 = ~n28210 & ~n28212;
  assign n28214 = ~n28206 & n28213;
  assign n28215 = ~n27017 & n27058;
  assign n28216 = n28214 & ~n28215;
  assign n28217 = ~n26992 & ~n28216;
  assign n28218 = n27027 & ~n28211;
  assign n28219 = ~n27046 & ~n27061;
  assign n28220 = ~n27031 & ~n27058;
  assign n28221 = n28219 & n28220;
  assign n28222 = n27017 & ~n28221;
  assign n28223 = ~n28218 & ~n28222;
  assign n28224 = ~n27243 & n28223;
  assign n28225 = n26992 & ~n28224;
  assign n28226 = ~n28217 & ~n28225;
  assign n28227 = n27017 & n27252;
  assign n28228 = ~n28215 & ~n28227;
  assign n28229 = n27023 & ~n28228;
  assign n28230 = n28226 & ~n28229;
  assign n28231 = pi0417 & ~n28230;
  assign n28232 = ~pi0417 & ~n28229;
  assign n28233 = ~n28225 & n28232;
  assign n28234 = ~n28217 & n28233;
  assign po0479 = n28231 | n28234;
  assign n28236 = ~n26848 & n26883;
  assign n28237 = n26897 & ~n27856;
  assign n28238 = ~n26885 & ~n28237;
  assign n28239 = ~n26933 & n28238;
  assign n28240 = n26848 & ~n28239;
  assign n28241 = n26842 & n26861;
  assign n28242 = ~n28240 & ~n28241;
  assign n28243 = ~n26856 & n26884;
  assign n28244 = ~n26842 & n26940;
  assign n28245 = ~n28243 & ~n28244;
  assign n28246 = ~n27859 & n28245;
  assign n28247 = ~n26848 & ~n28246;
  assign n28248 = n28242 & ~n28247;
  assign n28249 = n26823 & ~n28248;
  assign n28250 = ~n28236 & ~n28249;
  assign n28251 = ~n26842 & n26860;
  assign n28252 = ~n26932 & ~n28251;
  assign n28253 = ~n26848 & ~n28252;
  assign n28254 = ~n26886 & ~n28253;
  assign n28255 = ~n26878 & ~n26883;
  assign n28256 = n26842 & n26902;
  assign n28257 = ~n26940 & ~n28256;
  assign n28258 = ~n28243 & n28257;
  assign n28259 = n26848 & ~n28258;
  assign n28260 = ~n26842 & n26861;
  assign n28261 = ~n28259 & ~n28260;
  assign n28262 = n28255 & n28261;
  assign n28263 = n28254 & n28262;
  assign n28264 = ~n26823 & ~n28263;
  assign n28265 = ~n26907 & ~n27855;
  assign n28266 = n26848 & ~n28265;
  assign n28267 = ~n28264 & ~n28266;
  assign n28268 = n28250 & n28267;
  assign n28269 = pi0458 & n28268;
  assign n28270 = ~pi0458 & ~n28268;
  assign po0480 = n28269 | n28270;
  assign n28272 = ~n27588 & n27644;
  assign n28273 = ~n27607 & n27629;
  assign n28274 = ~n27628 & ~n28273;
  assign n28275 = ~n27588 & ~n28274;
  assign n28276 = n27588 & ~n28007;
  assign n28277 = ~n28275 & ~n28276;
  assign n28278 = ~n28018 & n28277;
  assign n28279 = n27625 & ~n28278;
  assign n28280 = ~n28272 & ~n28279;
  assign n28281 = n27613 & n27975;
  assign n28282 = ~n27987 & ~n28281;
  assign n28283 = ~n27594 & ~n28282;
  assign n28284 = ~n27615 & ~n28283;
  assign n28285 = ~n27988 & n28284;
  assign n28286 = n27607 & n27647;
  assign n28287 = n27588 & n27630;
  assign n28288 = ~n28286 & ~n28287;
  assign n28289 = n28285 & n28288;
  assign n28290 = ~n27625 & ~n28289;
  assign n28291 = ~n28033 & ~n28047;
  assign n28292 = n27588 & ~n28291;
  assign n28293 = ~n28290 & ~n28292;
  assign n28294 = n28280 & n28293;
  assign n28295 = ~pi0454 & ~n28294;
  assign n28296 = pi0454 & n28293;
  assign n28297 = ~n28279 & n28296;
  assign n28298 = ~n28272 & n28297;
  assign po0481 = n28295 | n28298;
  assign n28300 = pi3480 & pi9040;
  assign n28301 = pi3415 & ~pi9040;
  assign n28302 = ~n28300 & ~n28301;
  assign n28303 = ~pi0440 & n28302;
  assign n28304 = pi0440 & ~n28302;
  assign n28305 = ~n28303 & ~n28304;
  assign n28306 = pi3372 & pi9040;
  assign n28307 = pi3395 & ~pi9040;
  assign n28308 = ~n28306 & ~n28307;
  assign n28309 = ~pi0450 & n28308;
  assign n28310 = pi0450 & ~n28308;
  assign n28311 = ~n28309 & ~n28310;
  assign n28312 = pi3396 & pi9040;
  assign n28313 = pi3464 & ~pi9040;
  assign n28314 = ~n28312 & ~n28313;
  assign n28315 = ~pi0473 & n28314;
  assign n28316 = pi0473 & ~n28314;
  assign n28317 = ~n28315 & ~n28316;
  assign n28318 = pi3418 & pi9040;
  assign n28319 = pi3411 & ~pi9040;
  assign n28320 = ~n28318 & ~n28319;
  assign n28321 = ~pi0443 & n28320;
  assign n28322 = pi0443 & ~n28320;
  assign n28323 = ~n28321 & ~n28322;
  assign n28324 = ~n28317 & ~n28323;
  assign n28325 = n28311 & n28324;
  assign n28326 = pi3412 & pi9040;
  assign n28327 = pi3373 & ~pi9040;
  assign n28328 = ~n28326 & ~n28327;
  assign n28329 = pi0469 & n28328;
  assign n28330 = ~pi0469 & ~n28328;
  assign n28331 = ~n28329 & ~n28330;
  assign n28332 = n28325 & ~n28331;
  assign n28333 = n28317 & n28323;
  assign n28334 = n28311 & n28333;
  assign n28335 = ~n28331 & n28334;
  assign n28336 = ~n28332 & ~n28335;
  assign n28337 = ~n28311 & n28331;
  assign n28338 = n28333 & n28337;
  assign n28339 = ~n28317 & n28323;
  assign n28340 = n28311 & n28339;
  assign n28341 = n28331 & n28340;
  assign n28342 = ~n28338 & ~n28341;
  assign n28343 = n28336 & n28342;
  assign n28344 = ~n28305 & ~n28343;
  assign n28345 = n28311 & n28331;
  assign n28346 = ~n28323 & n28345;
  assign n28347 = n28317 & n28346;
  assign n28348 = ~n28340 & ~n28347;
  assign n28349 = ~n28305 & ~n28348;
  assign n28350 = ~n28323 & ~n28331;
  assign n28351 = n28305 & n28350;
  assign n28352 = ~n28311 & ~n28317;
  assign n28353 = n28331 & n28333;
  assign n28354 = ~n28352 & ~n28353;
  assign n28355 = n28305 & ~n28354;
  assign n28356 = ~n28351 & ~n28355;
  assign n28357 = n28317 & ~n28323;
  assign n28358 = ~n28311 & n28357;
  assign n28359 = ~n28331 & n28358;
  assign n28360 = n28356 & ~n28359;
  assign n28361 = ~n28323 & n28352;
  assign n28362 = n28331 & n28361;
  assign n28363 = n28360 & ~n28362;
  assign n28364 = ~n28349 & n28363;
  assign n28365 = pi3361 & ~pi9040;
  assign n28366 = ~pi3383 & pi9040;
  assign n28367 = ~n28365 & ~n28366;
  assign n28368 = pi0479 & n28367;
  assign n28369 = ~pi0479 & ~n28367;
  assign n28370 = ~n28368 & ~n28369;
  assign n28371 = ~n28364 & n28370;
  assign n28372 = n28311 & ~n28323;
  assign n28373 = n28305 & n28331;
  assign n28374 = ~n28370 & n28373;
  assign n28375 = n28372 & n28374;
  assign n28376 = n28311 & ~n28331;
  assign n28377 = n28323 & n28376;
  assign n28378 = n28305 & ~n28377;
  assign n28379 = n28317 & n28337;
  assign n28380 = ~n28311 & n28333;
  assign n28381 = ~n28324 & ~n28372;
  assign n28382 = ~n28331 & ~n28381;
  assign n28383 = ~n28380 & ~n28382;
  assign n28384 = ~n28305 & n28383;
  assign n28385 = ~n28379 & n28384;
  assign n28386 = ~n28378 & ~n28385;
  assign n28387 = ~n28311 & n28339;
  assign n28388 = n28331 & n28387;
  assign n28389 = ~n28386 & ~n28388;
  assign n28390 = ~n28370 & ~n28389;
  assign n28391 = ~n28375 & ~n28390;
  assign n28392 = ~n28371 & n28391;
  assign n28393 = ~n28344 & n28392;
  assign n28394 = n28305 & n28359;
  assign n28395 = n28393 & ~n28394;
  assign n28396 = pi0480 & ~n28395;
  assign n28397 = n28392 & ~n28394;
  assign n28398 = ~pi0480 & n28397;
  assign n28399 = ~n28344 & n28398;
  assign po0506 = n28396 | n28399;
  assign n28401 = pi3409 & pi9040;
  assign n28402 = pi3412 & ~pi9040;
  assign n28403 = ~n28401 & ~n28402;
  assign n28404 = pi0453 & n28403;
  assign n28405 = ~pi0453 & ~n28403;
  assign n28406 = ~n28404 & ~n28405;
  assign n28407 = pi3458 & ~pi9040;
  assign n28408 = pi3419 & pi9040;
  assign n28409 = ~n28407 & ~n28408;
  assign n28410 = ~pi0461 & ~n28409;
  assign n28411 = pi0461 & n28409;
  assign n28412 = ~n28410 & ~n28411;
  assign n28413 = ~n28406 & ~n28412;
  assign n28414 = pi3411 & pi9040;
  assign n28415 = pi3392 & ~pi9040;
  assign n28416 = ~n28414 & ~n28415;
  assign n28417 = ~pi0462 & ~n28416;
  assign n28418 = pi0462 & ~n28414;
  assign n28419 = ~n28415 & n28418;
  assign n28420 = ~n28417 & ~n28419;
  assign n28421 = pi3368 & pi9040;
  assign n28422 = pi3409 & ~pi9040;
  assign n28423 = ~n28421 & ~n28422;
  assign n28424 = ~pi0476 & ~n28423;
  assign n28425 = pi0476 & n28423;
  assign n28426 = ~n28424 & ~n28425;
  assign n28427 = pi3371 & pi9040;
  assign n28428 = pi3398 & ~pi9040;
  assign n28429 = ~n28427 & ~n28428;
  assign n28430 = ~pi0463 & ~n28429;
  assign n28431 = pi0463 & n28429;
  assign n28432 = ~n28430 & ~n28431;
  assign n28433 = n28426 & ~n28432;
  assign n28434 = ~n28420 & n28433;
  assign n28435 = pi3393 & pi9040;
  assign n28436 = pi3413 & ~pi9040;
  assign n28437 = ~n28435 & ~n28436;
  assign n28438 = ~pi0457 & ~n28437;
  assign n28439 = pi0457 & ~n28435;
  assign n28440 = ~n28436 & n28439;
  assign n28441 = ~n28438 & ~n28440;
  assign n28442 = n28432 & ~n28441;
  assign n28443 = n28426 & n28442;
  assign n28444 = n28420 & n28443;
  assign n28445 = n28432 & n28441;
  assign n28446 = ~n28420 & n28445;
  assign n28447 = ~n28444 & ~n28446;
  assign n28448 = ~n28434 & n28447;
  assign n28449 = n28413 & ~n28448;
  assign n28450 = ~n28420 & ~n28426;
  assign n28451 = ~n28441 & n28450;
  assign n28452 = ~n28432 & ~n28441;
  assign n28453 = n28426 & n28452;
  assign n28454 = n28420 & n28453;
  assign n28455 = ~n28451 & ~n28454;
  assign n28456 = ~n28426 & n28442;
  assign n28457 = n28426 & n28445;
  assign n28458 = ~n28456 & ~n28457;
  assign n28459 = n28455 & n28458;
  assign n28460 = n28406 & ~n28459;
  assign n28461 = ~n28432 & n28441;
  assign n28462 = ~n28426 & n28461;
  assign n28463 = n28420 & n28462;
  assign n28464 = ~n28460 & ~n28463;
  assign n28465 = ~n28412 & ~n28464;
  assign n28466 = ~n28449 & ~n28465;
  assign n28467 = n28406 & ~n28420;
  assign n28468 = n28426 & n28467;
  assign n28469 = n28441 & n28468;
  assign n28470 = ~n28420 & n28456;
  assign n28471 = ~n28469 & ~n28470;
  assign n28472 = ~n28426 & n28452;
  assign n28473 = ~n28445 & ~n28452;
  assign n28474 = n28420 & ~n28473;
  assign n28475 = ~n28472 & ~n28474;
  assign n28476 = ~n28406 & ~n28475;
  assign n28477 = n28426 & n28461;
  assign n28478 = ~n28434 & ~n28477;
  assign n28479 = ~n28444 & n28478;
  assign n28480 = n28406 & ~n28479;
  assign n28481 = ~n28476 & ~n28480;
  assign n28482 = ~n28406 & ~n28420;
  assign n28483 = n28442 & n28482;
  assign n28484 = n28420 & n28472;
  assign n28485 = ~n28426 & n28432;
  assign n28486 = n28441 & n28485;
  assign n28487 = n28420 & n28486;
  assign n28488 = ~n28484 & ~n28487;
  assign n28489 = n28441 & n28450;
  assign n28490 = ~n28432 & n28489;
  assign n28491 = n28488 & ~n28490;
  assign n28492 = ~n28483 & n28491;
  assign n28493 = n28481 & n28492;
  assign n28494 = n28412 & ~n28493;
  assign n28495 = n28471 & ~n28494;
  assign n28496 = n28466 & n28495;
  assign n28497 = pi0491 & ~n28496;
  assign n28498 = ~pi0491 & n28471;
  assign n28499 = n28466 & n28498;
  assign n28500 = ~n28494 & n28499;
  assign po0512 = n28497 | n28500;
  assign n28502 = pi3395 & pi9040;
  assign n28503 = pi3375 & ~pi9040;
  assign n28504 = ~n28502 & ~n28503;
  assign n28505 = pi0463 & n28504;
  assign n28506 = ~pi0463 & ~n28504;
  assign n28507 = ~n28505 & ~n28506;
  assign n28508 = pi3399 & pi9040;
  assign n28509 = pi3480 & ~pi9040;
  assign n28510 = ~n28508 & ~n28509;
  assign n28511 = ~pi0471 & n28510;
  assign n28512 = pi0471 & ~n28510;
  assign n28513 = ~n28511 & ~n28512;
  assign n28514 = pi3415 & pi9040;
  assign n28515 = pi3418 & ~pi9040;
  assign n28516 = ~n28514 & ~n28515;
  assign n28517 = ~pi0468 & ~n28516;
  assign n28518 = pi0468 & ~n28514;
  assign n28519 = ~n28515 & n28518;
  assign n28520 = ~n28517 & ~n28519;
  assign n28521 = pi3375 & pi9040;
  assign n28522 = pi3383 & ~pi9040;
  assign n28523 = ~n28521 & ~n28522;
  assign n28524 = pi0442 & n28523;
  assign n28525 = ~pi0442 & ~n28523;
  assign n28526 = ~n28524 & ~n28525;
  assign n28527 = pi3373 & pi9040;
  assign n28528 = pi3396 & ~pi9040;
  assign n28529 = ~n28527 & ~n28528;
  assign n28530 = pi0476 & n28529;
  assign n28531 = ~pi0476 & ~n28529;
  assign n28532 = ~n28530 & ~n28531;
  assign n28533 = n28526 & ~n28532;
  assign n28534 = n28520 & n28533;
  assign n28535 = ~n28513 & n28534;
  assign n28536 = n28513 & n28526;
  assign n28537 = n28532 & n28536;
  assign n28538 = pi3464 & pi9040;
  assign n28539 = pi3372 & ~pi9040;
  assign n28540 = ~n28538 & ~n28539;
  assign n28541 = pi0459 & n28540;
  assign n28542 = ~pi0459 & ~n28540;
  assign n28543 = ~n28541 & ~n28542;
  assign n28544 = ~n28520 & n28536;
  assign n28545 = n28520 & n28532;
  assign n28546 = ~n28526 & n28545;
  assign n28547 = ~n28544 & ~n28546;
  assign n28548 = ~n28543 & ~n28547;
  assign n28549 = ~n28537 & ~n28548;
  assign n28550 = n28526 & n28545;
  assign n28551 = ~n28520 & ~n28526;
  assign n28552 = ~n28526 & ~n28532;
  assign n28553 = n28513 & n28552;
  assign n28554 = ~n28520 & ~n28532;
  assign n28555 = ~n28513 & n28554;
  assign n28556 = ~n28553 & ~n28555;
  assign n28557 = ~n28551 & n28556;
  assign n28558 = ~n28550 & n28557;
  assign n28559 = n28543 & ~n28558;
  assign n28560 = n28549 & ~n28559;
  assign n28561 = ~n28535 & n28560;
  assign n28562 = n28507 & ~n28561;
  assign n28563 = ~n28520 & n28532;
  assign n28564 = ~n28526 & n28563;
  assign n28565 = n28513 & n28564;
  assign n28566 = ~n28526 & n28554;
  assign n28567 = ~n28513 & n28566;
  assign n28568 = ~n28535 & ~n28567;
  assign n28569 = ~n28565 & n28568;
  assign n28570 = n28543 & ~n28569;
  assign n28571 = ~n28562 & ~n28570;
  assign n28572 = n28513 & n28550;
  assign n28573 = n28520 & ~n28526;
  assign n28574 = ~n28543 & n28573;
  assign n28575 = ~n28513 & n28574;
  assign n28576 = n28526 & n28563;
  assign n28577 = ~n28513 & n28576;
  assign n28578 = n28533 & n28543;
  assign n28579 = n28513 & n28578;
  assign n28580 = ~n28577 & ~n28579;
  assign n28581 = ~n28520 & n28526;
  assign n28582 = ~n28513 & n28581;
  assign n28583 = n28520 & ~n28532;
  assign n28584 = ~n28526 & n28583;
  assign n28585 = ~n28582 & ~n28584;
  assign n28586 = ~n28543 & ~n28585;
  assign n28587 = ~n28543 & n28551;
  assign n28588 = n28513 & n28587;
  assign n28589 = ~n28586 & ~n28588;
  assign n28590 = n28580 & n28589;
  assign n28591 = ~n28507 & ~n28590;
  assign n28592 = ~n28575 & ~n28591;
  assign n28593 = ~n28572 & n28592;
  assign n28594 = n28571 & n28593;
  assign n28595 = ~pi0498 & ~n28594;
  assign n28596 = ~n28562 & ~n28572;
  assign n28597 = ~n28570 & n28596;
  assign n28598 = n28592 & n28597;
  assign n28599 = pi0498 & n28598;
  assign po0513 = n28595 | n28599;
  assign n28601 = pi3454 & ~pi9040;
  assign n28602 = pi3367 & pi9040;
  assign n28603 = ~n28601 & ~n28602;
  assign n28604 = ~pi0468 & ~n28603;
  assign n28605 = pi0468 & n28603;
  assign n28606 = ~n28604 & ~n28605;
  assign n28607 = pi3370 & pi9040;
  assign n28608 = pi3397 & ~pi9040;
  assign n28609 = ~n28607 & ~n28608;
  assign n28610 = ~pi0465 & n28609;
  assign n28611 = pi0465 & ~n28609;
  assign n28612 = ~n28610 & ~n28611;
  assign n28613 = pi3381 & pi9040;
  assign n28614 = pi3455 & ~pi9040;
  assign n28615 = ~n28613 & ~n28614;
  assign n28616 = ~pi0467 & n28615;
  assign n28617 = pi0467 & ~n28615;
  assign n28618 = ~n28616 & ~n28617;
  assign n28619 = pi3410 & pi9040;
  assign n28620 = pi3388 & ~pi9040;
  assign n28621 = ~n28619 & ~n28620;
  assign n28622 = ~pi0472 & ~n28621;
  assign n28623 = pi0472 & ~n28619;
  assign n28624 = ~n28620 & n28623;
  assign n28625 = ~n28622 & ~n28624;
  assign n28626 = pi3376 & pi9040;
  assign n28627 = pi3381 & ~pi9040;
  assign n28628 = ~n28626 & ~n28627;
  assign n28629 = ~pi0442 & n28628;
  assign n28630 = pi0442 & ~n28628;
  assign n28631 = ~n28629 & ~n28630;
  assign n28632 = ~n28625 & ~n28631;
  assign n28633 = ~n28618 & n28632;
  assign n28634 = ~n28612 & n28633;
  assign n28635 = pi3452 & pi9040;
  assign n28636 = pi3377 & ~pi9040;
  assign n28637 = ~n28635 & ~n28636;
  assign n28638 = pi0475 & n28637;
  assign n28639 = ~pi0475 & ~n28637;
  assign n28640 = ~n28638 & ~n28639;
  assign n28641 = n28625 & ~n28631;
  assign n28642 = ~n28612 & n28641;
  assign n28643 = n28618 & n28632;
  assign n28644 = n28612 & n28643;
  assign n28645 = ~n28642 & ~n28644;
  assign n28646 = ~n28640 & ~n28645;
  assign n28647 = ~n28634 & ~n28646;
  assign n28648 = ~n28625 & n28631;
  assign n28649 = n28618 & n28648;
  assign n28650 = n28640 & n28649;
  assign n28651 = n28632 & n28640;
  assign n28652 = ~n28612 & n28651;
  assign n28653 = ~n28650 & ~n28652;
  assign n28654 = n28647 & n28653;
  assign n28655 = n28625 & n28631;
  assign n28656 = ~n28618 & n28655;
  assign n28657 = ~n28612 & n28656;
  assign n28658 = ~n28618 & n28648;
  assign n28659 = n28612 & n28658;
  assign n28660 = ~n28657 & ~n28659;
  assign n28661 = n28654 & n28660;
  assign n28662 = n28606 & ~n28661;
  assign n28663 = ~n28606 & ~n28640;
  assign n28664 = ~n28612 & n28618;
  assign n28665 = ~n28625 & n28664;
  assign n28666 = n28618 & n28631;
  assign n28667 = ~n28665 & ~n28666;
  assign n28668 = n28663 & ~n28667;
  assign n28669 = n28618 & n28655;
  assign n28670 = n28612 & ~n28640;
  assign n28671 = n28669 & n28670;
  assign n28672 = ~n28618 & n28641;
  assign n28673 = n28612 & n28672;
  assign n28674 = ~n28659 & ~n28673;
  assign n28675 = ~n28640 & ~n28674;
  assign n28676 = ~n28671 & ~n28675;
  assign n28677 = n28612 & n28625;
  assign n28678 = n28618 & n28677;
  assign n28679 = n28612 & ~n28618;
  assign n28680 = ~n28631 & n28679;
  assign n28681 = ~n28625 & n28680;
  assign n28682 = ~n28678 & ~n28681;
  assign n28683 = ~n28612 & n28640;
  assign n28684 = ~n28618 & n28683;
  assign n28685 = ~n28632 & n28684;
  assign n28686 = n28640 & n28656;
  assign n28687 = ~n28685 & ~n28686;
  assign n28688 = n28682 & n28687;
  assign n28689 = ~n28606 & ~n28688;
  assign n28690 = n28640 & n28681;
  assign n28691 = ~n28689 & ~n28690;
  assign n28692 = n28676 & n28691;
  assign n28693 = ~n28668 & n28692;
  assign n28694 = ~n28662 & n28693;
  assign n28695 = n28618 & n28641;
  assign n28696 = n28612 & n28640;
  assign n28697 = n28695 & n28696;
  assign n28698 = n28694 & ~n28697;
  assign n28699 = ~pi0489 & ~n28698;
  assign n28700 = pi0489 & ~n28697;
  assign n28701 = n28693 & n28700;
  assign n28702 = ~n28662 & n28701;
  assign po0514 = n28699 | n28702;
  assign n28704 = n28513 & ~n28543;
  assign n28705 = n28520 & n28704;
  assign n28706 = n28526 & n28554;
  assign n28707 = ~n28513 & n28706;
  assign n28708 = ~n28513 & n28564;
  assign n28709 = ~n28707 & ~n28708;
  assign n28710 = n28513 & ~n28526;
  assign n28711 = ~n28532 & n28710;
  assign n28712 = ~n28520 & n28711;
  assign n28713 = ~n28546 & ~n28712;
  assign n28714 = n28543 & ~n28713;
  assign n28715 = n28709 & ~n28714;
  assign n28716 = ~n28705 & n28715;
  assign n28717 = n28507 & ~n28716;
  assign n28718 = ~n28513 & n28520;
  assign n28719 = ~n28526 & n28718;
  assign n28720 = ~n28532 & n28719;
  assign n28721 = ~n28543 & n28720;
  assign n28722 = n28513 & n28543;
  assign n28723 = n28584 & n28722;
  assign n28724 = ~n28544 & ~n28723;
  assign n28725 = ~n28546 & ~n28576;
  assign n28726 = n28513 & n28563;
  assign n28727 = n28725 & ~n28726;
  assign n28728 = ~n28543 & ~n28727;
  assign n28729 = n28543 & n28550;
  assign n28730 = n28568 & ~n28729;
  assign n28731 = ~n28728 & n28730;
  assign n28732 = n28724 & n28731;
  assign n28733 = ~n28507 & ~n28732;
  assign n28734 = ~n28721 & ~n28733;
  assign n28735 = ~n28717 & n28734;
  assign n28736 = n28576 & n28722;
  assign n28737 = ~n28513 & n28578;
  assign n28738 = ~n28736 & ~n28737;
  assign n28739 = n28543 & n28708;
  assign n28740 = n28738 & ~n28739;
  assign n28741 = n28735 & n28740;
  assign n28742 = ~pi0490 & ~n28741;
  assign n28743 = pi0490 & n28740;
  assign n28744 = n28734 & n28743;
  assign n28745 = ~n28717 & n28744;
  assign po0516 = n28742 | n28745;
  assign n28747 = pi3392 & pi9040;
  assign n28748 = pi3419 & ~pi9040;
  assign n28749 = ~n28747 & ~n28748;
  assign n28750 = pi0477 & n28749;
  assign n28751 = ~pi0477 & ~n28749;
  assign n28752 = ~n28750 & ~n28751;
  assign n28753 = pi3407 & pi9040;
  assign n28754 = pi3406 & ~pi9040;
  assign n28755 = ~n28753 & ~n28754;
  assign n28756 = pi0456 & n28755;
  assign n28757 = ~pi0456 & ~n28755;
  assign n28758 = ~n28756 & ~n28757;
  assign n28759 = pi3379 & pi9040;
  assign n28760 = pi3363 & ~pi9040;
  assign n28761 = ~n28759 & ~n28760;
  assign n28762 = ~pi0457 & ~n28761;
  assign n28763 = pi0457 & n28761;
  assign n28764 = ~n28762 & ~n28763;
  assign n28765 = pi3406 & pi9040;
  assign n28766 = pi3379 & ~pi9040;
  assign n28767 = ~n28765 & ~n28766;
  assign n28768 = ~pi0461 & n28767;
  assign n28769 = pi0461 & ~n28767;
  assign n28770 = ~n28768 & ~n28769;
  assign n28771 = pi3413 & pi9040;
  assign n28772 = pi3371 & ~pi9040;
  assign n28773 = ~n28771 & ~n28772;
  assign n28774 = ~pi0450 & n28773;
  assign n28775 = pi0450 & ~n28773;
  assign n28776 = ~n28774 & ~n28775;
  assign n28777 = n28770 & ~n28776;
  assign n28778 = ~n28764 & n28777;
  assign n28779 = n28758 & n28778;
  assign n28780 = ~n28770 & n28776;
  assign n28781 = ~n28764 & n28780;
  assign n28782 = n28770 & n28776;
  assign n28783 = n28764 & n28782;
  assign n28784 = n28758 & n28783;
  assign n28785 = ~n28781 & ~n28784;
  assign n28786 = ~n28779 & n28785;
  assign n28787 = n28752 & ~n28786;
  assign n28788 = n28764 & n28770;
  assign n28789 = ~n28758 & n28788;
  assign n28790 = n28764 & ~n28770;
  assign n28791 = n28758 & n28790;
  assign n28792 = ~n28789 & ~n28791;
  assign n28793 = ~n28752 & ~n28792;
  assign n28794 = ~n28787 & ~n28793;
  assign n28795 = ~pi3361 & pi9040;
  assign n28796 = pi3407 & ~pi9040;
  assign n28797 = ~n28795 & ~n28796;
  assign n28798 = pi0443 & n28797;
  assign n28799 = ~pi0443 & ~n28797;
  assign n28800 = ~n28798 & ~n28799;
  assign n28801 = n28764 & n28777;
  assign n28802 = ~n28758 & ~n28764;
  assign n28803 = ~n28776 & n28802;
  assign n28804 = ~n28770 & n28803;
  assign n28805 = ~n28801 & ~n28804;
  assign n28806 = ~n28752 & ~n28805;
  assign n28807 = n28776 & n28802;
  assign n28808 = n28770 & n28807;
  assign n28809 = ~n28779 & ~n28808;
  assign n28810 = n28758 & ~n28764;
  assign n28811 = ~n28770 & n28810;
  assign n28812 = ~n28770 & ~n28776;
  assign n28813 = n28764 & n28812;
  assign n28814 = ~n28758 & n28813;
  assign n28815 = ~n28811 & ~n28814;
  assign n28816 = n28752 & ~n28815;
  assign n28817 = n28809 & ~n28816;
  assign n28818 = ~n28806 & n28817;
  assign n28819 = n28800 & ~n28818;
  assign n28820 = ~n28752 & ~n28758;
  assign n28821 = n28777 & n28820;
  assign n28822 = n28764 & n28780;
  assign n28823 = n28776 & n28810;
  assign n28824 = n28770 & n28823;
  assign n28825 = ~n28822 & ~n28824;
  assign n28826 = n28758 & n28812;
  assign n28827 = n28825 & ~n28826;
  assign n28828 = ~n28752 & ~n28827;
  assign n28829 = ~n28764 & ~n28770;
  assign n28830 = n28752 & ~n28758;
  assign n28831 = n28829 & n28830;
  assign n28832 = ~n28770 & n28807;
  assign n28833 = ~n28831 & ~n28832;
  assign n28834 = ~n28828 & n28833;
  assign n28835 = ~n28821 & n28834;
  assign n28836 = ~n28758 & n28801;
  assign n28837 = n28764 & ~n28776;
  assign n28838 = n28758 & n28837;
  assign n28839 = ~n28770 & n28838;
  assign n28840 = ~n28836 & ~n28839;
  assign n28841 = n28835 & n28840;
  assign n28842 = ~n28800 & ~n28841;
  assign n28843 = ~n28764 & n28776;
  assign n28844 = n28752 & n28843;
  assign n28845 = ~n28758 & n28844;
  assign n28846 = ~n28842 & ~n28845;
  assign n28847 = ~n28819 & n28846;
  assign n28848 = n28794 & n28847;
  assign n28849 = ~pi0485 & ~n28848;
  assign n28850 = pi0485 & n28848;
  assign po0517 = n28849 | n28850;
  assign n28852 = n28420 & n28433;
  assign n28853 = ~n28457 & ~n28852;
  assign n28854 = ~n28470 & n28853;
  assign n28855 = n28406 & ~n28854;
  assign n28856 = ~n28420 & n28441;
  assign n28857 = n28485 & n28856;
  assign n28858 = ~n28420 & n28477;
  assign n28859 = ~n28426 & ~n28432;
  assign n28860 = ~n28442 & ~n28859;
  assign n28861 = n28420 & ~n28860;
  assign n28862 = ~n28858 & ~n28861;
  assign n28863 = ~n28857 & n28862;
  assign n28864 = ~n28406 & ~n28863;
  assign n28865 = ~n28855 & ~n28864;
  assign n28866 = n28412 & ~n28865;
  assign n28867 = ~n28432 & n28467;
  assign n28868 = ~n28420 & n28426;
  assign n28869 = n28432 & n28868;
  assign n28870 = ~n28852 & ~n28869;
  assign n28871 = ~n28406 & ~n28870;
  assign n28872 = ~n28483 & ~n28871;
  assign n28873 = ~n28420 & n28443;
  assign n28874 = ~n28487 & ~n28873;
  assign n28875 = n28406 & n28420;
  assign n28876 = n28485 & n28875;
  assign n28877 = n28406 & n28462;
  assign n28878 = ~n28876 & ~n28877;
  assign n28879 = n28874 & n28878;
  assign n28880 = n28872 & n28879;
  assign n28881 = ~n28867 & n28880;
  assign n28882 = ~n28412 & ~n28881;
  assign n28883 = n28472 & n28482;
  assign n28884 = n28426 & n28483;
  assign n28885 = ~n28883 & ~n28884;
  assign n28886 = n28406 & n28490;
  assign n28887 = n28885 & ~n28886;
  assign n28888 = n28420 & n28445;
  assign n28889 = ~n28420 & n28453;
  assign n28890 = ~n28888 & ~n28889;
  assign n28891 = n28406 & ~n28890;
  assign n28892 = n28887 & ~n28891;
  assign n28893 = ~n28882 & n28892;
  assign n28894 = ~n28866 & n28893;
  assign n28895 = ~pi0496 & ~n28894;
  assign n28896 = pi0496 & n28894;
  assign po0518 = n28895 | n28896;
  assign n28898 = pi3384 & pi9040;
  assign n28899 = pi3394 & ~pi9040;
  assign n28900 = ~n28898 & ~n28899;
  assign n28901 = ~pi0478 & n28900;
  assign n28902 = pi0478 & ~n28900;
  assign n28903 = ~n28901 & ~n28902;
  assign n28904 = pi3369 & pi9040;
  assign n28905 = pi3408 & ~pi9040;
  assign n28906 = ~n28904 & ~n28905;
  assign n28907 = ~pi0466 & ~n28906;
  assign n28908 = pi0466 & ~n28904;
  assign n28909 = ~n28905 & n28908;
  assign n28910 = ~n28907 & ~n28909;
  assign n28911 = pi3456 & pi9040;
  assign n28912 = pi3365 & ~pi9040;
  assign n28913 = ~n28911 & ~n28912;
  assign n28914 = pi0455 & n28913;
  assign n28915 = ~pi0455 & ~n28913;
  assign n28916 = ~n28914 & ~n28915;
  assign n28917 = n28910 & ~n28916;
  assign n28918 = pi3365 & pi9040;
  assign n28919 = pi3452 & ~pi9040;
  assign n28920 = ~n28918 & ~n28919;
  assign n28921 = pi0474 & n28920;
  assign n28922 = ~pi0474 & ~n28920;
  assign n28923 = ~n28921 & ~n28922;
  assign n28924 = pi3416 & pi9040;
  assign n28925 = pi3389 & ~pi9040;
  assign n28926 = ~n28924 & ~n28925;
  assign n28927 = pi0448 & n28926;
  assign n28928 = ~pi0448 & ~n28926;
  assign n28929 = ~n28927 & ~n28928;
  assign n28930 = n28923 & n28929;
  assign n28931 = n28917 & n28930;
  assign n28932 = n28923 & ~n28929;
  assign n28933 = ~n28910 & n28932;
  assign n28934 = ~n28931 & ~n28933;
  assign n28935 = n28903 & ~n28934;
  assign n28936 = pi3388 & pi9040;
  assign n28937 = pi3390 & ~pi9040;
  assign n28938 = ~n28936 & ~n28937;
  assign n28939 = pi0460 & n28938;
  assign n28940 = ~pi0460 & ~n28938;
  assign n28941 = ~n28939 & ~n28940;
  assign n28942 = ~n28903 & ~n28923;
  assign n28943 = n28910 & n28942;
  assign n28944 = n28917 & ~n28929;
  assign n28945 = n28910 & n28916;
  assign n28946 = n28929 & n28945;
  assign n28947 = ~n28944 & ~n28946;
  assign n28948 = ~n28910 & ~n28916;
  assign n28949 = n28929 & n28948;
  assign n28950 = n28923 & n28949;
  assign n28951 = n28947 & ~n28950;
  assign n28952 = ~n28903 & ~n28951;
  assign n28953 = ~n28943 & ~n28952;
  assign n28954 = ~n28910 & n28916;
  assign n28955 = ~n28929 & n28954;
  assign n28956 = n28923 & n28955;
  assign n28957 = n28953 & ~n28956;
  assign n28958 = ~n28923 & n28948;
  assign n28959 = ~n28910 & n28929;
  assign n28960 = n28916 & n28959;
  assign n28961 = ~n28958 & ~n28960;
  assign n28962 = n28903 & ~n28961;
  assign n28963 = ~n28929 & n28945;
  assign n28964 = ~n28923 & n28963;
  assign n28965 = ~n28962 & ~n28964;
  assign n28966 = n28957 & n28965;
  assign n28967 = n28941 & ~n28966;
  assign n28968 = ~n28935 & ~n28967;
  assign n28969 = ~n28903 & ~n28941;
  assign n28970 = ~n28961 & n28969;
  assign n28971 = ~n28929 & n28948;
  assign n28972 = ~n28963 & ~n28971;
  assign n28973 = n28923 & ~n28972;
  assign n28974 = ~n28931 & ~n28973;
  assign n28975 = ~n28941 & ~n28974;
  assign n28976 = ~n28970 & ~n28975;
  assign n28977 = n28903 & ~n28941;
  assign n28978 = n28917 & ~n28923;
  assign n28979 = ~n28955 & ~n28978;
  assign n28980 = n28910 & n28929;
  assign n28981 = n28979 & ~n28980;
  assign n28982 = n28977 & ~n28981;
  assign n28983 = n28976 & ~n28982;
  assign n28984 = n28968 & n28983;
  assign n28985 = ~pi0482 & ~n28984;
  assign n28986 = pi0482 & n28976;
  assign n28987 = n28968 & n28986;
  assign n28988 = ~n28982 & n28987;
  assign po0519 = n28985 | n28988;
  assign n28990 = n28612 & n28649;
  assign n28991 = ~n28612 & n28669;
  assign n28992 = ~n28990 & ~n28991;
  assign n28993 = n28640 & ~n28992;
  assign n28994 = ~n28640 & n28681;
  assign n28995 = ~n28681 & ~n28686;
  assign n28996 = ~n28625 & n28679;
  assign n28997 = ~n28678 & ~n28996;
  assign n28998 = ~n28640 & ~n28997;
  assign n28999 = ~n28612 & ~n28640;
  assign n29000 = n28648 & n28999;
  assign n29001 = n28618 & n29000;
  assign n29002 = ~n28612 & ~n28618;
  assign n29003 = ~n28631 & n29002;
  assign n29004 = n28625 & n29003;
  assign n29005 = n28618 & n28640;
  assign n29006 = ~n28631 & n29005;
  assign n29007 = ~n28625 & n29006;
  assign n29008 = ~n29004 & ~n29007;
  assign n29009 = ~n29001 & n29008;
  assign n29010 = ~n28998 & n29009;
  assign n29011 = n28995 & n29010;
  assign n29012 = n28606 & ~n29011;
  assign n29013 = n28612 & n28686;
  assign n29014 = ~n29012 & ~n29013;
  assign n29015 = ~n28994 & n29014;
  assign n29016 = ~n28993 & n29015;
  assign n29017 = ~n28618 & ~n28625;
  assign n29018 = n28683 & n29017;
  assign n29019 = ~n28650 & ~n29018;
  assign n29020 = n28640 & n28672;
  assign n29021 = n28612 & n28695;
  assign n29022 = ~n29020 & ~n29021;
  assign n29023 = ~n28612 & n28658;
  assign n29024 = ~n28990 & ~n29023;
  assign n29025 = ~n28612 & n28655;
  assign n29026 = n28618 & ~n28631;
  assign n29027 = ~n29025 & ~n29026;
  assign n29028 = ~n28640 & ~n29027;
  assign n29029 = n29024 & ~n29028;
  assign n29030 = n29022 & n29029;
  assign n29031 = n29019 & n29030;
  assign n29032 = ~n28606 & ~n29031;
  assign n29033 = n29016 & ~n29032;
  assign n29034 = ~pi0487 & ~n29033;
  assign n29035 = pi0487 & n29016;
  assign n29036 = ~n29032 & n29035;
  assign po0521 = n29034 | n29036;
  assign n29038 = n28916 & n28929;
  assign n29039 = ~n28910 & n29038;
  assign n29040 = n28923 & n29039;
  assign n29041 = ~n28923 & n28955;
  assign n29042 = ~n29040 & ~n29041;
  assign n29043 = n28903 & ~n29042;
  assign n29044 = n28903 & n28923;
  assign n29045 = ~n28948 & ~n28963;
  assign n29046 = n29044 & ~n29045;
  assign n29047 = n28903 & ~n28929;
  assign n29048 = n28948 & n29047;
  assign n29049 = ~n29046 & ~n29048;
  assign n29050 = n28941 & ~n29049;
  assign n29051 = ~n28923 & n28929;
  assign n29052 = n28916 & n29051;
  assign n29053 = n28910 & n29052;
  assign n29054 = ~n28980 & ~n29051;
  assign n29055 = ~n28903 & ~n29054;
  assign n29056 = ~n28923 & ~n28929;
  assign n29057 = ~n28916 & n29056;
  assign n29058 = n28910 & n29057;
  assign n29059 = ~n29055 & ~n29058;
  assign n29060 = ~n29053 & n29059;
  assign n29061 = n28941 & ~n29060;
  assign n29062 = ~n29050 & ~n29061;
  assign n29063 = ~n28903 & n28923;
  assign n29064 = n28945 & n29063;
  assign n29065 = ~n28929 & n29064;
  assign n29066 = ~n28917 & ~n28980;
  assign n29067 = n28923 & ~n29066;
  assign n29068 = ~n28955 & ~n29067;
  assign n29069 = n28903 & ~n29068;
  assign n29070 = n28916 & ~n28923;
  assign n29071 = n28903 & n29070;
  assign n29072 = ~n28929 & n29071;
  assign n29073 = ~n29040 & ~n29072;
  assign n29074 = ~n28916 & n28929;
  assign n29075 = ~n28955 & ~n29074;
  assign n29076 = ~n28923 & ~n29075;
  assign n29077 = n29073 & ~n29076;
  assign n29078 = ~n29069 & n29077;
  assign n29079 = ~n29065 & n29078;
  assign n29080 = ~n28941 & ~n29079;
  assign n29081 = n28923 & n28971;
  assign n29082 = ~n28923 & n28980;
  assign n29083 = ~n29081 & ~n29082;
  assign n29084 = ~n28903 & ~n29083;
  assign n29085 = ~n29080 & ~n29084;
  assign n29086 = n29062 & n29085;
  assign n29087 = ~n29043 & n29086;
  assign n29088 = pi0492 & n29087;
  assign n29089 = ~pi0492 & ~n29087;
  assign po0522 = n29088 | n29089;
  assign n29091 = ~n29013 & ~n29018;
  assign n29092 = ~n28669 & ~n28681;
  assign n29093 = ~n29025 & n29092;
  assign n29094 = ~n28640 & ~n29093;
  assign n29095 = ~n28612 & n28643;
  assign n29096 = ~n29004 & ~n29095;
  assign n29097 = ~n28697 & n29096;
  assign n29098 = n28640 & n28658;
  assign n29099 = n29097 & ~n29098;
  assign n29100 = ~n29094 & n29099;
  assign n29101 = n28606 & ~n29100;
  assign n29102 = n28612 & n28651;
  assign n29103 = n28625 & n28664;
  assign n29104 = ~n28669 & ~n29103;
  assign n29105 = n28640 & ~n29104;
  assign n29106 = ~n29102 & ~n29105;
  assign n29107 = n28641 & n28670;
  assign n29108 = ~n28640 & n28649;
  assign n29109 = ~n29107 & ~n29108;
  assign n29110 = n29106 & n29109;
  assign n29111 = n28625 & n28679;
  assign n29112 = ~n28990 & ~n29111;
  assign n29113 = ~n29023 & n29112;
  assign n29114 = n29110 & n29113;
  assign n29115 = ~n28606 & ~n29114;
  assign n29116 = ~n28990 & n29096;
  assign n29117 = ~n28640 & ~n29116;
  assign n29118 = ~n29115 & ~n29117;
  assign n29119 = ~n29101 & n29118;
  assign n29120 = n29091 & n29119;
  assign n29121 = pi0504 & ~n29120;
  assign n29122 = ~pi0504 & n29120;
  assign po0523 = n29121 | n29122;
  assign n29124 = n28513 & n28706;
  assign n29125 = ~n28564 & ~n28572;
  assign n29126 = ~n28513 & n28533;
  assign n29127 = n28513 & n28584;
  assign n29128 = ~n29126 & ~n29127;
  assign n29129 = n29125 & n29128;
  assign n29130 = ~n28543 & ~n29129;
  assign n29131 = ~n28513 & n28545;
  assign n29132 = ~n28544 & ~n29131;
  assign n29133 = ~n28566 & n29132;
  assign n29134 = n28543 & ~n29133;
  assign n29135 = ~n28513 & ~n28526;
  assign n29136 = n28532 & n29135;
  assign n29137 = n28520 & n29136;
  assign n29138 = ~n29134 & ~n29137;
  assign n29139 = ~n29130 & n29138;
  assign n29140 = ~n29124 & n29139;
  assign n29141 = ~n28507 & ~n29140;
  assign n29142 = ~n28513 & ~n28543;
  assign n29143 = n28550 & n29142;
  assign n29144 = ~n28543 & n28566;
  assign n29145 = ~n28543 & n28576;
  assign n29146 = ~n29144 & ~n29145;
  assign n29147 = n28513 & ~n29146;
  assign n29148 = ~n29143 & ~n29147;
  assign n29149 = n28513 & n28534;
  assign n29150 = ~n28720 & ~n29149;
  assign n29151 = ~n28513 & n28563;
  assign n29152 = n28513 & n28545;
  assign n29153 = ~n29151 & ~n29152;
  assign n29154 = ~n28534 & n29153;
  assign n29155 = ~n28564 & n29154;
  assign n29156 = n28543 & ~n29155;
  assign n29157 = n28513 & n28546;
  assign n29158 = ~n29156 & ~n29157;
  assign n29159 = n29150 & n29158;
  assign n29160 = n29148 & n29159;
  assign n29161 = n28507 & ~n29160;
  assign n29162 = ~n28543 & ~n28709;
  assign n29163 = ~n29161 & ~n29162;
  assign n29164 = ~n28567 & ~n29149;
  assign n29165 = n28543 & ~n29164;
  assign n29166 = n29163 & ~n29165;
  assign n29167 = ~n29141 & n29166;
  assign n29168 = pi0511 & ~n29167;
  assign n29169 = ~pi0511 & n29167;
  assign po0524 = n29168 | n29169;
  assign n29171 = n28758 & n28781;
  assign n29172 = ~n28790 & ~n28808;
  assign n29173 = n28752 & ~n29172;
  assign n29174 = ~n29171 & ~n29173;
  assign n29175 = ~n28804 & n29174;
  assign n29176 = ~n28752 & n28758;
  assign n29177 = n28778 & n29176;
  assign n29178 = ~n28836 & ~n29177;
  assign n29179 = ~n28784 & n29178;
  assign n29180 = n29175 & n29179;
  assign n29181 = n28800 & ~n29180;
  assign n29182 = ~n28764 & n28812;
  assign n29183 = n28758 & n29182;
  assign n29184 = ~n28824 & ~n29183;
  assign n29185 = n28752 & n28778;
  assign n29186 = n28758 & n28801;
  assign n29187 = ~n29185 & ~n29186;
  assign n29188 = n28758 & ~n28770;
  assign n29189 = ~n28837 & ~n29188;
  assign n29190 = ~n28843 & n29189;
  assign n29191 = ~n28752 & ~n29190;
  assign n29192 = ~n28758 & n28783;
  assign n29193 = ~n28832 & ~n29192;
  assign n29194 = ~n29191 & n29193;
  assign n29195 = n29187 & n29194;
  assign n29196 = n29184 & n29195;
  assign n29197 = ~n28800 & ~n29196;
  assign n29198 = ~n29181 & ~n29197;
  assign n29199 = pi0481 & ~n29198;
  assign n29200 = ~pi0481 & ~n29181;
  assign n29201 = ~n29197 & n29200;
  assign po0525 = n29199 | n29201;
  assign n29203 = ~n28472 & ~n28477;
  assign n29204 = ~n28406 & ~n29203;
  assign n29205 = n28420 & n28457;
  assign n29206 = ~n29204 & ~n29205;
  assign n29207 = n28420 & n28432;
  assign n29208 = ~n28485 & ~n29207;
  assign n29209 = ~n28453 & n29208;
  assign n29210 = n28406 & ~n29209;
  assign n29211 = n29206 & ~n29210;
  assign n29212 = ~n28412 & ~n29211;
  assign n29213 = ~n28420 & n28486;
  assign n29214 = ~n28406 & n29213;
  assign n29215 = ~n28884 & ~n29214;
  assign n29216 = ~n28886 & n29215;
  assign n29217 = n28406 & n28432;
  assign n29218 = n28868 & n29217;
  assign n29219 = n28420 & n28477;
  assign n29220 = ~n28406 & n28485;
  assign n29221 = ~n29219 & ~n29220;
  assign n29222 = ~n28484 & n29221;
  assign n29223 = ~n29218 & n29222;
  assign n29224 = ~n28441 & n28868;
  assign n29225 = ~n28490 & ~n29224;
  assign n29226 = n29223 & n29225;
  assign n29227 = ~n28877 & n29226;
  assign n29228 = n28412 & ~n29227;
  assign n29229 = n29216 & ~n29228;
  assign n29230 = ~n29212 & n29229;
  assign n29231 = ~pi0503 & ~n29230;
  assign n29232 = pi0503 & n29216;
  assign n29233 = ~n29212 & n29232;
  assign n29234 = ~n29228 & n29233;
  assign po0526 = n29231 | n29234;
  assign n29236 = ~n28331 & n28361;
  assign n29237 = n28331 & n28372;
  assign n29238 = ~n28358 & ~n29237;
  assign n29239 = ~n28305 & ~n29238;
  assign n29240 = ~n29236 & ~n29239;
  assign n29241 = n28305 & ~n28331;
  assign n29242 = ~n28323 & n29241;
  assign n29243 = ~n28317 & n29242;
  assign n29244 = n28339 & n28373;
  assign n29245 = ~n29243 & ~n29244;
  assign n29246 = n28305 & n28380;
  assign n29247 = n29245 & ~n29246;
  assign n29248 = ~n28335 & ~n28347;
  assign n29249 = n28323 & n28337;
  assign n29250 = n29248 & ~n29249;
  assign n29251 = n29247 & n29250;
  assign n29252 = n29240 & n29251;
  assign n29253 = n28370 & ~n29252;
  assign n29254 = ~n28334 & ~n28358;
  assign n29255 = n28331 & ~n29254;
  assign n29256 = ~n28317 & n28376;
  assign n29257 = ~n28387 & ~n29256;
  assign n29258 = ~n28311 & ~n28323;
  assign n29259 = n28331 & n29258;
  assign n29260 = n29257 & ~n29259;
  assign n29261 = ~n28305 & ~n29260;
  assign n29262 = ~n28331 & n28357;
  assign n29263 = ~n28317 & n28346;
  assign n29264 = ~n29262 & ~n29263;
  assign n29265 = n28305 & ~n29264;
  assign n29266 = ~n28331 & n28340;
  assign n29267 = ~n29265 & ~n29266;
  assign n29268 = ~n29261 & n29267;
  assign n29269 = ~n29255 & n29268;
  assign n29270 = ~n28370 & ~n29269;
  assign n29271 = ~n28305 & n28377;
  assign n29272 = ~n29270 & ~n29271;
  assign n29273 = n28352 & n29241;
  assign n29274 = ~n28323 & n29273;
  assign n29275 = n29272 & ~n29274;
  assign n29276 = ~n29253 & n29275;
  assign n29277 = ~pi0493 & ~n29276;
  assign n29278 = pi0493 & n29272;
  assign n29279 = ~n29253 & n29278;
  assign n29280 = ~n29274 & n29279;
  assign po0527 = n29277 | n29280;
  assign n29282 = pi3382 & pi9040;
  assign n29283 = pi3457 & ~pi9040;
  assign n29284 = ~n29282 & ~n29283;
  assign n29285 = pi0455 & n29284;
  assign n29286 = ~pi0455 & ~n29284;
  assign n29287 = ~n29285 & ~n29286;
  assign n29288 = pi3362 & pi9040;
  assign n29289 = pi3416 & ~pi9040;
  assign n29290 = ~n29288 & ~n29289;
  assign n29291 = ~pi0460 & n29290;
  assign n29292 = pi0460 & ~n29290;
  assign n29293 = ~n29291 & ~n29292;
  assign n29294 = pi3408 & pi9040;
  assign n29295 = pi3367 & ~pi9040;
  assign n29296 = ~n29294 & ~n29295;
  assign n29297 = ~pi0467 & n29296;
  assign n29298 = pi0467 & ~n29296;
  assign n29299 = ~n29297 & ~n29298;
  assign n29300 = ~n29293 & ~n29299;
  assign n29301 = n29287 & n29300;
  assign n29302 = ~pi0467 & ~n29296;
  assign n29303 = pi0467 & n29296;
  assign n29304 = ~n29302 & ~n29303;
  assign n29305 = ~n29293 & ~n29304;
  assign n29306 = ~n29287 & n29305;
  assign n29307 = ~n29301 & ~n29306;
  assign n29308 = pi3455 & pi9040;
  assign n29309 = pi3391 & ~pi9040;
  assign n29310 = ~n29308 & ~n29309;
  assign n29311 = pi0464 & n29310;
  assign n29312 = ~pi0464 & ~n29310;
  assign n29313 = ~n29311 & ~n29312;
  assign n29314 = n29287 & ~n29313;
  assign n29315 = n29304 & n29314;
  assign n29316 = n29307 & ~n29315;
  assign n29317 = pi3397 & pi9040;
  assign n29318 = pi3366 & ~pi9040;
  assign n29319 = ~n29317 & ~n29318;
  assign n29320 = pi0446 & n29319;
  assign n29321 = ~pi0446 & ~n29319;
  assign n29322 = ~n29320 & ~n29321;
  assign n29323 = pi3390 & pi9040;
  assign n29324 = pi3369 & ~pi9040;
  assign n29325 = ~n29323 & ~n29324;
  assign n29326 = ~pi0472 & n29325;
  assign n29327 = pi0472 & ~n29325;
  assign n29328 = ~n29326 & ~n29327;
  assign n29329 = ~n29322 & ~n29328;
  assign n29330 = ~n29316 & n29329;
  assign n29331 = n29293 & ~n29304;
  assign n29332 = n29287 & n29331;
  assign n29333 = ~n29328 & n29332;
  assign n29334 = n29313 & n29333;
  assign n29335 = n29287 & n29305;
  assign n29336 = n29322 & n29335;
  assign n29337 = ~n29287 & n29304;
  assign n29338 = n29293 & ~n29299;
  assign n29339 = n29313 & n29338;
  assign n29340 = ~n29337 & ~n29339;
  assign n29341 = n29322 & ~n29340;
  assign n29342 = ~n29336 & ~n29341;
  assign n29343 = ~n29328 & ~n29342;
  assign n29344 = ~n29334 & ~n29343;
  assign n29345 = ~n29287 & n29313;
  assign n29346 = n29304 & n29345;
  assign n29347 = ~n29287 & ~n29313;
  assign n29348 = ~n29304 & n29347;
  assign n29349 = n29293 & n29348;
  assign n29350 = ~n29346 & ~n29349;
  assign n29351 = n29322 & ~n29350;
  assign n29352 = n29344 & ~n29351;
  assign n29353 = n29313 & ~n29322;
  assign n29354 = n29338 & n29353;
  assign n29355 = n29287 & n29354;
  assign n29356 = ~n29300 & ~n29331;
  assign n29357 = n29314 & ~n29356;
  assign n29358 = ~n29293 & n29348;
  assign n29359 = ~n29357 & ~n29358;
  assign n29360 = ~n29287 & n29338;
  assign n29361 = ~n29313 & ~n29322;
  assign n29362 = n29360 & n29361;
  assign n29363 = n29345 & ~n29356;
  assign n29364 = n29313 & n29335;
  assign n29365 = ~n29363 & ~n29364;
  assign n29366 = ~n29362 & n29365;
  assign n29367 = n29359 & n29366;
  assign n29368 = ~n29355 & n29367;
  assign n29369 = ~n29313 & n29322;
  assign n29370 = n29287 & n29369;
  assign n29371 = n29293 & n29370;
  assign n29372 = n29368 & ~n29371;
  assign n29373 = n29328 & ~n29372;
  assign n29374 = n29352 & ~n29373;
  assign n29375 = ~n29330 & n29374;
  assign n29376 = ~pi0500 & ~n29375;
  assign n29377 = pi0500 & n29352;
  assign n29378 = ~n29330 & n29377;
  assign n29379 = ~n29373 & n29378;
  assign po0529 = n29376 | n29379;
  assign n29381 = n29287 & n29338;
  assign n29382 = n29322 & n29381;
  assign n29383 = ~n29313 & n29382;
  assign n29384 = n29305 & n29369;
  assign n29385 = ~n29287 & n29384;
  assign n29386 = ~n29383 & ~n29385;
  assign n29387 = ~n29358 & ~n29362;
  assign n29388 = ~n29293 & n29313;
  assign n29389 = n29287 & n29388;
  assign n29390 = ~n29339 & ~n29389;
  assign n29391 = n29322 & ~n29390;
  assign n29392 = ~n29322 & ~n29347;
  assign n29393 = ~n29356 & n29392;
  assign n29394 = ~n29287 & ~n29338;
  assign n29395 = n29322 & n29394;
  assign n29396 = ~n29313 & n29395;
  assign n29397 = ~n29393 & ~n29396;
  assign n29398 = ~n29391 & n29397;
  assign n29399 = n29387 & n29398;
  assign n29400 = ~n29328 & ~n29399;
  assign n29401 = n29386 & ~n29400;
  assign n29402 = n29301 & ~n29322;
  assign n29403 = n29313 & n29402;
  assign n29404 = ~n29322 & n29328;
  assign n29405 = n29347 & ~n29356;
  assign n29406 = ~n29339 & ~n29405;
  assign n29407 = ~n29335 & n29406;
  assign n29408 = n29404 & ~n29407;
  assign n29409 = n29306 & n29313;
  assign n29410 = ~n29287 & n29388;
  assign n29411 = n29313 & n29331;
  assign n29412 = ~n29410 & ~n29411;
  assign n29413 = ~n29313 & n29338;
  assign n29414 = ~n29332 & ~n29413;
  assign n29415 = n29412 & n29414;
  assign n29416 = n29322 & ~n29415;
  assign n29417 = ~n29409 & ~n29416;
  assign n29418 = n29328 & ~n29417;
  assign n29419 = ~n29408 & ~n29418;
  assign n29420 = ~n29403 & n29419;
  assign n29421 = n29401 & n29420;
  assign n29422 = pi0501 & ~n29421;
  assign n29423 = ~pi0501 & n29401;
  assign n29424 = n29420 & n29423;
  assign po0530 = n29422 | n29424;
  assign n29426 = ~n29332 & ~n29388;
  assign n29427 = n29329 & ~n29426;
  assign n29428 = n29287 & n29313;
  assign n29429 = ~n29300 & n29428;
  assign n29430 = ~n29328 & n29429;
  assign n29431 = n29322 & n29345;
  assign n29432 = n29300 & n29431;
  assign n29433 = n29287 & n29353;
  assign n29434 = ~n29304 & n29433;
  assign n29435 = ~n29432 & ~n29434;
  assign n29436 = ~n29430 & n29435;
  assign n29437 = ~n29411 & ~n29413;
  assign n29438 = n29322 & ~n29437;
  assign n29439 = ~n29385 & ~n29438;
  assign n29440 = ~n29328 & ~n29439;
  assign n29441 = ~n29287 & ~n29293;
  assign n29442 = ~n29300 & ~n29441;
  assign n29443 = ~n29313 & ~n29442;
  assign n29444 = ~n29381 & ~n29443;
  assign n29445 = ~n29322 & ~n29444;
  assign n29446 = ~n29405 & ~n29445;
  assign n29447 = n29313 & n29360;
  assign n29448 = ~n29304 & n29314;
  assign n29449 = n29313 & ~n29442;
  assign n29450 = ~n29448 & ~n29449;
  assign n29451 = n29322 & ~n29450;
  assign n29452 = ~n29447 & ~n29451;
  assign n29453 = n29446 & n29452;
  assign n29454 = n29328 & ~n29453;
  assign n29455 = ~n29440 & ~n29454;
  assign n29456 = n29436 & n29455;
  assign n29457 = ~n29427 & n29456;
  assign n29458 = pi0508 & ~n29457;
  assign n29459 = ~pi0508 & n29436;
  assign n29460 = ~n29427 & n29459;
  assign n29461 = n29455 & n29460;
  assign po0531 = n29458 | n29461;
  assign n29463 = pi3457 & pi9040;
  assign n29464 = pi3374 & ~pi9040;
  assign n29465 = ~n29463 & ~n29464;
  assign n29466 = ~pi0470 & n29465;
  assign n29467 = pi0470 & ~n29465;
  assign n29468 = ~n29466 & ~n29467;
  assign n29469 = pi3389 & pi9040;
  assign n29470 = pi3456 & ~pi9040;
  assign n29471 = ~n29469 & ~n29470;
  assign n29472 = ~pi0448 & n29471;
  assign n29473 = pi0448 & ~n29471;
  assign n29474 = ~n29472 & ~n29473;
  assign n29475 = pi3391 & pi9040;
  assign n29476 = pi3378 & ~pi9040;
  assign n29477 = ~n29475 & ~n29476;
  assign n29478 = pi0473 & n29477;
  assign n29479 = ~pi0473 & ~n29477;
  assign n29480 = ~n29478 & ~n29479;
  assign n29481 = pi3394 & pi9040;
  assign n29482 = pi3410 & ~pi9040;
  assign n29483 = ~n29481 & ~n29482;
  assign n29484 = pi0451 & n29483;
  assign n29485 = ~pi0451 & ~n29483;
  assign n29486 = ~n29484 & ~n29485;
  assign n29487 = n29480 & ~n29486;
  assign n29488 = n29474 & n29487;
  assign n29489 = pi3420 & pi9040;
  assign n29490 = pi3382 & ~pi9040;
  assign n29491 = ~n29489 & ~n29490;
  assign n29492 = pi0479 & n29491;
  assign n29493 = ~pi0479 & ~n29491;
  assign n29494 = ~n29492 & ~n29493;
  assign n29495 = n29480 & n29494;
  assign n29496 = ~n29474 & n29495;
  assign n29497 = n29486 & n29496;
  assign n29498 = ~n29488 & ~n29497;
  assign n29499 = ~n29474 & ~n29494;
  assign n29500 = ~n29480 & n29499;
  assign n29501 = n29486 & n29500;
  assign n29502 = n29498 & ~n29501;
  assign n29503 = n29468 & ~n29502;
  assign n29504 = pi3374 & pi9040;
  assign n29505 = pi3384 & ~pi9040;
  assign n29506 = ~n29504 & ~n29505;
  assign n29507 = ~pi0466 & ~n29506;
  assign n29508 = pi0466 & n29506;
  assign n29509 = ~n29507 & ~n29508;
  assign n29510 = ~n29468 & n29486;
  assign n29511 = n29499 & n29510;
  assign n29512 = n29480 & n29511;
  assign n29513 = ~n29468 & ~n29486;
  assign n29514 = ~n29474 & n29494;
  assign n29515 = n29513 & n29514;
  assign n29516 = n29474 & n29494;
  assign n29517 = n29480 & n29516;
  assign n29518 = ~n29468 & n29517;
  assign n29519 = n29486 & n29518;
  assign n29520 = n29480 & ~n29494;
  assign n29521 = n29474 & n29520;
  assign n29522 = ~n29486 & n29521;
  assign n29523 = ~n29519 & ~n29522;
  assign n29524 = ~n29515 & n29523;
  assign n29525 = ~n29512 & n29524;
  assign n29526 = ~n29480 & ~n29486;
  assign n29527 = n29514 & n29526;
  assign n29528 = n29525 & ~n29527;
  assign n29529 = ~n29509 & ~n29528;
  assign n29530 = n29474 & ~n29480;
  assign n29531 = n29494 & n29530;
  assign n29532 = n29468 & n29531;
  assign n29533 = n29486 & n29532;
  assign n29534 = n29487 & ~n29494;
  assign n29535 = n29474 & ~n29494;
  assign n29536 = ~n29486 & n29535;
  assign n29537 = ~n29534 & ~n29536;
  assign n29538 = n29468 & ~n29537;
  assign n29539 = ~n29533 & ~n29538;
  assign n29540 = ~n29509 & ~n29539;
  assign n29541 = ~n29529 & ~n29540;
  assign n29542 = ~n29503 & n29541;
  assign n29543 = ~n29480 & n29486;
  assign n29544 = ~n29468 & n29543;
  assign n29545 = n29535 & n29544;
  assign n29546 = ~n29480 & n29494;
  assign n29547 = n29513 & n29546;
  assign n29548 = n29468 & n29495;
  assign n29549 = n29486 & ~n29494;
  assign n29550 = ~n29480 & n29549;
  assign n29551 = ~n29500 & ~n29550;
  assign n29552 = ~n29548 & n29551;
  assign n29553 = ~n29486 & n29531;
  assign n29554 = n29552 & ~n29553;
  assign n29555 = ~n29468 & n29499;
  assign n29556 = ~n29486 & n29555;
  assign n29557 = ~n29474 & ~n29480;
  assign n29558 = n29486 & n29535;
  assign n29559 = ~n29557 & ~n29558;
  assign n29560 = ~n29468 & ~n29559;
  assign n29561 = ~n29556 & ~n29560;
  assign n29562 = n29554 & n29561;
  assign n29563 = n29509 & ~n29562;
  assign n29564 = ~n29547 & ~n29563;
  assign n29565 = ~n29545 & n29564;
  assign n29566 = n29542 & n29565;
  assign n29567 = pi0484 & n29566;
  assign n29568 = ~pi0484 & ~n29566;
  assign po0532 = n29567 | n29568;
  assign n29570 = ~n29520 & ~n29527;
  assign n29571 = ~n29549 & n29570;
  assign n29572 = ~n29468 & ~n29571;
  assign n29573 = n29468 & n29486;
  assign n29574 = n29494 & n29573;
  assign n29575 = n29480 & n29486;
  assign n29576 = ~n29474 & n29575;
  assign n29577 = ~n29486 & n29517;
  assign n29578 = ~n29576 & ~n29577;
  assign n29579 = ~n29480 & ~n29494;
  assign n29580 = n29468 & ~n29486;
  assign n29581 = n29579 & n29580;
  assign n29582 = n29578 & ~n29581;
  assign n29583 = ~n29574 & n29582;
  assign n29584 = ~n29572 & n29583;
  assign n29585 = n29509 & ~n29584;
  assign n29586 = n29480 & n29499;
  assign n29587 = ~n29486 & n29586;
  assign n29588 = n29486 & n29521;
  assign n29589 = ~n29587 & ~n29588;
  assign n29590 = ~n29468 & ~n29589;
  assign n29591 = ~n29585 & ~n29590;
  assign n29592 = n29486 & n29517;
  assign n29593 = ~n29496 & ~n29531;
  assign n29594 = ~n29468 & ~n29593;
  assign n29595 = ~n29592 & ~n29594;
  assign n29596 = ~n29501 & n29595;
  assign n29597 = ~n29509 & ~n29596;
  assign n29598 = ~n29514 & ~n29535;
  assign n29599 = ~n29480 & ~n29598;
  assign n29600 = ~n29536 & ~n29599;
  assign n29601 = n29468 & ~n29600;
  assign n29602 = ~n29509 & n29601;
  assign n29603 = ~n29597 & ~n29602;
  assign n29604 = n29591 & n29603;
  assign n29605 = pi0486 & ~n29604;
  assign n29606 = ~pi0486 & n29591;
  assign n29607 = n29603 & n29606;
  assign po0533 = n29605 | n29607;
  assign n29609 = ~n28420 & ~n28432;
  assign n29610 = ~n29224 & ~n29609;
  assign n29611 = ~n28406 & ~n29610;
  assign n29612 = n28420 & n28426;
  assign n29613 = n28441 & n29612;
  assign n29614 = ~n29611 & ~n29613;
  assign n29615 = n28406 & n28445;
  assign n29616 = ~n28420 & n29615;
  assign n29617 = ~n28889 & ~n29616;
  assign n29618 = n29614 & n29617;
  assign n29619 = n28412 & ~n29618;
  assign n29620 = ~n28443 & ~n28487;
  assign n29621 = ~n28420 & n28461;
  assign n29622 = n29620 & ~n29621;
  assign n29623 = n28406 & ~n29622;
  assign n29624 = n28445 & n28482;
  assign n29625 = ~n28470 & ~n29624;
  assign n29626 = ~n29623 & n29625;
  assign n29627 = ~n28453 & ~n28463;
  assign n29628 = ~n28406 & ~n29627;
  assign n29629 = n29626 & ~n29628;
  assign n29630 = ~n28412 & ~n29629;
  assign n29631 = ~n29619 & ~n29630;
  assign n29632 = ~n28420 & n28452;
  assign n29633 = n28420 & ~n28458;
  assign n29634 = ~n29632 & ~n29633;
  assign n29635 = ~n28406 & ~n29634;
  assign n29636 = ~n28443 & n29203;
  assign n29637 = n28875 & ~n29636;
  assign n29638 = ~n29635 & ~n29637;
  assign n29639 = n29631 & n29638;
  assign n29640 = ~pi0502 & ~n29639;
  assign n29641 = pi0502 & n29638;
  assign n29642 = ~n29630 & n29641;
  assign n29643 = ~n29619 & n29642;
  assign po0534 = n29640 | n29643;
  assign n29645 = n28656 & n28999;
  assign n29646 = ~n29001 & ~n29645;
  assign n29647 = ~n28678 & ~n29026;
  assign n29648 = n28640 & ~n29647;
  assign n29649 = n28606 & n29648;
  assign n29650 = n29646 & ~n29649;
  assign n29651 = ~n28657 & ~n28665;
  assign n29652 = n28606 & ~n29651;
  assign n29653 = n28633 & ~n28640;
  assign n29654 = ~n28680 & ~n28996;
  assign n29655 = ~n28640 & ~n29654;
  assign n29656 = ~n29653 & ~n29655;
  assign n29657 = n28606 & ~n29656;
  assign n29658 = ~n29652 & ~n29657;
  assign n29659 = n28631 & n28679;
  assign n29660 = n28625 & n29659;
  assign n29661 = n28612 & n28648;
  assign n29662 = ~n28991 & ~n29661;
  assign n29663 = n28640 & ~n29662;
  assign n29664 = ~n28681 & ~n29004;
  assign n29665 = n28612 & n28655;
  assign n29666 = ~n28695 & ~n29665;
  assign n29667 = ~n28640 & ~n29666;
  assign n29668 = n29664 & ~n29667;
  assign n29669 = ~n29663 & n29668;
  assign n29670 = ~n29660 & n29669;
  assign n29671 = ~n28606 & ~n29670;
  assign n29672 = ~n29023 & n29096;
  assign n29673 = n28640 & ~n29672;
  assign n29674 = ~n29671 & ~n29673;
  assign n29675 = n29658 & n29674;
  assign n29676 = n29650 & n29675;
  assign n29677 = ~pi0505 & ~n29676;
  assign n29678 = pi0505 & n29650;
  assign n29679 = n29658 & n29678;
  assign n29680 = n29674 & n29679;
  assign po0535 = n29677 | n29680;
  assign n29682 = ~n28332 & ~n28338;
  assign n29683 = n28305 & ~n29682;
  assign n29684 = ~n28394 & ~n29683;
  assign n29685 = n28311 & n28317;
  assign n29686 = ~n28305 & n29685;
  assign n29687 = n28331 & n29686;
  assign n29688 = n28305 & n28324;
  assign n29689 = n28331 & n29688;
  assign n29690 = ~n29246 & ~n29689;
  assign n29691 = ~n28311 & ~n28331;
  assign n29692 = ~n28317 & n29691;
  assign n29693 = n28331 & n28357;
  assign n29694 = ~n29692 & ~n29693;
  assign n29695 = ~n29685 & n29694;
  assign n29696 = ~n28305 & ~n29695;
  assign n29697 = ~n28341 & ~n29696;
  assign n29698 = n29690 & n29697;
  assign n29699 = n28370 & ~n29698;
  assign n29700 = ~n29687 & ~n29699;
  assign n29701 = ~n28358 & ~n28377;
  assign n29702 = ~n28387 & n29701;
  assign n29703 = n28305 & ~n29702;
  assign n29704 = n28333 & n29691;
  assign n29705 = ~n28361 & ~n29704;
  assign n29706 = ~n28305 & ~n29705;
  assign n29707 = ~n29703 & ~n29706;
  assign n29708 = ~n29256 & n29707;
  assign n29709 = ~n28347 & ~n28388;
  assign n29710 = n29708 & n29709;
  assign n29711 = ~n28370 & ~n29710;
  assign n29712 = n29700 & ~n29711;
  assign n29713 = n29684 & n29712;
  assign n29714 = ~pi0499 & ~n29713;
  assign n29715 = pi0499 & n29700;
  assign n29716 = n29684 & n29715;
  assign n29717 = ~n29711 & n29716;
  assign po0536 = n29714 | n29717;
  assign n29719 = ~n28712 & ~n29149;
  assign n29720 = ~n29137 & n29719;
  assign n29721 = ~n28543 & ~n29720;
  assign n29722 = ~n28723 & ~n28739;
  assign n29723 = ~n28572 & ~n28720;
  assign n29724 = ~n29145 & n29723;
  assign n29725 = n28507 & n29724;
  assign n29726 = ~n28706 & ~n29152;
  assign n29727 = n28543 & ~n29726;
  assign n29728 = n29725 & ~n29727;
  assign n29729 = ~n28513 & n28532;
  assign n29730 = ~n28546 & ~n29729;
  assign n29731 = ~n28554 & n29730;
  assign n29732 = ~n28543 & ~n29731;
  assign n29733 = ~n28526 & n28532;
  assign n29734 = ~n28551 & ~n29733;
  assign n29735 = ~n28513 & ~n29734;
  assign n29736 = ~n28534 & ~n28726;
  assign n29737 = n28543 & ~n29736;
  assign n29738 = ~n29735 & ~n29737;
  assign n29739 = ~n29732 & n29738;
  assign n29740 = ~n28507 & n29739;
  assign n29741 = ~n29728 & ~n29740;
  assign n29742 = n29722 & ~n29741;
  assign n29743 = ~n29721 & n29742;
  assign n29744 = ~pi0522 & ~n29743;
  assign n29745 = pi0522 & n29722;
  assign n29746 = ~n29721 & n29745;
  assign n29747 = ~n29741 & n29746;
  assign po0537 = n29744 | n29747;
  assign n29749 = ~n29287 & n29411;
  assign n29750 = ~n29364 & ~n29749;
  assign n29751 = n29322 & ~n29750;
  assign n29752 = ~n29287 & n29300;
  assign n29753 = ~n29381 & ~n29752;
  assign n29754 = n29322 & ~n29753;
  assign n29755 = ~n29313 & n29331;
  assign n29756 = ~n29301 & ~n29755;
  assign n29757 = ~n29360 & n29756;
  assign n29758 = ~n29322 & ~n29757;
  assign n29759 = ~n29754 & ~n29758;
  assign n29760 = ~n29336 & ~n29349;
  assign n29761 = n29759 & n29760;
  assign n29762 = n29328 & ~n29761;
  assign n29763 = n29313 & n29381;
  assign n29764 = n29305 & ~n29313;
  assign n29765 = ~n29411 & ~n29764;
  assign n29766 = ~n29322 & ~n29765;
  assign n29767 = ~n29763 & ~n29766;
  assign n29768 = n29322 & n29332;
  assign n29769 = n29307 & ~n29768;
  assign n29770 = ~n29360 & n29769;
  assign n29771 = ~n29313 & ~n29770;
  assign n29772 = n29767 & ~n29771;
  assign n29773 = ~n29328 & ~n29772;
  assign n29774 = ~n29762 & ~n29773;
  assign n29775 = n29353 & n29441;
  assign n29776 = n29774 & ~n29775;
  assign n29777 = ~n29751 & n29776;
  assign n29778 = ~pi0495 & ~n29777;
  assign n29779 = pi0495 & ~n29751;
  assign n29780 = n29774 & n29779;
  assign n29781 = ~n29775 & n29780;
  assign po0538 = n29778 | n29781;
  assign n29783 = ~n28923 & n28949;
  assign n29784 = ~n29072 & ~n29783;
  assign n29785 = ~n28916 & n28932;
  assign n29786 = ~n28963 & ~n29785;
  assign n29787 = n28903 & ~n29786;
  assign n29788 = n28923 & n28954;
  assign n29789 = ~n29057 & ~n29788;
  assign n29790 = ~n28903 & ~n29789;
  assign n29791 = ~n29787 & ~n29790;
  assign n29792 = ~n28931 & n29791;
  assign n29793 = n29784 & n29792;
  assign n29794 = ~n29040 & ~n29053;
  assign n29795 = n29793 & n29794;
  assign n29796 = n28941 & ~n29795;
  assign n29797 = n28917 & n29051;
  assign n29798 = n28972 & ~n29797;
  assign n29799 = ~n28903 & ~n29798;
  assign n29800 = ~n28923 & n28960;
  assign n29801 = ~n29799 & ~n29800;
  assign n29802 = n28910 & n28932;
  assign n29803 = n28923 & n28945;
  assign n29804 = ~n29802 & ~n29803;
  assign n29805 = ~n28903 & ~n29804;
  assign n29806 = ~n28903 & n28954;
  assign n29807 = ~n28923 & n29806;
  assign n29808 = ~n29805 & ~n29807;
  assign n29809 = n29801 & n29808;
  assign n29810 = ~n28941 & ~n29809;
  assign n29811 = ~n28949 & ~n28956;
  assign n29812 = ~n29058 & n29811;
  assign n29813 = n28977 & ~n29812;
  assign n29814 = ~n29810 & ~n29813;
  assign n29815 = ~n28931 & ~n29053;
  assign n29816 = n28903 & ~n29815;
  assign n29817 = n29814 & ~n29816;
  assign n29818 = ~n29796 & n29817;
  assign n29819 = ~pi0506 & n29818;
  assign n29820 = pi0506 & ~n29818;
  assign po0539 = n29819 | n29820;
  assign n29822 = n28311 & ~n28317;
  assign n29823 = n28305 & n29822;
  assign n29824 = n28331 & n29823;
  assign n29825 = ~n28331 & n29258;
  assign n29826 = ~n28338 & ~n29825;
  assign n29827 = ~n29263 & n29826;
  assign n29828 = ~n29824 & n29827;
  assign n29829 = ~n28305 & n28334;
  assign n29830 = n29828 & ~n29829;
  assign n29831 = ~n28370 & ~n29830;
  assign n29832 = ~n28388 & ~n29266;
  assign n29833 = ~n28305 & ~n29832;
  assign n29834 = n28370 & n28372;
  assign n29835 = n28305 & n29834;
  assign n29836 = n28317 & n29691;
  assign n29837 = ~n29258 & ~n29836;
  assign n29838 = ~n28340 & n29837;
  assign n29839 = ~n28305 & ~n29838;
  assign n29840 = n28311 & n28357;
  assign n29841 = ~n28331 & n29840;
  assign n29842 = ~n29839 & ~n29841;
  assign n29843 = n28370 & ~n29842;
  assign n29844 = ~n29835 & ~n29843;
  assign n29845 = ~n29833 & n29844;
  assign n29846 = ~n28331 & n28387;
  assign n29847 = ~n28335 & ~n29846;
  assign n29848 = ~n28338 & n29847;
  assign n29849 = ~n29237 & n29848;
  assign n29850 = n28305 & ~n29849;
  assign n29851 = n29845 & ~n29850;
  assign n29852 = ~n29831 & n29851;
  assign n29853 = ~pi0497 & ~n29852;
  assign n29854 = pi0497 & n29845;
  assign n29855 = ~n29831 & n29854;
  assign n29856 = ~n29850 & n29855;
  assign po0540 = n29853 | n29856;
  assign n29858 = ~n29486 & n29500;
  assign n29859 = ~n29577 & ~n29858;
  assign n29860 = n29468 & ~n29859;
  assign n29861 = n29496 & n29573;
  assign n29862 = ~n29860 & ~n29861;
  assign n29863 = ~n29547 & n29862;
  assign n29864 = n29486 & n29531;
  assign n29865 = ~n29521 & ~n29864;
  assign n29866 = ~n29500 & n29865;
  assign n29867 = n29468 & ~n29866;
  assign n29868 = n29509 & n29867;
  assign n29869 = ~n29468 & n29480;
  assign n29870 = ~n29474 & n29869;
  assign n29871 = ~n29494 & n29870;
  assign n29872 = ~n29527 & ~n29545;
  assign n29873 = ~n29519 & n29872;
  assign n29874 = ~n29871 & n29873;
  assign n29875 = n29509 & ~n29874;
  assign n29876 = n29474 & n29869;
  assign n29877 = ~n29494 & n29876;
  assign n29878 = n29486 & n29555;
  assign n29879 = ~n29877 & ~n29878;
  assign n29880 = ~n29576 & n29879;
  assign n29881 = n29474 & n29526;
  assign n29882 = n29486 & n29514;
  assign n29883 = ~n29495 & ~n29882;
  assign n29884 = n29468 & ~n29883;
  assign n29885 = ~n29881 & ~n29884;
  assign n29886 = n29880 & n29885;
  assign n29887 = ~n29509 & ~n29886;
  assign n29888 = ~n29486 & n29877;
  assign n29889 = ~n29887 & ~n29888;
  assign n29890 = ~n29875 & n29889;
  assign n29891 = ~n29868 & n29890;
  assign n29892 = n29863 & n29891;
  assign n29893 = pi0488 & ~n29892;
  assign n29894 = ~pi0488 & n29863;
  assign n29895 = n29891 & n29894;
  assign po0541 = n29893 | n29895;
  assign n29897 = ~n28758 & n28812;
  assign n29898 = ~n29192 & ~n29897;
  assign n29899 = n28752 & n29898;
  assign n29900 = n28758 & n28788;
  assign n29901 = ~n28777 & ~n28780;
  assign n29902 = n28764 & ~n29901;
  assign n29903 = n28770 & n28802;
  assign n29904 = n28758 & n28780;
  assign n29905 = ~n29903 & ~n29904;
  assign n29906 = ~n28752 & n29905;
  assign n29907 = ~n29902 & n29906;
  assign n29908 = ~n29900 & n29907;
  assign n29909 = ~n29899 & ~n29908;
  assign n29910 = n28758 & n29902;
  assign n29911 = ~n29183 & ~n29910;
  assign n29912 = ~n29909 & n29911;
  assign n29913 = n28800 & ~n29912;
  assign n29914 = n28752 & ~n29901;
  assign n29915 = ~n28758 & n29914;
  assign n29916 = n28758 & n28782;
  assign n29917 = ~n28839 & ~n29916;
  assign n29918 = n28752 & ~n29917;
  assign n29919 = ~n28764 & n29914;
  assign n29920 = ~n29918 & ~n29919;
  assign n29921 = ~n29915 & n29920;
  assign n29922 = ~n28800 & ~n29921;
  assign n29923 = ~n29913 & ~n29922;
  assign n29924 = n28752 & n28824;
  assign n29925 = ~n28752 & ~n29911;
  assign n29926 = ~n29924 & ~n29925;
  assign n29927 = ~n28752 & ~n29898;
  assign n29928 = ~n28824 & ~n29927;
  assign n29929 = ~n28800 & ~n29928;
  assign n29930 = n29926 & ~n29929;
  assign n29931 = n29923 & n29930;
  assign n29932 = pi0507 & ~n29931;
  assign n29933 = ~pi0507 & n29930;
  assign n29934 = ~n29922 & n29933;
  assign n29935 = ~n29913 & n29934;
  assign po0542 = n29932 | n29935;
  assign n29937 = n29486 & ~n29598;
  assign n29938 = ~n29480 & n29937;
  assign n29939 = n29474 & n29575;
  assign n29940 = ~n29557 & ~n29939;
  assign n29941 = ~n29521 & n29940;
  assign n29942 = ~n29468 & ~n29941;
  assign n29943 = ~n29530 & ~n29586;
  assign n29944 = n29468 & ~n29943;
  assign n29945 = ~n29942 & ~n29944;
  assign n29946 = ~n29938 & n29945;
  assign n29947 = ~n29486 & n29496;
  assign n29948 = n29946 & ~n29947;
  assign n29949 = ~n29509 & ~n29948;
  assign n29950 = ~n29500 & ~n29531;
  assign n29951 = ~n29496 & ~n29521;
  assign n29952 = n29950 & n29951;
  assign n29953 = n29486 & ~n29952;
  assign n29954 = n29513 & ~n29943;
  assign n29955 = ~n29953 & ~n29954;
  assign n29956 = ~n29577 & n29955;
  assign n29957 = n29509 & ~n29956;
  assign n29958 = ~n29949 & ~n29957;
  assign n29959 = n29486 & n29586;
  assign n29960 = ~n29947 & ~n29959;
  assign n29961 = n29468 & ~n29960;
  assign n29962 = n29958 & ~n29961;
  assign n29963 = pi0483 & ~n29962;
  assign n29964 = ~pi0483 & ~n29961;
  assign n29965 = ~n29957 & n29964;
  assign n29966 = ~n29949 & n29965;
  assign po0543 = n29963 | n29966;
  assign n29968 = n28903 & n28960;
  assign n29969 = ~n28923 & n28945;
  assign n29970 = ~n28944 & ~n29969;
  assign n29971 = n28903 & ~n29970;
  assign n29972 = ~n28903 & ~n29075;
  assign n29973 = ~n29971 & ~n29972;
  assign n29974 = ~n29081 & n29973;
  assign n29975 = n28941 & ~n29974;
  assign n29976 = ~n29968 & ~n29975;
  assign n29977 = n28929 & n29044;
  assign n29978 = ~n29056 & ~n29977;
  assign n29979 = ~n28910 & ~n29978;
  assign n29980 = ~n28931 & ~n29979;
  assign n29981 = ~n29057 & n29980;
  assign n29982 = ~n28903 & n28946;
  assign n29983 = n28923 & n28963;
  assign n29984 = ~n29982 & ~n29983;
  assign n29985 = n29981 & n29984;
  assign n29986 = ~n28941 & ~n29985;
  assign n29987 = ~n29783 & ~n29803;
  assign n29988 = ~n28903 & ~n29987;
  assign n29989 = ~n29986 & ~n29988;
  assign n29990 = n29976 & n29989;
  assign n29991 = ~pi0523 & ~n29990;
  assign n29992 = pi0523 & n29989;
  assign n29993 = ~n29975 & n29992;
  assign n29994 = ~n29968 & n29993;
  assign po0544 = n29991 | n29994;
  assign n29996 = n28752 & n28779;
  assign n29997 = n28802 & ~n29901;
  assign n29998 = ~n28783 & ~n29183;
  assign n29999 = ~n29997 & n29998;
  assign n30000 = ~n28752 & ~n29999;
  assign n30001 = n28758 & n28822;
  assign n30002 = ~n30000 & ~n30001;
  assign n30003 = ~n28764 & n28782;
  assign n30004 = ~n28758 & n28837;
  assign n30005 = ~n30003 & ~n30004;
  assign n30006 = ~n29904 & n30005;
  assign n30007 = n28752 & ~n30006;
  assign n30008 = n30002 & ~n30007;
  assign n30009 = n28800 & ~n30008;
  assign n30010 = ~n29996 & ~n30009;
  assign n30011 = ~n28779 & ~n28784;
  assign n30012 = ~n28758 & n28780;
  assign n30013 = ~n29182 & ~n30012;
  assign n30014 = n28752 & ~n30013;
  assign n30015 = n30011 & ~n30014;
  assign n30016 = ~n28758 & n28822;
  assign n30017 = n28758 & n28843;
  assign n30018 = ~n28837 & ~n30017;
  assign n30019 = ~n30003 & n30018;
  assign n30020 = ~n28752 & ~n30019;
  assign n30021 = ~n30016 & ~n30020;
  assign n30022 = ~n28839 & n30021;
  assign n30023 = n30015 & n30022;
  assign n30024 = ~n28800 & ~n30023;
  assign n30025 = ~n28814 & ~n29900;
  assign n30026 = ~n28752 & ~n30025;
  assign n30027 = ~n30024 & ~n30026;
  assign n30028 = n30010 & n30027;
  assign n30029 = pi0516 & n30028;
  assign n30030 = ~pi0516 & ~n30028;
  assign po0545 = n30029 | n30030;
  assign n30032 = pi3428 & ~pi9040;
  assign n30033 = pi3460 & pi9040;
  assign n30034 = ~n30032 & ~n30033;
  assign n30035 = ~pi0540 & ~n30034;
  assign n30036 = pi0540 & n30034;
  assign n30037 = ~n30035 & ~n30036;
  assign n30038 = pi3440 & pi9040;
  assign n30039 = pi3508 & ~pi9040;
  assign n30040 = ~n30038 & ~n30039;
  assign n30041 = pi0535 & n30040;
  assign n30042 = ~pi0535 & ~n30040;
  assign n30043 = ~n30041 & ~n30042;
  assign n30044 = pi3473 & pi9040;
  assign n30045 = pi3453 & ~pi9040;
  assign n30046 = ~n30044 & ~n30045;
  assign n30047 = ~pi0542 & n30046;
  assign n30048 = pi0542 & ~n30046;
  assign n30049 = ~n30047 & ~n30048;
  assign n30050 = pi3445 & pi9040;
  assign n30051 = pi3474 & ~pi9040;
  assign n30052 = ~n30050 & ~n30051;
  assign n30053 = pi0494 & n30052;
  assign n30054 = ~pi0494 & ~n30052;
  assign n30055 = ~n30053 & ~n30054;
  assign n30056 = n30049 & n30055;
  assign n30057 = pi3459 & pi9040;
  assign n30058 = pi3476 & ~pi9040;
  assign n30059 = ~n30057 & ~n30058;
  assign n30060 = ~pi0519 & n30059;
  assign n30061 = pi0519 & ~n30059;
  assign n30062 = ~n30060 & ~n30061;
  assign n30063 = pi3461 & pi9040;
  assign n30064 = pi3449 & ~pi9040;
  assign n30065 = ~n30063 & ~n30064;
  assign n30066 = ~pi0543 & n30065;
  assign n30067 = pi0543 & ~n30065;
  assign n30068 = ~n30066 & ~n30067;
  assign n30069 = ~n30062 & ~n30068;
  assign n30070 = n30056 & n30069;
  assign n30071 = n30043 & n30070;
  assign n30072 = n30062 & ~n30068;
  assign n30073 = ~n30049 & n30055;
  assign n30074 = n30072 & n30073;
  assign n30075 = n30043 & n30062;
  assign n30076 = ~n30055 & n30075;
  assign n30077 = n30049 & n30076;
  assign n30078 = ~n30049 & ~n30055;
  assign n30079 = n30043 & n30078;
  assign n30080 = ~n30068 & n30079;
  assign n30081 = ~n30062 & n30080;
  assign n30082 = ~n30077 & ~n30081;
  assign n30083 = ~n30074 & n30082;
  assign n30084 = ~n30071 & n30083;
  assign n30085 = n30062 & n30073;
  assign n30086 = ~n30043 & n30085;
  assign n30087 = n30084 & ~n30086;
  assign n30088 = ~n30037 & ~n30087;
  assign n30089 = n30043 & ~n30049;
  assign n30090 = n30055 & n30089;
  assign n30091 = ~n30062 & n30090;
  assign n30092 = ~n30076 & ~n30091;
  assign n30093 = ~n30043 & n30056;
  assign n30094 = ~n30062 & n30093;
  assign n30095 = n30092 & ~n30094;
  assign n30096 = n30068 & ~n30095;
  assign n30097 = ~n30043 & ~n30055;
  assign n30098 = ~n30049 & n30097;
  assign n30099 = n30068 & n30098;
  assign n30100 = ~n30062 & n30099;
  assign n30101 = n30049 & n30075;
  assign n30102 = n30049 & ~n30055;
  assign n30103 = n30062 & n30102;
  assign n30104 = ~n30101 & ~n30103;
  assign n30105 = n30068 & ~n30104;
  assign n30106 = ~n30100 & ~n30105;
  assign n30107 = ~n30037 & ~n30106;
  assign n30108 = ~n30096 & ~n30107;
  assign n30109 = ~n30088 & n30108;
  assign n30110 = ~n30043 & ~n30062;
  assign n30111 = ~n30068 & n30110;
  assign n30112 = n30102 & n30111;
  assign n30113 = ~n30043 & ~n30049;
  assign n30114 = n30072 & n30113;
  assign n30115 = ~n30043 & n30055;
  assign n30116 = ~n30062 & n30102;
  assign n30117 = ~n30115 & ~n30116;
  assign n30118 = ~n30068 & ~n30117;
  assign n30119 = n30056 & ~n30068;
  assign n30120 = n30062 & n30119;
  assign n30121 = ~n30118 & ~n30120;
  assign n30122 = n30068 & n30089;
  assign n30123 = n30049 & ~n30062;
  assign n30124 = ~n30043 & n30123;
  assign n30125 = ~n30093 & ~n30124;
  assign n30126 = ~n30122 & n30125;
  assign n30127 = n30062 & n30098;
  assign n30128 = n30126 & ~n30127;
  assign n30129 = n30121 & n30128;
  assign n30130 = n30037 & ~n30129;
  assign n30131 = ~n30114 & ~n30130;
  assign n30132 = ~n30112 & n30131;
  assign n30133 = n30109 & n30132;
  assign n30134 = pi0553 & n30133;
  assign n30135 = ~pi0553 & ~n30133;
  assign po0570 = n30134 | n30135;
  assign n30137 = n30043 & n30049;
  assign n30138 = ~n30086 & ~n30137;
  assign n30139 = ~n30123 & n30138;
  assign n30140 = ~n30068 & ~n30139;
  assign n30141 = ~n30062 & n30068;
  assign n30142 = ~n30049 & n30141;
  assign n30143 = n30043 & ~n30062;
  assign n30144 = n30055 & n30143;
  assign n30145 = n30062 & n30079;
  assign n30146 = ~n30144 & ~n30145;
  assign n30147 = ~n30043 & n30049;
  assign n30148 = n30062 & n30068;
  assign n30149 = n30147 & n30148;
  assign n30150 = n30146 & ~n30149;
  assign n30151 = ~n30142 & n30150;
  assign n30152 = ~n30140 & n30151;
  assign n30153 = n30037 & ~n30152;
  assign n30154 = n30043 & n30056;
  assign n30155 = n30062 & n30154;
  assign n30156 = n30043 & n30102;
  assign n30157 = ~n30062 & n30156;
  assign n30158 = ~n30155 & ~n30157;
  assign n30159 = ~n30068 & ~n30158;
  assign n30160 = ~n30153 & ~n30159;
  assign n30161 = ~n30062 & n30079;
  assign n30162 = ~n30090 & ~n30098;
  assign n30163 = ~n30068 & ~n30162;
  assign n30164 = ~n30161 & ~n30163;
  assign n30165 = ~n30094 & n30164;
  assign n30166 = ~n30037 & ~n30165;
  assign n30167 = ~n30073 & ~n30102;
  assign n30168 = ~n30043 & ~n30167;
  assign n30169 = ~n30103 & ~n30168;
  assign n30170 = n30068 & ~n30169;
  assign n30171 = ~n30037 & n30170;
  assign n30172 = ~n30166 & ~n30171;
  assign n30173 = n30160 & n30172;
  assign n30174 = pi0555 & ~n30173;
  assign n30175 = ~pi0555 & n30160;
  assign n30176 = n30172 & n30175;
  assign po0572 = n30174 | n30176;
  assign n30178 = pi3474 & pi9040;
  assign n30179 = pi3438 & ~pi9040;
  assign n30180 = ~n30178 & ~n30179;
  assign n30181 = pi0536 & n30180;
  assign n30182 = ~pi0536 & ~n30180;
  assign n30183 = ~n30181 & ~n30182;
  assign n30184 = pi3434 & pi9040;
  assign n30185 = pi3462 & ~pi9040;
  assign n30186 = ~n30184 & ~n30185;
  assign n30187 = pi0540 & n30186;
  assign n30188 = ~pi0540 & ~n30186;
  assign n30189 = ~n30187 & ~n30188;
  assign n30190 = pi3511 & pi9040;
  assign n30191 = pi3459 & ~pi9040;
  assign n30192 = ~n30190 & ~n30191;
  assign n30193 = pi0524 & n30192;
  assign n30194 = ~pi0524 & ~n30192;
  assign n30195 = ~n30193 & ~n30194;
  assign n30196 = n30189 & ~n30195;
  assign n30197 = pi3453 & pi9040;
  assign n30198 = pi3512 & ~pi9040;
  assign n30199 = ~n30197 & ~n30198;
  assign n30200 = ~pi0530 & n30199;
  assign n30201 = pi0530 & ~n30199;
  assign n30202 = ~n30200 & ~n30201;
  assign n30203 = pi3443 & pi9040;
  assign n30204 = pi3460 & ~pi9040;
  assign n30205 = ~n30203 & ~n30204;
  assign n30206 = pi0494 & n30205;
  assign n30207 = ~pi0494 & ~n30205;
  assign n30208 = ~n30206 & ~n30207;
  assign n30209 = ~n30202 & n30208;
  assign n30210 = n30196 & n30209;
  assign n30211 = ~n30202 & ~n30208;
  assign n30212 = ~n30189 & n30211;
  assign n30213 = ~n30210 & ~n30212;
  assign n30214 = ~n30183 & ~n30213;
  assign n30215 = pi3469 & ~pi9040;
  assign n30216 = pi3430 & pi9040;
  assign n30217 = ~n30215 & ~n30216;
  assign n30218 = ~pi0528 & ~n30217;
  assign n30219 = pi0528 & n30217;
  assign n30220 = ~n30218 & ~n30219;
  assign n30221 = n30183 & n30202;
  assign n30222 = n30189 & n30221;
  assign n30223 = n30196 & ~n30208;
  assign n30224 = n30189 & n30195;
  assign n30225 = n30208 & n30224;
  assign n30226 = ~n30223 & ~n30225;
  assign n30227 = ~n30189 & ~n30195;
  assign n30228 = n30208 & n30227;
  assign n30229 = ~n30202 & n30228;
  assign n30230 = n30226 & ~n30229;
  assign n30231 = n30183 & ~n30230;
  assign n30232 = ~n30222 & ~n30231;
  assign n30233 = ~n30189 & n30195;
  assign n30234 = ~n30208 & n30233;
  assign n30235 = ~n30202 & n30234;
  assign n30236 = n30232 & ~n30235;
  assign n30237 = n30202 & n30227;
  assign n30238 = ~n30189 & n30208;
  assign n30239 = n30195 & n30238;
  assign n30240 = ~n30237 & ~n30239;
  assign n30241 = ~n30183 & ~n30240;
  assign n30242 = ~n30208 & n30224;
  assign n30243 = n30202 & n30242;
  assign n30244 = ~n30241 & ~n30243;
  assign n30245 = n30236 & n30244;
  assign n30246 = n30220 & ~n30245;
  assign n30247 = ~n30214 & ~n30246;
  assign n30248 = n30183 & ~n30220;
  assign n30249 = ~n30240 & n30248;
  assign n30250 = ~n30208 & n30227;
  assign n30251 = ~n30242 & ~n30250;
  assign n30252 = ~n30202 & ~n30251;
  assign n30253 = ~n30210 & ~n30252;
  assign n30254 = ~n30220 & ~n30253;
  assign n30255 = ~n30249 & ~n30254;
  assign n30256 = ~n30183 & ~n30220;
  assign n30257 = n30196 & n30202;
  assign n30258 = ~n30234 & ~n30257;
  assign n30259 = n30189 & n30208;
  assign n30260 = n30258 & ~n30259;
  assign n30261 = n30256 & ~n30260;
  assign n30262 = n30255 & ~n30261;
  assign n30263 = n30247 & n30262;
  assign n30264 = ~pi0551 & ~n30263;
  assign n30265 = pi0551 & n30255;
  assign n30266 = n30247 & n30265;
  assign n30267 = ~n30261 & n30266;
  assign po0573 = n30264 | n30267;
  assign n30269 = pi3510 & ~pi9040;
  assign n30270 = pi3447 & pi9040;
  assign n30271 = ~n30269 & ~n30270;
  assign n30272 = ~pi0531 & ~n30271;
  assign n30273 = pi0531 & n30271;
  assign n30274 = ~n30272 & ~n30273;
  assign n30275 = pi3448 & pi9040;
  assign n30276 = pi3431 & ~pi9040;
  assign n30277 = ~n30275 & ~n30276;
  assign n30278 = ~pi0513 & n30277;
  assign n30279 = pi0513 & ~n30277;
  assign n30280 = ~n30278 & ~n30279;
  assign n30281 = pi3479 & pi9040;
  assign n30282 = pi3439 & ~pi9040;
  assign n30283 = ~n30281 & ~n30282;
  assign n30284 = pi0510 & n30283;
  assign n30285 = ~pi0510 & ~n30283;
  assign n30286 = ~n30284 & ~n30285;
  assign n30287 = pi3442 & pi9040;
  assign n30288 = pi3481 & ~pi9040;
  assign n30289 = ~n30287 & ~n30288;
  assign n30290 = ~pi0521 & ~n30289;
  assign n30291 = pi0521 & n30289;
  assign n30292 = ~n30290 & ~n30291;
  assign n30293 = pi3463 & pi9040;
  assign n30294 = pi3468 & ~pi9040;
  assign n30295 = ~n30293 & ~n30294;
  assign n30296 = ~pi0517 & ~n30295;
  assign n30297 = pi0517 & n30295;
  assign n30298 = ~n30296 & ~n30297;
  assign n30299 = n30292 & ~n30298;
  assign n30300 = n30286 & n30299;
  assign n30301 = pi3467 & pi9040;
  assign n30302 = pi3470 & ~pi9040;
  assign n30303 = ~n30301 & ~n30302;
  assign n30304 = ~pi0527 & ~n30303;
  assign n30305 = pi0527 & n30303;
  assign n30306 = ~n30304 & ~n30305;
  assign n30307 = n30298 & n30306;
  assign n30308 = n30292 & n30307;
  assign n30309 = ~n30300 & ~n30308;
  assign n30310 = n30298 & ~n30306;
  assign n30311 = ~n30292 & n30310;
  assign n30312 = ~n30286 & n30311;
  assign n30313 = n30309 & ~n30312;
  assign n30314 = ~n30280 & ~n30313;
  assign n30315 = ~n30292 & n30298;
  assign n30316 = n30306 & n30315;
  assign n30317 = ~n30286 & n30316;
  assign n30318 = ~n30298 & n30306;
  assign n30319 = n30292 & n30318;
  assign n30320 = ~n30286 & n30319;
  assign n30321 = ~n30292 & ~n30298;
  assign n30322 = ~n30310 & ~n30321;
  assign n30323 = n30286 & ~n30322;
  assign n30324 = ~n30320 & ~n30323;
  assign n30325 = ~n30317 & n30324;
  assign n30326 = n30280 & ~n30325;
  assign n30327 = ~n30314 & ~n30326;
  assign n30328 = n30274 & ~n30327;
  assign n30329 = ~n30280 & ~n30286;
  assign n30330 = ~n30298 & n30329;
  assign n30331 = n30280 & n30310;
  assign n30332 = ~n30286 & n30331;
  assign n30333 = ~n30286 & n30292;
  assign n30334 = n30298 & n30333;
  assign n30335 = ~n30300 & ~n30334;
  assign n30336 = n30280 & ~n30335;
  assign n30337 = ~n30332 & ~n30336;
  assign n30338 = n30292 & n30310;
  assign n30339 = ~n30286 & n30338;
  assign n30340 = n30286 & n30316;
  assign n30341 = ~n30339 & ~n30340;
  assign n30342 = ~n30280 & n30286;
  assign n30343 = n30315 & n30342;
  assign n30344 = ~n30292 & n30318;
  assign n30345 = ~n30280 & n30344;
  assign n30346 = ~n30343 & ~n30345;
  assign n30347 = n30341 & n30346;
  assign n30348 = n30337 & n30347;
  assign n30349 = ~n30330 & n30348;
  assign n30350 = ~n30274 & ~n30349;
  assign n30351 = ~n30298 & ~n30306;
  assign n30352 = ~n30292 & n30351;
  assign n30353 = n30280 & ~n30286;
  assign n30354 = n30352 & n30353;
  assign n30355 = n30310 & n30353;
  assign n30356 = n30292 & n30355;
  assign n30357 = ~n30354 & ~n30356;
  assign n30358 = ~n30286 & ~n30292;
  assign n30359 = n30306 & n30358;
  assign n30360 = ~n30298 & n30359;
  assign n30361 = ~n30280 & n30360;
  assign n30362 = n30357 & ~n30361;
  assign n30363 = n30286 & n30307;
  assign n30364 = n30292 & n30351;
  assign n30365 = ~n30286 & n30364;
  assign n30366 = ~n30363 & ~n30365;
  assign n30367 = ~n30280 & ~n30366;
  assign n30368 = n30362 & ~n30367;
  assign n30369 = ~n30350 & n30368;
  assign n30370 = ~n30328 & n30369;
  assign n30371 = ~pi0549 & ~n30370;
  assign n30372 = pi0549 & n30370;
  assign po0576 = n30371 | n30372;
  assign n30374 = pi3471 & pi9040;
  assign n30375 = pi3466 & ~pi9040;
  assign n30376 = ~n30374 & ~n30375;
  assign n30377 = pi0509 & n30376;
  assign n30378 = ~pi0509 & ~n30376;
  assign n30379 = ~n30377 & ~n30378;
  assign n30380 = pi3477 & pi9040;
  assign n30381 = pi3478 & ~pi9040;
  assign n30382 = ~n30380 & ~n30381;
  assign n30383 = pi0518 & n30382;
  assign n30384 = ~pi0518 & ~n30382;
  assign n30385 = ~n30383 & ~n30384;
  assign n30386 = pi3425 & pi9040;
  assign n30387 = pi3447 & ~pi9040;
  assign n30388 = ~n30386 & ~n30387;
  assign n30389 = ~pi0535 & ~n30388;
  assign n30390 = pi0535 & ~n30386;
  assign n30391 = ~n30387 & n30390;
  assign n30392 = ~n30389 & ~n30391;
  assign n30393 = pi3431 & pi9040;
  assign n30394 = pi3450 & ~pi9040;
  assign n30395 = ~n30393 & ~n30394;
  assign n30396 = ~pi0515 & n30395;
  assign n30397 = pi0515 & ~n30395;
  assign n30398 = ~n30396 & ~n30397;
  assign n30399 = n30392 & ~n30398;
  assign n30400 = ~n30385 & n30399;
  assign n30401 = pi3432 & pi9040;
  assign n30402 = pi3479 & ~pi9040;
  assign n30403 = ~n30401 & ~n30402;
  assign n30404 = pi0539 & n30403;
  assign n30405 = ~pi0539 & ~n30403;
  assign n30406 = ~n30404 & ~n30405;
  assign n30407 = n30400 & ~n30406;
  assign n30408 = ~n30392 & n30398;
  assign n30409 = ~n30385 & n30408;
  assign n30410 = ~n30406 & n30409;
  assign n30411 = ~n30407 & ~n30410;
  assign n30412 = n30385 & n30408;
  assign n30413 = n30406 & n30412;
  assign n30414 = n30392 & n30398;
  assign n30415 = ~n30385 & n30414;
  assign n30416 = n30406 & n30415;
  assign n30417 = ~n30413 & ~n30416;
  assign n30418 = n30411 & n30417;
  assign n30419 = n30379 & ~n30418;
  assign n30420 = ~n30385 & n30406;
  assign n30421 = ~n30398 & n30420;
  assign n30422 = ~n30392 & n30421;
  assign n30423 = ~n30415 & ~n30422;
  assign n30424 = n30379 & ~n30423;
  assign n30425 = ~n30398 & ~n30406;
  assign n30426 = ~n30379 & n30425;
  assign n30427 = n30385 & n30392;
  assign n30428 = n30406 & n30408;
  assign n30429 = ~n30427 & ~n30428;
  assign n30430 = ~n30379 & ~n30429;
  assign n30431 = ~n30426 & ~n30430;
  assign n30432 = ~n30392 & ~n30398;
  assign n30433 = n30385 & n30432;
  assign n30434 = ~n30406 & n30433;
  assign n30435 = n30431 & ~n30434;
  assign n30436 = ~n30398 & n30427;
  assign n30437 = n30406 & n30436;
  assign n30438 = n30435 & ~n30437;
  assign n30439 = ~n30424 & n30438;
  assign n30440 = pi3463 & ~pi9040;
  assign n30441 = pi3433 & pi9040;
  assign n30442 = ~n30440 & ~n30441;
  assign n30443 = ~pi0542 & ~n30442;
  assign n30444 = pi0542 & n30442;
  assign n30445 = ~n30443 & ~n30444;
  assign n30446 = ~n30439 & ~n30445;
  assign n30447 = ~n30385 & ~n30398;
  assign n30448 = ~n30379 & n30406;
  assign n30449 = n30445 & n30448;
  assign n30450 = n30447 & n30449;
  assign n30451 = n30398 & ~n30406;
  assign n30452 = ~n30385 & n30451;
  assign n30453 = ~n30379 & ~n30452;
  assign n30454 = n30385 & n30406;
  assign n30455 = ~n30392 & n30454;
  assign n30456 = ~n30399 & ~n30447;
  assign n30457 = ~n30406 & ~n30456;
  assign n30458 = n30379 & ~n30412;
  assign n30459 = ~n30457 & n30458;
  assign n30460 = ~n30455 & n30459;
  assign n30461 = ~n30453 & ~n30460;
  assign n30462 = n30385 & n30414;
  assign n30463 = n30406 & n30462;
  assign n30464 = ~n30461 & ~n30463;
  assign n30465 = n30445 & ~n30464;
  assign n30466 = ~n30450 & ~n30465;
  assign n30467 = ~n30446 & n30466;
  assign n30468 = ~n30419 & n30467;
  assign n30469 = ~n30379 & n30434;
  assign n30470 = n30468 & ~n30469;
  assign n30471 = pi0544 & ~n30470;
  assign n30472 = n30467 & ~n30469;
  assign n30473 = ~pi0544 & n30472;
  assign n30474 = ~n30419 & n30473;
  assign po0578 = n30471 | n30474;
  assign n30476 = ~n30274 & n30280;
  assign n30477 = ~n30286 & n30299;
  assign n30478 = n30286 & n30338;
  assign n30479 = ~n30286 & n30307;
  assign n30480 = ~n30478 & ~n30479;
  assign n30481 = ~n30477 & n30480;
  assign n30482 = n30476 & ~n30481;
  assign n30483 = ~n30306 & n30358;
  assign n30484 = n30286 & n30364;
  assign n30485 = ~n30483 & ~n30484;
  assign n30486 = ~n30308 & ~n30311;
  assign n30487 = n30485 & n30486;
  assign n30488 = ~n30280 & ~n30487;
  assign n30489 = n30286 & n30344;
  assign n30490 = ~n30488 & ~n30489;
  assign n30491 = ~n30274 & ~n30490;
  assign n30492 = ~n30482 & ~n30491;
  assign n30493 = n30292 & n30329;
  assign n30494 = n30306 & n30493;
  assign n30495 = ~n30312 & ~n30494;
  assign n30496 = ~n30307 & ~n30351;
  assign n30497 = n30286 & ~n30496;
  assign n30498 = ~n30352 & ~n30497;
  assign n30499 = n30280 & ~n30498;
  assign n30500 = ~n30319 & ~n30477;
  assign n30501 = ~n30478 & n30500;
  assign n30502 = ~n30280 & ~n30501;
  assign n30503 = ~n30499 & ~n30502;
  assign n30504 = n30286 & n30352;
  assign n30505 = ~n30340 & ~n30504;
  assign n30506 = ~n30360 & n30505;
  assign n30507 = ~n30332 & n30506;
  assign n30508 = n30503 & n30507;
  assign n30509 = n30274 & ~n30508;
  assign n30510 = n30495 & ~n30509;
  assign n30511 = n30492 & n30510;
  assign n30512 = pi0547 & ~n30511;
  assign n30513 = ~pi0547 & n30495;
  assign n30514 = n30492 & n30513;
  assign n30515 = ~n30509 & n30514;
  assign po0580 = n30512 | n30515;
  assign n30517 = ~n30183 & ~n30202;
  assign n30518 = ~n30227 & ~n30242;
  assign n30519 = n30517 & ~n30518;
  assign n30520 = ~n30183 & ~n30208;
  assign n30521 = n30227 & n30520;
  assign n30522 = ~n30519 & ~n30521;
  assign n30523 = n30220 & ~n30522;
  assign n30524 = n30202 & n30208;
  assign n30525 = n30195 & n30524;
  assign n30526 = n30189 & n30525;
  assign n30527 = ~n30259 & ~n30524;
  assign n30528 = n30183 & ~n30527;
  assign n30529 = n30202 & ~n30208;
  assign n30530 = ~n30195 & n30529;
  assign n30531 = n30189 & n30530;
  assign n30532 = ~n30528 & ~n30531;
  assign n30533 = ~n30526 & n30532;
  assign n30534 = n30220 & ~n30533;
  assign n30535 = ~n30523 & ~n30534;
  assign n30536 = n30195 & n30209;
  assign n30537 = ~n30189 & n30536;
  assign n30538 = n30202 & n30234;
  assign n30539 = ~n30537 & ~n30538;
  assign n30540 = ~n30183 & ~n30539;
  assign n30541 = ~n30196 & ~n30259;
  assign n30542 = ~n30202 & ~n30541;
  assign n30543 = ~n30234 & ~n30542;
  assign n30544 = ~n30183 & ~n30543;
  assign n30545 = n30195 & n30202;
  assign n30546 = ~n30183 & n30545;
  assign n30547 = ~n30208 & n30546;
  assign n30548 = ~n30195 & n30208;
  assign n30549 = ~n30234 & ~n30548;
  assign n30550 = n30202 & ~n30549;
  assign n30551 = n30183 & ~n30202;
  assign n30552 = n30224 & n30551;
  assign n30553 = ~n30208 & n30552;
  assign n30554 = ~n30550 & ~n30553;
  assign n30555 = ~n30547 & n30554;
  assign n30556 = ~n30544 & n30555;
  assign n30557 = ~n30537 & n30556;
  assign n30558 = ~n30220 & ~n30557;
  assign n30559 = ~n30202 & n30250;
  assign n30560 = n30202 & n30259;
  assign n30561 = ~n30559 & ~n30560;
  assign n30562 = n30183 & ~n30561;
  assign n30563 = ~n30558 & ~n30562;
  assign n30564 = ~n30540 & n30563;
  assign n30565 = n30535 & n30564;
  assign n30566 = pi0563 & n30565;
  assign n30567 = ~pi0563 & ~n30565;
  assign po0581 = n30566 | n30567;
  assign n30569 = n30062 & n30093;
  assign n30570 = ~n30145 & ~n30569;
  assign n30571 = n30068 & ~n30570;
  assign n30572 = n30090 & n30141;
  assign n30573 = ~n30571 & ~n30572;
  assign n30574 = ~n30114 & n30573;
  assign n30575 = ~n30049 & ~n30062;
  assign n30576 = n30097 & n30575;
  assign n30577 = ~n30156 & ~n30576;
  assign n30578 = ~n30093 & n30577;
  assign n30579 = n30068 & ~n30578;
  assign n30580 = n30037 & n30579;
  assign n30581 = ~n30068 & n30154;
  assign n30582 = ~n30086 & ~n30112;
  assign n30583 = ~n30081 & n30582;
  assign n30584 = ~n30581 & n30583;
  assign n30585 = n30037 & ~n30584;
  assign n30586 = n30043 & ~n30068;
  assign n30587 = ~n30055 & n30586;
  assign n30588 = n30049 & n30587;
  assign n30589 = n30062 & n30588;
  assign n30590 = ~n30062 & n30119;
  assign n30591 = ~n30588 & ~n30590;
  assign n30592 = ~n30144 & n30591;
  assign n30593 = ~n30043 & n30062;
  assign n30594 = ~n30055 & n30593;
  assign n30595 = ~n30062 & n30073;
  assign n30596 = ~n30089 & ~n30595;
  assign n30597 = n30068 & ~n30596;
  assign n30598 = ~n30594 & ~n30597;
  assign n30599 = n30592 & n30598;
  assign n30600 = ~n30037 & ~n30599;
  assign n30601 = ~n30589 & ~n30600;
  assign n30602 = ~n30585 & n30601;
  assign n30603 = ~n30580 & n30602;
  assign n30604 = n30574 & n30603;
  assign n30605 = pi0565 & ~n30604;
  assign n30606 = ~pi0565 & n30574;
  assign n30607 = n30603 & n30606;
  assign po0583 = n30605 | n30607;
  assign n30609 = ~n30062 & ~n30167;
  assign n30610 = ~n30043 & n30609;
  assign n30611 = ~n30055 & n30143;
  assign n30612 = ~n30115 & ~n30611;
  assign n30613 = ~n30156 & n30612;
  assign n30614 = ~n30068 & ~n30613;
  assign n30615 = ~n30097 & ~n30154;
  assign n30616 = n30068 & ~n30615;
  assign n30617 = ~n30614 & ~n30616;
  assign n30618 = ~n30610 & n30617;
  assign n30619 = n30062 & n30090;
  assign n30620 = n30618 & ~n30619;
  assign n30621 = ~n30037 & ~n30620;
  assign n30622 = n30072 & ~n30615;
  assign n30623 = ~n30093 & ~n30098;
  assign n30624 = ~n30090 & ~n30156;
  assign n30625 = n30623 & n30624;
  assign n30626 = ~n30062 & ~n30625;
  assign n30627 = ~n30622 & ~n30626;
  assign n30628 = ~n30145 & n30627;
  assign n30629 = n30037 & ~n30628;
  assign n30630 = ~n30621 & ~n30629;
  assign n30631 = ~n30062 & n30154;
  assign n30632 = ~n30619 & ~n30631;
  assign n30633 = n30068 & ~n30632;
  assign n30634 = n30630 & ~n30633;
  assign n30635 = pi0561 & ~n30634;
  assign n30636 = ~pi0561 & ~n30633;
  assign n30637 = ~n30629 & n30636;
  assign n30638 = ~n30621 & n30637;
  assign po0585 = n30635 | n30638;
  assign n30640 = pi3473 & ~pi9040;
  assign n30641 = pi3436 & pi9040;
  assign n30642 = ~n30640 & ~n30641;
  assign n30643 = ~pi0537 & ~n30642;
  assign n30644 = pi0537 & n30642;
  assign n30645 = ~n30643 & ~n30644;
  assign n30646 = pi3437 & pi9040;
  assign n30647 = pi3443 & ~pi9040;
  assign n30648 = ~n30646 & ~n30647;
  assign n30649 = ~pi0541 & n30648;
  assign n30650 = pi0541 & ~n30648;
  assign n30651 = ~n30649 & ~n30650;
  assign n30652 = pi3438 & pi9040;
  assign n30653 = pi3509 & ~pi9040;
  assign n30654 = ~n30652 & ~n30653;
  assign n30655 = ~pi0532 & ~n30654;
  assign n30656 = pi0532 & ~n30652;
  assign n30657 = ~n30653 & n30656;
  assign n30658 = ~n30655 & ~n30657;
  assign n30659 = pi3512 & pi9040;
  assign n30660 = pi3440 & ~pi9040;
  assign n30661 = ~n30659 & ~n30660;
  assign n30662 = ~pi0520 & ~n30661;
  assign n30663 = pi0520 & n30661;
  assign n30664 = ~n30662 & ~n30663;
  assign n30665 = pi3428 & pi9040;
  assign n30666 = pi3434 & ~pi9040;
  assign n30667 = ~n30665 & ~n30666;
  assign n30668 = ~pi0512 & n30667;
  assign n30669 = pi0512 & ~n30667;
  assign n30670 = ~n30668 & ~n30669;
  assign n30671 = n30664 & n30670;
  assign n30672 = n30658 & n30671;
  assign n30673 = ~n30651 & n30672;
  assign n30674 = ~n30664 & n30670;
  assign n30675 = n30658 & n30674;
  assign n30676 = n30651 & n30675;
  assign n30677 = ~n30673 & ~n30676;
  assign n30678 = ~n30664 & ~n30670;
  assign n30679 = n30658 & n30678;
  assign n30680 = ~n30651 & n30679;
  assign n30681 = pi3444 & pi9040;
  assign n30682 = pi3430 & ~pi9040;
  assign n30683 = ~n30681 & ~n30682;
  assign n30684 = pi0526 & n30683;
  assign n30685 = ~pi0526 & ~n30683;
  assign n30686 = ~n30684 & ~n30685;
  assign n30687 = n30664 & ~n30670;
  assign n30688 = ~n30651 & n30687;
  assign n30689 = ~n30658 & n30678;
  assign n30690 = n30651 & n30689;
  assign n30691 = ~n30688 & ~n30690;
  assign n30692 = ~n30686 & ~n30691;
  assign n30693 = ~n30680 & ~n30692;
  assign n30694 = ~n30658 & n30674;
  assign n30695 = n30686 & n30694;
  assign n30696 = n30678 & n30686;
  assign n30697 = ~n30651 & n30696;
  assign n30698 = ~n30695 & ~n30697;
  assign n30699 = n30693 & n30698;
  assign n30700 = n30677 & n30699;
  assign n30701 = n30645 & ~n30700;
  assign n30702 = ~n30645 & ~n30686;
  assign n30703 = ~n30651 & ~n30658;
  assign n30704 = ~n30664 & n30703;
  assign n30705 = ~n30658 & n30670;
  assign n30706 = ~n30704 & ~n30705;
  assign n30707 = n30702 & ~n30706;
  assign n30708 = n30651 & n30658;
  assign n30709 = ~n30670 & n30708;
  assign n30710 = ~n30664 & n30709;
  assign n30711 = n30651 & n30664;
  assign n30712 = ~n30658 & n30711;
  assign n30713 = ~n30710 & ~n30712;
  assign n30714 = ~n30651 & n30686;
  assign n30715 = n30658 & n30714;
  assign n30716 = ~n30678 & n30715;
  assign n30717 = n30672 & n30686;
  assign n30718 = ~n30716 & ~n30717;
  assign n30719 = n30713 & n30718;
  assign n30720 = ~n30645 & ~n30719;
  assign n30721 = ~n30658 & n30671;
  assign n30722 = n30651 & ~n30686;
  assign n30723 = n30721 & n30722;
  assign n30724 = n30658 & n30687;
  assign n30725 = n30651 & n30724;
  assign n30726 = ~n30676 & ~n30725;
  assign n30727 = ~n30686 & ~n30726;
  assign n30728 = ~n30723 & ~n30727;
  assign n30729 = n30686 & n30710;
  assign n30730 = n30728 & ~n30729;
  assign n30731 = ~n30720 & n30730;
  assign n30732 = ~n30707 & n30731;
  assign n30733 = ~n30701 & n30732;
  assign n30734 = ~n30658 & n30687;
  assign n30735 = n30651 & n30686;
  assign n30736 = n30734 & n30735;
  assign n30737 = n30733 & ~n30736;
  assign n30738 = ~pi0557 & ~n30737;
  assign n30739 = pi0557 & ~n30736;
  assign n30740 = n30732 & n30739;
  assign n30741 = ~n30701 & n30740;
  assign po0586 = n30738 | n30741;
  assign n30743 = pi3450 & pi9040;
  assign n30744 = pi3467 & ~pi9040;
  assign n30745 = ~n30743 & ~n30744;
  assign n30746 = pi0517 & n30745;
  assign n30747 = ~pi0517 & ~n30745;
  assign n30748 = ~n30746 & ~n30747;
  assign n30749 = pi3468 & pi9040;
  assign n30750 = pi3425 & ~pi9040;
  assign n30751 = ~n30749 & ~n30750;
  assign n30752 = pi0538 & n30751;
  assign n30753 = ~pi0538 & ~n30751;
  assign n30754 = ~n30752 & ~n30753;
  assign n30755 = pi3481 & pi9040;
  assign n30756 = pi3477 & ~pi9040;
  assign n30757 = ~n30755 & ~n30756;
  assign n30758 = ~pi0537 & ~n30757;
  assign n30759 = pi0537 & ~n30755;
  assign n30760 = ~n30756 & n30759;
  assign n30761 = ~n30758 & ~n30760;
  assign n30762 = pi3439 & pi9040;
  assign n30763 = pi3427 & ~pi9040;
  assign n30764 = ~n30762 & ~n30763;
  assign n30765 = ~pi0512 & n30764;
  assign n30766 = pi0512 & ~n30764;
  assign n30767 = ~n30765 & ~n30766;
  assign n30768 = pi3429 & pi9040;
  assign n30769 = pi3426 & ~pi9040;
  assign n30770 = ~n30768 & ~n30769;
  assign n30771 = ~pi0521 & ~n30770;
  assign n30772 = pi0521 & ~n30768;
  assign n30773 = ~n30769 & n30772;
  assign n30774 = ~n30771 & ~n30773;
  assign n30775 = ~n30767 & ~n30774;
  assign n30776 = n30761 & n30775;
  assign n30777 = n30754 & n30776;
  assign n30778 = ~n30754 & ~n30767;
  assign n30779 = n30774 & n30778;
  assign n30780 = pi3466 & pi9040;
  assign n30781 = pi3435 & ~pi9040;
  assign n30782 = ~n30780 & ~n30781;
  assign n30783 = ~pi0534 & n30782;
  assign n30784 = pi0534 & ~n30782;
  assign n30785 = ~n30783 & ~n30784;
  assign n30786 = ~n30761 & n30778;
  assign n30787 = n30761 & n30774;
  assign n30788 = n30767 & n30787;
  assign n30789 = ~n30786 & ~n30788;
  assign n30790 = n30785 & ~n30789;
  assign n30791 = ~n30779 & ~n30790;
  assign n30792 = ~n30761 & ~n30774;
  assign n30793 = n30754 & n30792;
  assign n30794 = ~n30767 & n30787;
  assign n30795 = ~n30761 & n30767;
  assign n30796 = ~n30754 & n30767;
  assign n30797 = ~n30774 & n30796;
  assign n30798 = ~n30795 & ~n30797;
  assign n30799 = ~n30794 & n30798;
  assign n30800 = ~n30793 & n30799;
  assign n30801 = ~n30785 & ~n30800;
  assign n30802 = n30791 & ~n30801;
  assign n30803 = ~n30777 & n30802;
  assign n30804 = n30748 & ~n30803;
  assign n30805 = ~n30761 & n30774;
  assign n30806 = n30767 & n30805;
  assign n30807 = ~n30754 & n30806;
  assign n30808 = n30767 & n30792;
  assign n30809 = n30754 & n30808;
  assign n30810 = ~n30777 & ~n30809;
  assign n30811 = ~n30807 & n30810;
  assign n30812 = ~n30785 & ~n30811;
  assign n30813 = ~n30804 & ~n30812;
  assign n30814 = ~n30754 & n30794;
  assign n30815 = n30761 & n30767;
  assign n30816 = n30785 & n30815;
  assign n30817 = n30754 & n30816;
  assign n30818 = ~n30754 & ~n30785;
  assign n30819 = n30775 & n30818;
  assign n30820 = ~n30767 & n30805;
  assign n30821 = n30754 & n30820;
  assign n30822 = ~n30819 & ~n30821;
  assign n30823 = ~n30761 & ~n30767;
  assign n30824 = n30754 & n30823;
  assign n30825 = n30761 & ~n30774;
  assign n30826 = n30767 & n30825;
  assign n30827 = ~n30824 & ~n30826;
  assign n30828 = n30785 & ~n30827;
  assign n30829 = ~n30761 & n30785;
  assign n30830 = n30767 & n30829;
  assign n30831 = ~n30754 & n30830;
  assign n30832 = ~n30828 & ~n30831;
  assign n30833 = n30822 & n30832;
  assign n30834 = ~n30748 & ~n30833;
  assign n30835 = ~n30817 & ~n30834;
  assign n30836 = ~n30814 & n30835;
  assign n30837 = n30813 & n30836;
  assign n30838 = ~pi0556 & ~n30837;
  assign n30839 = ~n30804 & ~n30814;
  assign n30840 = ~n30812 & n30839;
  assign n30841 = n30835 & n30840;
  assign n30842 = pi0556 & n30841;
  assign po0587 = n30838 | n30842;
  assign n30844 = ~n30319 & ~n30352;
  assign n30845 = n30280 & ~n30844;
  assign n30846 = n30286 & n30308;
  assign n30847 = ~n30845 & ~n30846;
  assign n30848 = n30286 & n30298;
  assign n30849 = ~n30315 & ~n30848;
  assign n30850 = ~n30364 & n30849;
  assign n30851 = ~n30280 & ~n30850;
  assign n30852 = n30847 & ~n30851;
  assign n30853 = ~n30274 & ~n30852;
  assign n30854 = n30280 & n30317;
  assign n30855 = ~n30356 & ~n30854;
  assign n30856 = ~n30361 & n30855;
  assign n30857 = ~n30280 & n30298;
  assign n30858 = n30333 & n30857;
  assign n30859 = n30286 & n30319;
  assign n30860 = n30280 & n30315;
  assign n30861 = ~n30859 & ~n30860;
  assign n30862 = ~n30504 & n30861;
  assign n30863 = ~n30858 & n30862;
  assign n30864 = ~n30306 & n30333;
  assign n30865 = ~n30360 & ~n30864;
  assign n30866 = n30863 & n30865;
  assign n30867 = ~n30345 & n30866;
  assign n30868 = n30274 & ~n30867;
  assign n30869 = n30856 & ~n30868;
  assign n30870 = ~n30853 & n30869;
  assign n30871 = ~pi0559 & ~n30870;
  assign n30872 = pi0559 & n30856;
  assign n30873 = ~n30853 & n30872;
  assign n30874 = ~n30868 & n30873;
  assign po0589 = n30871 | n30874;
  assign n30876 = ~n30754 & n30785;
  assign n30877 = n30761 & n30876;
  assign n30878 = ~n30767 & n30792;
  assign n30879 = n30754 & n30878;
  assign n30880 = n30754 & n30806;
  assign n30881 = ~n30879 & ~n30880;
  assign n30882 = ~n30754 & n30808;
  assign n30883 = ~n30788 & ~n30882;
  assign n30884 = ~n30785 & ~n30883;
  assign n30885 = n30881 & ~n30884;
  assign n30886 = ~n30877 & n30885;
  assign n30887 = n30748 & ~n30886;
  assign n30888 = n30754 & n30761;
  assign n30889 = n30767 & n30888;
  assign n30890 = ~n30774 & n30889;
  assign n30891 = n30785 & n30890;
  assign n30892 = n30818 & n30826;
  assign n30893 = ~n30786 & ~n30892;
  assign n30894 = ~n30788 & ~n30820;
  assign n30895 = ~n30754 & n30805;
  assign n30896 = n30894 & ~n30895;
  assign n30897 = n30785 & ~n30896;
  assign n30898 = ~n30785 & n30794;
  assign n30899 = n30810 & ~n30898;
  assign n30900 = ~n30897 & n30899;
  assign n30901 = n30893 & n30900;
  assign n30902 = ~n30748 & ~n30901;
  assign n30903 = ~n30891 & ~n30902;
  assign n30904 = ~n30887 & n30903;
  assign n30905 = n30818 & n30820;
  assign n30906 = n30775 & ~n30785;
  assign n30907 = n30754 & n30906;
  assign n30908 = ~n30905 & ~n30907;
  assign n30909 = ~n30785 & n30880;
  assign n30910 = n30908 & ~n30909;
  assign n30911 = n30904 & n30910;
  assign n30912 = ~pi0545 & ~n30911;
  assign n30913 = pi0545 & n30910;
  assign n30914 = n30903 & n30913;
  assign n30915 = ~n30887 & n30914;
  assign po0590 = n30912 | n30915;
  assign n30917 = pi3476 & pi9040;
  assign n30918 = pi3436 & ~pi9040;
  assign n30919 = ~n30917 & ~n30918;
  assign n30920 = pi0533 & n30919;
  assign n30921 = ~pi0533 & ~n30919;
  assign n30922 = ~n30920 & ~n30921;
  assign n30923 = pi3462 & pi9040;
  assign n30924 = pi3445 & ~pi9040;
  assign n30925 = ~n30923 & ~n30924;
  assign n30926 = pi0525 & n30925;
  assign n30927 = ~pi0525 & ~n30925;
  assign n30928 = ~n30926 & ~n30927;
  assign n30929 = pi3424 & pi9040;
  assign n30930 = pi3444 & ~pi9040;
  assign n30931 = ~n30929 & ~n30930;
  assign n30932 = ~pi0524 & ~n30931;
  assign n30933 = pi0524 & n30931;
  assign n30934 = ~n30932 & ~n30933;
  assign n30935 = pi3446 & pi9040;
  assign n30936 = pi3461 & ~pi9040;
  assign n30937 = ~n30935 & ~n30936;
  assign n30938 = pi0528 & n30937;
  assign n30939 = ~pi0528 & ~n30937;
  assign n30940 = ~n30938 & ~n30939;
  assign n30941 = pi3509 & pi9040;
  assign n30942 = pi3441 & ~pi9040;
  assign n30943 = ~n30941 & ~n30942;
  assign n30944 = ~pi0532 & n30943;
  assign n30945 = pi0532 & ~n30943;
  assign n30946 = ~n30944 & ~n30945;
  assign n30947 = ~n30940 & ~n30946;
  assign n30948 = n30934 & n30947;
  assign n30949 = n30928 & n30948;
  assign n30950 = ~n30922 & n30949;
  assign n30951 = n30940 & n30946;
  assign n30952 = ~n30922 & n30928;
  assign n30953 = n30951 & n30952;
  assign n30954 = ~n30934 & n30953;
  assign n30955 = ~n30950 & ~n30954;
  assign n30956 = ~n30934 & n30947;
  assign n30957 = ~n30928 & n30956;
  assign n30958 = ~n30922 & n30957;
  assign n30959 = ~n30934 & n30951;
  assign n30960 = ~n30922 & n30959;
  assign n30961 = ~n30958 & ~n30960;
  assign n30962 = n30922 & n30940;
  assign n30963 = n30934 & n30962;
  assign n30964 = n30922 & n30947;
  assign n30965 = ~n30963 & ~n30964;
  assign n30966 = n30928 & ~n30965;
  assign n30967 = n30940 & ~n30946;
  assign n30968 = ~n30940 & n30946;
  assign n30969 = ~n30967 & ~n30968;
  assign n30970 = ~n30922 & ~n30934;
  assign n30971 = ~n30928 & ~n30970;
  assign n30972 = ~n30969 & n30971;
  assign n30973 = ~n30934 & ~n30947;
  assign n30974 = n30928 & n30973;
  assign n30975 = ~n30922 & n30974;
  assign n30976 = ~n30972 & ~n30975;
  assign n30977 = ~n30966 & n30976;
  assign n30978 = n30961 & n30977;
  assign n30979 = pi3472 & pi9040;
  assign n30980 = pi3437 & ~pi9040;
  assign n30981 = ~n30979 & ~n30980;
  assign n30982 = ~pi0520 & n30981;
  assign n30983 = pi0520 & ~n30981;
  assign n30984 = ~n30982 & ~n30983;
  assign n30985 = ~n30978 & ~n30984;
  assign n30986 = n30955 & ~n30985;
  assign n30987 = n30934 & n30967;
  assign n30988 = ~n30928 & n30987;
  assign n30989 = n30922 & n30988;
  assign n30990 = ~n30928 & n30984;
  assign n30991 = n30934 & n30951;
  assign n30992 = ~n30969 & n30970;
  assign n30993 = ~n30964 & ~n30992;
  assign n30994 = ~n30991 & n30993;
  assign n30995 = n30990 & ~n30994;
  assign n30996 = n30922 & n30959;
  assign n30997 = ~n30934 & n30962;
  assign n30998 = n30922 & n30968;
  assign n30999 = ~n30997 & ~n30998;
  assign n31000 = ~n30922 & n30947;
  assign n31001 = n30934 & n30968;
  assign n31002 = ~n31000 & ~n31001;
  assign n31003 = n30999 & n31002;
  assign n31004 = n30928 & ~n31003;
  assign n31005 = ~n30996 & ~n31004;
  assign n31006 = n30984 & ~n31005;
  assign n31007 = ~n30995 & ~n31006;
  assign n31008 = ~n30989 & n31007;
  assign n31009 = n30986 & n31008;
  assign n31010 = pi0574 & ~n31009;
  assign n31011 = ~pi0574 & n30986;
  assign n31012 = n31008 & n31011;
  assign po0591 = n31010 | n31012;
  assign n31014 = pi3426 & pi9040;
  assign n31015 = pi3433 & ~pi9040;
  assign n31016 = ~n31014 & ~n31015;
  assign n31017 = ~pi0529 & n31016;
  assign n31018 = pi0529 & ~n31016;
  assign n31019 = ~n31017 & ~n31018;
  assign n31020 = pi3475 & pi9040;
  assign n31021 = pi3442 & ~pi9040;
  assign n31022 = ~n31020 & ~n31021;
  assign n31023 = pi0514 & n31022;
  assign n31024 = ~pi0514 & ~n31022;
  assign n31025 = ~n31023 & ~n31024;
  assign n31026 = pi3470 & pi9040;
  assign n31027 = pi3432 & ~pi9040;
  assign n31028 = ~n31026 & ~n31027;
  assign n31029 = ~pi0527 & ~n31028;
  assign n31030 = pi0527 & ~n31026;
  assign n31031 = ~n31027 & n31030;
  assign n31032 = ~n31029 & ~n31031;
  assign n31033 = pi3465 & pi9040;
  assign n31034 = pi3448 & ~pi9040;
  assign n31035 = ~n31033 & ~n31034;
  assign n31036 = ~pi0531 & n31035;
  assign n31037 = pi0531 & ~n31035;
  assign n31038 = ~n31036 & ~n31037;
  assign n31039 = pi3427 & pi9040;
  assign n31040 = pi3451 & ~pi9040;
  assign n31041 = ~n31039 & ~n31040;
  assign n31042 = ~pi0518 & n31041;
  assign n31043 = pi0518 & ~n31041;
  assign n31044 = ~n31042 & ~n31043;
  assign n31045 = n31038 & ~n31044;
  assign n31046 = ~n31032 & n31045;
  assign n31047 = n31025 & n31046;
  assign n31048 = ~n31038 & n31044;
  assign n31049 = ~n31032 & n31048;
  assign n31050 = n31038 & n31044;
  assign n31051 = n31032 & n31050;
  assign n31052 = n31025 & n31051;
  assign n31053 = ~n31049 & ~n31052;
  assign n31054 = ~n31047 & n31053;
  assign n31055 = ~n31019 & ~n31054;
  assign n31056 = n31032 & n31038;
  assign n31057 = ~n31025 & n31056;
  assign n31058 = n31032 & ~n31038;
  assign n31059 = n31025 & n31058;
  assign n31060 = ~n31057 & ~n31059;
  assign n31061 = n31019 & ~n31060;
  assign n31062 = ~n31055 & ~n31061;
  assign n31063 = pi3510 & pi9040;
  assign n31064 = pi3482 & ~pi9040;
  assign n31065 = ~n31063 & ~n31064;
  assign n31066 = pi0515 & n31065;
  assign n31067 = ~pi0515 & ~n31065;
  assign n31068 = ~n31066 & ~n31067;
  assign n31069 = n31032 & n31045;
  assign n31070 = ~n31032 & ~n31044;
  assign n31071 = ~n31025 & n31070;
  assign n31072 = ~n31038 & n31071;
  assign n31073 = ~n31069 & ~n31072;
  assign n31074 = n31019 & ~n31073;
  assign n31075 = ~n31025 & ~n31032;
  assign n31076 = n31044 & n31075;
  assign n31077 = n31038 & n31076;
  assign n31078 = ~n31047 & ~n31077;
  assign n31079 = n31025 & ~n31032;
  assign n31080 = ~n31038 & n31079;
  assign n31081 = ~n31038 & ~n31044;
  assign n31082 = n31032 & n31081;
  assign n31083 = ~n31025 & n31082;
  assign n31084 = ~n31080 & ~n31083;
  assign n31085 = ~n31019 & ~n31084;
  assign n31086 = n31078 & ~n31085;
  assign n31087 = ~n31074 & n31086;
  assign n31088 = n31068 & ~n31087;
  assign n31089 = n31019 & ~n31025;
  assign n31090 = n31045 & n31089;
  assign n31091 = n31032 & n31048;
  assign n31092 = n31044 & n31079;
  assign n31093 = n31038 & n31092;
  assign n31094 = ~n31091 & ~n31093;
  assign n31095 = n31025 & n31081;
  assign n31096 = n31094 & ~n31095;
  assign n31097 = n31019 & ~n31096;
  assign n31098 = ~n31032 & ~n31038;
  assign n31099 = ~n31019 & ~n31025;
  assign n31100 = n31098 & n31099;
  assign n31101 = ~n31025 & n31049;
  assign n31102 = ~n31100 & ~n31101;
  assign n31103 = ~n31097 & n31102;
  assign n31104 = ~n31090 & n31103;
  assign n31105 = ~n31025 & n31069;
  assign n31106 = n31025 & n31082;
  assign n31107 = ~n31105 & ~n31106;
  assign n31108 = n31104 & n31107;
  assign n31109 = ~n31068 & ~n31108;
  assign n31110 = ~n31032 & n31044;
  assign n31111 = ~n31019 & n31110;
  assign n31112 = ~n31025 & n31111;
  assign n31113 = ~n31109 & ~n31112;
  assign n31114 = ~n31088 & n31113;
  assign n31115 = n31062 & n31114;
  assign n31116 = ~pi0548 & ~n31115;
  assign n31117 = pi0548 & n31115;
  assign po0592 = n31116 | n31117;
  assign n31119 = n30651 & n30694;
  assign n31120 = n30670 & n30703;
  assign n31121 = n30664 & n31120;
  assign n31122 = ~n31119 & ~n31121;
  assign n31123 = n30686 & ~n31122;
  assign n31124 = ~n30710 & ~n30717;
  assign n31125 = ~n30664 & n30708;
  assign n31126 = ~n30712 & ~n31125;
  assign n31127 = ~n30686 & ~n31126;
  assign n31128 = ~n30651 & ~n30686;
  assign n31129 = n30674 & n31128;
  assign n31130 = ~n30658 & n31129;
  assign n31131 = ~n30651 & n30658;
  assign n31132 = ~n30670 & n31131;
  assign n31133 = n30664 & n31132;
  assign n31134 = n30686 & n30689;
  assign n31135 = ~n31133 & ~n31134;
  assign n31136 = ~n31130 & n31135;
  assign n31137 = ~n31127 & n31136;
  assign n31138 = n31124 & n31137;
  assign n31139 = n30645 & ~n31138;
  assign n31140 = ~n30686 & n30710;
  assign n31141 = n30651 & n30717;
  assign n31142 = ~n31140 & ~n31141;
  assign n31143 = ~n31139 & n31142;
  assign n31144 = ~n31123 & n31143;
  assign n31145 = n30658 & ~n30664;
  assign n31146 = n30714 & n31145;
  assign n31147 = ~n30695 & ~n31146;
  assign n31148 = n30686 & n30724;
  assign n31149 = n30651 & n30734;
  assign n31150 = ~n31148 & ~n31149;
  assign n31151 = ~n30651 & n30675;
  assign n31152 = ~n31119 & ~n31151;
  assign n31153 = ~n30651 & n30671;
  assign n31154 = ~n30658 & ~n30670;
  assign n31155 = ~n31153 & ~n31154;
  assign n31156 = ~n30686 & ~n31155;
  assign n31157 = n31152 & ~n31156;
  assign n31158 = n31150 & n31157;
  assign n31159 = n31147 & n31158;
  assign n31160 = ~n30645 & ~n31159;
  assign n31161 = n31144 & ~n31160;
  assign n31162 = ~pi0554 & ~n31161;
  assign n31163 = pi0554 & n31144;
  assign n31164 = ~n31160 & n31163;
  assign po0593 = n31162 | n31164;
  assign n31166 = ~n31141 & ~n31146;
  assign n31167 = n30651 & n30696;
  assign n31168 = n30664 & n30703;
  assign n31169 = ~n30721 & ~n31168;
  assign n31170 = n30686 & ~n31169;
  assign n31171 = ~n31167 & ~n31170;
  assign n31172 = n30687 & n30722;
  assign n31173 = ~n30686 & n30694;
  assign n31174 = ~n31172 & ~n31173;
  assign n31175 = n31171 & n31174;
  assign n31176 = n30664 & n30708;
  assign n31177 = ~n31119 & ~n31176;
  assign n31178 = ~n31151 & n31177;
  assign n31179 = n31175 & n31178;
  assign n31180 = ~n30645 & ~n31179;
  assign n31181 = ~n30710 & ~n30721;
  assign n31182 = ~n31153 & n31181;
  assign n31183 = ~n30686 & ~n31182;
  assign n31184 = ~n30651 & n30689;
  assign n31185 = ~n31133 & ~n31184;
  assign n31186 = ~n30736 & n31185;
  assign n31187 = n30675 & n30686;
  assign n31188 = n31186 & ~n31187;
  assign n31189 = ~n31183 & n31188;
  assign n31190 = n30645 & ~n31189;
  assign n31191 = ~n31119 & n31185;
  assign n31192 = ~n30686 & ~n31191;
  assign n31193 = ~n31190 & ~n31192;
  assign n31194 = ~n31180 & n31193;
  assign n31195 = n31166 & n31194;
  assign n31196 = pi0570 & ~n31195;
  assign n31197 = ~pi0570 & n31195;
  assign po0594 = n31196 | n31197;
  assign n31199 = ~n30754 & n30878;
  assign n31200 = ~n30806 & ~n30814;
  assign n31201 = n30754 & n30775;
  assign n31202 = ~n30754 & n30826;
  assign n31203 = ~n31201 & ~n31202;
  assign n31204 = n31200 & n31203;
  assign n31205 = n30785 & ~n31204;
  assign n31206 = n30754 & n30787;
  assign n31207 = ~n30786 & ~n31206;
  assign n31208 = ~n30808 & n31207;
  assign n31209 = ~n30785 & ~n31208;
  assign n31210 = n30754 & n30767;
  assign n31211 = n30774 & n31210;
  assign n31212 = n30761 & n31211;
  assign n31213 = ~n31209 & ~n31212;
  assign n31214 = ~n31205 & n31213;
  assign n31215 = ~n31199 & n31214;
  assign n31216 = ~n30748 & ~n31215;
  assign n31217 = n30754 & n30785;
  assign n31218 = n30794 & n31217;
  assign n31219 = n30785 & n30808;
  assign n31220 = n30785 & n30820;
  assign n31221 = ~n31219 & ~n31220;
  assign n31222 = ~n30754 & ~n31221;
  assign n31223 = ~n31218 & ~n31222;
  assign n31224 = ~n30754 & n30776;
  assign n31225 = ~n30890 & ~n31224;
  assign n31226 = n30754 & n30805;
  assign n31227 = ~n30754 & n30787;
  assign n31228 = ~n31226 & ~n31227;
  assign n31229 = ~n30776 & n31228;
  assign n31230 = ~n30806 & n31229;
  assign n31231 = ~n30785 & ~n31230;
  assign n31232 = ~n30754 & n30788;
  assign n31233 = ~n31231 & ~n31232;
  assign n31234 = n31225 & n31233;
  assign n31235 = n31223 & n31234;
  assign n31236 = n30748 & ~n31235;
  assign n31237 = n30785 & ~n30881;
  assign n31238 = ~n31236 & ~n31237;
  assign n31239 = ~n30809 & ~n31224;
  assign n31240 = ~n30785 & ~n31239;
  assign n31241 = n31238 & ~n31240;
  assign n31242 = ~n31216 & n31241;
  assign n31243 = pi0550 & ~n31242;
  assign n31244 = ~pi0550 & n31242;
  assign po0595 = n31243 | n31244;
  assign n31246 = ~n30338 & ~n30340;
  assign n31247 = ~n30286 & n30318;
  assign n31248 = n31246 & ~n31247;
  assign n31249 = ~n30280 & ~n31248;
  assign n31250 = n30280 & n30307;
  assign n31251 = ~n30286 & n31250;
  assign n31252 = ~n30312 & ~n31251;
  assign n31253 = ~n31249 & n31252;
  assign n31254 = ~n30364 & ~n30489;
  assign n31255 = n30280 & ~n31254;
  assign n31256 = n31253 & ~n31255;
  assign n31257 = ~n30274 & ~n31256;
  assign n31258 = n30286 & n30292;
  assign n31259 = n30306 & n31258;
  assign n31260 = ~n30280 & n30307;
  assign n31261 = ~n30286 & n31260;
  assign n31262 = ~n30365 & ~n31261;
  assign n31263 = ~n31259 & n31262;
  assign n31264 = ~n30286 & ~n30298;
  assign n31265 = ~n30864 & ~n31264;
  assign n31266 = n30280 & ~n31265;
  assign n31267 = n31263 & ~n31266;
  assign n31268 = n30274 & ~n31267;
  assign n31269 = ~n31257 & ~n31268;
  assign n31270 = ~n30286 & n30351;
  assign n31271 = n30286 & ~n30486;
  assign n31272 = ~n31270 & ~n31271;
  assign n31273 = n30280 & ~n31272;
  assign n31274 = ~n30338 & n30844;
  assign n31275 = n30342 & ~n31274;
  assign n31276 = ~n31273 & ~n31275;
  assign n31277 = n31269 & n31276;
  assign n31278 = ~pi0552 & ~n31277;
  assign n31279 = pi0552 & n31276;
  assign n31280 = ~n31257 & n31279;
  assign n31281 = ~n31268 & n31280;
  assign po0596 = n31278 | n31281;
  assign n31283 = ~n30195 & n30211;
  assign n31284 = ~n30242 & ~n31283;
  assign n31285 = ~n30183 & ~n31284;
  assign n31286 = ~n30202 & n30233;
  assign n31287 = ~n30530 & ~n31286;
  assign n31288 = n30183 & ~n31287;
  assign n31289 = n30202 & n30228;
  assign n31290 = ~n30547 & ~n31289;
  assign n31291 = ~n30210 & n31290;
  assign n31292 = ~n31288 & n31291;
  assign n31293 = ~n31285 & n31292;
  assign n31294 = ~n30526 & ~n30537;
  assign n31295 = n31293 & n31294;
  assign n31296 = n30220 & ~n31295;
  assign n31297 = n30196 & n30524;
  assign n31298 = n30251 & ~n31297;
  assign n31299 = n30183 & ~n31298;
  assign n31300 = n30202 & n30239;
  assign n31301 = ~n31299 & ~n31300;
  assign n31302 = n30189 & n30211;
  assign n31303 = ~n30202 & n30224;
  assign n31304 = ~n31302 & ~n31303;
  assign n31305 = n30183 & ~n31304;
  assign n31306 = n30183 & n30233;
  assign n31307 = n30202 & n31306;
  assign n31308 = ~n31305 & ~n31307;
  assign n31309 = n31301 & n31308;
  assign n31310 = ~n30220 & ~n31309;
  assign n31311 = ~n30228 & ~n30235;
  assign n31312 = ~n30531 & n31311;
  assign n31313 = n30256 & ~n31312;
  assign n31314 = ~n31310 & ~n31313;
  assign n31315 = ~n30210 & ~n30526;
  assign n31316 = ~n30183 & ~n31315;
  assign n31317 = n31314 & ~n31316;
  assign n31318 = ~n31296 & n31317;
  assign n31319 = ~pi0564 & n31318;
  assign n31320 = pi0564 & ~n31318;
  assign po0597 = n31319 | n31320;
  assign n31322 = ~n30934 & n30940;
  assign n31323 = ~n30928 & n31322;
  assign n31324 = n30922 & n31323;
  assign n31325 = ~n30922 & n30968;
  assign n31326 = ~n30956 & ~n31325;
  assign n31327 = ~n30987 & n31326;
  assign n31328 = ~n30928 & ~n31327;
  assign n31329 = ~n30934 & n30967;
  assign n31330 = ~n30948 & ~n31329;
  assign n31331 = n30928 & ~n31330;
  assign n31332 = ~n31328 & ~n31331;
  assign n31333 = n30928 & n30991;
  assign n31334 = ~n30934 & n31325;
  assign n31335 = ~n31333 & ~n31334;
  assign n31336 = n31332 & n31335;
  assign n31337 = n30984 & ~n31336;
  assign n31338 = n30922 & n30948;
  assign n31339 = ~n30922 & n30951;
  assign n31340 = ~n30998 & ~n31339;
  assign n31341 = ~n30928 & ~n31340;
  assign n31342 = ~n31338 & ~n31341;
  assign n31343 = n30928 & n31001;
  assign n31344 = ~n30959 & ~n30987;
  assign n31345 = ~n31343 & n31344;
  assign n31346 = ~n30956 & n31345;
  assign n31347 = ~n30922 & ~n31346;
  assign n31348 = n31342 & ~n31347;
  assign n31349 = ~n30984 & ~n31348;
  assign n31350 = ~n31337 & ~n31349;
  assign n31351 = ~n31324 & n31350;
  assign n31352 = n30922 & n30934;
  assign n31353 = n30946 & n31352;
  assign n31354 = n30940 & n31353;
  assign n31355 = ~n30934 & n30998;
  assign n31356 = ~n31354 & ~n31355;
  assign n31357 = n30928 & ~n31356;
  assign n31358 = n31351 & ~n31357;
  assign n31359 = ~pi0568 & ~n31358;
  assign n31360 = pi0568 & ~n31357;
  assign n31361 = n31350 & n31360;
  assign n31362 = ~n31324 & n31361;
  assign po0598 = n31359 | n31362;
  assign n31364 = ~n30998 & ~n31000;
  assign n31365 = n30928 & ~n31364;
  assign n31366 = ~n30954 & ~n31365;
  assign n31367 = ~n30984 & ~n31366;
  assign n31368 = ~n30967 & ~n31322;
  assign n31369 = ~n30922 & ~n31368;
  assign n31370 = ~n30948 & ~n31369;
  assign n31371 = ~n30928 & ~n31370;
  assign n31372 = ~n30992 & ~n31371;
  assign n31373 = n30922 & n30956;
  assign n31374 = ~n30922 & n30934;
  assign n31375 = n30946 & n31374;
  assign n31376 = n30922 & ~n31368;
  assign n31377 = ~n31375 & ~n31376;
  assign n31378 = n30928 & ~n31377;
  assign n31379 = ~n31373 & ~n31378;
  assign n31380 = n31372 & n31379;
  assign n31381 = n30984 & ~n31380;
  assign n31382 = ~n30967 & n31352;
  assign n31383 = ~n30984 & n31382;
  assign n31384 = n30922 & ~n30934;
  assign n31385 = n30928 & n31384;
  assign n31386 = n30967 & n31385;
  assign n31387 = n30922 & ~n30928;
  assign n31388 = n30934 & n31387;
  assign n31389 = n30946 & n31388;
  assign n31390 = ~n31386 & ~n31389;
  assign n31391 = ~n31383 & n31390;
  assign n31392 = ~n30962 & ~n31001;
  assign n31393 = ~n30928 & ~n30984;
  assign n31394 = ~n31392 & n31393;
  assign n31395 = n31391 & ~n31394;
  assign n31396 = ~n31381 & n31395;
  assign n31397 = ~n31367 & n31396;
  assign n31398 = pi0580 & ~n31397;
  assign n31399 = ~pi0580 & n31397;
  assign po0599 = n31398 | n31399;
  assign n31401 = ~n30882 & ~n31224;
  assign n31402 = ~n31212 & n31401;
  assign n31403 = n30785 & ~n31402;
  assign n31404 = ~n30892 & ~n30909;
  assign n31405 = ~n30890 & ~n31220;
  assign n31406 = ~n30878 & ~n31227;
  assign n31407 = ~n30785 & ~n31406;
  assign n31408 = ~n30814 & ~n31407;
  assign n31409 = n31405 & n31408;
  assign n31410 = n30748 & ~n31409;
  assign n31411 = n30767 & n30774;
  assign n31412 = ~n30795 & ~n31411;
  assign n31413 = n30754 & ~n31412;
  assign n31414 = ~n30776 & ~n30895;
  assign n31415 = ~n30785 & ~n31414;
  assign n31416 = n30754 & n30774;
  assign n31417 = ~n30788 & ~n31416;
  assign n31418 = ~n30792 & n31417;
  assign n31419 = n30785 & ~n31418;
  assign n31420 = ~n31415 & ~n31419;
  assign n31421 = ~n31413 & n31420;
  assign n31422 = ~n30748 & ~n31421;
  assign n31423 = ~n31410 & ~n31422;
  assign n31424 = n31404 & n31423;
  assign n31425 = ~n31403 & n31424;
  assign n31426 = ~pi0569 & ~n31425;
  assign n31427 = pi0569 & n31404;
  assign n31428 = ~n31403 & n31427;
  assign n31429 = n31423 & n31428;
  assign po0600 = n31426 | n31429;
  assign n31431 = ~n30183 & n30239;
  assign n31432 = n30202 & n30224;
  assign n31433 = ~n30223 & ~n31432;
  assign n31434 = ~n30183 & ~n31433;
  assign n31435 = n30183 & ~n30549;
  assign n31436 = ~n31434 & ~n31435;
  assign n31437 = ~n30559 & n31436;
  assign n31438 = n30220 & ~n31437;
  assign n31439 = ~n31431 & ~n31438;
  assign n31440 = n30208 & n30517;
  assign n31441 = ~n30529 & ~n31440;
  assign n31442 = ~n30189 & ~n31441;
  assign n31443 = ~n30210 & ~n31442;
  assign n31444 = ~n30530 & n31443;
  assign n31445 = ~n30202 & n30242;
  assign n31446 = n30183 & n30225;
  assign n31447 = ~n31445 & ~n31446;
  assign n31448 = n31444 & n31447;
  assign n31449 = ~n30220 & ~n31448;
  assign n31450 = ~n31289 & ~n31303;
  assign n31451 = n30183 & ~n31450;
  assign n31452 = ~n31449 & ~n31451;
  assign n31453 = n31439 & n31452;
  assign n31454 = ~pi0589 & ~n31453;
  assign n31455 = pi0589 & n31452;
  assign n31456 = ~n31438 & n31455;
  assign n31457 = ~n31431 & n31456;
  assign po0601 = n31454 | n31457;
  assign n31459 = ~n31038 & n31092;
  assign n31460 = ~n31058 & ~n31077;
  assign n31461 = ~n31019 & ~n31460;
  assign n31462 = ~n31459 & ~n31461;
  assign n31463 = ~n31072 & n31462;
  assign n31464 = n31019 & n31025;
  assign n31465 = n31046 & n31464;
  assign n31466 = ~n31105 & ~n31465;
  assign n31467 = ~n31052 & n31466;
  assign n31468 = n31463 & n31467;
  assign n31469 = n31068 & ~n31468;
  assign n31470 = ~n31032 & n31081;
  assign n31471 = n31025 & n31470;
  assign n31472 = ~n31093 & ~n31471;
  assign n31473 = ~n31025 & n31051;
  assign n31474 = ~n31101 & ~n31473;
  assign n31475 = n31032 & ~n31044;
  assign n31476 = n31025 & ~n31038;
  assign n31477 = ~n31475 & ~n31476;
  assign n31478 = ~n31110 & n31477;
  assign n31479 = n31019 & ~n31478;
  assign n31480 = ~n31019 & n31046;
  assign n31481 = n31025 & n31069;
  assign n31482 = ~n31480 & ~n31481;
  assign n31483 = ~n31479 & n31482;
  assign n31484 = n31474 & n31483;
  assign n31485 = n31472 & n31484;
  assign n31486 = ~n31068 & ~n31485;
  assign n31487 = ~n31469 & ~n31486;
  assign n31488 = pi0546 & ~n31487;
  assign n31489 = ~pi0546 & ~n31469;
  assign n31490 = ~n31486 & n31489;
  assign po0602 = n31488 | n31490;
  assign n31492 = ~n30673 & ~n30704;
  assign n31493 = n30645 & ~n31492;
  assign n31494 = n30679 & ~n30686;
  assign n31495 = ~n30709 & ~n31125;
  assign n31496 = ~n30686 & ~n31495;
  assign n31497 = ~n31494 & ~n31496;
  assign n31498 = n30645 & ~n31497;
  assign n31499 = ~n31493 & ~n31498;
  assign n31500 = n30672 & n31128;
  assign n31501 = ~n31130 & ~n31500;
  assign n31502 = ~n30712 & ~n31154;
  assign n31503 = n30686 & ~n31502;
  assign n31504 = n30645 & n31503;
  assign n31505 = n31501 & ~n31504;
  assign n31506 = n30670 & n30708;
  assign n31507 = n30664 & n31506;
  assign n31508 = n30651 & n30674;
  assign n31509 = ~n31121 & ~n31508;
  assign n31510 = n30686 & ~n31509;
  assign n31511 = ~n30710 & ~n31133;
  assign n31512 = n30651 & n30671;
  assign n31513 = ~n30734 & ~n31512;
  assign n31514 = ~n30686 & ~n31513;
  assign n31515 = n31511 & ~n31514;
  assign n31516 = ~n31510 & n31515;
  assign n31517 = ~n31507 & n31516;
  assign n31518 = ~n30645 & ~n31517;
  assign n31519 = ~n31151 & n31185;
  assign n31520 = n30686 & ~n31519;
  assign n31521 = ~n31518 & ~n31520;
  assign n31522 = n31505 & n31521;
  assign n31523 = n31499 & n31522;
  assign n31524 = ~pi0578 & ~n31523;
  assign n31525 = pi0578 & n31505;
  assign n31526 = n31499 & n31525;
  assign n31527 = n31521 & n31526;
  assign po0603 = n31524 | n31527;
  assign n31529 = ~n30946 & n31374;
  assign n31530 = n31344 & ~n31529;
  assign n31531 = n31393 & ~n31530;
  assign n31532 = ~n30984 & n31001;
  assign n31533 = n30922 & n31532;
  assign n31534 = ~n30934 & ~n30946;
  assign n31535 = ~n30964 & ~n31534;
  assign n31536 = n30928 & ~n31535;
  assign n31537 = ~n31333 & ~n31536;
  assign n31538 = ~n30984 & ~n31537;
  assign n31539 = ~n31533 & ~n31538;
  assign n31540 = ~n30946 & n31384;
  assign n31541 = ~n31334 & ~n31540;
  assign n31542 = n30928 & ~n31541;
  assign n31543 = n31539 & ~n31542;
  assign n31544 = n30947 & n31387;
  assign n31545 = n30934 & n31544;
  assign n31546 = ~n30969 & n31384;
  assign n31547 = ~n31545 & ~n31546;
  assign n31548 = ~n31354 & n31547;
  assign n31549 = ~n30969 & n31374;
  assign n31550 = ~n30960 & ~n31549;
  assign n31551 = n30934 & ~n30940;
  assign n31552 = n30952 & n31551;
  assign n31553 = ~n30958 & ~n31552;
  assign n31554 = n31550 & n31553;
  assign n31555 = n31548 & n31554;
  assign n31556 = n30984 & ~n31555;
  assign n31557 = n31543 & ~n31556;
  assign n31558 = ~n31531 & n31557;
  assign n31559 = ~pi0573 & ~n31558;
  assign n31560 = pi0573 & n31543;
  assign n31561 = ~n31531 & n31560;
  assign n31562 = ~n31556 & n31561;
  assign po0604 = n31559 | n31562;
  assign n31564 = ~n30385 & n30392;
  assign n31565 = ~n30379 & n31564;
  assign n31566 = n30406 & n31565;
  assign n31567 = n30392 & n30421;
  assign n31568 = n30385 & ~n30398;
  assign n31569 = ~n30406 & n31568;
  assign n31570 = ~n30413 & ~n31569;
  assign n31571 = ~n31567 & n31570;
  assign n31572 = ~n31566 & n31571;
  assign n31573 = n30379 & n30409;
  assign n31574 = n31572 & ~n31573;
  assign n31575 = n30445 & ~n31574;
  assign n31576 = ~n30406 & n30415;
  assign n31577 = ~n30463 & ~n31576;
  assign n31578 = n30379 & ~n31577;
  assign n31579 = ~n30445 & n30447;
  assign n31580 = ~n30379 & n31579;
  assign n31581 = n30385 & ~n30406;
  assign n31582 = ~n30392 & n31581;
  assign n31583 = ~n31568 & ~n31582;
  assign n31584 = ~n30415 & n31583;
  assign n31585 = n30379 & ~n31584;
  assign n31586 = ~n30385 & n30432;
  assign n31587 = ~n30406 & n31586;
  assign n31588 = ~n31585 & ~n31587;
  assign n31589 = ~n30445 & ~n31588;
  assign n31590 = ~n31580 & ~n31589;
  assign n31591 = ~n31578 & n31590;
  assign n31592 = ~n30410 & ~n30413;
  assign n31593 = n30406 & n30447;
  assign n31594 = ~n30406 & n30462;
  assign n31595 = ~n31593 & ~n31594;
  assign n31596 = n31592 & n31595;
  assign n31597 = ~n30379 & ~n31596;
  assign n31598 = n31591 & ~n31597;
  assign n31599 = ~n31575 & n31598;
  assign n31600 = ~pi0571 & ~n31599;
  assign n31601 = pi0571 & n31591;
  assign n31602 = ~n31575 & n31601;
  assign n31603 = ~n31597 & n31602;
  assign po0605 = n31600 | n31603;
  assign n31605 = ~n30406 & n30436;
  assign n31606 = ~n30433 & ~n31593;
  assign n31607 = n30379 & ~n31606;
  assign n31608 = ~n31605 & ~n31607;
  assign n31609 = ~n30379 & ~n30406;
  assign n31610 = ~n30398 & n31609;
  assign n31611 = n30392 & n31610;
  assign n31612 = n30414 & n30448;
  assign n31613 = ~n31611 & ~n31612;
  assign n31614 = ~n30379 & n30412;
  assign n31615 = n31613 & ~n31614;
  assign n31616 = ~n30410 & ~n30422;
  assign n31617 = n30398 & n30454;
  assign n31618 = n31616 & ~n31617;
  assign n31619 = n31615 & n31618;
  assign n31620 = n31608 & n31619;
  assign n31621 = ~n30445 & ~n31620;
  assign n31622 = ~n30409 & ~n30433;
  assign n31623 = n30406 & ~n31622;
  assign n31624 = ~n30385 & ~n30406;
  assign n31625 = n30392 & n31624;
  assign n31626 = ~n30462 & ~n31625;
  assign n31627 = n30406 & n31568;
  assign n31628 = n31626 & ~n31627;
  assign n31629 = n30379 & ~n31628;
  assign n31630 = ~n30406 & n30432;
  assign n31631 = ~n31567 & ~n31630;
  assign n31632 = ~n30379 & ~n31631;
  assign n31633 = ~n31576 & ~n31632;
  assign n31634 = ~n31629 & n31633;
  assign n31635 = ~n31623 & n31634;
  assign n31636 = n30445 & ~n31635;
  assign n31637 = n30379 & n30452;
  assign n31638 = ~n31636 & ~n31637;
  assign n31639 = n30427 & n31609;
  assign n31640 = ~n30398 & n31639;
  assign n31641 = n31638 & ~n31640;
  assign n31642 = ~n31621 & n31641;
  assign n31643 = ~pi0562 & ~n31642;
  assign n31644 = pi0562 & n31638;
  assign n31645 = ~n31621 & n31644;
  assign n31646 = ~n31640 & n31645;
  assign po0606 = n31643 | n31646;
  assign n31648 = ~n30407 & ~n30413;
  assign n31649 = ~n30379 & ~n31648;
  assign n31650 = ~n30469 & ~n31649;
  assign n31651 = ~n30385 & ~n30392;
  assign n31652 = n30379 & n31651;
  assign n31653 = n30406 & n31652;
  assign n31654 = ~n30379 & n30399;
  assign n31655 = n30406 & n31654;
  assign n31656 = ~n31614 & ~n31655;
  assign n31657 = n30392 & n31581;
  assign n31658 = n30406 & n30432;
  assign n31659 = ~n31657 & ~n31658;
  assign n31660 = ~n31651 & n31659;
  assign n31661 = n30379 & ~n31660;
  assign n31662 = ~n30416 & ~n31661;
  assign n31663 = n31656 & n31662;
  assign n31664 = ~n30445 & ~n31663;
  assign n31665 = ~n31653 & ~n31664;
  assign n31666 = ~n30433 & ~n30452;
  assign n31667 = ~n30462 & n31666;
  assign n31668 = ~n30379 & ~n31667;
  assign n31669 = ~n30406 & n30412;
  assign n31670 = ~n30436 & ~n31669;
  assign n31671 = n30379 & ~n31670;
  assign n31672 = ~n31625 & ~n31671;
  assign n31673 = ~n31668 & n31672;
  assign n31674 = ~n30422 & ~n30463;
  assign n31675 = n31673 & n31674;
  assign n31676 = n30445 & ~n31675;
  assign n31677 = n31665 & ~n31676;
  assign n31678 = n31650 & n31677;
  assign n31679 = ~pi0566 & ~n31678;
  assign n31680 = pi0566 & n31665;
  assign n31681 = n31650 & n31680;
  assign n31682 = ~n31676 & n31681;
  assign po0607 = n31679 | n31682;
  assign n31684 = ~n31025 & n31081;
  assign n31685 = ~n31473 & ~n31684;
  assign n31686 = ~n31019 & n31685;
  assign n31687 = n31025 & n31056;
  assign n31688 = ~n31045 & ~n31048;
  assign n31689 = n31032 & ~n31688;
  assign n31690 = n31038 & n31075;
  assign n31691 = n31025 & n31048;
  assign n31692 = ~n31690 & ~n31691;
  assign n31693 = ~n31689 & n31692;
  assign n31694 = n31019 & n31693;
  assign n31695 = ~n31687 & n31694;
  assign n31696 = ~n31686 & ~n31695;
  assign n31697 = n31025 & n31689;
  assign n31698 = ~n31471 & ~n31697;
  assign n31699 = ~n31696 & n31698;
  assign n31700 = n31068 & ~n31699;
  assign n31701 = ~n31019 & ~n31688;
  assign n31702 = ~n31025 & n31701;
  assign n31703 = n31025 & n31050;
  assign n31704 = ~n31106 & ~n31703;
  assign n31705 = ~n31019 & ~n31704;
  assign n31706 = ~n31032 & n31701;
  assign n31707 = ~n31705 & ~n31706;
  assign n31708 = ~n31702 & n31707;
  assign n31709 = ~n31068 & ~n31708;
  assign n31710 = ~n31700 & ~n31709;
  assign n31711 = n31019 & ~n31685;
  assign n31712 = ~n31093 & ~n31711;
  assign n31713 = ~n31068 & ~n31712;
  assign n31714 = ~n31019 & n31093;
  assign n31715 = n31019 & ~n31698;
  assign n31716 = ~n31714 & ~n31715;
  assign n31717 = ~n31713 & n31716;
  assign n31718 = n31710 & n31717;
  assign n31719 = pi0560 & ~n31718;
  assign n31720 = ~pi0560 & n31717;
  assign n31721 = ~n31709 & n31720;
  assign n31722 = ~n31700 & n31721;
  assign po0608 = n31719 | n31722;
  assign n31724 = ~n31019 & n31047;
  assign n31725 = n31075 & ~n31688;
  assign n31726 = ~n31051 & ~n31725;
  assign n31727 = ~n31471 & n31726;
  assign n31728 = n31019 & ~n31727;
  assign n31729 = n31025 & n31091;
  assign n31730 = ~n31728 & ~n31729;
  assign n31731 = ~n31032 & n31050;
  assign n31732 = ~n31025 & n31475;
  assign n31733 = ~n31731 & ~n31732;
  assign n31734 = ~n31691 & n31733;
  assign n31735 = ~n31019 & ~n31734;
  assign n31736 = n31730 & ~n31735;
  assign n31737 = n31068 & ~n31736;
  assign n31738 = ~n31724 & ~n31737;
  assign n31739 = ~n31025 & n31048;
  assign n31740 = ~n31470 & ~n31739;
  assign n31741 = ~n31019 & ~n31740;
  assign n31742 = ~n31052 & ~n31741;
  assign n31743 = ~n31047 & ~n31106;
  assign n31744 = n31025 & n31110;
  assign n31745 = ~n31475 & ~n31744;
  assign n31746 = ~n31731 & n31745;
  assign n31747 = n31019 & ~n31746;
  assign n31748 = ~n31025 & n31091;
  assign n31749 = ~n31747 & ~n31748;
  assign n31750 = n31743 & n31749;
  assign n31751 = n31742 & n31750;
  assign n31752 = ~n31068 & ~n31751;
  assign n31753 = ~n31083 & ~n31687;
  assign n31754 = n31019 & ~n31753;
  assign n31755 = ~n31752 & ~n31754;
  assign n31756 = n31738 & n31755;
  assign n31757 = pi0567 & n31756;
  assign n31758 = ~pi0567 & ~n31756;
  assign po0609 = n31757 | n31758;
  assign n31760 = pi3526 & pi9040;
  assign n31761 = pi3532 & ~pi9040;
  assign n31762 = ~n31760 & ~n31761;
  assign n31763 = pi0581 & n31762;
  assign n31764 = ~pi0581 & ~n31762;
  assign n31765 = ~n31763 & ~n31764;
  assign n31766 = pi3536 & pi9040;
  assign n31767 = pi3531 & ~pi9040;
  assign n31768 = ~n31766 & ~n31767;
  assign n31769 = ~pi0572 & ~n31768;
  assign n31770 = pi0572 & ~n31766;
  assign n31771 = ~n31767 & n31770;
  assign n31772 = ~n31769 & ~n31771;
  assign n31773 = pi3501 & pi9040;
  assign n31774 = pi3519 & ~pi9040;
  assign n31775 = ~n31773 & ~n31774;
  assign n31776 = ~pi0604 & ~n31775;
  assign n31777 = pi0604 & ~n31773;
  assign n31778 = ~n31774 & n31777;
  assign n31779 = ~n31776 & ~n31778;
  assign n31780 = pi3521 & pi9040;
  assign n31781 = pi3523 & ~pi9040;
  assign n31782 = ~n31780 & ~n31781;
  assign n31783 = ~pi0584 & n31782;
  assign n31784 = pi0584 & ~n31782;
  assign n31785 = ~n31783 & ~n31784;
  assign n31786 = n31779 & ~n31785;
  assign n31787 = ~n31772 & n31786;
  assign n31788 = pi3529 & pi9040;
  assign n31789 = pi3488 & ~pi9040;
  assign n31790 = ~n31788 & ~n31789;
  assign n31791 = pi0607 & n31790;
  assign n31792 = ~pi0607 & ~n31790;
  assign n31793 = ~n31791 & ~n31792;
  assign n31794 = n31787 & ~n31793;
  assign n31795 = ~n31779 & n31785;
  assign n31796 = ~n31772 & n31795;
  assign n31797 = ~n31793 & n31796;
  assign n31798 = ~n31794 & ~n31797;
  assign n31799 = n31772 & n31795;
  assign n31800 = n31793 & n31799;
  assign n31801 = n31779 & n31785;
  assign n31802 = ~n31772 & n31801;
  assign n31803 = n31793 & n31802;
  assign n31804 = ~n31800 & ~n31803;
  assign n31805 = n31798 & n31804;
  assign n31806 = n31765 & ~n31805;
  assign n31807 = ~n31772 & n31793;
  assign n31808 = ~n31785 & n31807;
  assign n31809 = ~n31779 & n31808;
  assign n31810 = ~n31802 & ~n31809;
  assign n31811 = n31765 & ~n31810;
  assign n31812 = ~n31785 & ~n31793;
  assign n31813 = ~n31765 & n31812;
  assign n31814 = n31772 & n31779;
  assign n31815 = n31793 & n31795;
  assign n31816 = ~n31814 & ~n31815;
  assign n31817 = ~n31765 & ~n31816;
  assign n31818 = ~n31813 & ~n31817;
  assign n31819 = ~n31779 & ~n31785;
  assign n31820 = n31772 & n31819;
  assign n31821 = ~n31793 & n31820;
  assign n31822 = n31818 & ~n31821;
  assign n31823 = ~n31785 & n31814;
  assign n31824 = n31793 & n31823;
  assign n31825 = n31822 & ~n31824;
  assign n31826 = ~n31811 & n31825;
  assign n31827 = ~pi3515 & ~pi9040;
  assign n31828 = ~pi3499 & pi9040;
  assign n31829 = ~n31827 & ~n31828;
  assign n31830 = ~pi0599 & n31829;
  assign n31831 = pi0599 & ~n31829;
  assign n31832 = ~n31830 & ~n31831;
  assign n31833 = ~n31826 & ~n31832;
  assign n31834 = ~n31772 & ~n31785;
  assign n31835 = ~n31765 & n31793;
  assign n31836 = n31832 & n31835;
  assign n31837 = n31834 & n31836;
  assign n31838 = ~n31772 & ~n31793;
  assign n31839 = n31785 & n31838;
  assign n31840 = ~n31765 & ~n31839;
  assign n31841 = n31772 & n31793;
  assign n31842 = ~n31779 & n31841;
  assign n31843 = ~n31786 & ~n31834;
  assign n31844 = ~n31793 & ~n31843;
  assign n31845 = ~n31799 & ~n31844;
  assign n31846 = n31765 & n31845;
  assign n31847 = ~n31842 & n31846;
  assign n31848 = ~n31840 & ~n31847;
  assign n31849 = n31772 & n31801;
  assign n31850 = n31793 & n31849;
  assign n31851 = ~n31848 & ~n31850;
  assign n31852 = n31832 & ~n31851;
  assign n31853 = ~n31837 & ~n31852;
  assign n31854 = ~n31833 & n31853;
  assign n31855 = ~n31806 & n31854;
  assign n31856 = ~n31765 & n31821;
  assign n31857 = n31855 & ~n31856;
  assign n31858 = pi0608 & ~n31857;
  assign n31859 = n31854 & ~n31856;
  assign n31860 = ~pi0608 & n31859;
  assign n31861 = ~n31806 & n31860;
  assign po0624 = n31858 | n31861;
  assign n31863 = pi3498 & pi9040;
  assign n31864 = pi3514 & ~pi9040;
  assign n31865 = ~n31863 & ~n31864;
  assign n31866 = pi0592 & n31865;
  assign n31867 = ~pi0592 & ~n31865;
  assign n31868 = ~n31866 & ~n31867;
  assign n31869 = pi3562 & pi9040;
  assign n31870 = pi3504 & ~pi9040;
  assign n31871 = ~n31869 & ~n31870;
  assign n31872 = ~pi0604 & n31871;
  assign n31873 = pi0604 & ~n31871;
  assign n31874 = ~n31872 & ~n31873;
  assign n31875 = pi3528 & pi9040;
  assign n31876 = pi3492 & ~pi9040;
  assign n31877 = ~n31875 & ~n31876;
  assign n31878 = pi0558 & n31877;
  assign n31879 = ~pi0558 & ~n31877;
  assign n31880 = ~n31878 & ~n31879;
  assign n31881 = pi3494 & pi9040;
  assign n31882 = pi3525 & ~pi9040;
  assign n31883 = ~n31881 & ~n31882;
  assign n31884 = ~pi0599 & ~n31883;
  assign n31885 = pi0599 & n31883;
  assign n31886 = ~n31884 & ~n31885;
  assign n31887 = n31880 & ~n31886;
  assign n31888 = pi3527 & pi9040;
  assign n31889 = pi3491 & ~pi9040;
  assign n31890 = ~n31888 & ~n31889;
  assign n31891 = pi0591 & n31890;
  assign n31892 = ~pi0591 & ~n31890;
  assign n31893 = ~n31891 & ~n31892;
  assign n31894 = pi3495 & pi9040;
  assign n31895 = pi3507 & ~pi9040;
  assign n31896 = ~n31894 & ~n31895;
  assign n31897 = ~pi0595 & n31896;
  assign n31898 = pi0595 & ~n31896;
  assign n31899 = ~n31897 & ~n31898;
  assign n31900 = n31893 & ~n31899;
  assign n31901 = n31887 & n31900;
  assign n31902 = ~n31874 & n31901;
  assign n31903 = ~n31893 & ~n31899;
  assign n31904 = ~pi0599 & n31883;
  assign n31905 = pi0599 & ~n31883;
  assign n31906 = ~n31904 & ~n31905;
  assign n31907 = n31880 & ~n31906;
  assign n31908 = n31903 & n31907;
  assign n31909 = ~n31880 & ~n31906;
  assign n31910 = ~n31874 & n31909;
  assign n31911 = ~n31899 & n31910;
  assign n31912 = n31893 & n31911;
  assign n31913 = ~n31874 & ~n31893;
  assign n31914 = ~n31880 & n31913;
  assign n31915 = ~n31886 & n31914;
  assign n31916 = ~n31912 & ~n31915;
  assign n31917 = ~n31908 & n31916;
  assign n31918 = ~n31902 & n31917;
  assign n31919 = n31874 & ~n31893;
  assign n31920 = n31907 & n31919;
  assign n31921 = n31918 & ~n31920;
  assign n31922 = ~n31868 & ~n31921;
  assign n31923 = ~n31874 & ~n31906;
  assign n31924 = n31880 & n31923;
  assign n31925 = n31893 & n31924;
  assign n31926 = ~n31914 & ~n31925;
  assign n31927 = n31874 & n31887;
  assign n31928 = n31893 & n31927;
  assign n31929 = n31926 & ~n31928;
  assign n31930 = n31899 & ~n31929;
  assign n31931 = n31874 & ~n31880;
  assign n31932 = ~n31906 & n31931;
  assign n31933 = n31899 & n31932;
  assign n31934 = n31893 & n31933;
  assign n31935 = ~n31886 & n31913;
  assign n31936 = ~n31880 & ~n31886;
  assign n31937 = ~n31893 & n31936;
  assign n31938 = ~n31935 & ~n31937;
  assign n31939 = n31899 & ~n31938;
  assign n31940 = ~n31934 & ~n31939;
  assign n31941 = ~n31868 & ~n31940;
  assign n31942 = ~n31930 & ~n31941;
  assign n31943 = ~n31922 & n31942;
  assign n31944 = n31874 & n31893;
  assign n31945 = ~n31899 & n31944;
  assign n31946 = n31936 & n31945;
  assign n31947 = n31874 & ~n31906;
  assign n31948 = n31903 & n31947;
  assign n31949 = n31899 & n31923;
  assign n31950 = n31893 & n31906;
  assign n31951 = n31874 & n31950;
  assign n31952 = ~n31927 & ~n31951;
  assign n31953 = ~n31949 & n31952;
  assign n31954 = ~n31893 & n31932;
  assign n31955 = n31953 & ~n31954;
  assign n31956 = n31887 & ~n31899;
  assign n31957 = ~n31893 & n31956;
  assign n31958 = n31874 & n31880;
  assign n31959 = n31893 & n31936;
  assign n31960 = ~n31958 & ~n31959;
  assign n31961 = ~n31899 & ~n31960;
  assign n31962 = ~n31957 & ~n31961;
  assign n31963 = n31955 & n31962;
  assign n31964 = n31868 & ~n31963;
  assign n31965 = ~n31948 & ~n31964;
  assign n31966 = ~n31946 & n31965;
  assign n31967 = n31943 & n31966;
  assign n31968 = pi0616 & n31967;
  assign n31969 = ~pi0616 & ~n31967;
  assign po0639 = n31968 | n31969;
  assign n31971 = pi3515 & pi9040;
  assign n31972 = pi3520 & ~pi9040;
  assign n31973 = ~n31971 & ~n31972;
  assign n31974 = ~pi0594 & n31973;
  assign n31975 = pi0594 & ~n31973;
  assign n31976 = ~n31974 & ~n31975;
  assign n31977 = pi3518 & pi9040;
  assign n31978 = pi3534 & ~pi9040;
  assign n31979 = ~n31977 & ~n31978;
  assign n31980 = pi0586 & n31979;
  assign n31981 = ~pi0586 & ~n31979;
  assign n31982 = ~n31980 & ~n31981;
  assign n31983 = pi3500 & pi9040;
  assign n31984 = pi3537 & ~pi9040;
  assign n31985 = ~n31983 & ~n31984;
  assign n31986 = ~pi0601 & n31985;
  assign n31987 = pi0601 & ~n31985;
  assign n31988 = ~n31986 & ~n31987;
  assign n31989 = pi3497 & pi9040;
  assign n31990 = pi3517 & ~pi9040;
  assign n31991 = ~n31989 & ~n31990;
  assign n31992 = ~pi0572 & n31991;
  assign n31993 = pi0572 & ~n31991;
  assign n31994 = ~n31992 & ~n31993;
  assign n31995 = n31988 & ~n31994;
  assign n31996 = pi3488 & pi9040;
  assign n31997 = pi3538 & ~pi9040;
  assign n31998 = ~n31996 & ~n31997;
  assign n31999 = ~pi0585 & ~n31998;
  assign n32000 = pi0585 & ~n31996;
  assign n32001 = ~n31997 & n32000;
  assign n32002 = ~n31999 & ~n32001;
  assign n32003 = n31995 & ~n32002;
  assign n32004 = n31982 & n32003;
  assign n32005 = ~n31988 & n31994;
  assign n32006 = ~n32002 & n32005;
  assign n32007 = n31988 & n31994;
  assign n32008 = n32002 & n32007;
  assign n32009 = n31982 & n32008;
  assign n32010 = ~n32006 & ~n32009;
  assign n32011 = ~n32004 & n32010;
  assign n32012 = ~n31976 & ~n32011;
  assign n32013 = n31994 & ~n32002;
  assign n32014 = ~n31976 & n32013;
  assign n32015 = ~n31982 & n32014;
  assign n32016 = n31988 & n32002;
  assign n32017 = ~n31982 & n32016;
  assign n32018 = ~n31988 & n32002;
  assign n32019 = n31982 & n32018;
  assign n32020 = ~n32017 & ~n32019;
  assign n32021 = n31976 & ~n32020;
  assign n32022 = ~n32015 & ~n32021;
  assign n32023 = pi3535 & ~pi9040;
  assign n32024 = ~pi3524 & pi9040;
  assign n32025 = ~n32023 & ~n32024;
  assign n32026 = pi0584 & n32025;
  assign n32027 = ~pi0584 & ~n32025;
  assign n32028 = ~n32026 & ~n32027;
  assign n32029 = n31976 & ~n31982;
  assign n32030 = n31995 & n32029;
  assign n32031 = n32002 & n32005;
  assign n32032 = n31982 & ~n32002;
  assign n32033 = n31994 & n32032;
  assign n32034 = n31988 & n32033;
  assign n32035 = ~n32031 & ~n32034;
  assign n32036 = ~n31988 & ~n31994;
  assign n32037 = n31982 & n32036;
  assign n32038 = n32035 & ~n32037;
  assign n32039 = n31976 & ~n32038;
  assign n32040 = ~n32030 & ~n32039;
  assign n32041 = n32002 & n32036;
  assign n32042 = n31982 & n32041;
  assign n32043 = n31995 & n32002;
  assign n32044 = ~n31982 & n32043;
  assign n32045 = ~n31988 & ~n32002;
  assign n32046 = ~n31976 & ~n31982;
  assign n32047 = n32045 & n32046;
  assign n32048 = ~n31982 & n32006;
  assign n32049 = ~n32047 & ~n32048;
  assign n32050 = ~n32044 & n32049;
  assign n32051 = ~n32042 & n32050;
  assign n32052 = n32040 & n32051;
  assign n32053 = ~n32028 & ~n32052;
  assign n32054 = ~n31994 & ~n32002;
  assign n32055 = ~n31982 & n32054;
  assign n32056 = ~n31988 & n32055;
  assign n32057 = ~n32043 & ~n32056;
  assign n32058 = n31976 & ~n32057;
  assign n32059 = ~n31982 & ~n32002;
  assign n32060 = n31994 & n32059;
  assign n32061 = n31988 & n32060;
  assign n32062 = ~n32004 & ~n32061;
  assign n32063 = ~n31988 & n32032;
  assign n32064 = ~n31982 & n32041;
  assign n32065 = ~n32063 & ~n32064;
  assign n32066 = ~n31976 & ~n32065;
  assign n32067 = n32062 & ~n32066;
  assign n32068 = ~n32058 & n32067;
  assign n32069 = n32028 & ~n32068;
  assign n32070 = ~n32053 & ~n32069;
  assign n32071 = n32022 & n32070;
  assign n32072 = ~n32012 & n32071;
  assign n32073 = ~pi0624 & ~n32072;
  assign n32074 = pi0624 & n32072;
  assign po0640 = n32073 | n32074;
  assign n32076 = ~n31874 & n31906;
  assign n32077 = ~n31920 & ~n32076;
  assign n32078 = ~n31950 & n32077;
  assign n32079 = ~n31899 & ~n32078;
  assign n32080 = n31893 & n31899;
  assign n32081 = n31886 & n32080;
  assign n32082 = ~n31874 & n31893;
  assign n32083 = n31880 & n32082;
  assign n32084 = ~n31893 & n31910;
  assign n32085 = ~n32083 & ~n32084;
  assign n32086 = n31874 & ~n31886;
  assign n32087 = ~n31893 & n31899;
  assign n32088 = n32086 & n32087;
  assign n32089 = n32085 & ~n32088;
  assign n32090 = ~n32081 & n32089;
  assign n32091 = ~n32079 & n32090;
  assign n32092 = n31868 & ~n32091;
  assign n32093 = ~n31874 & n31887;
  assign n32094 = ~n31893 & n32093;
  assign n32095 = ~n31874 & n31936;
  assign n32096 = n31893 & n32095;
  assign n32097 = ~n32094 & ~n32096;
  assign n32098 = ~n31899 & ~n32097;
  assign n32099 = ~n32092 & ~n32098;
  assign n32100 = n31893 & n31910;
  assign n32101 = ~n31924 & ~n31932;
  assign n32102 = ~n31899 & ~n32101;
  assign n32103 = ~n32100 & ~n32102;
  assign n32104 = ~n31928 & n32103;
  assign n32105 = ~n31868 & ~n32104;
  assign n32106 = ~n31907 & ~n31936;
  assign n32107 = n31874 & ~n32106;
  assign n32108 = ~n31937 & ~n32107;
  assign n32109 = n31899 & ~n32108;
  assign n32110 = ~n31868 & n32109;
  assign n32111 = ~n32105 & ~n32110;
  assign n32112 = n32099 & n32111;
  assign n32113 = pi0617 & ~n32112;
  assign n32114 = ~pi0617 & n32099;
  assign n32115 = n32111 & n32114;
  assign po0642 = n32113 | n32115;
  assign n32117 = ~n31893 & n31927;
  assign n32118 = ~n32084 & ~n32117;
  assign n32119 = n31899 & ~n32118;
  assign n32120 = n31924 & n32080;
  assign n32121 = ~n32119 & ~n32120;
  assign n32122 = ~n31948 & n32121;
  assign n32123 = n31893 & ~n31906;
  assign n32124 = n31931 & n32123;
  assign n32125 = ~n32095 & ~n32124;
  assign n32126 = ~n31927 & n32125;
  assign n32127 = n31899 & ~n32126;
  assign n32128 = n31868 & n32127;
  assign n32129 = ~n31899 & n32093;
  assign n32130 = ~n31920 & ~n31946;
  assign n32131 = ~n31912 & n32130;
  assign n32132 = ~n32129 & n32131;
  assign n32133 = n31868 & ~n32132;
  assign n32134 = ~n31874 & ~n31899;
  assign n32135 = ~n31880 & n32134;
  assign n32136 = ~n31886 & n32135;
  assign n32137 = ~n31893 & n32136;
  assign n32138 = n31893 & n31956;
  assign n32139 = ~n32136 & ~n32138;
  assign n32140 = ~n32083 & n32139;
  assign n32141 = ~n31880 & n31919;
  assign n32142 = n31893 & n31907;
  assign n32143 = ~n31923 & ~n32142;
  assign n32144 = n31899 & ~n32143;
  assign n32145 = ~n32141 & ~n32144;
  assign n32146 = n32140 & n32145;
  assign n32147 = ~n31868 & ~n32146;
  assign n32148 = ~n32137 & ~n32147;
  assign n32149 = ~n32133 & n32148;
  assign n32150 = ~n32128 & n32149;
  assign n32151 = n32122 & n32150;
  assign n32152 = pi0629 & ~n32151;
  assign n32153 = ~pi0629 & n32122;
  assign n32154 = n32150 & n32153;
  assign po0643 = n32152 | n32154;
  assign n32156 = pi3513 & ~pi9040;
  assign n32157 = pi3525 & pi9040;
  assign n32158 = ~n32156 & ~n32157;
  assign n32159 = ~pi0606 & ~n32158;
  assign n32160 = pi0606 & n32158;
  assign n32161 = ~n32159 & ~n32160;
  assign n32162 = pi3483 & pi9040;
  assign n32163 = pi3503 & ~pi9040;
  assign n32164 = ~n32162 & ~n32163;
  assign n32165 = ~pi0579 & ~n32164;
  assign n32166 = pi0579 & n32164;
  assign n32167 = ~n32165 & ~n32166;
  assign n32168 = pi3559 & pi9040;
  assign n32169 = pi3487 & ~pi9040;
  assign n32170 = ~n32168 & ~n32169;
  assign n32171 = ~pi0605 & n32170;
  assign n32172 = pi0605 & ~n32170;
  assign n32173 = ~n32171 & ~n32172;
  assign n32174 = pi3504 & pi9040;
  assign n32175 = pi3567 & ~pi9040;
  assign n32176 = ~n32174 & ~n32175;
  assign n32177 = pi0582 & n32176;
  assign n32178 = ~pi0582 & ~n32176;
  assign n32179 = ~n32177 & ~n32178;
  assign n32180 = pi3489 & pi9040;
  assign n32181 = pi3498 & ~pi9040;
  assign n32182 = ~n32180 & ~n32181;
  assign n32183 = ~pi0583 & ~n32182;
  assign n32184 = pi0583 & n32182;
  assign n32185 = ~n32183 & ~n32184;
  assign n32186 = ~n32179 & n32185;
  assign n32187 = ~n32173 & n32186;
  assign n32188 = n32167 & n32187;
  assign n32189 = pi3485 & pi9040;
  assign n32190 = pi3493 & ~pi9040;
  assign n32191 = ~n32189 & ~n32190;
  assign n32192 = pi0598 & n32191;
  assign n32193 = ~pi0598 & ~n32191;
  assign n32194 = ~n32192 & ~n32193;
  assign n32195 = n32179 & n32185;
  assign n32196 = n32167 & n32195;
  assign n32197 = n32173 & n32186;
  assign n32198 = ~n32167 & n32197;
  assign n32199 = ~n32196 & ~n32198;
  assign n32200 = ~n32194 & ~n32199;
  assign n32201 = ~n32188 & ~n32200;
  assign n32202 = ~n32179 & ~n32185;
  assign n32203 = n32173 & n32202;
  assign n32204 = n32194 & n32203;
  assign n32205 = n32186 & n32194;
  assign n32206 = n32167 & n32205;
  assign n32207 = ~n32204 & ~n32206;
  assign n32208 = n32201 & n32207;
  assign n32209 = n32179 & ~n32185;
  assign n32210 = ~n32173 & n32209;
  assign n32211 = n32167 & n32210;
  assign n32212 = ~n32173 & n32202;
  assign n32213 = ~n32167 & n32212;
  assign n32214 = ~n32211 & ~n32213;
  assign n32215 = n32208 & n32214;
  assign n32216 = n32161 & ~n32215;
  assign n32217 = ~n32161 & ~n32194;
  assign n32218 = n32167 & n32173;
  assign n32219 = ~n32179 & n32218;
  assign n32220 = n32173 & ~n32185;
  assign n32221 = ~n32219 & ~n32220;
  assign n32222 = n32217 & ~n32221;
  assign n32223 = ~n32167 & ~n32173;
  assign n32224 = n32185 & n32223;
  assign n32225 = ~n32179 & n32224;
  assign n32226 = ~n32167 & n32179;
  assign n32227 = n32173 & n32226;
  assign n32228 = ~n32225 & ~n32227;
  assign n32229 = n32167 & n32194;
  assign n32230 = ~n32173 & n32229;
  assign n32231 = ~n32186 & n32230;
  assign n32232 = n32194 & n32210;
  assign n32233 = ~n32231 & ~n32232;
  assign n32234 = n32228 & n32233;
  assign n32235 = ~n32161 & ~n32234;
  assign n32236 = n32173 & n32209;
  assign n32237 = ~n32167 & ~n32194;
  assign n32238 = n32236 & n32237;
  assign n32239 = ~n32173 & n32195;
  assign n32240 = ~n32167 & n32239;
  assign n32241 = ~n32213 & ~n32240;
  assign n32242 = ~n32194 & ~n32241;
  assign n32243 = ~n32238 & ~n32242;
  assign n32244 = n32194 & n32225;
  assign n32245 = n32243 & ~n32244;
  assign n32246 = ~n32235 & n32245;
  assign n32247 = ~n32222 & n32246;
  assign n32248 = ~n32216 & n32247;
  assign n32249 = n32173 & n32195;
  assign n32250 = ~n32167 & n32194;
  assign n32251 = n32249 & n32250;
  assign n32252 = n32248 & ~n32251;
  assign n32253 = ~pi0621 & ~n32252;
  assign n32254 = n32247 & ~n32251;
  assign n32255 = pi0621 & n32254;
  assign n32256 = ~n32216 & n32255;
  assign po0644 = n32253 | n32256;
  assign n32258 = pi3567 & pi9040;
  assign n32259 = pi3494 & ~pi9040;
  assign n32260 = ~n32258 & ~n32259;
  assign n32261 = ~pi0600 & ~n32260;
  assign n32262 = pi0600 & ~n32258;
  assign n32263 = ~n32259 & n32262;
  assign n32264 = ~n32261 & ~n32263;
  assign n32265 = pi3506 & pi9040;
  assign n32266 = pi3489 & ~pi9040;
  assign n32267 = ~n32265 & ~n32266;
  assign n32268 = pi0592 & n32267;
  assign n32269 = ~pi0592 & ~n32267;
  assign n32270 = ~n32268 & ~n32269;
  assign n32271 = pi3491 & pi9040;
  assign n32272 = pi3580 & ~pi9040;
  assign n32273 = ~n32271 & ~n32272;
  assign n32274 = pi0602 & n32273;
  assign n32275 = ~pi0602 & ~n32273;
  assign n32276 = ~n32274 & ~n32275;
  assign n32277 = ~n32270 & ~n32276;
  assign n32278 = ~n32264 & n32277;
  assign n32279 = pi3514 & pi9040;
  assign n32280 = pi3483 & ~pi9040;
  assign n32281 = ~n32279 & ~n32280;
  assign n32282 = ~pi0558 & n32281;
  assign n32283 = pi0558 & ~n32281;
  assign n32284 = ~n32282 & ~n32283;
  assign n32285 = ~n32270 & ~n32284;
  assign n32286 = n32276 & n32285;
  assign n32287 = ~n32278 & ~n32286;
  assign n32288 = pi3487 & pi9040;
  assign n32289 = pi3528 & ~pi9040;
  assign n32290 = ~n32288 & ~n32289;
  assign n32291 = ~pi0588 & n32290;
  assign n32292 = pi0588 & ~n32290;
  assign n32293 = ~n32291 & ~n32292;
  assign n32294 = pi3486 & pi9040;
  assign n32295 = pi3485 & ~pi9040;
  assign n32296 = ~n32294 & ~n32295;
  assign n32297 = ~pi0575 & ~n32296;
  assign n32298 = pi0575 & n32296;
  assign n32299 = ~n32297 & ~n32298;
  assign n32300 = ~n32293 & ~n32299;
  assign n32301 = ~n32287 & n32300;
  assign n32302 = n32270 & ~n32276;
  assign n32303 = n32264 & ~n32284;
  assign n32304 = n32302 & n32303;
  assign n32305 = n32270 & n32276;
  assign n32306 = n32284 & n32305;
  assign n32307 = n32277 & n32284;
  assign n32308 = ~n32306 & ~n32307;
  assign n32309 = n32264 & ~n32308;
  assign n32310 = ~n32304 & ~n32309;
  assign n32311 = ~n32299 & ~n32310;
  assign n32312 = ~n32301 & ~n32311;
  assign n32313 = n32264 & n32284;
  assign n32314 = ~n32270 & n32313;
  assign n32315 = ~n32304 & ~n32314;
  assign n32316 = n32293 & ~n32315;
  assign n32317 = ~n32264 & ~n32293;
  assign n32318 = n32270 & n32317;
  assign n32319 = n32284 & n32302;
  assign n32320 = ~n32284 & n32305;
  assign n32321 = ~n32319 & ~n32320;
  assign n32322 = n32277 & ~n32284;
  assign n32323 = n32264 & n32322;
  assign n32324 = n32321 & ~n32323;
  assign n32325 = ~n32293 & ~n32324;
  assign n32326 = ~n32318 & ~n32325;
  assign n32327 = ~n32270 & n32276;
  assign n32328 = n32284 & n32327;
  assign n32329 = n32264 & n32328;
  assign n32330 = n32326 & ~n32329;
  assign n32331 = ~n32287 & n32293;
  assign n32332 = ~n32264 & n32306;
  assign n32333 = ~n32331 & ~n32332;
  assign n32334 = n32330 & n32333;
  assign n32335 = n32299 & ~n32334;
  assign n32336 = ~n32316 & ~n32335;
  assign n32337 = n32293 & ~n32299;
  assign n32338 = ~n32264 & n32302;
  assign n32339 = ~n32328 & ~n32338;
  assign n32340 = n32270 & ~n32284;
  assign n32341 = n32339 & ~n32340;
  assign n32342 = n32337 & ~n32341;
  assign n32343 = n32336 & ~n32342;
  assign n32344 = n32312 & n32343;
  assign n32345 = ~pi0610 & ~n32344;
  assign n32346 = pi0610 & n32312;
  assign n32347 = n32336 & n32346;
  assign n32348 = ~n32342 & n32347;
  assign po0645 = n32345 | n32348;
  assign n32350 = ~n32167 & n32220;
  assign n32351 = ~n32179 & n32350;
  assign n32352 = ~n32185 & n32218;
  assign n32353 = n32179 & n32352;
  assign n32354 = ~n32351 & ~n32353;
  assign n32355 = n32194 & ~n32354;
  assign n32356 = ~n32225 & ~n32232;
  assign n32357 = n32167 & ~n32173;
  assign n32358 = n32185 & n32357;
  assign n32359 = n32179 & n32358;
  assign n32360 = n32167 & ~n32194;
  assign n32361 = n32202 & n32360;
  assign n32362 = n32173 & n32361;
  assign n32363 = ~n32179 & n32223;
  assign n32364 = ~n32227 & ~n32363;
  assign n32365 = ~n32194 & ~n32364;
  assign n32366 = n32173 & n32194;
  assign n32367 = n32185 & n32366;
  assign n32368 = ~n32179 & n32367;
  assign n32369 = ~n32365 & ~n32368;
  assign n32370 = ~n32362 & n32369;
  assign n32371 = ~n32359 & n32370;
  assign n32372 = n32356 & n32371;
  assign n32373 = n32161 & ~n32372;
  assign n32374 = ~n32194 & n32225;
  assign n32375 = ~n32167 & n32232;
  assign n32376 = ~n32374 & ~n32375;
  assign n32377 = ~n32373 & n32376;
  assign n32378 = ~n32355 & n32377;
  assign n32379 = ~n32173 & ~n32179;
  assign n32380 = n32229 & n32379;
  assign n32381 = ~n32204 & ~n32380;
  assign n32382 = n32194 & n32239;
  assign n32383 = ~n32167 & n32249;
  assign n32384 = ~n32382 & ~n32383;
  assign n32385 = n32167 & n32212;
  assign n32386 = ~n32351 & ~n32385;
  assign n32387 = n32167 & n32209;
  assign n32388 = n32173 & n32185;
  assign n32389 = ~n32387 & ~n32388;
  assign n32390 = ~n32194 & ~n32389;
  assign n32391 = n32386 & ~n32390;
  assign n32392 = n32384 & n32391;
  assign n32393 = n32381 & n32392;
  assign n32394 = ~n32161 & ~n32393;
  assign n32395 = n32378 & ~n32394;
  assign n32396 = ~pi0618 & ~n32395;
  assign n32397 = pi0618 & n32378;
  assign n32398 = ~n32394 & n32397;
  assign po0647 = n32396 | n32398;
  assign n32400 = pi3523 & pi9040;
  assign n32401 = pi3500 & ~pi9040;
  assign n32402 = ~n32400 & ~n32401;
  assign n32403 = ~pi0593 & n32402;
  assign n32404 = pi0593 & ~n32402;
  assign n32405 = ~n32403 & ~n32404;
  assign n32406 = pi3501 & ~pi9040;
  assign n32407 = pi3535 & pi9040;
  assign n32408 = ~n32406 & ~n32407;
  assign n32409 = ~pi0601 & ~n32408;
  assign n32410 = pi0601 & n32408;
  assign n32411 = ~n32409 & ~n32410;
  assign n32412 = n32405 & ~n32411;
  assign n32413 = pi3484 & pi9040;
  assign n32414 = pi3529 & ~pi9040;
  assign n32415 = ~n32413 & ~n32414;
  assign n32416 = pi0576 & n32415;
  assign n32417 = ~pi0576 & ~n32415;
  assign n32418 = ~n32416 & ~n32417;
  assign n32419 = pi3539 & pi9040;
  assign n32420 = pi3518 & ~pi9040;
  assign n32421 = ~n32419 & ~n32420;
  assign n32422 = ~pi0590 & n32421;
  assign n32423 = pi0590 & ~n32421;
  assign n32424 = ~n32422 & ~n32423;
  assign n32425 = pi3533 & pi9040;
  assign n32426 = pi3499 & ~pi9040;
  assign n32427 = ~n32425 & ~n32426;
  assign n32428 = ~pi0596 & ~n32427;
  assign n32429 = pi0596 & ~n32425;
  assign n32430 = ~n32426 & n32429;
  assign n32431 = ~n32428 & ~n32430;
  assign n32432 = ~n32424 & ~n32431;
  assign n32433 = ~n32418 & n32432;
  assign n32434 = pi3538 & pi9040;
  assign n32435 = pi3530 & ~pi9040;
  assign n32436 = ~n32434 & ~n32435;
  assign n32437 = ~pi0585 & n32436;
  assign n32438 = pi0585 & ~n32436;
  assign n32439 = ~n32437 & ~n32438;
  assign n32440 = n32431 & n32439;
  assign n32441 = ~n32424 & n32440;
  assign n32442 = n32418 & n32441;
  assign n32443 = n32431 & ~n32439;
  assign n32444 = ~n32418 & n32443;
  assign n32445 = ~n32442 & ~n32444;
  assign n32446 = ~n32433 & n32445;
  assign n32447 = n32412 & ~n32446;
  assign n32448 = ~n32418 & n32424;
  assign n32449 = n32439 & n32448;
  assign n32450 = ~n32431 & n32439;
  assign n32451 = ~n32424 & n32450;
  assign n32452 = n32418 & n32451;
  assign n32453 = ~n32449 & ~n32452;
  assign n32454 = n32424 & n32440;
  assign n32455 = ~n32424 & n32443;
  assign n32456 = ~n32454 & ~n32455;
  assign n32457 = n32453 & n32456;
  assign n32458 = ~n32405 & ~n32457;
  assign n32459 = ~n32431 & ~n32439;
  assign n32460 = n32424 & n32459;
  assign n32461 = n32418 & n32460;
  assign n32462 = ~n32458 & ~n32461;
  assign n32463 = ~n32411 & ~n32462;
  assign n32464 = ~n32447 & ~n32463;
  assign n32465 = ~n32405 & ~n32418;
  assign n32466 = ~n32424 & n32465;
  assign n32467 = ~n32439 & n32466;
  assign n32468 = ~n32418 & n32454;
  assign n32469 = ~n32467 & ~n32468;
  assign n32470 = ~n32443 & ~n32450;
  assign n32471 = n32418 & ~n32470;
  assign n32472 = n32424 & n32450;
  assign n32473 = ~n32471 & ~n32472;
  assign n32474 = n32405 & ~n32473;
  assign n32475 = ~n32424 & n32459;
  assign n32476 = ~n32433 & ~n32475;
  assign n32477 = ~n32442 & n32476;
  assign n32478 = ~n32405 & ~n32477;
  assign n32479 = ~n32474 & ~n32478;
  assign n32480 = n32405 & ~n32418;
  assign n32481 = n32440 & n32480;
  assign n32482 = n32418 & n32424;
  assign n32483 = n32439 & n32482;
  assign n32484 = ~n32431 & n32483;
  assign n32485 = n32424 & n32431;
  assign n32486 = ~n32439 & n32485;
  assign n32487 = n32418 & n32486;
  assign n32488 = ~n32484 & ~n32487;
  assign n32489 = ~n32439 & n32448;
  assign n32490 = ~n32431 & n32489;
  assign n32491 = n32488 & ~n32490;
  assign n32492 = ~n32481 & n32491;
  assign n32493 = n32479 & n32492;
  assign n32494 = n32411 & ~n32493;
  assign n32495 = n32469 & ~n32494;
  assign n32496 = n32464 & n32495;
  assign n32497 = pi0613 & ~n32496;
  assign n32498 = ~pi0613 & n32469;
  assign n32499 = n32464 & n32498;
  assign n32500 = ~n32494 & n32499;
  assign po0648 = n32497 | n32500;
  assign n32502 = n32264 & n32293;
  assign n32503 = ~n32277 & ~n32306;
  assign n32504 = n32502 & ~n32503;
  assign n32505 = n32284 & n32293;
  assign n32506 = n32277 & n32505;
  assign n32507 = ~n32504 & ~n32506;
  assign n32508 = n32299 & ~n32507;
  assign n32509 = ~n32264 & ~n32284;
  assign n32510 = n32276 & n32509;
  assign n32511 = n32270 & n32510;
  assign n32512 = ~n32340 & ~n32509;
  assign n32513 = ~n32293 & ~n32512;
  assign n32514 = ~n32264 & n32284;
  assign n32515 = ~n32276 & n32514;
  assign n32516 = n32270 & n32515;
  assign n32517 = ~n32513 & ~n32516;
  assign n32518 = ~n32511 & n32517;
  assign n32519 = n32299 & ~n32518;
  assign n32520 = ~n32508 & ~n32519;
  assign n32521 = n32276 & n32303;
  assign n32522 = ~n32270 & n32521;
  assign n32523 = ~n32264 & n32328;
  assign n32524 = ~n32522 & ~n32523;
  assign n32525 = n32293 & ~n32524;
  assign n32526 = n32264 & n32307;
  assign n32527 = ~n32264 & n32340;
  assign n32528 = ~n32526 & ~n32527;
  assign n32529 = ~n32293 & ~n32528;
  assign n32530 = ~n32302 & ~n32340;
  assign n32531 = n32264 & ~n32530;
  assign n32532 = ~n32328 & ~n32531;
  assign n32533 = n32293 & ~n32532;
  assign n32534 = ~n32264 & n32276;
  assign n32535 = n32293 & n32534;
  assign n32536 = n32284 & n32535;
  assign n32537 = ~n32276 & ~n32284;
  assign n32538 = ~n32328 & ~n32537;
  assign n32539 = ~n32264 & ~n32538;
  assign n32540 = n32264 & ~n32293;
  assign n32541 = n32305 & n32540;
  assign n32542 = n32284 & n32541;
  assign n32543 = ~n32539 & ~n32542;
  assign n32544 = ~n32536 & n32543;
  assign n32545 = ~n32533 & n32544;
  assign n32546 = ~n32522 & n32545;
  assign n32547 = ~n32299 & ~n32546;
  assign n32548 = ~n32529 & ~n32547;
  assign n32549 = ~n32525 & n32548;
  assign n32550 = n32520 & n32549;
  assign n32551 = pi0619 & n32550;
  assign n32552 = ~pi0619 & ~n32550;
  assign po0649 = n32551 | n32552;
  assign n32554 = ~n31988 & n32033;
  assign n32555 = ~n32018 & ~n32061;
  assign n32556 = ~n31976 & ~n32555;
  assign n32557 = ~n32554 & ~n32556;
  assign n32558 = ~n32056 & n32557;
  assign n32559 = n31976 & n31982;
  assign n32560 = n32003 & n32559;
  assign n32561 = ~n32044 & ~n32560;
  assign n32562 = ~n32009 & n32561;
  assign n32563 = n32558 & n32562;
  assign n32564 = n32028 & ~n32563;
  assign n32565 = ~n32002 & n32036;
  assign n32566 = n31982 & n32565;
  assign n32567 = ~n32034 & ~n32566;
  assign n32568 = ~n31976 & n32003;
  assign n32569 = n31982 & n32043;
  assign n32570 = ~n32568 & ~n32569;
  assign n32571 = ~n31982 & n32008;
  assign n32572 = ~n32048 & ~n32571;
  assign n32573 = ~n31994 & n32002;
  assign n32574 = n31982 & ~n31988;
  assign n32575 = ~n32573 & ~n32574;
  assign n32576 = ~n32013 & n32575;
  assign n32577 = n31976 & ~n32576;
  assign n32578 = n32572 & ~n32577;
  assign n32579 = n32570 & n32578;
  assign n32580 = n32567 & n32579;
  assign n32581 = ~n32028 & ~n32580;
  assign n32582 = ~n32564 & ~n32581;
  assign n32583 = pi0626 & ~n32582;
  assign n32584 = ~pi0626 & ~n32564;
  assign n32585 = ~n32581 & n32584;
  assign po0650 = n32583 | n32585;
  assign n32587 = ~n31793 & n31823;
  assign n32588 = n31793 & n31834;
  assign n32589 = ~n31820 & ~n32588;
  assign n32590 = n31765 & ~n32589;
  assign n32591 = ~n32587 & ~n32590;
  assign n32592 = ~n31765 & ~n31793;
  assign n32593 = ~n31785 & n32592;
  assign n32594 = n31779 & n32593;
  assign n32595 = n31801 & n31835;
  assign n32596 = ~n32594 & ~n32595;
  assign n32597 = ~n31765 & n31799;
  assign n32598 = n32596 & ~n32597;
  assign n32599 = ~n31797 & ~n31809;
  assign n32600 = n31785 & n31841;
  assign n32601 = n32599 & ~n32600;
  assign n32602 = n32598 & n32601;
  assign n32603 = n32591 & n32602;
  assign n32604 = ~n31832 & ~n32603;
  assign n32605 = ~n31796 & ~n31820;
  assign n32606 = n31793 & ~n32605;
  assign n32607 = n31779 & n31838;
  assign n32608 = ~n31849 & ~n32607;
  assign n32609 = n31772 & ~n31785;
  assign n32610 = n31793 & n32609;
  assign n32611 = n32608 & ~n32610;
  assign n32612 = n31765 & ~n32611;
  assign n32613 = ~n31793 & n31819;
  assign n32614 = n31779 & n31808;
  assign n32615 = ~n32613 & ~n32614;
  assign n32616 = ~n31765 & ~n32615;
  assign n32617 = ~n31793 & n31802;
  assign n32618 = ~n32616 & ~n32617;
  assign n32619 = ~n32612 & n32618;
  assign n32620 = ~n32606 & n32619;
  assign n32621 = n31832 & ~n32620;
  assign n32622 = n31765 & n31839;
  assign n32623 = ~n32621 & ~n32622;
  assign n32624 = n31814 & n32592;
  assign n32625 = ~n31785 & n32624;
  assign n32626 = n32623 & ~n32625;
  assign n32627 = ~n32604 & n32626;
  assign n32628 = ~pi0628 & ~n32627;
  assign n32629 = pi0628 & n32623;
  assign n32630 = ~n32604 & n32629;
  assign n32631 = ~n32625 & n32630;
  assign po0651 = n32628 | n32631;
  assign n32633 = ~n31931 & ~n32093;
  assign n32634 = n31903 & ~n32633;
  assign n32635 = ~n31927 & ~n31932;
  assign n32636 = ~n31924 & ~n32095;
  assign n32637 = n32635 & n32636;
  assign n32638 = n31893 & ~n32637;
  assign n32639 = ~n32634 & ~n32638;
  assign n32640 = ~n32084 & n32639;
  assign n32641 = n31868 & ~n32640;
  assign n32642 = ~n31893 & n31924;
  assign n32643 = n31893 & n32093;
  assign n32644 = ~n32642 & ~n32643;
  assign n32645 = n31899 & ~n32644;
  assign n32646 = n31899 & ~n32633;
  assign n32647 = ~n32642 & ~n32646;
  assign n32648 = ~n31880 & n32082;
  assign n32649 = ~n31958 & ~n32648;
  assign n32650 = ~n32095 & n32649;
  assign n32651 = ~n31899 & ~n32650;
  assign n32652 = n31893 & n32107;
  assign n32653 = ~n32651 & ~n32652;
  assign n32654 = n32647 & n32653;
  assign n32655 = ~n31868 & ~n32654;
  assign n32656 = ~n32645 & ~n32655;
  assign n32657 = ~n32641 & n32656;
  assign n32658 = ~pi0623 & ~n32657;
  assign n32659 = pi0623 & ~n32645;
  assign n32660 = ~n32641 & n32659;
  assign n32661 = ~n32655 & n32660;
  assign po0654 = n32658 | n32661;
  assign n32663 = n32418 & n32432;
  assign n32664 = ~n32455 & ~n32663;
  assign n32665 = ~n32468 & n32664;
  assign n32666 = ~n32405 & ~n32665;
  assign n32667 = ~n32418 & n32485;
  assign n32668 = ~n32439 & n32667;
  assign n32669 = ~n32418 & n32475;
  assign n32670 = n32424 & ~n32431;
  assign n32671 = ~n32440 & ~n32670;
  assign n32672 = n32418 & ~n32671;
  assign n32673 = ~n32669 & ~n32672;
  assign n32674 = ~n32668 & n32673;
  assign n32675 = n32405 & ~n32674;
  assign n32676 = ~n32666 & ~n32675;
  assign n32677 = n32411 & ~n32676;
  assign n32678 = ~n32431 & n32465;
  assign n32679 = ~n32418 & ~n32424;
  assign n32680 = n32431 & n32679;
  assign n32681 = ~n32663 & ~n32680;
  assign n32682 = n32405 & ~n32681;
  assign n32683 = ~n32481 & ~n32682;
  assign n32684 = ~n32418 & n32441;
  assign n32685 = ~n32487 & ~n32684;
  assign n32686 = ~n32405 & n32418;
  assign n32687 = n32485 & n32686;
  assign n32688 = ~n32405 & n32460;
  assign n32689 = ~n32687 & ~n32688;
  assign n32690 = n32685 & n32689;
  assign n32691 = n32683 & n32690;
  assign n32692 = ~n32678 & n32691;
  assign n32693 = ~n32411 & ~n32692;
  assign n32694 = n32472 & n32480;
  assign n32695 = ~n32424 & n32481;
  assign n32696 = ~n32694 & ~n32695;
  assign n32697 = ~n32405 & n32490;
  assign n32698 = n32696 & ~n32697;
  assign n32699 = n32418 & n32443;
  assign n32700 = ~n32418 & n32451;
  assign n32701 = ~n32699 & ~n32700;
  assign n32702 = ~n32405 & ~n32701;
  assign n32703 = n32698 & ~n32702;
  assign n32704 = ~n32693 & n32703;
  assign n32705 = ~n32677 & n32704;
  assign n32706 = ~pi0612 & ~n32705;
  assign n32707 = pi0612 & n32705;
  assign po0655 = n32706 | n32707;
  assign n32709 = ~n31772 & n31779;
  assign n32710 = ~n31765 & n32709;
  assign n32711 = n31793 & n32710;
  assign n32712 = ~n31793 & n32609;
  assign n32713 = ~n31800 & ~n32712;
  assign n32714 = ~n32614 & n32713;
  assign n32715 = ~n32711 & n32714;
  assign n32716 = n31765 & n31796;
  assign n32717 = n32715 & ~n32716;
  assign n32718 = n31832 & ~n32717;
  assign n32719 = ~n31850 & ~n32617;
  assign n32720 = n31765 & ~n32719;
  assign n32721 = ~n31832 & n31834;
  assign n32722 = ~n31765 & n32721;
  assign n32723 = n31772 & ~n31793;
  assign n32724 = ~n31779 & n32723;
  assign n32725 = ~n32609 & ~n32724;
  assign n32726 = ~n31802 & n32725;
  assign n32727 = n31765 & ~n32726;
  assign n32728 = ~n31772 & n31819;
  assign n32729 = ~n31793 & n32728;
  assign n32730 = ~n32727 & ~n32729;
  assign n32731 = ~n31832 & ~n32730;
  assign n32732 = ~n32722 & ~n32731;
  assign n32733 = ~n32720 & n32732;
  assign n32734 = ~n31793 & n31849;
  assign n32735 = ~n32588 & ~n32734;
  assign n32736 = ~n31797 & ~n31800;
  assign n32737 = n32735 & n32736;
  assign n32738 = ~n31765 & ~n32737;
  assign n32739 = n32733 & ~n32738;
  assign n32740 = ~n32718 & n32739;
  assign n32741 = ~pi0637 & ~n32740;
  assign n32742 = pi0637 & n32733;
  assign n32743 = ~n32718 & n32742;
  assign n32744 = ~n32738 & n32743;
  assign po0656 = n32741 | n32744;
  assign n32746 = pi3521 & ~pi9040;
  assign n32747 = pi3530 & pi9040;
  assign n32748 = ~n32746 & ~n32747;
  assign n32749 = ~pi0596 & ~n32748;
  assign n32750 = pi0596 & n32748;
  assign n32751 = ~n32749 & ~n32750;
  assign n32752 = pi3519 & pi9040;
  assign n32753 = pi3533 & ~pi9040;
  assign n32754 = ~n32752 & ~n32753;
  assign n32755 = ~pi0603 & n32754;
  assign n32756 = pi0603 & ~n32754;
  assign n32757 = ~n32755 & ~n32756;
  assign n32758 = pi3531 & pi9040;
  assign n32759 = pi3539 & ~pi9040;
  assign n32760 = ~n32758 & ~n32759;
  assign n32761 = ~pi0606 & ~n32760;
  assign n32762 = pi0606 & ~n32758;
  assign n32763 = ~n32759 & n32762;
  assign n32764 = ~n32761 & ~n32763;
  assign n32765 = pi3517 & pi9040;
  assign n32766 = pi3484 & ~pi9040;
  assign n32767 = ~n32765 & ~n32766;
  assign n32768 = pi0583 & n32767;
  assign n32769 = ~pi0583 & ~n32767;
  assign n32770 = ~n32768 & ~n32769;
  assign n32771 = pi3520 & pi9040;
  assign n32772 = pi3522 & ~pi9040;
  assign n32773 = ~n32771 & ~n32772;
  assign n32774 = pi0590 & n32773;
  assign n32775 = ~pi0590 & ~n32773;
  assign n32776 = ~n32774 & ~n32775;
  assign n32777 = n32770 & ~n32776;
  assign n32778 = n32764 & n32777;
  assign n32779 = ~n32757 & n32778;
  assign n32780 = n32757 & n32770;
  assign n32781 = n32776 & n32780;
  assign n32782 = pi3516 & pi9040;
  assign n32783 = pi3526 & ~pi9040;
  assign n32784 = ~n32782 & ~n32783;
  assign n32785 = pi0587 & n32784;
  assign n32786 = ~pi0587 & ~n32784;
  assign n32787 = ~n32785 & ~n32786;
  assign n32788 = ~n32764 & n32780;
  assign n32789 = n32764 & n32776;
  assign n32790 = ~n32770 & n32789;
  assign n32791 = ~n32788 & ~n32790;
  assign n32792 = ~n32787 & ~n32791;
  assign n32793 = ~n32781 & ~n32792;
  assign n32794 = n32770 & n32789;
  assign n32795 = ~n32764 & ~n32770;
  assign n32796 = ~n32770 & ~n32776;
  assign n32797 = n32757 & n32796;
  assign n32798 = ~n32764 & ~n32776;
  assign n32799 = ~n32757 & n32798;
  assign n32800 = ~n32797 & ~n32799;
  assign n32801 = ~n32795 & n32800;
  assign n32802 = ~n32794 & n32801;
  assign n32803 = n32787 & ~n32802;
  assign n32804 = n32793 & ~n32803;
  assign n32805 = ~n32779 & n32804;
  assign n32806 = n32751 & ~n32805;
  assign n32807 = ~n32764 & n32776;
  assign n32808 = ~n32770 & n32807;
  assign n32809 = n32757 & n32808;
  assign n32810 = ~n32770 & n32798;
  assign n32811 = ~n32757 & n32810;
  assign n32812 = ~n32779 & ~n32811;
  assign n32813 = ~n32809 & n32812;
  assign n32814 = n32787 & ~n32813;
  assign n32815 = ~n32806 & ~n32814;
  assign n32816 = n32757 & n32794;
  assign n32817 = ~n32757 & ~n32770;
  assign n32818 = ~n32787 & n32817;
  assign n32819 = n32764 & n32818;
  assign n32820 = n32770 & n32807;
  assign n32821 = ~n32757 & n32820;
  assign n32822 = n32777 & n32787;
  assign n32823 = n32757 & n32822;
  assign n32824 = ~n32821 & ~n32823;
  assign n32825 = ~n32764 & n32770;
  assign n32826 = ~n32757 & n32825;
  assign n32827 = n32764 & ~n32776;
  assign n32828 = ~n32770 & n32827;
  assign n32829 = ~n32826 & ~n32828;
  assign n32830 = ~n32787 & ~n32829;
  assign n32831 = ~n32787 & n32795;
  assign n32832 = n32757 & n32831;
  assign n32833 = ~n32830 & ~n32832;
  assign n32834 = n32824 & n32833;
  assign n32835 = ~n32751 & ~n32834;
  assign n32836 = ~n32819 & ~n32835;
  assign n32837 = ~n32816 & n32836;
  assign n32838 = n32815 & n32837;
  assign n32839 = ~pi0609 & ~n32838;
  assign n32840 = ~n32806 & ~n32816;
  assign n32841 = ~n32814 & n32840;
  assign n32842 = n32836 & n32841;
  assign n32843 = pi0609 & n32842;
  assign po0657 = n32839 | n32843;
  assign n32845 = n32757 & ~n32787;
  assign n32846 = n32764 & n32845;
  assign n32847 = n32770 & n32798;
  assign n32848 = ~n32757 & n32847;
  assign n32849 = ~n32757 & n32808;
  assign n32850 = ~n32848 & ~n32849;
  assign n32851 = n32757 & ~n32770;
  assign n32852 = ~n32776 & n32851;
  assign n32853 = ~n32764 & n32852;
  assign n32854 = ~n32790 & ~n32853;
  assign n32855 = n32787 & ~n32854;
  assign n32856 = n32850 & ~n32855;
  assign n32857 = ~n32846 & n32856;
  assign n32858 = n32751 & ~n32857;
  assign n32859 = ~n32757 & n32764;
  assign n32860 = ~n32770 & n32859;
  assign n32861 = ~n32776 & n32860;
  assign n32862 = ~n32787 & n32861;
  assign n32863 = n32757 & n32787;
  assign n32864 = n32828 & n32863;
  assign n32865 = ~n32788 & ~n32864;
  assign n32866 = ~n32790 & ~n32820;
  assign n32867 = n32757 & n32807;
  assign n32868 = n32866 & ~n32867;
  assign n32869 = ~n32787 & ~n32868;
  assign n32870 = n32787 & n32794;
  assign n32871 = n32812 & ~n32870;
  assign n32872 = ~n32869 & n32871;
  assign n32873 = n32865 & n32872;
  assign n32874 = ~n32751 & ~n32873;
  assign n32875 = ~n32862 & ~n32874;
  assign n32876 = ~n32858 & n32875;
  assign n32877 = n32820 & n32863;
  assign n32878 = ~n32757 & n32822;
  assign n32879 = ~n32877 & ~n32878;
  assign n32880 = n32787 & n32849;
  assign n32881 = n32879 & ~n32880;
  assign n32882 = n32876 & n32881;
  assign n32883 = ~pi0615 & ~n32882;
  assign n32884 = pi0615 & n32881;
  assign n32885 = n32875 & n32884;
  assign n32886 = ~n32858 & n32885;
  assign po0658 = n32883 | n32886;
  assign n32888 = ~n31794 & ~n31800;
  assign n32889 = ~n31765 & ~n32888;
  assign n32890 = ~n31856 & ~n32889;
  assign n32891 = ~n31772 & ~n31779;
  assign n32892 = n31765 & n32891;
  assign n32893 = n31793 & n32892;
  assign n32894 = ~n31765 & n31786;
  assign n32895 = n31793 & n32894;
  assign n32896 = ~n32597 & ~n32895;
  assign n32897 = n31779 & n32723;
  assign n32898 = n31793 & n31819;
  assign n32899 = ~n32897 & ~n32898;
  assign n32900 = ~n32891 & n32899;
  assign n32901 = n31765 & ~n32900;
  assign n32902 = ~n31803 & ~n32901;
  assign n32903 = n32896 & n32902;
  assign n32904 = ~n31832 & ~n32903;
  assign n32905 = ~n32893 & ~n32904;
  assign n32906 = ~n31820 & ~n31839;
  assign n32907 = ~n31849 & n32906;
  assign n32908 = ~n31765 & ~n32907;
  assign n32909 = ~n31793 & n31799;
  assign n32910 = ~n31823 & ~n32909;
  assign n32911 = n31765 & ~n32910;
  assign n32912 = ~n32908 & ~n32911;
  assign n32913 = ~n32607 & n32912;
  assign n32914 = ~n31809 & ~n31850;
  assign n32915 = n32913 & n32914;
  assign n32916 = n31832 & ~n32915;
  assign n32917 = n32905 & ~n32916;
  assign n32918 = n32890 & n32917;
  assign n32919 = ~pi0635 & ~n32918;
  assign n32920 = pi0635 & n32905;
  assign n32921 = n32890 & n32920;
  assign n32922 = ~n32916 & n32921;
  assign po0659 = n32919 | n32922;
  assign n32924 = pi3493 & pi9040;
  assign n32925 = pi3502 & ~pi9040;
  assign n32926 = ~n32924 & ~n32925;
  assign n32927 = pi0602 & n32926;
  assign n32928 = ~pi0602 & ~n32926;
  assign n32929 = ~n32927 & ~n32928;
  assign n32930 = pi3507 & pi9040;
  assign n32931 = pi3505 & ~pi9040;
  assign n32932 = ~n32930 & ~n32931;
  assign n32933 = ~pi0575 & n32932;
  assign n32934 = pi0575 & ~n32932;
  assign n32935 = ~n32933 & ~n32934;
  assign n32936 = pi3496 & pi9040;
  assign n32937 = pi3559 & ~pi9040;
  assign n32938 = ~n32936 & ~n32937;
  assign n32939 = ~pi0605 & n32938;
  assign n32940 = pi0605 & ~n32938;
  assign n32941 = ~n32939 & ~n32940;
  assign n32942 = ~n32935 & ~n32941;
  assign n32943 = n32929 & n32942;
  assign n32944 = ~pi0605 & ~n32938;
  assign n32945 = pi0605 & n32938;
  assign n32946 = ~n32944 & ~n32945;
  assign n32947 = ~n32935 & ~n32946;
  assign n32948 = ~n32929 & n32947;
  assign n32949 = ~n32943 & ~n32948;
  assign n32950 = pi3513 & pi9040;
  assign n32951 = pi3527 & ~pi9040;
  assign n32952 = ~n32950 & ~n32951;
  assign n32953 = pi0597 & n32952;
  assign n32954 = ~pi0597 & ~n32952;
  assign n32955 = ~n32953 & ~n32954;
  assign n32956 = n32929 & ~n32955;
  assign n32957 = n32946 & n32956;
  assign n32958 = n32949 & ~n32957;
  assign n32959 = pi3492 & pi9040;
  assign n32960 = pi3506 & ~pi9040;
  assign n32961 = ~n32959 & ~n32960;
  assign n32962 = pi0577 & n32961;
  assign n32963 = ~pi0577 & ~n32961;
  assign n32964 = ~n32962 & ~n32963;
  assign n32965 = pi3503 & pi9040;
  assign n32966 = pi3490 & ~pi9040;
  assign n32967 = ~n32965 & ~n32966;
  assign n32968 = ~pi0582 & n32967;
  assign n32969 = pi0582 & ~n32967;
  assign n32970 = ~n32968 & ~n32969;
  assign n32971 = ~n32964 & ~n32970;
  assign n32972 = ~n32958 & n32971;
  assign n32973 = n32935 & ~n32946;
  assign n32974 = n32929 & n32973;
  assign n32975 = ~n32970 & n32974;
  assign n32976 = n32955 & n32975;
  assign n32977 = n32929 & n32947;
  assign n32978 = n32964 & n32977;
  assign n32979 = ~n32929 & n32946;
  assign n32980 = n32935 & ~n32941;
  assign n32981 = n32955 & n32980;
  assign n32982 = ~n32979 & ~n32981;
  assign n32983 = n32964 & ~n32982;
  assign n32984 = ~n32978 & ~n32983;
  assign n32985 = ~n32970 & ~n32984;
  assign n32986 = ~n32976 & ~n32985;
  assign n32987 = ~n32929 & n32955;
  assign n32988 = n32946 & n32987;
  assign n32989 = ~n32929 & ~n32955;
  assign n32990 = ~n32946 & n32989;
  assign n32991 = n32935 & n32990;
  assign n32992 = ~n32988 & ~n32991;
  assign n32993 = n32964 & ~n32992;
  assign n32994 = n32986 & ~n32993;
  assign n32995 = n32955 & ~n32964;
  assign n32996 = n32980 & n32995;
  assign n32997 = n32929 & n32996;
  assign n32998 = ~n32942 & ~n32973;
  assign n32999 = n32956 & ~n32998;
  assign n33000 = ~n32935 & n32990;
  assign n33001 = ~n32999 & ~n33000;
  assign n33002 = ~n32929 & n32980;
  assign n33003 = ~n32955 & ~n32964;
  assign n33004 = n33002 & n33003;
  assign n33005 = n32987 & ~n32998;
  assign n33006 = n32955 & n32977;
  assign n33007 = ~n33005 & ~n33006;
  assign n33008 = ~n33004 & n33007;
  assign n33009 = n33001 & n33008;
  assign n33010 = ~n32997 & n33009;
  assign n33011 = ~n32955 & n32964;
  assign n33012 = n32929 & n33011;
  assign n33013 = n32935 & n33012;
  assign n33014 = n33010 & ~n33013;
  assign n33015 = n32970 & ~n33014;
  assign n33016 = n32994 & ~n33015;
  assign n33017 = ~n32972 & n33016;
  assign n33018 = ~pi0622 & ~n33017;
  assign n33019 = pi0622 & n32994;
  assign n33020 = ~n32972 & n33019;
  assign n33021 = ~n33015 & n33020;
  assign po0660 = n33018 | n33021;
  assign n33023 = n32929 & n32980;
  assign n33024 = n32964 & n33023;
  assign n33025 = ~n32955 & n33024;
  assign n33026 = n32947 & n33011;
  assign n33027 = ~n32929 & n33026;
  assign n33028 = ~n33025 & ~n33027;
  assign n33029 = ~n33000 & ~n33004;
  assign n33030 = ~n32935 & n32955;
  assign n33031 = n32929 & n33030;
  assign n33032 = ~n32981 & ~n33031;
  assign n33033 = n32964 & ~n33032;
  assign n33034 = ~n32964 & ~n32989;
  assign n33035 = ~n32998 & n33034;
  assign n33036 = ~n32929 & ~n32980;
  assign n33037 = n32964 & n33036;
  assign n33038 = ~n32955 & n33037;
  assign n33039 = ~n33035 & ~n33038;
  assign n33040 = ~n33033 & n33039;
  assign n33041 = n33029 & n33040;
  assign n33042 = ~n32970 & ~n33041;
  assign n33043 = n33028 & ~n33042;
  assign n33044 = n32943 & ~n32964;
  assign n33045 = n32955 & n33044;
  assign n33046 = ~n32964 & n32970;
  assign n33047 = n32989 & ~n32998;
  assign n33048 = ~n32981 & ~n33047;
  assign n33049 = ~n32977 & n33048;
  assign n33050 = n33046 & ~n33049;
  assign n33051 = n32948 & n32955;
  assign n33052 = ~n32929 & n33030;
  assign n33053 = n32955 & n32973;
  assign n33054 = ~n33052 & ~n33053;
  assign n33055 = ~n32955 & n32980;
  assign n33056 = ~n32974 & ~n33055;
  assign n33057 = n33054 & n33056;
  assign n33058 = n32964 & ~n33057;
  assign n33059 = ~n33051 & ~n33058;
  assign n33060 = n32970 & ~n33059;
  assign n33061 = ~n33050 & ~n33060;
  assign n33062 = ~n33045 & n33061;
  assign n33063 = n33043 & n33062;
  assign n33064 = pi0630 & ~n33063;
  assign n33065 = ~pi0630 & n33043;
  assign n33066 = n33062 & n33065;
  assign po0661 = n33064 | n33066;
  assign n33068 = n32264 & ~n32276;
  assign n33069 = n32284 & n33068;
  assign n33070 = ~n32306 & ~n33069;
  assign n33071 = n32293 & ~n33070;
  assign n33072 = n32264 & n32327;
  assign n33073 = ~n32515 & ~n33072;
  assign n33074 = ~n32293 & ~n33073;
  assign n33075 = ~n32264 & n32322;
  assign n33076 = ~n32536 & ~n33075;
  assign n33077 = ~n32304 & n33076;
  assign n33078 = ~n33074 & n33077;
  assign n33079 = ~n33071 & n33078;
  assign n33080 = ~n32511 & ~n32522;
  assign n33081 = n33079 & n33080;
  assign n33082 = n32299 & ~n33081;
  assign n33083 = n32302 & n32509;
  assign n33084 = n32308 & ~n33083;
  assign n33085 = ~n32293 & ~n33084;
  assign n33086 = ~n32264 & n32286;
  assign n33087 = ~n33085 & ~n33086;
  assign n33088 = n32270 & n32313;
  assign n33089 = n32264 & n32305;
  assign n33090 = ~n33088 & ~n33089;
  assign n33091 = ~n32293 & ~n33090;
  assign n33092 = ~n32293 & n32327;
  assign n33093 = ~n32264 & n33092;
  assign n33094 = ~n33091 & ~n33093;
  assign n33095 = n33087 & n33094;
  assign n33096 = ~n32299 & ~n33095;
  assign n33097 = ~n32322 & ~n32329;
  assign n33098 = ~n32516 & n33097;
  assign n33099 = n32337 & ~n33098;
  assign n33100 = ~n33096 & ~n33099;
  assign n33101 = ~n32304 & ~n32511;
  assign n33102 = n32293 & ~n33101;
  assign n33103 = n33100 & ~n33102;
  assign n33104 = ~n33082 & n33103;
  assign n33105 = ~pi0627 & n33104;
  assign n33106 = pi0627 & ~n33104;
  assign po0662 = n33105 | n33106;
  assign n33108 = ~n32167 & n32205;
  assign n33109 = n32179 & n32218;
  assign n33110 = ~n32236 & ~n33109;
  assign n33111 = n32194 & ~n33110;
  assign n33112 = ~n33108 & ~n33111;
  assign n33113 = n32195 & n32237;
  assign n33114 = ~n32194 & n32203;
  assign n33115 = ~n33113 & ~n33114;
  assign n33116 = n33112 & n33115;
  assign n33117 = n32179 & n32223;
  assign n33118 = ~n32351 & ~n33117;
  assign n33119 = ~n32385 & n33118;
  assign n33120 = n33116 & n33119;
  assign n33121 = ~n32161 & ~n33120;
  assign n33122 = ~n32225 & ~n32236;
  assign n33123 = ~n32387 & n33122;
  assign n33124 = ~n32194 & ~n33123;
  assign n33125 = n32167 & n32197;
  assign n33126 = ~n32359 & ~n33125;
  assign n33127 = ~n32251 & n33126;
  assign n33128 = n32194 & n32212;
  assign n33129 = n33127 & ~n33128;
  assign n33130 = ~n33124 & n33129;
  assign n33131 = n32161 & ~n33130;
  assign n33132 = ~n32375 & ~n32380;
  assign n33133 = ~n32351 & n33126;
  assign n33134 = ~n32194 & ~n33133;
  assign n33135 = n33132 & ~n33134;
  assign n33136 = ~n33131 & n33135;
  assign n33137 = ~n33121 & n33136;
  assign n33138 = pi0625 & ~n33137;
  assign n33139 = ~pi0625 & n33137;
  assign po0663 = n33138 | n33139;
  assign n33141 = ~n32472 & ~n32475;
  assign n33142 = n32405 & ~n33141;
  assign n33143 = n32418 & n32455;
  assign n33144 = ~n33142 & ~n33143;
  assign n33145 = n32418 & n32431;
  assign n33146 = ~n32485 & ~n33145;
  assign n33147 = ~n32451 & n33146;
  assign n33148 = ~n32405 & ~n33147;
  assign n33149 = n33144 & ~n33148;
  assign n33150 = ~n32411 & ~n33149;
  assign n33151 = ~n32418 & n32486;
  assign n33152 = n32405 & n33151;
  assign n33153 = ~n32695 & ~n33152;
  assign n33154 = ~n32697 & n33153;
  assign n33155 = ~n32405 & n32431;
  assign n33156 = n32679 & n33155;
  assign n33157 = n32418 & n32475;
  assign n33158 = n32405 & n32485;
  assign n33159 = ~n33157 & ~n33158;
  assign n33160 = ~n32484 & n33159;
  assign n33161 = ~n33156 & n33160;
  assign n33162 = n32439 & n32679;
  assign n33163 = ~n32490 & ~n33162;
  assign n33164 = n33161 & n33163;
  assign n33165 = ~n32688 & n33164;
  assign n33166 = n32411 & ~n33165;
  assign n33167 = n33154 & ~n33166;
  assign n33168 = ~n33150 & n33167;
  assign n33169 = ~pi0620 & ~n33168;
  assign n33170 = pi0620 & n33154;
  assign n33171 = ~n33150 & n33170;
  assign n33172 = ~n33166 & n33171;
  assign po0664 = n33169 | n33172;
  assign n33174 = ~n32211 & ~n32219;
  assign n33175 = n32161 & ~n33174;
  assign n33176 = n32187 & ~n32194;
  assign n33177 = ~n32224 & ~n32363;
  assign n33178 = ~n32194 & ~n33177;
  assign n33179 = ~n33176 & ~n33178;
  assign n33180 = n32161 & ~n33179;
  assign n33181 = ~n33175 & ~n33180;
  assign n33182 = n32210 & n32360;
  assign n33183 = ~n32362 & ~n33182;
  assign n33184 = ~n32227 & ~n32388;
  assign n33185 = n32194 & ~n33184;
  assign n33186 = n32161 & n33185;
  assign n33187 = n33183 & ~n33186;
  assign n33188 = ~n32167 & n32210;
  assign n33189 = ~n32167 & n32202;
  assign n33190 = ~n32353 & ~n33189;
  assign n33191 = n32194 & ~n33190;
  assign n33192 = ~n32225 & ~n32359;
  assign n33193 = ~n32167 & n32209;
  assign n33194 = ~n32249 & ~n33193;
  assign n33195 = ~n32194 & ~n33194;
  assign n33196 = n33192 & ~n33195;
  assign n33197 = ~n33191 & n33196;
  assign n33198 = ~n33188 & n33197;
  assign n33199 = ~n32161 & ~n33198;
  assign n33200 = ~n32385 & n33126;
  assign n33201 = n32194 & ~n33200;
  assign n33202 = ~n33199 & ~n33201;
  assign n33203 = n33187 & n33202;
  assign n33204 = n33181 & n33203;
  assign n33205 = ~pi0633 & ~n33204;
  assign n33206 = pi0633 & n33187;
  assign n33207 = n33181 & n33206;
  assign n33208 = n33202 & n33207;
  assign po0665 = n33205 | n33208;
  assign n33210 = ~n31982 & n32036;
  assign n33211 = ~n32571 & ~n33210;
  assign n33212 = ~n31976 & n33211;
  assign n33213 = n31982 & n32016;
  assign n33214 = ~n31995 & ~n32005;
  assign n33215 = n32002 & ~n33214;
  assign n33216 = n31988 & n32059;
  assign n33217 = n31982 & n32005;
  assign n33218 = ~n33216 & ~n33217;
  assign n33219 = ~n33215 & n33218;
  assign n33220 = n31976 & n33219;
  assign n33221 = ~n33213 & n33220;
  assign n33222 = ~n33212 & ~n33221;
  assign n33223 = n31982 & n33215;
  assign n33224 = ~n32566 & ~n33223;
  assign n33225 = ~n33222 & n33224;
  assign n33226 = n32028 & ~n33225;
  assign n33227 = ~n31976 & ~n33214;
  assign n33228 = ~n31982 & n33227;
  assign n33229 = n31982 & n32007;
  assign n33230 = ~n32042 & ~n33229;
  assign n33231 = ~n31976 & ~n33230;
  assign n33232 = ~n32002 & n33227;
  assign n33233 = ~n33231 & ~n33232;
  assign n33234 = ~n33228 & n33233;
  assign n33235 = ~n32028 & ~n33234;
  assign n33236 = ~n33226 & ~n33235;
  assign n33237 = n31976 & ~n33211;
  assign n33238 = ~n32034 & ~n33237;
  assign n33239 = ~n32028 & ~n33238;
  assign n33240 = ~n31976 & n32034;
  assign n33241 = n31976 & ~n33224;
  assign n33242 = ~n33240 & ~n33241;
  assign n33243 = ~n33239 & n33242;
  assign n33244 = n33236 & n33243;
  assign n33245 = pi0641 & ~n33244;
  assign n33246 = ~pi0641 & n33243;
  assign n33247 = ~n33235 & n33246;
  assign n33248 = ~n33226 & n33247;
  assign po0666 = n33245 | n33248;
  assign n33250 = ~n32929 & n32942;
  assign n33251 = ~n33023 & ~n33250;
  assign n33252 = n32964 & ~n33251;
  assign n33253 = ~n32955 & n32973;
  assign n33254 = ~n32943 & ~n33253;
  assign n33255 = ~n33002 & n33254;
  assign n33256 = ~n32964 & ~n33255;
  assign n33257 = ~n33252 & ~n33256;
  assign n33258 = ~n32978 & ~n32991;
  assign n33259 = n33257 & n33258;
  assign n33260 = n32970 & ~n33259;
  assign n33261 = n32955 & n33023;
  assign n33262 = n32947 & ~n32955;
  assign n33263 = ~n33053 & ~n33262;
  assign n33264 = ~n32964 & ~n33263;
  assign n33265 = ~n33261 & ~n33264;
  assign n33266 = n32964 & n32974;
  assign n33267 = n32949 & ~n33266;
  assign n33268 = ~n33002 & n33267;
  assign n33269 = ~n32955 & ~n33268;
  assign n33270 = n33265 & ~n33269;
  assign n33271 = ~n32970 & ~n33270;
  assign n33272 = ~n33260 & ~n33271;
  assign n33273 = ~n32929 & n33053;
  assign n33274 = ~n33006 & ~n33273;
  assign n33275 = n32964 & ~n33274;
  assign n33276 = ~n32929 & ~n32935;
  assign n33277 = n32995 & n33276;
  assign n33278 = ~n33275 & ~n33277;
  assign n33279 = n33272 & n33278;
  assign n33280 = ~pi0611 & ~n33279;
  assign n33281 = pi0611 & ~n33275;
  assign n33282 = n33272 & n33281;
  assign n33283 = ~n33277 & n33282;
  assign po0667 = n33280 | n33283;
  assign n33285 = n32286 & n32293;
  assign n33286 = ~n32264 & n32305;
  assign n33287 = ~n32319 & ~n33286;
  assign n33288 = n32293 & ~n33287;
  assign n33289 = ~n32293 & ~n32538;
  assign n33290 = ~n33288 & ~n33289;
  assign n33291 = ~n32526 & n33290;
  assign n33292 = n32299 & ~n33291;
  assign n33293 = ~n33285 & ~n33292;
  assign n33294 = ~n32284 & n32502;
  assign n33295 = ~n32514 & ~n33294;
  assign n33296 = ~n32270 & ~n33295;
  assign n33297 = ~n32304 & ~n33296;
  assign n33298 = ~n32515 & n33297;
  assign n33299 = ~n32293 & n32320;
  assign n33300 = n32264 & n32306;
  assign n33301 = ~n33299 & ~n33300;
  assign n33302 = n33298 & n33301;
  assign n33303 = ~n32299 & ~n33302;
  assign n33304 = ~n33075 & ~n33089;
  assign n33305 = ~n32293 & ~n33304;
  assign n33306 = ~n33303 & ~n33305;
  assign n33307 = n33293 & n33306;
  assign n33308 = ~pi0649 & ~n33307;
  assign n33309 = pi0649 & n33306;
  assign n33310 = ~n33292 & n33309;
  assign n33311 = ~n33285 & n33310;
  assign po0668 = n33308 | n33311;
  assign n33313 = ~n32974 & ~n33030;
  assign n33314 = n32971 & ~n33313;
  assign n33315 = ~n33053 & ~n33055;
  assign n33316 = n32964 & ~n33315;
  assign n33317 = ~n33027 & ~n33316;
  assign n33318 = ~n32970 & ~n33317;
  assign n33319 = n32955 & n33002;
  assign n33320 = ~n32946 & n32956;
  assign n33321 = ~n32942 & ~n33276;
  assign n33322 = n32955 & ~n33321;
  assign n33323 = ~n33320 & ~n33322;
  assign n33324 = n32964 & ~n33323;
  assign n33325 = ~n33319 & ~n33324;
  assign n33326 = ~n32955 & ~n33321;
  assign n33327 = ~n33023 & ~n33326;
  assign n33328 = ~n32964 & ~n33327;
  assign n33329 = ~n33047 & ~n33328;
  assign n33330 = n33325 & n33329;
  assign n33331 = n32970 & ~n33330;
  assign n33332 = ~n33318 & ~n33331;
  assign n33333 = n32964 & n32987;
  assign n33334 = n32942 & n33333;
  assign n33335 = n32929 & n32995;
  assign n33336 = ~n32946 & n33335;
  assign n33337 = ~n33334 & ~n33336;
  assign n33338 = n32929 & n32955;
  assign n33339 = ~n32942 & n33338;
  assign n33340 = ~n32970 & n33339;
  assign n33341 = n33337 & ~n33340;
  assign n33342 = n33332 & n33341;
  assign n33343 = ~n33314 & n33342;
  assign n33344 = pi0631 & ~n33343;
  assign n33345 = ~pi0631 & n33341;
  assign n33346 = ~n33314 & n33345;
  assign n33347 = n33332 & n33346;
  assign po0669 = n33344 | n33347;
  assign n33349 = ~n32418 & ~n32431;
  assign n33350 = ~n33162 & ~n33349;
  assign n33351 = n32405 & ~n33350;
  assign n33352 = n32418 & ~n32424;
  assign n33353 = ~n32439 & n33352;
  assign n33354 = ~n33351 & ~n33353;
  assign n33355 = ~n32405 & n32443;
  assign n33356 = ~n32418 & n33355;
  assign n33357 = ~n32700 & ~n33356;
  assign n33358 = n33354 & n33357;
  assign n33359 = n32411 & ~n33358;
  assign n33360 = ~n32441 & ~n32487;
  assign n33361 = ~n32418 & n32459;
  assign n33362 = n33360 & ~n33361;
  assign n33363 = ~n32405 & ~n33362;
  assign n33364 = n32443 & n32480;
  assign n33365 = ~n32468 & ~n33364;
  assign n33366 = ~n33363 & n33365;
  assign n33367 = ~n32451 & ~n32461;
  assign n33368 = n32405 & ~n33367;
  assign n33369 = n33366 & ~n33368;
  assign n33370 = ~n32411 & ~n33369;
  assign n33371 = ~n33359 & ~n33370;
  assign n33372 = ~n32418 & n32450;
  assign n33373 = n32418 & ~n32456;
  assign n33374 = ~n33372 & ~n33373;
  assign n33375 = n32405 & ~n33374;
  assign n33376 = ~n32441 & n33141;
  assign n33377 = n32686 & ~n33376;
  assign n33378 = ~n33375 & ~n33377;
  assign n33379 = n33371 & n33378;
  assign n33380 = ~pi0614 & ~n33379;
  assign n33381 = ~n33370 & n33378;
  assign n33382 = pi0614 & n33381;
  assign n33383 = ~n33359 & n33382;
  assign po0670 = n33380 | n33383;
  assign n33385 = n32757 & n32847;
  assign n33386 = ~n32808 & ~n32816;
  assign n33387 = ~n32757 & n32777;
  assign n33388 = n32757 & n32828;
  assign n33389 = ~n33387 & ~n33388;
  assign n33390 = n33386 & n33389;
  assign n33391 = ~n32787 & ~n33390;
  assign n33392 = ~n32757 & n32789;
  assign n33393 = ~n32788 & ~n33392;
  assign n33394 = ~n32810 & n33393;
  assign n33395 = n32787 & ~n33394;
  assign n33396 = n32776 & n32817;
  assign n33397 = n32764 & n33396;
  assign n33398 = ~n33395 & ~n33397;
  assign n33399 = ~n33391 & n33398;
  assign n33400 = ~n33385 & n33399;
  assign n33401 = ~n32751 & ~n33400;
  assign n33402 = ~n32757 & ~n32787;
  assign n33403 = n32794 & n33402;
  assign n33404 = ~n32787 & n32810;
  assign n33405 = ~n32787 & n32820;
  assign n33406 = ~n33404 & ~n33405;
  assign n33407 = n32757 & ~n33406;
  assign n33408 = ~n33403 & ~n33407;
  assign n33409 = n32757 & n32778;
  assign n33410 = ~n32861 & ~n33409;
  assign n33411 = ~n32757 & n32807;
  assign n33412 = n32757 & n32789;
  assign n33413 = ~n33411 & ~n33412;
  assign n33414 = ~n32778 & n33413;
  assign n33415 = ~n32808 & n33414;
  assign n33416 = n32787 & ~n33415;
  assign n33417 = n32757 & n32790;
  assign n33418 = ~n33416 & ~n33417;
  assign n33419 = n33410 & n33418;
  assign n33420 = n33408 & n33419;
  assign n33421 = n32751 & ~n33420;
  assign n33422 = ~n32787 & ~n32850;
  assign n33423 = ~n33421 & ~n33422;
  assign n33424 = ~n32811 & ~n33409;
  assign n33425 = n32787 & ~n33424;
  assign n33426 = n33423 & ~n33425;
  assign n33427 = ~n33401 & n33426;
  assign n33428 = pi0632 & ~n33427;
  assign n33429 = ~pi0632 & n33427;
  assign po0671 = n33428 | n33429;
  assign n33431 = ~n31976 & n32004;
  assign n33432 = n32059 & ~n33214;
  assign n33433 = ~n32008 & ~n33432;
  assign n33434 = ~n32566 & n33433;
  assign n33435 = n31976 & ~n33434;
  assign n33436 = n31982 & n32031;
  assign n33437 = ~n33435 & ~n33436;
  assign n33438 = ~n32002 & n32007;
  assign n33439 = ~n31982 & n32573;
  assign n33440 = ~n33438 & ~n33439;
  assign n33441 = ~n33217 & n33440;
  assign n33442 = ~n31976 & ~n33441;
  assign n33443 = n33437 & ~n33442;
  assign n33444 = n32028 & ~n33443;
  assign n33445 = ~n33431 & ~n33444;
  assign n33446 = ~n31982 & n32005;
  assign n33447 = ~n32565 & ~n33446;
  assign n33448 = ~n31976 & ~n33447;
  assign n33449 = ~n32009 & ~n33448;
  assign n33450 = ~n32004 & ~n32042;
  assign n33451 = n31982 & n32013;
  assign n33452 = ~n32573 & ~n33451;
  assign n33453 = ~n33438 & n33452;
  assign n33454 = n31976 & ~n33453;
  assign n33455 = ~n31982 & n32031;
  assign n33456 = ~n33454 & ~n33455;
  assign n33457 = n33450 & n33456;
  assign n33458 = n33449 & n33457;
  assign n33459 = ~n32028 & ~n33458;
  assign n33460 = ~n32064 & ~n33213;
  assign n33461 = n31976 & ~n33460;
  assign n33462 = ~n33459 & ~n33461;
  assign n33463 = n33445 & n33462;
  assign n33464 = pi0659 & n33463;
  assign n33465 = ~pi0659 & ~n33463;
  assign po0672 = n33464 | n33465;
  assign n33467 = ~n32853 & ~n33409;
  assign n33468 = ~n33397 & n33467;
  assign n33469 = ~n32787 & ~n33468;
  assign n33470 = ~n32864 & ~n32880;
  assign n33471 = ~n32778 & ~n32867;
  assign n33472 = n32787 & ~n33471;
  assign n33473 = ~n32770 & n32776;
  assign n33474 = ~n32795 & ~n33473;
  assign n33475 = ~n32757 & ~n33474;
  assign n33476 = ~n32757 & n32776;
  assign n33477 = ~n32790 & ~n33476;
  assign n33478 = ~n32798 & n33477;
  assign n33479 = ~n32787 & ~n33478;
  assign n33480 = ~n33475 & ~n33479;
  assign n33481 = ~n33472 & n33480;
  assign n33482 = ~n32751 & n33481;
  assign n33483 = ~n32847 & ~n33412;
  assign n33484 = n32787 & ~n33483;
  assign n33485 = ~n32816 & ~n32861;
  assign n33486 = ~n33405 & n33485;
  assign n33487 = n32751 & n33486;
  assign n33488 = ~n33484 & n33487;
  assign n33489 = ~n33482 & ~n33488;
  assign n33490 = n33470 & ~n33489;
  assign n33491 = ~n33469 & n33490;
  assign n33492 = ~pi0640 & ~n33491;
  assign n33493 = pi0640 & n33470;
  assign n33494 = ~n33469 & n33493;
  assign n33495 = ~n33489 & n33494;
  assign po0673 = n33492 | n33495;
  assign n33497 = pi3582 & pi9040;
  assign n33498 = pi3594 & ~pi9040;
  assign n33499 = ~n33497 & ~n33498;
  assign n33500 = pi0642 & n33499;
  assign n33501 = ~pi0642 & ~n33499;
  assign n33502 = ~n33500 & ~n33501;
  assign n33503 = pi3546 & pi9040;
  assign n33504 = pi3572 & ~pi9040;
  assign n33505 = ~n33503 & ~n33504;
  assign n33506 = ~pi0638 & ~n33505;
  assign n33507 = pi0638 & ~n33503;
  assign n33508 = ~n33504 & n33507;
  assign n33509 = ~n33506 & ~n33508;
  assign n33510 = pi3596 & pi9040;
  assign n33511 = pi3592 & ~pi9040;
  assign n33512 = ~n33510 & ~n33511;
  assign n33513 = ~pi0639 & n33512;
  assign n33514 = pi0639 & ~n33512;
  assign n33515 = ~n33513 & ~n33514;
  assign n33516 = pi3595 & pi9040;
  assign n33517 = pi3566 & ~pi9040;
  assign n33518 = ~n33516 & ~n33517;
  assign n33519 = pi0668 & n33518;
  assign n33520 = ~pi0668 & ~n33518;
  assign n33521 = ~n33519 & ~n33520;
  assign n33522 = ~n33515 & n33521;
  assign n33523 = ~n33509 & n33522;
  assign n33524 = pi3563 & pi9040;
  assign n33525 = pi3584 & ~pi9040;
  assign n33526 = ~n33524 & ~n33525;
  assign n33527 = ~pi0661 & n33526;
  assign n33528 = pi0661 & ~n33526;
  assign n33529 = ~n33527 & ~n33528;
  assign n33530 = n33523 & n33529;
  assign n33531 = n33515 & ~n33521;
  assign n33532 = ~n33509 & n33531;
  assign n33533 = n33529 & n33532;
  assign n33534 = ~n33530 & ~n33533;
  assign n33535 = n33509 & n33531;
  assign n33536 = ~n33529 & n33535;
  assign n33537 = n33515 & n33521;
  assign n33538 = ~n33509 & n33537;
  assign n33539 = ~n33529 & n33538;
  assign n33540 = ~n33536 & ~n33539;
  assign n33541 = n33534 & n33540;
  assign n33542 = n33502 & ~n33541;
  assign n33543 = ~n33509 & ~n33529;
  assign n33544 = ~n33515 & n33543;
  assign n33545 = ~n33521 & n33544;
  assign n33546 = ~n33538 & ~n33545;
  assign n33547 = n33502 & ~n33546;
  assign n33548 = ~n33515 & n33529;
  assign n33549 = ~n33502 & n33548;
  assign n33550 = n33509 & n33521;
  assign n33551 = ~n33529 & n33531;
  assign n33552 = ~n33550 & ~n33551;
  assign n33553 = ~n33502 & ~n33552;
  assign n33554 = ~n33549 & ~n33553;
  assign n33555 = ~n33515 & ~n33521;
  assign n33556 = n33509 & n33555;
  assign n33557 = n33529 & n33556;
  assign n33558 = n33554 & ~n33557;
  assign n33559 = ~n33515 & n33550;
  assign n33560 = ~n33529 & n33559;
  assign n33561 = n33558 & ~n33560;
  assign n33562 = ~n33547 & n33561;
  assign n33563 = ~pi3574 & ~pi9040;
  assign n33564 = ~pi3554 & pi9040;
  assign n33565 = ~n33563 & ~n33564;
  assign n33566 = ~pi0671 & n33565;
  assign n33567 = pi0671 & ~n33565;
  assign n33568 = ~n33566 & ~n33567;
  assign n33569 = ~n33562 & ~n33568;
  assign n33570 = ~n33509 & ~n33515;
  assign n33571 = ~n33502 & ~n33529;
  assign n33572 = n33568 & n33571;
  assign n33573 = n33570 & n33572;
  assign n33574 = ~n33509 & n33529;
  assign n33575 = n33515 & n33574;
  assign n33576 = ~n33502 & ~n33575;
  assign n33577 = n33509 & ~n33529;
  assign n33578 = ~n33521 & n33577;
  assign n33579 = ~n33522 & ~n33570;
  assign n33580 = n33529 & ~n33579;
  assign n33581 = n33502 & ~n33535;
  assign n33582 = ~n33580 & n33581;
  assign n33583 = ~n33578 & n33582;
  assign n33584 = ~n33576 & ~n33583;
  assign n33585 = n33509 & n33537;
  assign n33586 = ~n33529 & n33585;
  assign n33587 = ~n33584 & ~n33586;
  assign n33588 = n33568 & ~n33587;
  assign n33589 = ~n33573 & ~n33588;
  assign n33590 = ~n33569 & n33589;
  assign n33591 = ~n33542 & n33590;
  assign n33592 = ~n33502 & n33557;
  assign n33593 = n33591 & ~n33592;
  assign n33594 = pi0672 & ~n33593;
  assign n33595 = n33590 & ~n33592;
  assign n33596 = ~pi0672 & n33595;
  assign n33597 = ~n33542 & n33596;
  assign po0688 = n33594 | n33597;
  assign n33599 = pi3584 & pi9040;
  assign n33600 = pi3589 & ~pi9040;
  assign n33601 = ~n33599 & ~n33600;
  assign n33602 = pi0658 & n33601;
  assign n33603 = ~pi0658 & ~n33601;
  assign n33604 = ~n33602 & ~n33603;
  assign n33605 = pi3591 & ~pi9040;
  assign n33606 = pi3557 & pi9040;
  assign n33607 = ~n33605 & ~n33606;
  assign n33608 = ~pi0660 & ~n33607;
  assign n33609 = pi0660 & n33607;
  assign n33610 = ~n33608 & ~n33609;
  assign n33611 = ~n33604 & ~n33610;
  assign n33612 = pi3555 & pi9040;
  assign n33613 = pi3596 & ~pi9040;
  assign n33614 = ~n33612 & ~n33613;
  assign n33615 = ~pi0652 & ~n33614;
  assign n33616 = pi0652 & ~n33612;
  assign n33617 = ~n33613 & n33616;
  assign n33618 = ~n33615 & ~n33617;
  assign n33619 = pi3589 & pi9040;
  assign n33620 = pi3573 & ~pi9040;
  assign n33621 = ~n33619 & ~n33620;
  assign n33622 = ~pi0657 & ~n33621;
  assign n33623 = pi0657 & n33621;
  assign n33624 = ~n33622 & ~n33623;
  assign n33625 = pi3544 & pi9040;
  assign n33626 = pi3578 & ~pi9040;
  assign n33627 = ~n33625 & ~n33626;
  assign n33628 = ~pi0653 & ~n33627;
  assign n33629 = pi0653 & n33627;
  assign n33630 = ~n33628 & ~n33629;
  assign n33631 = n33624 & ~n33630;
  assign n33632 = ~n33618 & n33631;
  assign n33633 = pi3585 & pi9040;
  assign n33634 = pi3561 & ~pi9040;
  assign n33635 = ~n33633 & ~n33634;
  assign n33636 = ~pi0646 & ~n33635;
  assign n33637 = pi0646 & ~n33633;
  assign n33638 = ~n33634 & n33637;
  assign n33639 = ~n33636 & ~n33638;
  assign n33640 = n33630 & ~n33639;
  assign n33641 = n33624 & n33640;
  assign n33642 = n33618 & n33641;
  assign n33643 = n33630 & n33639;
  assign n33644 = ~n33618 & n33643;
  assign n33645 = ~n33642 & ~n33644;
  assign n33646 = ~n33632 & n33645;
  assign n33647 = n33611 & ~n33646;
  assign n33648 = ~n33618 & ~n33624;
  assign n33649 = ~n33639 & n33648;
  assign n33650 = ~n33630 & ~n33639;
  assign n33651 = n33624 & n33650;
  assign n33652 = n33618 & n33651;
  assign n33653 = ~n33649 & ~n33652;
  assign n33654 = ~n33624 & n33640;
  assign n33655 = n33624 & n33643;
  assign n33656 = ~n33654 & ~n33655;
  assign n33657 = n33653 & n33656;
  assign n33658 = n33604 & ~n33657;
  assign n33659 = ~n33630 & n33639;
  assign n33660 = ~n33624 & n33659;
  assign n33661 = n33618 & n33660;
  assign n33662 = ~n33658 & ~n33661;
  assign n33663 = ~n33610 & ~n33662;
  assign n33664 = ~n33647 & ~n33663;
  assign n33665 = n33604 & ~n33618;
  assign n33666 = n33624 & n33665;
  assign n33667 = n33639 & n33666;
  assign n33668 = ~n33618 & n33654;
  assign n33669 = ~n33667 & ~n33668;
  assign n33670 = ~n33624 & n33650;
  assign n33671 = ~n33643 & ~n33650;
  assign n33672 = n33618 & ~n33671;
  assign n33673 = ~n33670 & ~n33672;
  assign n33674 = ~n33604 & ~n33673;
  assign n33675 = n33624 & n33659;
  assign n33676 = ~n33632 & ~n33675;
  assign n33677 = ~n33642 & n33676;
  assign n33678 = n33604 & ~n33677;
  assign n33679 = ~n33674 & ~n33678;
  assign n33680 = ~n33604 & ~n33618;
  assign n33681 = n33640 & n33680;
  assign n33682 = n33618 & n33670;
  assign n33683 = ~n33624 & n33630;
  assign n33684 = n33639 & n33683;
  assign n33685 = n33618 & n33684;
  assign n33686 = ~n33682 & ~n33685;
  assign n33687 = n33639 & n33648;
  assign n33688 = ~n33630 & n33687;
  assign n33689 = n33686 & ~n33688;
  assign n33690 = ~n33681 & n33689;
  assign n33691 = n33679 & n33690;
  assign n33692 = n33610 & ~n33691;
  assign n33693 = n33669 & ~n33692;
  assign n33694 = n33664 & n33693;
  assign n33695 = pi0685 & ~n33694;
  assign n33696 = ~pi0685 & n33669;
  assign n33697 = n33664 & n33696;
  assign n33698 = ~n33692 & n33697;
  assign po0702 = n33695 | n33698;
  assign n33700 = pi3551 & pi9040;
  assign n33701 = pi3546 & ~pi9040;
  assign n33702 = ~n33700 & ~n33701;
  assign n33703 = ~pi0653 & ~n33702;
  assign n33704 = pi0653 & n33702;
  assign n33705 = ~n33703 & ~n33704;
  assign n33706 = pi3594 & pi9040;
  assign n33707 = pi3547 & ~pi9040;
  assign n33708 = ~n33706 & ~n33707;
  assign n33709 = pi0665 & n33708;
  assign n33710 = ~pi0665 & ~n33708;
  assign n33711 = ~n33709 & ~n33710;
  assign n33712 = pi3572 & pi9040;
  assign n33713 = pi3595 & ~pi9040;
  assign n33714 = ~n33712 & ~n33713;
  assign n33715 = ~pi0645 & n33714;
  assign n33716 = pi0645 & ~n33714;
  assign n33717 = ~n33715 & ~n33716;
  assign n33718 = ~n33711 & n33717;
  assign n33719 = pi3592 & pi9040;
  assign n33720 = pi3582 & ~pi9040;
  assign n33721 = ~n33719 & ~n33720;
  assign n33722 = ~pi0651 & ~n33721;
  assign n33723 = pi0651 & ~n33719;
  assign n33724 = ~n33720 & n33723;
  assign n33725 = ~n33722 & ~n33724;
  assign n33726 = n33718 & n33725;
  assign n33727 = pi3574 & pi9040;
  assign n33728 = pi3551 & ~pi9040;
  assign n33729 = ~n33727 & ~n33728;
  assign n33730 = ~pi0643 & n33729;
  assign n33731 = pi0643 & ~n33729;
  assign n33732 = ~n33730 & ~n33731;
  assign n33733 = pi3566 & pi9040;
  assign n33734 = pi3563 & ~pi9040;
  assign n33735 = ~n33733 & ~n33734;
  assign n33736 = ~pi0657 & ~n33735;
  assign n33737 = pi0657 & ~n33733;
  assign n33738 = ~n33734 & n33737;
  assign n33739 = ~n33736 & ~n33738;
  assign n33740 = ~n33725 & ~n33739;
  assign n33741 = ~n33732 & n33740;
  assign n33742 = n33711 & n33741;
  assign n33743 = ~n33725 & n33739;
  assign n33744 = n33732 & n33743;
  assign n33745 = n33711 & n33744;
  assign n33746 = ~n33742 & ~n33745;
  assign n33747 = n33725 & n33739;
  assign n33748 = n33732 & n33747;
  assign n33749 = ~n33711 & n33732;
  assign n33750 = ~n33739 & n33749;
  assign n33751 = ~n33725 & n33750;
  assign n33752 = ~n33748 & ~n33751;
  assign n33753 = ~n33717 & ~n33752;
  assign n33754 = n33746 & ~n33753;
  assign n33755 = ~n33726 & n33754;
  assign n33756 = n33705 & ~n33755;
  assign n33757 = n33711 & n33725;
  assign n33758 = n33732 & n33757;
  assign n33759 = ~n33739 & n33758;
  assign n33760 = n33717 & n33759;
  assign n33761 = ~n33711 & ~n33717;
  assign n33762 = n33725 & ~n33739;
  assign n33763 = n33732 & n33762;
  assign n33764 = n33761 & n33763;
  assign n33765 = ~n33711 & ~n33732;
  assign n33766 = ~n33725 & n33765;
  assign n33767 = ~n33764 & ~n33766;
  assign n33768 = ~n33732 & n33743;
  assign n33769 = ~n33748 & ~n33768;
  assign n33770 = ~n33711 & n33743;
  assign n33771 = n33769 & ~n33770;
  assign n33772 = n33717 & ~n33771;
  assign n33773 = ~n33732 & ~n33739;
  assign n33774 = n33725 & n33773;
  assign n33775 = n33711 & n33774;
  assign n33776 = n33732 & n33740;
  assign n33777 = n33711 & n33776;
  assign n33778 = ~n33775 & ~n33777;
  assign n33779 = ~n33732 & n33747;
  assign n33780 = ~n33717 & n33779;
  assign n33781 = n33778 & ~n33780;
  assign n33782 = ~n33772 & n33781;
  assign n33783 = n33767 & n33782;
  assign n33784 = ~n33705 & ~n33783;
  assign n33785 = ~n33760 & ~n33784;
  assign n33786 = ~n33756 & n33785;
  assign n33787 = n33761 & n33768;
  assign n33788 = ~n33717 & n33773;
  assign n33789 = n33711 & n33788;
  assign n33790 = ~n33787 & ~n33789;
  assign n33791 = ~n33717 & n33745;
  assign n33792 = n33790 & ~n33791;
  assign n33793 = n33786 & n33792;
  assign n33794 = ~pi0674 & ~n33793;
  assign n33795 = pi0674 & n33792;
  assign n33796 = n33785 & n33795;
  assign n33797 = ~n33756 & n33796;
  assign po0705 = n33794 | n33797;
  assign n33799 = pi3586 & pi9040;
  assign n33800 = pi3554 & ~pi9040;
  assign n33801 = ~n33799 & ~n33800;
  assign n33802 = pi0639 & n33801;
  assign n33803 = ~pi0639 & ~n33801;
  assign n33804 = ~n33802 & ~n33803;
  assign n33805 = pi3558 & pi9040;
  assign n33806 = pi3593 & ~pi9040;
  assign n33807 = ~n33805 & ~n33806;
  assign n33808 = ~pi0660 & n33807;
  assign n33809 = pi0660 & ~n33807;
  assign n33810 = ~n33808 & ~n33809;
  assign n33811 = pi3578 & pi9040;
  assign n33812 = pi3585 & ~pi9040;
  assign n33813 = ~n33811 & ~n33812;
  assign n33814 = ~pi0638 & n33813;
  assign n33815 = pi0638 & ~n33813;
  assign n33816 = ~n33814 & ~n33815;
  assign n33817 = n33810 & ~n33816;
  assign n33818 = pi3593 & pi9040;
  assign n33819 = pi3586 & ~pi9040;
  assign n33820 = ~n33818 & ~n33819;
  assign n33821 = ~pi0647 & n33820;
  assign n33822 = pi0647 & ~n33820;
  assign n33823 = ~n33821 & ~n33822;
  assign n33824 = pi3591 & pi9040;
  assign n33825 = pi3555 & ~pi9040;
  assign n33826 = ~n33824 & ~n33825;
  assign n33827 = ~pi0663 & n33826;
  assign n33828 = pi0663 & ~n33826;
  assign n33829 = ~n33827 & ~n33828;
  assign n33830 = n33823 & n33829;
  assign n33831 = n33817 & n33830;
  assign n33832 = pi3552 & pi9040;
  assign n33833 = pi3558 & ~pi9040;
  assign n33834 = ~n33832 & ~n33833;
  assign n33835 = ~pi0646 & ~n33834;
  assign n33836 = pi0646 & n33834;
  assign n33837 = ~n33835 & ~n33836;
  assign n33838 = ~n33810 & n33816;
  assign n33839 = n33837 & n33838;
  assign n33840 = n33810 & ~n33837;
  assign n33841 = n33816 & n33840;
  assign n33842 = ~n33823 & n33841;
  assign n33843 = ~n33839 & ~n33842;
  assign n33844 = ~n33810 & ~n33816;
  assign n33845 = ~n33823 & n33844;
  assign n33846 = n33843 & ~n33845;
  assign n33847 = n33829 & ~n33846;
  assign n33848 = ~n33810 & ~n33837;
  assign n33849 = n33823 & ~n33829;
  assign n33850 = n33848 & n33849;
  assign n33851 = ~n33837 & n33838;
  assign n33852 = n33823 & n33851;
  assign n33853 = ~n33850 & ~n33852;
  assign n33854 = ~n33847 & n33853;
  assign n33855 = ~n33831 & n33854;
  assign n33856 = n33817 & n33837;
  assign n33857 = n33823 & n33856;
  assign n33858 = n33837 & n33844;
  assign n33859 = ~n33823 & n33858;
  assign n33860 = ~n33857 & ~n33859;
  assign n33861 = n33855 & n33860;
  assign n33862 = ~n33804 & ~n33861;
  assign n33863 = n33823 & ~n33837;
  assign n33864 = ~n33816 & n33863;
  assign n33865 = ~n33810 & n33864;
  assign n33866 = ~n33856 & ~n33865;
  assign n33867 = n33829 & ~n33866;
  assign n33868 = n33817 & ~n33837;
  assign n33869 = ~n33823 & n33868;
  assign n33870 = n33816 & n33863;
  assign n33871 = n33810 & n33870;
  assign n33872 = ~n33869 & ~n33871;
  assign n33873 = ~n33823 & ~n33837;
  assign n33874 = ~n33810 & n33873;
  assign n33875 = n33823 & n33858;
  assign n33876 = ~n33874 & ~n33875;
  assign n33877 = ~n33829 & ~n33876;
  assign n33878 = n33872 & ~n33877;
  assign n33879 = ~n33867 & n33878;
  assign n33880 = n33804 & ~n33879;
  assign n33881 = n33810 & n33816;
  assign n33882 = n33837 & n33881;
  assign n33883 = ~n33823 & n33882;
  assign n33884 = ~n33851 & ~n33883;
  assign n33885 = ~n33869 & n33884;
  assign n33886 = ~n33829 & ~n33885;
  assign n33887 = n33810 & n33837;
  assign n33888 = n33823 & n33887;
  assign n33889 = ~n33810 & n33837;
  assign n33890 = ~n33823 & n33889;
  assign n33891 = ~n33888 & ~n33890;
  assign n33892 = n33829 & ~n33891;
  assign n33893 = ~n33886 & ~n33892;
  assign n33894 = n33816 & ~n33837;
  assign n33895 = ~n33829 & n33894;
  assign n33896 = n33823 & n33895;
  assign n33897 = n33893 & ~n33896;
  assign n33898 = ~n33880 & n33897;
  assign n33899 = ~n33862 & n33898;
  assign n33900 = ~pi0681 & ~n33899;
  assign n33901 = pi0681 & n33899;
  assign po0706 = n33900 | n33901;
  assign n33903 = n33618 & n33631;
  assign n33904 = ~n33655 & ~n33903;
  assign n33905 = ~n33668 & n33904;
  assign n33906 = n33604 & ~n33905;
  assign n33907 = ~n33618 & n33639;
  assign n33908 = n33683 & n33907;
  assign n33909 = ~n33618 & n33675;
  assign n33910 = ~n33624 & ~n33630;
  assign n33911 = ~n33640 & ~n33910;
  assign n33912 = n33618 & ~n33911;
  assign n33913 = ~n33909 & ~n33912;
  assign n33914 = ~n33908 & n33913;
  assign n33915 = ~n33604 & ~n33914;
  assign n33916 = ~n33906 & ~n33915;
  assign n33917 = n33610 & ~n33916;
  assign n33918 = n33670 & n33680;
  assign n33919 = n33624 & n33681;
  assign n33920 = ~n33918 & ~n33919;
  assign n33921 = n33604 & n33688;
  assign n33922 = n33920 & ~n33921;
  assign n33923 = ~n33630 & n33665;
  assign n33924 = ~n33618 & n33624;
  assign n33925 = n33630 & n33924;
  assign n33926 = ~n33903 & ~n33925;
  assign n33927 = ~n33604 & ~n33926;
  assign n33928 = ~n33681 & ~n33927;
  assign n33929 = ~n33618 & n33641;
  assign n33930 = ~n33685 & ~n33929;
  assign n33931 = n33604 & n33618;
  assign n33932 = n33683 & n33931;
  assign n33933 = n33604 & n33660;
  assign n33934 = ~n33932 & ~n33933;
  assign n33935 = n33930 & n33934;
  assign n33936 = n33928 & n33935;
  assign n33937 = ~n33923 & n33936;
  assign n33938 = ~n33610 & ~n33937;
  assign n33939 = n33618 & n33643;
  assign n33940 = ~n33618 & n33651;
  assign n33941 = ~n33939 & ~n33940;
  assign n33942 = n33604 & ~n33941;
  assign n33943 = ~n33938 & ~n33942;
  assign n33944 = n33922 & n33943;
  assign n33945 = ~n33917 & n33944;
  assign n33946 = ~pi0682 & ~n33945;
  assign n33947 = pi0682 & n33945;
  assign po0707 = n33946 | n33947;
  assign n33949 = ~n33711 & n33741;
  assign n33950 = ~n33711 & n33779;
  assign n33951 = ~n33744 & ~n33950;
  assign n33952 = n33711 & n33773;
  assign n33953 = ~n33711 & n33763;
  assign n33954 = ~n33952 & ~n33953;
  assign n33955 = n33951 & n33954;
  assign n33956 = n33717 & ~n33955;
  assign n33957 = n33711 & n33747;
  assign n33958 = ~n33766 & ~n33957;
  assign n33959 = ~n33776 & n33958;
  assign n33960 = ~n33717 & ~n33959;
  assign n33961 = n33711 & n33748;
  assign n33962 = ~n33960 & ~n33961;
  assign n33963 = ~n33956 & n33962;
  assign n33964 = ~n33949 & n33963;
  assign n33965 = ~n33705 & ~n33964;
  assign n33966 = n33711 & n33717;
  assign n33967 = n33779 & n33966;
  assign n33968 = n33717 & n33776;
  assign n33969 = n33717 & n33768;
  assign n33970 = ~n33968 & ~n33969;
  assign n33971 = ~n33711 & ~n33970;
  assign n33972 = ~n33967 & ~n33971;
  assign n33973 = ~n33711 & n33774;
  assign n33974 = ~n33759 & ~n33973;
  assign n33975 = n33711 & n33743;
  assign n33976 = ~n33711 & n33747;
  assign n33977 = ~n33975 & ~n33976;
  assign n33978 = ~n33774 & n33977;
  assign n33979 = ~n33744 & n33978;
  assign n33980 = ~n33717 & ~n33979;
  assign n33981 = ~n33711 & n33748;
  assign n33982 = ~n33980 & ~n33981;
  assign n33983 = n33974 & n33982;
  assign n33984 = n33972 & n33983;
  assign n33985 = n33705 & ~n33984;
  assign n33986 = n33717 & ~n33746;
  assign n33987 = ~n33985 & ~n33986;
  assign n33988 = ~n33777 & ~n33973;
  assign n33989 = ~n33717 & ~n33988;
  assign n33990 = n33987 & ~n33989;
  assign n33991 = ~n33965 & n33990;
  assign n33992 = pi0689 & ~n33991;
  assign n33993 = ~pi0689 & n33991;
  assign po0709 = n33992 | n33993;
  assign n33995 = pi3570 & pi9040;
  assign n33996 = pi3571 & ~pi9040;
  assign n33997 = ~n33995 & ~n33996;
  assign n33998 = ~pi0654 & ~n33997;
  assign n33999 = pi0654 & n33997;
  assign n34000 = ~n33998 & ~n33999;
  assign n34001 = pi3576 & pi9040;
  assign n34002 = pi3540 & ~pi9040;
  assign n34003 = ~n34001 & ~n34002;
  assign n34004 = ~pi0668 & n34003;
  assign n34005 = pi0668 & ~n34003;
  assign n34006 = ~n34004 & ~n34005;
  assign n34007 = pi3541 & pi9040;
  assign n34008 = pi3587 & ~pi9040;
  assign n34009 = ~n34007 & ~n34008;
  assign n34010 = ~pi0671 & n34009;
  assign n34011 = pi0671 & ~n34009;
  assign n34012 = ~n34010 & ~n34011;
  assign n34013 = pi3613 & pi9040;
  assign n34014 = pi3579 & ~pi9040;
  assign n34015 = ~n34013 & ~n34014;
  assign n34016 = ~pi0634 & n34015;
  assign n34017 = pi0634 & ~n34015;
  assign n34018 = ~n34016 & ~n34017;
  assign n34019 = n34012 & ~n34018;
  assign n34020 = pi3590 & pi9040;
  assign n34021 = pi3556 & ~pi9040;
  assign n34022 = ~n34020 & ~n34021;
  assign n34023 = ~pi0644 & n34022;
  assign n34024 = pi0644 & ~n34022;
  assign n34025 = ~n34023 & ~n34024;
  assign n34026 = pi3571 & pi9040;
  assign n34027 = pi3543 & ~pi9040;
  assign n34028 = ~n34026 & ~n34027;
  assign n34029 = ~pi0669 & n34028;
  assign n34030 = pi0669 & ~n34028;
  assign n34031 = ~n34029 & ~n34030;
  assign n34032 = ~n34025 & ~n34031;
  assign n34033 = n34019 & n34032;
  assign n34034 = ~n34006 & n34033;
  assign n34035 = n34025 & ~n34031;
  assign n34036 = ~n34012 & ~n34018;
  assign n34037 = n34035 & n34036;
  assign n34038 = ~n34006 & n34025;
  assign n34039 = n34018 & n34038;
  assign n34040 = n34012 & n34039;
  assign n34041 = ~n34012 & n34018;
  assign n34042 = ~n34006 & n34041;
  assign n34043 = ~n34031 & n34042;
  assign n34044 = ~n34025 & n34043;
  assign n34045 = ~n34040 & ~n34044;
  assign n34046 = ~n34037 & n34045;
  assign n34047 = ~n34034 & n34046;
  assign n34048 = n34006 & n34025;
  assign n34049 = n34036 & n34048;
  assign n34050 = n34047 & ~n34049;
  assign n34051 = ~n34000 & ~n34050;
  assign n34052 = ~n34006 & ~n34012;
  assign n34053 = ~n34018 & n34052;
  assign n34054 = ~n34025 & n34053;
  assign n34055 = ~n34039 & ~n34054;
  assign n34056 = n34006 & n34019;
  assign n34057 = ~n34025 & n34056;
  assign n34058 = n34055 & ~n34057;
  assign n34059 = n34031 & ~n34058;
  assign n34060 = n34006 & n34018;
  assign n34061 = ~n34012 & n34060;
  assign n34062 = n34031 & n34061;
  assign n34063 = ~n34025 & n34062;
  assign n34064 = n34012 & n34038;
  assign n34065 = n34012 & n34018;
  assign n34066 = n34025 & n34065;
  assign n34067 = ~n34064 & ~n34066;
  assign n34068 = n34031 & ~n34067;
  assign n34069 = ~n34063 & ~n34068;
  assign n34070 = ~n34000 & ~n34069;
  assign n34071 = ~n34059 & ~n34070;
  assign n34072 = ~n34051 & n34071;
  assign n34073 = n34006 & ~n34025;
  assign n34074 = ~n34031 & n34073;
  assign n34075 = n34065 & n34074;
  assign n34076 = n34006 & ~n34012;
  assign n34077 = n34035 & n34076;
  assign n34078 = n34031 & n34052;
  assign n34079 = n34012 & ~n34025;
  assign n34080 = n34006 & n34079;
  assign n34081 = ~n34056 & ~n34080;
  assign n34082 = ~n34078 & n34081;
  assign n34083 = n34025 & n34061;
  assign n34084 = n34082 & ~n34083;
  assign n34085 = n34006 & ~n34018;
  assign n34086 = ~n34025 & n34065;
  assign n34087 = ~n34085 & ~n34086;
  assign n34088 = ~n34031 & ~n34087;
  assign n34089 = n34019 & ~n34031;
  assign n34090 = n34025 & n34089;
  assign n34091 = ~n34088 & ~n34090;
  assign n34092 = n34084 & n34091;
  assign n34093 = n34000 & ~n34092;
  assign n34094 = ~n34077 & ~n34093;
  assign n34095 = ~n34075 & n34094;
  assign n34096 = n34072 & n34095;
  assign n34097 = pi0675 & n34096;
  assign n34098 = ~pi0675 & ~n34096;
  assign po0711 = n34097 | n34098;
  assign n34100 = ~n33871 & ~n33889;
  assign n34101 = ~n33829 & ~n34100;
  assign n34102 = ~n33823 & n33851;
  assign n34103 = ~n34101 & ~n34102;
  assign n34104 = ~n33865 & n34103;
  assign n34105 = ~n33823 & n33829;
  assign n34106 = n33868 & n34105;
  assign n34107 = ~n33857 & ~n34106;
  assign n34108 = ~n33883 & n34107;
  assign n34109 = n34104 & n34108;
  assign n34110 = n33804 & ~n34109;
  assign n34111 = ~n33816 & n33848;
  assign n34112 = ~n33823 & n34111;
  assign n34113 = ~n33842 & ~n34112;
  assign n34114 = n33823 & n33882;
  assign n34115 = ~n33852 & ~n34114;
  assign n34116 = ~n33829 & n33868;
  assign n34117 = ~n33823 & n33856;
  assign n34118 = ~n34116 & ~n34117;
  assign n34119 = ~n33816 & n33837;
  assign n34120 = ~n33810 & ~n33823;
  assign n34121 = ~n34119 & ~n34120;
  assign n34122 = ~n33894 & n34121;
  assign n34123 = n33829 & ~n34122;
  assign n34124 = n34118 & ~n34123;
  assign n34125 = n34115 & n34124;
  assign n34126 = n34113 & n34125;
  assign n34127 = ~n33804 & ~n34126;
  assign n34128 = ~n34110 & ~n34127;
  assign n34129 = pi0677 & ~n34128;
  assign n34130 = ~pi0677 & ~n34110;
  assign n34131 = ~n34127 & n34130;
  assign po0712 = n34129 | n34131;
  assign n34133 = ~n34006 & n34012;
  assign n34134 = ~n34049 & ~n34133;
  assign n34135 = ~n34079 & n34134;
  assign n34136 = ~n34031 & ~n34135;
  assign n34137 = ~n34025 & n34031;
  assign n34138 = ~n34012 & n34137;
  assign n34139 = ~n34006 & ~n34025;
  assign n34140 = ~n34018 & n34139;
  assign n34141 = n34025 & n34042;
  assign n34142 = ~n34140 & ~n34141;
  assign n34143 = n34006 & n34012;
  assign n34144 = n34025 & n34031;
  assign n34145 = n34143 & n34144;
  assign n34146 = n34142 & ~n34145;
  assign n34147 = ~n34138 & n34146;
  assign n34148 = ~n34136 & n34147;
  assign n34149 = n34000 & ~n34148;
  assign n34150 = ~n34006 & n34019;
  assign n34151 = n34025 & n34150;
  assign n34152 = ~n34006 & n34065;
  assign n34153 = ~n34025 & n34152;
  assign n34154 = ~n34151 & ~n34153;
  assign n34155 = ~n34031 & ~n34154;
  assign n34156 = ~n34149 & ~n34155;
  assign n34157 = ~n34025 & n34042;
  assign n34158 = ~n34053 & ~n34061;
  assign n34159 = ~n34031 & ~n34158;
  assign n34160 = ~n34157 & ~n34159;
  assign n34161 = ~n34057 & n34160;
  assign n34162 = ~n34000 & ~n34161;
  assign n34163 = ~n34036 & ~n34065;
  assign n34164 = n34006 & ~n34163;
  assign n34165 = ~n34066 & ~n34164;
  assign n34166 = n34031 & ~n34165;
  assign n34167 = ~n34000 & n34166;
  assign n34168 = ~n34162 & ~n34167;
  assign n34169 = n34156 & n34168;
  assign n34170 = pi0678 & ~n34169;
  assign n34171 = ~pi0678 & n34156;
  assign n34172 = n34168 & n34171;
  assign po0713 = n34170 | n34172;
  assign n34174 = pi3556 & pi9040;
  assign n34175 = pi3570 & ~pi9040;
  assign n34176 = ~n34174 & ~n34175;
  assign n34177 = ~pi0670 & n34176;
  assign n34178 = pi0670 & ~n34176;
  assign n34179 = ~n34177 & ~n34178;
  assign n34180 = pi3583 & pi9040;
  assign n34181 = pi3569 & ~pi9040;
  assign n34182 = ~n34180 & ~n34181;
  assign n34183 = ~pi0654 & ~n34182;
  assign n34184 = pi0654 & ~n34180;
  assign n34185 = ~n34181 & n34184;
  assign n34186 = ~n34183 & ~n34185;
  assign n34187 = pi3542 & pi9040;
  assign n34188 = pi3613 & ~pi9040;
  assign n34189 = ~n34187 & ~n34188;
  assign n34190 = pi0664 & n34189;
  assign n34191 = ~pi0664 & ~n34189;
  assign n34192 = ~n34190 & ~n34191;
  assign n34193 = n34186 & ~n34192;
  assign n34194 = pi3616 & pi9040;
  assign n34195 = pi3542 & ~pi9040;
  assign n34196 = ~n34194 & ~n34195;
  assign n34197 = ~pi0650 & ~n34196;
  assign n34198 = pi0650 & ~n34194;
  assign n34199 = ~n34195 & n34198;
  assign n34200 = ~n34197 & ~n34199;
  assign n34201 = pi3579 & pi9040;
  assign n34202 = pi3568 & ~pi9040;
  assign n34203 = ~n34201 & ~n34202;
  assign n34204 = ~pi0634 & n34203;
  assign n34205 = pi0634 & ~n34203;
  assign n34206 = ~n34204 & ~n34205;
  assign n34207 = n34200 & ~n34206;
  assign n34208 = n34193 & n34207;
  assign n34209 = n34200 & n34206;
  assign n34210 = ~n34186 & n34209;
  assign n34211 = ~n34208 & ~n34210;
  assign n34212 = n34179 & ~n34211;
  assign n34213 = pi3550 & pi9040;
  assign n34214 = pi3548 & ~pi9040;
  assign n34215 = ~n34213 & ~n34214;
  assign n34216 = ~pi0648 & ~n34215;
  assign n34217 = pi0648 & n34215;
  assign n34218 = ~n34216 & ~n34217;
  assign n34219 = ~n34179 & ~n34200;
  assign n34220 = n34186 & n34219;
  assign n34221 = n34193 & n34206;
  assign n34222 = n34186 & n34192;
  assign n34223 = ~n34206 & n34222;
  assign n34224 = ~n34221 & ~n34223;
  assign n34225 = ~n34186 & ~n34192;
  assign n34226 = ~n34206 & n34225;
  assign n34227 = n34200 & n34226;
  assign n34228 = n34224 & ~n34227;
  assign n34229 = ~n34179 & ~n34228;
  assign n34230 = ~n34220 & ~n34229;
  assign n34231 = ~n34186 & n34192;
  assign n34232 = n34206 & n34231;
  assign n34233 = n34200 & n34232;
  assign n34234 = n34230 & ~n34233;
  assign n34235 = ~n34200 & n34225;
  assign n34236 = ~n34186 & ~n34206;
  assign n34237 = n34192 & n34236;
  assign n34238 = ~n34235 & ~n34237;
  assign n34239 = n34179 & ~n34238;
  assign n34240 = n34206 & n34222;
  assign n34241 = ~n34200 & n34240;
  assign n34242 = ~n34239 & ~n34241;
  assign n34243 = n34234 & n34242;
  assign n34244 = n34218 & ~n34243;
  assign n34245 = ~n34212 & ~n34244;
  assign n34246 = ~n34179 & ~n34218;
  assign n34247 = ~n34238 & n34246;
  assign n34248 = n34206 & n34225;
  assign n34249 = ~n34240 & ~n34248;
  assign n34250 = n34200 & ~n34249;
  assign n34251 = ~n34208 & ~n34250;
  assign n34252 = ~n34218 & ~n34251;
  assign n34253 = ~n34247 & ~n34252;
  assign n34254 = n34179 & ~n34218;
  assign n34255 = n34193 & ~n34200;
  assign n34256 = ~n34232 & ~n34255;
  assign n34257 = n34186 & ~n34206;
  assign n34258 = n34256 & ~n34257;
  assign n34259 = n34254 & ~n34258;
  assign n34260 = n34253 & ~n34259;
  assign n34261 = n34245 & n34260;
  assign n34262 = ~pi0673 & ~n34261;
  assign n34263 = pi0673 & n34253;
  assign n34264 = n34245 & n34263;
  assign n34265 = ~n34259 & n34264;
  assign po0714 = n34262 | n34265;
  assign n34267 = n33739 & n33765;
  assign n34268 = ~n33775 & ~n34267;
  assign n34269 = ~n33725 & n33732;
  assign n34270 = ~n33779 & ~n34269;
  assign n34271 = n33732 & ~n33739;
  assign n34272 = ~n33711 & n34271;
  assign n34273 = n33711 & n33740;
  assign n34274 = ~n34272 & ~n34273;
  assign n34275 = n34270 & n34274;
  assign n34276 = ~n33717 & ~n34275;
  assign n34277 = ~n33748 & ~n33766;
  assign n34278 = n33717 & ~n34277;
  assign n34279 = ~n34276 & ~n34278;
  assign n34280 = n34268 & n34279;
  assign n34281 = n33705 & ~n34280;
  assign n34282 = ~n33711 & n33744;
  assign n34283 = n33778 & ~n34282;
  assign n34284 = ~n33717 & ~n34283;
  assign n34285 = ~n34281 & ~n34284;
  assign n34286 = n33725 & n33732;
  assign n34287 = n33717 & n34286;
  assign n34288 = n33711 & n34287;
  assign n34289 = n33761 & n33773;
  assign n34290 = n33711 & n33768;
  assign n34291 = ~n34289 & ~n34290;
  assign n34292 = ~n33725 & ~n33732;
  assign n34293 = n33711 & n34292;
  assign n34294 = ~n33763 & ~n34293;
  assign n34295 = n33717 & ~n34294;
  assign n34296 = n33717 & ~n33725;
  assign n34297 = n33732 & n34296;
  assign n34298 = ~n33711 & n34297;
  assign n34299 = ~n34295 & ~n34298;
  assign n34300 = n34291 & n34299;
  assign n34301 = ~n33705 & ~n34300;
  assign n34302 = ~n34288 & ~n34301;
  assign n34303 = ~n33950 & n34302;
  assign n34304 = n34285 & n34303;
  assign n34305 = ~pi0684 & ~n34304;
  assign n34306 = ~n33950 & ~n34281;
  assign n34307 = ~n34284 & n34306;
  assign n34308 = n34302 & n34307;
  assign n34309 = pi0684 & n34308;
  assign po0715 = n34305 | n34309;
  assign n34311 = pi3545 & ~pi9040;
  assign n34312 = pi3588 & pi9040;
  assign n34313 = ~n34311 & ~n34312;
  assign n34314 = ~pi0651 & ~n34313;
  assign n34315 = pi0651 & n34313;
  assign n34316 = ~n34314 & ~n34315;
  assign n34317 = pi3564 & pi9040;
  assign n34318 = pi3565 & ~pi9040;
  assign n34319 = ~n34317 & ~n34318;
  assign n34320 = ~pi0662 & n34319;
  assign n34321 = pi0662 & ~n34319;
  assign n34322 = ~n34320 & ~n34321;
  assign n34323 = pi3615 & pi9040;
  assign n34324 = pi3560 & ~pi9040;
  assign n34325 = ~n34323 & ~n34324;
  assign n34326 = ~pi0655 & n34325;
  assign n34327 = pi0655 & ~n34325;
  assign n34328 = ~n34326 & ~n34327;
  assign n34329 = pi3548 & pi9040;
  assign n34330 = pi3590 & ~pi9040;
  assign n34331 = ~n34329 & ~n34330;
  assign n34332 = ~pi0666 & ~n34331;
  assign n34333 = pi0666 & n34331;
  assign n34334 = ~n34332 & ~n34333;
  assign n34335 = pi3560 & pi9040;
  assign n34336 = pi3553 & ~pi9040;
  assign n34337 = ~n34335 & ~n34336;
  assign n34338 = ~pi0643 & n34337;
  assign n34339 = pi0643 & ~n34337;
  assign n34340 = ~n34338 & ~n34339;
  assign n34341 = ~n34334 & ~n34340;
  assign n34342 = ~n34328 & n34341;
  assign n34343 = ~n34322 & n34342;
  assign n34344 = pi3577 & pi9040;
  assign n34345 = pi3616 & ~pi9040;
  assign n34346 = ~n34344 & ~n34345;
  assign n34347 = ~pi0667 & ~n34346;
  assign n34348 = pi0667 & n34346;
  assign n34349 = ~n34347 & ~n34348;
  assign n34350 = n34334 & ~n34340;
  assign n34351 = ~n34322 & n34350;
  assign n34352 = n34328 & n34341;
  assign n34353 = n34322 & n34352;
  assign n34354 = ~n34351 & ~n34353;
  assign n34355 = ~n34349 & ~n34354;
  assign n34356 = ~n34343 & ~n34355;
  assign n34357 = ~n34334 & n34340;
  assign n34358 = n34328 & n34357;
  assign n34359 = n34349 & n34358;
  assign n34360 = n34341 & n34349;
  assign n34361 = ~n34322 & n34360;
  assign n34362 = ~n34359 & ~n34361;
  assign n34363 = n34356 & n34362;
  assign n34364 = n34334 & n34340;
  assign n34365 = ~n34328 & n34364;
  assign n34366 = ~n34322 & n34365;
  assign n34367 = ~n34328 & n34357;
  assign n34368 = n34322 & n34367;
  assign n34369 = ~n34366 & ~n34368;
  assign n34370 = n34363 & n34369;
  assign n34371 = n34316 & ~n34370;
  assign n34372 = ~n34316 & ~n34349;
  assign n34373 = ~n34322 & n34328;
  assign n34374 = ~n34334 & n34373;
  assign n34375 = n34328 & n34340;
  assign n34376 = ~n34374 & ~n34375;
  assign n34377 = n34372 & ~n34376;
  assign n34378 = n34322 & ~n34328;
  assign n34379 = ~n34340 & n34378;
  assign n34380 = ~n34334 & n34379;
  assign n34381 = n34322 & n34334;
  assign n34382 = n34328 & n34381;
  assign n34383 = ~n34380 & ~n34382;
  assign n34384 = ~n34322 & n34349;
  assign n34385 = ~n34328 & n34384;
  assign n34386 = ~n34341 & n34385;
  assign n34387 = n34349 & n34365;
  assign n34388 = ~n34386 & ~n34387;
  assign n34389 = n34383 & n34388;
  assign n34390 = ~n34316 & ~n34389;
  assign n34391 = n34328 & n34364;
  assign n34392 = n34322 & ~n34349;
  assign n34393 = n34391 & n34392;
  assign n34394 = ~n34328 & n34350;
  assign n34395 = n34322 & n34394;
  assign n34396 = ~n34368 & ~n34395;
  assign n34397 = ~n34349 & ~n34396;
  assign n34398 = ~n34393 & ~n34397;
  assign n34399 = n34349 & n34380;
  assign n34400 = n34398 & ~n34399;
  assign n34401 = ~n34390 & n34400;
  assign n34402 = ~n34377 & n34401;
  assign n34403 = ~n34371 & n34402;
  assign n34404 = n34328 & n34350;
  assign n34405 = n34322 & n34349;
  assign n34406 = n34404 & n34405;
  assign n34407 = n34403 & ~n34406;
  assign n34408 = ~pi0690 & ~n34407;
  assign n34409 = pi0690 & ~n34406;
  assign n34410 = n34402 & n34409;
  assign n34411 = ~n34371 & n34410;
  assign po0716 = n34408 | n34411;
  assign n34413 = ~n33670 & ~n33675;
  assign n34414 = ~n33604 & ~n34413;
  assign n34415 = n33618 & n33655;
  assign n34416 = ~n34414 & ~n34415;
  assign n34417 = n33618 & n33630;
  assign n34418 = ~n33683 & ~n34417;
  assign n34419 = ~n33651 & n34418;
  assign n34420 = n33604 & ~n34419;
  assign n34421 = n34416 & ~n34420;
  assign n34422 = ~n33610 & ~n34421;
  assign n34423 = ~n33618 & n33684;
  assign n34424 = ~n33604 & n34423;
  assign n34425 = ~n33919 & ~n34424;
  assign n34426 = ~n33921 & n34425;
  assign n34427 = n33604 & n33630;
  assign n34428 = n33924 & n34427;
  assign n34429 = n33618 & n33675;
  assign n34430 = ~n33604 & n33683;
  assign n34431 = ~n34429 & ~n34430;
  assign n34432 = ~n33682 & n34431;
  assign n34433 = ~n34428 & n34432;
  assign n34434 = ~n33639 & n33924;
  assign n34435 = ~n33688 & ~n34434;
  assign n34436 = n34433 & n34435;
  assign n34437 = ~n33933 & n34436;
  assign n34438 = n33610 & ~n34437;
  assign n34439 = n34426 & ~n34438;
  assign n34440 = ~n34422 & n34439;
  assign n34441 = ~pi0692 & ~n34440;
  assign n34442 = pi0692 & n34426;
  assign n34443 = ~n34422 & n34442;
  assign n34444 = ~n34438 & n34443;
  assign po0717 = n34441 | n34444;
  assign n34446 = n33823 & n33844;
  assign n34447 = ~n34114 & ~n34446;
  assign n34448 = ~n33829 & n34447;
  assign n34449 = n33804 & ~n34448;
  assign n34450 = ~n33817 & ~n33838;
  assign n34451 = n33837 & ~n34450;
  assign n34452 = n33810 & n33863;
  assign n34453 = ~n33823 & n33838;
  assign n34454 = ~n34452 & ~n34453;
  assign n34455 = ~n33823 & n33887;
  assign n34456 = n34454 & ~n34455;
  assign n34457 = ~n34451 & n34456;
  assign n34458 = n33829 & n34457;
  assign n34459 = n34449 & ~n34458;
  assign n34460 = ~n33823 & n34451;
  assign n34461 = ~n34112 & ~n34460;
  assign n34462 = n33804 & ~n34461;
  assign n34463 = ~n34459 & ~n34462;
  assign n34464 = ~n33829 & ~n34450;
  assign n34465 = n33823 & n34464;
  assign n34466 = ~n33823 & n33881;
  assign n34467 = ~n33859 & ~n34466;
  assign n34468 = ~n33829 & ~n34467;
  assign n34469 = ~n33837 & n34464;
  assign n34470 = ~n34468 & ~n34469;
  assign n34471 = ~n34465 & n34470;
  assign n34472 = ~n33804 & ~n34471;
  assign n34473 = n34463 & ~n34472;
  assign n34474 = n33829 & ~n34447;
  assign n34475 = ~n33842 & ~n34474;
  assign n34476 = ~n33804 & ~n34475;
  assign n34477 = ~n33829 & n33842;
  assign n34478 = n33829 & ~n34461;
  assign n34479 = ~n34477 & ~n34478;
  assign n34480 = ~n34476 & n34479;
  assign n34481 = n34473 & n34480;
  assign n34482 = pi0700 & ~n34481;
  assign n34483 = ~pi0700 & n34480;
  assign n34484 = ~n34472 & n34483;
  assign n34485 = n34463 & n34484;
  assign po0718 = n34482 | n34485;
  assign n34487 = n33529 & n33559;
  assign n34488 = ~n33515 & ~n33529;
  assign n34489 = ~n33509 & n34488;
  assign n34490 = ~n33556 & ~n34489;
  assign n34491 = n33502 & ~n34490;
  assign n34492 = ~n34487 & ~n34491;
  assign n34493 = ~n33502 & n33529;
  assign n34494 = ~n33515 & n34493;
  assign n34495 = n33521 & n34494;
  assign n34496 = n33537 & n33571;
  assign n34497 = ~n34495 & ~n34496;
  assign n34498 = ~n33502 & n33509;
  assign n34499 = n33531 & n34498;
  assign n34500 = n34497 & ~n34499;
  assign n34501 = ~n33533 & ~n33545;
  assign n34502 = n33515 & n33577;
  assign n34503 = n34501 & ~n34502;
  assign n34504 = n34500 & n34503;
  assign n34505 = n34492 & n34504;
  assign n34506 = ~n33568 & ~n34505;
  assign n34507 = ~n33532 & ~n33556;
  assign n34508 = ~n33529 & ~n34507;
  assign n34509 = n33521 & n33529;
  assign n34510 = ~n33509 & n34509;
  assign n34511 = ~n33585 & ~n34510;
  assign n34512 = n33509 & ~n33515;
  assign n34513 = ~n33529 & n34512;
  assign n34514 = n34511 & ~n34513;
  assign n34515 = n33502 & ~n34514;
  assign n34516 = n33529 & n33555;
  assign n34517 = n33521 & n33544;
  assign n34518 = ~n34516 & ~n34517;
  assign n34519 = ~n33502 & ~n34518;
  assign n34520 = n33529 & n33538;
  assign n34521 = ~n34519 & ~n34520;
  assign n34522 = ~n34515 & n34521;
  assign n34523 = ~n34508 & n34522;
  assign n34524 = n33568 & ~n34523;
  assign n34525 = n33502 & n33575;
  assign n34526 = ~n34524 & ~n34525;
  assign n34527 = n33550 & n34493;
  assign n34528 = ~n33515 & n34527;
  assign n34529 = n34526 & ~n34528;
  assign n34530 = ~n34506 & n34529;
  assign n34531 = ~pi0697 & ~n34530;
  assign n34532 = pi0697 & n34526;
  assign n34533 = ~n34506 & n34532;
  assign n34534 = ~n34528 & n34533;
  assign po0720 = n34531 | n34534;
  assign n34536 = n34192 & n34207;
  assign n34537 = ~n34186 & n34536;
  assign n34538 = ~n34193 & ~n34257;
  assign n34539 = n34200 & ~n34538;
  assign n34540 = ~n34232 & ~n34539;
  assign n34541 = n34179 & ~n34540;
  assign n34542 = n34192 & ~n34200;
  assign n34543 = n34179 & n34542;
  assign n34544 = n34206 & n34543;
  assign n34545 = ~n34192 & ~n34206;
  assign n34546 = ~n34232 & ~n34545;
  assign n34547 = ~n34200 & ~n34546;
  assign n34548 = ~n34179 & n34200;
  assign n34549 = n34222 & n34548;
  assign n34550 = n34206 & n34549;
  assign n34551 = ~n34547 & ~n34550;
  assign n34552 = ~n34544 & n34551;
  assign n34553 = ~n34541 & n34552;
  assign n34554 = ~n34537 & n34553;
  assign n34555 = ~n34218 & ~n34554;
  assign n34556 = n34179 & n34200;
  assign n34557 = ~n34225 & ~n34240;
  assign n34558 = n34556 & ~n34557;
  assign n34559 = n34179 & n34206;
  assign n34560 = n34225 & n34559;
  assign n34561 = ~n34558 & ~n34560;
  assign n34562 = n34218 & ~n34561;
  assign n34563 = ~n34200 & n34257;
  assign n34564 = n34200 & n34248;
  assign n34565 = ~n34563 & ~n34564;
  assign n34566 = ~n34179 & ~n34565;
  assign n34567 = ~n34562 & ~n34566;
  assign n34568 = ~n34200 & ~n34206;
  assign n34569 = n34192 & n34568;
  assign n34570 = n34186 & n34569;
  assign n34571 = ~n34257 & ~n34568;
  assign n34572 = ~n34179 & ~n34571;
  assign n34573 = ~n34200 & n34206;
  assign n34574 = ~n34192 & n34573;
  assign n34575 = n34186 & n34574;
  assign n34576 = ~n34572 & ~n34575;
  assign n34577 = ~n34570 & n34576;
  assign n34578 = n34218 & ~n34577;
  assign n34579 = ~n34200 & n34232;
  assign n34580 = ~n34537 & ~n34579;
  assign n34581 = n34179 & ~n34580;
  assign n34582 = ~n34578 & ~n34581;
  assign n34583 = n34567 & n34582;
  assign n34584 = ~n34555 & n34583;
  assign n34585 = pi0679 & n34584;
  assign n34586 = ~pi0679 & ~n34584;
  assign po0721 = n34585 | n34586;
  assign n34588 = ~n33618 & ~n33630;
  assign n34589 = ~n34434 & ~n34588;
  assign n34590 = ~n33604 & ~n34589;
  assign n34591 = n33618 & n33624;
  assign n34592 = n33639 & n34591;
  assign n34593 = ~n34590 & ~n34592;
  assign n34594 = n33604 & n33643;
  assign n34595 = ~n33618 & n34594;
  assign n34596 = ~n33940 & ~n34595;
  assign n34597 = n34593 & n34596;
  assign n34598 = n33610 & ~n34597;
  assign n34599 = ~n33641 & ~n33685;
  assign n34600 = ~n33618 & n33659;
  assign n34601 = n34599 & ~n34600;
  assign n34602 = n33604 & ~n34601;
  assign n34603 = n33643 & n33680;
  assign n34604 = ~n33668 & ~n34603;
  assign n34605 = ~n34602 & n34604;
  assign n34606 = ~n33651 & ~n33661;
  assign n34607 = ~n33604 & ~n34606;
  assign n34608 = n34605 & ~n34607;
  assign n34609 = ~n33610 & ~n34608;
  assign n34610 = ~n34598 & ~n34609;
  assign n34611 = ~n33618 & n33650;
  assign n34612 = n33618 & ~n33656;
  assign n34613 = ~n34611 & ~n34612;
  assign n34614 = ~n33604 & ~n34613;
  assign n34615 = ~n33641 & n34413;
  assign n34616 = n33931 & ~n34615;
  assign n34617 = ~n34614 & ~n34616;
  assign n34618 = n34610 & n34617;
  assign n34619 = ~pi0686 & ~n34618;
  assign n34620 = ~n34609 & n34617;
  assign n34621 = pi0686 & n34620;
  assign n34622 = ~n34598 & n34621;
  assign po0722 = n34619 | n34622;
  assign n34624 = n34025 & n34056;
  assign n34625 = ~n34141 & ~n34624;
  assign n34626 = n34031 & ~n34625;
  assign n34627 = n34053 & n34137;
  assign n34628 = ~n34626 & ~n34627;
  assign n34629 = ~n34077 & n34628;
  assign n34630 = ~n34012 & ~n34025;
  assign n34631 = n34006 & n34630;
  assign n34632 = n34018 & n34631;
  assign n34633 = ~n34152 & ~n34632;
  assign n34634 = ~n34056 & n34633;
  assign n34635 = n34031 & ~n34634;
  assign n34636 = n34000 & n34635;
  assign n34637 = ~n34006 & n34018;
  assign n34638 = ~n34031 & n34637;
  assign n34639 = n34012 & n34638;
  assign n34640 = n34025 & n34639;
  assign n34641 = ~n34031 & n34150;
  assign n34642 = ~n34049 & ~n34075;
  assign n34643 = ~n34044 & n34642;
  assign n34644 = ~n34641 & n34643;
  assign n34645 = n34000 & ~n34644;
  assign n34646 = ~n34025 & n34089;
  assign n34647 = ~n34639 & ~n34646;
  assign n34648 = ~n34140 & n34647;
  assign n34649 = n34018 & n34048;
  assign n34650 = ~n34025 & n34036;
  assign n34651 = ~n34052 & ~n34650;
  assign n34652 = n34031 & ~n34651;
  assign n34653 = ~n34649 & ~n34652;
  assign n34654 = n34648 & n34653;
  assign n34655 = ~n34000 & ~n34654;
  assign n34656 = ~n34645 & ~n34655;
  assign n34657 = ~n34640 & n34656;
  assign n34658 = ~n34636 & n34657;
  assign n34659 = n34629 & n34658;
  assign n34660 = pi0688 & ~n34659;
  assign n34661 = ~pi0688 & n34629;
  assign n34662 = n34658 & n34661;
  assign po0723 = n34660 | n34662;
  assign n34664 = ~n33530 & ~n33536;
  assign n34665 = ~n33502 & ~n34664;
  assign n34666 = ~n33592 & ~n34665;
  assign n34667 = ~n33509 & ~n33521;
  assign n34668 = n33502 & n34667;
  assign n34669 = ~n33529 & n34668;
  assign n34670 = ~n33502 & n33522;
  assign n34671 = ~n33529 & n34670;
  assign n34672 = ~n34499 & ~n34671;
  assign n34673 = n33509 & n33529;
  assign n34674 = n33521 & n34673;
  assign n34675 = ~n33529 & n33555;
  assign n34676 = ~n34674 & ~n34675;
  assign n34677 = ~n34667 & n34676;
  assign n34678 = n33502 & ~n34677;
  assign n34679 = ~n33539 & ~n34678;
  assign n34680 = n34672 & n34679;
  assign n34681 = ~n33568 & ~n34680;
  assign n34682 = ~n34669 & ~n34681;
  assign n34683 = ~n33556 & ~n33575;
  assign n34684 = ~n33585 & n34683;
  assign n34685 = ~n33502 & ~n34684;
  assign n34686 = n33529 & n33535;
  assign n34687 = ~n33559 & ~n34686;
  assign n34688 = n33502 & ~n34687;
  assign n34689 = ~n34510 & ~n34688;
  assign n34690 = ~n34685 & n34689;
  assign n34691 = ~n33545 & ~n33586;
  assign n34692 = n34690 & n34691;
  assign n34693 = n33568 & ~n34692;
  assign n34694 = n34682 & ~n34693;
  assign n34695 = n34666 & n34694;
  assign n34696 = ~pi0698 & ~n34695;
  assign n34697 = pi0698 & n34682;
  assign n34698 = n34666 & n34697;
  assign n34699 = ~n34693 & n34698;
  assign po0724 = n34696 | n34699;
  assign n34701 = ~n33751 & ~n33973;
  assign n34702 = ~n33961 & n34701;
  assign n34703 = n33717 & ~n34702;
  assign n34704 = ~n33764 & ~n33791;
  assign n34705 = ~n33759 & ~n33969;
  assign n34706 = ~n33741 & ~n33976;
  assign n34707 = ~n33717 & ~n34706;
  assign n34708 = ~n33950 & ~n34707;
  assign n34709 = n34705 & n34708;
  assign n34710 = n33705 & ~n34709;
  assign n34711 = n33732 & n33739;
  assign n34712 = ~n34269 & ~n34711;
  assign n34713 = n33711 & ~n34712;
  assign n34714 = ~n33770 & ~n33774;
  assign n34715 = ~n33717 & ~n34714;
  assign n34716 = n33711 & n33739;
  assign n34717 = ~n33748 & ~n34716;
  assign n34718 = ~n33740 & n34717;
  assign n34719 = n33717 & ~n34718;
  assign n34720 = ~n34715 & ~n34719;
  assign n34721 = ~n34713 & n34720;
  assign n34722 = ~n33705 & ~n34721;
  assign n34723 = ~n34710 & ~n34722;
  assign n34724 = n34704 & n34723;
  assign n34725 = ~n34703 & n34724;
  assign n34726 = ~pi0693 & ~n34725;
  assign n34727 = pi0693 & n34704;
  assign n34728 = ~n34703 & n34727;
  assign n34729 = n34723 & n34728;
  assign po0725 = n34726 | n34729;
  assign n34731 = n34322 & n34358;
  assign n34732 = ~n34322 & n34391;
  assign n34733 = ~n34731 & ~n34732;
  assign n34734 = n34349 & ~n34733;
  assign n34735 = ~n34380 & ~n34387;
  assign n34736 = ~n34334 & n34378;
  assign n34737 = ~n34382 & ~n34736;
  assign n34738 = ~n34349 & ~n34737;
  assign n34739 = ~n34322 & ~n34349;
  assign n34740 = n34357 & n34739;
  assign n34741 = n34328 & n34740;
  assign n34742 = ~n34322 & ~n34328;
  assign n34743 = ~n34340 & n34742;
  assign n34744 = n34334 & n34743;
  assign n34745 = n34349 & n34352;
  assign n34746 = ~n34744 & ~n34745;
  assign n34747 = ~n34741 & n34746;
  assign n34748 = ~n34738 & n34747;
  assign n34749 = n34735 & n34748;
  assign n34750 = n34316 & ~n34749;
  assign n34751 = ~n34349 & n34380;
  assign n34752 = n34364 & n34405;
  assign n34753 = ~n34328 & n34752;
  assign n34754 = ~n34751 & ~n34753;
  assign n34755 = ~n34750 & n34754;
  assign n34756 = ~n34734 & n34755;
  assign n34757 = ~n34328 & ~n34334;
  assign n34758 = n34384 & n34757;
  assign n34759 = ~n34359 & ~n34758;
  assign n34760 = n34349 & n34394;
  assign n34761 = n34322 & n34404;
  assign n34762 = ~n34760 & ~n34761;
  assign n34763 = ~n34322 & n34367;
  assign n34764 = ~n34731 & ~n34763;
  assign n34765 = ~n34322 & n34364;
  assign n34766 = n34328 & ~n34340;
  assign n34767 = ~n34765 & ~n34766;
  assign n34768 = ~n34349 & ~n34767;
  assign n34769 = n34764 & ~n34768;
  assign n34770 = n34762 & n34769;
  assign n34771 = n34759 & n34770;
  assign n34772 = ~n34316 & ~n34771;
  assign n34773 = n34756 & ~n34772;
  assign n34774 = ~pi0676 & ~n34773;
  assign n34775 = pi0676 & n34756;
  assign n34776 = ~n34772 & n34775;
  assign po0726 = n34774 | n34776;
  assign n34778 = ~n34753 & ~n34758;
  assign n34779 = ~n34380 & ~n34391;
  assign n34780 = ~n34765 & n34779;
  assign n34781 = ~n34349 & ~n34780;
  assign n34782 = ~n34340 & n34373;
  assign n34783 = ~n34334 & n34782;
  assign n34784 = ~n34744 & ~n34783;
  assign n34785 = ~n34406 & n34784;
  assign n34786 = n34349 & n34367;
  assign n34787 = n34785 & ~n34786;
  assign n34788 = ~n34781 & n34787;
  assign n34789 = n34316 & ~n34788;
  assign n34790 = n34322 & n34360;
  assign n34791 = n34334 & n34373;
  assign n34792 = ~n34391 & ~n34791;
  assign n34793 = n34349 & ~n34792;
  assign n34794 = ~n34790 & ~n34793;
  assign n34795 = n34350 & n34392;
  assign n34796 = ~n34349 & n34358;
  assign n34797 = ~n34795 & ~n34796;
  assign n34798 = n34794 & n34797;
  assign n34799 = n34334 & n34378;
  assign n34800 = ~n34731 & ~n34799;
  assign n34801 = ~n34763 & n34800;
  assign n34802 = n34798 & n34801;
  assign n34803 = ~n34316 & ~n34802;
  assign n34804 = ~n34731 & n34784;
  assign n34805 = ~n34349 & ~n34804;
  assign n34806 = ~n34803 & ~n34805;
  assign n34807 = ~n34789 & n34806;
  assign n34808 = n34778 & n34807;
  assign n34809 = pi0683 & ~n34808;
  assign n34810 = ~pi0683 & n34808;
  assign po0727 = n34809 | n34810;
  assign n34812 = ~n33509 & n33521;
  assign n34813 = ~n33502 & n34812;
  assign n34814 = ~n33529 & n34813;
  assign n34815 = n33529 & n34512;
  assign n34816 = ~n33536 & ~n34815;
  assign n34817 = ~n34517 & n34816;
  assign n34818 = ~n34814 & n34817;
  assign n34819 = n33502 & n33532;
  assign n34820 = n34818 & ~n34819;
  assign n34821 = n33568 & ~n34820;
  assign n34822 = ~n33586 & ~n34520;
  assign n34823 = n33502 & ~n34822;
  assign n34824 = ~n33568 & n33570;
  assign n34825 = ~n33502 & n34824;
  assign n34826 = ~n33521 & n34673;
  assign n34827 = ~n34512 & ~n34826;
  assign n34828 = ~n33538 & n34827;
  assign n34829 = n33502 & ~n34828;
  assign n34830 = ~n33509 & n33555;
  assign n34831 = n33529 & n34830;
  assign n34832 = ~n34829 & ~n34831;
  assign n34833 = ~n33568 & ~n34832;
  assign n34834 = ~n34825 & ~n34833;
  assign n34835 = ~n34823 & n34834;
  assign n34836 = ~n33533 & ~n33536;
  assign n34837 = n33529 & n33585;
  assign n34838 = ~n34489 & ~n34837;
  assign n34839 = n34836 & n34838;
  assign n34840 = ~n33502 & ~n34839;
  assign n34841 = n34835 & ~n34840;
  assign n34842 = ~n34821 & n34841;
  assign n34843 = ~pi0695 & ~n34842;
  assign n34844 = pi0695 & n34835;
  assign n34845 = ~n34821 & n34844;
  assign n34846 = ~n34840 & n34845;
  assign po0728 = n34843 | n34846;
  assign n34848 = ~n33829 & n33869;
  assign n34849 = n33863 & ~n34450;
  assign n34850 = ~n33882 & ~n34849;
  assign n34851 = ~n34112 & n34850;
  assign n34852 = n33829 & ~n34851;
  assign n34853 = ~n33823 & n33839;
  assign n34854 = ~n34852 & ~n34853;
  assign n34855 = ~n33837 & n33881;
  assign n34856 = n33823 & n34119;
  assign n34857 = ~n34855 & ~n34856;
  assign n34858 = ~n34453 & n34857;
  assign n34859 = ~n33829 & ~n34858;
  assign n34860 = n34854 & ~n34859;
  assign n34861 = n33804 & ~n34860;
  assign n34862 = ~n34848 & ~n34861;
  assign n34863 = n33823 & n33838;
  assign n34864 = ~n33837 & n33844;
  assign n34865 = ~n34863 & ~n34864;
  assign n34866 = ~n33829 & ~n34865;
  assign n34867 = ~n33883 & ~n34866;
  assign n34868 = ~n33859 & ~n33869;
  assign n34869 = ~n33823 & n33894;
  assign n34870 = ~n34119 & ~n34869;
  assign n34871 = ~n34855 & n34870;
  assign n34872 = n33829 & ~n34871;
  assign n34873 = n33823 & n33839;
  assign n34874 = ~n34872 & ~n34873;
  assign n34875 = n34868 & n34874;
  assign n34876 = n34867 & n34875;
  assign n34877 = ~n33804 & ~n34876;
  assign n34878 = ~n33875 & ~n34455;
  assign n34879 = n33829 & ~n34878;
  assign n34880 = ~n34877 & ~n34879;
  assign n34881 = n34862 & n34880;
  assign n34882 = pi0699 & n34881;
  assign n34883 = ~pi0699 & ~n34881;
  assign po0729 = n34882 | n34883;
  assign n34885 = pi3543 & pi9040;
  assign n34886 = pi3541 & ~pi9040;
  assign n34887 = ~n34885 & ~n34886;
  assign n34888 = pi0664 & n34887;
  assign n34889 = ~pi0664 & ~n34887;
  assign n34890 = ~n34888 & ~n34889;
  assign n34891 = pi3545 & pi9040;
  assign n34892 = pi3583 & ~pi9040;
  assign n34893 = ~n34891 & ~n34892;
  assign n34894 = pi0655 & n34893;
  assign n34895 = ~pi0655 & ~n34893;
  assign n34896 = ~n34894 & ~n34895;
  assign n34897 = pi3568 & pi9040;
  assign n34898 = pi3575 & ~pi9040;
  assign n34899 = ~n34897 & ~n34898;
  assign n34900 = ~pi0648 & n34899;
  assign n34901 = pi0648 & ~n34899;
  assign n34902 = ~n34900 & ~n34901;
  assign n34903 = ~n34896 & ~n34902;
  assign n34904 = ~n34890 & n34903;
  assign n34905 = n34896 & ~n34902;
  assign n34906 = n34890 & n34905;
  assign n34907 = ~n34904 & ~n34906;
  assign n34908 = pi3540 & pi9040;
  assign n34909 = pi3615 & ~pi9040;
  assign n34910 = ~n34908 & ~n34909;
  assign n34911 = pi0656 & n34910;
  assign n34912 = ~pi0656 & ~n34910;
  assign n34913 = ~n34911 & ~n34912;
  assign n34914 = n34890 & ~n34913;
  assign n34915 = n34896 & n34914;
  assign n34916 = n34907 & ~n34915;
  assign n34917 = pi3549 & pi9040;
  assign n34918 = pi3564 & ~pi9040;
  assign n34919 = ~n34917 & ~n34918;
  assign n34920 = ~pi0636 & n34919;
  assign n34921 = pi0636 & ~n34919;
  assign n34922 = ~n34920 & ~n34921;
  assign n34923 = pi3569 & pi9040;
  assign n34924 = pi3550 & ~pi9040;
  assign n34925 = ~n34923 & ~n34924;
  assign n34926 = ~pi0666 & n34925;
  assign n34927 = pi0666 & ~n34925;
  assign n34928 = ~n34926 & ~n34927;
  assign n34929 = n34922 & ~n34928;
  assign n34930 = ~n34916 & n34929;
  assign n34931 = ~n34896 & n34902;
  assign n34932 = n34890 & n34931;
  assign n34933 = ~n34928 & n34932;
  assign n34934 = n34913 & n34933;
  assign n34935 = n34890 & n34903;
  assign n34936 = ~n34922 & n34935;
  assign n34937 = ~n34890 & n34896;
  assign n34938 = n34896 & n34902;
  assign n34939 = n34913 & n34938;
  assign n34940 = ~n34937 & ~n34939;
  assign n34941 = ~n34922 & ~n34940;
  assign n34942 = ~n34936 & ~n34941;
  assign n34943 = ~n34928 & ~n34942;
  assign n34944 = ~n34934 & ~n34943;
  assign n34945 = ~n34890 & n34913;
  assign n34946 = n34896 & n34945;
  assign n34947 = ~n34890 & ~n34913;
  assign n34948 = ~n34896 & n34947;
  assign n34949 = n34902 & n34948;
  assign n34950 = ~n34946 & ~n34949;
  assign n34951 = ~n34922 & ~n34950;
  assign n34952 = n34944 & ~n34951;
  assign n34953 = n34913 & n34922;
  assign n34954 = n34938 & n34953;
  assign n34955 = n34890 & n34954;
  assign n34956 = ~n34905 & ~n34931;
  assign n34957 = n34914 & ~n34956;
  assign n34958 = n34904 & ~n34913;
  assign n34959 = ~n34957 & ~n34958;
  assign n34960 = ~n34890 & n34938;
  assign n34961 = n34922 & n34960;
  assign n34962 = ~n34913 & n34961;
  assign n34963 = n34945 & ~n34956;
  assign n34964 = n34913 & n34935;
  assign n34965 = ~n34963 & ~n34964;
  assign n34966 = ~n34962 & n34965;
  assign n34967 = n34959 & n34966;
  assign n34968 = ~n34955 & n34967;
  assign n34969 = ~n34913 & ~n34922;
  assign n34970 = n34890 & n34969;
  assign n34971 = n34902 & n34970;
  assign n34972 = n34968 & ~n34971;
  assign n34973 = n34928 & ~n34972;
  assign n34974 = n34952 & ~n34973;
  assign n34975 = ~n34930 & n34974;
  assign n34976 = ~pi0714 & ~n34975;
  assign n34977 = pi0714 & n34952;
  assign n34978 = ~n34930 & n34977;
  assign n34979 = ~n34973 & n34978;
  assign po0730 = n34976 | n34979;
  assign n34981 = n34890 & n34938;
  assign n34982 = ~n34922 & n34981;
  assign n34983 = ~n34913 & n34982;
  assign n34984 = n34903 & n34969;
  assign n34985 = ~n34890 & n34984;
  assign n34986 = ~n34983 & ~n34985;
  assign n34987 = ~n34958 & ~n34962;
  assign n34988 = ~n34902 & n34913;
  assign n34989 = n34890 & n34988;
  assign n34990 = ~n34939 & ~n34989;
  assign n34991 = ~n34922 & ~n34990;
  assign n34992 = n34922 & ~n34947;
  assign n34993 = ~n34956 & n34992;
  assign n34994 = ~n34890 & ~n34938;
  assign n34995 = ~n34922 & n34994;
  assign n34996 = ~n34913 & n34995;
  assign n34997 = ~n34993 & ~n34996;
  assign n34998 = ~n34991 & n34997;
  assign n34999 = n34987 & n34998;
  assign n35000 = ~n34928 & ~n34999;
  assign n35001 = n34986 & ~n35000;
  assign n35002 = n34906 & n34922;
  assign n35003 = n34913 & n35002;
  assign n35004 = n34922 & n34928;
  assign n35005 = n34947 & ~n34956;
  assign n35006 = ~n34939 & ~n35005;
  assign n35007 = ~n34935 & n35006;
  assign n35008 = n35004 & ~n35007;
  assign n35009 = n34904 & n34913;
  assign n35010 = ~n34890 & n34988;
  assign n35011 = n34913 & n34931;
  assign n35012 = ~n35010 & ~n35011;
  assign n35013 = ~n34913 & n34938;
  assign n35014 = ~n34932 & ~n35013;
  assign n35015 = n35012 & n35014;
  assign n35016 = ~n34922 & ~n35015;
  assign n35017 = ~n35009 & ~n35016;
  assign n35018 = n34928 & ~n35017;
  assign n35019 = ~n35008 & ~n35018;
  assign n35020 = ~n35003 & n35019;
  assign n35021 = n35001 & n35020;
  assign n35022 = pi0702 & ~n35021;
  assign n35023 = ~pi0702 & n35001;
  assign n35024 = n35020 & n35023;
  assign po0731 = n35022 | n35024;
  assign n35026 = ~n34025 & ~n34163;
  assign n35027 = n34006 & n35026;
  assign n35028 = n34018 & n34139;
  assign n35029 = ~n34085 & ~n35028;
  assign n35030 = ~n34152 & n35029;
  assign n35031 = ~n34031 & ~n35030;
  assign n35032 = ~n34060 & ~n34150;
  assign n35033 = n34031 & ~n35032;
  assign n35034 = ~n35031 & ~n35033;
  assign n35035 = ~n35027 & n35034;
  assign n35036 = n34025 & n34053;
  assign n35037 = n35035 & ~n35036;
  assign n35038 = ~n34000 & ~n35037;
  assign n35039 = n34035 & ~n35032;
  assign n35040 = ~n34056 & ~n34061;
  assign n35041 = ~n34053 & ~n34152;
  assign n35042 = n35040 & n35041;
  assign n35043 = ~n34025 & ~n35042;
  assign n35044 = ~n35039 & ~n35043;
  assign n35045 = ~n34141 & n35044;
  assign n35046 = n34000 & ~n35045;
  assign n35047 = ~n35038 & ~n35046;
  assign n35048 = ~n34025 & n34150;
  assign n35049 = ~n35036 & ~n35048;
  assign n35050 = n34031 & ~n35049;
  assign n35051 = n35047 & ~n35050;
  assign n35052 = pi0680 & ~n35051;
  assign n35053 = ~pi0680 & ~n35050;
  assign n35054 = ~n35046 & n35053;
  assign n35055 = ~n35038 & n35054;
  assign po0732 = n35052 | n35055;
  assign n35057 = n34179 & n34237;
  assign n35058 = ~n34200 & n34222;
  assign n35059 = ~n34221 & ~n35058;
  assign n35060 = n34179 & ~n35059;
  assign n35061 = ~n34179 & ~n34546;
  assign n35062 = ~n35060 & ~n35061;
  assign n35063 = ~n34564 & n35062;
  assign n35064 = n34218 & ~n35063;
  assign n35065 = ~n35057 & ~n35064;
  assign n35066 = ~n34206 & n34556;
  assign n35067 = ~n34573 & ~n35066;
  assign n35068 = ~n34186 & ~n35067;
  assign n35069 = ~n34208 & ~n35068;
  assign n35070 = ~n34574 & n35069;
  assign n35071 = n34200 & n34240;
  assign n35072 = ~n34179 & n34223;
  assign n35073 = ~n35071 & ~n35072;
  assign n35074 = n35070 & n35073;
  assign n35075 = ~n34218 & ~n35074;
  assign n35076 = ~n34200 & n34226;
  assign n35077 = n34200 & n34222;
  assign n35078 = ~n35076 & ~n35077;
  assign n35079 = ~n34179 & ~n35078;
  assign n35080 = ~n35075 & ~n35079;
  assign n35081 = n35065 & n35080;
  assign n35082 = ~pi0694 & ~n35081;
  assign n35083 = ~n35064 & n35080;
  assign n35084 = pi0694 & n35083;
  assign n35085 = ~n35057 & n35084;
  assign po0733 = n35082 | n35085;
  assign n35087 = ~n34366 & ~n34374;
  assign n35088 = n34316 & ~n35087;
  assign n35089 = n34342 & ~n34349;
  assign n35090 = ~n34379 & ~n34736;
  assign n35091 = ~n34349 & ~n35090;
  assign n35092 = ~n35089 & ~n35091;
  assign n35093 = n34316 & ~n35092;
  assign n35094 = ~n35088 & ~n35093;
  assign n35095 = n34365 & n34739;
  assign n35096 = ~n34741 & ~n35095;
  assign n35097 = ~n34382 & ~n34766;
  assign n35098 = n34349 & ~n35097;
  assign n35099 = n34316 & n35098;
  assign n35100 = n35096 & ~n35099;
  assign n35101 = ~n34380 & ~n34744;
  assign n35102 = n34322 & n34357;
  assign n35103 = ~n34732 & ~n35102;
  assign n35104 = n34349 & ~n35103;
  assign n35105 = n34322 & n34365;
  assign n35106 = n34322 & n34364;
  assign n35107 = ~n34404 & ~n35106;
  assign n35108 = ~n34349 & ~n35107;
  assign n35109 = ~n35105 & ~n35108;
  assign n35110 = ~n35104 & n35109;
  assign n35111 = n35101 & n35110;
  assign n35112 = ~n34316 & ~n35111;
  assign n35113 = ~n34763 & n34784;
  assign n35114 = n34349 & ~n35113;
  assign n35115 = ~n35112 & ~n35114;
  assign n35116 = n35100 & n35115;
  assign n35117 = n35094 & n35116;
  assign n35118 = ~pi0696 & ~n35117;
  assign n35119 = pi0696 & n35100;
  assign n35120 = n35094 & n35119;
  assign n35121 = n35115 & n35120;
  assign po0734 = n35118 | n35121;
  assign n35123 = ~n34192 & n34209;
  assign n35124 = ~n34240 & ~n35123;
  assign n35125 = n34179 & ~n35124;
  assign n35126 = n34200 & n34231;
  assign n35127 = ~n34574 & ~n35126;
  assign n35128 = ~n34179 & ~n35127;
  assign n35129 = ~n34544 & ~n35076;
  assign n35130 = ~n34208 & n35129;
  assign n35131 = ~n35128 & n35130;
  assign n35132 = ~n35125 & n35131;
  assign n35133 = ~n34537 & ~n34570;
  assign n35134 = n35132 & n35133;
  assign n35135 = n34218 & ~n35134;
  assign n35136 = n34193 & n34568;
  assign n35137 = n34249 & ~n35136;
  assign n35138 = ~n34179 & ~n35137;
  assign n35139 = ~n34200 & n34237;
  assign n35140 = ~n35138 & ~n35139;
  assign n35141 = n34186 & n34209;
  assign n35142 = ~n35077 & ~n35141;
  assign n35143 = ~n34179 & ~n35142;
  assign n35144 = ~n34179 & n34231;
  assign n35145 = ~n34200 & n35144;
  assign n35146 = ~n35143 & ~n35145;
  assign n35147 = n35140 & n35146;
  assign n35148 = ~n34218 & ~n35147;
  assign n35149 = ~n34226 & ~n34233;
  assign n35150 = ~n34575 & n35149;
  assign n35151 = n34254 & ~n35150;
  assign n35152 = ~n35148 & ~n35151;
  assign n35153 = ~n34208 & ~n34570;
  assign n35154 = n34179 & ~n35153;
  assign n35155 = n35152 & ~n35154;
  assign n35156 = ~n35135 & n35155;
  assign n35157 = ~pi0687 & n35156;
  assign n35158 = pi0687 & ~n35156;
  assign po0735 = n35157 | n35158;
  assign n35160 = ~n34890 & n35011;
  assign n35161 = ~n34964 & ~n35160;
  assign n35162 = ~n34922 & ~n35161;
  assign n35163 = ~n34890 & n34905;
  assign n35164 = ~n34981 & ~n35163;
  assign n35165 = ~n34922 & ~n35164;
  assign n35166 = ~n34913 & n34931;
  assign n35167 = ~n34906 & ~n35166;
  assign n35168 = ~n34960 & n35167;
  assign n35169 = n34922 & ~n35168;
  assign n35170 = ~n35165 & ~n35169;
  assign n35171 = ~n34936 & ~n34949;
  assign n35172 = n35170 & n35171;
  assign n35173 = n34928 & ~n35172;
  assign n35174 = n34913 & n34981;
  assign n35175 = n34903 & ~n34913;
  assign n35176 = ~n35011 & ~n35175;
  assign n35177 = n34922 & ~n35176;
  assign n35178 = ~n35174 & ~n35177;
  assign n35179 = n34890 & ~n34922;
  assign n35180 = ~n34896 & n35179;
  assign n35181 = n34902 & n35180;
  assign n35182 = n34907 & ~n35181;
  assign n35183 = ~n34960 & n35182;
  assign n35184 = ~n34913 & ~n35183;
  assign n35185 = n35178 & ~n35184;
  assign n35186 = ~n34928 & ~n35185;
  assign n35187 = ~n35173 & ~n35186;
  assign n35188 = ~n34890 & ~n34902;
  assign n35189 = n34953 & n35188;
  assign n35190 = n35187 & ~n35189;
  assign n35191 = ~n35162 & n35190;
  assign n35192 = ~pi0701 & ~n35191;
  assign n35193 = pi0701 & ~n35162;
  assign n35194 = n35187 & n35193;
  assign n35195 = ~n35189 & n35194;
  assign po0736 = n35192 | n35195;
  assign n35197 = ~n34932 & ~n34988;
  assign n35198 = n34929 & ~n35197;
  assign n35199 = n34890 & n34913;
  assign n35200 = ~n34905 & n35199;
  assign n35201 = ~n34928 & n35200;
  assign n35202 = ~n34922 & n34945;
  assign n35203 = n34905 & n35202;
  assign n35204 = n34890 & n34953;
  assign n35205 = ~n34896 & n35204;
  assign n35206 = ~n35203 & ~n35205;
  assign n35207 = ~n35201 & n35206;
  assign n35208 = ~n35011 & ~n35013;
  assign n35209 = ~n34922 & ~n35208;
  assign n35210 = ~n34985 & ~n35209;
  assign n35211 = ~n34928 & ~n35210;
  assign n35212 = ~n34905 & ~n35188;
  assign n35213 = ~n34913 & ~n35212;
  assign n35214 = ~n34981 & ~n35213;
  assign n35215 = n34922 & ~n35214;
  assign n35216 = ~n35005 & ~n35215;
  assign n35217 = n34913 & n34960;
  assign n35218 = ~n34896 & n34914;
  assign n35219 = n34913 & ~n35212;
  assign n35220 = ~n35218 & ~n35219;
  assign n35221 = ~n34922 & ~n35220;
  assign n35222 = ~n35217 & ~n35221;
  assign n35223 = n35216 & n35222;
  assign n35224 = n34928 & ~n35223;
  assign n35225 = ~n35211 & ~n35224;
  assign n35226 = n35207 & n35225;
  assign n35227 = ~n35198 & n35226;
  assign n35228 = pi0707 & ~n35227;
  assign n35229 = ~pi0707 & n35207;
  assign n35230 = ~n35198 & n35229;
  assign n35231 = n35225 & n35230;
  assign po0737 = n35228 | n35231;
  assign n35233 = pi3642 & pi9040;
  assign n35234 = pi3601 & ~pi9040;
  assign n35235 = ~n35233 & ~n35234;
  assign n35236 = pi0704 & n35235;
  assign n35237 = ~pi0704 & ~n35235;
  assign n35238 = ~n35236 & ~n35237;
  assign n35239 = pi3614 & pi9040;
  assign n35240 = pi3603 & ~pi9040;
  assign n35241 = ~n35239 & ~n35240;
  assign n35242 = ~pi0713 & ~n35241;
  assign n35243 = pi0713 & ~n35239;
  assign n35244 = ~n35240 & n35243;
  assign n35245 = ~n35242 & ~n35244;
  assign n35246 = pi3647 & pi9040;
  assign n35247 = pi3607 & ~pi9040;
  assign n35248 = ~n35246 & ~n35247;
  assign n35249 = ~pi0726 & ~n35248;
  assign n35250 = pi0726 & ~n35246;
  assign n35251 = ~n35247 & n35250;
  assign n35252 = ~n35249 & ~n35251;
  assign n35253 = pi3648 & pi9040;
  assign n35254 = pi3652 & ~pi9040;
  assign n35255 = ~n35253 & ~n35254;
  assign n35256 = ~pi0703 & n35255;
  assign n35257 = pi0703 & ~n35255;
  assign n35258 = ~n35256 & ~n35257;
  assign n35259 = n35252 & ~n35258;
  assign n35260 = ~n35245 & n35259;
  assign n35261 = pi3605 & pi9040;
  assign n35262 = pi3624 & ~pi9040;
  assign n35263 = ~n35261 & ~n35262;
  assign n35264 = pi0732 & n35263;
  assign n35265 = ~pi0732 & ~n35263;
  assign n35266 = ~n35264 & ~n35265;
  assign n35267 = n35260 & ~n35266;
  assign n35268 = ~n35252 & n35258;
  assign n35269 = ~n35266 & n35268;
  assign n35270 = ~n35245 & n35269;
  assign n35271 = ~n35267 & ~n35270;
  assign n35272 = n35245 & n35266;
  assign n35273 = n35268 & n35272;
  assign n35274 = n35252 & n35258;
  assign n35275 = ~n35245 & n35274;
  assign n35276 = n35266 & n35275;
  assign n35277 = ~n35273 & ~n35276;
  assign n35278 = n35271 & n35277;
  assign n35279 = n35238 & ~n35278;
  assign n35280 = ~n35245 & n35266;
  assign n35281 = ~n35258 & n35280;
  assign n35282 = ~n35252 & n35281;
  assign n35283 = ~n35275 & ~n35282;
  assign n35284 = n35238 & ~n35283;
  assign n35285 = ~n35258 & ~n35266;
  assign n35286 = ~n35238 & n35285;
  assign n35287 = n35245 & n35252;
  assign n35288 = n35266 & n35268;
  assign n35289 = ~n35287 & ~n35288;
  assign n35290 = ~n35238 & ~n35289;
  assign n35291 = ~n35286 & ~n35290;
  assign n35292 = ~n35252 & ~n35258;
  assign n35293 = n35245 & n35292;
  assign n35294 = ~n35266 & n35293;
  assign n35295 = n35291 & ~n35294;
  assign n35296 = ~n35258 & n35287;
  assign n35297 = n35266 & n35296;
  assign n35298 = n35295 & ~n35297;
  assign n35299 = ~n35284 & n35298;
  assign n35300 = pi3640 & pi9040;
  assign n35301 = pi3619 & ~pi9040;
  assign n35302 = ~n35300 & ~n35301;
  assign n35303 = ~pi0731 & ~n35302;
  assign n35304 = pi0731 & n35302;
  assign n35305 = ~n35303 & ~n35304;
  assign n35306 = ~n35299 & ~n35305;
  assign n35307 = ~n35245 & ~n35258;
  assign n35308 = ~n35238 & n35266;
  assign n35309 = n35305 & n35308;
  assign n35310 = n35307 & n35309;
  assign n35311 = ~n35245 & ~n35266;
  assign n35312 = n35258 & n35311;
  assign n35313 = ~n35238 & ~n35312;
  assign n35314 = ~n35252 & n35272;
  assign n35315 = ~n35259 & ~n35307;
  assign n35316 = ~n35266 & ~n35315;
  assign n35317 = n35245 & n35268;
  assign n35318 = ~n35316 & ~n35317;
  assign n35319 = n35238 & n35318;
  assign n35320 = ~n35314 & n35319;
  assign n35321 = ~n35313 & ~n35320;
  assign n35322 = n35245 & n35274;
  assign n35323 = n35266 & n35322;
  assign n35324 = ~n35321 & ~n35323;
  assign n35325 = n35305 & ~n35324;
  assign n35326 = ~n35310 & ~n35325;
  assign n35327 = ~n35306 & n35326;
  assign n35328 = ~n35279 & n35327;
  assign n35329 = ~n35238 & n35294;
  assign n35330 = n35328 & ~n35329;
  assign n35331 = pi0736 & ~n35330;
  assign n35332 = n35327 & ~n35329;
  assign n35333 = ~pi0736 & n35332;
  assign n35334 = ~n35279 & n35333;
  assign po0764 = n35331 | n35334;
  assign n35336 = pi3600 & ~pi9040;
  assign n35337 = pi3603 & pi9040;
  assign n35338 = ~n35336 & ~n35337;
  assign n35339 = ~pi0735 & ~n35338;
  assign n35340 = pi0735 & n35338;
  assign n35341 = ~n35339 & ~n35340;
  assign n35342 = pi3617 & pi9040;
  assign n35343 = pi3642 & ~pi9040;
  assign n35344 = ~n35342 & ~n35343;
  assign n35345 = ~pi0716 & n35344;
  assign n35346 = pi0716 & ~n35344;
  assign n35347 = ~n35345 & ~n35346;
  assign n35348 = pi3607 & pi9040;
  assign n35349 = pi3614 & ~pi9040;
  assign n35350 = ~n35348 & ~n35349;
  assign n35351 = ~pi0708 & ~n35350;
  assign n35352 = pi0708 & ~n35348;
  assign n35353 = ~n35349 & n35352;
  assign n35354 = ~n35351 & ~n35353;
  assign n35355 = pi3631 & pi9040;
  assign n35356 = pi3608 & ~pi9040;
  assign n35357 = ~n35355 & ~n35356;
  assign n35358 = ~pi0727 & ~n35357;
  assign n35359 = pi0727 & n35357;
  assign n35360 = ~n35358 & ~n35359;
  assign n35361 = pi3643 & pi9040;
  assign n35362 = pi3599 & ~pi9040;
  assign n35363 = ~n35361 & ~n35362;
  assign n35364 = ~pi0710 & ~n35363;
  assign n35365 = pi0710 & n35363;
  assign n35366 = ~n35364 & ~n35365;
  assign n35367 = n35360 & ~n35366;
  assign n35368 = n35354 & n35367;
  assign n35369 = pi3619 & pi9040;
  assign n35370 = pi3646 & ~pi9040;
  assign n35371 = ~n35369 & ~n35370;
  assign n35372 = ~pi0712 & ~n35371;
  assign n35373 = pi0712 & ~n35369;
  assign n35374 = ~n35370 & n35373;
  assign n35375 = ~n35372 & ~n35374;
  assign n35376 = n35366 & n35375;
  assign n35377 = n35360 & n35376;
  assign n35378 = ~n35368 & ~n35377;
  assign n35379 = n35366 & ~n35375;
  assign n35380 = ~n35360 & n35379;
  assign n35381 = ~n35354 & n35380;
  assign n35382 = n35378 & ~n35381;
  assign n35383 = ~n35347 & ~n35382;
  assign n35384 = ~n35360 & n35366;
  assign n35385 = ~n35354 & n35375;
  assign n35386 = n35384 & n35385;
  assign n35387 = ~n35366 & n35375;
  assign n35388 = n35360 & n35387;
  assign n35389 = ~n35354 & n35388;
  assign n35390 = ~n35360 & ~n35366;
  assign n35391 = ~n35379 & ~n35390;
  assign n35392 = n35354 & ~n35391;
  assign n35393 = ~n35389 & ~n35392;
  assign n35394 = ~n35386 & n35393;
  assign n35395 = n35347 & ~n35394;
  assign n35396 = ~n35383 & ~n35395;
  assign n35397 = n35341 & ~n35396;
  assign n35398 = ~n35366 & ~n35375;
  assign n35399 = ~n35360 & n35398;
  assign n35400 = n35347 & ~n35354;
  assign n35401 = n35399 & n35400;
  assign n35402 = n35379 & n35400;
  assign n35403 = n35360 & n35402;
  assign n35404 = ~n35401 & ~n35403;
  assign n35405 = ~n35354 & ~n35360;
  assign n35406 = n35375 & n35405;
  assign n35407 = ~n35366 & n35406;
  assign n35408 = ~n35347 & n35407;
  assign n35409 = n35404 & ~n35408;
  assign n35410 = ~n35347 & ~n35354;
  assign n35411 = ~n35366 & n35410;
  assign n35412 = n35347 & n35379;
  assign n35413 = ~n35354 & n35412;
  assign n35414 = ~n35354 & n35360;
  assign n35415 = n35366 & n35414;
  assign n35416 = ~n35368 & ~n35415;
  assign n35417 = n35347 & ~n35416;
  assign n35418 = ~n35413 & ~n35417;
  assign n35419 = n35360 & n35379;
  assign n35420 = ~n35354 & n35419;
  assign n35421 = n35375 & n35384;
  assign n35422 = n35354 & n35421;
  assign n35423 = ~n35420 & ~n35422;
  assign n35424 = ~n35347 & n35354;
  assign n35425 = n35384 & n35424;
  assign n35426 = ~n35360 & n35387;
  assign n35427 = ~n35347 & n35426;
  assign n35428 = ~n35425 & ~n35427;
  assign n35429 = n35423 & n35428;
  assign n35430 = n35418 & n35429;
  assign n35431 = ~n35411 & n35430;
  assign n35432 = ~n35341 & ~n35431;
  assign n35433 = n35354 & n35376;
  assign n35434 = n35360 & n35398;
  assign n35435 = ~n35354 & n35434;
  assign n35436 = ~n35433 & ~n35435;
  assign n35437 = ~n35347 & ~n35436;
  assign n35438 = ~n35432 & ~n35437;
  assign n35439 = n35409 & n35438;
  assign n35440 = ~n35397 & n35439;
  assign n35441 = ~pi0748 & ~n35440;
  assign n35442 = pi0748 & n35440;
  assign po0766 = n35441 | n35442;
  assign n35444 = ~n35341 & n35347;
  assign n35445 = ~n35354 & n35367;
  assign n35446 = n35354 & n35419;
  assign n35447 = ~n35354 & n35376;
  assign n35448 = ~n35446 & ~n35447;
  assign n35449 = ~n35445 & n35448;
  assign n35450 = n35444 & ~n35449;
  assign n35451 = ~n35375 & n35405;
  assign n35452 = n35354 & n35434;
  assign n35453 = ~n35451 & ~n35452;
  assign n35454 = ~n35377 & ~n35380;
  assign n35455 = n35453 & n35454;
  assign n35456 = ~n35347 & ~n35455;
  assign n35457 = n35354 & n35426;
  assign n35458 = ~n35456 & ~n35457;
  assign n35459 = ~n35341 & ~n35458;
  assign n35460 = ~n35450 & ~n35459;
  assign n35461 = n35360 & n35410;
  assign n35462 = n35375 & n35461;
  assign n35463 = ~n35381 & ~n35462;
  assign n35464 = ~n35376 & ~n35398;
  assign n35465 = n35354 & ~n35464;
  assign n35466 = ~n35399 & ~n35465;
  assign n35467 = n35347 & ~n35466;
  assign n35468 = ~n35388 & ~n35445;
  assign n35469 = ~n35446 & n35468;
  assign n35470 = ~n35347 & ~n35469;
  assign n35471 = ~n35467 & ~n35470;
  assign n35472 = n35354 & n35399;
  assign n35473 = ~n35422 & ~n35472;
  assign n35474 = ~n35407 & n35473;
  assign n35475 = ~n35413 & n35474;
  assign n35476 = n35471 & n35475;
  assign n35477 = n35341 & ~n35476;
  assign n35478 = n35463 & ~n35477;
  assign n35479 = n35460 & n35478;
  assign n35480 = pi0739 & ~n35479;
  assign n35481 = ~pi0739 & n35463;
  assign n35482 = n35460 & n35481;
  assign n35483 = ~n35477 & n35482;
  assign po0768 = n35480 | n35483;
  assign n35485 = pi3622 & pi9040;
  assign n35486 = pi3597 & ~pi9040;
  assign n35487 = ~n35485 & ~n35486;
  assign n35488 = ~pi0730 & n35487;
  assign n35489 = pi0730 & ~n35487;
  assign n35490 = ~n35488 & ~n35489;
  assign n35491 = pi3654 & pi9040;
  assign n35492 = pi3628 & ~pi9040;
  assign n35493 = ~n35491 & ~n35492;
  assign n35494 = ~pi0728 & ~n35493;
  assign n35495 = pi0728 & ~n35491;
  assign n35496 = ~n35492 & n35495;
  assign n35497 = ~n35494 & ~n35496;
  assign n35498 = pi3621 & pi9040;
  assign n35499 = pi3649 & ~pi9040;
  assign n35500 = ~n35498 & ~n35499;
  assign n35501 = pi0723 & n35500;
  assign n35502 = ~pi0723 & ~n35500;
  assign n35503 = ~n35501 & ~n35502;
  assign n35504 = n35497 & ~n35503;
  assign n35505 = pi3626 & pi9040;
  assign n35506 = pi3622 & ~pi9040;
  assign n35507 = ~n35505 & ~n35506;
  assign n35508 = pi0733 & n35507;
  assign n35509 = ~pi0733 & ~n35507;
  assign n35510 = ~n35508 & ~n35509;
  assign n35511 = pi3629 & pi9040;
  assign n35512 = pi3635 & ~pi9040;
  assign n35513 = ~n35511 & ~n35512;
  assign n35514 = ~pi0691 & ~n35513;
  assign n35515 = pi0691 & ~n35511;
  assign n35516 = ~n35512 & n35515;
  assign n35517 = ~n35514 & ~n35516;
  assign n35518 = n35510 & n35517;
  assign n35519 = n35504 & n35518;
  assign n35520 = n35510 & ~n35517;
  assign n35521 = ~n35497 & n35520;
  assign n35522 = ~n35519 & ~n35521;
  assign n35523 = n35490 & ~n35522;
  assign n35524 = pi3609 & ~pi9040;
  assign n35525 = pi3630 & pi9040;
  assign n35526 = ~n35524 & ~n35525;
  assign n35527 = ~pi0717 & ~n35526;
  assign n35528 = pi0717 & n35526;
  assign n35529 = ~n35527 & ~n35528;
  assign n35530 = ~n35490 & ~n35510;
  assign n35531 = n35497 & n35530;
  assign n35532 = n35504 & ~n35517;
  assign n35533 = n35497 & n35503;
  assign n35534 = n35517 & n35533;
  assign n35535 = ~n35532 & ~n35534;
  assign n35536 = ~n35497 & ~n35503;
  assign n35537 = n35517 & n35536;
  assign n35538 = n35510 & n35537;
  assign n35539 = n35535 & ~n35538;
  assign n35540 = ~n35490 & ~n35539;
  assign n35541 = ~n35531 & ~n35540;
  assign n35542 = ~n35497 & n35503;
  assign n35543 = ~n35517 & n35542;
  assign n35544 = n35510 & n35543;
  assign n35545 = n35541 & ~n35544;
  assign n35546 = ~n35510 & n35536;
  assign n35547 = ~n35497 & n35517;
  assign n35548 = n35503 & n35547;
  assign n35549 = ~n35546 & ~n35548;
  assign n35550 = n35490 & ~n35549;
  assign n35551 = ~n35517 & n35533;
  assign n35552 = ~n35510 & n35551;
  assign n35553 = ~n35550 & ~n35552;
  assign n35554 = n35545 & n35553;
  assign n35555 = n35529 & ~n35554;
  assign n35556 = ~n35523 & ~n35555;
  assign n35557 = ~n35490 & ~n35529;
  assign n35558 = ~n35549 & n35557;
  assign n35559 = ~n35517 & n35536;
  assign n35560 = ~n35551 & ~n35559;
  assign n35561 = n35510 & ~n35560;
  assign n35562 = ~n35519 & ~n35561;
  assign n35563 = ~n35529 & ~n35562;
  assign n35564 = ~n35558 & ~n35563;
  assign n35565 = n35490 & ~n35529;
  assign n35566 = n35504 & ~n35510;
  assign n35567 = ~n35543 & ~n35566;
  assign n35568 = n35497 & n35517;
  assign n35569 = n35567 & ~n35568;
  assign n35570 = n35565 & ~n35569;
  assign n35571 = n35564 & ~n35570;
  assign n35572 = n35556 & n35571;
  assign n35573 = ~pi0740 & ~n35572;
  assign n35574 = pi0740 & n35564;
  assign n35575 = n35556 & n35574;
  assign n35576 = ~n35570 & n35575;
  assign po0769 = n35573 | n35576;
  assign n35578 = pi3612 & pi9040;
  assign n35579 = pi3626 & ~pi9040;
  assign n35580 = ~n35578 & ~n35579;
  assign n35581 = ~pi0722 & n35580;
  assign n35582 = pi0722 & ~n35580;
  assign n35583 = ~n35581 & ~n35582;
  assign n35584 = pi3698 & pi9040;
  assign n35585 = pi3612 & ~pi9040;
  assign n35586 = ~n35584 & ~n35585;
  assign n35587 = ~pi0691 & n35586;
  assign n35588 = pi0691 & ~n35586;
  assign n35589 = ~n35587 & ~n35588;
  assign n35590 = pi3627 & pi9040;
  assign n35591 = pi3620 & ~pi9040;
  assign n35592 = ~n35590 & ~n35591;
  assign n35593 = ~pi0726 & n35592;
  assign n35594 = pi0726 & ~n35592;
  assign n35595 = ~n35593 & ~n35594;
  assign n35596 = pi3653 & pi9040;
  assign n35597 = pi3604 & ~pi9040;
  assign n35598 = ~n35596 & ~n35597;
  assign n35599 = pi0706 & n35598;
  assign n35600 = ~pi0706 & ~n35598;
  assign n35601 = ~n35599 & ~n35600;
  assign n35602 = ~n35595 & ~n35601;
  assign n35603 = n35589 & n35602;
  assign n35604 = pi3625 & pi9040;
  assign n35605 = pi3698 & ~pi9040;
  assign n35606 = ~n35604 & ~n35605;
  assign n35607 = ~pi0731 & n35606;
  assign n35608 = pi0731 & ~n35606;
  assign n35609 = ~n35607 & ~n35608;
  assign n35610 = ~n35595 & ~n35609;
  assign n35611 = ~n35589 & n35610;
  assign n35612 = n35601 & n35611;
  assign n35613 = ~n35603 & ~n35612;
  assign n35614 = ~n35589 & n35609;
  assign n35615 = n35595 & n35614;
  assign n35616 = n35601 & n35615;
  assign n35617 = n35613 & ~n35616;
  assign n35618 = n35583 & ~n35617;
  assign n35619 = pi3649 & pi9040;
  assign n35620 = pi3602 & ~pi9040;
  assign n35621 = ~n35619 & ~n35620;
  assign n35622 = ~pi0728 & ~n35621;
  assign n35623 = pi0728 & n35621;
  assign n35624 = ~n35622 & ~n35623;
  assign n35625 = ~n35583 & n35601;
  assign n35626 = n35614 & n35625;
  assign n35627 = ~n35595 & n35626;
  assign n35628 = ~n35583 & ~n35601;
  assign n35629 = ~n35589 & ~n35609;
  assign n35630 = n35628 & n35629;
  assign n35631 = n35589 & ~n35609;
  assign n35632 = ~n35595 & n35631;
  assign n35633 = ~n35583 & n35632;
  assign n35634 = n35601 & n35633;
  assign n35635 = n35589 & n35609;
  assign n35636 = ~n35595 & n35635;
  assign n35637 = ~n35601 & n35636;
  assign n35638 = ~n35634 & ~n35637;
  assign n35639 = ~n35630 & n35638;
  assign n35640 = ~n35627 & n35639;
  assign n35641 = n35595 & ~n35601;
  assign n35642 = ~n35589 & n35641;
  assign n35643 = ~n35609 & n35642;
  assign n35644 = n35640 & ~n35643;
  assign n35645 = ~n35624 & ~n35644;
  assign n35646 = n35589 & n35595;
  assign n35647 = ~n35609 & n35646;
  assign n35648 = n35583 & n35647;
  assign n35649 = n35601 & n35648;
  assign n35650 = n35602 & n35609;
  assign n35651 = ~n35601 & n35635;
  assign n35652 = ~n35650 & ~n35651;
  assign n35653 = n35583 & ~n35652;
  assign n35654 = ~n35649 & ~n35653;
  assign n35655 = ~n35624 & ~n35654;
  assign n35656 = ~n35645 & ~n35655;
  assign n35657 = ~n35618 & n35656;
  assign n35658 = n35595 & n35601;
  assign n35659 = ~n35583 & n35658;
  assign n35660 = n35635 & n35659;
  assign n35661 = n35595 & ~n35609;
  assign n35662 = n35628 & n35661;
  assign n35663 = n35583 & n35610;
  assign n35664 = n35601 & n35609;
  assign n35665 = n35595 & n35664;
  assign n35666 = ~n35615 & ~n35665;
  assign n35667 = ~n35663 & n35666;
  assign n35668 = ~n35601 & n35647;
  assign n35669 = n35667 & ~n35668;
  assign n35670 = ~n35583 & n35614;
  assign n35671 = ~n35601 & n35670;
  assign n35672 = ~n35589 & n35595;
  assign n35673 = n35601 & n35635;
  assign n35674 = ~n35672 & ~n35673;
  assign n35675 = ~n35583 & ~n35674;
  assign n35676 = ~n35671 & ~n35675;
  assign n35677 = n35669 & n35676;
  assign n35678 = n35624 & ~n35677;
  assign n35679 = ~n35662 & ~n35678;
  assign n35680 = ~n35660 & n35679;
  assign n35681 = n35657 & n35680;
  assign n35682 = pi0742 & n35681;
  assign n35683 = ~pi0742 & ~n35681;
  assign po0772 = n35682 | n35683;
  assign n35685 = ~n35595 & n35609;
  assign n35686 = ~n35643 & ~n35685;
  assign n35687 = ~n35664 & n35686;
  assign n35688 = ~n35583 & ~n35687;
  assign n35689 = n35583 & n35601;
  assign n35690 = ~n35609 & n35689;
  assign n35691 = ~n35595 & n35601;
  assign n35692 = ~n35589 & n35691;
  assign n35693 = ~n35601 & n35632;
  assign n35694 = ~n35692 & ~n35693;
  assign n35695 = n35595 & n35609;
  assign n35696 = n35583 & ~n35601;
  assign n35697 = n35695 & n35696;
  assign n35698 = n35694 & ~n35697;
  assign n35699 = ~n35690 & n35698;
  assign n35700 = ~n35688 & n35699;
  assign n35701 = n35624 & ~n35700;
  assign n35702 = ~n35595 & n35614;
  assign n35703 = ~n35601 & n35702;
  assign n35704 = n35601 & n35636;
  assign n35705 = ~n35703 & ~n35704;
  assign n35706 = ~n35583 & ~n35705;
  assign n35707 = ~n35701 & ~n35706;
  assign n35708 = n35601 & n35632;
  assign n35709 = ~n35611 & ~n35647;
  assign n35710 = ~n35583 & ~n35709;
  assign n35711 = ~n35708 & ~n35710;
  assign n35712 = ~n35616 & n35711;
  assign n35713 = ~n35624 & ~n35712;
  assign n35714 = ~n35629 & ~n35635;
  assign n35715 = n35595 & ~n35714;
  assign n35716 = ~n35651 & ~n35715;
  assign n35717 = n35583 & ~n35716;
  assign n35718 = ~n35624 & n35717;
  assign n35719 = ~n35713 & ~n35718;
  assign n35720 = n35707 & n35719;
  assign n35721 = pi0749 & ~n35720;
  assign n35722 = ~pi0749 & n35707;
  assign n35723 = n35719 & n35722;
  assign po0773 = n35721 | n35723;
  assign n35725 = n35490 & n35510;
  assign n35726 = ~n35536 & ~n35551;
  assign n35727 = n35725 & ~n35726;
  assign n35728 = n35490 & ~n35517;
  assign n35729 = n35536 & n35728;
  assign n35730 = ~n35727 & ~n35729;
  assign n35731 = n35529 & ~n35730;
  assign n35732 = ~n35510 & n35517;
  assign n35733 = n35503 & n35732;
  assign n35734 = n35497 & n35733;
  assign n35735 = ~n35568 & ~n35732;
  assign n35736 = ~n35490 & ~n35735;
  assign n35737 = ~n35510 & ~n35517;
  assign n35738 = ~n35503 & n35737;
  assign n35739 = n35497 & n35738;
  assign n35740 = ~n35736 & ~n35739;
  assign n35741 = ~n35734 & n35740;
  assign n35742 = n35529 & ~n35741;
  assign n35743 = ~n35731 & ~n35742;
  assign n35744 = n35503 & n35518;
  assign n35745 = ~n35497 & n35744;
  assign n35746 = ~n35510 & n35543;
  assign n35747 = ~n35745 & ~n35746;
  assign n35748 = n35490 & ~n35747;
  assign n35749 = n35510 & n35559;
  assign n35750 = ~n35510 & n35568;
  assign n35751 = ~n35749 & ~n35750;
  assign n35752 = ~n35490 & ~n35751;
  assign n35753 = ~n35504 & ~n35568;
  assign n35754 = n35510 & ~n35753;
  assign n35755 = ~n35543 & ~n35754;
  assign n35756 = n35490 & ~n35755;
  assign n35757 = n35503 & ~n35510;
  assign n35758 = n35490 & n35757;
  assign n35759 = ~n35517 & n35758;
  assign n35760 = ~n35503 & n35517;
  assign n35761 = ~n35543 & ~n35760;
  assign n35762 = ~n35510 & ~n35761;
  assign n35763 = ~n35490 & n35510;
  assign n35764 = n35533 & n35763;
  assign n35765 = ~n35517 & n35764;
  assign n35766 = ~n35762 & ~n35765;
  assign n35767 = ~n35759 & n35766;
  assign n35768 = ~n35756 & n35767;
  assign n35769 = ~n35745 & n35768;
  assign n35770 = ~n35529 & ~n35769;
  assign n35771 = ~n35752 & ~n35770;
  assign n35772 = ~n35748 & n35771;
  assign n35773 = n35743 & n35772;
  assign n35774 = pi0750 & n35773;
  assign n35775 = ~pi0750 & ~n35773;
  assign po0774 = n35774 | n35775;
  assign n35777 = ~n35388 & ~n35399;
  assign n35778 = n35347 & ~n35777;
  assign n35779 = n35354 & n35377;
  assign n35780 = ~n35778 & ~n35779;
  assign n35781 = n35354 & n35366;
  assign n35782 = ~n35384 & ~n35781;
  assign n35783 = ~n35434 & n35782;
  assign n35784 = ~n35347 & ~n35783;
  assign n35785 = n35780 & ~n35784;
  assign n35786 = ~n35341 & ~n35785;
  assign n35787 = ~n35354 & n35421;
  assign n35788 = n35347 & n35787;
  assign n35789 = ~n35403 & ~n35788;
  assign n35790 = ~n35408 & n35789;
  assign n35791 = ~n35347 & n35366;
  assign n35792 = n35414 & n35791;
  assign n35793 = n35354 & n35388;
  assign n35794 = n35347 & n35384;
  assign n35795 = ~n35793 & ~n35794;
  assign n35796 = ~n35472 & n35795;
  assign n35797 = ~n35792 & n35796;
  assign n35798 = ~n35375 & n35414;
  assign n35799 = ~n35407 & ~n35798;
  assign n35800 = n35797 & n35799;
  assign n35801 = ~n35427 & n35800;
  assign n35802 = n35341 & ~n35801;
  assign n35803 = n35790 & ~n35802;
  assign n35804 = ~n35786 & n35803;
  assign n35805 = ~pi0746 & ~n35804;
  assign n35806 = pi0746 & n35790;
  assign n35807 = ~n35786 & n35806;
  assign n35808 = ~n35802 & n35807;
  assign po0775 = n35805 | n35808;
  assign n35810 = pi3636 & pi9040;
  assign n35811 = pi3606 & ~pi9040;
  assign n35812 = ~n35810 & ~n35811;
  assign n35813 = pi0710 & n35812;
  assign n35814 = ~pi0710 & ~n35812;
  assign n35815 = ~n35813 & ~n35814;
  assign n35816 = pi3608 & pi9040;
  assign n35817 = pi3605 & ~pi9040;
  assign n35818 = ~n35816 & ~n35817;
  assign n35819 = ~pi0724 & n35818;
  assign n35820 = pi0724 & ~n35818;
  assign n35821 = ~n35819 & ~n35820;
  assign n35822 = pi3624 & pi9040;
  assign n35823 = pi3647 & ~pi9040;
  assign n35824 = ~n35822 & ~n35823;
  assign n35825 = ~pi0734 & ~n35824;
  assign n35826 = pi0734 & ~n35822;
  assign n35827 = ~n35823 & n35826;
  assign n35828 = ~n35825 & ~n35827;
  assign n35829 = pi3600 & pi9040;
  assign n35830 = pi3651 & ~pi9040;
  assign n35831 = ~n35829 & ~n35830;
  assign n35832 = pi0705 & n35831;
  assign n35833 = ~pi0705 & ~n35831;
  assign n35834 = ~n35832 & ~n35833;
  assign n35835 = pi3601 & pi9040;
  assign n35836 = pi3648 & ~pi9040;
  assign n35837 = ~n35835 & ~n35836;
  assign n35838 = pi0727 & n35837;
  assign n35839 = ~pi0727 & ~n35837;
  assign n35840 = ~n35838 & ~n35839;
  assign n35841 = n35834 & ~n35840;
  assign n35842 = n35828 & n35841;
  assign n35843 = ~n35821 & n35842;
  assign n35844 = pi3652 & pi9040;
  assign n35845 = pi3610 & ~pi9040;
  assign n35846 = ~n35844 & ~n35845;
  assign n35847 = pi0721 & n35846;
  assign n35848 = ~pi0721 & ~n35846;
  assign n35849 = ~n35847 & ~n35848;
  assign n35850 = n35828 & n35840;
  assign n35851 = n35834 & n35850;
  assign n35852 = ~n35828 & ~n35834;
  assign n35853 = ~n35834 & ~n35840;
  assign n35854 = n35821 & n35853;
  assign n35855 = ~n35828 & ~n35840;
  assign n35856 = ~n35821 & n35855;
  assign n35857 = ~n35854 & ~n35856;
  assign n35858 = ~n35852 & n35857;
  assign n35859 = ~n35851 & n35858;
  assign n35860 = n35849 & ~n35859;
  assign n35861 = n35821 & n35834;
  assign n35862 = n35840 & n35861;
  assign n35863 = ~n35828 & n35861;
  assign n35864 = ~n35834 & n35850;
  assign n35865 = ~n35863 & ~n35864;
  assign n35866 = ~n35849 & ~n35865;
  assign n35867 = ~n35862 & ~n35866;
  assign n35868 = ~n35860 & n35867;
  assign n35869 = ~n35843 & n35868;
  assign n35870 = n35815 & ~n35869;
  assign n35871 = ~n35828 & n35840;
  assign n35872 = ~n35834 & n35871;
  assign n35873 = n35821 & n35872;
  assign n35874 = ~n35834 & n35855;
  assign n35875 = ~n35821 & n35874;
  assign n35876 = ~n35843 & ~n35875;
  assign n35877 = ~n35873 & n35876;
  assign n35878 = n35849 & ~n35877;
  assign n35879 = ~n35870 & ~n35878;
  assign n35880 = n35821 & n35851;
  assign n35881 = ~n35821 & ~n35834;
  assign n35882 = ~n35849 & n35881;
  assign n35883 = n35828 & n35882;
  assign n35884 = n35834 & n35871;
  assign n35885 = ~n35821 & n35884;
  assign n35886 = n35841 & n35849;
  assign n35887 = n35821 & n35886;
  assign n35888 = ~n35885 & ~n35887;
  assign n35889 = ~n35828 & n35834;
  assign n35890 = ~n35821 & n35889;
  assign n35891 = n35828 & ~n35840;
  assign n35892 = ~n35834 & n35891;
  assign n35893 = ~n35890 & ~n35892;
  assign n35894 = ~n35849 & ~n35893;
  assign n35895 = ~n35849 & n35852;
  assign n35896 = n35821 & n35895;
  assign n35897 = ~n35894 & ~n35896;
  assign n35898 = n35888 & n35897;
  assign n35899 = ~n35815 & ~n35898;
  assign n35900 = ~n35883 & ~n35899;
  assign n35901 = ~n35880 & n35900;
  assign n35902 = n35879 & n35901;
  assign n35903 = ~pi0756 & ~n35902;
  assign n35904 = ~n35870 & ~n35880;
  assign n35905 = ~n35878 & n35904;
  assign n35906 = n35900 & n35905;
  assign n35907 = pi0756 & n35906;
  assign po0776 = n35903 | n35907;
  assign n35909 = pi3618 & ~pi9040;
  assign n35910 = pi3644 & pi9040;
  assign n35911 = ~n35909 & ~n35910;
  assign n35912 = ~pi0734 & ~n35911;
  assign n35913 = pi0734 & n35911;
  assign n35914 = ~n35912 & ~n35913;
  assign n35915 = pi3637 & pi9040;
  assign n35916 = pi3623 & ~pi9040;
  assign n35917 = ~n35915 & ~n35916;
  assign n35918 = ~pi0719 & n35917;
  assign n35919 = pi0719 & ~n35917;
  assign n35920 = ~n35918 & ~n35919;
  assign n35921 = pi3650 & pi9040;
  assign n35922 = pi3633 & ~pi9040;
  assign n35923 = ~n35921 & ~n35922;
  assign n35924 = ~pi0715 & n35923;
  assign n35925 = pi0715 & ~n35923;
  assign n35926 = ~n35924 & ~n35925;
  assign n35927 = pi3632 & pi9040;
  assign n35928 = pi3650 & ~pi9040;
  assign n35929 = ~n35927 & ~n35928;
  assign n35930 = ~pi0718 & ~n35929;
  assign n35931 = pi0718 & n35929;
  assign n35932 = ~n35930 & ~n35931;
  assign n35933 = pi3604 & pi9040;
  assign n35934 = pi3630 & ~pi9040;
  assign n35935 = ~n35933 & ~n35934;
  assign n35936 = ~pi0705 & n35935;
  assign n35937 = pi0705 & ~n35935;
  assign n35938 = ~n35936 & ~n35937;
  assign n35939 = ~n35932 & ~n35938;
  assign n35940 = ~n35926 & n35939;
  assign n35941 = ~n35920 & n35940;
  assign n35942 = pi3602 & pi9040;
  assign n35943 = pi3653 & ~pi9040;
  assign n35944 = ~n35942 & ~n35943;
  assign n35945 = pi0725 & n35944;
  assign n35946 = ~pi0725 & ~n35944;
  assign n35947 = ~n35945 & ~n35946;
  assign n35948 = n35932 & ~n35938;
  assign n35949 = ~n35920 & n35948;
  assign n35950 = n35926 & n35939;
  assign n35951 = n35920 & n35950;
  assign n35952 = ~n35949 & ~n35951;
  assign n35953 = ~n35947 & ~n35952;
  assign n35954 = ~n35941 & ~n35953;
  assign n35955 = n35926 & ~n35932;
  assign n35956 = n35938 & n35955;
  assign n35957 = n35947 & n35956;
  assign n35958 = n35939 & n35947;
  assign n35959 = ~n35920 & n35958;
  assign n35960 = ~n35957 & ~n35959;
  assign n35961 = n35954 & n35960;
  assign n35962 = n35932 & n35938;
  assign n35963 = ~n35926 & n35962;
  assign n35964 = ~n35920 & n35963;
  assign n35965 = ~n35932 & n35938;
  assign n35966 = ~n35926 & n35965;
  assign n35967 = n35920 & n35966;
  assign n35968 = ~n35964 & ~n35967;
  assign n35969 = n35961 & n35968;
  assign n35970 = n35914 & ~n35969;
  assign n35971 = ~n35914 & ~n35947;
  assign n35972 = ~n35920 & n35926;
  assign n35973 = ~n35932 & n35972;
  assign n35974 = n35926 & n35938;
  assign n35975 = ~n35973 & ~n35974;
  assign n35976 = n35971 & ~n35975;
  assign n35977 = n35920 & ~n35926;
  assign n35978 = ~n35938 & n35977;
  assign n35979 = ~n35932 & n35978;
  assign n35980 = n35920 & n35932;
  assign n35981 = n35926 & n35980;
  assign n35982 = ~n35979 & ~n35981;
  assign n35983 = ~n35920 & n35947;
  assign n35984 = ~n35926 & n35983;
  assign n35985 = ~n35939 & n35984;
  assign n35986 = n35947 & n35963;
  assign n35987 = ~n35985 & ~n35986;
  assign n35988 = n35982 & n35987;
  assign n35989 = ~n35914 & ~n35988;
  assign n35990 = n35926 & n35962;
  assign n35991 = n35920 & ~n35947;
  assign n35992 = n35990 & n35991;
  assign n35993 = ~n35926 & n35948;
  assign n35994 = n35920 & n35993;
  assign n35995 = ~n35967 & ~n35994;
  assign n35996 = ~n35947 & ~n35995;
  assign n35997 = ~n35992 & ~n35996;
  assign n35998 = n35947 & n35979;
  assign n35999 = n35997 & ~n35998;
  assign n36000 = ~n35989 & n35999;
  assign n36001 = ~n35976 & n36000;
  assign n36002 = ~n35970 & n36001;
  assign n36003 = n35926 & n35948;
  assign n36004 = n35920 & n35947;
  assign n36005 = n36003 & n36004;
  assign n36006 = n36002 & ~n36005;
  assign n36007 = ~pi0757 & ~n36006;
  assign n36008 = pi0757 & ~n36005;
  assign n36009 = n36001 & n36008;
  assign n36010 = ~n35970 & n36009;
  assign po0777 = n36007 | n36010;
  assign n36012 = n35821 & ~n35849;
  assign n36013 = n35828 & n36012;
  assign n36014 = n35834 & n35855;
  assign n36015 = ~n35821 & n36014;
  assign n36016 = ~n35821 & n35872;
  assign n36017 = ~n36015 & ~n36016;
  assign n36018 = n35821 & ~n35834;
  assign n36019 = ~n35840 & n36018;
  assign n36020 = ~n35828 & n36019;
  assign n36021 = ~n35864 & ~n36020;
  assign n36022 = n35849 & ~n36021;
  assign n36023 = n36017 & ~n36022;
  assign n36024 = ~n36013 & n36023;
  assign n36025 = n35815 & ~n36024;
  assign n36026 = ~n35821 & n35828;
  assign n36027 = ~n35834 & n36026;
  assign n36028 = ~n35840 & n36027;
  assign n36029 = ~n35849 & n36028;
  assign n36030 = n35821 & n35849;
  assign n36031 = n35892 & n36030;
  assign n36032 = ~n35863 & ~n36031;
  assign n36033 = ~n35864 & ~n35884;
  assign n36034 = n35821 & n35871;
  assign n36035 = n36033 & ~n36034;
  assign n36036 = ~n35849 & ~n36035;
  assign n36037 = n35849 & n35851;
  assign n36038 = n35876 & ~n36037;
  assign n36039 = ~n36036 & n36038;
  assign n36040 = n36032 & n36039;
  assign n36041 = ~n35815 & ~n36040;
  assign n36042 = ~n36029 & ~n36041;
  assign n36043 = ~n36025 & n36042;
  assign n36044 = n35884 & n36030;
  assign n36045 = ~n35821 & n35886;
  assign n36046 = ~n36044 & ~n36045;
  assign n36047 = n35849 & n36016;
  assign n36048 = n36046 & ~n36047;
  assign n36049 = n36043 & n36048;
  assign n36050 = ~pi0752 & ~n36049;
  assign n36051 = pi0752 & n36048;
  assign n36052 = n36042 & n36051;
  assign n36053 = ~n36025 & n36052;
  assign po0778 = n36050 | n36053;
  assign n36055 = pi3620 & pi9040;
  assign n36056 = pi3637 & ~pi9040;
  assign n36057 = ~n36055 & ~n36056;
  assign n36058 = ~pi0715 & n36057;
  assign n36059 = pi0715 & ~n36057;
  assign n36060 = ~n36058 & ~n36059;
  assign n36061 = pi3609 & pi9040;
  assign n36062 = pi3654 & ~pi9040;
  assign n36063 = ~n36061 & ~n36062;
  assign n36064 = pi0711 & n36063;
  assign n36065 = ~pi0711 & ~n36063;
  assign n36066 = ~n36064 & ~n36065;
  assign n36067 = pi3635 & pi9040;
  assign n36068 = pi3621 & ~pi9040;
  assign n36069 = ~n36067 & ~n36068;
  assign n36070 = ~pi0723 & ~n36069;
  assign n36071 = pi0723 & n36069;
  assign n36072 = ~n36070 & ~n36071;
  assign n36073 = ~n36066 & n36072;
  assign n36074 = ~n36060 & n36073;
  assign n36075 = pi3634 & pi9040;
  assign n36076 = pi3625 & ~pi9040;
  assign n36077 = ~n36075 & ~n36076;
  assign n36078 = ~pi0717 & ~n36077;
  assign n36079 = pi0717 & ~n36075;
  assign n36080 = ~n36076 & n36079;
  assign n36081 = ~n36078 & ~n36080;
  assign n36082 = ~n36060 & n36081;
  assign n36083 = n36072 & n36082;
  assign n36084 = n36060 & n36081;
  assign n36085 = ~n36072 & n36084;
  assign n36086 = ~n36083 & ~n36085;
  assign n36087 = ~n36074 & n36086;
  assign n36088 = pi3618 & pi9040;
  assign n36089 = pi3634 & ~pi9040;
  assign n36090 = ~n36088 & ~n36089;
  assign n36091 = ~pi0709 & n36090;
  assign n36092 = pi0709 & ~n36090;
  assign n36093 = ~n36091 & ~n36092;
  assign n36094 = pi3633 & pi9040;
  assign n36095 = pi3627 & ~pi9040;
  assign n36096 = ~n36094 & ~n36095;
  assign n36097 = ~pi0718 & n36096;
  assign n36098 = pi0718 & ~n36096;
  assign n36099 = ~n36097 & ~n36098;
  assign n36100 = n36093 & ~n36099;
  assign n36101 = ~n36087 & n36100;
  assign n36102 = n36060 & ~n36081;
  assign n36103 = n36072 & n36102;
  assign n36104 = ~n36099 & n36103;
  assign n36105 = n36066 & n36104;
  assign n36106 = ~n36060 & ~n36072;
  assign n36107 = ~n36060 & ~n36081;
  assign n36108 = n36066 & n36107;
  assign n36109 = ~n36106 & ~n36108;
  assign n36110 = ~n36093 & ~n36109;
  assign n36111 = n36072 & n36084;
  assign n36112 = ~n36093 & n36111;
  assign n36113 = ~n36110 & ~n36112;
  assign n36114 = ~n36099 & ~n36113;
  assign n36115 = ~n36105 & ~n36114;
  assign n36116 = n36066 & ~n36072;
  assign n36117 = ~n36060 & n36116;
  assign n36118 = ~n36066 & n36102;
  assign n36119 = ~n36072 & n36118;
  assign n36120 = ~n36117 & ~n36119;
  assign n36121 = ~n36093 & ~n36120;
  assign n36122 = n36115 & ~n36121;
  assign n36123 = n36066 & n36072;
  assign n36124 = n36060 & n36123;
  assign n36125 = n36081 & n36124;
  assign n36126 = n36066 & n36093;
  assign n36127 = n36107 & n36126;
  assign n36128 = n36072 & n36127;
  assign n36129 = ~n36082 & ~n36102;
  assign n36130 = n36116 & ~n36129;
  assign n36131 = ~n36128 & ~n36130;
  assign n36132 = ~n36125 & n36131;
  assign n36133 = n36073 & ~n36129;
  assign n36134 = ~n36066 & ~n36072;
  assign n36135 = n36060 & n36134;
  assign n36136 = n36081 & n36135;
  assign n36137 = ~n36133 & ~n36136;
  assign n36138 = ~n36066 & ~n36093;
  assign n36139 = n36072 & ~n36081;
  assign n36140 = n36138 & n36139;
  assign n36141 = ~n36066 & n36093;
  assign n36142 = n36107 & n36141;
  assign n36143 = ~n36072 & n36142;
  assign n36144 = ~n36140 & ~n36143;
  assign n36145 = n36137 & n36144;
  assign n36146 = n36132 & n36145;
  assign n36147 = n36099 & ~n36146;
  assign n36148 = n36122 & ~n36147;
  assign n36149 = ~n36101 & n36148;
  assign n36150 = ~pi0759 & ~n36149;
  assign n36151 = pi0759 & n36122;
  assign n36152 = ~n36101 & n36151;
  assign n36153 = ~n36147 & n36152;
  assign po0780 = n36150 | n36153;
  assign n36155 = ~n36072 & n36081;
  assign n36156 = n36093 & n36155;
  assign n36157 = n36066 & n36156;
  assign n36158 = ~n36072 & n36107;
  assign n36159 = ~n36118 & ~n36158;
  assign n36160 = ~n36083 & n36159;
  assign n36161 = n36093 & ~n36160;
  assign n36162 = n36072 & n36107;
  assign n36163 = ~n36072 & n36082;
  assign n36164 = ~n36162 & ~n36163;
  assign n36165 = ~n36093 & ~n36164;
  assign n36166 = ~n36161 & ~n36165;
  assign n36167 = ~n36112 & ~n36119;
  assign n36168 = n36166 & n36167;
  assign n36169 = n36099 & ~n36168;
  assign n36170 = n36066 & n36162;
  assign n36171 = ~n36066 & n36084;
  assign n36172 = n36066 & n36102;
  assign n36173 = ~n36171 & ~n36172;
  assign n36174 = n36093 & ~n36173;
  assign n36175 = ~n36170 & ~n36174;
  assign n36176 = ~n36093 & n36103;
  assign n36177 = n36086 & ~n36176;
  assign n36178 = ~n36158 & n36177;
  assign n36179 = ~n36066 & ~n36178;
  assign n36180 = n36175 & ~n36179;
  assign n36181 = ~n36099 & ~n36180;
  assign n36182 = ~n36169 & ~n36181;
  assign n36183 = ~n36157 & n36182;
  assign n36184 = ~n36072 & n36172;
  assign n36185 = ~n36125 & ~n36184;
  assign n36186 = ~n36093 & ~n36185;
  assign n36187 = n36183 & ~n36186;
  assign n36188 = ~pi0753 & ~n36187;
  assign n36189 = n36182 & ~n36186;
  assign n36190 = pi0753 & n36189;
  assign n36191 = ~n36157 & n36190;
  assign po0781 = n36188 | n36191;
  assign n36193 = pi3641 & pi9040;
  assign n36194 = pi3598 & ~pi9040;
  assign n36195 = ~n36193 & ~n36194;
  assign n36196 = ~pi0703 & ~n36195;
  assign n36197 = pi0703 & n36195;
  assign n36198 = ~n36196 & ~n36197;
  assign n36199 = pi3645 & pi9040;
  assign n36200 = pi3638 & ~pi9040;
  assign n36201 = ~n36199 & ~n36200;
  assign n36202 = ~pi0735 & ~n36201;
  assign n36203 = pi0735 & n36201;
  assign n36204 = ~n36202 & ~n36203;
  assign n36205 = pi3598 & pi9040;
  assign n36206 = pi3645 & ~pi9040;
  assign n36207 = ~n36205 & ~n36206;
  assign n36208 = ~pi0713 & n36207;
  assign n36209 = pi0713 & ~n36207;
  assign n36210 = ~n36208 & ~n36209;
  assign n36211 = ~n36204 & ~n36210;
  assign n36212 = pi3646 & pi9040;
  assign n36213 = pi3643 & ~pi9040;
  assign n36214 = ~n36212 & ~n36213;
  assign n36215 = pi0720 & n36214;
  assign n36216 = ~pi0720 & ~n36214;
  assign n36217 = ~n36215 & ~n36216;
  assign n36218 = pi3610 & pi9040;
  assign n36219 = pi3636 & ~pi9040;
  assign n36220 = ~n36218 & ~n36219;
  assign n36221 = ~pi0729 & n36220;
  assign n36222 = pi0729 & ~n36220;
  assign n36223 = ~n36221 & ~n36222;
  assign n36224 = ~n36217 & n36223;
  assign n36225 = n36211 & n36224;
  assign n36226 = pi3599 & pi9040;
  assign n36227 = pi3631 & ~pi9040;
  assign n36228 = ~n36226 & ~n36227;
  assign n36229 = ~pi0712 & ~n36228;
  assign n36230 = pi0712 & n36228;
  assign n36231 = ~n36229 & ~n36230;
  assign n36232 = n36204 & n36210;
  assign n36233 = n36231 & n36232;
  assign n36234 = n36217 & ~n36231;
  assign n36235 = n36210 & n36234;
  assign n36236 = ~n36204 & n36235;
  assign n36237 = ~n36233 & ~n36236;
  assign n36238 = n36204 & ~n36210;
  assign n36239 = n36217 & n36238;
  assign n36240 = n36237 & ~n36239;
  assign n36241 = n36223 & ~n36240;
  assign n36242 = n36204 & ~n36231;
  assign n36243 = ~n36217 & ~n36223;
  assign n36244 = n36242 & n36243;
  assign n36245 = ~n36231 & n36232;
  assign n36246 = ~n36217 & n36245;
  assign n36247 = ~n36244 & ~n36246;
  assign n36248 = ~n36241 & n36247;
  assign n36249 = ~n36225 & n36248;
  assign n36250 = n36211 & n36231;
  assign n36251 = ~n36217 & n36250;
  assign n36252 = n36231 & n36238;
  assign n36253 = n36217 & n36252;
  assign n36254 = ~n36251 & ~n36253;
  assign n36255 = n36249 & n36254;
  assign n36256 = ~n36198 & ~n36255;
  assign n36257 = n36211 & ~n36231;
  assign n36258 = n36217 & n36257;
  assign n36259 = ~n36204 & n36210;
  assign n36260 = n36231 & n36259;
  assign n36261 = n36217 & n36260;
  assign n36262 = ~n36245 & ~n36261;
  assign n36263 = ~n36258 & n36262;
  assign n36264 = ~n36223 & ~n36263;
  assign n36265 = ~n36204 & n36231;
  assign n36266 = ~n36217 & n36265;
  assign n36267 = n36204 & n36231;
  assign n36268 = n36217 & n36267;
  assign n36269 = ~n36266 & ~n36268;
  assign n36270 = n36223 & ~n36269;
  assign n36271 = ~n36264 & ~n36270;
  assign n36272 = ~n36217 & ~n36231;
  assign n36273 = ~n36210 & n36272;
  assign n36274 = n36204 & n36273;
  assign n36275 = ~n36250 & ~n36274;
  assign n36276 = n36223 & ~n36275;
  assign n36277 = ~n36231 & n36259;
  assign n36278 = ~n36217 & n36277;
  assign n36279 = ~n36258 & ~n36278;
  assign n36280 = n36204 & n36234;
  assign n36281 = ~n36217 & n36252;
  assign n36282 = ~n36280 & ~n36281;
  assign n36283 = ~n36223 & ~n36282;
  assign n36284 = n36279 & ~n36283;
  assign n36285 = ~n36276 & n36284;
  assign n36286 = n36198 & ~n36285;
  assign n36287 = n36210 & ~n36231;
  assign n36288 = ~n36223 & n36287;
  assign n36289 = ~n36217 & n36288;
  assign n36290 = ~n36286 & ~n36289;
  assign n36291 = n36271 & n36290;
  assign n36292 = ~n36256 & n36291;
  assign n36293 = ~pi0738 & ~n36292;
  assign n36294 = pi0738 & n36292;
  assign po0782 = n36293 | n36294;
  assign n36296 = n35920 & n35956;
  assign n36297 = ~n35920 & n35990;
  assign n36298 = ~n36296 & ~n36297;
  assign n36299 = n35947 & ~n36298;
  assign n36300 = ~n35979 & ~n35986;
  assign n36301 = ~n35932 & n35977;
  assign n36302 = ~n35981 & ~n36301;
  assign n36303 = ~n35947 & ~n36302;
  assign n36304 = ~n35920 & ~n35947;
  assign n36305 = n35965 & n36304;
  assign n36306 = n35926 & n36305;
  assign n36307 = ~n35920 & ~n35926;
  assign n36308 = ~n35938 & n36307;
  assign n36309 = n35932 & n36308;
  assign n36310 = n35947 & n35950;
  assign n36311 = ~n36309 & ~n36310;
  assign n36312 = ~n36306 & n36311;
  assign n36313 = ~n36303 & n36312;
  assign n36314 = n36300 & n36313;
  assign n36315 = n35914 & ~n36314;
  assign n36316 = ~n35947 & n35979;
  assign n36317 = n35920 & n35986;
  assign n36318 = ~n36316 & ~n36317;
  assign n36319 = ~n36315 & n36318;
  assign n36320 = ~n36299 & n36319;
  assign n36321 = ~n35926 & ~n35932;
  assign n36322 = n35983 & n36321;
  assign n36323 = ~n35957 & ~n36322;
  assign n36324 = n35947 & n35993;
  assign n36325 = n35920 & n36003;
  assign n36326 = ~n36324 & ~n36325;
  assign n36327 = ~n35920 & n35966;
  assign n36328 = ~n36296 & ~n36327;
  assign n36329 = ~n35920 & n35962;
  assign n36330 = n35926 & ~n35938;
  assign n36331 = ~n36329 & ~n36330;
  assign n36332 = ~n35947 & ~n36331;
  assign n36333 = n36328 & ~n36332;
  assign n36334 = n36326 & n36333;
  assign n36335 = n36323 & n36334;
  assign n36336 = ~n35914 & ~n36335;
  assign n36337 = n36320 & ~n36336;
  assign n36338 = ~pi0743 & ~n36337;
  assign n36339 = pi0743 & n36320;
  assign n36340 = ~n36336 & n36339;
  assign po0783 = n36338 | n36340;
  assign n36342 = ~n35354 & ~n35366;
  assign n36343 = ~n35798 & ~n36342;
  assign n36344 = n35347 & ~n36343;
  assign n36345 = n35354 & n35360;
  assign n36346 = n35375 & n36345;
  assign n36347 = ~n36344 & ~n36346;
  assign n36348 = ~n35347 & n35376;
  assign n36349 = ~n35354 & n36348;
  assign n36350 = ~n35435 & ~n36349;
  assign n36351 = n36347 & n36350;
  assign n36352 = n35341 & ~n36351;
  assign n36353 = ~n35419 & ~n35422;
  assign n36354 = ~n35354 & n35387;
  assign n36355 = n36353 & ~n36354;
  assign n36356 = ~n35347 & ~n36355;
  assign n36357 = n35376 & n35400;
  assign n36358 = ~n35381 & ~n36357;
  assign n36359 = ~n36356 & n36358;
  assign n36360 = ~n35434 & ~n35457;
  assign n36361 = n35347 & ~n36360;
  assign n36362 = n36359 & ~n36361;
  assign n36363 = ~n35341 & ~n36362;
  assign n36364 = ~n36352 & ~n36363;
  assign n36365 = ~n35354 & n35398;
  assign n36366 = n35354 & ~n35454;
  assign n36367 = ~n36365 & ~n36366;
  assign n36368 = n35347 & ~n36367;
  assign n36369 = ~n35419 & n35777;
  assign n36370 = n35424 & ~n36369;
  assign n36371 = ~n36368 & ~n36370;
  assign n36372 = n36364 & n36371;
  assign n36373 = ~pi0741 & ~n36372;
  assign n36374 = pi0741 & n36371;
  assign n36375 = ~n36363 & n36374;
  assign n36376 = ~n36352 & n36375;
  assign po0784 = n36373 | n36376;
  assign n36378 = ~n35503 & n35520;
  assign n36379 = ~n35551 & ~n36378;
  assign n36380 = n35490 & ~n36379;
  assign n36381 = n35510 & n35542;
  assign n36382 = ~n35738 & ~n36381;
  assign n36383 = ~n35490 & ~n36382;
  assign n36384 = ~n35510 & n35537;
  assign n36385 = ~n35759 & ~n36384;
  assign n36386 = ~n35519 & n36385;
  assign n36387 = ~n36383 & n36386;
  assign n36388 = ~n36380 & n36387;
  assign n36389 = ~n35734 & ~n35745;
  assign n36390 = n36388 & n36389;
  assign n36391 = n35529 & ~n36390;
  assign n36392 = n35504 & n35732;
  assign n36393 = n35560 & ~n36392;
  assign n36394 = ~n35490 & ~n36393;
  assign n36395 = ~n35510 & n35548;
  assign n36396 = ~n36394 & ~n36395;
  assign n36397 = n35497 & n35520;
  assign n36398 = n35510 & n35533;
  assign n36399 = ~n36397 & ~n36398;
  assign n36400 = ~n35490 & ~n36399;
  assign n36401 = ~n35490 & n35542;
  assign n36402 = ~n35510 & n36401;
  assign n36403 = ~n36400 & ~n36402;
  assign n36404 = n36396 & n36403;
  assign n36405 = ~n35529 & ~n36404;
  assign n36406 = ~n35537 & ~n35544;
  assign n36407 = ~n35739 & n36406;
  assign n36408 = n35565 & ~n36407;
  assign n36409 = ~n36405 & ~n36408;
  assign n36410 = ~n35519 & ~n35734;
  assign n36411 = n35490 & ~n36410;
  assign n36412 = n36409 & ~n36411;
  assign n36413 = ~n36391 & n36412;
  assign n36414 = ~pi0765 & n36413;
  assign n36415 = pi0765 & ~n36413;
  assign po0785 = n36414 | n36415;
  assign n36417 = ~n36317 & ~n36322;
  assign n36418 = ~n35979 & ~n35990;
  assign n36419 = ~n36329 & n36418;
  assign n36420 = ~n35947 & ~n36419;
  assign n36421 = ~n35938 & n35972;
  assign n36422 = ~n35932 & n36421;
  assign n36423 = ~n36309 & ~n36422;
  assign n36424 = ~n36005 & n36423;
  assign n36425 = n35947 & n35966;
  assign n36426 = n36424 & ~n36425;
  assign n36427 = ~n36420 & n36426;
  assign n36428 = n35914 & ~n36427;
  assign n36429 = n35920 & n35958;
  assign n36430 = n35932 & n35972;
  assign n36431 = ~n35990 & ~n36430;
  assign n36432 = n35947 & ~n36431;
  assign n36433 = ~n36429 & ~n36432;
  assign n36434 = n35948 & n35991;
  assign n36435 = ~n35947 & n35956;
  assign n36436 = ~n36434 & ~n36435;
  assign n36437 = n36433 & n36436;
  assign n36438 = n35932 & n35977;
  assign n36439 = ~n36296 & ~n36438;
  assign n36440 = ~n36327 & n36439;
  assign n36441 = n36437 & n36440;
  assign n36442 = ~n35914 & ~n36441;
  assign n36443 = ~n36296 & n36423;
  assign n36444 = ~n35947 & ~n36443;
  assign n36445 = ~n36442 & ~n36444;
  assign n36446 = ~n36428 & n36445;
  assign n36447 = n36417 & n36446;
  assign n36448 = pi0763 & ~n36447;
  assign n36449 = ~pi0763 & n36447;
  assign po0786 = n36448 | n36449;
  assign n36451 = ~n35266 & n35296;
  assign n36452 = n35266 & n35307;
  assign n36453 = ~n35293 & ~n36452;
  assign n36454 = n35238 & ~n36453;
  assign n36455 = ~n36451 & ~n36454;
  assign n36456 = ~n35238 & ~n35266;
  assign n36457 = ~n35258 & n36456;
  assign n36458 = n35252 & n36457;
  assign n36459 = n35274 & n35308;
  assign n36460 = ~n36458 & ~n36459;
  assign n36461 = ~n35238 & n35317;
  assign n36462 = n36460 & ~n36461;
  assign n36463 = ~n35270 & ~n35282;
  assign n36464 = n35258 & n35272;
  assign n36465 = n36463 & ~n36464;
  assign n36466 = n36462 & n36465;
  assign n36467 = n36455 & n36466;
  assign n36468 = ~n35305 & ~n36467;
  assign n36469 = ~n35245 & n35268;
  assign n36470 = ~n35293 & ~n36469;
  assign n36471 = n35266 & ~n36470;
  assign n36472 = n35252 & n35311;
  assign n36473 = ~n35322 & ~n36472;
  assign n36474 = n35245 & ~n35258;
  assign n36475 = n35266 & n36474;
  assign n36476 = n36473 & ~n36475;
  assign n36477 = n35238 & ~n36476;
  assign n36478 = ~n35266 & n35292;
  assign n36479 = n35252 & n35281;
  assign n36480 = ~n36478 & ~n36479;
  assign n36481 = ~n35238 & ~n36480;
  assign n36482 = ~n35266 & n35275;
  assign n36483 = ~n36481 & ~n36482;
  assign n36484 = ~n36477 & n36483;
  assign n36485 = ~n36471 & n36484;
  assign n36486 = n35305 & ~n36485;
  assign n36487 = n35238 & n35312;
  assign n36488 = ~n36486 & ~n36487;
  assign n36489 = n35287 & n36456;
  assign n36490 = ~n35258 & n36489;
  assign n36491 = n36488 & ~n36490;
  assign n36492 = ~n36468 & n36491;
  assign n36493 = ~pi0744 & ~n36492;
  assign n36494 = pi0744 & n36488;
  assign n36495 = ~n36468 & n36494;
  assign n36496 = ~n36490 & n36495;
  assign po0787 = n36493 | n36496;
  assign n36498 = ~n35601 & n35615;
  assign n36499 = ~n35693 & ~n36498;
  assign n36500 = n35583 & ~n36499;
  assign n36501 = n35611 & n35689;
  assign n36502 = ~n36500 & ~n36501;
  assign n36503 = ~n35662 & n36502;
  assign n36504 = n35601 & ~n35609;
  assign n36505 = n35595 & n36504;
  assign n36506 = n35589 & n36505;
  assign n36507 = ~n35636 & ~n36506;
  assign n36508 = ~n35615 & n36507;
  assign n36509 = n35583 & ~n36508;
  assign n36510 = n35624 & n36509;
  assign n36511 = ~n35583 & n35702;
  assign n36512 = ~n35643 & ~n35660;
  assign n36513 = ~n35634 & n36512;
  assign n36514 = ~n36511 & n36513;
  assign n36515 = n35624 & ~n36514;
  assign n36516 = ~n35583 & ~n35595;
  assign n36517 = n35589 & n36516;
  assign n36518 = n35609 & n36517;
  assign n36519 = ~n35601 & n36518;
  assign n36520 = n35601 & n35670;
  assign n36521 = ~n36518 & ~n36520;
  assign n36522 = ~n35692 & n36521;
  assign n36523 = n35589 & n35641;
  assign n36524 = n35601 & n35629;
  assign n36525 = ~n35610 & ~n36524;
  assign n36526 = n35583 & ~n36525;
  assign n36527 = ~n36523 & ~n36526;
  assign n36528 = n36522 & n36527;
  assign n36529 = ~n35624 & ~n36528;
  assign n36530 = ~n36519 & ~n36529;
  assign n36531 = ~n36515 & n36530;
  assign n36532 = ~n36510 & n36531;
  assign n36533 = n36503 & n36532;
  assign n36534 = pi0755 & ~n36533;
  assign n36535 = ~pi0755 & n36503;
  assign n36536 = n36532 & n36535;
  assign po0788 = n36534 | n36536;
  assign n36538 = ~n36093 & n36162;
  assign n36539 = ~n36066 & n36538;
  assign n36540 = n36084 & n36138;
  assign n36541 = ~n36072 & n36540;
  assign n36542 = ~n36539 & ~n36541;
  assign n36543 = ~n36136 & ~n36143;
  assign n36544 = n36066 & n36081;
  assign n36545 = n36072 & n36544;
  assign n36546 = ~n36108 & ~n36545;
  assign n36547 = ~n36093 & ~n36546;
  assign n36548 = n36093 & ~n36134;
  assign n36549 = ~n36129 & n36548;
  assign n36550 = ~n36072 & ~n36107;
  assign n36551 = ~n36093 & n36550;
  assign n36552 = ~n36066 & n36551;
  assign n36553 = ~n36549 & ~n36552;
  assign n36554 = ~n36547 & n36553;
  assign n36555 = n36543 & n36554;
  assign n36556 = ~n36099 & ~n36555;
  assign n36557 = n36542 & ~n36556;
  assign n36558 = n36083 & n36093;
  assign n36559 = n36066 & n36558;
  assign n36560 = n36093 & n36099;
  assign n36561 = ~n36129 & n36134;
  assign n36562 = ~n36108 & ~n36561;
  assign n36563 = ~n36111 & n36562;
  assign n36564 = n36560 & ~n36563;
  assign n36565 = n36066 & n36085;
  assign n36566 = ~n36072 & n36544;
  assign n36567 = ~n36172 & ~n36566;
  assign n36568 = ~n36066 & n36107;
  assign n36569 = ~n36103 & ~n36568;
  assign n36570 = n36567 & n36569;
  assign n36571 = ~n36093 & ~n36570;
  assign n36572 = ~n36565 & ~n36571;
  assign n36573 = n36099 & ~n36572;
  assign n36574 = ~n36564 & ~n36573;
  assign n36575 = ~n36559 & n36574;
  assign n36576 = n36557 & n36575;
  assign n36577 = pi0761 & ~n36576;
  assign n36578 = ~pi0761 & n36557;
  assign n36579 = n36575 & n36578;
  assign po0790 = n36577 | n36579;
  assign n36581 = ~n36172 & ~n36568;
  assign n36582 = ~n36093 & ~n36581;
  assign n36583 = ~n36541 & ~n36582;
  assign n36584 = ~n36099 & ~n36583;
  assign n36585 = ~n36082 & ~n36155;
  assign n36586 = ~n36066 & ~n36585;
  assign n36587 = ~n36162 & ~n36586;
  assign n36588 = n36093 & ~n36587;
  assign n36589 = ~n36561 & ~n36588;
  assign n36590 = n36066 & n36158;
  assign n36591 = n36060 & n36073;
  assign n36592 = n36066 & ~n36585;
  assign n36593 = ~n36591 & ~n36592;
  assign n36594 = ~n36093 & ~n36593;
  assign n36595 = ~n36590 & ~n36594;
  assign n36596 = n36589 & n36595;
  assign n36597 = n36099 & ~n36596;
  assign n36598 = ~n36082 & n36123;
  assign n36599 = ~n36099 & n36598;
  assign n36600 = n36082 & n36116;
  assign n36601 = ~n36093 & n36600;
  assign n36602 = n36072 & n36126;
  assign n36603 = n36060 & n36602;
  assign n36604 = ~n36601 & ~n36603;
  assign n36605 = ~n36599 & n36604;
  assign n36606 = ~n36103 & ~n36544;
  assign n36607 = n36100 & ~n36606;
  assign n36608 = n36605 & ~n36607;
  assign n36609 = ~n36597 & n36608;
  assign n36610 = ~n36584 & n36609;
  assign n36611 = pi0769 & ~n36610;
  assign n36612 = ~pi0769 & n36610;
  assign po0791 = n36611 | n36612;
  assign n36614 = n35821 & n36014;
  assign n36615 = ~n35872 & ~n35880;
  assign n36616 = ~n35821 & n35841;
  assign n36617 = n35821 & n35892;
  assign n36618 = ~n36616 & ~n36617;
  assign n36619 = n36615 & n36618;
  assign n36620 = ~n35849 & ~n36619;
  assign n36621 = ~n35821 & n35850;
  assign n36622 = ~n35863 & ~n36621;
  assign n36623 = ~n35874 & n36622;
  assign n36624 = n35849 & ~n36623;
  assign n36625 = n35840 & n35881;
  assign n36626 = n35828 & n36625;
  assign n36627 = ~n36624 & ~n36626;
  assign n36628 = ~n36620 & n36627;
  assign n36629 = ~n36614 & n36628;
  assign n36630 = ~n35815 & ~n36629;
  assign n36631 = n35821 & n35842;
  assign n36632 = ~n36028 & ~n36631;
  assign n36633 = ~n35821 & ~n35849;
  assign n36634 = n35851 & n36633;
  assign n36635 = ~n35849 & n35874;
  assign n36636 = ~n35849 & n35884;
  assign n36637 = ~n36635 & ~n36636;
  assign n36638 = n35821 & ~n36637;
  assign n36639 = ~n36634 & ~n36638;
  assign n36640 = ~n35821 & n35871;
  assign n36641 = n35821 & n35850;
  assign n36642 = ~n36640 & ~n36641;
  assign n36643 = ~n35842 & n36642;
  assign n36644 = ~n35872 & n36643;
  assign n36645 = n35849 & ~n36644;
  assign n36646 = n35821 & n35864;
  assign n36647 = ~n36645 & ~n36646;
  assign n36648 = n36639 & n36647;
  assign n36649 = n36632 & n36648;
  assign n36650 = n35815 & ~n36649;
  assign n36651 = ~n35849 & ~n36017;
  assign n36652 = ~n36650 & ~n36651;
  assign n36653 = ~n35875 & ~n36631;
  assign n36654 = n35849 & ~n36653;
  assign n36655 = n36652 & ~n36654;
  assign n36656 = ~n36630 & n36655;
  assign n36657 = pi0754 & ~n36656;
  assign n36658 = ~pi0754 & n36656;
  assign po0792 = n36657 | n36658;
  assign n36660 = ~n35267 & ~n35273;
  assign n36661 = ~n35238 & ~n36660;
  assign n36662 = ~n35329 & ~n36661;
  assign n36663 = ~n35245 & ~n35252;
  assign n36664 = n35238 & n36663;
  assign n36665 = n35266 & n36664;
  assign n36666 = ~n35238 & n35259;
  assign n36667 = n35266 & n36666;
  assign n36668 = ~n36461 & ~n36667;
  assign n36669 = n35245 & ~n35266;
  assign n36670 = n35252 & n36669;
  assign n36671 = n35266 & n35292;
  assign n36672 = ~n36670 & ~n36671;
  assign n36673 = ~n36663 & n36672;
  assign n36674 = n35238 & ~n36673;
  assign n36675 = ~n35276 & ~n36674;
  assign n36676 = n36668 & n36675;
  assign n36677 = ~n35305 & ~n36676;
  assign n36678 = ~n36665 & ~n36677;
  assign n36679 = ~n35293 & ~n35312;
  assign n36680 = ~n35322 & n36679;
  assign n36681 = ~n35238 & ~n36680;
  assign n36682 = ~n35266 & n35317;
  assign n36683 = ~n35296 & ~n36682;
  assign n36684 = n35238 & ~n36683;
  assign n36685 = ~n36681 & ~n36684;
  assign n36686 = ~n36472 & n36685;
  assign n36687 = ~n35282 & ~n35323;
  assign n36688 = n36686 & n36687;
  assign n36689 = n35305 & ~n36688;
  assign n36690 = n36678 & ~n36689;
  assign n36691 = n36662 & n36690;
  assign n36692 = ~pi0758 & ~n36691;
  assign n36693 = pi0758 & n36678;
  assign n36694 = n36662 & n36693;
  assign n36695 = ~n36689 & n36694;
  assign po0793 = n36692 | n36695;
  assign n36697 = n35601 & ~n35714;
  assign n36698 = n35595 & n36697;
  assign n36699 = n35589 & n35691;
  assign n36700 = ~n35672 & ~n36699;
  assign n36701 = ~n35636 & n36700;
  assign n36702 = ~n35583 & ~n36701;
  assign n36703 = ~n35646 & ~n35702;
  assign n36704 = n35583 & ~n36703;
  assign n36705 = ~n36702 & ~n36704;
  assign n36706 = ~n36698 & n36705;
  assign n36707 = ~n35601 & n35611;
  assign n36708 = n36706 & ~n36707;
  assign n36709 = ~n35624 & ~n36708;
  assign n36710 = n35628 & ~n36703;
  assign n36711 = ~n35615 & ~n35647;
  assign n36712 = ~n35611 & ~n35636;
  assign n36713 = n36711 & n36712;
  assign n36714 = n35601 & ~n36713;
  assign n36715 = ~n36710 & ~n36714;
  assign n36716 = ~n35693 & n36715;
  assign n36717 = n35624 & ~n36716;
  assign n36718 = ~n36709 & ~n36717;
  assign n36719 = n35601 & n35702;
  assign n36720 = ~n36707 & ~n36719;
  assign n36721 = n35583 & ~n36720;
  assign n36722 = n36718 & ~n36721;
  assign n36723 = pi0747 & ~n36722;
  assign n36724 = ~pi0747 & ~n36721;
  assign n36725 = ~n36717 & n36724;
  assign n36726 = ~n36709 & n36725;
  assign po0794 = n36723 | n36726;
  assign n36728 = n35490 & n35548;
  assign n36729 = ~n35510 & n35533;
  assign n36730 = ~n35532 & ~n36729;
  assign n36731 = n35490 & ~n36730;
  assign n36732 = ~n35490 & ~n35761;
  assign n36733 = ~n36731 & ~n36732;
  assign n36734 = ~n35749 & n36733;
  assign n36735 = n35529 & ~n36734;
  assign n36736 = ~n36728 & ~n36735;
  assign n36737 = n35517 & n35725;
  assign n36738 = ~n35737 & ~n36737;
  assign n36739 = ~n35497 & ~n36738;
  assign n36740 = ~n35519 & ~n36739;
  assign n36741 = ~n35738 & n36740;
  assign n36742 = ~n35490 & n35534;
  assign n36743 = n35510 & n35551;
  assign n36744 = ~n36742 & ~n36743;
  assign n36745 = n36741 & n36744;
  assign n36746 = ~n35529 & ~n36745;
  assign n36747 = ~n36384 & ~n36398;
  assign n36748 = ~n35490 & ~n36747;
  assign n36749 = ~n36746 & ~n36748;
  assign n36750 = n36736 & n36749;
  assign n36751 = ~pi0768 & ~n36750;
  assign n36752 = ~n36735 & n36749;
  assign n36753 = pi0768 & n36752;
  assign n36754 = ~n36728 & n36753;
  assign po0795 = n36751 | n36754;
  assign n36756 = n36204 & n36235;
  assign n36757 = ~n36267 & ~n36278;
  assign n36758 = ~n36223 & ~n36757;
  assign n36759 = ~n36756 & ~n36758;
  assign n36760 = ~n36274 & n36759;
  assign n36761 = n36217 & n36223;
  assign n36762 = n36257 & n36761;
  assign n36763 = ~n36251 & ~n36762;
  assign n36764 = ~n36261 & n36763;
  assign n36765 = n36760 & n36764;
  assign n36766 = n36198 & ~n36765;
  assign n36767 = ~n36210 & n36234;
  assign n36768 = n36204 & n36767;
  assign n36769 = ~n36236 & ~n36768;
  assign n36770 = ~n36217 & n36260;
  assign n36771 = ~n36246 & ~n36770;
  assign n36772 = ~n36223 & n36257;
  assign n36773 = n36217 & n36250;
  assign n36774 = ~n36772 & ~n36773;
  assign n36775 = ~n36210 & n36231;
  assign n36776 = n36204 & n36217;
  assign n36777 = ~n36775 & ~n36776;
  assign n36778 = ~n36287 & n36777;
  assign n36779 = n36223 & ~n36778;
  assign n36780 = n36774 & ~n36779;
  assign n36781 = n36771 & n36780;
  assign n36782 = n36769 & n36781;
  assign n36783 = ~n36198 & ~n36782;
  assign n36784 = ~n36766 & ~n36783;
  assign n36785 = pi0737 & ~n36784;
  assign n36786 = ~pi0737 & ~n36766;
  assign n36787 = ~n36783 & n36786;
  assign po0796 = n36785 | n36787;
  assign n36789 = ~n35245 & n35252;
  assign n36790 = ~n35238 & n36789;
  assign n36791 = n35266 & n36790;
  assign n36792 = ~n35266 & n36474;
  assign n36793 = ~n35273 & ~n36792;
  assign n36794 = ~n36479 & n36793;
  assign n36795 = ~n36791 & n36794;
  assign n36796 = n35238 & n36469;
  assign n36797 = n36795 & ~n36796;
  assign n36798 = n35305 & ~n36797;
  assign n36799 = ~n35323 & ~n36482;
  assign n36800 = n35238 & ~n36799;
  assign n36801 = ~n35305 & n35307;
  assign n36802 = ~n35238 & n36801;
  assign n36803 = ~n35252 & n36669;
  assign n36804 = ~n36474 & ~n36803;
  assign n36805 = ~n35275 & n36804;
  assign n36806 = n35238 & ~n36805;
  assign n36807 = ~n35245 & n35292;
  assign n36808 = ~n35266 & n36807;
  assign n36809 = ~n36806 & ~n36808;
  assign n36810 = ~n35305 & ~n36809;
  assign n36811 = ~n36802 & ~n36810;
  assign n36812 = ~n36800 & n36811;
  assign n36813 = ~n35266 & n35322;
  assign n36814 = ~n36452 & ~n36813;
  assign n36815 = ~n35270 & ~n35273;
  assign n36816 = n36814 & n36815;
  assign n36817 = ~n35238 & ~n36816;
  assign n36818 = n36812 & ~n36817;
  assign n36819 = ~n36798 & n36818;
  assign n36820 = ~pi0751 & ~n36819;
  assign n36821 = pi0751 & n36812;
  assign n36822 = ~n36798 & n36821;
  assign n36823 = ~n36817 & n36822;
  assign po0797 = n36820 | n36823;
  assign n36825 = ~n35964 & ~n35973;
  assign n36826 = n35914 & ~n36825;
  assign n36827 = n35940 & ~n35947;
  assign n36828 = ~n35978 & ~n36301;
  assign n36829 = ~n35947 & ~n36828;
  assign n36830 = ~n36827 & ~n36829;
  assign n36831 = n35914 & ~n36830;
  assign n36832 = ~n36826 & ~n36831;
  assign n36833 = n35963 & n36304;
  assign n36834 = ~n36306 & ~n36833;
  assign n36835 = ~n35981 & ~n36330;
  assign n36836 = n35947 & ~n36835;
  assign n36837 = n35914 & n36836;
  assign n36838 = n36834 & ~n36837;
  assign n36839 = n35938 & n35977;
  assign n36840 = n35932 & n36839;
  assign n36841 = n35920 & n35965;
  assign n36842 = ~n36297 & ~n36841;
  assign n36843 = n35947 & ~n36842;
  assign n36844 = ~n35979 & ~n36309;
  assign n36845 = n35920 & n35962;
  assign n36846 = ~n36003 & ~n36845;
  assign n36847 = ~n35947 & ~n36846;
  assign n36848 = n36844 & ~n36847;
  assign n36849 = ~n36843 & n36848;
  assign n36850 = ~n36840 & n36849;
  assign n36851 = ~n35914 & ~n36850;
  assign n36852 = ~n36327 & n36423;
  assign n36853 = n35947 & ~n36852;
  assign n36854 = ~n36851 & ~n36853;
  assign n36855 = n36838 & n36854;
  assign n36856 = n36832 & n36855;
  assign n36857 = ~pi0764 & ~n36856;
  assign n36858 = pi0764 & n36838;
  assign n36859 = n36832 & n36858;
  assign n36860 = n36854 & n36859;
  assign po0798 = n36857 | n36860;
  assign n36862 = ~n36020 & ~n36631;
  assign n36863 = ~n36626 & n36862;
  assign n36864 = ~n35849 & ~n36863;
  assign n36865 = ~n36031 & ~n36047;
  assign n36866 = ~n36028 & ~n36636;
  assign n36867 = ~n36014 & ~n36641;
  assign n36868 = n35849 & ~n36867;
  assign n36869 = ~n35880 & ~n36868;
  assign n36870 = n36866 & n36869;
  assign n36871 = n35815 & ~n36870;
  assign n36872 = ~n35834 & n35840;
  assign n36873 = ~n35852 & ~n36872;
  assign n36874 = ~n35821 & ~n36873;
  assign n36875 = ~n35842 & ~n36034;
  assign n36876 = n35849 & ~n36875;
  assign n36877 = ~n35821 & n35840;
  assign n36878 = ~n35864 & ~n36877;
  assign n36879 = ~n35855 & n36878;
  assign n36880 = ~n35849 & ~n36879;
  assign n36881 = ~n36876 & ~n36880;
  assign n36882 = ~n36874 & n36881;
  assign n36883 = ~n35815 & ~n36882;
  assign n36884 = ~n36871 & ~n36883;
  assign n36885 = n36865 & n36884;
  assign n36886 = ~n36864 & n36885;
  assign n36887 = ~pi0770 & ~n36886;
  assign n36888 = pi0770 & n36865;
  assign n36889 = ~n36864 & n36888;
  assign n36890 = n36884 & n36889;
  assign po0799 = n36887 | n36890;
  assign n36892 = ~n36217 & n36238;
  assign n36893 = ~n36770 & ~n36892;
  assign n36894 = ~n36223 & n36893;
  assign n36895 = ~n36211 & ~n36232;
  assign n36896 = n36231 & ~n36895;
  assign n36897 = n36217 & n36265;
  assign n36898 = ~n36204 & n36272;
  assign n36899 = n36217 & n36232;
  assign n36900 = ~n36898 & ~n36899;
  assign n36901 = ~n36897 & n36900;
  assign n36902 = ~n36896 & n36901;
  assign n36903 = n36223 & n36902;
  assign n36904 = ~n36894 & ~n36903;
  assign n36905 = n36217 & n36896;
  assign n36906 = ~n36768 & ~n36905;
  assign n36907 = ~n36904 & n36906;
  assign n36908 = n36198 & ~n36907;
  assign n36909 = ~n36223 & ~n36895;
  assign n36910 = ~n36217 & n36909;
  assign n36911 = n36217 & n36259;
  assign n36912 = ~n36253 & ~n36911;
  assign n36913 = ~n36223 & ~n36912;
  assign n36914 = ~n36231 & n36909;
  assign n36915 = ~n36913 & ~n36914;
  assign n36916 = ~n36910 & n36915;
  assign n36917 = ~n36198 & ~n36916;
  assign n36918 = ~n36908 & ~n36917;
  assign n36919 = ~n36223 & n36236;
  assign n36920 = n36223 & ~n36906;
  assign n36921 = ~n36919 & ~n36920;
  assign n36922 = n36223 & ~n36893;
  assign n36923 = ~n36236 & ~n36922;
  assign n36924 = ~n36198 & ~n36923;
  assign n36925 = n36921 & ~n36924;
  assign n36926 = n36918 & n36925;
  assign n36927 = pi0760 & ~n36926;
  assign n36928 = ~pi0760 & n36925;
  assign n36929 = ~n36917 & n36928;
  assign n36930 = ~n36908 & n36929;
  assign po0800 = n36927 | n36930;
  assign n36932 = ~n36223 & n36258;
  assign n36933 = n36272 & ~n36895;
  assign n36934 = ~n36260 & ~n36933;
  assign n36935 = ~n36768 & n36934;
  assign n36936 = n36223 & ~n36935;
  assign n36937 = n36217 & n36233;
  assign n36938 = ~n36936 & ~n36937;
  assign n36939 = ~n36217 & n36775;
  assign n36940 = ~n36277 & ~n36939;
  assign n36941 = ~n36899 & n36940;
  assign n36942 = ~n36223 & ~n36941;
  assign n36943 = n36938 & ~n36942;
  assign n36944 = n36198 & ~n36943;
  assign n36945 = ~n36932 & ~n36944;
  assign n36946 = ~n36217 & n36232;
  assign n36947 = ~n36231 & n36238;
  assign n36948 = ~n36946 & ~n36947;
  assign n36949 = ~n36223 & ~n36948;
  assign n36950 = ~n36261 & ~n36949;
  assign n36951 = n36217 & n36287;
  assign n36952 = ~n36775 & ~n36951;
  assign n36953 = ~n36277 & n36952;
  assign n36954 = n36223 & ~n36953;
  assign n36955 = ~n36253 & ~n36258;
  assign n36956 = ~n36217 & n36233;
  assign n36957 = n36955 & ~n36956;
  assign n36958 = ~n36954 & n36957;
  assign n36959 = n36950 & n36958;
  assign n36960 = ~n36198 & ~n36959;
  assign n36961 = ~n36281 & ~n36897;
  assign n36962 = n36223 & ~n36961;
  assign n36963 = ~n36960 & ~n36962;
  assign n36964 = n36945 & n36963;
  assign n36965 = pi0767 & n36964;
  assign n36966 = ~pi0767 & ~n36964;
  assign po0801 = n36965 | n36966;
  assign n36968 = pi3677 & pi9040;
  assign n36969 = pi3682 & ~pi9040;
  assign n36970 = ~n36968 & ~n36969;
  assign n36971 = pi0771 & n36970;
  assign n36972 = ~pi0771 & ~n36970;
  assign n36973 = ~n36971 & ~n36972;
  assign n36974 = pi3672 & pi9040;
  assign n36975 = pi3702 & ~pi9040;
  assign n36976 = ~n36974 & ~n36975;
  assign n36977 = pi0798 & n36976;
  assign n36978 = ~pi0798 & ~n36976;
  assign n36979 = ~n36977 & ~n36978;
  assign n36980 = pi3701 & pi9040;
  assign n36981 = pi3668 & ~pi9040;
  assign n36982 = ~n36980 & ~n36981;
  assign n36983 = ~pi0766 & ~n36982;
  assign n36984 = pi0766 & n36982;
  assign n36985 = ~n36983 & ~n36984;
  assign n36986 = pi3657 & pi9040;
  assign n36987 = pi3658 & ~pi9040;
  assign n36988 = ~n36986 & ~n36987;
  assign n36989 = ~pi0795 & ~n36988;
  assign n36990 = pi0795 & ~n36986;
  assign n36991 = ~n36987 & n36990;
  assign n36992 = ~n36989 & ~n36991;
  assign n36993 = pi3690 & pi9040;
  assign n36994 = pi3684 & ~pi9040;
  assign n36995 = ~n36993 & ~n36994;
  assign n36996 = ~pi0774 & n36995;
  assign n36997 = pi0774 & ~n36995;
  assign n36998 = ~n36996 & ~n36997;
  assign n36999 = ~n36992 & n36998;
  assign n37000 = n36985 & n36999;
  assign n37001 = n36979 & n37000;
  assign n37002 = n36992 & n36998;
  assign n37003 = ~n36985 & n37002;
  assign n37004 = n36979 & n37003;
  assign n37005 = ~n37001 & ~n37004;
  assign n37006 = n36992 & ~n36998;
  assign n37007 = ~n36985 & n37006;
  assign n37008 = ~n36979 & n37007;
  assign n37009 = ~n36985 & n36999;
  assign n37010 = ~n36979 & n37009;
  assign n37011 = ~n37008 & ~n37010;
  assign n37012 = n37005 & n37011;
  assign n37013 = n36973 & ~n37012;
  assign n37014 = n36979 & ~n36985;
  assign n37015 = ~n36998 & n37014;
  assign n37016 = ~n36992 & n37015;
  assign n37017 = ~n37003 & ~n37016;
  assign n37018 = n36973 & ~n37017;
  assign n37019 = ~n36979 & ~n36998;
  assign n37020 = ~n36973 & n37019;
  assign n37021 = n36985 & n36992;
  assign n37022 = n36979 & n36999;
  assign n37023 = ~n37021 & ~n37022;
  assign n37024 = ~n36973 & ~n37023;
  assign n37025 = ~n37020 & ~n37024;
  assign n37026 = ~n36992 & ~n36998;
  assign n37027 = n36985 & n37026;
  assign n37028 = ~n36979 & n37027;
  assign n37029 = n37025 & ~n37028;
  assign n37030 = ~n36998 & n37021;
  assign n37031 = n36979 & n37030;
  assign n37032 = n37029 & ~n37031;
  assign n37033 = ~n37018 & n37032;
  assign n37034 = ~pi3705 & ~pi9040;
  assign n37035 = ~pi3668 & pi9040;
  assign n37036 = ~n37034 & ~n37035;
  assign n37037 = ~pi0796 & n37036;
  assign n37038 = pi0796 & ~n37036;
  assign n37039 = ~n37037 & ~n37038;
  assign n37040 = ~n37033 & ~n37039;
  assign n37041 = ~n36985 & ~n36998;
  assign n37042 = ~n36973 & n36979;
  assign n37043 = n37039 & n37042;
  assign n37044 = n37041 & n37043;
  assign n37045 = ~n36979 & ~n36985;
  assign n37046 = n36998 & n37045;
  assign n37047 = ~n36973 & ~n37046;
  assign n37048 = n36979 & n36985;
  assign n37049 = ~n36992 & n37048;
  assign n37050 = ~n37006 & ~n37041;
  assign n37051 = ~n36979 & ~n37050;
  assign n37052 = ~n37000 & ~n37051;
  assign n37053 = n36973 & n37052;
  assign n37054 = ~n37049 & n37053;
  assign n37055 = ~n37047 & ~n37054;
  assign n37056 = n36985 & n37002;
  assign n37057 = n36979 & n37056;
  assign n37058 = ~n37055 & ~n37057;
  assign n37059 = n37039 & ~n37058;
  assign n37060 = ~n37044 & ~n37059;
  assign n37061 = ~n37040 & n37060;
  assign n37062 = ~n37013 & n37061;
  assign n37063 = ~n36973 & n37028;
  assign n37064 = n37062 & ~n37063;
  assign n37065 = pi0800 & ~n37064;
  assign n37066 = n37061 & ~n37063;
  assign n37067 = ~pi0800 & n37066;
  assign n37068 = ~n37013 & n37067;
  assign po0821 = n37065 | n37068;
  assign n37070 = pi3660 & pi9040;
  assign n37071 = pi3656 & ~pi9040;
  assign n37072 = ~n37070 & ~n37071;
  assign n37073 = ~pi0790 & n37072;
  assign n37074 = pi0790 & ~n37072;
  assign n37075 = ~n37073 & ~n37074;
  assign n37076 = pi3752 & pi9040;
  assign n37077 = pi3692 & ~pi9040;
  assign n37078 = ~n37076 & ~n37077;
  assign n37079 = ~pi0781 & ~n37078;
  assign n37080 = pi0781 & ~n37076;
  assign n37081 = ~n37077 & n37080;
  assign n37082 = ~n37079 & ~n37081;
  assign n37083 = pi3696 & pi9040;
  assign n37084 = pi3686 & ~pi9040;
  assign n37085 = ~n37083 & ~n37084;
  assign n37086 = pi0791 & n37085;
  assign n37087 = ~pi0791 & ~n37085;
  assign n37088 = ~n37086 & ~n37087;
  assign n37089 = n37082 & ~n37088;
  assign n37090 = pi3678 & pi9040;
  assign n37091 = pi3669 & ~pi9040;
  assign n37092 = ~n37090 & ~n37091;
  assign n37093 = pi0789 & n37092;
  assign n37094 = ~pi0789 & ~n37092;
  assign n37095 = ~n37093 & ~n37094;
  assign n37096 = pi3673 & pi9040;
  assign n37097 = pi3678 & ~pi9040;
  assign n37098 = ~n37096 & ~n37097;
  assign n37099 = ~pi0745 & ~n37098;
  assign n37100 = pi0745 & ~n37096;
  assign n37101 = ~n37097 & n37100;
  assign n37102 = ~n37099 & ~n37101;
  assign n37103 = n37095 & n37102;
  assign n37104 = n37089 & n37103;
  assign n37105 = n37095 & ~n37102;
  assign n37106 = ~n37082 & n37105;
  assign n37107 = ~n37104 & ~n37106;
  assign n37108 = n37075 & ~n37107;
  assign n37109 = pi3661 & ~pi9040;
  assign n37110 = pi3656 & pi9040;
  assign n37111 = ~n37109 & ~n37110;
  assign n37112 = ~pi0782 & ~n37111;
  assign n37113 = pi0782 & n37111;
  assign n37114 = ~n37112 & ~n37113;
  assign n37115 = ~n37075 & ~n37095;
  assign n37116 = n37082 & n37115;
  assign n37117 = n37089 & ~n37102;
  assign n37118 = n37082 & n37088;
  assign n37119 = n37102 & n37118;
  assign n37120 = ~n37117 & ~n37119;
  assign n37121 = ~n37082 & ~n37088;
  assign n37122 = n37102 & n37121;
  assign n37123 = n37095 & n37122;
  assign n37124 = n37120 & ~n37123;
  assign n37125 = ~n37075 & ~n37124;
  assign n37126 = ~n37116 & ~n37125;
  assign n37127 = ~n37082 & n37088;
  assign n37128 = ~n37102 & n37127;
  assign n37129 = n37095 & n37128;
  assign n37130 = n37126 & ~n37129;
  assign n37131 = ~n37095 & n37121;
  assign n37132 = ~n37082 & n37102;
  assign n37133 = n37088 & n37132;
  assign n37134 = ~n37131 & ~n37133;
  assign n37135 = n37075 & ~n37134;
  assign n37136 = ~n37102 & n37118;
  assign n37137 = ~n37095 & n37136;
  assign n37138 = ~n37135 & ~n37137;
  assign n37139 = n37130 & n37138;
  assign n37140 = n37114 & ~n37139;
  assign n37141 = ~n37108 & ~n37140;
  assign n37142 = ~n37075 & ~n37114;
  assign n37143 = ~n37134 & n37142;
  assign n37144 = ~n37102 & n37121;
  assign n37145 = ~n37136 & ~n37144;
  assign n37146 = n37095 & ~n37145;
  assign n37147 = ~n37104 & ~n37146;
  assign n37148 = ~n37114 & ~n37147;
  assign n37149 = ~n37143 & ~n37148;
  assign n37150 = n37075 & ~n37114;
  assign n37151 = n37089 & ~n37095;
  assign n37152 = ~n37128 & ~n37151;
  assign n37153 = n37082 & n37102;
  assign n37154 = n37152 & ~n37153;
  assign n37155 = n37150 & ~n37154;
  assign n37156 = n37149 & ~n37155;
  assign n37157 = n37141 & n37156;
  assign n37158 = ~pi0804 & ~n37157;
  assign n37159 = pi0804 & n37149;
  assign n37160 = n37141 & n37159;
  assign n37161 = ~n37155 & n37160;
  assign po0833 = n37158 | n37161;
  assign n37163 = pi3755 & pi9040;
  assign n37164 = pi3662 & ~pi9040;
  assign n37165 = ~n37163 & ~n37164;
  assign n37166 = ~pi0781 & ~n37165;
  assign n37167 = pi0781 & n37165;
  assign n37168 = ~n37166 & ~n37167;
  assign n37169 = pi3680 & pi9040;
  assign n37170 = pi3665 & ~pi9040;
  assign n37171 = ~n37169 & ~n37170;
  assign n37172 = ~pi0795 & n37171;
  assign n37173 = pi0795 & ~n37171;
  assign n37174 = ~n37172 & ~n37173;
  assign n37175 = pi3697 & pi9040;
  assign n37176 = pi3755 & ~pi9040;
  assign n37177 = ~n37175 & ~n37176;
  assign n37178 = ~pi0796 & n37177;
  assign n37179 = pi0796 & ~n37177;
  assign n37180 = ~n37178 & ~n37179;
  assign n37181 = pi3703 & pi9040;
  assign n37182 = pi3683 & ~pi9040;
  assign n37183 = ~n37181 & ~n37182;
  assign n37184 = ~pi0745 & n37183;
  assign n37185 = pi0745 & ~n37183;
  assign n37186 = ~n37184 & ~n37185;
  assign n37187 = n37180 & ~n37186;
  assign n37188 = pi3708 & pi9040;
  assign n37189 = pi3679 & ~pi9040;
  assign n37190 = ~n37188 & ~n37189;
  assign n37191 = pi0779 & n37190;
  assign n37192 = ~pi0779 & ~n37190;
  assign n37193 = ~n37191 & ~n37192;
  assign n37194 = pi3699 & pi9040;
  assign n37195 = pi3708 & ~pi9040;
  assign n37196 = ~n37194 & ~n37195;
  assign n37197 = ~pi0799 & n37196;
  assign n37198 = pi0799 & ~n37196;
  assign n37199 = ~n37197 & ~n37198;
  assign n37200 = n37193 & ~n37199;
  assign n37201 = n37187 & n37200;
  assign n37202 = ~n37174 & n37201;
  assign n37203 = ~n37193 & ~n37199;
  assign n37204 = ~n37180 & ~n37186;
  assign n37205 = n37203 & n37204;
  assign n37206 = n37180 & n37186;
  assign n37207 = ~n37174 & n37206;
  assign n37208 = ~n37193 & n37207;
  assign n37209 = ~n37180 & n37186;
  assign n37210 = ~n37174 & n37209;
  assign n37211 = ~n37199 & n37210;
  assign n37212 = n37193 & n37211;
  assign n37213 = ~n37208 & ~n37212;
  assign n37214 = ~n37205 & n37213;
  assign n37215 = ~n37202 & n37214;
  assign n37216 = n37174 & ~n37193;
  assign n37217 = ~n37186 & n37216;
  assign n37218 = ~n37180 & n37217;
  assign n37219 = n37215 & ~n37218;
  assign n37220 = ~n37168 & ~n37219;
  assign n37221 = ~n37174 & ~n37193;
  assign n37222 = n37186 & n37221;
  assign n37223 = ~n37174 & ~n37180;
  assign n37224 = ~n37186 & n37223;
  assign n37225 = n37193 & n37224;
  assign n37226 = ~n37222 & ~n37225;
  assign n37227 = n37174 & n37187;
  assign n37228 = n37193 & n37227;
  assign n37229 = n37226 & ~n37228;
  assign n37230 = n37199 & ~n37229;
  assign n37231 = n37174 & n37186;
  assign n37232 = ~n37180 & n37231;
  assign n37233 = n37199 & n37232;
  assign n37234 = n37193 & n37233;
  assign n37235 = n37180 & n37221;
  assign n37236 = ~n37193 & n37206;
  assign n37237 = ~n37235 & ~n37236;
  assign n37238 = n37199 & ~n37237;
  assign n37239 = ~n37234 & ~n37238;
  assign n37240 = ~n37168 & ~n37239;
  assign n37241 = ~n37230 & ~n37240;
  assign n37242 = ~n37220 & n37241;
  assign n37243 = n37174 & n37193;
  assign n37244 = ~n37199 & n37243;
  assign n37245 = n37206 & n37244;
  assign n37246 = n37174 & ~n37180;
  assign n37247 = n37203 & n37246;
  assign n37248 = n37199 & n37223;
  assign n37249 = n37180 & n37193;
  assign n37250 = n37174 & n37249;
  assign n37251 = ~n37227 & ~n37250;
  assign n37252 = ~n37248 & n37251;
  assign n37253 = ~n37193 & n37232;
  assign n37254 = n37252 & ~n37253;
  assign n37255 = n37174 & ~n37186;
  assign n37256 = n37193 & n37206;
  assign n37257 = ~n37255 & ~n37256;
  assign n37258 = ~n37199 & ~n37257;
  assign n37259 = n37187 & ~n37199;
  assign n37260 = ~n37193 & n37259;
  assign n37261 = ~n37258 & ~n37260;
  assign n37262 = n37254 & n37261;
  assign n37263 = n37168 & ~n37262;
  assign n37264 = ~n37247 & ~n37263;
  assign n37265 = ~n37245 & n37264;
  assign n37266 = n37242 & n37265;
  assign n37267 = pi0811 & n37266;
  assign n37268 = ~pi0811 & ~n37266;
  assign po0834 = n37267 | n37268;
  assign n37270 = ~n37174 & n37180;
  assign n37271 = ~n37218 & ~n37270;
  assign n37272 = ~n37249 & n37271;
  assign n37273 = ~n37199 & ~n37272;
  assign n37274 = n37193 & n37199;
  assign n37275 = ~n37180 & n37274;
  assign n37276 = ~n37174 & n37193;
  assign n37277 = ~n37186 & n37276;
  assign n37278 = ~n37193 & n37210;
  assign n37279 = ~n37277 & ~n37278;
  assign n37280 = n37174 & n37180;
  assign n37281 = ~n37193 & n37199;
  assign n37282 = n37280 & n37281;
  assign n37283 = n37279 & ~n37282;
  assign n37284 = ~n37275 & n37283;
  assign n37285 = ~n37273 & n37284;
  assign n37286 = n37168 & ~n37285;
  assign n37287 = ~n37174 & n37187;
  assign n37288 = ~n37193 & n37287;
  assign n37289 = n37193 & n37207;
  assign n37290 = ~n37288 & ~n37289;
  assign n37291 = ~n37199 & ~n37290;
  assign n37292 = ~n37286 & ~n37291;
  assign n37293 = n37193 & n37210;
  assign n37294 = ~n37224 & ~n37232;
  assign n37295 = ~n37199 & ~n37294;
  assign n37296 = ~n37293 & ~n37295;
  assign n37297 = ~n37228 & n37296;
  assign n37298 = ~n37168 & ~n37297;
  assign n37299 = ~n37204 & ~n37206;
  assign n37300 = n37174 & ~n37299;
  assign n37301 = ~n37236 & ~n37300;
  assign n37302 = n37199 & ~n37301;
  assign n37303 = ~n37168 & n37302;
  assign n37304 = ~n37298 & ~n37303;
  assign n37305 = n37292 & n37304;
  assign n37306 = pi0818 & ~n37305;
  assign n37307 = ~pi0818 & n37292;
  assign n37308 = n37304 & n37307;
  assign po0835 = n37306 | n37308;
  assign n37310 = n37075 & n37095;
  assign n37311 = ~n37121 & ~n37136;
  assign n37312 = n37310 & ~n37311;
  assign n37313 = n37075 & ~n37102;
  assign n37314 = n37121 & n37313;
  assign n37315 = ~n37312 & ~n37314;
  assign n37316 = n37114 & ~n37315;
  assign n37317 = ~n37095 & n37102;
  assign n37318 = n37088 & n37317;
  assign n37319 = n37082 & n37318;
  assign n37320 = ~n37153 & ~n37317;
  assign n37321 = ~n37075 & ~n37320;
  assign n37322 = ~n37095 & ~n37102;
  assign n37323 = ~n37088 & n37322;
  assign n37324 = n37082 & n37323;
  assign n37325 = ~n37321 & ~n37324;
  assign n37326 = ~n37319 & n37325;
  assign n37327 = n37114 & ~n37326;
  assign n37328 = ~n37316 & ~n37327;
  assign n37329 = n37088 & n37103;
  assign n37330 = ~n37082 & n37329;
  assign n37331 = ~n37095 & n37128;
  assign n37332 = ~n37330 & ~n37331;
  assign n37333 = n37075 & ~n37332;
  assign n37334 = n37095 & n37144;
  assign n37335 = ~n37095 & n37153;
  assign n37336 = ~n37334 & ~n37335;
  assign n37337 = ~n37075 & ~n37336;
  assign n37338 = ~n37089 & ~n37153;
  assign n37339 = n37095 & ~n37338;
  assign n37340 = ~n37128 & ~n37339;
  assign n37341 = n37075 & ~n37340;
  assign n37342 = n37088 & ~n37095;
  assign n37343 = n37075 & n37342;
  assign n37344 = ~n37102 & n37343;
  assign n37345 = ~n37088 & n37102;
  assign n37346 = ~n37128 & ~n37345;
  assign n37347 = ~n37095 & ~n37346;
  assign n37348 = ~n37075 & n37095;
  assign n37349 = n37118 & n37348;
  assign n37350 = ~n37102 & n37349;
  assign n37351 = ~n37347 & ~n37350;
  assign n37352 = ~n37344 & n37351;
  assign n37353 = ~n37341 & n37352;
  assign n37354 = ~n37330 & n37353;
  assign n37355 = ~n37114 & ~n37354;
  assign n37356 = ~n37337 & ~n37355;
  assign n37357 = ~n37333 & n37356;
  assign n37358 = n37328 & n37357;
  assign n37359 = pi0813 & n37358;
  assign n37360 = ~pi0813 & ~n37358;
  assign po0836 = n37359 | n37360;
  assign n37362 = ~pi3689 & pi9040;
  assign n37363 = pi3675 & ~pi9040;
  assign n37364 = ~n37362 & ~n37363;
  assign n37365 = ~pi0774 & ~n37364;
  assign n37366 = pi0774 & n37364;
  assign n37367 = ~n37365 & ~n37366;
  assign n37368 = pi3705 & pi9040;
  assign n37369 = pi3664 & ~pi9040;
  assign n37370 = ~n37368 & ~n37369;
  assign n37371 = ~pi0792 & n37370;
  assign n37372 = pi0792 & ~n37370;
  assign n37373 = ~n37371 & ~n37372;
  assign n37374 = pi3670 & pi9040;
  assign n37375 = pi3663 & ~pi9040;
  assign n37376 = ~n37374 & ~n37375;
  assign n37377 = ~pi0766 & n37376;
  assign n37378 = pi0766 & ~n37376;
  assign n37379 = ~n37377 & ~n37378;
  assign n37380 = n37373 & ~n37379;
  assign n37381 = pi3695 & pi9040;
  assign n37382 = pi3671 & ~pi9040;
  assign n37383 = ~n37381 & ~n37382;
  assign n37384 = ~pi0787 & n37383;
  assign n37385 = pi0787 & ~n37383;
  assign n37386 = ~n37384 & ~n37385;
  assign n37387 = pi3706 & pi9040;
  assign n37388 = pi3681 & ~pi9040;
  assign n37389 = ~n37387 & ~n37388;
  assign n37390 = ~pi0788 & n37389;
  assign n37391 = pi0788 & ~n37389;
  assign n37392 = ~n37390 & ~n37391;
  assign n37393 = n37386 & n37392;
  assign n37394 = n37380 & n37393;
  assign n37395 = pi3675 & pi9040;
  assign n37396 = pi3677 & ~pi9040;
  assign n37397 = ~n37395 & ~n37396;
  assign n37398 = ~pi0786 & ~n37397;
  assign n37399 = pi0786 & ~n37395;
  assign n37400 = ~n37396 & n37399;
  assign n37401 = ~n37398 & ~n37400;
  assign n37402 = ~n37373 & n37379;
  assign n37403 = n37401 & n37402;
  assign n37404 = ~n37386 & ~n37401;
  assign n37405 = n37379 & n37404;
  assign n37406 = n37373 & n37405;
  assign n37407 = ~n37403 & ~n37406;
  assign n37408 = ~n37373 & ~n37379;
  assign n37409 = ~n37386 & n37408;
  assign n37410 = n37407 & ~n37409;
  assign n37411 = n37392 & ~n37410;
  assign n37412 = ~n37373 & ~n37401;
  assign n37413 = n37386 & ~n37392;
  assign n37414 = n37412 & n37413;
  assign n37415 = ~n37401 & n37402;
  assign n37416 = n37386 & n37415;
  assign n37417 = ~n37414 & ~n37416;
  assign n37418 = ~n37411 & n37417;
  assign n37419 = ~n37394 & n37418;
  assign n37420 = n37380 & n37401;
  assign n37421 = n37386 & n37420;
  assign n37422 = ~n37379 & n37401;
  assign n37423 = ~n37386 & n37422;
  assign n37424 = ~n37373 & n37423;
  assign n37425 = ~n37421 & ~n37424;
  assign n37426 = n37419 & n37425;
  assign n37427 = ~n37367 & ~n37426;
  assign n37428 = ~n37379 & ~n37401;
  assign n37429 = n37386 & n37428;
  assign n37430 = ~n37373 & n37429;
  assign n37431 = ~n37420 & ~n37430;
  assign n37432 = n37392 & ~n37431;
  assign n37433 = n37380 & ~n37401;
  assign n37434 = ~n37386 & n37433;
  assign n37435 = n37379 & ~n37401;
  assign n37436 = n37386 & n37435;
  assign n37437 = n37373 & n37436;
  assign n37438 = ~n37434 & ~n37437;
  assign n37439 = ~n37373 & n37404;
  assign n37440 = n37401 & n37408;
  assign n37441 = n37386 & n37440;
  assign n37442 = ~n37439 & ~n37441;
  assign n37443 = ~n37392 & ~n37442;
  assign n37444 = n37438 & ~n37443;
  assign n37445 = ~n37432 & n37444;
  assign n37446 = n37367 & ~n37445;
  assign n37447 = n37373 & n37379;
  assign n37448 = n37401 & n37447;
  assign n37449 = ~n37386 & n37448;
  assign n37450 = ~n37415 & ~n37449;
  assign n37451 = ~n37434 & n37450;
  assign n37452 = ~n37392 & ~n37451;
  assign n37453 = n37373 & n37401;
  assign n37454 = n37386 & n37453;
  assign n37455 = ~n37373 & n37401;
  assign n37456 = ~n37386 & n37455;
  assign n37457 = ~n37454 & ~n37456;
  assign n37458 = n37392 & ~n37457;
  assign n37459 = ~n37452 & ~n37458;
  assign n37460 = ~n37392 & n37435;
  assign n37461 = n37386 & n37460;
  assign n37462 = n37459 & ~n37461;
  assign n37463 = ~n37446 & n37462;
  assign n37464 = ~n37427 & n37463;
  assign n37465 = ~pi0805 & ~n37464;
  assign n37466 = pi0805 & n37464;
  assign po0838 = n37465 | n37466;
  assign n37468 = pi3685 & ~pi9040;
  assign n37469 = pi3684 & pi9040;
  assign n37470 = ~n37468 & ~n37469;
  assign n37471 = ~pi0792 & ~n37470;
  assign n37472 = pi0792 & n37470;
  assign n37473 = ~n37471 & ~n37472;
  assign n37474 = pi3674 & pi9040;
  assign n37475 = pi3657 & ~pi9040;
  assign n37476 = ~n37474 & ~n37475;
  assign n37477 = ~pi0785 & n37476;
  assign n37478 = pi0785 & ~n37476;
  assign n37479 = ~n37477 & ~n37478;
  assign n37480 = pi3682 & pi9040;
  assign n37481 = pi3676 & ~pi9040;
  assign n37482 = ~n37480 & ~n37481;
  assign n37483 = ~pi0762 & ~n37482;
  assign n37484 = pi0762 & ~n37480;
  assign n37485 = ~n37481 & n37484;
  assign n37486 = ~n37483 & ~n37485;
  assign n37487 = pi3663 & pi9040;
  assign n37488 = pi3655 & ~pi9040;
  assign n37489 = ~n37487 & ~n37488;
  assign n37490 = pi0773 & n37489;
  assign n37491 = ~pi0773 & ~n37489;
  assign n37492 = ~n37490 & ~n37491;
  assign n37493 = pi3704 & pi9040;
  assign n37494 = pi3674 & ~pi9040;
  assign n37495 = ~n37493 & ~n37494;
  assign n37496 = ~pi0778 & ~n37495;
  assign n37497 = pi0778 & n37495;
  assign n37498 = ~n37496 & ~n37497;
  assign n37499 = n37492 & ~n37498;
  assign n37500 = n37486 & n37499;
  assign n37501 = pi3685 & pi9040;
  assign n37502 = pi3707 & ~pi9040;
  assign n37503 = ~n37501 & ~n37502;
  assign n37504 = ~pi0786 & ~n37503;
  assign n37505 = pi0786 & ~n37501;
  assign n37506 = ~n37502 & n37505;
  assign n37507 = ~n37504 & ~n37506;
  assign n37508 = n37498 & n37507;
  assign n37509 = n37492 & n37508;
  assign n37510 = ~n37500 & ~n37509;
  assign n37511 = n37498 & ~n37507;
  assign n37512 = ~n37492 & n37511;
  assign n37513 = ~n37486 & n37512;
  assign n37514 = n37510 & ~n37513;
  assign n37515 = ~n37479 & ~n37514;
  assign n37516 = ~n37492 & n37498;
  assign n37517 = ~n37486 & n37507;
  assign n37518 = n37516 & n37517;
  assign n37519 = ~n37498 & n37507;
  assign n37520 = n37492 & n37519;
  assign n37521 = ~n37486 & n37520;
  assign n37522 = ~n37492 & ~n37498;
  assign n37523 = ~n37511 & ~n37522;
  assign n37524 = n37486 & ~n37523;
  assign n37525 = ~n37521 & ~n37524;
  assign n37526 = ~n37518 & n37525;
  assign n37527 = n37479 & ~n37526;
  assign n37528 = ~n37515 & ~n37527;
  assign n37529 = n37473 & ~n37528;
  assign n37530 = ~n37498 & ~n37507;
  assign n37531 = ~n37492 & n37530;
  assign n37532 = n37479 & ~n37486;
  assign n37533 = n37531 & n37532;
  assign n37534 = n37511 & n37532;
  assign n37535 = n37492 & n37534;
  assign n37536 = ~n37533 & ~n37535;
  assign n37537 = ~n37486 & ~n37492;
  assign n37538 = n37507 & n37537;
  assign n37539 = ~n37498 & n37538;
  assign n37540 = ~n37479 & n37539;
  assign n37541 = n37536 & ~n37540;
  assign n37542 = ~n37479 & ~n37486;
  assign n37543 = ~n37498 & n37542;
  assign n37544 = n37479 & n37511;
  assign n37545 = ~n37486 & n37544;
  assign n37546 = ~n37486 & n37492;
  assign n37547 = n37498 & n37546;
  assign n37548 = ~n37500 & ~n37547;
  assign n37549 = n37479 & ~n37548;
  assign n37550 = ~n37545 & ~n37549;
  assign n37551 = n37492 & n37511;
  assign n37552 = ~n37486 & n37551;
  assign n37553 = n37507 & n37516;
  assign n37554 = n37486 & n37553;
  assign n37555 = ~n37552 & ~n37554;
  assign n37556 = ~n37479 & n37486;
  assign n37557 = n37516 & n37556;
  assign n37558 = ~n37492 & n37519;
  assign n37559 = ~n37479 & n37558;
  assign n37560 = ~n37557 & ~n37559;
  assign n37561 = n37555 & n37560;
  assign n37562 = n37550 & n37561;
  assign n37563 = ~n37543 & n37562;
  assign n37564 = ~n37473 & ~n37563;
  assign n37565 = n37486 & n37508;
  assign n37566 = n37492 & n37530;
  assign n37567 = ~n37486 & n37566;
  assign n37568 = ~n37565 & ~n37567;
  assign n37569 = ~n37479 & ~n37568;
  assign n37570 = ~n37564 & ~n37569;
  assign n37571 = n37541 & n37570;
  assign n37572 = ~n37529 & n37571;
  assign n37573 = ~pi0801 & ~n37572;
  assign n37574 = pi0801 & n37572;
  assign po0839 = n37573 | n37574;
  assign n37576 = pi3683 & pi9040;
  assign n37577 = pi3687 & ~pi9040;
  assign n37578 = ~n37576 & ~n37577;
  assign n37579 = pi0780 & n37578;
  assign n37580 = ~pi0780 & ~n37578;
  assign n37581 = ~n37579 & ~n37580;
  assign n37582 = pi3700 & pi9040;
  assign n37583 = pi3697 & ~pi9040;
  assign n37584 = ~n37582 & ~n37583;
  assign n37585 = pi0784 & n37584;
  assign n37586 = ~pi0784 & ~n37584;
  assign n37587 = ~n37585 & ~n37586;
  assign n37588 = pi3687 & pi9040;
  assign n37589 = pi3694 & ~pi9040;
  assign n37590 = ~n37588 & ~n37589;
  assign n37591 = ~pi0793 & ~n37590;
  assign n37592 = pi0793 & n37590;
  assign n37593 = ~n37591 & ~n37592;
  assign n37594 = pi3662 & pi9040;
  assign n37595 = pi3752 & ~pi9040;
  assign n37596 = ~n37594 & ~n37595;
  assign n37597 = ~pi0772 & ~n37596;
  assign n37598 = pi0772 & ~n37594;
  assign n37599 = ~n37595 & n37598;
  assign n37600 = ~n37597 & ~n37599;
  assign n37601 = pi3669 & pi9040;
  assign n37602 = pi3680 & ~pi9040;
  assign n37603 = ~n37601 & ~n37602;
  assign n37604 = ~pi0777 & n37603;
  assign n37605 = pi0777 & ~n37603;
  assign n37606 = ~n37604 & ~n37605;
  assign n37607 = ~n37600 & n37606;
  assign n37608 = ~n37593 & n37607;
  assign n37609 = ~n37587 & n37608;
  assign n37610 = n37587 & ~n37593;
  assign n37611 = n37606 & n37610;
  assign n37612 = n37600 & n37611;
  assign n37613 = ~n37609 & ~n37612;
  assign n37614 = n37581 & ~n37613;
  assign n37615 = ~n37587 & n37593;
  assign n37616 = ~n37606 & n37615;
  assign n37617 = ~n37600 & n37616;
  assign n37618 = ~n37581 & n37617;
  assign n37619 = pi3673 & ~pi9040;
  assign n37620 = pi3659 & pi9040;
  assign n37621 = ~n37619 & ~n37620;
  assign n37622 = ~pi0797 & ~n37621;
  assign n37623 = pi0797 & n37621;
  assign n37624 = ~n37622 & ~n37623;
  assign n37625 = n37600 & n37606;
  assign n37626 = n37593 & n37625;
  assign n37627 = n37581 & n37626;
  assign n37628 = ~n37617 & ~n37627;
  assign n37629 = ~n37587 & n37600;
  assign n37630 = ~n37593 & n37629;
  assign n37631 = ~n37600 & n37615;
  assign n37632 = ~n37630 & ~n37631;
  assign n37633 = ~n37581 & ~n37632;
  assign n37634 = ~n37581 & ~n37593;
  assign n37635 = n37607 & n37634;
  assign n37636 = n37587 & n37635;
  assign n37637 = n37587 & n37593;
  assign n37638 = ~n37606 & n37637;
  assign n37639 = n37600 & n37638;
  assign n37640 = n37581 & ~n37593;
  assign n37641 = ~n37606 & n37640;
  assign n37642 = ~n37600 & n37641;
  assign n37643 = ~n37639 & ~n37642;
  assign n37644 = ~n37636 & n37643;
  assign n37645 = ~n37633 & n37644;
  assign n37646 = n37628 & n37645;
  assign n37647 = n37624 & ~n37646;
  assign n37648 = ~n37587 & n37627;
  assign n37649 = ~n37647 & ~n37648;
  assign n37650 = ~n37618 & n37649;
  assign n37651 = ~n37614 & n37650;
  assign n37652 = n37581 & n37587;
  assign n37653 = n37593 & ~n37600;
  assign n37654 = n37652 & n37653;
  assign n37655 = n37581 & n37608;
  assign n37656 = ~n37654 & ~n37655;
  assign n37657 = n37600 & ~n37606;
  assign n37658 = n37593 & n37657;
  assign n37659 = n37581 & n37658;
  assign n37660 = ~n37593 & n37657;
  assign n37661 = ~n37587 & n37660;
  assign n37662 = ~n37659 & ~n37661;
  assign n37663 = n37593 & n37607;
  assign n37664 = n37587 & n37663;
  assign n37665 = ~n37609 & ~n37664;
  assign n37666 = n37587 & n37625;
  assign n37667 = ~n37593 & ~n37606;
  assign n37668 = ~n37666 & ~n37667;
  assign n37669 = ~n37581 & ~n37668;
  assign n37670 = n37665 & ~n37669;
  assign n37671 = n37662 & n37670;
  assign n37672 = n37656 & n37671;
  assign n37673 = ~n37624 & ~n37672;
  assign n37674 = n37651 & ~n37673;
  assign n37675 = ~pi0806 & ~n37674;
  assign n37676 = pi0806 & n37651;
  assign n37677 = ~n37673 & n37676;
  assign po0840 = n37675 | n37677;
  assign n37679 = ~n37648 & ~n37654;
  assign n37680 = ~n37606 & n37610;
  assign n37681 = ~n37600 & n37680;
  assign n37682 = ~n37639 & ~n37681;
  assign n37683 = ~n37609 & n37682;
  assign n37684 = ~n37581 & ~n37683;
  assign n37685 = ~n37600 & ~n37606;
  assign n37686 = n37581 & n37685;
  assign n37687 = ~n37587 & n37686;
  assign n37688 = n37600 & n37610;
  assign n37689 = ~n37593 & n37625;
  assign n37690 = ~n37688 & ~n37689;
  assign n37691 = n37581 & ~n37690;
  assign n37692 = ~n37687 & ~n37691;
  assign n37693 = ~n37581 & ~n37587;
  assign n37694 = n37657 & n37693;
  assign n37695 = ~n37581 & n37608;
  assign n37696 = ~n37694 & ~n37695;
  assign n37697 = n37692 & n37696;
  assign n37698 = n37600 & n37615;
  assign n37699 = ~n37609 & ~n37698;
  assign n37700 = ~n37664 & n37699;
  assign n37701 = n37697 & n37700;
  assign n37702 = ~n37624 & ~n37701;
  assign n37703 = ~n37617 & ~n37689;
  assign n37704 = ~n37666 & n37703;
  assign n37705 = ~n37581 & ~n37704;
  assign n37706 = n37581 & ~n37587;
  assign n37707 = n37660 & n37706;
  assign n37708 = n37682 & ~n37707;
  assign n37709 = n37581 & n37663;
  assign n37710 = n37708 & ~n37709;
  assign n37711 = ~n37705 & n37710;
  assign n37712 = n37624 & ~n37711;
  assign n37713 = ~n37702 & ~n37712;
  assign n37714 = ~n37684 & n37713;
  assign n37715 = n37679 & n37714;
  assign n37716 = pi0814 & ~n37715;
  assign n37717 = ~pi0814 & n37715;
  assign po0841 = n37716 | n37717;
  assign n37719 = pi3658 & pi9040;
  assign n37720 = ~pi3689 & ~pi9040;
  assign n37721 = ~n37719 & ~n37720;
  assign n37722 = ~pi0778 & ~n37721;
  assign n37723 = pi0778 & n37721;
  assign n37724 = ~n37722 & ~n37723;
  assign n37725 = pi3664 & pi9040;
  assign n37726 = pi3690 & ~pi9040;
  assign n37727 = ~n37725 & ~n37726;
  assign n37728 = pi0783 & n37727;
  assign n37729 = ~pi0783 & ~n37727;
  assign n37730 = ~n37728 & ~n37729;
  assign n37731 = pi3709 & pi9040;
  assign n37732 = pi3706 & ~pi9040;
  assign n37733 = ~n37731 & ~n37732;
  assign n37734 = ~pi0797 & ~n37733;
  assign n37735 = pi0797 & ~n37731;
  assign n37736 = ~n37732 & n37735;
  assign n37737 = ~n37734 & ~n37736;
  assign n37738 = pi3667 & pi9040;
  assign n37739 = pi3695 & ~pi9040;
  assign n37740 = ~n37738 & ~n37739;
  assign n37741 = ~pi0777 & n37740;
  assign n37742 = pi0777 & ~n37740;
  assign n37743 = ~n37741 & ~n37742;
  assign n37744 = pi3655 & pi9040;
  assign n37745 = pi3701 & ~pi9040;
  assign n37746 = ~n37744 & ~n37745;
  assign n37747 = ~pi0773 & ~n37746;
  assign n37748 = pi0773 & ~n37744;
  assign n37749 = ~n37745 & n37748;
  assign n37750 = ~n37747 & ~n37749;
  assign n37751 = ~n37743 & ~n37750;
  assign n37752 = n37737 & n37751;
  assign n37753 = n37730 & n37752;
  assign n37754 = ~n37730 & ~n37743;
  assign n37755 = n37750 & n37754;
  assign n37756 = pi3702 & pi9040;
  assign n37757 = pi3667 & ~pi9040;
  assign n37758 = ~n37756 & ~n37757;
  assign n37759 = ~pi0775 & n37758;
  assign n37760 = pi0775 & ~n37758;
  assign n37761 = ~n37759 & ~n37760;
  assign n37762 = ~n37737 & n37754;
  assign n37763 = n37737 & n37750;
  assign n37764 = n37743 & n37763;
  assign n37765 = ~n37762 & ~n37764;
  assign n37766 = n37761 & ~n37765;
  assign n37767 = ~n37755 & ~n37766;
  assign n37768 = ~n37737 & ~n37750;
  assign n37769 = n37730 & n37768;
  assign n37770 = ~n37743 & n37763;
  assign n37771 = ~n37737 & n37743;
  assign n37772 = ~n37730 & n37743;
  assign n37773 = ~n37750 & n37772;
  assign n37774 = ~n37771 & ~n37773;
  assign n37775 = ~n37770 & n37774;
  assign n37776 = ~n37769 & n37775;
  assign n37777 = ~n37761 & ~n37776;
  assign n37778 = n37767 & ~n37777;
  assign n37779 = ~n37753 & n37778;
  assign n37780 = n37724 & ~n37779;
  assign n37781 = ~n37737 & n37750;
  assign n37782 = n37743 & n37781;
  assign n37783 = ~n37730 & n37782;
  assign n37784 = n37743 & n37768;
  assign n37785 = n37730 & n37784;
  assign n37786 = ~n37753 & ~n37785;
  assign n37787 = ~n37783 & n37786;
  assign n37788 = ~n37761 & ~n37787;
  assign n37789 = ~n37780 & ~n37788;
  assign n37790 = ~n37730 & n37770;
  assign n37791 = n37737 & n37743;
  assign n37792 = n37761 & n37791;
  assign n37793 = n37730 & n37792;
  assign n37794 = ~n37730 & ~n37761;
  assign n37795 = n37751 & n37794;
  assign n37796 = ~n37743 & n37781;
  assign n37797 = n37730 & n37796;
  assign n37798 = ~n37795 & ~n37797;
  assign n37799 = ~n37737 & ~n37743;
  assign n37800 = n37730 & n37799;
  assign n37801 = n37737 & ~n37750;
  assign n37802 = n37743 & n37801;
  assign n37803 = ~n37800 & ~n37802;
  assign n37804 = n37761 & ~n37803;
  assign n37805 = ~n37737 & n37761;
  assign n37806 = n37743 & n37805;
  assign n37807 = ~n37730 & n37806;
  assign n37808 = ~n37804 & ~n37807;
  assign n37809 = n37798 & n37808;
  assign n37810 = ~n37724 & ~n37809;
  assign n37811 = ~n37793 & ~n37810;
  assign n37812 = ~n37790 & n37811;
  assign n37813 = n37789 & n37812;
  assign n37814 = ~pi0809 & ~n37813;
  assign n37815 = ~n37780 & ~n37790;
  assign n37816 = ~n37788 & n37815;
  assign n37817 = n37811 & n37816;
  assign n37818 = pi0809 & n37817;
  assign po0842 = n37814 | n37818;
  assign n37820 = ~n37473 & n37479;
  assign n37821 = ~n37486 & n37499;
  assign n37822 = n37486 & n37551;
  assign n37823 = ~n37486 & n37508;
  assign n37824 = ~n37822 & ~n37823;
  assign n37825 = ~n37821 & n37824;
  assign n37826 = n37820 & ~n37825;
  assign n37827 = ~n37507 & n37537;
  assign n37828 = n37486 & n37566;
  assign n37829 = ~n37827 & ~n37828;
  assign n37830 = ~n37509 & ~n37512;
  assign n37831 = n37829 & n37830;
  assign n37832 = ~n37479 & ~n37831;
  assign n37833 = n37486 & n37558;
  assign n37834 = ~n37832 & ~n37833;
  assign n37835 = ~n37473 & ~n37834;
  assign n37836 = ~n37826 & ~n37835;
  assign n37837 = n37492 & n37542;
  assign n37838 = n37507 & n37837;
  assign n37839 = ~n37513 & ~n37838;
  assign n37840 = ~n37508 & ~n37530;
  assign n37841 = n37486 & ~n37840;
  assign n37842 = ~n37531 & ~n37841;
  assign n37843 = n37479 & ~n37842;
  assign n37844 = ~n37520 & ~n37821;
  assign n37845 = ~n37822 & n37844;
  assign n37846 = ~n37479 & ~n37845;
  assign n37847 = ~n37843 & ~n37846;
  assign n37848 = n37486 & n37531;
  assign n37849 = ~n37554 & ~n37848;
  assign n37850 = ~n37539 & n37849;
  assign n37851 = ~n37545 & n37850;
  assign n37852 = n37847 & n37851;
  assign n37853 = n37473 & ~n37852;
  assign n37854 = n37839 & ~n37853;
  assign n37855 = n37836 & n37854;
  assign n37856 = pi0802 & ~n37855;
  assign n37857 = ~pi0802 & n37839;
  assign n37858 = n37836 & n37857;
  assign n37859 = ~n37853 & n37858;
  assign po0843 = n37856 | n37859;
  assign n37861 = ~n37088 & n37105;
  assign n37862 = ~n37136 & ~n37861;
  assign n37863 = n37075 & ~n37862;
  assign n37864 = n37095 & n37127;
  assign n37865 = ~n37323 & ~n37864;
  assign n37866 = ~n37075 & ~n37865;
  assign n37867 = ~n37095 & n37122;
  assign n37868 = ~n37344 & ~n37867;
  assign n37869 = ~n37104 & n37868;
  assign n37870 = ~n37866 & n37869;
  assign n37871 = ~n37863 & n37870;
  assign n37872 = ~n37319 & ~n37330;
  assign n37873 = n37871 & n37872;
  assign n37874 = n37114 & ~n37873;
  assign n37875 = n37089 & n37317;
  assign n37876 = n37145 & ~n37875;
  assign n37877 = ~n37075 & ~n37876;
  assign n37878 = ~n37095 & n37133;
  assign n37879 = ~n37877 & ~n37878;
  assign n37880 = n37082 & n37105;
  assign n37881 = n37095 & n37118;
  assign n37882 = ~n37880 & ~n37881;
  assign n37883 = ~n37075 & ~n37882;
  assign n37884 = ~n37075 & n37127;
  assign n37885 = ~n37095 & n37884;
  assign n37886 = ~n37883 & ~n37885;
  assign n37887 = n37879 & n37886;
  assign n37888 = ~n37114 & ~n37887;
  assign n37889 = ~n37122 & ~n37129;
  assign n37890 = ~n37324 & n37889;
  assign n37891 = n37150 & ~n37890;
  assign n37892 = ~n37888 & ~n37891;
  assign n37893 = ~n37104 & ~n37319;
  assign n37894 = n37075 & ~n37893;
  assign n37895 = n37892 & ~n37894;
  assign n37896 = ~n37874 & n37895;
  assign n37897 = ~pi0807 & n37896;
  assign n37898 = pi0807 & ~n37896;
  assign po0845 = n37897 | n37898;
  assign n37900 = ~n37193 & n37227;
  assign n37901 = ~n37278 & ~n37900;
  assign n37902 = n37199 & ~n37901;
  assign n37903 = n37224 & n37274;
  assign n37904 = ~n37902 & ~n37903;
  assign n37905 = ~n37247 & n37904;
  assign n37906 = ~n37180 & n37193;
  assign n37907 = n37174 & n37906;
  assign n37908 = n37186 & n37907;
  assign n37909 = ~n37207 & ~n37908;
  assign n37910 = ~n37227 & n37909;
  assign n37911 = n37199 & ~n37910;
  assign n37912 = n37168 & n37911;
  assign n37913 = ~n37199 & n37287;
  assign n37914 = ~n37218 & ~n37245;
  assign n37915 = ~n37212 & n37914;
  assign n37916 = ~n37913 & n37915;
  assign n37917 = n37168 & ~n37916;
  assign n37918 = ~n37174 & ~n37199;
  assign n37919 = n37186 & n37918;
  assign n37920 = n37180 & n37919;
  assign n37921 = ~n37193 & n37920;
  assign n37922 = n37193 & n37259;
  assign n37923 = ~n37920 & ~n37922;
  assign n37924 = ~n37277 & n37923;
  assign n37925 = n37186 & n37216;
  assign n37926 = n37193 & n37204;
  assign n37927 = ~n37223 & ~n37926;
  assign n37928 = n37199 & ~n37927;
  assign n37929 = ~n37925 & ~n37928;
  assign n37930 = n37924 & n37929;
  assign n37931 = ~n37168 & ~n37930;
  assign n37932 = ~n37921 & ~n37931;
  assign n37933 = ~n37917 & n37932;
  assign n37934 = ~n37912 & n37933;
  assign n37935 = n37905 & n37934;
  assign n37936 = pi0830 & ~n37935;
  assign n37937 = ~pi0830 & n37905;
  assign n37938 = n37934 & n37937;
  assign po0846 = n37936 | n37938;
  assign n37940 = ~n37730 & n37761;
  assign n37941 = n37737 & n37940;
  assign n37942 = ~n37743 & n37768;
  assign n37943 = n37730 & n37942;
  assign n37944 = n37730 & n37782;
  assign n37945 = ~n37943 & ~n37944;
  assign n37946 = ~n37730 & n37784;
  assign n37947 = ~n37764 & ~n37946;
  assign n37948 = ~n37761 & ~n37947;
  assign n37949 = n37945 & ~n37948;
  assign n37950 = ~n37941 & n37949;
  assign n37951 = n37724 & ~n37950;
  assign n37952 = n37730 & n37737;
  assign n37953 = n37743 & n37952;
  assign n37954 = ~n37750 & n37953;
  assign n37955 = n37761 & n37954;
  assign n37956 = n37794 & n37802;
  assign n37957 = ~n37762 & ~n37956;
  assign n37958 = ~n37764 & ~n37796;
  assign n37959 = ~n37730 & n37781;
  assign n37960 = n37958 & ~n37959;
  assign n37961 = n37761 & ~n37960;
  assign n37962 = ~n37761 & n37770;
  assign n37963 = n37786 & ~n37962;
  assign n37964 = ~n37961 & n37963;
  assign n37965 = n37957 & n37964;
  assign n37966 = ~n37724 & ~n37965;
  assign n37967 = ~n37955 & ~n37966;
  assign n37968 = ~n37951 & n37967;
  assign n37969 = n37794 & n37796;
  assign n37970 = n37751 & ~n37761;
  assign n37971 = n37730 & n37970;
  assign n37972 = ~n37969 & ~n37971;
  assign n37973 = ~n37761 & n37944;
  assign n37974 = n37972 & ~n37973;
  assign n37975 = n37968 & n37974;
  assign n37976 = ~pi0810 & ~n37975;
  assign n37977 = pi0810 & n37974;
  assign n37978 = n37967 & n37977;
  assign n37979 = ~n37951 & n37978;
  assign po0847 = n37976 | n37979;
  assign n37981 = ~n37386 & n37415;
  assign n37982 = ~n37437 & ~n37455;
  assign n37983 = ~n37392 & ~n37982;
  assign n37984 = ~n37981 & ~n37983;
  assign n37985 = ~n37430 & n37984;
  assign n37986 = ~n37386 & n37392;
  assign n37987 = n37433 & n37986;
  assign n37988 = ~n37421 & ~n37987;
  assign n37989 = ~n37449 & n37988;
  assign n37990 = n37985 & n37989;
  assign n37991 = n37367 & ~n37990;
  assign n37992 = ~n37401 & n37408;
  assign n37993 = ~n37386 & n37992;
  assign n37994 = ~n37406 & ~n37993;
  assign n37995 = n37386 & n37448;
  assign n37996 = ~n37416 & ~n37995;
  assign n37997 = ~n37373 & ~n37386;
  assign n37998 = ~n37422 & ~n37997;
  assign n37999 = ~n37435 & n37998;
  assign n38000 = n37392 & ~n37999;
  assign n38001 = ~n37392 & n37433;
  assign n38002 = ~n37386 & n37420;
  assign n38003 = ~n38001 & ~n38002;
  assign n38004 = ~n38000 & n38003;
  assign n38005 = n37996 & n38004;
  assign n38006 = n37994 & n38005;
  assign n38007 = ~n37367 & ~n38006;
  assign n38008 = ~n37991 & ~n38007;
  assign n38009 = pi0812 & ~n38008;
  assign n38010 = ~pi0812 & ~n37991;
  assign n38011 = ~n38007 & n38010;
  assign po0848 = n38009 | n38011;
  assign n38013 = ~n37730 & n37942;
  assign n38014 = ~n37782 & ~n37790;
  assign n38015 = n37730 & n37751;
  assign n38016 = ~n37730 & n37802;
  assign n38017 = ~n38015 & ~n38016;
  assign n38018 = n38014 & n38017;
  assign n38019 = n37761 & ~n38018;
  assign n38020 = n37730 & n37763;
  assign n38021 = ~n37762 & ~n38020;
  assign n38022 = ~n37784 & n38021;
  assign n38023 = ~n37761 & ~n38022;
  assign n38024 = n37730 & n37743;
  assign n38025 = n37750 & n38024;
  assign n38026 = n37737 & n38025;
  assign n38027 = ~n38023 & ~n38026;
  assign n38028 = ~n38019 & n38027;
  assign n38029 = ~n38013 & n38028;
  assign n38030 = ~n37724 & ~n38029;
  assign n38031 = n37730 & n37761;
  assign n38032 = n37770 & n38031;
  assign n38033 = n37761 & n37784;
  assign n38034 = n37761 & n37796;
  assign n38035 = ~n38033 & ~n38034;
  assign n38036 = ~n37730 & ~n38035;
  assign n38037 = ~n38032 & ~n38036;
  assign n38038 = ~n37730 & n37752;
  assign n38039 = ~n37954 & ~n38038;
  assign n38040 = n37730 & n37781;
  assign n38041 = ~n37730 & n37763;
  assign n38042 = ~n38040 & ~n38041;
  assign n38043 = ~n37752 & n38042;
  assign n38044 = ~n37782 & n38043;
  assign n38045 = ~n37761 & ~n38044;
  assign n38046 = ~n37730 & n37764;
  assign n38047 = ~n38045 & ~n38046;
  assign n38048 = n38039 & n38047;
  assign n38049 = n38037 & n38048;
  assign n38050 = n37724 & ~n38049;
  assign n38051 = n37761 & ~n37945;
  assign n38052 = ~n38050 & ~n38051;
  assign n38053 = ~n37785 & ~n38038;
  assign n38054 = ~n37761 & ~n38053;
  assign n38055 = n38052 & ~n38054;
  assign n38056 = ~n38030 & n38055;
  assign n38057 = pi0820 & ~n38056;
  assign n38058 = ~pi0820 & n38056;
  assign po0849 = n38057 | n38058;
  assign n38060 = n37593 & n37685;
  assign n38061 = n37587 & n38060;
  assign n38062 = n37587 & n37657;
  assign n38063 = ~n37593 & n37685;
  assign n38064 = ~n37587 & n38063;
  assign n38065 = ~n38062 & ~n38064;
  assign n38066 = ~n37581 & ~n38065;
  assign n38067 = ~n38061 & ~n38066;
  assign n38068 = n37587 & n37686;
  assign n38069 = ~n37655 & ~n38068;
  assign n38070 = n38067 & n38069;
  assign n38071 = n37587 & n37626;
  assign n38072 = ~n37587 & n37663;
  assign n38073 = ~n38071 & ~n38072;
  assign n38074 = n38070 & n38073;
  assign n38075 = n37624 & ~n38074;
  assign n38076 = ~n37581 & ~n37624;
  assign n38077 = ~n37600 & n37610;
  assign n38078 = ~n37593 & n37606;
  assign n38079 = ~n38077 & ~n38078;
  assign n38080 = n38076 & ~n38079;
  assign n38081 = ~n37617 & ~n37630;
  assign n38082 = n37593 & n37652;
  assign n38083 = ~n37685 & n38082;
  assign n38084 = ~n37627 & ~n38083;
  assign n38085 = n38081 & n38084;
  assign n38086 = ~n37624 & ~n38085;
  assign n38087 = n37689 & n37693;
  assign n38088 = ~n37587 & n37658;
  assign n38089 = ~n38072 & ~n38088;
  assign n38090 = ~n37581 & ~n38089;
  assign n38091 = ~n38087 & ~n38090;
  assign n38092 = n37581 & n37617;
  assign n38093 = n38091 & ~n38092;
  assign n38094 = ~n38086 & n38093;
  assign n38095 = ~n38080 & n38094;
  assign n38096 = ~n38075 & n38095;
  assign n38097 = ~n37707 & n38096;
  assign n38098 = ~pi0815 & ~n38097;
  assign n38099 = ~n37707 & n38095;
  assign n38100 = pi0815 & n38099;
  assign n38101 = ~n38075 & n38100;
  assign po0850 = n38098 | n38101;
  assign n38103 = ~n37520 & ~n37531;
  assign n38104 = n37479 & ~n38103;
  assign n38105 = n37486 & n37509;
  assign n38106 = ~n38104 & ~n38105;
  assign n38107 = n37486 & n37498;
  assign n38108 = ~n37516 & ~n38107;
  assign n38109 = ~n37566 & n38108;
  assign n38110 = ~n37479 & ~n38109;
  assign n38111 = n38106 & ~n38110;
  assign n38112 = ~n37473 & ~n38111;
  assign n38113 = ~n37486 & n37553;
  assign n38114 = n37479 & n38113;
  assign n38115 = ~n37535 & ~n38114;
  assign n38116 = ~n37540 & n38115;
  assign n38117 = ~n37479 & n37498;
  assign n38118 = n37546 & n38117;
  assign n38119 = n37486 & n37520;
  assign n38120 = n37479 & n37516;
  assign n38121 = ~n38119 & ~n38120;
  assign n38122 = ~n37848 & n38121;
  assign n38123 = ~n38118 & n38122;
  assign n38124 = ~n37507 & n37546;
  assign n38125 = ~n37539 & ~n38124;
  assign n38126 = n38123 & n38125;
  assign n38127 = ~n37559 & n38126;
  assign n38128 = n37473 & ~n38127;
  assign n38129 = n38116 & ~n38128;
  assign n38130 = ~n38112 & n38129;
  assign n38131 = ~pi0808 & ~n38130;
  assign n38132 = pi0808 & n38116;
  assign n38133 = ~n38112 & n38132;
  assign n38134 = ~n38128 & n38133;
  assign po0851 = n38131 | n38134;
  assign n38136 = ~n37946 & ~n38038;
  assign n38137 = ~n38026 & n38136;
  assign n38138 = n37761 & ~n38137;
  assign n38139 = ~n37956 & ~n37973;
  assign n38140 = ~n37954 & ~n38034;
  assign n38141 = ~n37942 & ~n38041;
  assign n38142 = ~n37761 & ~n38141;
  assign n38143 = ~n37790 & ~n38142;
  assign n38144 = n38140 & n38143;
  assign n38145 = n37724 & ~n38144;
  assign n38146 = n37743 & n37750;
  assign n38147 = ~n37771 & ~n38146;
  assign n38148 = n37730 & ~n38147;
  assign n38149 = ~n37752 & ~n37959;
  assign n38150 = ~n37761 & ~n38149;
  assign n38151 = n37730 & n37750;
  assign n38152 = ~n37764 & ~n38151;
  assign n38153 = ~n37768 & n38152;
  assign n38154 = n37761 & ~n38153;
  assign n38155 = ~n38150 & ~n38154;
  assign n38156 = ~n38148 & n38155;
  assign n38157 = ~n37724 & ~n38156;
  assign n38158 = ~n38145 & ~n38157;
  assign n38159 = n38139 & n38158;
  assign n38160 = ~n38138 & n38159;
  assign n38161 = ~pi0833 & ~n38160;
  assign n38162 = pi0833 & n38139;
  assign n38163 = ~n38138 & n38162;
  assign n38164 = n38158 & n38163;
  assign po0852 = n38161 | n38164;
  assign n38166 = n37193 & ~n37299;
  assign n38167 = n37174 & n38166;
  assign n38168 = n37186 & n37276;
  assign n38169 = ~n37255 & ~n38168;
  assign n38170 = ~n37207 & n38169;
  assign n38171 = ~n37199 & ~n38170;
  assign n38172 = ~n37231 & ~n37287;
  assign n38173 = n37199 & ~n38172;
  assign n38174 = ~n38171 & ~n38173;
  assign n38175 = ~n38167 & n38174;
  assign n38176 = ~n37193 & n37224;
  assign n38177 = n38175 & ~n38176;
  assign n38178 = ~n37168 & ~n38177;
  assign n38179 = n37203 & ~n38172;
  assign n38180 = ~n37227 & ~n37232;
  assign n38181 = ~n37207 & ~n37224;
  assign n38182 = n38180 & n38181;
  assign n38183 = n37193 & ~n38182;
  assign n38184 = ~n38179 & ~n38183;
  assign n38185 = ~n37278 & n38184;
  assign n38186 = n37168 & ~n38185;
  assign n38187 = ~n38178 & ~n38186;
  assign n38188 = n37193 & n37287;
  assign n38189 = ~n38176 & ~n38188;
  assign n38190 = n37199 & ~n38189;
  assign n38191 = n38187 & ~n38190;
  assign n38192 = pi0817 & ~n38191;
  assign n38193 = ~pi0817 & ~n38190;
  assign n38194 = ~n38186 & n38193;
  assign n38195 = ~n38178 & n38194;
  assign po0853 = n38192 | n38195;
  assign n38197 = n37075 & n37133;
  assign n38198 = ~n37095 & n37118;
  assign n38199 = ~n37117 & ~n38198;
  assign n38200 = n37075 & ~n38199;
  assign n38201 = ~n37075 & ~n37346;
  assign n38202 = ~n38200 & ~n38201;
  assign n38203 = ~n37334 & n38202;
  assign n38204 = n37114 & ~n38203;
  assign n38205 = ~n38197 & ~n38204;
  assign n38206 = n37102 & n37310;
  assign n38207 = ~n37322 & ~n38206;
  assign n38208 = ~n37082 & ~n38207;
  assign n38209 = ~n37104 & ~n38208;
  assign n38210 = ~n37323 & n38209;
  assign n38211 = ~n37075 & n37119;
  assign n38212 = n37095 & n37136;
  assign n38213 = ~n38211 & ~n38212;
  assign n38214 = n38210 & n38213;
  assign n38215 = ~n37114 & ~n38214;
  assign n38216 = ~n37867 & ~n37881;
  assign n38217 = ~n37075 & ~n38216;
  assign n38218 = ~n38215 & ~n38217;
  assign n38219 = n38205 & n38218;
  assign n38220 = ~pi0846 & ~n38219;
  assign n38221 = ~n38204 & n38218;
  assign n38222 = pi0846 & n38221;
  assign n38223 = ~n38197 & n38222;
  assign po0854 = n38220 | n38223;
  assign n38225 = ~n36985 & n36992;
  assign n38226 = ~n36973 & n38225;
  assign n38227 = n36979 & n38226;
  assign n38228 = n36992 & n37015;
  assign n38229 = n36985 & ~n36998;
  assign n38230 = ~n36979 & n38229;
  assign n38231 = ~n37001 & ~n38230;
  assign n38232 = ~n38228 & n38231;
  assign n38233 = ~n38227 & n38232;
  assign n38234 = n36973 & n37009;
  assign n38235 = n38233 & ~n38234;
  assign n38236 = n37039 & ~n38235;
  assign n38237 = ~n36979 & n37003;
  assign n38238 = ~n37057 & ~n38237;
  assign n38239 = n36973 & ~n38238;
  assign n38240 = ~n37039 & n37041;
  assign n38241 = ~n36973 & n38240;
  assign n38242 = ~n36979 & n36985;
  assign n38243 = ~n36992 & n38242;
  assign n38244 = ~n38229 & ~n38243;
  assign n38245 = ~n37003 & n38244;
  assign n38246 = n36973 & ~n38245;
  assign n38247 = ~n36985 & n37026;
  assign n38248 = ~n36979 & n38247;
  assign n38249 = ~n38246 & ~n38248;
  assign n38250 = ~n37039 & ~n38249;
  assign n38251 = ~n38241 & ~n38250;
  assign n38252 = ~n38239 & n38251;
  assign n38253 = ~n37001 & ~n37010;
  assign n38254 = n36979 & ~n36998;
  assign n38255 = ~n36985 & n38254;
  assign n38256 = ~n36979 & n37056;
  assign n38257 = ~n38255 & ~n38256;
  assign n38258 = n38253 & n38257;
  assign n38259 = ~n36973 & ~n38258;
  assign n38260 = n38252 & ~n38259;
  assign n38261 = ~n38236 & n38260;
  assign n38262 = ~pi0827 & ~n38261;
  assign n38263 = pi0827 & n38252;
  assign n38264 = ~n38236 & n38263;
  assign n38265 = ~n38259 & n38264;
  assign po0855 = n38262 | n38265;
  assign n38267 = ~n38071 & ~n38077;
  assign n38268 = n37624 & ~n38267;
  assign n38269 = ~n37581 & n38060;
  assign n38270 = ~n37616 & ~n37631;
  assign n38271 = ~n37581 & ~n38270;
  assign n38272 = ~n38269 & ~n38271;
  assign n38273 = n37624 & ~n38272;
  assign n38274 = ~n38268 & ~n38273;
  assign n38275 = ~n37587 & n37626;
  assign n38276 = ~n37617 & ~n37639;
  assign n38277 = ~n37587 & n37607;
  assign n38278 = ~n37612 & ~n38277;
  assign n38279 = n37581 & ~n38278;
  assign n38280 = ~n37587 & n37625;
  assign n38281 = ~n37660 & ~n38280;
  assign n38282 = ~n37581 & ~n38281;
  assign n38283 = ~n38279 & ~n38282;
  assign n38284 = n38276 & n38283;
  assign n38285 = ~n38275 & n38284;
  assign n38286 = ~n37624 & ~n38285;
  assign n38287 = ~n37664 & n37682;
  assign n38288 = n37581 & ~n38287;
  assign n38289 = ~n38286 & ~n38288;
  assign n38290 = ~n37581 & n37587;
  assign n38291 = n37626 & n38290;
  assign n38292 = ~n37636 & ~n38291;
  assign n38293 = ~n37630 & ~n37667;
  assign n38294 = n37581 & ~n38293;
  assign n38295 = n37624 & n38294;
  assign n38296 = n38292 & ~n38295;
  assign n38297 = n38289 & n38296;
  assign n38298 = n38274 & n38297;
  assign n38299 = ~pi0821 & ~n38298;
  assign n38300 = pi0821 & n38296;
  assign n38301 = n38274 & n38300;
  assign n38302 = n38289 & n38301;
  assign po0856 = n38299 | n38302;
  assign n38304 = ~n36979 & n37030;
  assign n38305 = ~n37027 & ~n38255;
  assign n38306 = n36973 & ~n38305;
  assign n38307 = ~n38304 & ~n38306;
  assign n38308 = ~n36973 & ~n36979;
  assign n38309 = ~n36998 & n38308;
  assign n38310 = n36992 & n38309;
  assign n38311 = n37002 & n37042;
  assign n38312 = ~n38310 & ~n38311;
  assign n38313 = ~n36973 & n37000;
  assign n38314 = n38312 & ~n38313;
  assign n38315 = ~n37010 & ~n37016;
  assign n38316 = n36998 & n37048;
  assign n38317 = n38315 & ~n38316;
  assign n38318 = n38314 & n38317;
  assign n38319 = n38307 & n38318;
  assign n38320 = ~n37039 & ~n38319;
  assign n38321 = ~n37009 & ~n37027;
  assign n38322 = n36979 & ~n38321;
  assign n38323 = n36992 & n37045;
  assign n38324 = ~n37056 & ~n38323;
  assign n38325 = n36979 & n38229;
  assign n38326 = n38324 & ~n38325;
  assign n38327 = n36973 & ~n38326;
  assign n38328 = ~n36979 & n37026;
  assign n38329 = ~n38228 & ~n38328;
  assign n38330 = ~n36973 & ~n38329;
  assign n38331 = ~n38237 & ~n38330;
  assign n38332 = ~n38327 & n38331;
  assign n38333 = ~n38322 & n38332;
  assign n38334 = n37039 & ~n38333;
  assign n38335 = n36973 & n37046;
  assign n38336 = ~n38334 & ~n38335;
  assign n38337 = n37021 & n38308;
  assign n38338 = ~n36998 & n38337;
  assign n38339 = n38336 & ~n38338;
  assign n38340 = ~n38320 & n38339;
  assign n38341 = ~pi0822 & ~n38340;
  assign n38342 = pi0822 & n38336;
  assign n38343 = ~n38320 & n38342;
  assign n38344 = ~n38338 & n38343;
  assign po0857 = n38341 | n38344;
  assign n38346 = ~n37479 & n37508;
  assign n38347 = ~n37486 & n38346;
  assign n38348 = ~n37567 & ~n38347;
  assign n38349 = ~n37486 & ~n37498;
  assign n38350 = ~n38124 & ~n38349;
  assign n38351 = n37479 & ~n38350;
  assign n38352 = n37486 & n37492;
  assign n38353 = n37507 & n38352;
  assign n38354 = ~n38351 & ~n38353;
  assign n38355 = n38348 & n38354;
  assign n38356 = n37473 & ~n38355;
  assign n38357 = ~n37551 & ~n37554;
  assign n38358 = ~n37486 & n37519;
  assign n38359 = n38357 & ~n38358;
  assign n38360 = ~n37479 & ~n38359;
  assign n38361 = n37508 & n37532;
  assign n38362 = ~n37513 & ~n38361;
  assign n38363 = ~n38360 & n38362;
  assign n38364 = ~n37566 & ~n37833;
  assign n38365 = n37479 & ~n38364;
  assign n38366 = n38363 & ~n38365;
  assign n38367 = ~n37473 & ~n38366;
  assign n38368 = ~n38356 & ~n38367;
  assign n38369 = ~n37486 & n37530;
  assign n38370 = n37486 & ~n37830;
  assign n38371 = ~n38369 & ~n38370;
  assign n38372 = n37479 & ~n38371;
  assign n38373 = ~n37551 & n38103;
  assign n38374 = n37556 & ~n38373;
  assign n38375 = ~n38372 & ~n38374;
  assign n38376 = n38368 & n38375;
  assign n38377 = ~pi0803 & ~n38376;
  assign n38378 = pi0803 & n38375;
  assign n38379 = ~n38367 & n38378;
  assign n38380 = ~n38356 & n38379;
  assign po0858 = n38377 | n38380;
  assign n38382 = ~n37001 & ~n37008;
  assign n38383 = ~n36973 & ~n38382;
  assign n38384 = ~n37063 & ~n38383;
  assign n38385 = ~n36985 & ~n36992;
  assign n38386 = n36973 & n38385;
  assign n38387 = n36979 & n38386;
  assign n38388 = ~n36973 & n37006;
  assign n38389 = n36979 & n38388;
  assign n38390 = ~n38313 & ~n38389;
  assign n38391 = n36992 & n38242;
  assign n38392 = n36979 & n37026;
  assign n38393 = ~n38391 & ~n38392;
  assign n38394 = ~n38385 & n38393;
  assign n38395 = n36973 & ~n38394;
  assign n38396 = ~n37004 & ~n38395;
  assign n38397 = n38390 & n38396;
  assign n38398 = ~n37039 & ~n38397;
  assign n38399 = ~n38387 & ~n38398;
  assign n38400 = ~n37027 & ~n37046;
  assign n38401 = ~n37056 & n38400;
  assign n38402 = ~n36973 & ~n38401;
  assign n38403 = n36999 & n38242;
  assign n38404 = ~n37030 & ~n38403;
  assign n38405 = n36973 & ~n38404;
  assign n38406 = ~n38402 & ~n38405;
  assign n38407 = ~n38323 & n38406;
  assign n38408 = ~n37016 & ~n37057;
  assign n38409 = n38407 & n38408;
  assign n38410 = n37039 & ~n38409;
  assign n38411 = n38399 & ~n38410;
  assign n38412 = n38384 & n38411;
  assign n38413 = ~pi0823 & ~n38412;
  assign n38414 = pi0823 & n38399;
  assign n38415 = n38384 & n38414;
  assign n38416 = ~n38410 & n38415;
  assign po0859 = n38413 | n38416;
  assign n38418 = n37386 & n37408;
  assign n38419 = ~n37995 & ~n38418;
  assign n38420 = ~n37392 & n38419;
  assign n38421 = ~n37386 & n37453;
  assign n38422 = ~n37380 & ~n37402;
  assign n38423 = n37401 & ~n38422;
  assign n38424 = n37386 & ~n37401;
  assign n38425 = n37373 & n38424;
  assign n38426 = ~n37386 & n37402;
  assign n38427 = ~n38425 & ~n38426;
  assign n38428 = n37392 & n38427;
  assign n38429 = ~n38423 & n38428;
  assign n38430 = ~n38421 & n38429;
  assign n38431 = ~n38420 & ~n38430;
  assign n38432 = ~n37386 & n38423;
  assign n38433 = ~n37993 & ~n38432;
  assign n38434 = ~n38431 & n38433;
  assign n38435 = n37367 & ~n38434;
  assign n38436 = ~n37392 & ~n38422;
  assign n38437 = n37386 & n38436;
  assign n38438 = ~n37386 & n37447;
  assign n38439 = ~n37424 & ~n38438;
  assign n38440 = ~n37392 & ~n38439;
  assign n38441 = ~n37401 & n38436;
  assign n38442 = ~n38440 & ~n38441;
  assign n38443 = ~n38437 & n38442;
  assign n38444 = ~n37367 & ~n38443;
  assign n38445 = ~n38435 & ~n38444;
  assign n38446 = n37392 & ~n38419;
  assign n38447 = ~n37406 & ~n38446;
  assign n38448 = ~n37367 & ~n38447;
  assign n38449 = ~n37392 & n37406;
  assign n38450 = n37392 & ~n38433;
  assign n38451 = ~n38449 & ~n38450;
  assign n38452 = ~n38448 & n38451;
  assign n38453 = n38445 & n38452;
  assign n38454 = pi0824 & ~n38453;
  assign n38455 = ~pi0824 & n38452;
  assign n38456 = ~n38444 & n38455;
  assign n38457 = ~n38435 & n38456;
  assign po0860 = n38454 | n38457;
  assign n38459 = ~n37392 & n37434;
  assign n38460 = ~n38422 & n38424;
  assign n38461 = ~n37448 & ~n38460;
  assign n38462 = ~n37993 & n38461;
  assign n38463 = n37392 & ~n38462;
  assign n38464 = ~n37386 & n37403;
  assign n38465 = ~n38463 & ~n38464;
  assign n38466 = ~n37401 & n37447;
  assign n38467 = n37386 & n37422;
  assign n38468 = ~n38466 & ~n38467;
  assign n38469 = ~n38426 & n38468;
  assign n38470 = ~n37392 & ~n38469;
  assign n38471 = n38465 & ~n38470;
  assign n38472 = n37367 & ~n38471;
  assign n38473 = ~n38459 & ~n38472;
  assign n38474 = n37386 & n37402;
  assign n38475 = ~n37992 & ~n38474;
  assign n38476 = ~n37392 & ~n38475;
  assign n38477 = ~n37449 & ~n38476;
  assign n38478 = ~n37424 & ~n37434;
  assign n38479 = ~n37386 & n37435;
  assign n38480 = ~n37422 & ~n38479;
  assign n38481 = ~n38466 & n38480;
  assign n38482 = n37392 & ~n38481;
  assign n38483 = n37386 & n37403;
  assign n38484 = ~n38482 & ~n38483;
  assign n38485 = n38478 & n38484;
  assign n38486 = n38477 & n38485;
  assign n38487 = ~n37367 & ~n38486;
  assign n38488 = ~n37441 & ~n38421;
  assign n38489 = n37392 & ~n38488;
  assign n38490 = ~n38487 & ~n38489;
  assign n38491 = n38473 & n38490;
  assign n38492 = pi0829 & n38491;
  assign n38493 = ~pi0829 & ~n38491;
  assign po0861 = n38492 | n38493;
  assign n38495 = pi3666 & pi9040;
  assign n38496 = pi3700 & ~pi9040;
  assign n38497 = ~n38495 & ~n38496;
  assign n38498 = ~pi0794 & n38497;
  assign n38499 = pi0794 & ~n38497;
  assign n38500 = ~n38498 & ~n38499;
  assign n38501 = pi3693 & pi9040;
  assign n38502 = pi3696 & ~pi9040;
  assign n38503 = ~n38501 & ~n38502;
  assign n38504 = ~pi0782 & n38503;
  assign n38505 = pi0782 & ~n38503;
  assign n38506 = ~n38504 & ~n38505;
  assign n38507 = ~n38500 & ~n38506;
  assign n38508 = pi3691 & pi9040;
  assign n38509 = pi3660 & ~pi9040;
  assign n38510 = ~n38508 & ~n38509;
  assign n38511 = pi0791 & n38510;
  assign n38512 = ~pi0791 & ~n38510;
  assign n38513 = ~n38511 & ~n38512;
  assign n38514 = pi3661 & pi9040;
  assign n38515 = pi3693 & ~pi9040;
  assign n38516 = ~n38514 & ~n38515;
  assign n38517 = pi0793 & n38516;
  assign n38518 = ~pi0793 & ~n38516;
  assign n38519 = ~n38517 & ~n38518;
  assign n38520 = n38506 & ~n38519;
  assign n38521 = n38513 & n38520;
  assign n38522 = ~n38507 & ~n38521;
  assign n38523 = pi3659 & ~pi9040;
  assign n38524 = pi3679 & pi9040;
  assign n38525 = ~n38523 & ~n38524;
  assign n38526 = ~pi0772 & n38525;
  assign n38527 = pi0772 & ~n38525;
  assign n38528 = ~n38526 & ~n38527;
  assign n38529 = pi3665 & pi9040;
  assign n38530 = pi3691 & ~pi9040;
  assign n38531 = ~n38529 & ~n38530;
  assign n38532 = pi0776 & n38531;
  assign n38533 = ~pi0776 & ~n38531;
  assign n38534 = ~n38532 & ~n38533;
  assign n38535 = ~n38528 & ~n38534;
  assign n38536 = ~n38522 & n38535;
  assign n38537 = ~n38506 & n38519;
  assign n38538 = ~n38500 & n38513;
  assign n38539 = ~n38537 & n38538;
  assign n38540 = ~n38528 & n38539;
  assign n38541 = ~n38500 & ~n38513;
  assign n38542 = n38534 & n38541;
  assign n38543 = n38537 & n38542;
  assign n38544 = ~n38500 & ~n38534;
  assign n38545 = n38513 & n38544;
  assign n38546 = ~n38519 & n38545;
  assign n38547 = ~n38543 & ~n38546;
  assign n38548 = ~n38540 & n38547;
  assign n38549 = ~n38500 & n38520;
  assign n38550 = n38506 & n38519;
  assign n38551 = n38500 & n38550;
  assign n38552 = ~n38549 & ~n38551;
  assign n38553 = n38534 & ~n38552;
  assign n38554 = ~n38506 & ~n38519;
  assign n38555 = n38500 & n38534;
  assign n38556 = n38554 & n38555;
  assign n38557 = ~n38513 & n38556;
  assign n38558 = ~n38553 & ~n38557;
  assign n38559 = ~n38528 & ~n38558;
  assign n38560 = n38500 & ~n38513;
  assign n38561 = ~n38520 & ~n38537;
  assign n38562 = n38560 & ~n38561;
  assign n38563 = ~n38506 & ~n38513;
  assign n38564 = ~n38537 & ~n38563;
  assign n38565 = n38500 & ~n38564;
  assign n38566 = n38513 & n38550;
  assign n38567 = ~n38565 & ~n38566;
  assign n38568 = ~n38534 & ~n38567;
  assign n38569 = ~n38562 & ~n38568;
  assign n38570 = ~n38513 & n38550;
  assign n38571 = ~n38500 & n38570;
  assign n38572 = n38500 & n38513;
  assign n38573 = ~n38519 & n38572;
  assign n38574 = ~n38500 & ~n38564;
  assign n38575 = ~n38573 & ~n38574;
  assign n38576 = n38534 & ~n38575;
  assign n38577 = ~n38571 & ~n38576;
  assign n38578 = n38569 & n38577;
  assign n38579 = n38528 & ~n38578;
  assign n38580 = ~n38559 & ~n38579;
  assign n38581 = n38548 & n38580;
  assign n38582 = ~n38536 & n38581;
  assign n38583 = pi0825 & ~n38582;
  assign n38584 = ~pi0825 & n38548;
  assign n38585 = ~n38536 & n38584;
  assign n38586 = n38580 & n38585;
  assign po0862 = n38583 | n38586;
  assign n38588 = ~n38513 & n38554;
  assign n38589 = n38513 & n38537;
  assign n38590 = ~n38588 & ~n38589;
  assign n38591 = n38519 & n38572;
  assign n38592 = n38590 & ~n38591;
  assign n38593 = n38535 & ~n38592;
  assign n38594 = n38521 & ~n38528;
  assign n38595 = ~n38500 & n38594;
  assign n38596 = n38513 & n38554;
  assign n38597 = n38534 & n38596;
  assign n38598 = ~n38513 & n38519;
  assign n38599 = ~n38500 & n38550;
  assign n38600 = ~n38598 & ~n38599;
  assign n38601 = n38534 & ~n38600;
  assign n38602 = ~n38597 & ~n38601;
  assign n38603 = ~n38528 & ~n38602;
  assign n38604 = ~n38595 & ~n38603;
  assign n38605 = n38519 & n38541;
  assign n38606 = ~n38519 & n38560;
  assign n38607 = n38506 & n38606;
  assign n38608 = ~n38605 & ~n38607;
  assign n38609 = n38534 & ~n38608;
  assign n38610 = n38604 & ~n38609;
  assign n38611 = n38544 & n38550;
  assign n38612 = n38513 & n38611;
  assign n38613 = ~n38561 & n38572;
  assign n38614 = n38500 & n38588;
  assign n38615 = ~n38613 & ~n38614;
  assign n38616 = n38500 & ~n38534;
  assign n38617 = n38570 & n38616;
  assign n38618 = n38541 & ~n38561;
  assign n38619 = ~n38500 & n38596;
  assign n38620 = ~n38618 & ~n38619;
  assign n38621 = ~n38617 & n38620;
  assign n38622 = n38615 & n38621;
  assign n38623 = ~n38612 & n38622;
  assign n38624 = n38513 & n38555;
  assign n38625 = n38506 & n38624;
  assign n38626 = n38623 & ~n38625;
  assign n38627 = n38528 & ~n38626;
  assign n38628 = n38610 & ~n38627;
  assign n38629 = ~n38593 & n38628;
  assign n38630 = ~pi0831 & ~n38629;
  assign n38631 = pi0831 & n38610;
  assign n38632 = ~n38593 & n38631;
  assign n38633 = ~n38627 & n38632;
  assign po0863 = n38630 | n38633;
  assign n38635 = ~n38513 & n38537;
  assign n38636 = ~n38566 & ~n38635;
  assign n38637 = n38534 & ~n38636;
  assign n38638 = n38500 & n38520;
  assign n38639 = ~n38589 & ~n38638;
  assign n38640 = ~n38570 & n38639;
  assign n38641 = ~n38534 & ~n38640;
  assign n38642 = ~n38637 & ~n38641;
  assign n38643 = ~n38597 & ~n38607;
  assign n38644 = n38642 & n38643;
  assign n38645 = n38528 & ~n38644;
  assign n38646 = n38513 & n38534;
  assign n38647 = ~n38519 & n38646;
  assign n38648 = n38506 & n38647;
  assign n38649 = n38590 & ~n38648;
  assign n38650 = ~n38570 & n38649;
  assign n38651 = n38500 & ~n38650;
  assign n38652 = ~n38500 & n38566;
  assign n38653 = n38500 & n38554;
  assign n38654 = ~n38549 & ~n38653;
  assign n38655 = ~n38534 & ~n38654;
  assign n38656 = ~n38652 & ~n38655;
  assign n38657 = ~n38651 & n38656;
  assign n38658 = ~n38528 & ~n38657;
  assign n38659 = ~n38645 & ~n38658;
  assign n38660 = ~n38513 & n38549;
  assign n38661 = ~n38619 & ~n38660;
  assign n38662 = n38534 & ~n38661;
  assign n38663 = n38544 & n38563;
  assign n38664 = ~n38662 & ~n38663;
  assign n38665 = n38659 & n38664;
  assign n38666 = ~pi0816 & ~n38665;
  assign n38667 = pi0816 & ~n38662;
  assign n38668 = n38659 & n38667;
  assign n38669 = ~n38663 & n38668;
  assign po0864 = n38666 | n38669;
  assign n38671 = n38534 & n38566;
  assign n38672 = n38500 & n38671;
  assign n38673 = ~n38557 & ~n38672;
  assign n38674 = ~n38614 & ~n38617;
  assign n38675 = n38507 & n38513;
  assign n38676 = ~n38599 & ~n38675;
  assign n38677 = n38534 & ~n38676;
  assign n38678 = ~n38534 & ~n38560;
  assign n38679 = ~n38561 & n38678;
  assign n38680 = ~n38513 & ~n38550;
  assign n38681 = n38534 & n38680;
  assign n38682 = n38500 & n38681;
  assign n38683 = ~n38679 & ~n38682;
  assign n38684 = ~n38677 & n38683;
  assign n38685 = n38674 & n38684;
  assign n38686 = ~n38528 & ~n38685;
  assign n38687 = n38673 & ~n38686;
  assign n38688 = ~n38534 & n38589;
  assign n38689 = ~n38500 & n38688;
  assign n38690 = n38528 & ~n38534;
  assign n38691 = ~n38562 & ~n38599;
  assign n38692 = ~n38596 & n38691;
  assign n38693 = n38690 & ~n38692;
  assign n38694 = ~n38500 & n38588;
  assign n38695 = n38507 & ~n38513;
  assign n38696 = ~n38549 & ~n38695;
  assign n38697 = ~n38521 & ~n38551;
  assign n38698 = n38696 & n38697;
  assign n38699 = n38534 & ~n38698;
  assign n38700 = ~n38694 & ~n38699;
  assign n38701 = n38528 & ~n38700;
  assign n38702 = ~n38693 & ~n38701;
  assign n38703 = ~n38689 & n38702;
  assign n38704 = n38687 & n38703;
  assign n38705 = pi0832 & ~n38704;
  assign n38706 = ~pi0832 & n38687;
  assign n38707 = n38703 & n38706;
  assign po0865 = n38705 | n38707;
  assign n38709 = pi3725 & pi9040;
  assign n38710 = pi3735 & ~pi9040;
  assign n38711 = ~n38709 & ~n38710;
  assign n38712 = pi0838 & n38711;
  assign n38713 = ~pi0838 & ~n38711;
  assign n38714 = ~n38712 & ~n38713;
  assign n38715 = pi3738 & pi9040;
  assign n38716 = pi3712 & ~pi9040;
  assign n38717 = ~n38715 & ~n38716;
  assign n38718 = ~pi0850 & ~n38717;
  assign n38719 = pi0850 & ~n38715;
  assign n38720 = ~n38716 & n38719;
  assign n38721 = ~n38718 & ~n38720;
  assign n38722 = pi3717 & pi9040;
  assign n38723 = pi3750 & ~pi9040;
  assign n38724 = ~n38722 & ~n38723;
  assign n38725 = ~pi0835 & n38724;
  assign n38726 = pi0835 & ~n38724;
  assign n38727 = ~n38725 & ~n38726;
  assign n38728 = ~n38721 & n38727;
  assign n38729 = pi3768 & pi9040;
  assign n38730 = pi3722 & ~pi9040;
  assign n38731 = ~n38729 & ~n38730;
  assign n38732 = ~pi0828 & ~n38731;
  assign n38733 = pi0828 & ~n38729;
  assign n38734 = ~n38730 & n38733;
  assign n38735 = ~n38732 & ~n38734;
  assign n38736 = pi3716 & pi9040;
  assign n38737 = pi3774 & ~pi9040;
  assign n38738 = ~n38736 & ~n38737;
  assign n38739 = pi0854 & n38738;
  assign n38740 = ~pi0854 & ~n38738;
  assign n38741 = ~n38739 & ~n38740;
  assign n38742 = n38735 & n38741;
  assign n38743 = n38728 & n38742;
  assign n38744 = n38721 & n38727;
  assign n38745 = ~n38735 & n38744;
  assign n38746 = n38741 & n38745;
  assign n38747 = ~n38743 & ~n38746;
  assign n38748 = n38721 & ~n38727;
  assign n38749 = ~n38735 & n38748;
  assign n38750 = ~n38741 & n38749;
  assign n38751 = n38728 & ~n38741;
  assign n38752 = ~n38735 & n38751;
  assign n38753 = ~n38750 & ~n38752;
  assign n38754 = n38747 & n38753;
  assign n38755 = n38714 & ~n38754;
  assign n38756 = ~n38727 & ~n38735;
  assign n38757 = pi3750 & pi9040;
  assign n38758 = pi3769 & ~pi9040;
  assign n38759 = ~n38757 & ~n38758;
  assign n38760 = ~pi0863 & ~n38759;
  assign n38761 = pi0863 & n38759;
  assign n38762 = ~n38760 & ~n38761;
  assign n38763 = ~n38714 & n38741;
  assign n38764 = n38762 & n38763;
  assign n38765 = n38756 & n38764;
  assign n38766 = ~n38735 & ~n38741;
  assign n38767 = n38727 & n38766;
  assign n38768 = ~n38714 & ~n38767;
  assign n38769 = ~n38721 & n38742;
  assign n38770 = ~n38748 & ~n38756;
  assign n38771 = ~n38741 & ~n38770;
  assign n38772 = n38728 & n38735;
  assign n38773 = ~n38771 & ~n38772;
  assign n38774 = n38714 & n38773;
  assign n38775 = ~n38769 & n38774;
  assign n38776 = ~n38768 & ~n38775;
  assign n38777 = n38735 & n38744;
  assign n38778 = n38741 & n38777;
  assign n38779 = ~n38776 & ~n38778;
  assign n38780 = n38762 & ~n38779;
  assign n38781 = ~n38765 & ~n38780;
  assign n38782 = ~n38721 & n38741;
  assign n38783 = ~n38727 & n38782;
  assign n38784 = ~n38735 & n38783;
  assign n38785 = ~n38745 & ~n38784;
  assign n38786 = n38714 & ~n38785;
  assign n38787 = ~n38727 & ~n38741;
  assign n38788 = ~n38714 & n38787;
  assign n38789 = n38721 & n38735;
  assign n38790 = n38728 & n38741;
  assign n38791 = ~n38789 & ~n38790;
  assign n38792 = ~n38714 & ~n38791;
  assign n38793 = ~n38788 & ~n38792;
  assign n38794 = ~n38721 & ~n38727;
  assign n38795 = n38735 & n38794;
  assign n38796 = ~n38741 & n38795;
  assign n38797 = n38793 & ~n38796;
  assign n38798 = ~n38727 & n38789;
  assign n38799 = n38741 & n38798;
  assign n38800 = n38797 & ~n38799;
  assign n38801 = ~n38786 & n38800;
  assign n38802 = ~n38762 & ~n38801;
  assign n38803 = n38781 & ~n38802;
  assign n38804 = ~n38755 & n38803;
  assign n38805 = ~n38714 & n38796;
  assign n38806 = n38804 & ~n38805;
  assign n38807 = pi0866 & ~n38806;
  assign n38808 = ~pi0866 & ~n38805;
  assign n38809 = ~n38802 & n38808;
  assign n38810 = n38781 & n38809;
  assign n38811 = ~n38755 & n38810;
  assign po0875 = n38807 | n38811;
  assign n38813 = pi3773 & pi9040;
  assign n38814 = pi3716 & ~pi9040;
  assign n38815 = ~n38813 & ~n38814;
  assign n38816 = pi0844 & n38815;
  assign n38817 = ~pi0844 & ~n38815;
  assign n38818 = ~n38816 & ~n38817;
  assign n38819 = pi3766 & pi9040;
  assign n38820 = pi3773 & ~pi9040;
  assign n38821 = ~n38819 & ~n38820;
  assign n38822 = ~pi0852 & n38821;
  assign n38823 = pi0852 & ~n38821;
  assign n38824 = ~n38822 & ~n38823;
  assign n38825 = pi3749 & pi9040;
  assign n38826 = pi3738 & ~pi9040;
  assign n38827 = ~n38825 & ~n38826;
  assign n38828 = ~pi0837 & ~n38827;
  assign n38829 = pi0837 & ~n38825;
  assign n38830 = ~n38826 & n38829;
  assign n38831 = ~n38828 & ~n38830;
  assign n38832 = pi3722 & pi9040;
  assign n38833 = pi3725 & ~pi9040;
  assign n38834 = ~n38832 & ~n38833;
  assign n38835 = ~pi0828 & n38834;
  assign n38836 = pi0828 & ~n38834;
  assign n38837 = ~n38835 & ~n38836;
  assign n38838 = ~n38831 & n38837;
  assign n38839 = ~n38824 & n38838;
  assign n38840 = ~n38818 & n38839;
  assign n38841 = pi3754 & pi9040;
  assign n38842 = pi3743 & ~pi9040;
  assign n38843 = ~n38841 & ~n38842;
  assign n38844 = pi0859 & n38843;
  assign n38845 = ~pi0859 & ~n38843;
  assign n38846 = ~n38844 & ~n38845;
  assign n38847 = n38831 & ~n38846;
  assign n38848 = ~n38818 & n38847;
  assign n38849 = n38831 & n38846;
  assign n38850 = n38818 & n38849;
  assign n38851 = ~n38848 & ~n38850;
  assign n38852 = n38824 & ~n38851;
  assign n38853 = ~n38837 & ~n38846;
  assign n38854 = ~n38831 & n38853;
  assign n38855 = n38818 & n38854;
  assign n38856 = n38837 & n38846;
  assign n38857 = ~n38831 & n38856;
  assign n38858 = n38837 & ~n38846;
  assign n38859 = n38831 & n38858;
  assign n38860 = n38818 & n38859;
  assign n38861 = ~n38857 & ~n38860;
  assign n38862 = ~n38855 & n38861;
  assign n38863 = ~n38824 & ~n38862;
  assign n38864 = ~n38852 & ~n38863;
  assign n38865 = ~n38818 & ~n38831;
  assign n38866 = ~n38837 & n38865;
  assign n38867 = n38846 & n38866;
  assign n38868 = n38831 & n38853;
  assign n38869 = ~n38867 & ~n38868;
  assign n38870 = n38824 & ~n38869;
  assign n38871 = n38837 & n38865;
  assign n38872 = ~n38846 & n38871;
  assign n38873 = ~n38855 & ~n38872;
  assign n38874 = n38818 & ~n38831;
  assign n38875 = n38846 & n38874;
  assign n38876 = ~n38837 & n38846;
  assign n38877 = n38831 & n38876;
  assign n38878 = ~n38818 & n38877;
  assign n38879 = ~n38875 & ~n38878;
  assign n38880 = ~n38824 & ~n38879;
  assign n38881 = n38873 & ~n38880;
  assign n38882 = ~n38870 & n38881;
  assign n38883 = pi3726 & pi9040;
  assign n38884 = pi3758 & ~pi9040;
  assign n38885 = ~n38883 & ~n38884;
  assign n38886 = pi0835 & n38885;
  assign n38887 = ~pi0835 & ~n38885;
  assign n38888 = ~n38886 & ~n38887;
  assign n38889 = ~n38882 & n38888;
  assign n38890 = ~n38818 & n38824;
  assign n38891 = n38853 & n38890;
  assign n38892 = n38831 & n38856;
  assign n38893 = n38837 & n38874;
  assign n38894 = ~n38846 & n38893;
  assign n38895 = ~n38892 & ~n38894;
  assign n38896 = n38818 & n38876;
  assign n38897 = n38895 & ~n38896;
  assign n38898 = n38824 & ~n38897;
  assign n38899 = ~n38891 & ~n38898;
  assign n38900 = n38818 & n38877;
  assign n38901 = ~n38818 & n38868;
  assign n38902 = ~n38831 & n38846;
  assign n38903 = ~n38818 & ~n38824;
  assign n38904 = n38902 & n38903;
  assign n38905 = ~n38818 & n38857;
  assign n38906 = ~n38904 & ~n38905;
  assign n38907 = ~n38901 & n38906;
  assign n38908 = ~n38900 & n38907;
  assign n38909 = n38899 & n38908;
  assign n38910 = ~n38888 & ~n38909;
  assign n38911 = ~n38889 & ~n38910;
  assign n38912 = n38864 & n38911;
  assign n38913 = ~n38840 & n38912;
  assign n38914 = ~pi0884 & ~n38913;
  assign n38915 = pi0884 & n38913;
  assign po0892 = n38914 | n38915;
  assign n38917 = pi3715 & pi9040;
  assign n38918 = pi3746 & ~pi9040;
  assign n38919 = ~n38917 & ~n38918;
  assign n38920 = ~pi0837 & ~n38919;
  assign n38921 = pi0837 & ~n38917;
  assign n38922 = ~n38918 & n38921;
  assign n38923 = ~n38920 & ~n38922;
  assign n38924 = pi3769 & pi9040;
  assign n38925 = pi3747 & ~pi9040;
  assign n38926 = ~n38924 & ~n38925;
  assign n38927 = ~pi0851 & n38926;
  assign n38928 = pi0851 & ~n38926;
  assign n38929 = ~n38927 & ~n38928;
  assign n38930 = pi3747 & pi9040;
  assign n38931 = pi3726 & ~pi9040;
  assign n38932 = ~n38930 & ~n38931;
  assign n38933 = pi0834 & n38932;
  assign n38934 = ~pi0834 & ~n38932;
  assign n38935 = ~n38933 & ~n38934;
  assign n38936 = pi3758 & pi9040;
  assign n38937 = pi3766 & ~pi9040;
  assign n38938 = ~n38936 & ~n38937;
  assign n38939 = ~pi0856 & n38938;
  assign n38940 = pi0856 & ~n38938;
  assign n38941 = ~n38939 & ~n38940;
  assign n38942 = ~n38935 & ~n38941;
  assign n38943 = ~n38929 & n38942;
  assign n38944 = n38923 & n38943;
  assign n38945 = pi3733 & pi9040;
  assign n38946 = pi3714 & ~pi9040;
  assign n38947 = ~n38945 & ~n38946;
  assign n38948 = pi0840 & n38947;
  assign n38949 = ~pi0840 & ~n38947;
  assign n38950 = ~n38948 & ~n38949;
  assign n38951 = ~n38923 & n38950;
  assign n38952 = n38929 & n38951;
  assign n38953 = ~n38935 & n38952;
  assign n38954 = ~n38944 & ~n38953;
  assign n38955 = ~n38923 & ~n38950;
  assign n38956 = n38929 & n38955;
  assign n38957 = n38923 & n38950;
  assign n38958 = ~n38955 & ~n38957;
  assign n38959 = n38935 & ~n38958;
  assign n38960 = ~n38956 & ~n38959;
  assign n38961 = n38941 & ~n38960;
  assign n38962 = ~n38929 & ~n38950;
  assign n38963 = ~n38935 & n38962;
  assign n38964 = n38923 & ~n38950;
  assign n38965 = ~n38929 & n38964;
  assign n38966 = ~n38963 & ~n38965;
  assign n38967 = ~n38929 & n38951;
  assign n38968 = n38935 & n38967;
  assign n38969 = n38966 & ~n38968;
  assign n38970 = ~n38941 & ~n38969;
  assign n38971 = ~n38961 & ~n38970;
  assign n38972 = ~n38935 & n38941;
  assign n38973 = n38951 & n38972;
  assign n38974 = n38935 & n38956;
  assign n38975 = n38929 & n38950;
  assign n38976 = n38923 & n38975;
  assign n38977 = n38935 & n38976;
  assign n38978 = ~n38974 & ~n38977;
  assign n38979 = n38929 & ~n38935;
  assign n38980 = n38923 & n38979;
  assign n38981 = ~n38950 & n38980;
  assign n38982 = n38978 & ~n38981;
  assign n38983 = ~n38973 & n38982;
  assign n38984 = n38971 & n38983;
  assign n38985 = pi3754 & ~pi9040;
  assign n38986 = pi3774 & pi9040;
  assign n38987 = ~n38985 & ~n38986;
  assign n38988 = ~pi0859 & ~n38987;
  assign n38989 = pi0859 & n38987;
  assign n38990 = ~n38988 & ~n38989;
  assign n38991 = ~n38984 & n38990;
  assign n38992 = n38941 & ~n38990;
  assign n38993 = ~n38935 & n38957;
  assign n38994 = ~n38968 & ~n38993;
  assign n38995 = ~n38963 & n38994;
  assign n38996 = n38992 & ~n38995;
  assign n38997 = ~n38923 & n38979;
  assign n38998 = ~n38929 & n38955;
  assign n38999 = n38935 & n38998;
  assign n39000 = ~n38997 & ~n38999;
  assign n39001 = ~n38929 & n38957;
  assign n39002 = ~n38952 & ~n39001;
  assign n39003 = n39000 & n39002;
  assign n39004 = ~n38941 & ~n39003;
  assign n39005 = n38929 & n38964;
  assign n39006 = n38935 & n39005;
  assign n39007 = ~n39004 & ~n39006;
  assign n39008 = ~n38990 & ~n39007;
  assign n39009 = ~n38996 & ~n39008;
  assign n39010 = ~n38991 & n39009;
  assign n39011 = n38954 & n39010;
  assign n39012 = pi0869 & ~n39011;
  assign n39013 = ~pi0869 & n38954;
  assign n39014 = n39009 & n39013;
  assign n39015 = ~n38991 & n39014;
  assign po0896 = n39012 | n39015;
  assign n39017 = pi3740 & pi9040;
  assign n39018 = pi3737 & ~pi9040;
  assign n39019 = ~n39017 & ~n39018;
  assign n39020 = ~pi0860 & n39019;
  assign n39021 = pi0860 & ~n39019;
  assign n39022 = ~n39020 & ~n39021;
  assign n39023 = pi3728 & pi9040;
  assign n39024 = pi3729 & ~pi9040;
  assign n39025 = ~n39023 & ~n39024;
  assign n39026 = ~pi0819 & n39025;
  assign n39027 = pi0819 & ~n39025;
  assign n39028 = ~n39026 & ~n39027;
  assign n39029 = pi3741 & pi9040;
  assign n39030 = pi3723 & ~pi9040;
  assign n39031 = ~n39029 & ~n39030;
  assign n39032 = ~pi0850 & ~n39031;
  assign n39033 = pi0850 & n39031;
  assign n39034 = ~n39032 & ~n39033;
  assign n39035 = pi3736 & ~pi9040;
  assign n39036 = pi3711 & pi9040;
  assign n39037 = ~n39035 & ~n39036;
  assign n39038 = pi0841 & n39037;
  assign n39039 = ~pi0841 & ~n39037;
  assign n39040 = ~n39038 & ~n39039;
  assign n39041 = n39034 & ~n39040;
  assign n39042 = n39028 & n39041;
  assign n39043 = pi3721 & pi9040;
  assign n39044 = pi3772 & ~pi9040;
  assign n39045 = ~n39043 & ~n39044;
  assign n39046 = pi0863 & n39045;
  assign n39047 = ~pi0863 & ~n39045;
  assign n39048 = ~n39046 & ~n39047;
  assign n39049 = n39034 & n39048;
  assign n39050 = ~n39028 & n39049;
  assign n39051 = n39040 & n39050;
  assign n39052 = ~n39042 & ~n39051;
  assign n39053 = ~n39028 & ~n39048;
  assign n39054 = ~n39034 & n39053;
  assign n39055 = n39040 & n39054;
  assign n39056 = n39052 & ~n39055;
  assign n39057 = n39022 & ~n39056;
  assign n39058 = pi3775 & pi9040;
  assign n39059 = pi3718 & ~pi9040;
  assign n39060 = ~n39058 & ~n39059;
  assign n39061 = ~pi0842 & ~n39060;
  assign n39062 = pi0842 & n39060;
  assign n39063 = ~n39061 & ~n39062;
  assign n39064 = ~n39022 & n39040;
  assign n39065 = n39053 & n39064;
  assign n39066 = n39034 & n39065;
  assign n39067 = ~n39022 & ~n39040;
  assign n39068 = ~n39028 & n39048;
  assign n39069 = n39067 & n39068;
  assign n39070 = n39028 & n39048;
  assign n39071 = n39034 & n39070;
  assign n39072 = ~n39022 & n39071;
  assign n39073 = n39040 & n39072;
  assign n39074 = n39042 & ~n39048;
  assign n39075 = ~n39073 & ~n39074;
  assign n39076 = ~n39069 & n39075;
  assign n39077 = ~n39066 & n39076;
  assign n39078 = ~n39034 & ~n39040;
  assign n39079 = ~n39028 & n39078;
  assign n39080 = n39048 & n39079;
  assign n39081 = n39077 & ~n39080;
  assign n39082 = ~n39063 & ~n39081;
  assign n39083 = n39028 & ~n39034;
  assign n39084 = n39048 & n39083;
  assign n39085 = n39022 & n39084;
  assign n39086 = n39040 & n39085;
  assign n39087 = n39041 & ~n39048;
  assign n39088 = n39028 & ~n39048;
  assign n39089 = ~n39040 & n39088;
  assign n39090 = ~n39087 & ~n39089;
  assign n39091 = n39022 & ~n39090;
  assign n39092 = ~n39086 & ~n39091;
  assign n39093 = ~n39063 & ~n39092;
  assign n39094 = ~n39082 & ~n39093;
  assign n39095 = ~n39057 & n39094;
  assign n39096 = ~n39034 & n39040;
  assign n39097 = ~n39022 & n39096;
  assign n39098 = n39088 & n39097;
  assign n39099 = ~n39034 & n39048;
  assign n39100 = n39067 & n39099;
  assign n39101 = n39022 & n39049;
  assign n39102 = n39040 & ~n39048;
  assign n39103 = ~n39034 & n39102;
  assign n39104 = ~n39054 & ~n39103;
  assign n39105 = ~n39101 & n39104;
  assign n39106 = ~n39040 & n39084;
  assign n39107 = n39105 & ~n39106;
  assign n39108 = ~n39022 & n39053;
  assign n39109 = ~n39040 & n39108;
  assign n39110 = ~n39028 & ~n39034;
  assign n39111 = n39040 & n39088;
  assign n39112 = ~n39110 & ~n39111;
  assign n39113 = ~n39022 & ~n39112;
  assign n39114 = ~n39109 & ~n39113;
  assign n39115 = n39107 & n39114;
  assign n39116 = n39063 & ~n39115;
  assign n39117 = ~n39100 & ~n39116;
  assign n39118 = ~n39098 & n39117;
  assign n39119 = n39095 & n39118;
  assign n39120 = pi0867 & n39119;
  assign n39121 = ~pi0867 & ~n39119;
  assign po0901 = n39120 | n39121;
  assign n39123 = n38846 & n38893;
  assign n39124 = ~n38849 & ~n38872;
  assign n39125 = ~n38824 & ~n39124;
  assign n39126 = ~n39123 & ~n39125;
  assign n39127 = ~n38867 & n39126;
  assign n39128 = n38818 & n38824;
  assign n39129 = n38854 & n39128;
  assign n39130 = ~n38901 & ~n39129;
  assign n39131 = ~n38860 & n39130;
  assign n39132 = n39127 & n39131;
  assign n39133 = n38888 & ~n39132;
  assign n39134 = ~n38831 & n38876;
  assign n39135 = n38818 & n39134;
  assign n39136 = ~n38894 & ~n39135;
  assign n39137 = ~n38818 & n38859;
  assign n39138 = ~n38905 & ~n39137;
  assign n39139 = ~n38824 & n38854;
  assign n39140 = n38818 & n38868;
  assign n39141 = ~n39139 & ~n39140;
  assign n39142 = n38831 & ~n38837;
  assign n39143 = n38818 & n38846;
  assign n39144 = ~n39142 & ~n39143;
  assign n39145 = ~n38838 & n39144;
  assign n39146 = n38824 & ~n39145;
  assign n39147 = n39141 & ~n39146;
  assign n39148 = n39138 & n39147;
  assign n39149 = n39136 & n39148;
  assign n39150 = ~n38888 & ~n39149;
  assign n39151 = ~n39133 & ~n39150;
  assign n39152 = pi0879 & ~n39151;
  assign n39153 = ~pi0879 & ~n39133;
  assign n39154 = ~n39150 & n39153;
  assign po0902 = n39152 | n39154;
  assign n39156 = ~n38741 & n38798;
  assign n39157 = n38741 & n38756;
  assign n39158 = ~n38795 & ~n39157;
  assign n39159 = n38714 & ~n39158;
  assign n39160 = ~n39156 & ~n39159;
  assign n39161 = ~n38714 & ~n38741;
  assign n39162 = ~n38727 & n39161;
  assign n39163 = n38721 & n39162;
  assign n39164 = n38744 & n38763;
  assign n39165 = ~n39163 & ~n39164;
  assign n39166 = ~n38714 & n38772;
  assign n39167 = n39165 & ~n39166;
  assign n39168 = ~n38752 & ~n38784;
  assign n39169 = n38727 & n38742;
  assign n39170 = n39168 & ~n39169;
  assign n39171 = n39167 & n39170;
  assign n39172 = n39160 & n39171;
  assign n39173 = ~n38762 & ~n39172;
  assign n39174 = n38728 & ~n38735;
  assign n39175 = ~n38795 & ~n39174;
  assign n39176 = n38741 & ~n39175;
  assign n39177 = n38721 & n38766;
  assign n39178 = ~n38777 & ~n39177;
  assign n39179 = ~n38727 & n38735;
  assign n39180 = n38741 & n39179;
  assign n39181 = n39178 & ~n39180;
  assign n39182 = n38714 & ~n39181;
  assign n39183 = ~n38741 & n38794;
  assign n39184 = ~n38735 & n38741;
  assign n39185 = ~n38727 & n39184;
  assign n39186 = n38721 & n39185;
  assign n39187 = ~n39183 & ~n39186;
  assign n39188 = ~n38714 & ~n39187;
  assign n39189 = ~n38741 & n38745;
  assign n39190 = ~n39188 & ~n39189;
  assign n39191 = ~n39182 & n39190;
  assign n39192 = ~n39176 & n39191;
  assign n39193 = n38762 & ~n39192;
  assign n39194 = n38714 & n38767;
  assign n39195 = ~n39193 & ~n39194;
  assign n39196 = n38789 & n39161;
  assign n39197 = ~n38727 & n39196;
  assign n39198 = n39195 & ~n39197;
  assign n39199 = ~n39173 & n39198;
  assign n39200 = ~pi0889 & ~n39199;
  assign n39201 = pi0889 & n39195;
  assign n39202 = ~n39173 & n39201;
  assign n39203 = ~n39197 & n39202;
  assign po0903 = n39200 | n39203;
  assign n39205 = pi3732 & pi9040;
  assign n39206 = pi3741 & ~pi9040;
  assign n39207 = ~n39205 & ~n39206;
  assign n39208 = ~pi0853 & n39207;
  assign n39209 = pi0853 & ~n39207;
  assign n39210 = ~n39208 & ~n39209;
  assign n39211 = pi3777 & pi9040;
  assign n39212 = pi3721 & ~pi9040;
  assign n39213 = ~n39211 & ~n39212;
  assign n39214 = pi0842 & n39213;
  assign n39215 = ~pi0842 & ~n39213;
  assign n39216 = ~n39214 & ~n39215;
  assign n39217 = pi3756 & pi9040;
  assign n39218 = pi3713 & ~pi9040;
  assign n39219 = ~n39217 & ~n39218;
  assign n39220 = pi0861 & n39219;
  assign n39221 = ~pi0861 & ~n39219;
  assign n39222 = ~n39220 & ~n39221;
  assign n39223 = n39216 & ~n39222;
  assign n39224 = pi3739 & pi9040;
  assign n39225 = pi3734 & ~pi9040;
  assign n39226 = ~n39224 & ~n39225;
  assign n39227 = pi0857 & n39226;
  assign n39228 = ~pi0857 & ~n39226;
  assign n39229 = ~n39227 & ~n39228;
  assign n39230 = pi3723 & pi9040;
  assign n39231 = pi3711 & ~pi9040;
  assign n39232 = ~n39230 & ~n39231;
  assign n39233 = ~pi0819 & n39232;
  assign n39234 = pi0819 & ~n39232;
  assign n39235 = ~n39233 & ~n39234;
  assign n39236 = n39229 & ~n39235;
  assign n39237 = n39223 & n39236;
  assign n39238 = n39229 & n39235;
  assign n39239 = ~n39216 & n39238;
  assign n39240 = ~n39237 & ~n39239;
  assign n39241 = n39210 & ~n39240;
  assign n39242 = pi3713 & pi9040;
  assign n39243 = pi3730 & ~pi9040;
  assign n39244 = ~n39242 & ~n39243;
  assign n39245 = ~pi0845 & ~n39244;
  assign n39246 = pi0845 & n39244;
  assign n39247 = ~n39245 & ~n39246;
  assign n39248 = ~n39210 & ~n39229;
  assign n39249 = n39216 & n39248;
  assign n39250 = n39223 & n39235;
  assign n39251 = n39216 & n39222;
  assign n39252 = ~n39235 & n39251;
  assign n39253 = ~n39250 & ~n39252;
  assign n39254 = ~n39216 & ~n39222;
  assign n39255 = ~n39235 & n39254;
  assign n39256 = n39229 & n39255;
  assign n39257 = n39253 & ~n39256;
  assign n39258 = ~n39210 & ~n39257;
  assign n39259 = ~n39249 & ~n39258;
  assign n39260 = ~n39216 & n39222;
  assign n39261 = n39235 & n39260;
  assign n39262 = n39229 & n39261;
  assign n39263 = n39259 & ~n39262;
  assign n39264 = ~n39229 & n39254;
  assign n39265 = ~n39216 & ~n39235;
  assign n39266 = n39222 & n39265;
  assign n39267 = ~n39264 & ~n39266;
  assign n39268 = n39210 & ~n39267;
  assign n39269 = n39235 & n39251;
  assign n39270 = ~n39229 & n39269;
  assign n39271 = ~n39268 & ~n39270;
  assign n39272 = n39263 & n39271;
  assign n39273 = n39247 & ~n39272;
  assign n39274 = ~n39241 & ~n39273;
  assign n39275 = ~n39210 & ~n39247;
  assign n39276 = ~n39267 & n39275;
  assign n39277 = n39235 & n39254;
  assign n39278 = ~n39269 & ~n39277;
  assign n39279 = n39229 & ~n39278;
  assign n39280 = ~n39237 & ~n39279;
  assign n39281 = ~n39247 & ~n39280;
  assign n39282 = ~n39276 & ~n39281;
  assign n39283 = n39210 & ~n39247;
  assign n39284 = n39223 & ~n39229;
  assign n39285 = ~n39261 & ~n39284;
  assign n39286 = n39216 & ~n39235;
  assign n39287 = n39285 & ~n39286;
  assign n39288 = n39283 & ~n39287;
  assign n39289 = n39282 & ~n39288;
  assign n39290 = n39274 & n39289;
  assign n39291 = ~pi0864 & ~n39290;
  assign n39292 = pi0864 & n39282;
  assign n39293 = n39274 & n39292;
  assign n39294 = ~n39288 & n39293;
  assign po0904 = n39291 | n39294;
  assign n39296 = ~n38956 & ~n38965;
  assign n39297 = n38941 & ~n39296;
  assign n39298 = n38935 & n39001;
  assign n39299 = ~n39297 & ~n39298;
  assign n39300 = n38935 & n38950;
  assign n39301 = ~n38975 & ~n39300;
  assign n39302 = ~n38998 & n39301;
  assign n39303 = ~n38941 & ~n39302;
  assign n39304 = n39299 & ~n39303;
  assign n39305 = ~n38990 & ~n39304;
  assign n39306 = ~n38935 & n38976;
  assign n39307 = n38941 & n39306;
  assign n39308 = ~n38929 & n38973;
  assign n39309 = ~n39307 & ~n39308;
  assign n39310 = ~n38941 & n38981;
  assign n39311 = n39309 & ~n39310;
  assign n39312 = ~n38941 & n39005;
  assign n39313 = ~n38929 & ~n38935;
  assign n39314 = ~n38923 & n39313;
  assign n39315 = ~n38981 & ~n39314;
  assign n39316 = ~n38941 & n38950;
  assign n39317 = n39313 & n39316;
  assign n39318 = n38935 & n38965;
  assign n39319 = n38941 & n38975;
  assign n39320 = ~n39318 & ~n39319;
  assign n39321 = ~n38974 & n39320;
  assign n39322 = ~n39317 & n39321;
  assign n39323 = n39315 & n39322;
  assign n39324 = ~n39312 & n39323;
  assign n39325 = n38990 & ~n39324;
  assign n39326 = n39311 & ~n39325;
  assign n39327 = ~n39305 & n39326;
  assign n39328 = ~pi0870 & ~n39327;
  assign n39329 = pi0870 & n39311;
  assign n39330 = ~n39305 & n39329;
  assign n39331 = ~n39325 & n39330;
  assign po0905 = n39328 | n39331;
  assign n39333 = n38935 & n38962;
  assign n39334 = ~n39001 & ~n39333;
  assign n39335 = ~n38953 & n39334;
  assign n39336 = ~n38941 & ~n39335;
  assign n39337 = n38923 & ~n38935;
  assign n39338 = n38975 & n39337;
  assign n39339 = ~n38935 & n38965;
  assign n39340 = n38929 & ~n38950;
  assign n39341 = ~n38951 & ~n39340;
  assign n39342 = n38935 & ~n39341;
  assign n39343 = ~n39339 & ~n39342;
  assign n39344 = ~n39338 & n39343;
  assign n39345 = n38941 & ~n39344;
  assign n39346 = ~n39336 & ~n39345;
  assign n39347 = n38990 & ~n39346;
  assign n39348 = n38942 & ~n38950;
  assign n39349 = ~n38935 & n38950;
  assign n39350 = ~n38929 & n39349;
  assign n39351 = ~n39333 & ~n39350;
  assign n39352 = n38941 & ~n39351;
  assign n39353 = ~n38973 & ~n39352;
  assign n39354 = ~n38935 & n38967;
  assign n39355 = ~n38977 & ~n39354;
  assign n39356 = ~n38941 & n38975;
  assign n39357 = n38935 & n39356;
  assign n39358 = ~n39312 & ~n39357;
  assign n39359 = n39355 & n39358;
  assign n39360 = n39353 & n39359;
  assign n39361 = ~n39348 & n39360;
  assign n39362 = ~n38990 & ~n39361;
  assign n39363 = n38941 & n38956;
  assign n39364 = ~n38935 & n39363;
  assign n39365 = ~n39308 & ~n39364;
  assign n39366 = ~n39310 & n39365;
  assign n39367 = ~n38935 & n38998;
  assign n39368 = n38935 & n38957;
  assign n39369 = ~n39367 & ~n39368;
  assign n39370 = ~n38941 & ~n39369;
  assign n39371 = n39366 & ~n39370;
  assign n39372 = ~n39362 & n39371;
  assign n39373 = ~n39347 & n39372;
  assign n39374 = ~pi0878 & n39373;
  assign n39375 = pi0878 & ~n39373;
  assign po0906 = n39374 | n39375;
  assign n39377 = n39034 & ~n39048;
  assign n39378 = ~n39080 & ~n39377;
  assign n39379 = ~n39102 & n39378;
  assign n39380 = ~n39022 & ~n39379;
  assign n39381 = n39022 & n39040;
  assign n39382 = n39048 & n39381;
  assign n39383 = ~n39034 & ~n39048;
  assign n39384 = n39022 & ~n39040;
  assign n39385 = n39383 & n39384;
  assign n39386 = n39034 & n39040;
  assign n39387 = ~n39028 & n39386;
  assign n39388 = ~n39040 & n39071;
  assign n39389 = ~n39387 & ~n39388;
  assign n39390 = ~n39385 & n39389;
  assign n39391 = ~n39382 & n39390;
  assign n39392 = ~n39380 & n39391;
  assign n39393 = n39063 & ~n39392;
  assign n39394 = n39034 & n39053;
  assign n39395 = ~n39040 & n39394;
  assign n39396 = n39034 & n39088;
  assign n39397 = n39040 & n39396;
  assign n39398 = ~n39395 & ~n39397;
  assign n39399 = ~n39022 & ~n39398;
  assign n39400 = ~n39393 & ~n39399;
  assign n39401 = n39040 & n39071;
  assign n39402 = ~n39050 & ~n39084;
  assign n39403 = ~n39022 & ~n39402;
  assign n39404 = ~n39401 & ~n39403;
  assign n39405 = ~n39055 & n39404;
  assign n39406 = ~n39063 & ~n39405;
  assign n39407 = ~n39068 & ~n39088;
  assign n39408 = ~n39034 & ~n39407;
  assign n39409 = ~n39089 & ~n39408;
  assign n39410 = n39022 & ~n39409;
  assign n39411 = ~n39063 & n39410;
  assign n39412 = ~n39406 & ~n39411;
  assign n39413 = n39400 & n39412;
  assign n39414 = pi0871 & ~n39413;
  assign n39415 = ~pi0871 & n39400;
  assign n39416 = n39412 & n39415;
  assign po0907 = n39414 | n39416;
  assign n39418 = pi3757 & pi9040;
  assign n39419 = pi3777 & ~pi9040;
  assign n39420 = ~n39418 & ~n39419;
  assign n39421 = pi0855 & n39420;
  assign n39422 = ~pi0855 & ~n39420;
  assign n39423 = ~n39421 & ~n39422;
  assign n39424 = pi3729 & pi9040;
  assign n39425 = pi3816 & ~pi9040;
  assign n39426 = ~n39424 & ~n39425;
  assign n39427 = ~pi0839 & n39426;
  assign n39428 = pi0839 & ~n39426;
  assign n39429 = ~n39427 & ~n39428;
  assign n39430 = pi3745 & pi9040;
  assign n39431 = pi3751 & ~pi9040;
  assign n39432 = ~n39430 & ~n39431;
  assign n39433 = ~pi0847 & n39432;
  assign n39434 = pi0847 & ~n39432;
  assign n39435 = ~n39433 & ~n39434;
  assign n39436 = pi3737 & pi9040;
  assign n39437 = pi3731 & ~pi9040;
  assign n39438 = ~n39436 & ~n39437;
  assign n39439 = ~pi0848 & n39438;
  assign n39440 = pi0848 & ~n39438;
  assign n39441 = ~n39439 & ~n39440;
  assign n39442 = pi3816 & pi9040;
  assign n39443 = pi3756 & ~pi9040;
  assign n39444 = ~n39442 & ~n39443;
  assign n39445 = ~pi0849 & ~n39444;
  assign n39446 = pi0849 & n39444;
  assign n39447 = ~n39445 & ~n39446;
  assign n39448 = n39441 & ~n39447;
  assign n39449 = n39435 & n39448;
  assign n39450 = n39429 & n39449;
  assign n39451 = n39441 & n39447;
  assign n39452 = n39435 & n39451;
  assign n39453 = ~n39429 & n39452;
  assign n39454 = ~n39450 & ~n39453;
  assign n39455 = n39423 & ~n39454;
  assign n39456 = ~n39441 & ~n39447;
  assign n39457 = ~n39435 & n39456;
  assign n39458 = n39429 & n39457;
  assign n39459 = ~n39423 & n39458;
  assign n39460 = pi3740 & ~pi9040;
  assign n39461 = pi3751 & pi9040;
  assign n39462 = ~n39460 & ~n39461;
  assign n39463 = ~pi0858 & ~n39462;
  assign n39464 = pi0858 & n39462;
  assign n39465 = ~n39463 & ~n39464;
  assign n39466 = ~n39429 & n39435;
  assign n39467 = ~n39441 & n39466;
  assign n39468 = n39423 & n39467;
  assign n39469 = ~n39458 & ~n39468;
  assign n39470 = ~n39429 & ~n39447;
  assign n39471 = n39441 & n39470;
  assign n39472 = n39429 & n39456;
  assign n39473 = ~n39471 & ~n39472;
  assign n39474 = ~n39423 & ~n39473;
  assign n39475 = n39429 & n39435;
  assign n39476 = ~n39423 & n39447;
  assign n39477 = n39475 & n39476;
  assign n39478 = n39441 & n39477;
  assign n39479 = ~n39441 & n39447;
  assign n39480 = ~n39435 & n39479;
  assign n39481 = ~n39429 & n39480;
  assign n39482 = n39429 & ~n39435;
  assign n39483 = n39441 & n39482;
  assign n39484 = n39423 & n39483;
  assign n39485 = ~n39481 & ~n39484;
  assign n39486 = ~n39478 & n39485;
  assign n39487 = ~n39474 & n39486;
  assign n39488 = n39469 & n39487;
  assign n39489 = n39465 & ~n39488;
  assign n39490 = ~n39447 & n39468;
  assign n39491 = ~n39489 & ~n39490;
  assign n39492 = ~n39459 & n39491;
  assign n39493 = ~n39455 & n39492;
  assign n39494 = n39423 & n39447;
  assign n39495 = n39429 & ~n39441;
  assign n39496 = n39494 & n39495;
  assign n39497 = n39441 & n39475;
  assign n39498 = n39423 & n39497;
  assign n39499 = ~n39496 & ~n39498;
  assign n39500 = ~n39429 & ~n39435;
  assign n39501 = ~n39441 & n39500;
  assign n39502 = n39423 & n39501;
  assign n39503 = n39441 & n39500;
  assign n39504 = ~n39447 & n39503;
  assign n39505 = ~n39502 & ~n39504;
  assign n39506 = ~n39441 & n39475;
  assign n39507 = n39447 & n39506;
  assign n39508 = ~n39450 & ~n39507;
  assign n39509 = n39447 & n39466;
  assign n39510 = ~n39435 & n39441;
  assign n39511 = ~n39509 & ~n39510;
  assign n39512 = ~n39423 & ~n39511;
  assign n39513 = n39508 & ~n39512;
  assign n39514 = n39505 & n39513;
  assign n39515 = n39499 & n39514;
  assign n39516 = ~n39465 & ~n39515;
  assign n39517 = n39493 & ~n39516;
  assign n39518 = ~pi0868 & ~n39517;
  assign n39519 = pi0868 & n39493;
  assign n39520 = ~n39516 & n39519;
  assign po0908 = n39518 | n39520;
  assign n39522 = n39210 & n39229;
  assign n39523 = ~n39254 & ~n39269;
  assign n39524 = n39522 & ~n39523;
  assign n39525 = n39210 & n39235;
  assign n39526 = n39254 & n39525;
  assign n39527 = ~n39524 & ~n39526;
  assign n39528 = n39247 & ~n39527;
  assign n39529 = ~n39229 & ~n39235;
  assign n39530 = n39222 & n39529;
  assign n39531 = n39216 & n39530;
  assign n39532 = ~n39286 & ~n39529;
  assign n39533 = ~n39210 & ~n39532;
  assign n39534 = ~n39229 & n39235;
  assign n39535 = ~n39222 & n39534;
  assign n39536 = n39216 & n39535;
  assign n39537 = ~n39533 & ~n39536;
  assign n39538 = ~n39531 & n39537;
  assign n39539 = n39247 & ~n39538;
  assign n39540 = ~n39528 & ~n39539;
  assign n39541 = n39222 & n39236;
  assign n39542 = ~n39216 & n39541;
  assign n39543 = ~n39229 & n39261;
  assign n39544 = ~n39542 & ~n39543;
  assign n39545 = n39210 & ~n39544;
  assign n39546 = n39229 & n39277;
  assign n39547 = ~n39229 & n39286;
  assign n39548 = ~n39546 & ~n39547;
  assign n39549 = ~n39210 & ~n39548;
  assign n39550 = ~n39223 & ~n39286;
  assign n39551 = n39229 & ~n39550;
  assign n39552 = ~n39261 & ~n39551;
  assign n39553 = n39210 & ~n39552;
  assign n39554 = n39222 & ~n39229;
  assign n39555 = n39210 & n39554;
  assign n39556 = n39235 & n39555;
  assign n39557 = ~n39222 & ~n39235;
  assign n39558 = ~n39261 & ~n39557;
  assign n39559 = ~n39229 & ~n39558;
  assign n39560 = ~n39210 & n39229;
  assign n39561 = n39251 & n39560;
  assign n39562 = n39235 & n39561;
  assign n39563 = ~n39559 & ~n39562;
  assign n39564 = ~n39556 & n39563;
  assign n39565 = ~n39553 & n39564;
  assign n39566 = ~n39542 & n39565;
  assign n39567 = ~n39247 & ~n39566;
  assign n39568 = ~n39549 & ~n39567;
  assign n39569 = ~n39545 & n39568;
  assign n39570 = n39540 & n39569;
  assign n39571 = pi0873 & n39570;
  assign n39572 = ~pi0873 & ~n39570;
  assign po0909 = n39571 | n39572;
  assign n39574 = n38721 & ~n38735;
  assign n39575 = ~n38714 & n39574;
  assign n39576 = n38741 & n39575;
  assign n39577 = ~n38741 & n39179;
  assign n39578 = ~n38743 & ~n39577;
  assign n39579 = ~n39186 & n39578;
  assign n39580 = ~n39576 & n39579;
  assign n39581 = n38714 & n39174;
  assign n39582 = n39580 & ~n39581;
  assign n39583 = n38762 & ~n39582;
  assign n39584 = ~n38778 & ~n39189;
  assign n39585 = n38714 & ~n39584;
  assign n39586 = n38756 & ~n38762;
  assign n39587 = ~n38714 & n39586;
  assign n39588 = n38735 & ~n38741;
  assign n39589 = ~n38721 & n39588;
  assign n39590 = ~n39179 & ~n39589;
  assign n39591 = ~n38745 & n39590;
  assign n39592 = n38714 & ~n39591;
  assign n39593 = ~n38735 & n38794;
  assign n39594 = ~n38741 & n39593;
  assign n39595 = ~n39592 & ~n39594;
  assign n39596 = ~n38762 & ~n39595;
  assign n39597 = ~n39587 & ~n39596;
  assign n39598 = ~n39585 & n39597;
  assign n39599 = ~n38741 & n38777;
  assign n39600 = ~n39157 & ~n39599;
  assign n39601 = ~n38743 & ~n38752;
  assign n39602 = n39600 & n39601;
  assign n39603 = ~n38714 & ~n39602;
  assign n39604 = n39598 & ~n39603;
  assign n39605 = ~n39583 & n39604;
  assign n39606 = ~pi0894 & ~n39605;
  assign n39607 = pi0894 & n39598;
  assign n39608 = ~n39583 & n39607;
  assign n39609 = ~n39603 & n39608;
  assign po0910 = n39606 | n39609;
  assign n39611 = ~n38941 & n38957;
  assign n39612 = ~n38935 & n39611;
  assign n39613 = ~n39367 & ~n39612;
  assign n39614 = ~n38935 & ~n38950;
  assign n39615 = ~n39314 & ~n39614;
  assign n39616 = n38941 & ~n39615;
  assign n39617 = ~n38929 & n38935;
  assign n39618 = n38923 & n39617;
  assign n39619 = ~n39616 & ~n39618;
  assign n39620 = n39613 & n39619;
  assign n39621 = n38990 & ~n39620;
  assign n39622 = ~n38967 & ~n38977;
  assign n39623 = ~n38935 & n38964;
  assign n39624 = n39622 & ~n39623;
  assign n39625 = ~n38941 & ~n39624;
  assign n39626 = n38957 & n38972;
  assign n39627 = ~n38953 & ~n39626;
  assign n39628 = ~n39625 & n39627;
  assign n39629 = ~n38998 & ~n39006;
  assign n39630 = n38941 & ~n39629;
  assign n39631 = n39628 & ~n39630;
  assign n39632 = ~n38990 & ~n39631;
  assign n39633 = ~n39621 & ~n39632;
  assign n39634 = n38935 & n39002;
  assign n39635 = ~n38935 & ~n38955;
  assign n39636 = ~n39634 & ~n39635;
  assign n39637 = n38941 & n39636;
  assign n39638 = n38935 & ~n38941;
  assign n39639 = ~n38967 & n39296;
  assign n39640 = n39638 & ~n39639;
  assign n39641 = ~n39637 & ~n39640;
  assign n39642 = n39633 & n39641;
  assign n39643 = ~pi0865 & ~n39642;
  assign n39644 = pi0865 & n39641;
  assign n39645 = ~n39632 & n39644;
  assign n39646 = ~n39621 & n39645;
  assign po0911 = n39643 | n39646;
  assign n39648 = pi3735 & pi9040;
  assign n39649 = pi3733 & ~pi9040;
  assign n39650 = ~n39648 & ~n39649;
  assign n39651 = ~pi0840 & ~n39650;
  assign n39652 = pi0840 & n39650;
  assign n39653 = ~n39651 & ~n39652;
  assign n39654 = pi3746 & pi9040;
  assign n39655 = pi3768 & ~pi9040;
  assign n39656 = ~n39654 & ~n39655;
  assign n39657 = pi0862 & n39656;
  assign n39658 = ~pi0862 & ~n39656;
  assign n39659 = ~n39657 & ~n39658;
  assign n39660 = pi3742 & pi9040;
  assign n39661 = pi3765 & ~pi9040;
  assign n39662 = ~n39660 & ~n39661;
  assign n39663 = ~pi0847 & n39662;
  assign n39664 = pi0847 & ~n39662;
  assign n39665 = ~n39663 & ~n39664;
  assign n39666 = pi3714 & pi9040;
  assign n39667 = pi3742 & ~pi9040;
  assign n39668 = ~n39666 & ~n39667;
  assign n39669 = ~pi0858 & ~n39668;
  assign n39670 = pi0858 & ~n39666;
  assign n39671 = ~n39667 & n39670;
  assign n39672 = ~n39669 & ~n39671;
  assign n39673 = pi3743 & pi9040;
  assign n39674 = pi3753 & ~pi9040;
  assign n39675 = ~n39673 & ~n39674;
  assign n39676 = ~pi0851 & ~n39675;
  assign n39677 = pi0851 & n39675;
  assign n39678 = ~n39676 & ~n39677;
  assign n39679 = ~n39672 & ~n39678;
  assign n39680 = ~n39665 & n39679;
  assign n39681 = n39659 & n39680;
  assign n39682 = ~n39672 & n39678;
  assign n39683 = n39665 & n39682;
  assign n39684 = n39659 & n39683;
  assign n39685 = ~n39681 & ~n39684;
  assign n39686 = n39672 & n39678;
  assign n39687 = n39665 & n39686;
  assign n39688 = n39665 & n39679;
  assign n39689 = ~n39659 & n39688;
  assign n39690 = ~n39687 & ~n39689;
  assign n39691 = pi3748 & pi9040;
  assign n39692 = pi3715 & ~pi9040;
  assign n39693 = ~n39691 & ~n39692;
  assign n39694 = ~pi0836 & n39693;
  assign n39695 = pi0836 & ~n39693;
  assign n39696 = ~n39694 & ~n39695;
  assign n39697 = ~n39690 & ~n39696;
  assign n39698 = n39685 & ~n39697;
  assign n39699 = ~n39659 & n39696;
  assign n39700 = n39672 & n39699;
  assign n39701 = n39698 & ~n39700;
  assign n39702 = n39653 & ~n39701;
  assign n39703 = n39659 & n39672;
  assign n39704 = n39665 & n39703;
  assign n39705 = ~n39678 & n39704;
  assign n39706 = n39696 & n39705;
  assign n39707 = ~n39659 & ~n39696;
  assign n39708 = n39672 & ~n39678;
  assign n39709 = n39665 & n39708;
  assign n39710 = n39707 & n39709;
  assign n39711 = ~n39659 & ~n39665;
  assign n39712 = ~n39672 & n39711;
  assign n39713 = ~n39710 & ~n39712;
  assign n39714 = ~n39665 & n39682;
  assign n39715 = ~n39687 & ~n39714;
  assign n39716 = ~n39659 & n39682;
  assign n39717 = n39715 & ~n39716;
  assign n39718 = n39696 & ~n39717;
  assign n39719 = ~n39665 & ~n39678;
  assign n39720 = n39672 & n39719;
  assign n39721 = n39659 & n39720;
  assign n39722 = n39659 & n39688;
  assign n39723 = ~n39721 & ~n39722;
  assign n39724 = ~n39665 & n39686;
  assign n39725 = ~n39696 & n39724;
  assign n39726 = n39723 & ~n39725;
  assign n39727 = ~n39718 & n39726;
  assign n39728 = n39713 & n39727;
  assign n39729 = ~n39653 & ~n39728;
  assign n39730 = ~n39706 & ~n39729;
  assign n39731 = ~n39702 & n39730;
  assign n39732 = n39707 & n39714;
  assign n39733 = ~n39696 & n39719;
  assign n39734 = n39659 & n39733;
  assign n39735 = ~n39732 & ~n39734;
  assign n39736 = n39684 & ~n39696;
  assign n39737 = n39735 & ~n39736;
  assign n39738 = n39731 & n39737;
  assign n39739 = ~pi0875 & ~n39738;
  assign n39740 = ~n39702 & n39737;
  assign n39741 = n39730 & n39740;
  assign n39742 = pi0875 & n39741;
  assign po0912 = n39739 | n39742;
  assign n39744 = n39210 & n39266;
  assign n39745 = ~n39229 & n39251;
  assign n39746 = ~n39250 & ~n39745;
  assign n39747 = n39210 & ~n39746;
  assign n39748 = ~n39210 & ~n39558;
  assign n39749 = ~n39747 & ~n39748;
  assign n39750 = ~n39546 & n39749;
  assign n39751 = n39247 & ~n39750;
  assign n39752 = ~n39744 & ~n39751;
  assign n39753 = ~n39235 & n39522;
  assign n39754 = ~n39534 & ~n39753;
  assign n39755 = ~n39216 & ~n39754;
  assign n39756 = ~n39237 & ~n39755;
  assign n39757 = ~n39535 & n39756;
  assign n39758 = ~n39210 & n39252;
  assign n39759 = n39229 & n39269;
  assign n39760 = ~n39758 & ~n39759;
  assign n39761 = n39757 & n39760;
  assign n39762 = ~n39247 & ~n39761;
  assign n39763 = ~n39229 & n39255;
  assign n39764 = n39229 & n39251;
  assign n39765 = ~n39763 & ~n39764;
  assign n39766 = ~n39210 & ~n39765;
  assign n39767 = ~n39762 & ~n39766;
  assign n39768 = n39752 & n39767;
  assign n39769 = ~pi0902 & ~n39768;
  assign n39770 = ~n39751 & n39767;
  assign n39771 = pi0902 & n39770;
  assign n39772 = ~n39744 & n39771;
  assign po0913 = n39769 | n39772;
  assign n39774 = ~n39678 & n39711;
  assign n39775 = ~n39672 & n39774;
  assign n39776 = ~n39659 & n39724;
  assign n39777 = ~n39683 & ~n39776;
  assign n39778 = n39659 & n39719;
  assign n39779 = ~n39659 & n39709;
  assign n39780 = ~n39778 & ~n39779;
  assign n39781 = n39777 & n39780;
  assign n39782 = n39696 & ~n39781;
  assign n39783 = n39659 & n39686;
  assign n39784 = ~n39712 & ~n39783;
  assign n39785 = ~n39688 & n39784;
  assign n39786 = ~n39696 & ~n39785;
  assign n39787 = n39659 & n39665;
  assign n39788 = n39678 & n39787;
  assign n39789 = n39672 & n39788;
  assign n39790 = ~n39786 & ~n39789;
  assign n39791 = ~n39782 & n39790;
  assign n39792 = ~n39775 & n39791;
  assign n39793 = ~n39653 & ~n39792;
  assign n39794 = n39659 & n39696;
  assign n39795 = n39724 & n39794;
  assign n39796 = n39688 & n39696;
  assign n39797 = n39696 & n39714;
  assign n39798 = ~n39796 & ~n39797;
  assign n39799 = ~n39659 & ~n39798;
  assign n39800 = ~n39795 & ~n39799;
  assign n39801 = n39659 & n39682;
  assign n39802 = ~n39659 & n39686;
  assign n39803 = ~n39801 & ~n39802;
  assign n39804 = ~n39720 & n39803;
  assign n39805 = ~n39683 & n39804;
  assign n39806 = ~n39696 & ~n39805;
  assign n39807 = ~n39659 & n39687;
  assign n39808 = ~n39806 & ~n39807;
  assign n39809 = ~n39659 & n39720;
  assign n39810 = ~n39705 & ~n39809;
  assign n39811 = n39808 & n39810;
  assign n39812 = n39800 & n39811;
  assign n39813 = n39653 & ~n39812;
  assign n39814 = ~n39685 & n39696;
  assign n39815 = ~n39813 & ~n39814;
  assign n39816 = ~n39722 & ~n39809;
  assign n39817 = ~n39696 & ~n39816;
  assign n39818 = n39815 & ~n39817;
  assign n39819 = ~n39793 & n39818;
  assign n39820 = pi0880 & ~n39819;
  assign n39821 = ~pi0880 & n39819;
  assign po0914 = n39820 | n39821;
  assign n39823 = ~n39040 & n39054;
  assign n39824 = ~n39388 & ~n39823;
  assign n39825 = n39022 & ~n39824;
  assign n39826 = n39050 & n39381;
  assign n39827 = ~n39825 & ~n39826;
  assign n39828 = ~n39100 & n39827;
  assign n39829 = n39040 & n39084;
  assign n39830 = ~n39396 & ~n39829;
  assign n39831 = ~n39054 & n39830;
  assign n39832 = n39022 & ~n39831;
  assign n39833 = n39063 & n39832;
  assign n39834 = ~n39022 & n39394;
  assign n39835 = ~n39080 & ~n39098;
  assign n39836 = ~n39073 & n39835;
  assign n39837 = ~n39834 & n39836;
  assign n39838 = n39063 & ~n39837;
  assign n39839 = ~n39022 & n39034;
  assign n39840 = n39028 & n39839;
  assign n39841 = ~n39048 & n39840;
  assign n39842 = ~n39040 & n39841;
  assign n39843 = n39040 & n39108;
  assign n39844 = ~n39841 & ~n39843;
  assign n39845 = ~n39387 & n39844;
  assign n39846 = n39028 & n39078;
  assign n39847 = n39040 & n39068;
  assign n39848 = ~n39049 & ~n39847;
  assign n39849 = n39022 & ~n39848;
  assign n39850 = ~n39846 & ~n39849;
  assign n39851 = n39845 & n39850;
  assign n39852 = ~n39063 & ~n39851;
  assign n39853 = ~n39842 & ~n39852;
  assign n39854 = ~n39838 & n39853;
  assign n39855 = ~n39833 & n39854;
  assign n39856 = n39828 & n39855;
  assign n39857 = pi0882 & ~n39856;
  assign n39858 = ~pi0882 & n39828;
  assign n39859 = n39855 & n39858;
  assign po0915 = n39857 | n39859;
  assign n39861 = n39678 & n39711;
  assign n39862 = ~n39687 & ~n39712;
  assign n39863 = n39696 & ~n39862;
  assign n39864 = ~n39861 & ~n39863;
  assign n39865 = n39665 & ~n39672;
  assign n39866 = n39665 & ~n39678;
  assign n39867 = ~n39659 & n39866;
  assign n39868 = n39659 & n39679;
  assign n39869 = ~n39867 & ~n39868;
  assign n39870 = ~n39865 & n39869;
  assign n39871 = ~n39724 & n39870;
  assign n39872 = ~n39696 & ~n39871;
  assign n39873 = n39864 & ~n39872;
  assign n39874 = ~n39721 & n39873;
  assign n39875 = n39653 & ~n39874;
  assign n39876 = ~n39659 & n39683;
  assign n39877 = n39723 & ~n39876;
  assign n39878 = ~n39696 & ~n39877;
  assign n39879 = ~n39875 & ~n39878;
  assign n39880 = n39665 & n39672;
  assign n39881 = n39696 & n39880;
  assign n39882 = n39659 & n39881;
  assign n39883 = n39707 & n39719;
  assign n39884 = n39659 & n39714;
  assign n39885 = ~n39883 & ~n39884;
  assign n39886 = ~n39665 & ~n39672;
  assign n39887 = n39659 & n39886;
  assign n39888 = ~n39709 & ~n39887;
  assign n39889 = n39696 & ~n39888;
  assign n39890 = n39696 & n39865;
  assign n39891 = ~n39659 & n39890;
  assign n39892 = ~n39889 & ~n39891;
  assign n39893 = n39885 & n39892;
  assign n39894 = ~n39653 & ~n39893;
  assign n39895 = ~n39882 & ~n39894;
  assign n39896 = ~n39776 & n39895;
  assign n39897 = n39879 & n39896;
  assign n39898 = ~pi0874 & ~n39897;
  assign n39899 = ~n39776 & ~n39875;
  assign n39900 = ~n39878 & n39899;
  assign n39901 = n39895 & n39900;
  assign n39902 = pi0874 & n39901;
  assign po0916 = n39898 | n39902;
  assign n39904 = n39447 & n39467;
  assign n39905 = ~n39447 & n39506;
  assign n39906 = ~n39904 & ~n39905;
  assign n39907 = ~n39441 & n39482;
  assign n39908 = n39447 & n39907;
  assign n39909 = n39447 & n39500;
  assign n39910 = ~n39447 & n39483;
  assign n39911 = ~n39909 & ~n39910;
  assign n39912 = ~n39423 & ~n39911;
  assign n39913 = ~n39908 & ~n39912;
  assign n39914 = n39423 & n39482;
  assign n39915 = n39447 & n39914;
  assign n39916 = ~n39498 & ~n39915;
  assign n39917 = n39913 & n39916;
  assign n39918 = n39906 & n39917;
  assign n39919 = n39465 & ~n39918;
  assign n39920 = ~n39423 & ~n39465;
  assign n39921 = n39429 & n39451;
  assign n39922 = n39435 & n39441;
  assign n39923 = ~n39921 & ~n39922;
  assign n39924 = n39920 & ~n39923;
  assign n39925 = ~n39458 & ~n39471;
  assign n39926 = ~n39441 & n39494;
  assign n39927 = ~n39482 & n39926;
  assign n39928 = ~n39468 & ~n39927;
  assign n39929 = n39925 & n39928;
  assign n39930 = ~n39465 & ~n39929;
  assign n39931 = n39441 & n39466;
  assign n39932 = ~n39423 & ~n39447;
  assign n39933 = n39931 & n39932;
  assign n39934 = ~n39447 & n39501;
  assign n39935 = ~n39905 & ~n39934;
  assign n39936 = ~n39423 & ~n39935;
  assign n39937 = ~n39933 & ~n39936;
  assign n39938 = n39423 & n39458;
  assign n39939 = n39937 & ~n39938;
  assign n39940 = ~n39930 & n39939;
  assign n39941 = ~n39924 & n39940;
  assign n39942 = ~n39919 & n39941;
  assign n39943 = n39423 & ~n39447;
  assign n39944 = n39503 & n39943;
  assign n39945 = n39942 & ~n39944;
  assign n39946 = ~pi0872 & ~n39945;
  assign n39947 = n39941 & ~n39944;
  assign n39948 = pi0872 & n39947;
  assign n39949 = ~n39919 & n39948;
  assign po0917 = n39946 | n39949;
  assign n39951 = ~n38743 & ~n38750;
  assign n39952 = ~n38714 & ~n39951;
  assign n39953 = ~n38805 & ~n39952;
  assign n39954 = ~n38721 & ~n38735;
  assign n39955 = n38714 & n39954;
  assign n39956 = n38741 & n39955;
  assign n39957 = ~n38714 & n38748;
  assign n39958 = n38741 & n39957;
  assign n39959 = ~n39166 & ~n39958;
  assign n39960 = n38721 & n39588;
  assign n39961 = n38741 & n38794;
  assign n39962 = ~n39960 & ~n39961;
  assign n39963 = ~n39954 & n39962;
  assign n39964 = n38714 & ~n39963;
  assign n39965 = ~n38746 & ~n39964;
  assign n39966 = n39959 & n39965;
  assign n39967 = ~n38762 & ~n39966;
  assign n39968 = ~n39956 & ~n39967;
  assign n39969 = ~n38767 & ~n38795;
  assign n39970 = ~n38777 & n39969;
  assign n39971 = ~n38714 & ~n39970;
  assign n39972 = ~n38741 & n38772;
  assign n39973 = ~n38798 & ~n39972;
  assign n39974 = n38714 & ~n39973;
  assign n39975 = ~n39177 & ~n39974;
  assign n39976 = ~n39971 & n39975;
  assign n39977 = ~n38778 & ~n38784;
  assign n39978 = n39976 & n39977;
  assign n39979 = n38762 & ~n39978;
  assign n39980 = n39968 & ~n39979;
  assign n39981 = n39953 & n39980;
  assign n39982 = ~pi0900 & ~n39981;
  assign n39983 = pi0900 & n39968;
  assign n39984 = n39953 & n39983;
  assign n39985 = ~n39979 & n39984;
  assign po0918 = n39982 | n39985;
  assign n39987 = pi3720 & pi9040;
  assign n39988 = pi3745 & ~pi9040;
  assign n39989 = ~n39987 & ~n39988;
  assign n39990 = pi0861 & n39989;
  assign n39991 = ~pi0861 & ~n39989;
  assign n39992 = ~n39990 & ~n39991;
  assign n39993 = pi3724 & pi9040;
  assign n39994 = pi3732 & ~pi9040;
  assign n39995 = ~n39993 & ~n39994;
  assign n39996 = ~pi0845 & n39995;
  assign n39997 = pi0845 & ~n39995;
  assign n39998 = ~n39996 & ~n39997;
  assign n39999 = pi3719 & pi9040;
  assign n40000 = pi3720 & ~pi9040;
  assign n40001 = ~n39999 & ~n40000;
  assign n40002 = ~pi0848 & n40001;
  assign n40003 = pi0848 & ~n40001;
  assign n40004 = ~n40002 & ~n40003;
  assign n40005 = ~n39998 & ~n40004;
  assign n40006 = n39992 & n40005;
  assign n40007 = ~pi0848 & ~n40001;
  assign n40008 = pi0848 & n40001;
  assign n40009 = ~n40007 & ~n40008;
  assign n40010 = ~n39998 & ~n40009;
  assign n40011 = ~n39992 & n40010;
  assign n40012 = ~n40006 & ~n40011;
  assign n40013 = pi3718 & pi9040;
  assign n40014 = pi3724 & ~pi9040;
  assign n40015 = ~n40013 & ~n40014;
  assign n40016 = pi0843 & n40015;
  assign n40017 = ~pi0843 & ~n40015;
  assign n40018 = ~n40016 & ~n40017;
  assign n40019 = n39992 & ~n40018;
  assign n40020 = n40009 & n40019;
  assign n40021 = n40012 & ~n40020;
  assign n40022 = pi3730 & pi9040;
  assign n40023 = pi3739 & ~pi9040;
  assign n40024 = ~n40022 & ~n40023;
  assign n40025 = pi0826 & n40024;
  assign n40026 = ~pi0826 & ~n40024;
  assign n40027 = ~n40025 & ~n40026;
  assign n40028 = pi3734 & pi9040;
  assign n40029 = pi3744 & ~pi9040;
  assign n40030 = ~n40028 & ~n40029;
  assign n40031 = ~pi0839 & n40030;
  assign n40032 = pi0839 & ~n40030;
  assign n40033 = ~n40031 & ~n40032;
  assign n40034 = ~n40027 & ~n40033;
  assign n40035 = ~n40021 & n40034;
  assign n40036 = n39998 & ~n40009;
  assign n40037 = n39992 & n40036;
  assign n40038 = ~n40033 & n40037;
  assign n40039 = n40018 & n40038;
  assign n40040 = n39992 & n40010;
  assign n40041 = n40027 & n40040;
  assign n40042 = ~n39992 & n40009;
  assign n40043 = n39998 & ~n40004;
  assign n40044 = n40018 & n40043;
  assign n40045 = ~n40042 & ~n40044;
  assign n40046 = n40027 & ~n40045;
  assign n40047 = ~n40041 & ~n40046;
  assign n40048 = ~n40033 & ~n40047;
  assign n40049 = ~n40039 & ~n40048;
  assign n40050 = ~n39992 & n40018;
  assign n40051 = n40009 & n40050;
  assign n40052 = ~n39992 & ~n40018;
  assign n40053 = ~n40009 & n40052;
  assign n40054 = n39998 & n40053;
  assign n40055 = ~n40051 & ~n40054;
  assign n40056 = n40027 & ~n40055;
  assign n40057 = n40049 & ~n40056;
  assign n40058 = n40018 & ~n40027;
  assign n40059 = n40043 & n40058;
  assign n40060 = n39992 & n40059;
  assign n40061 = ~n40005 & ~n40036;
  assign n40062 = n40019 & ~n40061;
  assign n40063 = ~n39998 & n40053;
  assign n40064 = ~n40062 & ~n40063;
  assign n40065 = ~n39992 & n40043;
  assign n40066 = ~n40018 & ~n40027;
  assign n40067 = n40065 & n40066;
  assign n40068 = n40050 & ~n40061;
  assign n40069 = n40018 & n40040;
  assign n40070 = ~n40068 & ~n40069;
  assign n40071 = ~n40067 & n40070;
  assign n40072 = n40064 & n40071;
  assign n40073 = ~n40060 & n40072;
  assign n40074 = ~n40018 & n40027;
  assign n40075 = n39992 & n40074;
  assign n40076 = n39998 & n40075;
  assign n40077 = n40073 & ~n40076;
  assign n40078 = n40033 & ~n40077;
  assign n40079 = n40057 & ~n40078;
  assign n40080 = ~n40035 & n40079;
  assign n40081 = ~pi0886 & ~n40080;
  assign n40082 = pi0886 & n40057;
  assign n40083 = ~n40035 & n40082;
  assign n40084 = ~n40078 & n40083;
  assign po0919 = n40081 | n40084;
  assign n40086 = ~n38853 & ~n38856;
  assign n40087 = n38831 & ~n40086;
  assign n40088 = n38818 & n40087;
  assign n40089 = ~n39135 & ~n40088;
  assign n40090 = ~n38818 & n38876;
  assign n40091 = ~n39137 & ~n40090;
  assign n40092 = ~n38824 & n40091;
  assign n40093 = n38818 & n38847;
  assign n40094 = ~n38846 & n38865;
  assign n40095 = n38818 & n38856;
  assign n40096 = ~n40094 & ~n40095;
  assign n40097 = n38824 & n40096;
  assign n40098 = ~n40087 & n40097;
  assign n40099 = ~n40093 & n40098;
  assign n40100 = ~n40092 & ~n40099;
  assign n40101 = n40089 & ~n40100;
  assign n40102 = n38888 & ~n40101;
  assign n40103 = ~n38824 & ~n40086;
  assign n40104 = ~n38818 & n40103;
  assign n40105 = n38818 & n38858;
  assign n40106 = ~n38900 & ~n40105;
  assign n40107 = ~n38824 & ~n40106;
  assign n40108 = ~n38831 & n40103;
  assign n40109 = ~n40107 & ~n40108;
  assign n40110 = ~n40104 & n40109;
  assign n40111 = ~n38888 & ~n40110;
  assign n40112 = ~n40102 & ~n40111;
  assign n40113 = n38824 & ~n40091;
  assign n40114 = ~n38894 & ~n40113;
  assign n40115 = ~n38888 & ~n40114;
  assign n40116 = ~n38824 & n38894;
  assign n40117 = n38824 & ~n40089;
  assign n40118 = ~n40116 & ~n40117;
  assign n40119 = ~n40115 & n40118;
  assign n40120 = n40112 & n40119;
  assign n40121 = pi0908 & ~n40120;
  assign n40122 = ~pi0908 & n40119;
  assign n40123 = ~n40111 & n40122;
  assign n40124 = ~n40102 & n40123;
  assign po0920 = n40121 | n40124;
  assign n40126 = n39040 & ~n39407;
  assign n40127 = ~n39034 & n40126;
  assign n40128 = n39028 & n39386;
  assign n40129 = ~n39110 & ~n40128;
  assign n40130 = ~n39396 & n40129;
  assign n40131 = ~n39022 & ~n40130;
  assign n40132 = ~n39083 & ~n39394;
  assign n40133 = n39022 & ~n40132;
  assign n40134 = ~n40131 & ~n40133;
  assign n40135 = ~n40127 & n40134;
  assign n40136 = ~n39040 & n39050;
  assign n40137 = n40135 & ~n40136;
  assign n40138 = ~n39063 & ~n40137;
  assign n40139 = ~n39054 & ~n39084;
  assign n40140 = ~n39050 & ~n39396;
  assign n40141 = n40139 & n40140;
  assign n40142 = n39040 & ~n40141;
  assign n40143 = n39067 & ~n40132;
  assign n40144 = ~n40142 & ~n40143;
  assign n40145 = ~n39388 & n40144;
  assign n40146 = n39063 & ~n40145;
  assign n40147 = ~n40138 & ~n40146;
  assign n40148 = n39040 & n39394;
  assign n40149 = ~n40136 & ~n40148;
  assign n40150 = n39022 & ~n40149;
  assign n40151 = n40147 & ~n40150;
  assign n40152 = pi0877 & ~n40151;
  assign n40153 = ~pi0877 & ~n40150;
  assign n40154 = ~n40146 & n40153;
  assign n40155 = ~n40138 & n40154;
  assign po0921 = n40152 | n40155;
  assign n40157 = n39992 & n40043;
  assign n40158 = n40027 & n40157;
  assign n40159 = ~n40018 & n40158;
  assign n40160 = n40010 & n40074;
  assign n40161 = ~n39992 & n40160;
  assign n40162 = ~n40159 & ~n40161;
  assign n40163 = ~n40063 & ~n40067;
  assign n40164 = ~n39998 & n40018;
  assign n40165 = n39992 & n40164;
  assign n40166 = ~n40044 & ~n40165;
  assign n40167 = n40027 & ~n40166;
  assign n40168 = ~n40027 & ~n40052;
  assign n40169 = ~n40061 & n40168;
  assign n40170 = ~n39992 & ~n40043;
  assign n40171 = n40027 & n40170;
  assign n40172 = ~n40018 & n40171;
  assign n40173 = ~n40169 & ~n40172;
  assign n40174 = ~n40167 & n40173;
  assign n40175 = n40163 & n40174;
  assign n40176 = ~n40033 & ~n40175;
  assign n40177 = n40162 & ~n40176;
  assign n40178 = n40006 & ~n40027;
  assign n40179 = n40018 & n40178;
  assign n40180 = ~n40027 & n40033;
  assign n40181 = n40052 & ~n40061;
  assign n40182 = ~n40044 & ~n40181;
  assign n40183 = ~n40040 & n40182;
  assign n40184 = n40180 & ~n40183;
  assign n40185 = n40011 & n40018;
  assign n40186 = ~n39992 & n40164;
  assign n40187 = n40018 & n40036;
  assign n40188 = ~n40186 & ~n40187;
  assign n40189 = ~n40018 & n40043;
  assign n40190 = ~n40037 & ~n40189;
  assign n40191 = n40188 & n40190;
  assign n40192 = n40027 & ~n40191;
  assign n40193 = ~n40185 & ~n40192;
  assign n40194 = n40033 & ~n40193;
  assign n40195 = ~n40184 & ~n40194;
  assign n40196 = ~n40179 & n40195;
  assign n40197 = n40177 & n40196;
  assign n40198 = pi0887 & ~n40197;
  assign n40199 = ~pi0887 & n40177;
  assign n40200 = n40196 & n40199;
  assign po0922 = n40198 | n40200;
  assign n40202 = ~n39222 & n39238;
  assign n40203 = ~n39269 & ~n40202;
  assign n40204 = n39210 & ~n40203;
  assign n40205 = n39229 & n39260;
  assign n40206 = ~n39535 & ~n40205;
  assign n40207 = ~n39210 & ~n40206;
  assign n40208 = ~n39556 & ~n39763;
  assign n40209 = ~n39237 & n40208;
  assign n40210 = ~n40207 & n40209;
  assign n40211 = ~n40204 & n40210;
  assign n40212 = ~n39531 & ~n39542;
  assign n40213 = n40211 & n40212;
  assign n40214 = n39247 & ~n40213;
  assign n40215 = n39223 & n39529;
  assign n40216 = n39278 & ~n40215;
  assign n40217 = ~n39210 & ~n40216;
  assign n40218 = ~n39229 & n39266;
  assign n40219 = ~n40217 & ~n40218;
  assign n40220 = n39216 & n39238;
  assign n40221 = ~n39764 & ~n40220;
  assign n40222 = ~n39210 & ~n40221;
  assign n40223 = ~n39210 & n39260;
  assign n40224 = ~n39229 & n40223;
  assign n40225 = ~n40222 & ~n40224;
  assign n40226 = n40219 & n40225;
  assign n40227 = ~n39247 & ~n40226;
  assign n40228 = ~n39255 & ~n39262;
  assign n40229 = ~n39536 & n40228;
  assign n40230 = n39283 & ~n40229;
  assign n40231 = ~n40227 & ~n40230;
  assign n40232 = ~n39237 & ~n39531;
  assign n40233 = n39210 & ~n40232;
  assign n40234 = n40231 & ~n40233;
  assign n40235 = ~n40214 & n40234;
  assign n40236 = ~pi0885 & n40235;
  assign n40237 = pi0885 & ~n40235;
  assign po0923 = n40236 | n40237;
  assign n40239 = ~n39447 & n39914;
  assign n40240 = ~n39429 & n39451;
  assign n40241 = ~n39931 & ~n40240;
  assign n40242 = n39423 & ~n40241;
  assign n40243 = ~n40239 & ~n40242;
  assign n40244 = n39500 & n39932;
  assign n40245 = ~n39423 & n39497;
  assign n40246 = ~n40244 & ~n40245;
  assign n40247 = n40243 & n40246;
  assign n40248 = ~n39429 & n39456;
  assign n40249 = ~n39450 & ~n40248;
  assign n40250 = ~n39507 & n40249;
  assign n40251 = n40247 & n40250;
  assign n40252 = ~n39465 & ~n40251;
  assign n40253 = ~n39458 & ~n39931;
  assign n40254 = ~n39509 & n40253;
  assign n40255 = ~n39423 & ~n40254;
  assign n40256 = n39447 & n39483;
  assign n40257 = ~n39481 & ~n40256;
  assign n40258 = ~n39944 & n40257;
  assign n40259 = n39423 & n39506;
  assign n40260 = n40258 & ~n40259;
  assign n40261 = ~n40255 & n40260;
  assign n40262 = n39465 & ~n40261;
  assign n40263 = ~n39490 & ~n39496;
  assign n40264 = ~n39450 & n40257;
  assign n40265 = ~n39423 & ~n40264;
  assign n40266 = n40263 & ~n40265;
  assign n40267 = ~n40262 & n40266;
  assign n40268 = ~n40252 & n40267;
  assign n40269 = pi0881 & ~n40268;
  assign n40270 = ~pi0881 & n40268;
  assign po0924 = n40269 | n40270;
  assign n40272 = ~n39904 & ~n39921;
  assign n40273 = n39465 & ~n40272;
  assign n40274 = ~n39423 & n39907;
  assign n40275 = ~n39457 & ~n39472;
  assign n40276 = ~n39423 & ~n40275;
  assign n40277 = ~n40274 & ~n40276;
  assign n40278 = n39465 & ~n40277;
  assign n40279 = ~n40273 & ~n40278;
  assign n40280 = n39467 & n39476;
  assign n40281 = ~n39478 & ~n40280;
  assign n40282 = ~n39471 & ~n39510;
  assign n40283 = n39423 & ~n40282;
  assign n40284 = n39465 & n40283;
  assign n40285 = n40281 & ~n40284;
  assign n40286 = ~n39447 & n39467;
  assign n40287 = ~n39447 & n39475;
  assign n40288 = ~n39453 & ~n40287;
  assign n40289 = n39423 & ~n40288;
  assign n40290 = ~n39458 & ~n39481;
  assign n40291 = ~n39447 & n39466;
  assign n40292 = ~n39503 & ~n40291;
  assign n40293 = ~n39423 & ~n40292;
  assign n40294 = n40290 & ~n40293;
  assign n40295 = ~n40289 & n40294;
  assign n40296 = ~n40286 & n40295;
  assign n40297 = ~n39465 & ~n40296;
  assign n40298 = ~n39507 & n40257;
  assign n40299 = n39423 & ~n40298;
  assign n40300 = ~n40297 & ~n40299;
  assign n40301 = n40285 & n40300;
  assign n40302 = n40279 & n40301;
  assign n40303 = ~pi0888 & ~n40302;
  assign n40304 = pi0888 & n40285;
  assign n40305 = n40279 & n40304;
  assign n40306 = n40300 & n40305;
  assign po0925 = n40303 | n40306;
  assign n40308 = ~n38824 & n38855;
  assign n40309 = n38865 & ~n40086;
  assign n40310 = ~n38859 & ~n39135;
  assign n40311 = ~n40309 & n40310;
  assign n40312 = n38824 & ~n40311;
  assign n40313 = n38818 & n38892;
  assign n40314 = ~n40312 & ~n40313;
  assign n40315 = ~n38831 & n38858;
  assign n40316 = ~n38818 & n39142;
  assign n40317 = ~n40315 & ~n40316;
  assign n40318 = ~n40095 & n40317;
  assign n40319 = ~n38824 & ~n40318;
  assign n40320 = n40314 & ~n40319;
  assign n40321 = n38888 & ~n40320;
  assign n40322 = ~n40308 & ~n40321;
  assign n40323 = ~n38818 & n38856;
  assign n40324 = ~n39134 & ~n40323;
  assign n40325 = ~n38824 & ~n40324;
  assign n40326 = ~n38860 & ~n40325;
  assign n40327 = ~n38855 & ~n38900;
  assign n40328 = n38818 & n38838;
  assign n40329 = ~n39142 & ~n40328;
  assign n40330 = ~n40315 & n40329;
  assign n40331 = n38824 & ~n40330;
  assign n40332 = ~n38818 & n38892;
  assign n40333 = ~n40331 & ~n40332;
  assign n40334 = n40327 & n40333;
  assign n40335 = n40326 & n40334;
  assign n40336 = ~n38888 & ~n40335;
  assign n40337 = ~n38878 & ~n40093;
  assign n40338 = n38824 & ~n40337;
  assign n40339 = ~n40336 & ~n40338;
  assign n40340 = n40322 & n40339;
  assign n40341 = pi0913 & n40340;
  assign n40342 = ~pi0913 & ~n40340;
  assign po0926 = n40341 | n40342;
  assign n40344 = ~n39992 & n40187;
  assign n40345 = ~n40069 & ~n40344;
  assign n40346 = n40027 & ~n40345;
  assign n40347 = ~n39992 & n40005;
  assign n40348 = ~n40157 & ~n40347;
  assign n40349 = n40027 & ~n40348;
  assign n40350 = ~n40018 & n40036;
  assign n40351 = ~n40006 & ~n40350;
  assign n40352 = ~n40065 & n40351;
  assign n40353 = ~n40027 & ~n40352;
  assign n40354 = ~n40349 & ~n40353;
  assign n40355 = ~n40041 & ~n40054;
  assign n40356 = n40354 & n40355;
  assign n40357 = n40033 & ~n40356;
  assign n40358 = n40018 & n40157;
  assign n40359 = n40010 & ~n40018;
  assign n40360 = ~n40187 & ~n40359;
  assign n40361 = ~n40027 & ~n40360;
  assign n40362 = ~n40358 & ~n40361;
  assign n40363 = n40027 & n40037;
  assign n40364 = n40012 & ~n40363;
  assign n40365 = ~n40065 & n40364;
  assign n40366 = ~n40018 & ~n40365;
  assign n40367 = n40362 & ~n40366;
  assign n40368 = ~n40033 & ~n40367;
  assign n40369 = ~n40357 & ~n40368;
  assign n40370 = ~n39992 & ~n39998;
  assign n40371 = n40058 & n40370;
  assign n40372 = n40369 & ~n40371;
  assign n40373 = ~n40346 & n40372;
  assign n40374 = ~pi0876 & ~n40373;
  assign n40375 = pi0876 & ~n40346;
  assign n40376 = n40369 & n40375;
  assign n40377 = ~n40371 & n40376;
  assign po0927 = n40374 | n40377;
  assign n40379 = ~n40037 & ~n40164;
  assign n40380 = n40034 & ~n40379;
  assign n40381 = n39992 & n40018;
  assign n40382 = ~n40005 & n40381;
  assign n40383 = ~n40033 & n40382;
  assign n40384 = n40027 & n40050;
  assign n40385 = n40005 & n40384;
  assign n40386 = n39992 & n40058;
  assign n40387 = ~n40009 & n40386;
  assign n40388 = ~n40385 & ~n40387;
  assign n40389 = ~n40383 & n40388;
  assign n40390 = ~n40187 & ~n40189;
  assign n40391 = n40027 & ~n40390;
  assign n40392 = ~n40161 & ~n40391;
  assign n40393 = ~n40033 & ~n40392;
  assign n40394 = ~n40005 & ~n40370;
  assign n40395 = ~n40018 & ~n40394;
  assign n40396 = ~n40157 & ~n40395;
  assign n40397 = ~n40027 & ~n40396;
  assign n40398 = ~n40181 & ~n40397;
  assign n40399 = n40018 & n40065;
  assign n40400 = ~n40009 & n40019;
  assign n40401 = n40018 & ~n40394;
  assign n40402 = ~n40400 & ~n40401;
  assign n40403 = n40027 & ~n40402;
  assign n40404 = ~n40399 & ~n40403;
  assign n40405 = n40398 & n40404;
  assign n40406 = n40033 & ~n40405;
  assign n40407 = ~n40393 & ~n40406;
  assign n40408 = n40389 & n40407;
  assign n40409 = ~n40380 & n40408;
  assign n40410 = pi0883 & ~n40409;
  assign n40411 = ~pi0883 & n40389;
  assign n40412 = ~n40380 & n40411;
  assign n40413 = n40407 & n40412;
  assign po0928 = n40410 | n40413;
  assign n40415 = ~n39689 & ~n39809;
  assign n40416 = ~n39789 & n40415;
  assign n40417 = n39696 & ~n40416;
  assign n40418 = ~n39710 & ~n39736;
  assign n40419 = ~n39705 & ~n39797;
  assign n40420 = ~n39680 & ~n39802;
  assign n40421 = ~n39696 & ~n40420;
  assign n40422 = ~n39776 & ~n40421;
  assign n40423 = n40419 & n40422;
  assign n40424 = n39653 & ~n40423;
  assign n40425 = n39665 & n39678;
  assign n40426 = ~n39865 & ~n40425;
  assign n40427 = n39659 & ~n40426;
  assign n40428 = ~n39716 & ~n39720;
  assign n40429 = ~n39696 & ~n40428;
  assign n40430 = n39659 & n39678;
  assign n40431 = ~n39687 & ~n40430;
  assign n40432 = ~n39679 & n40431;
  assign n40433 = n39696 & ~n40432;
  assign n40434 = ~n40429 & ~n40433;
  assign n40435 = ~n40427 & n40434;
  assign n40436 = ~n39653 & ~n40435;
  assign n40437 = ~n40424 & ~n40436;
  assign n40438 = n40418 & n40437;
  assign n40439 = ~n40417 & n40438;
  assign n40440 = ~pi0892 & ~n40439;
  assign n40441 = pi0892 & n40418;
  assign n40442 = ~n40417 & n40441;
  assign n40443 = n40437 & n40442;
  assign po0929 = n40440 | n40443;
  assign n40445 = pi3802 & pi9040;
  assign n40446 = pi3815 & ~pi9040;
  assign n40447 = ~n40445 & ~n40446;
  assign n40448 = pi0893 & n40447;
  assign n40449 = ~pi0893 & ~n40447;
  assign n40450 = ~n40448 & ~n40449;
  assign n40451 = pi3801 & pi9040;
  assign n40452 = pi3803 & ~pi9040;
  assign n40453 = ~n40451 & ~n40452;
  assign n40454 = ~pi0895 & n40453;
  assign n40455 = pi0895 & ~n40453;
  assign n40456 = ~n40454 & ~n40455;
  assign n40457 = pi3806 & pi9040;
  assign n40458 = pi3794 & ~pi9040;
  assign n40459 = ~n40457 & ~n40458;
  assign n40460 = ~pi0921 & ~n40459;
  assign n40461 = pi0921 & ~n40457;
  assign n40462 = ~n40458 & n40461;
  assign n40463 = ~n40460 & ~n40462;
  assign n40464 = pi3830 & pi9040;
  assign n40465 = pi3835 & ~pi9040;
  assign n40466 = ~n40464 & ~n40465;
  assign n40467 = ~pi0891 & n40466;
  assign n40468 = pi0891 & ~n40466;
  assign n40469 = ~n40467 & ~n40468;
  assign n40470 = n40463 & ~n40469;
  assign n40471 = n40456 & n40470;
  assign n40472 = pi3787 & pi9040;
  assign n40473 = pi3790 & ~pi9040;
  assign n40474 = ~n40472 & ~n40473;
  assign n40475 = ~pi0911 & n40474;
  assign n40476 = pi0911 & ~n40474;
  assign n40477 = ~n40475 & ~n40476;
  assign n40478 = n40471 & n40477;
  assign n40479 = ~n40463 & n40469;
  assign n40480 = n40456 & n40477;
  assign n40481 = n40479 & n40480;
  assign n40482 = ~n40478 & ~n40481;
  assign n40483 = ~n40456 & ~n40477;
  assign n40484 = n40479 & n40483;
  assign n40485 = n40463 & n40469;
  assign n40486 = n40456 & n40485;
  assign n40487 = ~n40477 & n40486;
  assign n40488 = ~n40484 & ~n40487;
  assign n40489 = n40482 & n40488;
  assign n40490 = n40450 & ~n40489;
  assign n40491 = n40456 & ~n40477;
  assign n40492 = ~n40469 & n40491;
  assign n40493 = ~n40463 & n40492;
  assign n40494 = ~n40486 & ~n40493;
  assign n40495 = n40450 & ~n40494;
  assign n40496 = ~n40469 & n40477;
  assign n40497 = ~n40450 & n40496;
  assign n40498 = ~n40456 & n40463;
  assign n40499 = ~n40477 & n40479;
  assign n40500 = ~n40498 & ~n40499;
  assign n40501 = ~n40450 & ~n40500;
  assign n40502 = ~n40497 & ~n40501;
  assign n40503 = ~n40463 & ~n40469;
  assign n40504 = ~n40456 & n40503;
  assign n40505 = n40477 & n40504;
  assign n40506 = n40502 & ~n40505;
  assign n40507 = ~n40469 & n40498;
  assign n40508 = ~n40477 & n40507;
  assign n40509 = n40506 & ~n40508;
  assign n40510 = ~n40495 & n40509;
  assign n40511 = pi3790 & pi9040;
  assign n40512 = pi3802 & ~pi9040;
  assign n40513 = ~n40511 & ~n40512;
  assign n40514 = ~pi0927 & n40513;
  assign n40515 = pi0927 & ~n40513;
  assign n40516 = ~n40514 & ~n40515;
  assign n40517 = ~n40510 & n40516;
  assign n40518 = n40456 & ~n40469;
  assign n40519 = ~n40450 & ~n40477;
  assign n40520 = ~n40516 & n40519;
  assign n40521 = n40518 & n40520;
  assign n40522 = n40469 & n40480;
  assign n40523 = ~n40450 & ~n40522;
  assign n40524 = ~n40463 & n40483;
  assign n40525 = ~n40470 & ~n40518;
  assign n40526 = n40477 & ~n40525;
  assign n40527 = ~n40456 & n40479;
  assign n40528 = n40450 & ~n40527;
  assign n40529 = ~n40526 & n40528;
  assign n40530 = ~n40524 & n40529;
  assign n40531 = ~n40523 & ~n40530;
  assign n40532 = ~n40456 & n40485;
  assign n40533 = ~n40477 & n40532;
  assign n40534 = ~n40531 & ~n40533;
  assign n40535 = ~n40516 & ~n40534;
  assign n40536 = ~n40521 & ~n40535;
  assign n40537 = ~n40517 & n40536;
  assign n40538 = ~n40490 & n40537;
  assign n40539 = ~n40450 & n40505;
  assign n40540 = n40538 & ~n40539;
  assign n40541 = pi0928 & ~n40540;
  assign n40542 = ~pi0928 & ~n40539;
  assign n40543 = n40537 & n40542;
  assign n40544 = ~n40490 & n40543;
  assign po0949 = n40541 | n40544;
  assign n40546 = pi3859 & ~pi9040;
  assign n40547 = pi3797 & pi9040;
  assign n40548 = ~n40546 & ~n40547;
  assign n40549 = ~pi0917 & ~n40548;
  assign n40550 = pi0917 & n40548;
  assign n40551 = ~n40549 & ~n40550;
  assign n40552 = pi3795 & pi9040;
  assign n40553 = pi3796 & ~pi9040;
  assign n40554 = ~n40552 & ~n40553;
  assign n40555 = ~pi0910 & n40554;
  assign n40556 = pi0910 & ~n40554;
  assign n40557 = ~n40555 & ~n40556;
  assign n40558 = pi3827 & pi9040;
  assign n40559 = pi3805 & ~pi9040;
  assign n40560 = ~n40558 & ~n40559;
  assign n40561 = pi0912 & n40560;
  assign n40562 = ~pi0912 & ~n40560;
  assign n40563 = ~n40561 & ~n40562;
  assign n40564 = pi3859 & pi9040;
  assign n40565 = pi3832 & ~pi9040;
  assign n40566 = ~n40564 & ~n40565;
  assign n40567 = ~pi0922 & n40566;
  assign n40568 = pi0922 & ~n40566;
  assign n40569 = ~n40567 & ~n40568;
  assign n40570 = pi3805 & pi9040;
  assign n40571 = pi3854 & ~pi9040;
  assign n40572 = ~n40570 & ~n40571;
  assign n40573 = ~pi0904 & ~n40572;
  assign n40574 = pi0904 & ~n40570;
  assign n40575 = ~n40571 & n40574;
  assign n40576 = ~n40573 & ~n40575;
  assign n40577 = ~n40569 & ~n40576;
  assign n40578 = n40563 & n40577;
  assign n40579 = pi3831 & pi9040;
  assign n40580 = pi3812 & ~pi9040;
  assign n40581 = ~n40579 & ~n40580;
  assign n40582 = ~pi0898 & n40581;
  assign n40583 = pi0898 & ~n40581;
  assign n40584 = ~n40582 & ~n40583;
  assign n40585 = n40576 & ~n40584;
  assign n40586 = ~n40569 & n40585;
  assign n40587 = ~n40578 & ~n40586;
  assign n40588 = n40576 & n40584;
  assign n40589 = n40569 & n40588;
  assign n40590 = ~n40563 & n40589;
  assign n40591 = n40587 & ~n40590;
  assign n40592 = ~n40557 & ~n40591;
  assign n40593 = n40569 & n40576;
  assign n40594 = ~n40563 & n40593;
  assign n40595 = ~n40584 & n40594;
  assign n40596 = ~n40576 & ~n40584;
  assign n40597 = ~n40569 & n40596;
  assign n40598 = ~n40563 & n40597;
  assign n40599 = n40569 & ~n40576;
  assign n40600 = ~n40588 & ~n40599;
  assign n40601 = n40563 & ~n40600;
  assign n40602 = ~n40598 & ~n40601;
  assign n40603 = ~n40595 & n40602;
  assign n40604 = n40557 & ~n40603;
  assign n40605 = ~n40592 & ~n40604;
  assign n40606 = n40551 & ~n40605;
  assign n40607 = ~n40557 & ~n40563;
  assign n40608 = ~n40576 & n40607;
  assign n40609 = n40557 & ~n40563;
  assign n40610 = n40588 & n40609;
  assign n40611 = ~n40563 & ~n40569;
  assign n40612 = n40576 & n40611;
  assign n40613 = ~n40578 & ~n40612;
  assign n40614 = n40557 & ~n40613;
  assign n40615 = ~n40610 & ~n40614;
  assign n40616 = ~n40569 & n40588;
  assign n40617 = ~n40563 & n40616;
  assign n40618 = ~n40584 & n40593;
  assign n40619 = n40563 & n40618;
  assign n40620 = ~n40617 & ~n40619;
  assign n40621 = ~n40557 & n40563;
  assign n40622 = n40593 & n40621;
  assign n40623 = n40569 & n40596;
  assign n40624 = ~n40557 & n40623;
  assign n40625 = ~n40622 & ~n40624;
  assign n40626 = n40620 & n40625;
  assign n40627 = n40615 & n40626;
  assign n40628 = ~n40608 & n40627;
  assign n40629 = ~n40551 & ~n40628;
  assign n40630 = ~n40576 & n40584;
  assign n40631 = n40569 & n40630;
  assign n40632 = n40609 & n40631;
  assign n40633 = ~n40569 & n40610;
  assign n40634 = ~n40632 & ~n40633;
  assign n40635 = ~n40584 & n40599;
  assign n40636 = ~n40563 & n40635;
  assign n40637 = ~n40557 & n40636;
  assign n40638 = n40634 & ~n40637;
  assign n40639 = n40563 & n40585;
  assign n40640 = ~n40569 & n40630;
  assign n40641 = ~n40563 & n40640;
  assign n40642 = ~n40639 & ~n40641;
  assign n40643 = ~n40557 & ~n40642;
  assign n40644 = n40638 & ~n40643;
  assign n40645 = ~n40629 & n40644;
  assign n40646 = ~n40606 & n40645;
  assign n40647 = pi0947 & n40646;
  assign n40648 = ~pi0947 & ~n40646;
  assign po0956 = n40647 | n40648;
  assign n40650 = ~n40551 & n40557;
  assign n40651 = ~n40563 & n40577;
  assign n40652 = n40563 & n40616;
  assign n40653 = ~n40563 & n40585;
  assign n40654 = ~n40652 & ~n40653;
  assign n40655 = ~n40651 & n40654;
  assign n40656 = n40650 & ~n40655;
  assign n40657 = ~n40563 & n40569;
  assign n40658 = n40584 & n40657;
  assign n40659 = n40563 & n40640;
  assign n40660 = ~n40658 & ~n40659;
  assign n40661 = ~n40586 & ~n40589;
  assign n40662 = n40660 & n40661;
  assign n40663 = ~n40557 & ~n40662;
  assign n40664 = n40563 & n40623;
  assign n40665 = ~n40663 & ~n40664;
  assign n40666 = ~n40551 & ~n40665;
  assign n40667 = ~n40656 & ~n40666;
  assign n40668 = ~n40569 & n40607;
  assign n40669 = ~n40584 & n40668;
  assign n40670 = ~n40590 & ~n40669;
  assign n40671 = ~n40585 & ~n40630;
  assign n40672 = n40563 & ~n40671;
  assign n40673 = ~n40631 & ~n40672;
  assign n40674 = n40557 & ~n40673;
  assign n40675 = ~n40597 & ~n40651;
  assign n40676 = ~n40652 & n40675;
  assign n40677 = ~n40557 & ~n40676;
  assign n40678 = ~n40674 & ~n40677;
  assign n40679 = n40584 & n40599;
  assign n40680 = n40563 & n40679;
  assign n40681 = ~n40619 & ~n40680;
  assign n40682 = ~n40636 & n40681;
  assign n40683 = ~n40610 & n40682;
  assign n40684 = n40678 & n40683;
  assign n40685 = n40551 & ~n40684;
  assign n40686 = n40670 & ~n40685;
  assign n40687 = n40667 & n40686;
  assign n40688 = pi0943 & ~n40687;
  assign n40689 = ~pi0943 & n40670;
  assign n40690 = n40667 & n40689;
  assign n40691 = ~n40685 & n40690;
  assign po0958 = n40688 | n40691;
  assign n40693 = pi3804 & pi9040;
  assign n40694 = pi3817 & ~pi9040;
  assign n40695 = ~n40693 & ~n40694;
  assign n40696 = ~pi0925 & n40695;
  assign n40697 = pi0925 & ~n40695;
  assign n40698 = ~n40696 & ~n40697;
  assign n40699 = pi3794 & pi9040;
  assign n40700 = pi3830 & ~pi9040;
  assign n40701 = ~n40699 & ~n40700;
  assign n40702 = pi0899 & n40701;
  assign n40703 = ~pi0899 & ~n40701;
  assign n40704 = ~n40702 & ~n40703;
  assign n40705 = pi3803 & pi9040;
  assign n40706 = pi3804 & ~pi9040;
  assign n40707 = ~n40705 & ~n40706;
  assign n40708 = ~pi0898 & ~n40707;
  assign n40709 = pi0898 & ~n40705;
  assign n40710 = ~n40706 & n40709;
  assign n40711 = ~n40708 & ~n40710;
  assign n40712 = pi3799 & pi9040;
  assign n40713 = pi3827 & ~pi9040;
  assign n40714 = ~n40712 & ~n40713;
  assign n40715 = ~pi0917 & n40714;
  assign n40716 = pi0917 & ~n40714;
  assign n40717 = ~n40715 & ~n40716;
  assign n40718 = pi3835 & pi9040;
  assign n40719 = pi3806 & ~pi9040;
  assign n40720 = ~n40718 & ~n40719;
  assign n40721 = ~pi0895 & n40720;
  assign n40722 = pi0895 & ~n40720;
  assign n40723 = ~n40721 & ~n40722;
  assign n40724 = n40717 & ~n40723;
  assign n40725 = ~n40711 & n40724;
  assign n40726 = n40704 & n40725;
  assign n40727 = ~n40717 & n40723;
  assign n40728 = ~n40711 & n40727;
  assign n40729 = n40717 & n40723;
  assign n40730 = n40711 & n40729;
  assign n40731 = n40704 & n40730;
  assign n40732 = ~n40728 & ~n40731;
  assign n40733 = ~n40726 & n40732;
  assign n40734 = ~n40698 & ~n40733;
  assign n40735 = n40711 & n40717;
  assign n40736 = ~n40704 & n40735;
  assign n40737 = n40711 & ~n40717;
  assign n40738 = n40704 & n40737;
  assign n40739 = ~n40736 & ~n40738;
  assign n40740 = n40698 & ~n40739;
  assign n40741 = ~n40734 & ~n40740;
  assign n40742 = pi3822 & pi9040;
  assign n40743 = pi3838 & ~pi9040;
  assign n40744 = ~n40742 & ~n40743;
  assign n40745 = ~pi0891 & ~n40744;
  assign n40746 = pi0891 & n40744;
  assign n40747 = ~n40745 & ~n40746;
  assign n40748 = n40711 & n40724;
  assign n40749 = ~n40711 & ~n40723;
  assign n40750 = ~n40704 & n40749;
  assign n40751 = ~n40717 & n40750;
  assign n40752 = ~n40748 & ~n40751;
  assign n40753 = n40698 & ~n40752;
  assign n40754 = ~n40704 & ~n40711;
  assign n40755 = n40723 & n40754;
  assign n40756 = n40717 & n40755;
  assign n40757 = ~n40726 & ~n40756;
  assign n40758 = n40704 & ~n40711;
  assign n40759 = ~n40717 & n40758;
  assign n40760 = ~n40717 & ~n40723;
  assign n40761 = n40711 & n40760;
  assign n40762 = ~n40704 & n40761;
  assign n40763 = ~n40759 & ~n40762;
  assign n40764 = ~n40698 & ~n40763;
  assign n40765 = n40757 & ~n40764;
  assign n40766 = ~n40753 & n40765;
  assign n40767 = n40747 & ~n40766;
  assign n40768 = n40698 & ~n40704;
  assign n40769 = n40724 & n40768;
  assign n40770 = n40711 & n40727;
  assign n40771 = n40723 & n40758;
  assign n40772 = n40717 & n40771;
  assign n40773 = ~n40770 & ~n40772;
  assign n40774 = n40704 & n40760;
  assign n40775 = n40773 & ~n40774;
  assign n40776 = n40698 & ~n40775;
  assign n40777 = ~n40711 & ~n40717;
  assign n40778 = ~n40698 & ~n40704;
  assign n40779 = n40777 & n40778;
  assign n40780 = ~n40704 & n40728;
  assign n40781 = ~n40779 & ~n40780;
  assign n40782 = ~n40776 & n40781;
  assign n40783 = ~n40769 & n40782;
  assign n40784 = ~n40704 & n40748;
  assign n40785 = n40704 & n40761;
  assign n40786 = ~n40784 & ~n40785;
  assign n40787 = n40783 & n40786;
  assign n40788 = ~n40747 & ~n40787;
  assign n40789 = ~n40711 & n40723;
  assign n40790 = ~n40698 & n40789;
  assign n40791 = ~n40704 & n40790;
  assign n40792 = ~n40788 & ~n40791;
  assign n40793 = ~n40767 & n40792;
  assign n40794 = n40741 & n40793;
  assign n40795 = ~pi0930 & ~n40794;
  assign n40796 = pi0930 & n40794;
  assign po0964 = n40795 | n40796;
  assign n40798 = pi3792 & pi9040;
  assign n40799 = pi3836 & ~pi9040;
  assign n40800 = ~n40798 & ~n40799;
  assign n40801 = pi0926 & n40800;
  assign n40802 = ~pi0926 & ~n40800;
  assign n40803 = ~n40801 & ~n40802;
  assign n40804 = pi3825 & pi9040;
  assign n40805 = pi3826 & ~pi9040;
  assign n40806 = ~n40804 & ~n40805;
  assign n40807 = ~pi0905 & ~n40806;
  assign n40808 = pi0905 & ~n40804;
  assign n40809 = ~n40805 & n40808;
  assign n40810 = ~n40807 & ~n40809;
  assign n40811 = pi3826 & pi9040;
  assign n40812 = pi3833 & ~pi9040;
  assign n40813 = ~n40811 & ~n40812;
  assign n40814 = pi0918 & n40813;
  assign n40815 = ~pi0918 & ~n40813;
  assign n40816 = ~n40814 & ~n40815;
  assign n40817 = n40810 & ~n40816;
  assign n40818 = pi3784 & pi9040;
  assign n40819 = pi3834 & ~pi9040;
  assign n40820 = ~n40818 & ~n40819;
  assign n40821 = pi0915 & n40820;
  assign n40822 = ~pi0915 & ~n40820;
  assign n40823 = ~n40821 & ~n40822;
  assign n40824 = pi3829 & pi9040;
  assign n40825 = pi3837 & ~pi9040;
  assign n40826 = ~n40824 & ~n40825;
  assign n40827 = pi0890 & n40826;
  assign n40828 = ~pi0890 & ~n40826;
  assign n40829 = ~n40827 & ~n40828;
  assign n40830 = n40823 & n40829;
  assign n40831 = n40817 & n40830;
  assign n40832 = n40823 & ~n40829;
  assign n40833 = ~n40810 & n40832;
  assign n40834 = ~n40831 & ~n40833;
  assign n40835 = ~n40803 & ~n40834;
  assign n40836 = pi3818 & pi9040;
  assign n40837 = pi3829 & ~pi9040;
  assign n40838 = ~n40836 & ~n40837;
  assign n40839 = ~pi0909 & ~n40838;
  assign n40840 = pi0909 & n40838;
  assign n40841 = ~n40839 & ~n40840;
  assign n40842 = n40803 & ~n40823;
  assign n40843 = n40810 & n40842;
  assign n40844 = n40817 & ~n40829;
  assign n40845 = n40810 & n40816;
  assign n40846 = n40829 & n40845;
  assign n40847 = ~n40844 & ~n40846;
  assign n40848 = ~n40810 & ~n40816;
  assign n40849 = n40829 & n40848;
  assign n40850 = n40823 & n40849;
  assign n40851 = n40847 & ~n40850;
  assign n40852 = n40803 & ~n40851;
  assign n40853 = ~n40843 & ~n40852;
  assign n40854 = ~n40810 & n40816;
  assign n40855 = ~n40829 & n40854;
  assign n40856 = n40823 & n40855;
  assign n40857 = n40853 & ~n40856;
  assign n40858 = ~n40823 & n40848;
  assign n40859 = ~n40810 & n40829;
  assign n40860 = n40816 & n40859;
  assign n40861 = ~n40858 & ~n40860;
  assign n40862 = ~n40803 & ~n40861;
  assign n40863 = ~n40829 & n40845;
  assign n40864 = ~n40823 & n40863;
  assign n40865 = ~n40862 & ~n40864;
  assign n40866 = n40857 & n40865;
  assign n40867 = n40841 & ~n40866;
  assign n40868 = ~n40835 & ~n40867;
  assign n40869 = n40803 & ~n40841;
  assign n40870 = ~n40861 & n40869;
  assign n40871 = ~n40829 & n40848;
  assign n40872 = ~n40863 & ~n40871;
  assign n40873 = n40823 & ~n40872;
  assign n40874 = ~n40831 & ~n40873;
  assign n40875 = ~n40841 & ~n40874;
  assign n40876 = ~n40870 & ~n40875;
  assign n40877 = ~n40803 & ~n40841;
  assign n40878 = n40817 & ~n40823;
  assign n40879 = ~n40855 & ~n40878;
  assign n40880 = n40810 & n40829;
  assign n40881 = n40879 & ~n40880;
  assign n40882 = n40877 & ~n40881;
  assign n40883 = n40876 & ~n40882;
  assign n40884 = n40868 & n40883;
  assign n40885 = ~pi0937 & ~n40884;
  assign n40886 = pi0937 & n40876;
  assign n40887 = n40868 & n40886;
  assign n40888 = ~n40882 & n40887;
  assign po0965 = n40885 | n40888;
  assign n40890 = ~n40597 & ~n40631;
  assign n40891 = n40557 & ~n40890;
  assign n40892 = n40563 & n40586;
  assign n40893 = ~n40891 & ~n40892;
  assign n40894 = n40563 & n40576;
  assign n40895 = ~n40593 & ~n40894;
  assign n40896 = ~n40640 & n40895;
  assign n40897 = ~n40557 & ~n40896;
  assign n40898 = n40893 & ~n40897;
  assign n40899 = ~n40551 & ~n40898;
  assign n40900 = ~n40563 & n40618;
  assign n40901 = n40557 & n40900;
  assign n40902 = ~n40633 & ~n40901;
  assign n40903 = ~n40637 & n40902;
  assign n40904 = ~n40557 & n40576;
  assign n40905 = n40611 & n40904;
  assign n40906 = n40563 & n40597;
  assign n40907 = n40557 & n40593;
  assign n40908 = ~n40906 & ~n40907;
  assign n40909 = ~n40680 & n40908;
  assign n40910 = ~n40905 & n40909;
  assign n40911 = n40584 & n40611;
  assign n40912 = ~n40636 & ~n40911;
  assign n40913 = n40910 & n40912;
  assign n40914 = ~n40624 & n40913;
  assign n40915 = n40551 & ~n40914;
  assign n40916 = n40903 & ~n40915;
  assign n40917 = ~n40899 & n40916;
  assign n40918 = ~pi0941 & ~n40917;
  assign n40919 = pi0941 & n40903;
  assign n40920 = ~n40899 & n40919;
  assign n40921 = ~n40915 & n40920;
  assign po0966 = n40918 | n40921;
  assign n40923 = pi3832 & pi9040;
  assign n40924 = pi3798 & ~pi9040;
  assign n40925 = ~n40923 & ~n40924;
  assign n40926 = pi0904 & n40925;
  assign n40927 = ~pi0904 & ~n40925;
  assign n40928 = ~n40926 & ~n40927;
  assign n40929 = pi3848 & pi9040;
  assign n40930 = pi3858 & ~pi9040;
  assign n40931 = ~n40929 & ~n40930;
  assign n40932 = pi0919 & n40931;
  assign n40933 = ~pi0919 & ~n40931;
  assign n40934 = ~n40932 & ~n40933;
  assign n40935 = pi3838 & pi9040;
  assign n40936 = pi3831 & ~pi9040;
  assign n40937 = ~n40935 & ~n40936;
  assign n40938 = ~pi0916 & ~n40937;
  assign n40939 = pi0916 & ~n40935;
  assign n40940 = ~n40936 & n40939;
  assign n40941 = ~n40938 & ~n40940;
  assign n40942 = pi3796 & pi9040;
  assign n40943 = pi3848 & ~pi9040;
  assign n40944 = ~n40942 & ~n40943;
  assign n40945 = ~pi0896 & n40944;
  assign n40946 = pi0896 & ~n40944;
  assign n40947 = ~n40945 & ~n40946;
  assign n40948 = pi3812 & pi9040;
  assign n40949 = pi3822 & ~pi9040;
  assign n40950 = ~n40948 & ~n40949;
  assign n40951 = pi0922 & n40950;
  assign n40952 = ~pi0922 & ~n40950;
  assign n40953 = ~n40951 & ~n40952;
  assign n40954 = ~n40947 & ~n40953;
  assign n40955 = n40941 & n40954;
  assign n40956 = n40934 & n40955;
  assign n40957 = ~n40934 & ~n40947;
  assign n40958 = n40953 & n40957;
  assign n40959 = pi3854 & pi9040;
  assign n40960 = pi3799 & ~pi9040;
  assign n40961 = ~n40959 & ~n40960;
  assign n40962 = pi0897 & n40961;
  assign n40963 = ~pi0897 & ~n40961;
  assign n40964 = ~n40962 & ~n40963;
  assign n40965 = ~n40941 & n40957;
  assign n40966 = n40941 & n40953;
  assign n40967 = n40947 & n40966;
  assign n40968 = ~n40965 & ~n40967;
  assign n40969 = ~n40964 & ~n40968;
  assign n40970 = ~n40958 & ~n40969;
  assign n40971 = ~n40947 & n40966;
  assign n40972 = ~n40941 & n40947;
  assign n40973 = n40947 & ~n40953;
  assign n40974 = ~n40934 & n40973;
  assign n40975 = ~n40941 & ~n40953;
  assign n40976 = n40934 & n40975;
  assign n40977 = ~n40974 & ~n40976;
  assign n40978 = ~n40972 & n40977;
  assign n40979 = ~n40971 & n40978;
  assign n40980 = n40964 & ~n40979;
  assign n40981 = n40970 & ~n40980;
  assign n40982 = ~n40956 & n40981;
  assign n40983 = n40928 & ~n40982;
  assign n40984 = ~n40941 & n40953;
  assign n40985 = n40947 & n40984;
  assign n40986 = ~n40934 & n40985;
  assign n40987 = n40947 & n40975;
  assign n40988 = n40934 & n40987;
  assign n40989 = ~n40956 & ~n40988;
  assign n40990 = ~n40986 & n40989;
  assign n40991 = n40964 & ~n40990;
  assign n40992 = ~n40983 & ~n40991;
  assign n40993 = ~n40934 & n40971;
  assign n40994 = n40941 & n40947;
  assign n40995 = ~n40964 & n40994;
  assign n40996 = n40934 & n40995;
  assign n40997 = ~n40947 & n40984;
  assign n40998 = n40934 & n40997;
  assign n40999 = n40954 & n40964;
  assign n41000 = ~n40934 & n40999;
  assign n41001 = ~n40998 & ~n41000;
  assign n41002 = ~n40941 & ~n40947;
  assign n41003 = n40934 & n41002;
  assign n41004 = n40941 & ~n40953;
  assign n41005 = n40947 & n41004;
  assign n41006 = ~n41003 & ~n41005;
  assign n41007 = ~n40964 & ~n41006;
  assign n41008 = ~n40964 & n40972;
  assign n41009 = ~n40934 & n41008;
  assign n41010 = ~n41007 & ~n41009;
  assign n41011 = n41001 & n41010;
  assign n41012 = ~n40928 & ~n41011;
  assign n41013 = ~n40996 & ~n41012;
  assign n41014 = ~n40993 & n41013;
  assign n41015 = n40992 & n41014;
  assign n41016 = ~pi0956 & ~n41015;
  assign n41017 = ~n40983 & ~n40993;
  assign n41018 = ~n40991 & n41017;
  assign n41019 = n41013 & n41018;
  assign n41020 = pi0956 & n41019;
  assign po0967 = n41016 | n41020;
  assign n41022 = pi3793 & pi9040;
  assign n41023 = pi3821 & ~pi9040;
  assign n41024 = ~n41022 & ~n41023;
  assign n41025 = ~pi0905 & ~n41024;
  assign n41026 = pi0905 & n41024;
  assign n41027 = ~n41025 & ~n41026;
  assign n41028 = pi3833 & pi9040;
  assign n41029 = pi3819 & ~pi9040;
  assign n41030 = ~n41028 & ~n41029;
  assign n41031 = ~pi0921 & n41030;
  assign n41032 = pi0921 & ~n41030;
  assign n41033 = ~n41031 & ~n41032;
  assign n41034 = pi3788 & pi9040;
  assign n41035 = pi3818 & ~pi9040;
  assign n41036 = ~n41034 & ~n41035;
  assign n41037 = ~pi0927 & n41036;
  assign n41038 = pi0927 & ~n41036;
  assign n41039 = ~n41037 & ~n41038;
  assign n41040 = pi3791 & pi9040;
  assign n41041 = pi3811 & ~pi9040;
  assign n41042 = ~n41040 & ~n41041;
  assign n41043 = ~pi0890 & n41042;
  assign n41044 = pi0890 & ~n41042;
  assign n41045 = ~n41043 & ~n41044;
  assign n41046 = n41039 & ~n41045;
  assign n41047 = pi3786 & pi9040;
  assign n41048 = pi3808 & ~pi9040;
  assign n41049 = ~n41047 & ~n41048;
  assign n41050 = pi0901 & n41049;
  assign n41051 = ~pi0901 & ~n41049;
  assign n41052 = ~n41050 & ~n41051;
  assign n41053 = pi3819 & pi9040;
  assign n41054 = pi3825 & ~pi9040;
  assign n41055 = ~n41053 & ~n41054;
  assign n41056 = ~pi0923 & n41055;
  assign n41057 = pi0923 & ~n41055;
  assign n41058 = ~n41056 & ~n41057;
  assign n41059 = n41052 & ~n41058;
  assign n41060 = n41046 & n41059;
  assign n41061 = ~n41033 & n41060;
  assign n41062 = ~n41052 & ~n41058;
  assign n41063 = ~n41039 & ~n41045;
  assign n41064 = n41062 & n41063;
  assign n41065 = ~n41039 & n41045;
  assign n41066 = ~n41033 & n41065;
  assign n41067 = ~n41058 & n41066;
  assign n41068 = n41052 & n41067;
  assign n41069 = ~n41033 & ~n41052;
  assign n41070 = n41045 & n41069;
  assign n41071 = n41039 & n41070;
  assign n41072 = ~n41068 & ~n41071;
  assign n41073 = ~n41064 & n41072;
  assign n41074 = ~n41061 & n41073;
  assign n41075 = n41033 & ~n41052;
  assign n41076 = ~n41045 & n41075;
  assign n41077 = ~n41039 & n41076;
  assign n41078 = n41074 & ~n41077;
  assign n41079 = ~n41027 & ~n41078;
  assign n41080 = ~n41033 & ~n41039;
  assign n41081 = ~n41045 & n41080;
  assign n41082 = n41052 & n41081;
  assign n41083 = ~n41070 & ~n41082;
  assign n41084 = n41033 & n41046;
  assign n41085 = n41052 & n41084;
  assign n41086 = n41083 & ~n41085;
  assign n41087 = n41058 & ~n41086;
  assign n41088 = n41033 & n41045;
  assign n41089 = ~n41039 & n41088;
  assign n41090 = n41058 & n41089;
  assign n41091 = n41052 & n41090;
  assign n41092 = n41039 & n41069;
  assign n41093 = n41039 & n41045;
  assign n41094 = ~n41052 & n41093;
  assign n41095 = ~n41092 & ~n41094;
  assign n41096 = n41058 & ~n41095;
  assign n41097 = ~n41091 & ~n41096;
  assign n41098 = ~n41027 & ~n41097;
  assign n41099 = ~n41087 & ~n41098;
  assign n41100 = ~n41079 & n41099;
  assign n41101 = n41033 & n41052;
  assign n41102 = ~n41058 & n41101;
  assign n41103 = n41093 & n41102;
  assign n41104 = n41033 & ~n41039;
  assign n41105 = n41062 & n41104;
  assign n41106 = n41058 & n41080;
  assign n41107 = n41039 & n41052;
  assign n41108 = n41033 & n41107;
  assign n41109 = ~n41084 & ~n41108;
  assign n41110 = ~n41106 & n41109;
  assign n41111 = ~n41052 & n41089;
  assign n41112 = n41110 & ~n41111;
  assign n41113 = n41046 & ~n41058;
  assign n41114 = ~n41052 & n41113;
  assign n41115 = n41033 & ~n41045;
  assign n41116 = n41052 & n41093;
  assign n41117 = ~n41115 & ~n41116;
  assign n41118 = ~n41058 & ~n41117;
  assign n41119 = ~n41114 & ~n41118;
  assign n41120 = n41112 & n41119;
  assign n41121 = n41027 & ~n41120;
  assign n41122 = ~n41105 & ~n41121;
  assign n41123 = ~n41103 & n41122;
  assign n41124 = n41100 & n41123;
  assign n41125 = pi0931 & n41124;
  assign n41126 = ~pi0931 & ~n41124;
  assign po0968 = n41125 | n41126;
  assign n41128 = ~n40717 & n40771;
  assign n41129 = ~n40737 & ~n40756;
  assign n41130 = ~n40698 & ~n41129;
  assign n41131 = ~n41128 & ~n41130;
  assign n41132 = ~n40751 & n41131;
  assign n41133 = n40698 & n40704;
  assign n41134 = n40725 & n41133;
  assign n41135 = ~n40784 & ~n41134;
  assign n41136 = ~n40731 & n41135;
  assign n41137 = n41132 & n41136;
  assign n41138 = n40747 & ~n41137;
  assign n41139 = ~n40711 & n40760;
  assign n41140 = n40704 & n41139;
  assign n41141 = ~n40772 & ~n41140;
  assign n41142 = ~n40704 & n40730;
  assign n41143 = ~n40780 & ~n41142;
  assign n41144 = n40711 & ~n40723;
  assign n41145 = n40704 & ~n40717;
  assign n41146 = ~n41144 & ~n41145;
  assign n41147 = ~n40789 & n41146;
  assign n41148 = n40698 & ~n41147;
  assign n41149 = ~n40698 & n40725;
  assign n41150 = n40704 & n40748;
  assign n41151 = ~n41149 & ~n41150;
  assign n41152 = ~n41148 & n41151;
  assign n41153 = n41143 & n41152;
  assign n41154 = n41141 & n41153;
  assign n41155 = ~n40747 & ~n41154;
  assign n41156 = ~n41138 & ~n41155;
  assign n41157 = pi0933 & ~n41156;
  assign n41158 = ~pi0933 & ~n41138;
  assign n41159 = ~n41155 & n41158;
  assign po0969 = n41157 | n41159;
  assign n41161 = pi3823 & pi9040;
  assign n41162 = pi3850 & ~pi9040;
  assign n41163 = ~n41161 & ~n41162;
  assign n41164 = ~pi0924 & n41163;
  assign n41165 = pi0924 & ~n41163;
  assign n41166 = ~n41164 & ~n41165;
  assign n41167 = pi3850 & pi9040;
  assign n41168 = pi3792 & ~pi9040;
  assign n41169 = ~n41167 & ~n41168;
  assign n41170 = ~pi0906 & n41169;
  assign n41171 = pi0906 & ~n41169;
  assign n41172 = ~n41170 & ~n41171;
  assign n41173 = pi3837 & pi9040;
  assign n41174 = pi3788 & ~pi9040;
  assign n41175 = ~n41173 & ~n41174;
  assign n41176 = ~pi0914 & ~n41175;
  assign n41177 = pi0914 & ~n41173;
  assign n41178 = ~n41174 & n41177;
  assign n41179 = ~n41176 & ~n41178;
  assign n41180 = pi3814 & pi9040;
  assign n41181 = pi3855 & ~pi9040;
  assign n41182 = ~n41180 & ~n41181;
  assign n41183 = ~pi0920 & ~n41182;
  assign n41184 = pi0920 & n41182;
  assign n41185 = ~n41183 & ~n41184;
  assign n41186 = pi3813 & pi9040;
  assign n41187 = pi3785 & ~pi9040;
  assign n41188 = ~n41186 & ~n41187;
  assign n41189 = ~pi0896 & ~n41188;
  assign n41190 = pi0896 & n41188;
  assign n41191 = ~n41189 & ~n41190;
  assign n41192 = ~n41185 & ~n41191;
  assign n41193 = ~n41179 & n41192;
  assign n41194 = n41172 & n41193;
  assign n41195 = n41185 & ~n41191;
  assign n41196 = ~n41179 & n41195;
  assign n41197 = ~n41172 & n41196;
  assign n41198 = ~n41194 & ~n41197;
  assign n41199 = ~n41166 & ~n41198;
  assign n41200 = ~pi0896 & n41188;
  assign n41201 = pi0896 & ~n41188;
  assign n41202 = ~n41200 & ~n41201;
  assign n41203 = n41172 & n41179;
  assign n41204 = ~n41202 & n41203;
  assign n41205 = ~n41185 & n41204;
  assign n41206 = n41166 & n41205;
  assign n41207 = pi3823 & ~pi9040;
  assign n41208 = pi3836 & pi9040;
  assign n41209 = ~n41207 & ~n41208;
  assign n41210 = ~pi0916 & ~n41209;
  assign n41211 = pi0916 & n41209;
  assign n41212 = ~n41210 & ~n41211;
  assign n41213 = n41179 & n41195;
  assign n41214 = ~n41166 & n41213;
  assign n41215 = ~n41205 & ~n41214;
  assign n41216 = n41172 & n41185;
  assign n41217 = ~n41179 & n41216;
  assign n41218 = ~n41185 & n41203;
  assign n41219 = ~n41217 & ~n41218;
  assign n41220 = n41166 & ~n41219;
  assign n41221 = n41166 & ~n41172;
  assign n41222 = n41192 & n41221;
  assign n41223 = ~n41179 & n41222;
  assign n41224 = ~n41172 & n41179;
  assign n41225 = ~n41202 & n41224;
  assign n41226 = n41185 & n41225;
  assign n41227 = ~n41185 & ~n41202;
  assign n41228 = ~n41179 & n41227;
  assign n41229 = ~n41166 & n41228;
  assign n41230 = ~n41226 & ~n41229;
  assign n41231 = ~n41223 & n41230;
  assign n41232 = ~n41220 & n41231;
  assign n41233 = n41215 & n41232;
  assign n41234 = n41212 & ~n41233;
  assign n41235 = n41172 & n41214;
  assign n41236 = ~n41234 & ~n41235;
  assign n41237 = ~n41206 & n41236;
  assign n41238 = ~n41199 & n41237;
  assign n41239 = ~n41166 & ~n41172;
  assign n41240 = n41179 & ~n41185;
  assign n41241 = n41239 & n41240;
  assign n41242 = ~n41166 & n41193;
  assign n41243 = ~n41241 & ~n41242;
  assign n41244 = n41185 & ~n41202;
  assign n41245 = n41179 & n41244;
  assign n41246 = ~n41166 & n41245;
  assign n41247 = ~n41179 & n41244;
  assign n41248 = n41172 & n41247;
  assign n41249 = ~n41246 & ~n41248;
  assign n41250 = n41179 & n41192;
  assign n41251 = ~n41172 & n41250;
  assign n41252 = ~n41194 & ~n41251;
  assign n41253 = ~n41172 & n41195;
  assign n41254 = ~n41179 & n41191;
  assign n41255 = ~n41253 & ~n41254;
  assign n41256 = n41166 & ~n41255;
  assign n41257 = n41252 & ~n41256;
  assign n41258 = n41249 & n41257;
  assign n41259 = n41243 & n41258;
  assign n41260 = ~n41212 & ~n41259;
  assign n41261 = n41238 & ~n41260;
  assign n41262 = ~pi0932 & ~n41261;
  assign n41263 = pi0932 & n41238;
  assign n41264 = ~n41260 & n41263;
  assign po0970 = n41262 | n41264;
  assign n41266 = ~n40803 & n40823;
  assign n41267 = ~n40848 & ~n40863;
  assign n41268 = n41266 & ~n41267;
  assign n41269 = ~n40803 & ~n40829;
  assign n41270 = n40848 & n41269;
  assign n41271 = ~n41268 & ~n41270;
  assign n41272 = n40841 & ~n41271;
  assign n41273 = ~n40823 & n40846;
  assign n41274 = ~n40823 & n40829;
  assign n41275 = ~n40880 & ~n41274;
  assign n41276 = n40803 & ~n41275;
  assign n41277 = ~n40823 & ~n40829;
  assign n41278 = ~n40816 & n41277;
  assign n41279 = n40810 & n41278;
  assign n41280 = ~n41276 & ~n41279;
  assign n41281 = ~n41273 & n41280;
  assign n41282 = n40841 & ~n41281;
  assign n41283 = ~n41272 & ~n41282;
  assign n41284 = n40816 & n40830;
  assign n41285 = ~n40810 & n41284;
  assign n41286 = ~n40823 & n40855;
  assign n41287 = ~n41285 & ~n41286;
  assign n41288 = ~n40803 & ~n41287;
  assign n41289 = n40823 & n40871;
  assign n41290 = ~n40823 & n40880;
  assign n41291 = ~n41289 & ~n41290;
  assign n41292 = n40803 & ~n41291;
  assign n41293 = ~n40817 & ~n40880;
  assign n41294 = n40823 & ~n41293;
  assign n41295 = ~n40855 & ~n41294;
  assign n41296 = ~n40803 & ~n41295;
  assign n41297 = n40816 & ~n40823;
  assign n41298 = ~n40803 & n41297;
  assign n41299 = ~n40829 & n41298;
  assign n41300 = ~n40816 & n40829;
  assign n41301 = ~n40855 & ~n41300;
  assign n41302 = ~n40823 & ~n41301;
  assign n41303 = n40803 & n40823;
  assign n41304 = n40845 & n41303;
  assign n41305 = ~n40829 & n41304;
  assign n41306 = ~n41302 & ~n41305;
  assign n41307 = ~n41299 & n41306;
  assign n41308 = ~n41296 & n41307;
  assign n41309 = ~n41285 & n41308;
  assign n41310 = ~n40841 & ~n41309;
  assign n41311 = ~n41292 & ~n41310;
  assign n41312 = ~n41288 & n41311;
  assign n41313 = n41283 & n41312;
  assign n41314 = pi0949 & n41313;
  assign n41315 = ~pi0949 & ~n41313;
  assign po0971 = n41314 | n41315;
  assign n41317 = ~n40563 & ~n40576;
  assign n41318 = ~n40911 & ~n41317;
  assign n41319 = n40557 & ~n41318;
  assign n41320 = n40563 & ~n40569;
  assign n41321 = ~n40584 & n41320;
  assign n41322 = ~n41319 & ~n41321;
  assign n41323 = ~n40557 & n40585;
  assign n41324 = ~n40563 & n41323;
  assign n41325 = ~n40641 & ~n41324;
  assign n41326 = n41322 & n41325;
  assign n41327 = n40551 & ~n41326;
  assign n41328 = ~n40616 & ~n40619;
  assign n41329 = ~n40563 & n40596;
  assign n41330 = n41328 & ~n41329;
  assign n41331 = ~n40557 & ~n41330;
  assign n41332 = n40585 & n40609;
  assign n41333 = ~n40590 & ~n41332;
  assign n41334 = ~n41331 & n41333;
  assign n41335 = ~n40640 & ~n40664;
  assign n41336 = n40557 & ~n41335;
  assign n41337 = n41334 & ~n41336;
  assign n41338 = ~n40551 & ~n41337;
  assign n41339 = ~n41327 & ~n41338;
  assign n41340 = ~n40563 & n40630;
  assign n41341 = n40563 & ~n40661;
  assign n41342 = ~n41340 & ~n41341;
  assign n41343 = n40557 & ~n41342;
  assign n41344 = ~n40616 & n40890;
  assign n41345 = n40621 & ~n41344;
  assign n41346 = ~n41343 & ~n41345;
  assign n41347 = n41339 & n41346;
  assign n41348 = ~pi0938 & ~n41347;
  assign n41349 = pi0938 & n41346;
  assign n41350 = ~n41338 & n41349;
  assign n41351 = ~n41327 & n41350;
  assign po0972 = n41348 | n41351;
  assign n41353 = ~n41235 & ~n41241;
  assign n41354 = ~n41196 & ~n41205;
  assign n41355 = ~n41253 & n41354;
  assign n41356 = n41166 & ~n41355;
  assign n41357 = ~n41172 & ~n41179;
  assign n41358 = ~n41202 & n41357;
  assign n41359 = ~n41185 & n41358;
  assign n41360 = ~n41226 & ~n41359;
  assign n41361 = ~n41166 & n41172;
  assign n41362 = n41247 & n41361;
  assign n41363 = n41360 & ~n41362;
  assign n41364 = ~n41166 & n41250;
  assign n41365 = n41363 & ~n41364;
  assign n41366 = ~n41356 & n41365;
  assign n41367 = n41212 & ~n41366;
  assign n41368 = ~n41166 & n41227;
  assign n41369 = n41172 & n41368;
  assign n41370 = n41185 & n41357;
  assign n41371 = ~n41196 & ~n41370;
  assign n41372 = ~n41166 & ~n41371;
  assign n41373 = ~n41369 & ~n41372;
  assign n41374 = n41166 & n41172;
  assign n41375 = n41244 & n41374;
  assign n41376 = n41166 & n41193;
  assign n41377 = ~n41375 & ~n41376;
  assign n41378 = n41373 & n41377;
  assign n41379 = n41185 & n41203;
  assign n41380 = ~n41194 & ~n41379;
  assign n41381 = ~n41251 & n41380;
  assign n41382 = n41378 & n41381;
  assign n41383 = ~n41212 & ~n41382;
  assign n41384 = ~n41194 & n41360;
  assign n41385 = n41166 & ~n41384;
  assign n41386 = ~n41383 & ~n41385;
  assign n41387 = ~n41367 & n41386;
  assign n41388 = n41353 & n41387;
  assign n41389 = pi0935 & ~n41388;
  assign n41390 = ~pi0935 & n41388;
  assign po0973 = n41389 | n41390;
  assign n41392 = n41179 & n41227;
  assign n41393 = ~n41172 & n41392;
  assign n41394 = ~n41172 & n41244;
  assign n41395 = n41172 & n41228;
  assign n41396 = ~n41394 & ~n41395;
  assign n41397 = n41166 & ~n41396;
  assign n41398 = ~n41393 & ~n41397;
  assign n41399 = ~n41172 & n41368;
  assign n41400 = ~n41242 & ~n41399;
  assign n41401 = n41398 & n41400;
  assign n41402 = ~n41172 & n41213;
  assign n41403 = n41172 & n41250;
  assign n41404 = ~n41402 & ~n41403;
  assign n41405 = n41401 & n41404;
  assign n41406 = n41212 & ~n41405;
  assign n41407 = n41166 & ~n41212;
  assign n41408 = ~n41185 & n41357;
  assign n41409 = ~n41179 & ~n41191;
  assign n41410 = ~n41408 & ~n41409;
  assign n41411 = n41407 & ~n41410;
  assign n41412 = n41166 & n41196;
  assign n41413 = n41172 & n41412;
  assign n41414 = n41172 & n41245;
  assign n41415 = ~n41403 & ~n41414;
  assign n41416 = n41166 & ~n41415;
  assign n41417 = ~n41413 & ~n41416;
  assign n41418 = ~n41205 & ~n41217;
  assign n41419 = n41179 & n41239;
  assign n41420 = ~n41227 & n41419;
  assign n41421 = ~n41214 & ~n41420;
  assign n41422 = n41418 & n41421;
  assign n41423 = ~n41212 & ~n41422;
  assign n41424 = ~n41166 & n41205;
  assign n41425 = ~n41423 & ~n41424;
  assign n41426 = n41417 & n41425;
  assign n41427 = ~n41411 & n41426;
  assign n41428 = ~n41406 & n41427;
  assign n41429 = ~n41362 & n41428;
  assign n41430 = ~pi0934 & ~n41429;
  assign n41431 = pi0934 & ~n41362;
  assign n41432 = n41427 & n41431;
  assign n41433 = ~n41406 & n41432;
  assign po0974 = n41430 | n41433;
  assign n41435 = ~n40947 & n40975;
  assign n41436 = n40934 & n41435;
  assign n41437 = n40934 & n40985;
  assign n41438 = ~n41436 & ~n41437;
  assign n41439 = ~n40934 & n40987;
  assign n41440 = ~n40967 & ~n41439;
  assign n41441 = n40964 & ~n41440;
  assign n41442 = n41438 & ~n41441;
  assign n41443 = ~n40934 & ~n40964;
  assign n41444 = n40941 & n41443;
  assign n41445 = n41442 & ~n41444;
  assign n41446 = n40928 & ~n41445;
  assign n41447 = n40934 & n40941;
  assign n41448 = n40947 & n41447;
  assign n41449 = ~n40953 & n41448;
  assign n41450 = ~n40964 & n41449;
  assign n41451 = ~n40934 & n40964;
  assign n41452 = n41005 & n41451;
  assign n41453 = ~n40965 & ~n41452;
  assign n41454 = ~n40967 & ~n40997;
  assign n41455 = ~n40934 & n40984;
  assign n41456 = n41454 & ~n41455;
  assign n41457 = ~n40964 & ~n41456;
  assign n41458 = n40964 & n40971;
  assign n41459 = n40989 & ~n41458;
  assign n41460 = ~n41457 & n41459;
  assign n41461 = n41453 & n41460;
  assign n41462 = ~n40928 & ~n41461;
  assign n41463 = ~n41450 & ~n41462;
  assign n41464 = ~n41446 & n41463;
  assign n41465 = n40997 & n41451;
  assign n41466 = n40934 & n40999;
  assign n41467 = ~n41465 & ~n41466;
  assign n41468 = n40964 & n41437;
  assign n41469 = n41467 & ~n41468;
  assign n41470 = n41464 & n41469;
  assign n41471 = ~pi0946 & ~n41470;
  assign n41472 = ~n41446 & n41469;
  assign n41473 = n41463 & n41472;
  assign n41474 = pi0946 & n41473;
  assign po0975 = n41471 | n41474;
  assign n41476 = ~n41033 & n41039;
  assign n41477 = ~n41077 & ~n41476;
  assign n41478 = ~n41107 & n41477;
  assign n41479 = ~n41058 & ~n41478;
  assign n41480 = n41052 & n41058;
  assign n41481 = ~n41039 & n41480;
  assign n41482 = ~n41033 & n41052;
  assign n41483 = ~n41045 & n41482;
  assign n41484 = ~n41052 & n41066;
  assign n41485 = ~n41483 & ~n41484;
  assign n41486 = n41033 & n41039;
  assign n41487 = ~n41052 & n41058;
  assign n41488 = n41486 & n41487;
  assign n41489 = n41485 & ~n41488;
  assign n41490 = ~n41481 & n41489;
  assign n41491 = ~n41479 & n41490;
  assign n41492 = n41027 & ~n41491;
  assign n41493 = ~n41033 & n41046;
  assign n41494 = ~n41052 & n41493;
  assign n41495 = ~n41033 & n41093;
  assign n41496 = n41052 & n41495;
  assign n41497 = ~n41494 & ~n41496;
  assign n41498 = ~n41058 & ~n41497;
  assign n41499 = ~n41492 & ~n41498;
  assign n41500 = n41052 & n41066;
  assign n41501 = ~n41081 & ~n41089;
  assign n41502 = ~n41058 & ~n41501;
  assign n41503 = ~n41500 & ~n41502;
  assign n41504 = ~n41085 & n41503;
  assign n41505 = ~n41027 & ~n41504;
  assign n41506 = ~n41063 & ~n41093;
  assign n41507 = n41033 & ~n41506;
  assign n41508 = ~n41094 & ~n41507;
  assign n41509 = n41058 & ~n41508;
  assign n41510 = ~n41027 & n41509;
  assign n41511 = ~n41505 & ~n41510;
  assign n41512 = n41499 & n41511;
  assign n41513 = pi0936 & ~n41512;
  assign n41514 = ~pi0936 & n41499;
  assign n41515 = n41511 & n41514;
  assign po0977 = n41513 | n41515;
  assign n41517 = ~n40816 & n40832;
  assign n41518 = ~n40863 & ~n41517;
  assign n41519 = ~n40803 & ~n41518;
  assign n41520 = n40823 & n40854;
  assign n41521 = ~n41278 & ~n41520;
  assign n41522 = n40803 & ~n41521;
  assign n41523 = ~n40823 & n40849;
  assign n41524 = ~n41299 & ~n41523;
  assign n41525 = ~n40831 & n41524;
  assign n41526 = ~n41522 & n41525;
  assign n41527 = ~n41519 & n41526;
  assign n41528 = ~n41273 & ~n41285;
  assign n41529 = n41527 & n41528;
  assign n41530 = n40841 & ~n41529;
  assign n41531 = n40817 & n41274;
  assign n41532 = n40872 & ~n41531;
  assign n41533 = n40803 & ~n41532;
  assign n41534 = ~n40823 & n40860;
  assign n41535 = ~n41533 & ~n41534;
  assign n41536 = n40810 & n40832;
  assign n41537 = n40823 & n40845;
  assign n41538 = ~n41536 & ~n41537;
  assign n41539 = n40803 & ~n41538;
  assign n41540 = n40803 & n40854;
  assign n41541 = ~n40823 & n41540;
  assign n41542 = ~n41539 & ~n41541;
  assign n41543 = n41535 & n41542;
  assign n41544 = ~n40841 & ~n41543;
  assign n41545 = ~n40849 & ~n40856;
  assign n41546 = ~n41279 & n41545;
  assign n41547 = n40877 & ~n41546;
  assign n41548 = ~n41544 & ~n41547;
  assign n41549 = ~n40831 & ~n41273;
  assign n41550 = ~n40803 & ~n41549;
  assign n41551 = n41548 & ~n41550;
  assign n41552 = ~n41530 & n41551;
  assign n41553 = ~pi0957 & n41552;
  assign n41554 = pi0957 & ~n41552;
  assign po0978 = n41553 | n41554;
  assign n41556 = ~n40953 & n40957;
  assign n41557 = ~n40941 & n41556;
  assign n41558 = ~n40985 & ~n40993;
  assign n41559 = n40934 & n40954;
  assign n41560 = ~n40934 & n41005;
  assign n41561 = ~n41559 & ~n41560;
  assign n41562 = n41558 & n41561;
  assign n41563 = ~n40964 & ~n41562;
  assign n41564 = n40934 & n40966;
  assign n41565 = ~n40965 & ~n41564;
  assign n41566 = ~n40987 & n41565;
  assign n41567 = n40964 & ~n41566;
  assign n41568 = n40934 & n40947;
  assign n41569 = n40953 & n41568;
  assign n41570 = n40941 & n41569;
  assign n41571 = ~n41567 & ~n41570;
  assign n41572 = ~n41563 & n41571;
  assign n41573 = ~n41557 & n41572;
  assign n41574 = ~n40928 & ~n41573;
  assign n41575 = n40934 & ~n40964;
  assign n41576 = n40971 & n41575;
  assign n41577 = ~n40964 & n40987;
  assign n41578 = ~n40964 & n40997;
  assign n41579 = ~n41577 & ~n41578;
  assign n41580 = ~n40934 & ~n41579;
  assign n41581 = ~n41576 & ~n41580;
  assign n41582 = n40934 & n40984;
  assign n41583 = ~n40934 & n40966;
  assign n41584 = ~n41582 & ~n41583;
  assign n41585 = ~n40955 & n41584;
  assign n41586 = ~n40985 & n41585;
  assign n41587 = n40964 & ~n41586;
  assign n41588 = ~n40934 & n40967;
  assign n41589 = ~n41587 & ~n41588;
  assign n41590 = ~n40934 & n40955;
  assign n41591 = ~n41449 & ~n41590;
  assign n41592 = n41589 & n41591;
  assign n41593 = n41581 & n41592;
  assign n41594 = n40928 & ~n41593;
  assign n41595 = ~n40964 & ~n41438;
  assign n41596 = ~n41594 & ~n41595;
  assign n41597 = ~n40988 & ~n41590;
  assign n41598 = n40964 & ~n41597;
  assign n41599 = n41596 & ~n41598;
  assign n41600 = ~n41574 & n41599;
  assign n41601 = pi0955 & ~n41600;
  assign n41602 = ~pi0955 & n41600;
  assign po0979 = n41601 | n41602;
  assign n41604 = ~n41402 & ~n41408;
  assign n41605 = n41212 & ~n41604;
  assign n41606 = n41191 & n41203;
  assign n41607 = ~n41218 & ~n41606;
  assign n41608 = n41166 & ~n41607;
  assign n41609 = n41166 & n41392;
  assign n41610 = ~n41608 & ~n41609;
  assign n41611 = n41212 & ~n41610;
  assign n41612 = ~n41605 & ~n41611;
  assign n41613 = n41213 & n41221;
  assign n41614 = ~n41223 & ~n41613;
  assign n41615 = ~n41217 & ~n41254;
  assign n41616 = ~n41166 & ~n41615;
  assign n41617 = n41212 & n41616;
  assign n41618 = n41614 & ~n41617;
  assign n41619 = ~n41191 & n41203;
  assign n41620 = n41185 & n41619;
  assign n41621 = n41172 & n41192;
  assign n41622 = ~n41197 & ~n41621;
  assign n41623 = ~n41166 & ~n41622;
  assign n41624 = ~n41205 & ~n41226;
  assign n41625 = n41172 & n41195;
  assign n41626 = ~n41247 & ~n41625;
  assign n41627 = n41166 & ~n41626;
  assign n41628 = n41624 & ~n41627;
  assign n41629 = ~n41623 & n41628;
  assign n41630 = ~n41620 & n41629;
  assign n41631 = ~n41212 & ~n41630;
  assign n41632 = ~n41251 & n41360;
  assign n41633 = ~n41166 & ~n41632;
  assign n41634 = ~n41631 & ~n41633;
  assign n41635 = n41618 & n41634;
  assign n41636 = n41612 & n41635;
  assign n41637 = ~pi0948 & ~n41636;
  assign n41638 = pi0948 & n41618;
  assign n41639 = n41612 & n41638;
  assign n41640 = n41634 & n41639;
  assign po0980 = n41637 | n41640;
  assign n41642 = n40477 & n40507;
  assign n41643 = ~n40469 & ~n40477;
  assign n41644 = n40456 & n41643;
  assign n41645 = ~n40504 & ~n41644;
  assign n41646 = n40450 & ~n41645;
  assign n41647 = ~n41642 & ~n41646;
  assign n41648 = ~n40450 & n40477;
  assign n41649 = ~n40469 & n41648;
  assign n41650 = n40463 & n41649;
  assign n41651 = n40485 & n40519;
  assign n41652 = ~n41650 & ~n41651;
  assign n41653 = ~n40450 & n40527;
  assign n41654 = n41652 & ~n41653;
  assign n41655 = ~n40481 & ~n40493;
  assign n41656 = n40469 & n40483;
  assign n41657 = n41655 & ~n41656;
  assign n41658 = n41654 & n41657;
  assign n41659 = n41647 & n41658;
  assign n41660 = n40516 & ~n41659;
  assign n41661 = n40456 & n40479;
  assign n41662 = ~n40504 & ~n41661;
  assign n41663 = ~n40477 & ~n41662;
  assign n41664 = n40463 & n40480;
  assign n41665 = ~n40532 & ~n41664;
  assign n41666 = ~n40456 & ~n40469;
  assign n41667 = ~n40477 & n41666;
  assign n41668 = n41665 & ~n41667;
  assign n41669 = n40450 & ~n41668;
  assign n41670 = n40477 & n40503;
  assign n41671 = n40463 & n40492;
  assign n41672 = ~n41670 & ~n41671;
  assign n41673 = ~n40450 & ~n41672;
  assign n41674 = n40477 & n40486;
  assign n41675 = ~n41673 & ~n41674;
  assign n41676 = ~n41669 & n41675;
  assign n41677 = ~n41663 & n41676;
  assign n41678 = ~n40516 & ~n41677;
  assign n41679 = n40450 & n40522;
  assign n41680 = ~n41678 & ~n41679;
  assign n41681 = n40498 & n41648;
  assign n41682 = ~n40469 & n41681;
  assign n41683 = n41680 & ~n41682;
  assign n41684 = ~n41660 & n41683;
  assign n41685 = ~pi0942 & ~n41684;
  assign n41686 = pi0942 & n41680;
  assign n41687 = ~n41660 & n41686;
  assign n41688 = ~n41682 & n41687;
  assign po0981 = n41685 | n41688;
  assign n41690 = ~n40478 & ~n40484;
  assign n41691 = ~n40450 & ~n41690;
  assign n41692 = ~n40539 & ~n41691;
  assign n41693 = n40456 & ~n40463;
  assign n41694 = n40450 & n41693;
  assign n41695 = ~n40477 & n41694;
  assign n41696 = ~n40456 & n40477;
  assign n41697 = n40463 & n41696;
  assign n41698 = ~n40477 & n40503;
  assign n41699 = ~n41697 & ~n41698;
  assign n41700 = ~n41693 & n41699;
  assign n41701 = n40450 & ~n41700;
  assign n41702 = ~n40487 & ~n41701;
  assign n41703 = ~n40450 & n40470;
  assign n41704 = ~n40477 & n41703;
  assign n41705 = ~n41653 & ~n41704;
  assign n41706 = n41702 & n41705;
  assign n41707 = n40516 & ~n41706;
  assign n41708 = ~n41695 & ~n41707;
  assign n41709 = ~n40504 & ~n40522;
  assign n41710 = ~n40532 & n41709;
  assign n41711 = ~n40450 & ~n41710;
  assign n41712 = n40477 & n40527;
  assign n41713 = ~n40507 & ~n41712;
  assign n41714 = n40450 & ~n41713;
  assign n41715 = ~n41664 & ~n41714;
  assign n41716 = ~n41711 & n41715;
  assign n41717 = ~n40493 & ~n40533;
  assign n41718 = n41716 & n41717;
  assign n41719 = ~n40516 & ~n41718;
  assign n41720 = n41708 & ~n41719;
  assign n41721 = n41692 & n41720;
  assign n41722 = ~pi0952 & ~n41721;
  assign n41723 = pi0952 & n41708;
  assign n41724 = n41692 & n41723;
  assign n41725 = ~n41719 & n41724;
  assign po0982 = n41722 | n41725;
  assign n41727 = ~n40704 & n40760;
  assign n41728 = ~n41142 & ~n41727;
  assign n41729 = ~n40698 & n41728;
  assign n41730 = n40704 & n40735;
  assign n41731 = ~n40724 & ~n40727;
  assign n41732 = n40711 & ~n41731;
  assign n41733 = n40717 & n40754;
  assign n41734 = n40704 & n40727;
  assign n41735 = ~n41733 & ~n41734;
  assign n41736 = ~n41732 & n41735;
  assign n41737 = n40698 & n41736;
  assign n41738 = ~n41730 & n41737;
  assign n41739 = ~n41729 & ~n41738;
  assign n41740 = n40704 & n41732;
  assign n41741 = ~n41140 & ~n41740;
  assign n41742 = ~n41739 & n41741;
  assign n41743 = n40747 & ~n41742;
  assign n41744 = ~n40698 & ~n41731;
  assign n41745 = ~n40704 & n41744;
  assign n41746 = n40704 & n40729;
  assign n41747 = ~n40785 & ~n41746;
  assign n41748 = ~n40698 & ~n41747;
  assign n41749 = ~n40711 & n41744;
  assign n41750 = ~n41748 & ~n41749;
  assign n41751 = ~n41745 & n41750;
  assign n41752 = ~n40747 & ~n41751;
  assign n41753 = ~n41743 & ~n41752;
  assign n41754 = n40698 & ~n41728;
  assign n41755 = ~n40772 & ~n41754;
  assign n41756 = ~n40747 & ~n41755;
  assign n41757 = ~n40698 & n40772;
  assign n41758 = n40698 & ~n41741;
  assign n41759 = ~n41757 & ~n41758;
  assign n41760 = ~n41756 & n41759;
  assign n41761 = n41753 & n41760;
  assign n41762 = pi0950 & ~n41761;
  assign n41763 = ~pi0950 & n41760;
  assign n41764 = ~n41752 & n41763;
  assign n41765 = ~n41743 & n41764;
  assign po0983 = n41762 | n41765;
  assign n41767 = pi3811 & pi9040;
  assign n41768 = pi3820 & ~pi9040;
  assign n41769 = ~n41767 & ~n41768;
  assign n41770 = ~pi0907 & n41769;
  assign n41771 = pi0907 & ~n41769;
  assign n41772 = ~n41770 & ~n41771;
  assign n41773 = pi3855 & pi9040;
  assign n41774 = pi3813 & ~pi9040;
  assign n41775 = ~n41773 & ~n41774;
  assign n41776 = ~pi0909 & n41775;
  assign n41777 = pi0909 & ~n41775;
  assign n41778 = ~n41776 & ~n41777;
  assign n41779 = ~n41772 & ~n41778;
  assign n41780 = pi3820 & pi9040;
  assign n41781 = pi3807 & ~pi9040;
  assign n41782 = ~n41780 & ~n41781;
  assign n41783 = pi0918 & n41782;
  assign n41784 = ~pi0918 & ~n41782;
  assign n41785 = ~n41783 & ~n41784;
  assign n41786 = pi3821 & pi9040;
  assign n41787 = pi3784 & ~pi9040;
  assign n41788 = ~n41786 & ~n41787;
  assign n41789 = pi0914 & n41788;
  assign n41790 = ~pi0914 & ~n41788;
  assign n41791 = ~n41789 & ~n41790;
  assign n41792 = n41778 & ~n41791;
  assign n41793 = n41785 & n41792;
  assign n41794 = ~n41779 & ~n41793;
  assign n41795 = pi3807 & pi9040;
  assign n41796 = pi3791 & ~pi9040;
  assign n41797 = ~n41795 & ~n41796;
  assign n41798 = ~pi0920 & n41797;
  assign n41799 = pi0920 & ~n41797;
  assign n41800 = ~n41798 & ~n41799;
  assign n41801 = pi3828 & pi9040;
  assign n41802 = pi3786 & ~pi9040;
  assign n41803 = ~n41801 & ~n41802;
  assign n41804 = pi0903 & n41803;
  assign n41805 = ~pi0903 & ~n41803;
  assign n41806 = ~n41804 & ~n41805;
  assign n41807 = ~n41800 & ~n41806;
  assign n41808 = ~n41794 & n41807;
  assign n41809 = ~n41778 & n41791;
  assign n41810 = ~n41772 & n41785;
  assign n41811 = ~n41809 & n41810;
  assign n41812 = ~n41800 & n41811;
  assign n41813 = ~n41772 & ~n41785;
  assign n41814 = n41806 & n41813;
  assign n41815 = n41809 & n41814;
  assign n41816 = ~n41772 & ~n41806;
  assign n41817 = n41785 & n41816;
  assign n41818 = ~n41791 & n41817;
  assign n41819 = ~n41815 & ~n41818;
  assign n41820 = ~n41812 & n41819;
  assign n41821 = ~n41772 & n41792;
  assign n41822 = n41778 & n41791;
  assign n41823 = n41772 & n41822;
  assign n41824 = ~n41821 & ~n41823;
  assign n41825 = n41806 & ~n41824;
  assign n41826 = ~n41778 & ~n41791;
  assign n41827 = n41772 & n41806;
  assign n41828 = n41826 & n41827;
  assign n41829 = ~n41785 & n41828;
  assign n41830 = ~n41825 & ~n41829;
  assign n41831 = ~n41800 & ~n41830;
  assign n41832 = n41772 & ~n41785;
  assign n41833 = ~n41792 & ~n41809;
  assign n41834 = n41832 & ~n41833;
  assign n41835 = ~n41778 & ~n41785;
  assign n41836 = ~n41809 & ~n41835;
  assign n41837 = n41772 & ~n41836;
  assign n41838 = n41785 & n41822;
  assign n41839 = ~n41837 & ~n41838;
  assign n41840 = ~n41806 & ~n41839;
  assign n41841 = ~n41834 & ~n41840;
  assign n41842 = ~n41785 & n41822;
  assign n41843 = ~n41772 & n41842;
  assign n41844 = n41772 & n41785;
  assign n41845 = ~n41791 & n41844;
  assign n41846 = ~n41772 & ~n41836;
  assign n41847 = ~n41845 & ~n41846;
  assign n41848 = n41806 & ~n41847;
  assign n41849 = ~n41843 & ~n41848;
  assign n41850 = n41841 & n41849;
  assign n41851 = n41800 & ~n41850;
  assign n41852 = ~n41831 & ~n41851;
  assign n41853 = n41820 & n41852;
  assign n41854 = ~n41808 & n41853;
  assign n41855 = pi0966 & ~n41854;
  assign n41856 = ~pi0966 & n41820;
  assign n41857 = ~n41808 & n41856;
  assign n41858 = n41852 & n41857;
  assign po0984 = n41855 | n41858;
  assign n41860 = n40456 & n40463;
  assign n41861 = ~n40450 & n41860;
  assign n41862 = ~n40477 & n41861;
  assign n41863 = n40477 & n41666;
  assign n41864 = ~n40484 & ~n41863;
  assign n41865 = ~n41671 & n41864;
  assign n41866 = ~n41862 & n41865;
  assign n41867 = n40450 & n41661;
  assign n41868 = n41866 & ~n41867;
  assign n41869 = ~n40516 & ~n41868;
  assign n41870 = ~n40533 & ~n41674;
  assign n41871 = n40450 & ~n41870;
  assign n41872 = n40516 & n40518;
  assign n41873 = ~n40450 & n41872;
  assign n41874 = ~n40463 & n41696;
  assign n41875 = ~n41666 & ~n41874;
  assign n41876 = ~n40486 & n41875;
  assign n41877 = n40450 & ~n41876;
  assign n41878 = n40456 & n40503;
  assign n41879 = n40477 & n41878;
  assign n41880 = ~n41877 & ~n41879;
  assign n41881 = n40516 & ~n41880;
  assign n41882 = ~n41873 & ~n41881;
  assign n41883 = ~n41871 & n41882;
  assign n41884 = ~n40481 & ~n40484;
  assign n41885 = n40477 & n40532;
  assign n41886 = ~n41644 & ~n41885;
  assign n41887 = n41884 & n41886;
  assign n41888 = ~n40450 & ~n41887;
  assign n41889 = n41883 & ~n41888;
  assign n41890 = ~n41869 & n41889;
  assign n41891 = ~pi0940 & ~n41890;
  assign n41892 = pi0940 & n41883;
  assign n41893 = ~n41869 & n41892;
  assign n41894 = ~n41888 & n41893;
  assign po0985 = n41891 | n41894;
  assign n41896 = ~n41052 & n41084;
  assign n41897 = ~n41484 & ~n41896;
  assign n41898 = n41058 & ~n41897;
  assign n41899 = n41081 & n41480;
  assign n41900 = ~n41898 & ~n41899;
  assign n41901 = ~n41105 & n41900;
  assign n41902 = ~n41039 & n41052;
  assign n41903 = n41033 & n41902;
  assign n41904 = n41045 & n41903;
  assign n41905 = ~n41495 & ~n41904;
  assign n41906 = ~n41084 & n41905;
  assign n41907 = n41058 & ~n41906;
  assign n41908 = n41027 & n41907;
  assign n41909 = ~n41058 & n41493;
  assign n41910 = ~n41077 & ~n41103;
  assign n41911 = ~n41068 & n41910;
  assign n41912 = ~n41909 & n41911;
  assign n41913 = n41027 & ~n41912;
  assign n41914 = ~n41033 & ~n41058;
  assign n41915 = n41045 & n41914;
  assign n41916 = n41039 & n41915;
  assign n41917 = n41052 & n41113;
  assign n41918 = ~n41916 & ~n41917;
  assign n41919 = ~n41483 & n41918;
  assign n41920 = n41045 & n41075;
  assign n41921 = n41052 & n41063;
  assign n41922 = ~n41080 & ~n41921;
  assign n41923 = n41058 & ~n41922;
  assign n41924 = ~n41920 & ~n41923;
  assign n41925 = n41919 & n41924;
  assign n41926 = ~n41027 & ~n41925;
  assign n41927 = ~n41052 & n41916;
  assign n41928 = ~n41926 & ~n41927;
  assign n41929 = ~n41913 & n41928;
  assign n41930 = ~n41908 & n41929;
  assign n41931 = n41901 & n41930;
  assign n41932 = pi0939 & ~n41931;
  assign n41933 = ~pi0939 & n41901;
  assign n41934 = n41930 & n41933;
  assign po0986 = n41932 | n41934;
  assign n41936 = ~n41785 & n41826;
  assign n41937 = n41785 & n41809;
  assign n41938 = ~n41936 & ~n41937;
  assign n41939 = n41791 & n41844;
  assign n41940 = n41938 & ~n41939;
  assign n41941 = n41807 & ~n41940;
  assign n41942 = n41793 & ~n41800;
  assign n41943 = ~n41772 & n41942;
  assign n41944 = n41785 & n41826;
  assign n41945 = n41806 & n41944;
  assign n41946 = ~n41785 & n41791;
  assign n41947 = ~n41772 & n41822;
  assign n41948 = ~n41946 & ~n41947;
  assign n41949 = n41806 & ~n41948;
  assign n41950 = ~n41945 & ~n41949;
  assign n41951 = ~n41800 & ~n41950;
  assign n41952 = ~n41943 & ~n41951;
  assign n41953 = n41791 & n41813;
  assign n41954 = ~n41791 & n41832;
  assign n41955 = n41778 & n41954;
  assign n41956 = ~n41953 & ~n41955;
  assign n41957 = n41806 & ~n41956;
  assign n41958 = n41952 & ~n41957;
  assign n41959 = n41816 & n41822;
  assign n41960 = n41785 & n41959;
  assign n41961 = ~n41833 & n41844;
  assign n41962 = n41772 & n41936;
  assign n41963 = ~n41961 & ~n41962;
  assign n41964 = n41772 & ~n41806;
  assign n41965 = n41842 & n41964;
  assign n41966 = n41813 & ~n41833;
  assign n41967 = ~n41772 & n41944;
  assign n41968 = ~n41966 & ~n41967;
  assign n41969 = ~n41965 & n41968;
  assign n41970 = n41963 & n41969;
  assign n41971 = ~n41960 & n41970;
  assign n41972 = n41785 & n41827;
  assign n41973 = n41778 & n41972;
  assign n41974 = n41971 & ~n41973;
  assign n41975 = n41800 & ~n41974;
  assign n41976 = n41958 & ~n41975;
  assign n41977 = ~n41941 & n41976;
  assign n41978 = ~pi0959 & ~n41977;
  assign n41979 = pi0959 & n41958;
  assign n41980 = ~n41941 & n41979;
  assign n41981 = ~n41975 & n41980;
  assign po0987 = n41978 | n41981;
  assign n41983 = ~n41785 & n41809;
  assign n41984 = ~n41838 & ~n41983;
  assign n41985 = n41806 & ~n41984;
  assign n41986 = n41772 & n41792;
  assign n41987 = ~n41937 & ~n41986;
  assign n41988 = ~n41842 & n41987;
  assign n41989 = ~n41806 & ~n41988;
  assign n41990 = ~n41985 & ~n41989;
  assign n41991 = ~n41945 & ~n41955;
  assign n41992 = n41990 & n41991;
  assign n41993 = n41800 & ~n41992;
  assign n41994 = n41785 & n41806;
  assign n41995 = ~n41791 & n41994;
  assign n41996 = n41778 & n41995;
  assign n41997 = n41938 & ~n41996;
  assign n41998 = ~n41842 & n41997;
  assign n41999 = n41772 & ~n41998;
  assign n42000 = ~n41772 & n41838;
  assign n42001 = n41772 & n41826;
  assign n42002 = ~n41821 & ~n42001;
  assign n42003 = ~n41806 & ~n42002;
  assign n42004 = ~n42000 & ~n42003;
  assign n42005 = ~n41999 & n42004;
  assign n42006 = ~n41800 & ~n42005;
  assign n42007 = ~n41993 & ~n42006;
  assign n42008 = ~n41785 & n41821;
  assign n42009 = ~n41967 & ~n42008;
  assign n42010 = n41806 & ~n42009;
  assign n42011 = n41816 & n41835;
  assign n42012 = ~n42010 & ~n42011;
  assign n42013 = n42007 & n42012;
  assign n42014 = ~pi0951 & ~n42013;
  assign n42015 = pi0951 & ~n42010;
  assign n42016 = n42007 & n42015;
  assign n42017 = ~n42011 & n42016;
  assign po0988 = n42014 | n42017;
  assign n42019 = n41806 & n41838;
  assign n42020 = n41772 & n42019;
  assign n42021 = ~n41829 & ~n42020;
  assign n42022 = ~n41962 & ~n41965;
  assign n42023 = n41779 & n41785;
  assign n42024 = ~n41947 & ~n42023;
  assign n42025 = n41806 & ~n42024;
  assign n42026 = ~n41806 & ~n41832;
  assign n42027 = ~n41833 & n42026;
  assign n42028 = ~n41785 & ~n41822;
  assign n42029 = n41806 & n42028;
  assign n42030 = n41772 & n42029;
  assign n42031 = ~n42027 & ~n42030;
  assign n42032 = ~n42025 & n42031;
  assign n42033 = n42022 & n42032;
  assign n42034 = ~n41800 & ~n42033;
  assign n42035 = n42021 & ~n42034;
  assign n42036 = ~n41806 & n41937;
  assign n42037 = ~n41772 & n42036;
  assign n42038 = n41800 & ~n41806;
  assign n42039 = ~n41834 & ~n41947;
  assign n42040 = ~n41944 & n42039;
  assign n42041 = n42038 & ~n42040;
  assign n42042 = ~n41772 & n41936;
  assign n42043 = n41779 & ~n41785;
  assign n42044 = ~n41821 & ~n42043;
  assign n42045 = ~n41793 & ~n41823;
  assign n42046 = n42044 & n42045;
  assign n42047 = n41806 & ~n42046;
  assign n42048 = ~n42042 & ~n42047;
  assign n42049 = n41800 & ~n42048;
  assign n42050 = ~n42041 & ~n42049;
  assign n42051 = ~n42037 & n42050;
  assign n42052 = n42035 & n42051;
  assign n42053 = pi0965 & ~n42052;
  assign n42054 = ~pi0965 & n42035;
  assign n42055 = n42051 & n42054;
  assign po0989 = n42053 | n42055;
  assign n42057 = ~n41439 & ~n41590;
  assign n42058 = ~n41570 & n42057;
  assign n42059 = ~n40964 & ~n42058;
  assign n42060 = ~n41452 & ~n41468;
  assign n42061 = ~n41449 & ~n41578;
  assign n42062 = ~n41435 & ~n41583;
  assign n42063 = n40964 & ~n42062;
  assign n42064 = ~n40993 & ~n42063;
  assign n42065 = n42061 & n42064;
  assign n42066 = n40928 & ~n42065;
  assign n42067 = n40947 & n40953;
  assign n42068 = ~n40972 & ~n42067;
  assign n42069 = n40934 & ~n42068;
  assign n42070 = ~n40955 & ~n41455;
  assign n42071 = n40964 & ~n42070;
  assign n42072 = n40934 & n40953;
  assign n42073 = ~n40967 & ~n42072;
  assign n42074 = ~n40975 & n42073;
  assign n42075 = ~n40964 & ~n42074;
  assign n42076 = ~n42071 & ~n42075;
  assign n42077 = ~n42069 & n42076;
  assign n42078 = ~n40928 & ~n42077;
  assign n42079 = ~n42066 & ~n42078;
  assign n42080 = n42060 & n42079;
  assign n42081 = ~n42059 & n42080;
  assign n42082 = ~pi0960 & ~n42081;
  assign n42083 = pi0960 & n42060;
  assign n42084 = ~n42059 & n42083;
  assign n42085 = n42079 & n42084;
  assign po0990 = n42082 | n42085;
  assign n42087 = n41052 & ~n41506;
  assign n42088 = n41033 & n42087;
  assign n42089 = n41045 & n41482;
  assign n42090 = ~n41115 & ~n42089;
  assign n42091 = ~n41495 & n42090;
  assign n42092 = ~n41058 & ~n42091;
  assign n42093 = ~n41088 & ~n41493;
  assign n42094 = n41058 & ~n42093;
  assign n42095 = ~n42092 & ~n42094;
  assign n42096 = ~n42088 & n42095;
  assign n42097 = ~n41052 & n41081;
  assign n42098 = n42096 & ~n42097;
  assign n42099 = ~n41027 & ~n42098;
  assign n42100 = ~n41084 & ~n41089;
  assign n42101 = ~n41081 & ~n41495;
  assign n42102 = n42100 & n42101;
  assign n42103 = n41052 & ~n42102;
  assign n42104 = n41062 & ~n42093;
  assign n42105 = ~n42103 & ~n42104;
  assign n42106 = ~n41484 & n42105;
  assign n42107 = n41027 & ~n42106;
  assign n42108 = ~n42099 & ~n42107;
  assign n42109 = n41052 & n41493;
  assign n42110 = ~n42097 & ~n42109;
  assign n42111 = n41058 & ~n42110;
  assign n42112 = n42108 & ~n42111;
  assign n42113 = pi0929 & ~n42112;
  assign n42114 = ~pi0929 & ~n42111;
  assign n42115 = ~n42107 & n42114;
  assign n42116 = ~n42099 & n42115;
  assign po0991 = n42113 | n42116;
  assign n42118 = ~n40803 & n40860;
  assign n42119 = ~n40823 & n40845;
  assign n42120 = ~n40844 & ~n42119;
  assign n42121 = ~n40803 & ~n42120;
  assign n42122 = n40803 & ~n41301;
  assign n42123 = ~n42121 & ~n42122;
  assign n42124 = ~n41289 & n42123;
  assign n42125 = n40841 & ~n42124;
  assign n42126 = ~n42118 & ~n42125;
  assign n42127 = n40829 & n41266;
  assign n42128 = ~n41277 & ~n42127;
  assign n42129 = ~n40810 & ~n42128;
  assign n42130 = ~n40831 & ~n42129;
  assign n42131 = ~n41278 & n42130;
  assign n42132 = n40823 & n40863;
  assign n42133 = n40803 & n40846;
  assign n42134 = ~n42132 & ~n42133;
  assign n42135 = n42131 & n42134;
  assign n42136 = ~n40841 & ~n42135;
  assign n42137 = ~n41523 & ~n41537;
  assign n42138 = n40803 & ~n42137;
  assign n42139 = ~n42136 & ~n42138;
  assign n42140 = n42126 & n42139;
  assign n42141 = ~pi0980 & ~n42140;
  assign n42142 = ~n42125 & n42139;
  assign n42143 = pi0980 & n42142;
  assign n42144 = ~n42118 & n42143;
  assign po0992 = n42141 | n42144;
  assign n42146 = ~n40698 & n40726;
  assign n42147 = n40754 & ~n41731;
  assign n42148 = ~n40730 & ~n42147;
  assign n42149 = ~n41140 & n42148;
  assign n42150 = n40698 & ~n42149;
  assign n42151 = n40704 & n40770;
  assign n42152 = ~n42150 & ~n42151;
  assign n42153 = ~n40711 & n40729;
  assign n42154 = ~n40704 & n41144;
  assign n42155 = ~n42153 & ~n42154;
  assign n42156 = ~n41734 & n42155;
  assign n42157 = ~n40698 & ~n42156;
  assign n42158 = n42152 & ~n42157;
  assign n42159 = n40747 & ~n42158;
  assign n42160 = ~n42146 & ~n42159;
  assign n42161 = ~n40704 & n40727;
  assign n42162 = ~n41139 & ~n42161;
  assign n42163 = ~n40698 & ~n42162;
  assign n42164 = ~n40731 & ~n42163;
  assign n42165 = ~n40726 & ~n40785;
  assign n42166 = n40704 & n40789;
  assign n42167 = ~n41144 & ~n42166;
  assign n42168 = ~n42153 & n42167;
  assign n42169 = n40698 & ~n42168;
  assign n42170 = ~n40704 & n40770;
  assign n42171 = ~n42169 & ~n42170;
  assign n42172 = n42165 & n42171;
  assign n42173 = n42164 & n42172;
  assign n42174 = ~n40747 & ~n42173;
  assign n42175 = ~n40762 & ~n41730;
  assign n42176 = n40698 & ~n42175;
  assign n42177 = ~n42174 & ~n42176;
  assign n42178 = n42160 & n42177;
  assign n42179 = pi0944 & n42178;
  assign n42180 = ~pi0944 & ~n42178;
  assign po0993 = n42179 | n42180;
  assign n42182 = pi3942 & pi9040;
  assign n42183 = pi3891 & ~pi9040;
  assign n42184 = ~n42182 & ~n42183;
  assign n42185 = pi0954 & n42184;
  assign n42186 = ~pi0954 & ~n42184;
  assign n42187 = ~n42185 & ~n42186;
  assign n42188 = pi3927 & pi9040;
  assign n42189 = pi3884 & ~pi9040;
  assign n42190 = ~n42188 & ~n42189;
  assign n42191 = ~pi0973 & ~n42190;
  assign n42192 = pi0973 & ~n42188;
  assign n42193 = ~n42189 & n42192;
  assign n42194 = ~n42191 & ~n42193;
  assign n42195 = pi3882 & pi9040;
  assign n42196 = pi3944 & ~pi9040;
  assign n42197 = ~n42195 & ~n42196;
  assign n42198 = ~pi0975 & ~n42197;
  assign n42199 = pi0975 & ~n42195;
  assign n42200 = ~n42196 & n42199;
  assign n42201 = ~n42198 & ~n42200;
  assign n42202 = pi3883 & pi9040;
  assign n42203 = pi3896 & ~pi9040;
  assign n42204 = ~n42202 & ~n42203;
  assign n42205 = ~pi0972 & n42204;
  assign n42206 = pi0972 & ~n42204;
  assign n42207 = ~n42205 & ~n42206;
  assign n42208 = n42201 & ~n42207;
  assign n42209 = ~n42194 & n42208;
  assign n42210 = pi3910 & pi9040;
  assign n42211 = pi3916 & ~pi9040;
  assign n42212 = ~n42210 & ~n42211;
  assign n42213 = pi0990 & n42212;
  assign n42214 = ~pi0990 & ~n42212;
  assign n42215 = ~n42213 & ~n42214;
  assign n42216 = n42209 & ~n42215;
  assign n42217 = ~n42201 & n42207;
  assign n42218 = ~n42215 & n42217;
  assign n42219 = ~n42194 & n42218;
  assign n42220 = ~n42216 & ~n42219;
  assign n42221 = n42194 & n42215;
  assign n42222 = n42217 & n42221;
  assign n42223 = n42201 & n42207;
  assign n42224 = ~n42194 & n42223;
  assign n42225 = n42215 & n42224;
  assign n42226 = ~n42222 & ~n42225;
  assign n42227 = n42220 & n42226;
  assign n42228 = n42187 & ~n42227;
  assign n42229 = ~n42194 & n42215;
  assign n42230 = ~n42207 & n42229;
  assign n42231 = ~n42201 & n42230;
  assign n42232 = ~n42224 & ~n42231;
  assign n42233 = n42187 & ~n42232;
  assign n42234 = ~n42207 & ~n42215;
  assign n42235 = ~n42187 & n42234;
  assign n42236 = n42194 & n42201;
  assign n42237 = n42215 & n42217;
  assign n42238 = ~n42236 & ~n42237;
  assign n42239 = ~n42187 & ~n42238;
  assign n42240 = ~n42235 & ~n42239;
  assign n42241 = ~n42201 & ~n42207;
  assign n42242 = n42194 & n42241;
  assign n42243 = ~n42215 & n42242;
  assign n42244 = n42240 & ~n42243;
  assign n42245 = ~n42207 & n42236;
  assign n42246 = n42215 & n42245;
  assign n42247 = n42244 & ~n42246;
  assign n42248 = ~n42233 & n42247;
  assign n42249 = pi3882 & ~pi9040;
  assign n42250 = pi3885 & pi9040;
  assign n42251 = ~n42249 & ~n42250;
  assign n42252 = ~pi0985 & ~n42251;
  assign n42253 = pi0985 & n42251;
  assign n42254 = ~n42252 & ~n42253;
  assign n42255 = ~n42248 & ~n42254;
  assign n42256 = ~n42194 & ~n42207;
  assign n42257 = ~n42187 & n42215;
  assign n42258 = n42254 & n42257;
  assign n42259 = n42256 & n42258;
  assign n42260 = ~n42194 & ~n42215;
  assign n42261 = n42207 & n42260;
  assign n42262 = ~n42187 & ~n42261;
  assign n42263 = ~n42201 & n42221;
  assign n42264 = ~n42208 & ~n42256;
  assign n42265 = ~n42215 & ~n42264;
  assign n42266 = n42194 & n42217;
  assign n42267 = ~n42265 & ~n42266;
  assign n42268 = n42187 & n42267;
  assign n42269 = ~n42263 & n42268;
  assign n42270 = ~n42262 & ~n42269;
  assign n42271 = n42194 & n42223;
  assign n42272 = n42215 & n42271;
  assign n42273 = ~n42270 & ~n42272;
  assign n42274 = n42254 & ~n42273;
  assign n42275 = ~n42259 & ~n42274;
  assign n42276 = ~n42255 & n42275;
  assign n42277 = ~n42228 & n42276;
  assign n42278 = ~n42187 & n42243;
  assign n42279 = n42277 & ~n42278;
  assign n42280 = pi1059 & ~n42279;
  assign n42281 = n42276 & ~n42278;
  assign n42282 = ~pi1059 & n42281;
  assign n42283 = ~n42228 & n42282;
  assign po1020 = n42280 | n42283;
  assign n42285 = pi3908 & pi9040;
  assign n42286 = pi3888 & ~pi9040;
  assign n42287 = ~n42285 & ~n42286;
  assign n42288 = pi0978 & n42287;
  assign n42289 = ~pi0978 & ~n42287;
  assign n42290 = ~n42288 & ~n42289;
  assign n42291 = pi3913 & pi9040;
  assign n42292 = pi3908 & ~pi9040;
  assign n42293 = ~n42291 & ~n42292;
  assign n42294 = pi0977 & n42293;
  assign n42295 = ~pi0977 & ~n42293;
  assign n42296 = ~n42294 & ~n42295;
  assign n42297 = pi3877 & pi9040;
  assign n42298 = pi3906 & ~pi9040;
  assign n42299 = ~n42297 & ~n42298;
  assign n42300 = pi0967 & n42299;
  assign n42301 = ~pi0967 & ~n42299;
  assign n42302 = ~n42300 & ~n42301;
  assign n42303 = n42296 & ~n42302;
  assign n42304 = pi3878 & pi9040;
  assign n42305 = pi3872 & ~pi9040;
  assign n42306 = ~n42304 & ~n42305;
  assign n42307 = ~pi0986 & n42306;
  assign n42308 = pi0986 & ~n42306;
  assign n42309 = ~n42307 & ~n42308;
  assign n42310 = pi3909 & pi9040;
  assign n42311 = pi3913 & ~pi9040;
  assign n42312 = ~n42310 & ~n42311;
  assign n42313 = pi0945 & n42312;
  assign n42314 = ~pi0945 & ~n42312;
  assign n42315 = ~n42313 & ~n42314;
  assign n42316 = ~n42309 & n42315;
  assign n42317 = n42303 & n42316;
  assign n42318 = ~n42309 & ~n42315;
  assign n42319 = ~n42296 & n42318;
  assign n42320 = ~n42317 & ~n42319;
  assign n42321 = ~n42290 & ~n42320;
  assign n42322 = pi3898 & pi9040;
  assign n42323 = pi3924 & ~pi9040;
  assign n42324 = ~n42322 & ~n42323;
  assign n42325 = ~pi0979 & ~n42324;
  assign n42326 = pi0979 & n42324;
  assign n42327 = ~n42325 & ~n42326;
  assign n42328 = n42290 & n42309;
  assign n42329 = n42296 & n42328;
  assign n42330 = n42303 & ~n42315;
  assign n42331 = n42296 & n42302;
  assign n42332 = n42315 & n42331;
  assign n42333 = ~n42330 & ~n42332;
  assign n42334 = ~n42296 & ~n42302;
  assign n42335 = n42315 & n42334;
  assign n42336 = ~n42309 & n42335;
  assign n42337 = n42333 & ~n42336;
  assign n42338 = n42290 & ~n42337;
  assign n42339 = ~n42329 & ~n42338;
  assign n42340 = ~n42296 & n42302;
  assign n42341 = ~n42315 & n42340;
  assign n42342 = ~n42309 & n42341;
  assign n42343 = n42339 & ~n42342;
  assign n42344 = n42309 & n42334;
  assign n42345 = ~n42296 & n42315;
  assign n42346 = n42302 & n42345;
  assign n42347 = ~n42344 & ~n42346;
  assign n42348 = ~n42290 & ~n42347;
  assign n42349 = ~n42315 & n42331;
  assign n42350 = n42309 & n42349;
  assign n42351 = ~n42348 & ~n42350;
  assign n42352 = n42343 & n42351;
  assign n42353 = n42327 & ~n42352;
  assign n42354 = ~n42321 & ~n42353;
  assign n42355 = n42290 & ~n42327;
  assign n42356 = ~n42347 & n42355;
  assign n42357 = ~n42315 & n42334;
  assign n42358 = ~n42349 & ~n42357;
  assign n42359 = ~n42309 & ~n42358;
  assign n42360 = ~n42317 & ~n42359;
  assign n42361 = ~n42327 & ~n42360;
  assign n42362 = ~n42356 & ~n42361;
  assign n42363 = ~n42290 & ~n42327;
  assign n42364 = n42303 & n42309;
  assign n42365 = ~n42341 & ~n42364;
  assign n42366 = n42296 & n42315;
  assign n42367 = n42365 & ~n42366;
  assign n42368 = n42363 & ~n42367;
  assign n42369 = n42362 & ~n42368;
  assign n42370 = n42354 & n42369;
  assign n42371 = ~pi1061 & ~n42370;
  assign n42372 = pi1061 & n42362;
  assign n42373 = n42354 & n42372;
  assign n42374 = ~n42368 & n42373;
  assign po1021 = n42371 | n42374;
  assign n42376 = pi3920 & pi9040;
  assign n42377 = pi3894 & ~pi9040;
  assign n42378 = ~n42376 & ~n42377;
  assign n42379 = ~pi0977 & ~n42378;
  assign n42380 = pi0977 & n42378;
  assign n42381 = ~n42379 & ~n42380;
  assign n42382 = pi3922 & pi9040;
  assign n42383 = pi3907 & ~pi9040;
  assign n42384 = ~n42382 & ~n42383;
  assign n42385 = ~pi0975 & n42384;
  assign n42386 = pi0975 & ~n42384;
  assign n42387 = ~n42385 & ~n42386;
  assign n42388 = pi3900 & pi9040;
  assign n42389 = pi3922 & ~pi9040;
  assign n42390 = ~n42388 & ~n42389;
  assign n42391 = ~pi0985 & ~n42390;
  assign n42392 = pi0985 & ~n42388;
  assign n42393 = ~n42389 & n42392;
  assign n42394 = ~n42391 & ~n42393;
  assign n42395 = pi3928 & pi9040;
  assign n42396 = pi3874 & ~pi9040;
  assign n42397 = ~n42395 & ~n42396;
  assign n42398 = ~pi0945 & n42397;
  assign n42399 = pi0945 & ~n42397;
  assign n42400 = ~n42398 & ~n42399;
  assign n42401 = ~n42394 & ~n42400;
  assign n42402 = pi3899 & pi9040;
  assign n42403 = pi3900 & ~pi9040;
  assign n42404 = ~n42402 & ~n42403;
  assign n42405 = pi0976 & n42404;
  assign n42406 = ~pi0976 & ~n42404;
  assign n42407 = ~n42405 & ~n42406;
  assign n42408 = pi3924 & pi9040;
  assign n42409 = pi3893 & ~pi9040;
  assign n42410 = ~n42408 & ~n42409;
  assign n42411 = ~pi0987 & n42410;
  assign n42412 = pi0987 & ~n42410;
  assign n42413 = ~n42411 & ~n42412;
  assign n42414 = n42407 & ~n42413;
  assign n42415 = n42401 & n42414;
  assign n42416 = ~n42387 & n42415;
  assign n42417 = ~n42407 & ~n42413;
  assign n42418 = n42394 & ~n42400;
  assign n42419 = n42417 & n42418;
  assign n42420 = ~n42394 & n42400;
  assign n42421 = ~n42387 & n42420;
  assign n42422 = ~n42407 & n42421;
  assign n42423 = n42394 & n42400;
  assign n42424 = ~n42387 & n42423;
  assign n42425 = ~n42413 & n42424;
  assign n42426 = n42407 & n42425;
  assign n42427 = ~n42422 & ~n42426;
  assign n42428 = ~n42419 & n42427;
  assign n42429 = ~n42416 & n42428;
  assign n42430 = n42387 & ~n42407;
  assign n42431 = ~n42400 & n42430;
  assign n42432 = n42394 & n42431;
  assign n42433 = n42429 & ~n42432;
  assign n42434 = ~n42381 & ~n42433;
  assign n42435 = ~n42387 & n42394;
  assign n42436 = ~n42400 & n42435;
  assign n42437 = n42407 & n42436;
  assign n42438 = ~n42387 & ~n42407;
  assign n42439 = n42400 & n42438;
  assign n42440 = ~n42437 & ~n42439;
  assign n42441 = n42387 & n42401;
  assign n42442 = n42407 & n42441;
  assign n42443 = n42440 & ~n42442;
  assign n42444 = n42413 & ~n42443;
  assign n42445 = n42387 & n42400;
  assign n42446 = n42394 & n42445;
  assign n42447 = n42413 & n42446;
  assign n42448 = n42407 & n42447;
  assign n42449 = ~n42394 & n42438;
  assign n42450 = ~n42407 & n42420;
  assign n42451 = ~n42449 & ~n42450;
  assign n42452 = n42413 & ~n42451;
  assign n42453 = ~n42448 & ~n42452;
  assign n42454 = ~n42381 & ~n42453;
  assign n42455 = ~n42444 & ~n42454;
  assign n42456 = ~n42434 & n42455;
  assign n42457 = n42387 & n42407;
  assign n42458 = ~n42413 & n42457;
  assign n42459 = n42420 & n42458;
  assign n42460 = n42387 & n42394;
  assign n42461 = n42417 & n42460;
  assign n42462 = n42413 & n42435;
  assign n42463 = ~n42394 & n42407;
  assign n42464 = n42387 & n42463;
  assign n42465 = ~n42441 & ~n42464;
  assign n42466 = ~n42462 & n42465;
  assign n42467 = ~n42407 & n42446;
  assign n42468 = n42466 & ~n42467;
  assign n42469 = n42387 & ~n42400;
  assign n42470 = n42407 & n42420;
  assign n42471 = ~n42469 & ~n42470;
  assign n42472 = ~n42413 & ~n42471;
  assign n42473 = n42401 & ~n42413;
  assign n42474 = ~n42407 & n42473;
  assign n42475 = ~n42472 & ~n42474;
  assign n42476 = n42468 & n42475;
  assign n42477 = n42381 & ~n42476;
  assign n42478 = ~n42461 & ~n42477;
  assign n42479 = ~n42459 & n42478;
  assign n42480 = n42456 & n42479;
  assign n42481 = pi1071 & n42480;
  assign n42482 = ~pi1071 & ~n42480;
  assign po1023 = n42481 | n42482;
  assign n42484 = pi3884 & pi9040;
  assign n42485 = pi3897 & ~pi9040;
  assign n42486 = ~n42484 & ~n42485;
  assign n42487 = ~pi0964 & n42486;
  assign n42488 = pi0964 & ~n42486;
  assign n42489 = ~n42487 & ~n42488;
  assign n42490 = pi3889 & pi9040;
  assign n42491 = pi3942 & ~pi9040;
  assign n42492 = ~n42490 & ~n42491;
  assign n42493 = ~pi0989 & n42492;
  assign n42494 = pi0989 & ~n42492;
  assign n42495 = ~n42493 & ~n42494;
  assign n42496 = n42489 & n42495;
  assign n42497 = pi3926 & pi9040;
  assign n42498 = pi3871 & ~pi9040;
  assign n42499 = ~n42497 & ~n42498;
  assign n42500 = pi0953 & n42499;
  assign n42501 = ~pi0953 & ~n42499;
  assign n42502 = ~n42500 & ~n42501;
  assign n42503 = pi3918 & pi9040;
  assign n42504 = pi3919 & ~pi9040;
  assign n42505 = ~n42503 & ~n42504;
  assign n42506 = ~pi0971 & n42505;
  assign n42507 = pi0971 & ~n42505;
  assign n42508 = ~n42506 & ~n42507;
  assign n42509 = pi3911 & pi9040;
  assign n42510 = pi3889 & ~pi9040;
  assign n42511 = ~n42509 & ~n42510;
  assign n42512 = ~pi0961 & ~n42511;
  assign n42513 = pi0961 & n42511;
  assign n42514 = ~n42512 & ~n42513;
  assign n42515 = ~n42508 & ~n42514;
  assign n42516 = ~n42502 & n42515;
  assign n42517 = pi3897 & pi9040;
  assign n42518 = pi3926 & ~pi9040;
  assign n42519 = ~n42517 & ~n42518;
  assign n42520 = ~pi0983 & ~n42519;
  assign n42521 = pi0983 & n42519;
  assign n42522 = ~n42520 & ~n42521;
  assign n42523 = n42514 & ~n42522;
  assign n42524 = ~n42508 & n42523;
  assign n42525 = n42502 & n42524;
  assign n42526 = n42514 & n42522;
  assign n42527 = ~n42502 & n42526;
  assign n42528 = ~n42525 & ~n42527;
  assign n42529 = ~n42516 & n42528;
  assign n42530 = n42496 & ~n42529;
  assign n42531 = ~n42502 & n42508;
  assign n42532 = ~n42522 & n42531;
  assign n42533 = ~n42514 & ~n42522;
  assign n42534 = ~n42508 & n42533;
  assign n42535 = n42502 & n42534;
  assign n42536 = ~n42532 & ~n42535;
  assign n42537 = n42508 & n42523;
  assign n42538 = ~n42508 & n42526;
  assign n42539 = ~n42537 & ~n42538;
  assign n42540 = n42536 & n42539;
  assign n42541 = ~n42489 & ~n42540;
  assign n42542 = ~n42514 & n42522;
  assign n42543 = n42508 & n42542;
  assign n42544 = n42502 & n42543;
  assign n42545 = ~n42541 & ~n42544;
  assign n42546 = n42495 & ~n42545;
  assign n42547 = ~n42530 & ~n42546;
  assign n42548 = ~n42526 & ~n42533;
  assign n42549 = n42502 & ~n42548;
  assign n42550 = n42508 & n42533;
  assign n42551 = ~n42549 & ~n42550;
  assign n42552 = n42489 & ~n42551;
  assign n42553 = ~n42508 & n42542;
  assign n42554 = ~n42516 & ~n42553;
  assign n42555 = ~n42525 & n42554;
  assign n42556 = ~n42489 & ~n42555;
  assign n42557 = ~n42552 & ~n42556;
  assign n42558 = n42489 & ~n42502;
  assign n42559 = n42523 & n42558;
  assign n42560 = n42502 & n42508;
  assign n42561 = ~n42522 & n42560;
  assign n42562 = ~n42514 & n42561;
  assign n42563 = n42508 & n42514;
  assign n42564 = n42522 & n42563;
  assign n42565 = n42502 & n42564;
  assign n42566 = ~n42562 & ~n42565;
  assign n42567 = n42522 & n42531;
  assign n42568 = ~n42514 & n42567;
  assign n42569 = n42566 & ~n42568;
  assign n42570 = ~n42559 & n42569;
  assign n42571 = n42557 & n42570;
  assign n42572 = ~n42495 & ~n42571;
  assign n42573 = ~n42489 & ~n42502;
  assign n42574 = ~n42508 & n42573;
  assign n42575 = n42522 & n42574;
  assign n42576 = ~n42502 & n42537;
  assign n42577 = ~n42575 & ~n42576;
  assign n42578 = ~n42572 & n42577;
  assign n42579 = n42547 & n42578;
  assign n42580 = pi1060 & ~n42579;
  assign n42581 = ~pi1060 & n42577;
  assign n42582 = n42547 & n42581;
  assign n42583 = ~n42572 & n42582;
  assign po1025 = n42580 | n42583;
  assign n42585 = ~n42387 & ~n42394;
  assign n42586 = ~n42432 & ~n42585;
  assign n42587 = ~n42463 & n42586;
  assign n42588 = ~n42413 & ~n42587;
  assign n42589 = n42407 & n42413;
  assign n42590 = n42394 & n42589;
  assign n42591 = ~n42387 & n42407;
  assign n42592 = ~n42400 & n42591;
  assign n42593 = ~n42407 & n42424;
  assign n42594 = ~n42592 & ~n42593;
  assign n42595 = n42387 & ~n42394;
  assign n42596 = ~n42407 & n42413;
  assign n42597 = n42595 & n42596;
  assign n42598 = n42594 & ~n42597;
  assign n42599 = ~n42590 & n42598;
  assign n42600 = ~n42588 & n42599;
  assign n42601 = n42381 & ~n42600;
  assign n42602 = ~n42387 & n42401;
  assign n42603 = ~n42407 & n42602;
  assign n42604 = n42407 & n42421;
  assign n42605 = ~n42603 & ~n42604;
  assign n42606 = ~n42413 & ~n42605;
  assign n42607 = ~n42601 & ~n42606;
  assign n42608 = n42407 & n42424;
  assign n42609 = ~n42436 & ~n42446;
  assign n42610 = ~n42413 & ~n42609;
  assign n42611 = ~n42608 & ~n42610;
  assign n42612 = ~n42442 & n42611;
  assign n42613 = ~n42381 & ~n42612;
  assign n42614 = ~n42418 & ~n42420;
  assign n42615 = n42387 & ~n42614;
  assign n42616 = ~n42450 & ~n42615;
  assign n42617 = n42413 & ~n42616;
  assign n42618 = ~n42381 & n42617;
  assign n42619 = ~n42613 & ~n42618;
  assign n42620 = n42607 & n42619;
  assign n42621 = pi1066 & ~n42620;
  assign n42622 = ~pi1066 & n42607;
  assign n42623 = n42619 & n42622;
  assign po1026 = n42621 | n42623;
  assign n42625 = ~n42550 & ~n42553;
  assign n42626 = n42489 & ~n42625;
  assign n42627 = n42502 & n42538;
  assign n42628 = ~n42626 & ~n42627;
  assign n42629 = n42502 & n42514;
  assign n42630 = ~n42563 & ~n42629;
  assign n42631 = ~n42534 & n42630;
  assign n42632 = ~n42489 & ~n42631;
  assign n42633 = n42628 & ~n42632;
  assign n42634 = n42495 & ~n42633;
  assign n42635 = ~n42502 & n42564;
  assign n42636 = n42489 & n42635;
  assign n42637 = ~n42508 & n42559;
  assign n42638 = ~n42636 & ~n42637;
  assign n42639 = ~n42489 & n42568;
  assign n42640 = n42638 & ~n42639;
  assign n42641 = ~n42489 & n42543;
  assign n42642 = ~n42502 & ~n42508;
  assign n42643 = ~n42522 & n42642;
  assign n42644 = ~n42568 & ~n42643;
  assign n42645 = ~n42489 & n42514;
  assign n42646 = n42642 & n42645;
  assign n42647 = n42502 & n42553;
  assign n42648 = n42489 & n42563;
  assign n42649 = ~n42647 & ~n42648;
  assign n42650 = ~n42562 & n42649;
  assign n42651 = ~n42646 & n42650;
  assign n42652 = n42644 & n42651;
  assign n42653 = ~n42641 & n42652;
  assign n42654 = ~n42495 & ~n42653;
  assign n42655 = n42640 & ~n42654;
  assign n42656 = ~n42634 & n42655;
  assign n42657 = ~pi1078 & ~n42656;
  assign n42658 = pi1078 & n42640;
  assign n42659 = ~n42634 & n42658;
  assign n42660 = ~n42654 & n42659;
  assign po1027 = n42657 | n42660;
  assign n42662 = pi3873 & pi9040;
  assign n42663 = pi3910 & ~pi9040;
  assign n42664 = ~n42662 & ~n42663;
  assign n42665 = pi0961 & n42664;
  assign n42666 = ~pi0961 & ~n42664;
  assign n42667 = ~n42665 & ~n42666;
  assign n42668 = pi3904 & pi9040;
  assign n42669 = pi3887 & ~pi9040;
  assign n42670 = ~n42668 & ~n42669;
  assign n42671 = ~pi0991 & n42670;
  assign n42672 = pi0991 & ~n42670;
  assign n42673 = ~n42671 & ~n42672;
  assign n42674 = pi3868 & pi9040;
  assign n42675 = pi3880 & ~pi9040;
  assign n42676 = ~n42674 & ~n42675;
  assign n42677 = pi0988 & n42676;
  assign n42678 = ~pi0988 & ~n42676;
  assign n42679 = ~n42677 & ~n42678;
  assign n42680 = pi3905 & pi9040;
  assign n42681 = pi3879 & ~pi9040;
  assign n42682 = ~n42680 & ~n42681;
  assign n42683 = ~pi0963 & ~n42682;
  assign n42684 = pi0963 & ~n42680;
  assign n42685 = ~n42681 & n42684;
  assign n42686 = ~n42683 & ~n42685;
  assign n42687 = pi3879 & pi9040;
  assign n42688 = pi3911 & ~pi9040;
  assign n42689 = ~n42687 & ~n42688;
  assign n42690 = ~pi0971 & ~n42689;
  assign n42691 = pi0971 & n42689;
  assign n42692 = ~n42690 & ~n42691;
  assign n42693 = n42686 & ~n42692;
  assign n42694 = n42679 & n42693;
  assign n42695 = ~n42673 & n42694;
  assign n42696 = n42673 & n42686;
  assign n42697 = n42692 & n42696;
  assign n42698 = pi3890 & pi9040;
  assign n42699 = pi3918 & ~pi9040;
  assign n42700 = ~n42698 & ~n42699;
  assign n42701 = ~pi0970 & n42700;
  assign n42702 = pi0970 & ~n42700;
  assign n42703 = ~n42701 & ~n42702;
  assign n42704 = ~n42679 & n42696;
  assign n42705 = n42679 & n42692;
  assign n42706 = ~n42686 & n42705;
  assign n42707 = ~n42704 & ~n42706;
  assign n42708 = n42703 & ~n42707;
  assign n42709 = ~n42697 & ~n42708;
  assign n42710 = n42686 & n42705;
  assign n42711 = ~n42679 & ~n42686;
  assign n42712 = ~n42686 & ~n42692;
  assign n42713 = n42673 & n42712;
  assign n42714 = ~n42679 & ~n42692;
  assign n42715 = ~n42673 & n42714;
  assign n42716 = ~n42713 & ~n42715;
  assign n42717 = ~n42711 & n42716;
  assign n42718 = ~n42710 & n42717;
  assign n42719 = ~n42703 & ~n42718;
  assign n42720 = n42709 & ~n42719;
  assign n42721 = ~n42695 & n42720;
  assign n42722 = n42667 & ~n42721;
  assign n42723 = ~n42679 & n42692;
  assign n42724 = ~n42686 & n42723;
  assign n42725 = n42673 & n42724;
  assign n42726 = ~n42686 & n42714;
  assign n42727 = ~n42673 & n42726;
  assign n42728 = ~n42695 & ~n42727;
  assign n42729 = ~n42725 & n42728;
  assign n42730 = ~n42703 & ~n42729;
  assign n42731 = ~n42722 & ~n42730;
  assign n42732 = n42673 & n42710;
  assign n42733 = n42679 & ~n42686;
  assign n42734 = n42703 & n42733;
  assign n42735 = ~n42673 & n42734;
  assign n42736 = n42686 & n42723;
  assign n42737 = ~n42673 & n42736;
  assign n42738 = ~n42679 & n42686;
  assign n42739 = ~n42673 & n42738;
  assign n42740 = n42679 & ~n42692;
  assign n42741 = ~n42686 & n42740;
  assign n42742 = ~n42739 & ~n42741;
  assign n42743 = n42703 & ~n42742;
  assign n42744 = ~n42737 & ~n42743;
  assign n42745 = n42693 & ~n42703;
  assign n42746 = n42673 & n42745;
  assign n42747 = n42703 & n42711;
  assign n42748 = n42673 & n42747;
  assign n42749 = ~n42746 & ~n42748;
  assign n42750 = n42744 & n42749;
  assign n42751 = ~n42667 & ~n42750;
  assign n42752 = ~n42735 & ~n42751;
  assign n42753 = ~n42732 & n42752;
  assign n42754 = n42731 & n42753;
  assign n42755 = ~pi1062 & ~n42754;
  assign n42756 = ~n42722 & ~n42732;
  assign n42757 = ~n42730 & n42756;
  assign n42758 = n42752 & n42757;
  assign n42759 = pi1062 & n42758;
  assign po1028 = n42755 | n42759;
  assign n42761 = pi3881 & ~pi9040;
  assign n42762 = pi3906 & pi9040;
  assign n42763 = ~n42761 & ~n42762;
  assign n42764 = ~pi0988 & ~n42763;
  assign n42765 = pi0988 & n42763;
  assign n42766 = ~n42764 & ~n42765;
  assign n42767 = pi3893 & pi9040;
  assign n42768 = pi3869 & ~pi9040;
  assign n42769 = ~n42767 & ~n42768;
  assign n42770 = pi0982 & n42769;
  assign n42771 = ~pi0982 & ~n42769;
  assign n42772 = ~n42770 & ~n42771;
  assign n42773 = pi3923 & pi9040;
  assign n42774 = pi3877 & ~pi9040;
  assign n42775 = ~n42773 & ~n42774;
  assign n42776 = ~pi0984 & n42775;
  assign n42777 = pi0984 & ~n42775;
  assign n42778 = ~n42776 & ~n42777;
  assign n42779 = pi3881 & pi9040;
  assign n42780 = pi3901 & ~pi9040;
  assign n42781 = ~n42779 & ~n42780;
  assign n42782 = ~pi0968 & ~n42781;
  assign n42783 = pi0968 & ~n42779;
  assign n42784 = ~n42780 & n42783;
  assign n42785 = ~n42782 & ~n42784;
  assign n42786 = pi3869 & pi9040;
  assign n42787 = pi3928 & ~pi9040;
  assign n42788 = ~n42786 & ~n42787;
  assign n42789 = ~pi0963 & n42788;
  assign n42790 = pi0963 & ~n42788;
  assign n42791 = ~n42789 & ~n42790;
  assign n42792 = ~n42785 & ~n42791;
  assign n42793 = ~n42778 & n42792;
  assign n42794 = n42772 & n42793;
  assign n42795 = pi3907 & pi9040;
  assign n42796 = pi3941 & ~pi9040;
  assign n42797 = ~n42795 & ~n42796;
  assign n42798 = ~pi0969 & n42797;
  assign n42799 = pi0969 & ~n42797;
  assign n42800 = ~n42798 & ~n42799;
  assign n42801 = n42785 & ~n42791;
  assign n42802 = n42772 & n42801;
  assign n42803 = n42778 & n42792;
  assign n42804 = ~n42772 & n42803;
  assign n42805 = ~n42802 & ~n42804;
  assign n42806 = n42800 & ~n42805;
  assign n42807 = ~n42794 & ~n42806;
  assign n42808 = ~n42785 & n42791;
  assign n42809 = n42778 & n42808;
  assign n42810 = ~n42800 & n42809;
  assign n42811 = n42792 & ~n42800;
  assign n42812 = n42772 & n42811;
  assign n42813 = ~n42810 & ~n42812;
  assign n42814 = n42807 & n42813;
  assign n42815 = n42785 & n42791;
  assign n42816 = ~n42778 & n42815;
  assign n42817 = n42772 & n42816;
  assign n42818 = ~n42778 & n42808;
  assign n42819 = ~n42772 & n42818;
  assign n42820 = ~n42817 & ~n42819;
  assign n42821 = n42814 & n42820;
  assign n42822 = n42766 & ~n42821;
  assign n42823 = ~n42766 & n42800;
  assign n42824 = n42772 & n42778;
  assign n42825 = ~n42785 & n42824;
  assign n42826 = n42778 & n42791;
  assign n42827 = ~n42825 & ~n42826;
  assign n42828 = n42823 & ~n42827;
  assign n42829 = ~n42772 & ~n42778;
  assign n42830 = ~n42791 & n42829;
  assign n42831 = ~n42785 & n42830;
  assign n42832 = ~n42772 & n42785;
  assign n42833 = n42778 & n42832;
  assign n42834 = ~n42831 & ~n42833;
  assign n42835 = n42772 & ~n42800;
  assign n42836 = ~n42778 & n42835;
  assign n42837 = ~n42792 & n42836;
  assign n42838 = ~n42800 & n42816;
  assign n42839 = ~n42837 & ~n42838;
  assign n42840 = n42834 & n42839;
  assign n42841 = ~n42766 & ~n42840;
  assign n42842 = n42778 & n42815;
  assign n42843 = n42800 & n42842;
  assign n42844 = ~n42772 & n42843;
  assign n42845 = ~n42778 & n42801;
  assign n42846 = ~n42772 & n42845;
  assign n42847 = ~n42819 & ~n42846;
  assign n42848 = n42800 & ~n42847;
  assign n42849 = ~n42844 & ~n42848;
  assign n42850 = ~n42800 & n42831;
  assign n42851 = n42849 & ~n42850;
  assign n42852 = ~n42841 & n42851;
  assign n42853 = ~n42828 & n42852;
  assign n42854 = ~n42822 & n42853;
  assign n42855 = n42778 & n42801;
  assign n42856 = ~n42772 & ~n42800;
  assign n42857 = n42855 & n42856;
  assign n42858 = n42854 & ~n42857;
  assign n42859 = ~pi1081 & ~n42858;
  assign n42860 = ~n42822 & ~n42857;
  assign n42861 = pi1081 & n42860;
  assign n42862 = n42853 & n42861;
  assign po1029 = n42859 | n42862;
  assign n42864 = ~n42290 & ~n42309;
  assign n42865 = ~n42334 & ~n42349;
  assign n42866 = n42864 & ~n42865;
  assign n42867 = ~n42290 & ~n42315;
  assign n42868 = n42334 & n42867;
  assign n42869 = ~n42866 & ~n42868;
  assign n42870 = n42327 & ~n42869;
  assign n42871 = n42309 & n42315;
  assign n42872 = n42302 & n42871;
  assign n42873 = n42296 & n42872;
  assign n42874 = ~n42366 & ~n42871;
  assign n42875 = n42290 & ~n42874;
  assign n42876 = n42309 & ~n42315;
  assign n42877 = ~n42302 & n42876;
  assign n42878 = n42296 & n42877;
  assign n42879 = ~n42875 & ~n42878;
  assign n42880 = ~n42873 & n42879;
  assign n42881 = n42327 & ~n42880;
  assign n42882 = ~n42870 & ~n42881;
  assign n42883 = n42302 & n42316;
  assign n42884 = ~n42296 & n42883;
  assign n42885 = n42309 & n42341;
  assign n42886 = ~n42884 & ~n42885;
  assign n42887 = ~n42290 & ~n42886;
  assign n42888 = ~n42309 & n42357;
  assign n42889 = n42309 & n42366;
  assign n42890 = ~n42888 & ~n42889;
  assign n42891 = n42290 & ~n42890;
  assign n42892 = ~n42303 & ~n42366;
  assign n42893 = ~n42309 & ~n42892;
  assign n42894 = ~n42341 & ~n42893;
  assign n42895 = ~n42290 & ~n42894;
  assign n42896 = n42302 & n42309;
  assign n42897 = ~n42290 & n42896;
  assign n42898 = ~n42315 & n42897;
  assign n42899 = ~n42302 & n42315;
  assign n42900 = ~n42341 & ~n42899;
  assign n42901 = n42309 & ~n42900;
  assign n42902 = n42290 & ~n42309;
  assign n42903 = n42331 & n42902;
  assign n42904 = ~n42315 & n42903;
  assign n42905 = ~n42901 & ~n42904;
  assign n42906 = ~n42898 & n42905;
  assign n42907 = ~n42895 & n42906;
  assign n42908 = ~n42884 & n42907;
  assign n42909 = ~n42327 & ~n42908;
  assign n42910 = ~n42891 & ~n42909;
  assign n42911 = ~n42887 & n42910;
  assign n42912 = n42882 & n42911;
  assign n42913 = pi1072 & n42912;
  assign n42914 = ~pi1072 & ~n42912;
  assign po1031 = n42913 | n42914;
  assign n42916 = n42502 & n42515;
  assign n42917 = ~n42538 & ~n42916;
  assign n42918 = ~n42576 & n42917;
  assign n42919 = ~n42489 & ~n42918;
  assign n42920 = ~n42502 & n42522;
  assign n42921 = n42563 & n42920;
  assign n42922 = ~n42502 & n42553;
  assign n42923 = n42508 & ~n42514;
  assign n42924 = ~n42523 & ~n42923;
  assign n42925 = n42502 & ~n42924;
  assign n42926 = ~n42922 & ~n42925;
  assign n42927 = ~n42921 & n42926;
  assign n42928 = n42489 & ~n42927;
  assign n42929 = ~n42919 & ~n42928;
  assign n42930 = ~n42495 & ~n42929;
  assign n42931 = n42489 & n42550;
  assign n42932 = ~n42502 & n42931;
  assign n42933 = ~n42637 & ~n42932;
  assign n42934 = ~n42639 & n42933;
  assign n42935 = ~n42514 & n42573;
  assign n42936 = n42514 & n42642;
  assign n42937 = ~n42916 & ~n42936;
  assign n42938 = n42489 & ~n42937;
  assign n42939 = ~n42559 & ~n42938;
  assign n42940 = ~n42502 & n42524;
  assign n42941 = ~n42565 & ~n42940;
  assign n42942 = ~n42489 & n42563;
  assign n42943 = n42502 & n42942;
  assign n42944 = ~n42641 & ~n42943;
  assign n42945 = n42941 & n42944;
  assign n42946 = n42939 & n42945;
  assign n42947 = ~n42935 & n42946;
  assign n42948 = n42495 & ~n42947;
  assign n42949 = ~n42502 & n42534;
  assign n42950 = n42502 & n42526;
  assign n42951 = ~n42949 & ~n42950;
  assign n42952 = ~n42489 & ~n42951;
  assign n42953 = ~n42948 & ~n42952;
  assign n42954 = n42934 & n42953;
  assign n42955 = ~n42930 & n42954;
  assign n42956 = ~pi1065 & n42955;
  assign n42957 = pi1065 & ~n42955;
  assign po1033 = n42956 | n42957;
  assign n42959 = ~n42772 & n42809;
  assign n42960 = n42791 & n42824;
  assign n42961 = n42785 & n42960;
  assign n42962 = ~n42959 & ~n42961;
  assign n42963 = ~n42800 & ~n42962;
  assign n42964 = ~n42831 & ~n42838;
  assign n42965 = ~n42785 & n42829;
  assign n42966 = ~n42833 & ~n42965;
  assign n42967 = n42800 & ~n42966;
  assign n42968 = n42772 & n42800;
  assign n42969 = n42808 & n42968;
  assign n42970 = n42778 & n42969;
  assign n42971 = n42772 & ~n42778;
  assign n42972 = ~n42791 & n42971;
  assign n42973 = n42785 & n42972;
  assign n42974 = ~n42800 & n42803;
  assign n42975 = ~n42973 & ~n42974;
  assign n42976 = ~n42970 & n42975;
  assign n42977 = ~n42967 & n42976;
  assign n42978 = n42964 & n42977;
  assign n42979 = n42766 & ~n42978;
  assign n42980 = n42800 & n42831;
  assign n42981 = ~n42772 & n42838;
  assign n42982 = ~n42980 & ~n42981;
  assign n42983 = ~n42979 & n42982;
  assign n42984 = ~n42963 & n42983;
  assign n42985 = ~n42778 & ~n42785;
  assign n42986 = n42835 & n42985;
  assign n42987 = ~n42810 & ~n42986;
  assign n42988 = ~n42800 & n42845;
  assign n42989 = ~n42772 & n42855;
  assign n42990 = ~n42988 & ~n42989;
  assign n42991 = n42772 & n42818;
  assign n42992 = ~n42959 & ~n42991;
  assign n42993 = n42772 & n42815;
  assign n42994 = n42778 & ~n42791;
  assign n42995 = ~n42993 & ~n42994;
  assign n42996 = n42800 & ~n42995;
  assign n42997 = n42992 & ~n42996;
  assign n42998 = n42990 & n42997;
  assign n42999 = n42987 & n42998;
  assign n43000 = ~n42766 & ~n42999;
  assign n43001 = n42984 & ~n43000;
  assign n43002 = ~pi1057 & ~n43001;
  assign n43003 = pi1057 & n42984;
  assign n43004 = ~n43000 & n43003;
  assign po1034 = n43002 | n43004;
  assign n43006 = ~n42489 & n42526;
  assign n43007 = ~n42502 & n43006;
  assign n43008 = ~n42949 & ~n43007;
  assign n43009 = ~n42502 & ~n42514;
  assign n43010 = ~n42643 & ~n43009;
  assign n43011 = n42489 & ~n43010;
  assign n43012 = n42502 & ~n42508;
  assign n43013 = n42522 & n43012;
  assign n43014 = ~n43011 & ~n43013;
  assign n43015 = n43008 & n43014;
  assign n43016 = ~n42495 & ~n43015;
  assign n43017 = ~n42524 & ~n42565;
  assign n43018 = ~n42502 & n42542;
  assign n43019 = n43017 & ~n43018;
  assign n43020 = ~n42489 & ~n43019;
  assign n43021 = n42526 & n42558;
  assign n43022 = ~n42576 & ~n43021;
  assign n43023 = ~n43020 & n43022;
  assign n43024 = ~n42534 & ~n42544;
  assign n43025 = n42489 & ~n43024;
  assign n43026 = n43023 & ~n43025;
  assign n43027 = n42495 & ~n43026;
  assign n43028 = ~n43016 & ~n43027;
  assign n43029 = n42502 & n42539;
  assign n43030 = ~n42502 & ~n42533;
  assign n43031 = ~n43029 & ~n43030;
  assign n43032 = n42489 & n43031;
  assign n43033 = ~n42489 & n42502;
  assign n43034 = ~n42524 & n42625;
  assign n43035 = n43033 & ~n43034;
  assign n43036 = ~n43032 & ~n43035;
  assign n43037 = n43028 & n43036;
  assign n43038 = ~pi1058 & ~n43037;
  assign n43039 = pi1058 & n43036;
  assign n43040 = ~n43027 & n43039;
  assign n43041 = ~n43016 & n43040;
  assign po1035 = n43038 | n43041;
  assign n43043 = n42673 & n42694;
  assign n43044 = ~n42673 & n42679;
  assign n43045 = ~n42686 & n43044;
  assign n43046 = ~n42692 & n43045;
  assign n43047 = ~n43043 & ~n43046;
  assign n43048 = ~n42673 & n42723;
  assign n43049 = n42673 & n42705;
  assign n43050 = ~n43048 & ~n43049;
  assign n43051 = ~n42694 & n43050;
  assign n43052 = ~n42724 & n43051;
  assign n43053 = ~n42703 & ~n43052;
  assign n43054 = n42673 & n42706;
  assign n43055 = ~n43053 & ~n43054;
  assign n43056 = ~n42673 & n42703;
  assign n43057 = n42710 & n43056;
  assign n43058 = n42703 & n42726;
  assign n43059 = n42703 & n42736;
  assign n43060 = ~n43058 & ~n43059;
  assign n43061 = n42673 & ~n43060;
  assign n43062 = ~n43057 & ~n43061;
  assign n43063 = n43055 & n43062;
  assign n43064 = n43047 & n43063;
  assign n43065 = n42667 & ~n43064;
  assign n43066 = ~n42727 & ~n43043;
  assign n43067 = ~n42703 & ~n43066;
  assign n43068 = n42686 & n42714;
  assign n43069 = ~n42673 & n43068;
  assign n43070 = ~n42673 & n42724;
  assign n43071 = ~n43069 & ~n43070;
  assign n43072 = n42703 & ~n43071;
  assign n43073 = ~n43067 & ~n43072;
  assign n43074 = ~n42692 & n42696;
  assign n43075 = ~n42679 & n43074;
  assign n43076 = ~n42724 & ~n42732;
  assign n43077 = ~n42673 & n42693;
  assign n43078 = n42673 & n42741;
  assign n43079 = ~n43077 & ~n43078;
  assign n43080 = n43076 & n43079;
  assign n43081 = n42703 & ~n43080;
  assign n43082 = ~n42673 & n42705;
  assign n43083 = ~n42704 & ~n43082;
  assign n43084 = ~n42726 & n43083;
  assign n43085 = ~n42703 & ~n43084;
  assign n43086 = ~n42673 & n42706;
  assign n43087 = ~n43085 & ~n43086;
  assign n43088 = ~n43081 & n43087;
  assign n43089 = ~n43075 & n43088;
  assign n43090 = ~n42667 & ~n43089;
  assign n43091 = n43073 & ~n43090;
  assign n43092 = ~n43065 & n43091;
  assign n43093 = pi1077 & ~n43092;
  assign n43094 = ~pi1077 & n43092;
  assign po1036 = n43093 | n43094;
  assign n43096 = ~n42772 & n42811;
  assign n43097 = n42785 & n42824;
  assign n43098 = ~n42842 & ~n43097;
  assign n43099 = ~n42800 & ~n43098;
  assign n43100 = ~n43096 & ~n43099;
  assign n43101 = ~n42772 & n42800;
  assign n43102 = n42801 & n43101;
  assign n43103 = n42800 & n42809;
  assign n43104 = ~n43102 & ~n43103;
  assign n43105 = n43100 & n43104;
  assign n43106 = n42785 & n42829;
  assign n43107 = ~n42959 & ~n43106;
  assign n43108 = ~n42991 & n43107;
  assign n43109 = n43105 & n43108;
  assign n43110 = ~n42766 & ~n43109;
  assign n43111 = ~n42831 & ~n42842;
  assign n43112 = ~n42993 & n43111;
  assign n43113 = n42800 & ~n43112;
  assign n43114 = ~n42791 & n42824;
  assign n43115 = ~n42785 & n43114;
  assign n43116 = ~n42973 & ~n43115;
  assign n43117 = ~n42857 & n43116;
  assign n43118 = ~n42800 & n42818;
  assign n43119 = n43117 & ~n43118;
  assign n43120 = ~n43113 & n43119;
  assign n43121 = n42766 & ~n43120;
  assign n43122 = ~n42981 & ~n42986;
  assign n43123 = ~n42959 & n43116;
  assign n43124 = n42800 & ~n43123;
  assign n43125 = n43122 & ~n43124;
  assign n43126 = ~n43121 & n43125;
  assign n43127 = ~n43110 & n43126;
  assign n43128 = pi1086 & ~n43127;
  assign n43129 = ~pi1086 & n43127;
  assign po1037 = n43128 | n43129;
  assign n43131 = n42673 & n42703;
  assign n43132 = n42679 & n43131;
  assign n43133 = n42673 & ~n42686;
  assign n43134 = ~n42692 & n43133;
  assign n43135 = ~n42679 & n43134;
  assign n43136 = ~n42706 & ~n43135;
  assign n43137 = ~n42703 & ~n43136;
  assign n43138 = n43071 & ~n43137;
  assign n43139 = ~n43132 & n43138;
  assign n43140 = n42667 & ~n43139;
  assign n43141 = n42703 & n43046;
  assign n43142 = n42673 & ~n42703;
  assign n43143 = n42741 & n43142;
  assign n43144 = ~n42704 & ~n43143;
  assign n43145 = ~n42706 & ~n42736;
  assign n43146 = n42673 & n42723;
  assign n43147 = n43145 & ~n43146;
  assign n43148 = n42703 & ~n43147;
  assign n43149 = ~n42703 & n42710;
  assign n43150 = n42728 & ~n43149;
  assign n43151 = ~n43148 & n43150;
  assign n43152 = n43144 & n43151;
  assign n43153 = ~n42667 & ~n43152;
  assign n43154 = ~n43141 & ~n43153;
  assign n43155 = ~n43140 & n43154;
  assign n43156 = n42736 & n43142;
  assign n43157 = ~n42673 & n42745;
  assign n43158 = ~n43156 & ~n43157;
  assign n43159 = ~n42703 & n43070;
  assign n43160 = n43158 & ~n43159;
  assign n43161 = n43155 & n43160;
  assign n43162 = ~pi1063 & ~n43161;
  assign n43163 = pi1063 & n43160;
  assign n43164 = n43154 & n43163;
  assign n43165 = ~n43140 & n43164;
  assign po1039 = n43162 | n43165;
  assign n43167 = ~n42407 & n42441;
  assign n43168 = ~n42593 & ~n43167;
  assign n43169 = n42413 & ~n43168;
  assign n43170 = n42436 & n42589;
  assign n43171 = ~n43169 & ~n43170;
  assign n43172 = ~n42461 & n43171;
  assign n43173 = n42394 & n42407;
  assign n43174 = n42387 & n43173;
  assign n43175 = n42400 & n43174;
  assign n43176 = ~n42421 & ~n43175;
  assign n43177 = ~n42441 & n43176;
  assign n43178 = n42413 & ~n43177;
  assign n43179 = n42381 & n43178;
  assign n43180 = ~n42413 & n42602;
  assign n43181 = ~n42432 & ~n42459;
  assign n43182 = ~n42426 & n43181;
  assign n43183 = ~n43180 & n43182;
  assign n43184 = n42381 & ~n43183;
  assign n43185 = ~n42387 & ~n42413;
  assign n43186 = n42400 & n43185;
  assign n43187 = ~n42394 & n43186;
  assign n43188 = ~n42407 & n43187;
  assign n43189 = n42407 & n42473;
  assign n43190 = ~n43187 & ~n43189;
  assign n43191 = ~n42592 & n43190;
  assign n43192 = n42400 & n42430;
  assign n43193 = n42407 & n42418;
  assign n43194 = ~n42435 & ~n43193;
  assign n43195 = n42413 & ~n43194;
  assign n43196 = ~n43192 & ~n43195;
  assign n43197 = n43191 & n43196;
  assign n43198 = ~n42381 & ~n43197;
  assign n43199 = ~n43188 & ~n43198;
  assign n43200 = ~n43184 & n43199;
  assign n43201 = ~n43179 & n43200;
  assign n43202 = n43172 & n43201;
  assign n43203 = pi1096 & ~n43202;
  assign n43204 = ~pi1096 & n43172;
  assign n43205 = n43201 & n43204;
  assign po1040 = n43203 | n43205;
  assign n43207 = pi3886 & pi9040;
  assign n43208 = pi3878 & ~pi9040;
  assign n43209 = ~n43207 & ~n43208;
  assign n43210 = ~pi0962 & n43209;
  assign n43211 = pi0962 & ~n43209;
  assign n43212 = ~n43210 & ~n43211;
  assign n43213 = pi3941 & pi9040;
  assign n43214 = pi3925 & ~pi9040;
  assign n43215 = ~n43213 & ~n43214;
  assign n43216 = ~pi0979 & n43215;
  assign n43217 = pi0979 & ~n43215;
  assign n43218 = ~n43216 & ~n43217;
  assign n43219 = ~n43212 & ~n43218;
  assign n43220 = pi3901 & pi9040;
  assign n43221 = pi3876 & ~pi9040;
  assign n43222 = ~n43220 & ~n43221;
  assign n43223 = pi0967 & n43222;
  assign n43224 = ~pi0967 & ~n43222;
  assign n43225 = ~n43223 & ~n43224;
  assign n43226 = pi3874 & pi9040;
  assign n43227 = pi3899 & ~pi9040;
  assign n43228 = ~n43226 & ~n43227;
  assign n43229 = pi0984 & n43228;
  assign n43230 = ~pi0984 & ~n43228;
  assign n43231 = ~n43229 & ~n43230;
  assign n43232 = n43218 & ~n43231;
  assign n43233 = n43225 & n43232;
  assign n43234 = ~n43219 & ~n43233;
  assign n43235 = pi3925 & pi9040;
  assign n43236 = pi3920 & ~pi9040;
  assign n43237 = ~n43235 & ~n43236;
  assign n43238 = ~pi0968 & n43237;
  assign n43239 = pi0968 & ~n43237;
  assign n43240 = ~n43238 & ~n43239;
  assign n43241 = pi3894 & pi9040;
  assign n43242 = pi3923 & ~pi9040;
  assign n43243 = ~n43241 & ~n43242;
  assign n43244 = pi0974 & n43243;
  assign n43245 = ~pi0974 & ~n43243;
  assign n43246 = ~n43244 & ~n43245;
  assign n43247 = ~n43240 & ~n43246;
  assign n43248 = ~n43234 & n43247;
  assign n43249 = ~n43218 & n43231;
  assign n43250 = ~n43212 & n43225;
  assign n43251 = ~n43249 & n43250;
  assign n43252 = ~n43240 & n43251;
  assign n43253 = ~n43212 & ~n43225;
  assign n43254 = n43246 & n43253;
  assign n43255 = n43249 & n43254;
  assign n43256 = ~n43212 & ~n43246;
  assign n43257 = n43225 & n43256;
  assign n43258 = ~n43231 & n43257;
  assign n43259 = ~n43255 & ~n43258;
  assign n43260 = ~n43252 & n43259;
  assign n43261 = ~n43212 & n43232;
  assign n43262 = n43218 & n43231;
  assign n43263 = n43212 & n43262;
  assign n43264 = ~n43261 & ~n43263;
  assign n43265 = n43246 & ~n43264;
  assign n43266 = ~n43218 & ~n43231;
  assign n43267 = n43212 & n43246;
  assign n43268 = n43266 & n43267;
  assign n43269 = ~n43225 & n43268;
  assign n43270 = ~n43265 & ~n43269;
  assign n43271 = ~n43240 & ~n43270;
  assign n43272 = n43212 & ~n43225;
  assign n43273 = ~n43232 & ~n43249;
  assign n43274 = n43272 & ~n43273;
  assign n43275 = ~n43218 & ~n43225;
  assign n43276 = ~n43249 & ~n43275;
  assign n43277 = n43212 & ~n43276;
  assign n43278 = n43225 & n43262;
  assign n43279 = ~n43277 & ~n43278;
  assign n43280 = ~n43246 & ~n43279;
  assign n43281 = ~n43274 & ~n43280;
  assign n43282 = ~n43225 & n43262;
  assign n43283 = ~n43212 & n43282;
  assign n43284 = n43212 & n43225;
  assign n43285 = ~n43231 & n43284;
  assign n43286 = ~n43212 & ~n43276;
  assign n43287 = ~n43285 & ~n43286;
  assign n43288 = n43246 & ~n43287;
  assign n43289 = ~n43283 & ~n43288;
  assign n43290 = n43281 & n43289;
  assign n43291 = n43240 & ~n43290;
  assign n43292 = ~n43271 & ~n43291;
  assign n43293 = n43260 & n43292;
  assign n43294 = ~n43248 & n43293;
  assign n43295 = pi1093 & ~n43294;
  assign n43296 = ~pi1093 & n43260;
  assign n43297 = ~n43248 & n43296;
  assign n43298 = n43292 & n43297;
  assign po1041 = n43295 | n43298;
  assign n43300 = pi3903 & pi9040;
  assign n43301 = pi3904 & ~pi9040;
  assign n43302 = ~n43300 & ~n43301;
  assign n43303 = pi0981 & n43302;
  assign n43304 = ~pi0981 & ~n43302;
  assign n43305 = ~n43303 & ~n43304;
  assign n43306 = pi3927 & ~pi9040;
  assign n43307 = pi3891 & pi9040;
  assign n43308 = ~n43306 & ~n43307;
  assign n43309 = ~pi0958 & n43308;
  assign n43310 = pi0958 & ~n43308;
  assign n43311 = ~n43309 & ~n43310;
  assign n43312 = pi3896 & pi9040;
  assign n43313 = pi3905 & ~pi9040;
  assign n43314 = ~n43312 & ~n43313;
  assign n43315 = ~pi0983 & ~n43314;
  assign n43316 = pi0983 & ~n43312;
  assign n43317 = ~n43313 & n43316;
  assign n43318 = ~n43315 & ~n43317;
  assign n43319 = pi3880 & pi9040;
  assign n43320 = pi3873 & ~pi9040;
  assign n43321 = ~n43319 & ~n43320;
  assign n43322 = ~pi0989 & n43321;
  assign n43323 = pi0989 & ~n43321;
  assign n43324 = ~n43322 & ~n43323;
  assign n43325 = pi3916 & pi9040;
  assign n43326 = pi3903 & ~pi9040;
  assign n43327 = ~n43325 & ~n43326;
  assign n43328 = ~pi0973 & n43327;
  assign n43329 = pi0973 & ~n43327;
  assign n43330 = ~n43328 & ~n43329;
  assign n43331 = n43324 & ~n43330;
  assign n43332 = ~n43318 & n43331;
  assign n43333 = ~n43311 & n43332;
  assign n43334 = ~n43324 & n43330;
  assign n43335 = ~n43318 & n43334;
  assign n43336 = n43324 & n43330;
  assign n43337 = n43318 & n43336;
  assign n43338 = ~n43311 & n43337;
  assign n43339 = ~n43335 & ~n43338;
  assign n43340 = ~n43333 & n43339;
  assign n43341 = n43305 & ~n43340;
  assign n43342 = n43318 & n43324;
  assign n43343 = n43311 & n43342;
  assign n43344 = n43318 & ~n43324;
  assign n43345 = ~n43311 & n43344;
  assign n43346 = ~n43343 & ~n43345;
  assign n43347 = ~n43305 & ~n43346;
  assign n43348 = ~n43341 & ~n43347;
  assign n43349 = pi3887 & pi9040;
  assign n43350 = pi3890 & ~pi9040;
  assign n43351 = ~n43349 & ~n43350;
  assign n43352 = ~pi0972 & ~n43351;
  assign n43353 = pi0972 & n43351;
  assign n43354 = ~n43352 & ~n43353;
  assign n43355 = n43318 & n43331;
  assign n43356 = ~n43318 & ~n43330;
  assign n43357 = n43311 & n43356;
  assign n43358 = ~n43324 & n43357;
  assign n43359 = ~n43355 & ~n43358;
  assign n43360 = ~n43305 & ~n43359;
  assign n43361 = n43311 & ~n43318;
  assign n43362 = n43330 & n43361;
  assign n43363 = n43324 & n43362;
  assign n43364 = ~n43333 & ~n43363;
  assign n43365 = ~n43311 & ~n43318;
  assign n43366 = ~n43324 & n43365;
  assign n43367 = ~n43324 & ~n43330;
  assign n43368 = n43318 & n43367;
  assign n43369 = n43311 & n43368;
  assign n43370 = ~n43366 & ~n43369;
  assign n43371 = n43305 & ~n43370;
  assign n43372 = n43364 & ~n43371;
  assign n43373 = ~n43360 & n43372;
  assign n43374 = n43354 & ~n43373;
  assign n43375 = ~n43305 & n43311;
  assign n43376 = n43331 & n43375;
  assign n43377 = n43318 & n43334;
  assign n43378 = n43330 & n43365;
  assign n43379 = n43324 & n43378;
  assign n43380 = ~n43377 & ~n43379;
  assign n43381 = ~n43311 & n43367;
  assign n43382 = n43380 & ~n43381;
  assign n43383 = ~n43305 & ~n43382;
  assign n43384 = ~n43318 & ~n43324;
  assign n43385 = n43305 & n43311;
  assign n43386 = n43384 & n43385;
  assign n43387 = n43311 & n43335;
  assign n43388 = ~n43386 & ~n43387;
  assign n43389 = ~n43383 & n43388;
  assign n43390 = ~n43376 & n43389;
  assign n43391 = n43311 & n43355;
  assign n43392 = ~n43311 & n43368;
  assign n43393 = ~n43391 & ~n43392;
  assign n43394 = n43390 & n43393;
  assign n43395 = ~n43354 & ~n43394;
  assign n43396 = ~n43318 & n43330;
  assign n43397 = n43305 & n43396;
  assign n43398 = n43311 & n43397;
  assign n43399 = ~n43395 & ~n43398;
  assign n43400 = ~n43374 & n43399;
  assign n43401 = n43348 & n43400;
  assign n43402 = ~pi1076 & ~n43401;
  assign n43403 = pi1076 & n43401;
  assign po1042 = n43402 | n43403;
  assign n43405 = ~n42302 & n42318;
  assign n43406 = ~n42349 & ~n43405;
  assign n43407 = ~n42290 & ~n43406;
  assign n43408 = ~n42309 & n42340;
  assign n43409 = ~n42877 & ~n43408;
  assign n43410 = n42290 & ~n43409;
  assign n43411 = n42309 & n42335;
  assign n43412 = ~n42898 & ~n43411;
  assign n43413 = ~n42317 & n43412;
  assign n43414 = ~n43410 & n43413;
  assign n43415 = ~n43407 & n43414;
  assign n43416 = ~n42873 & ~n42884;
  assign n43417 = n43415 & n43416;
  assign n43418 = n42327 & ~n43417;
  assign n43419 = n42303 & n42871;
  assign n43420 = n42358 & ~n43419;
  assign n43421 = n42290 & ~n43420;
  assign n43422 = n42309 & n42346;
  assign n43423 = ~n43421 & ~n43422;
  assign n43424 = n42296 & n42318;
  assign n43425 = ~n42309 & n42331;
  assign n43426 = ~n43424 & ~n43425;
  assign n43427 = n42290 & ~n43426;
  assign n43428 = n42290 & n42340;
  assign n43429 = n42309 & n43428;
  assign n43430 = ~n43427 & ~n43429;
  assign n43431 = n43423 & n43430;
  assign n43432 = ~n42327 & ~n43431;
  assign n43433 = ~n42335 & ~n42342;
  assign n43434 = ~n42878 & n43433;
  assign n43435 = n42363 & ~n43434;
  assign n43436 = ~n43432 & ~n43435;
  assign n43437 = ~n42317 & ~n42873;
  assign n43438 = ~n42290 & ~n43437;
  assign n43439 = n43436 & ~n43438;
  assign n43440 = ~n43418 & n43439;
  assign n43441 = ~pi1087 & n43440;
  assign n43442 = pi1087 & ~n43440;
  assign po1044 = n43441 | n43442;
  assign n43444 = ~n43225 & n43266;
  assign n43445 = n43225 & n43249;
  assign n43446 = ~n43444 & ~n43445;
  assign n43447 = n43231 & n43284;
  assign n43448 = n43446 & ~n43447;
  assign n43449 = n43247 & ~n43448;
  assign n43450 = n43233 & ~n43240;
  assign n43451 = ~n43212 & n43450;
  assign n43452 = n43225 & n43266;
  assign n43453 = n43246 & n43452;
  assign n43454 = ~n43225 & n43231;
  assign n43455 = ~n43212 & n43262;
  assign n43456 = ~n43454 & ~n43455;
  assign n43457 = n43246 & ~n43456;
  assign n43458 = ~n43453 & ~n43457;
  assign n43459 = ~n43240 & ~n43458;
  assign n43460 = ~n43451 & ~n43459;
  assign n43461 = n43231 & n43253;
  assign n43462 = ~n43231 & n43272;
  assign n43463 = n43218 & n43462;
  assign n43464 = ~n43461 & ~n43463;
  assign n43465 = n43246 & ~n43464;
  assign n43466 = n43460 & ~n43465;
  assign n43467 = n43256 & n43262;
  assign n43468 = n43225 & n43467;
  assign n43469 = n43212 & ~n43246;
  assign n43470 = n43282 & n43469;
  assign n43471 = ~n43273 & n43284;
  assign n43472 = n43212 & n43444;
  assign n43473 = ~n43471 & ~n43472;
  assign n43474 = n43253 & ~n43273;
  assign n43475 = ~n43212 & n43452;
  assign n43476 = ~n43474 & ~n43475;
  assign n43477 = n43473 & n43476;
  assign n43478 = ~n43470 & n43477;
  assign n43479 = ~n43468 & n43478;
  assign n43480 = n43225 & n43267;
  assign n43481 = n43218 & n43480;
  assign n43482 = n43479 & ~n43481;
  assign n43483 = n43240 & ~n43482;
  assign n43484 = n43466 & ~n43483;
  assign n43485 = ~n43449 & n43484;
  assign n43486 = ~pi1084 & ~n43485;
  assign n43487 = pi1084 & n43466;
  assign n43488 = ~n43449 & n43487;
  assign n43489 = ~n43483 & n43488;
  assign po1045 = n43486 | n43489;
  assign n43491 = ~n43225 & n43249;
  assign n43492 = ~n43278 & ~n43491;
  assign n43493 = n43246 & ~n43492;
  assign n43494 = n43212 & n43232;
  assign n43495 = ~n43445 & ~n43494;
  assign n43496 = ~n43282 & n43495;
  assign n43497 = ~n43246 & ~n43496;
  assign n43498 = ~n43493 & ~n43497;
  assign n43499 = ~n43453 & ~n43463;
  assign n43500 = n43498 & n43499;
  assign n43501 = n43240 & ~n43500;
  assign n43502 = n43225 & n43246;
  assign n43503 = ~n43231 & n43502;
  assign n43504 = n43218 & n43503;
  assign n43505 = n43446 & ~n43504;
  assign n43506 = ~n43282 & n43505;
  assign n43507 = n43212 & ~n43506;
  assign n43508 = ~n43212 & n43278;
  assign n43509 = n43212 & n43266;
  assign n43510 = ~n43261 & ~n43509;
  assign n43511 = ~n43246 & ~n43510;
  assign n43512 = ~n43508 & ~n43511;
  assign n43513 = ~n43507 & n43512;
  assign n43514 = ~n43240 & ~n43513;
  assign n43515 = ~n43501 & ~n43514;
  assign n43516 = ~n43225 & n43261;
  assign n43517 = ~n43475 & ~n43516;
  assign n43518 = n43246 & ~n43517;
  assign n43519 = n43256 & n43275;
  assign n43520 = ~n43518 & ~n43519;
  assign n43521 = n43515 & n43520;
  assign n43522 = ~pi1064 & ~n43521;
  assign n43523 = pi1064 & ~n43518;
  assign n43524 = n43515 & n43523;
  assign n43525 = ~n43519 & n43524;
  assign po1046 = n43522 | n43525;
  assign n43527 = n43246 & n43278;
  assign n43528 = n43212 & n43527;
  assign n43529 = ~n43269 & ~n43528;
  assign n43530 = ~n43470 & ~n43472;
  assign n43531 = n43219 & n43225;
  assign n43532 = ~n43455 & ~n43531;
  assign n43533 = n43246 & ~n43532;
  assign n43534 = ~n43246 & ~n43272;
  assign n43535 = ~n43273 & n43534;
  assign n43536 = ~n43225 & ~n43262;
  assign n43537 = n43246 & n43536;
  assign n43538 = n43212 & n43537;
  assign n43539 = ~n43535 & ~n43538;
  assign n43540 = ~n43533 & n43539;
  assign n43541 = n43530 & n43540;
  assign n43542 = ~n43240 & ~n43541;
  assign n43543 = n43529 & ~n43542;
  assign n43544 = ~n43246 & n43445;
  assign n43545 = ~n43212 & n43544;
  assign n43546 = n43240 & ~n43246;
  assign n43547 = ~n43274 & ~n43455;
  assign n43548 = ~n43452 & n43547;
  assign n43549 = n43546 & ~n43548;
  assign n43550 = ~n43212 & n43444;
  assign n43551 = n43219 & ~n43225;
  assign n43552 = ~n43261 & ~n43551;
  assign n43553 = ~n43233 & ~n43263;
  assign n43554 = n43552 & n43553;
  assign n43555 = n43246 & ~n43554;
  assign n43556 = ~n43550 & ~n43555;
  assign n43557 = n43240 & ~n43556;
  assign n43558 = ~n43549 & ~n43557;
  assign n43559 = ~n43545 & n43558;
  assign n43560 = n43543 & n43559;
  assign n43561 = pi1070 & ~n43560;
  assign n43562 = ~pi1070 & n43543;
  assign n43563 = n43559 & n43562;
  assign po1047 = n43561 | n43563;
  assign n43565 = n42407 & ~n42614;
  assign n43566 = n42387 & n43565;
  assign n43567 = n42400 & n42591;
  assign n43568 = ~n42469 & ~n43567;
  assign n43569 = ~n42421 & n43568;
  assign n43570 = ~n42413 & ~n43569;
  assign n43571 = ~n42445 & ~n42602;
  assign n43572 = n42413 & ~n43571;
  assign n43573 = ~n43570 & ~n43572;
  assign n43574 = ~n43566 & n43573;
  assign n43575 = ~n42407 & n42436;
  assign n43576 = n43574 & ~n43575;
  assign n43577 = ~n42381 & ~n43576;
  assign n43578 = n42417 & ~n43571;
  assign n43579 = ~n42441 & ~n42446;
  assign n43580 = ~n42421 & ~n42436;
  assign n43581 = n43579 & n43580;
  assign n43582 = n42407 & ~n43581;
  assign n43583 = ~n43578 & ~n43582;
  assign n43584 = ~n42593 & n43583;
  assign n43585 = n42381 & ~n43584;
  assign n43586 = ~n43577 & ~n43585;
  assign n43587 = n42407 & n42602;
  assign n43588 = ~n43575 & ~n43587;
  assign n43589 = n42413 & ~n43588;
  assign n43590 = n43586 & ~n43589;
  assign n43591 = pi1069 & ~n43590;
  assign n43592 = ~pi1069 & ~n43589;
  assign n43593 = ~n43585 & n43592;
  assign n43594 = ~n43577 & n43593;
  assign po1048 = n43591 | n43594;
  assign n43596 = ~n42290 & n42346;
  assign n43597 = n42309 & n42331;
  assign n43598 = ~n42330 & ~n43597;
  assign n43599 = ~n42290 & ~n43598;
  assign n43600 = n42290 & ~n42900;
  assign n43601 = ~n43599 & ~n43600;
  assign n43602 = ~n42888 & n43601;
  assign n43603 = n42327 & ~n43602;
  assign n43604 = ~n43596 & ~n43603;
  assign n43605 = n42315 & n42864;
  assign n43606 = ~n42876 & ~n43605;
  assign n43607 = ~n42296 & ~n43606;
  assign n43608 = ~n42317 & ~n43607;
  assign n43609 = ~n42877 & n43608;
  assign n43610 = ~n42309 & n42349;
  assign n43611 = n42290 & n42332;
  assign n43612 = ~n43610 & ~n43611;
  assign n43613 = n43609 & n43612;
  assign n43614 = ~n42327 & ~n43613;
  assign n43615 = ~n43411 & ~n43425;
  assign n43616 = n42290 & ~n43615;
  assign n43617 = ~n43614 & ~n43616;
  assign n43618 = n43604 & n43617;
  assign n43619 = ~pi1141 & ~n43618;
  assign n43620 = ~n43603 & n43617;
  assign n43621 = pi1141 & n43620;
  assign n43622 = ~n43596 & n43621;
  assign po1049 = n43619 | n43622;
  assign n43624 = ~n43344 & ~n43363;
  assign n43625 = n43305 & ~n43624;
  assign n43626 = ~n43324 & n43378;
  assign n43627 = ~n43625 & ~n43626;
  assign n43628 = ~n43358 & n43627;
  assign n43629 = ~n43305 & n43333;
  assign n43630 = ~n43391 & ~n43629;
  assign n43631 = ~n43338 & n43630;
  assign n43632 = n43628 & n43631;
  assign n43633 = n43354 & ~n43632;
  assign n43634 = ~n43318 & n43367;
  assign n43635 = ~n43311 & n43634;
  assign n43636 = ~n43379 & ~n43635;
  assign n43637 = n43311 & n43337;
  assign n43638 = ~n43387 & ~n43637;
  assign n43639 = n43318 & ~n43330;
  assign n43640 = ~n43311 & ~n43324;
  assign n43641 = ~n43639 & ~n43640;
  assign n43642 = ~n43396 & n43641;
  assign n43643 = ~n43305 & ~n43642;
  assign n43644 = n43305 & n43332;
  assign n43645 = ~n43311 & n43355;
  assign n43646 = ~n43644 & ~n43645;
  assign n43647 = ~n43643 & n43646;
  assign n43648 = n43638 & n43647;
  assign n43649 = n43636 & n43648;
  assign n43650 = ~n43354 & ~n43649;
  assign n43651 = ~n43633 & ~n43650;
  assign n43652 = pi1056 & ~n43651;
  assign n43653 = ~pi1056 & ~n43633;
  assign n43654 = ~n43650 & n43653;
  assign po1050 = n43652 | n43654;
  assign n43656 = ~n42817 & ~n42825;
  assign n43657 = n42766 & ~n43656;
  assign n43658 = ~n42830 & ~n42965;
  assign n43659 = n42800 & ~n43658;
  assign n43660 = n42793 & n42800;
  assign n43661 = ~n43659 & ~n43660;
  assign n43662 = n42766 & ~n43661;
  assign n43663 = ~n43657 & ~n43662;
  assign n43664 = n42816 & n42968;
  assign n43665 = ~n42970 & ~n43664;
  assign n43666 = ~n42833 & ~n42994;
  assign n43667 = ~n42800 & ~n43666;
  assign n43668 = n42766 & n43667;
  assign n43669 = n43665 & ~n43668;
  assign n43670 = ~n42772 & n42816;
  assign n43671 = ~n42772 & n42808;
  assign n43672 = ~n42961 & ~n43671;
  assign n43673 = ~n42800 & ~n43672;
  assign n43674 = ~n42831 & ~n42973;
  assign n43675 = ~n42772 & n42815;
  assign n43676 = ~n42855 & ~n43675;
  assign n43677 = n42800 & ~n43676;
  assign n43678 = n43674 & ~n43677;
  assign n43679 = ~n43673 & n43678;
  assign n43680 = ~n43670 & n43679;
  assign n43681 = ~n42766 & ~n43680;
  assign n43682 = ~n42991 & n43116;
  assign n43683 = ~n42800 & ~n43682;
  assign n43684 = ~n43681 & ~n43683;
  assign n43685 = n43669 & n43684;
  assign n43686 = n43663 & n43685;
  assign n43687 = ~pi1079 & ~n43686;
  assign n43688 = pi1079 & n43669;
  assign n43689 = n43663 & n43688;
  assign n43690 = n43684 & n43689;
  assign po1051 = n43687 | n43690;
  assign n43692 = ~n42215 & n42245;
  assign n43693 = n42215 & n42256;
  assign n43694 = ~n42242 & ~n43693;
  assign n43695 = n42187 & ~n43694;
  assign n43696 = ~n43692 & ~n43695;
  assign n43697 = ~n42187 & ~n42215;
  assign n43698 = ~n42207 & n43697;
  assign n43699 = n42201 & n43698;
  assign n43700 = n42223 & n42257;
  assign n43701 = ~n43699 & ~n43700;
  assign n43702 = ~n42187 & n42266;
  assign n43703 = n43701 & ~n43702;
  assign n43704 = ~n42219 & ~n42231;
  assign n43705 = n42207 & n42221;
  assign n43706 = n43704 & ~n43705;
  assign n43707 = n43703 & n43706;
  assign n43708 = n43696 & n43707;
  assign n43709 = ~n42254 & ~n43708;
  assign n43710 = ~n42194 & n42217;
  assign n43711 = ~n42242 & ~n43710;
  assign n43712 = n42215 & ~n43711;
  assign n43713 = n42201 & n42260;
  assign n43714 = ~n42271 & ~n43713;
  assign n43715 = n42194 & ~n42207;
  assign n43716 = n42215 & n43715;
  assign n43717 = n43714 & ~n43716;
  assign n43718 = n42187 & ~n43717;
  assign n43719 = ~n42215 & n42241;
  assign n43720 = n42201 & n42230;
  assign n43721 = ~n43719 & ~n43720;
  assign n43722 = ~n42187 & ~n43721;
  assign n43723 = ~n42215 & n42224;
  assign n43724 = ~n43722 & ~n43723;
  assign n43725 = ~n43718 & n43724;
  assign n43726 = ~n43712 & n43725;
  assign n43727 = n42254 & ~n43726;
  assign n43728 = n42187 & n42261;
  assign n43729 = ~n43727 & ~n43728;
  assign n43730 = n42236 & n43697;
  assign n43731 = ~n42207 & n43730;
  assign n43732 = n43729 & ~n43731;
  assign n43733 = ~n43709 & n43732;
  assign n43734 = ~pi1067 & ~n43733;
  assign n43735 = pi1067 & n43729;
  assign n43736 = ~n43709 & n43735;
  assign n43737 = ~n43731 & n43736;
  assign po1052 = n43734 | n43737;
  assign n43739 = ~n43043 & ~n43135;
  assign n43740 = ~n43086 & n43739;
  assign n43741 = n42703 & ~n43740;
  assign n43742 = ~n43143 & ~n43159;
  assign n43743 = ~n43046 & ~n43059;
  assign n43744 = ~n43049 & ~n43068;
  assign n43745 = ~n42703 & ~n43744;
  assign n43746 = ~n42732 & ~n43745;
  assign n43747 = n43743 & n43746;
  assign n43748 = n42667 & ~n43747;
  assign n43749 = ~n42686 & n42692;
  assign n43750 = ~n42711 & ~n43749;
  assign n43751 = ~n42673 & ~n43750;
  assign n43752 = ~n42694 & ~n43146;
  assign n43753 = ~n42703 & ~n43752;
  assign n43754 = ~n42673 & n42692;
  assign n43755 = ~n42706 & ~n43754;
  assign n43756 = ~n42714 & n43755;
  assign n43757 = n42703 & ~n43756;
  assign n43758 = ~n43753 & ~n43757;
  assign n43759 = ~n43751 & n43758;
  assign n43760 = ~n42667 & ~n43759;
  assign n43761 = ~n43748 & ~n43760;
  assign n43762 = n43742 & n43761;
  assign n43763 = ~n43741 & n43762;
  assign n43764 = ~pi1107 & ~n43763;
  assign n43765 = pi1107 & n43742;
  assign n43766 = ~n43741 & n43765;
  assign n43767 = n43761 & n43766;
  assign po1053 = n43764 | n43767;
  assign n43769 = ~n42194 & n42201;
  assign n43770 = ~n42187 & n43769;
  assign n43771 = n42215 & n43770;
  assign n43772 = ~n42215 & n43715;
  assign n43773 = ~n42222 & ~n43772;
  assign n43774 = ~n43720 & n43773;
  assign n43775 = ~n43771 & n43774;
  assign n43776 = n42187 & n43710;
  assign n43777 = n43775 & ~n43776;
  assign n43778 = n42254 & ~n43777;
  assign n43779 = ~n42272 & ~n43723;
  assign n43780 = n42187 & ~n43779;
  assign n43781 = ~n42254 & n42256;
  assign n43782 = ~n42187 & n43781;
  assign n43783 = n42194 & ~n42215;
  assign n43784 = ~n42201 & n43783;
  assign n43785 = ~n43715 & ~n43784;
  assign n43786 = ~n42224 & n43785;
  assign n43787 = n42187 & ~n43786;
  assign n43788 = ~n42194 & n42241;
  assign n43789 = ~n42215 & n43788;
  assign n43790 = ~n43787 & ~n43789;
  assign n43791 = ~n42254 & ~n43790;
  assign n43792 = ~n43782 & ~n43791;
  assign n43793 = ~n43780 & n43792;
  assign n43794 = ~n42215 & n42271;
  assign n43795 = ~n43693 & ~n43794;
  assign n43796 = ~n42219 & ~n42222;
  assign n43797 = n43795 & n43796;
  assign n43798 = ~n42187 & ~n43797;
  assign n43799 = n43793 & ~n43798;
  assign n43800 = ~n43778 & n43799;
  assign n43801 = ~pi1088 & ~n43800;
  assign n43802 = pi1088 & n43793;
  assign n43803 = ~n43778 & n43802;
  assign n43804 = ~n43798 & n43803;
  assign po1054 = n43801 | n43804;
  assign n43806 = ~n42216 & ~n42222;
  assign n43807 = ~n42187 & ~n43806;
  assign n43808 = ~n42278 & ~n43807;
  assign n43809 = ~n42194 & ~n42201;
  assign n43810 = n42187 & n43809;
  assign n43811 = n42215 & n43810;
  assign n43812 = ~n42187 & n42208;
  assign n43813 = n42215 & n43812;
  assign n43814 = ~n43702 & ~n43813;
  assign n43815 = n42201 & n43783;
  assign n43816 = n42215 & n42241;
  assign n43817 = ~n43815 & ~n43816;
  assign n43818 = ~n43809 & n43817;
  assign n43819 = n42187 & ~n43818;
  assign n43820 = ~n42225 & ~n43819;
  assign n43821 = n43814 & n43820;
  assign n43822 = ~n42254 & ~n43821;
  assign n43823 = ~n43811 & ~n43822;
  assign n43824 = ~n42242 & ~n42261;
  assign n43825 = ~n42271 & n43824;
  assign n43826 = ~n42187 & ~n43825;
  assign n43827 = ~n42215 & n42266;
  assign n43828 = ~n42245 & ~n43827;
  assign n43829 = n42187 & ~n43828;
  assign n43830 = ~n43713 & ~n43829;
  assign n43831 = ~n43826 & n43830;
  assign n43832 = ~n42231 & ~n42272;
  assign n43833 = n43831 & n43832;
  assign n43834 = n42254 & ~n43833;
  assign n43835 = n43823 & ~n43834;
  assign n43836 = n43808 & n43835;
  assign n43837 = ~pi1075 & ~n43836;
  assign n43838 = pi1075 & n43823;
  assign n43839 = n43808 & n43838;
  assign n43840 = ~n43834 & n43839;
  assign po1055 = n43837 | n43840;
  assign n43842 = n43311 & n43367;
  assign n43843 = ~n43637 & ~n43842;
  assign n43844 = n43305 & n43843;
  assign n43845 = ~n43311 & n43342;
  assign n43846 = ~n43331 & ~n43334;
  assign n43847 = n43318 & ~n43846;
  assign n43848 = n43324 & n43361;
  assign n43849 = ~n43311 & n43334;
  assign n43850 = ~n43848 & ~n43849;
  assign n43851 = ~n43847 & n43850;
  assign n43852 = ~n43305 & n43851;
  assign n43853 = ~n43845 & n43852;
  assign n43854 = ~n43844 & ~n43853;
  assign n43855 = ~n43311 & n43847;
  assign n43856 = ~n43635 & ~n43855;
  assign n43857 = ~n43854 & n43856;
  assign n43858 = n43354 & ~n43857;
  assign n43859 = n43305 & ~n43846;
  assign n43860 = n43311 & n43859;
  assign n43861 = ~n43311 & n43336;
  assign n43862 = ~n43392 & ~n43861;
  assign n43863 = n43305 & ~n43862;
  assign n43864 = ~n43318 & n43859;
  assign n43865 = ~n43863 & ~n43864;
  assign n43866 = ~n43860 & n43865;
  assign n43867 = ~n43354 & ~n43866;
  assign n43868 = ~n43858 & ~n43867;
  assign n43869 = n43305 & n43379;
  assign n43870 = ~n43305 & ~n43856;
  assign n43871 = ~n43869 & ~n43870;
  assign n43872 = ~n43305 & ~n43843;
  assign n43873 = ~n43379 & ~n43872;
  assign n43874 = ~n43354 & ~n43873;
  assign n43875 = n43871 & ~n43874;
  assign n43876 = n43868 & n43875;
  assign n43877 = pi1085 & ~n43876;
  assign n43878 = ~pi1085 & n43875;
  assign n43879 = ~n43867 & n43878;
  assign n43880 = ~n43858 & n43879;
  assign po1056 = n43877 | n43880;
  assign n43882 = n43305 & n43333;
  assign n43883 = n43361 & ~n43846;
  assign n43884 = ~n43337 & ~n43635;
  assign n43885 = ~n43883 & n43884;
  assign n43886 = ~n43305 & ~n43885;
  assign n43887 = ~n43311 & n43377;
  assign n43888 = ~n43886 & ~n43887;
  assign n43889 = ~n43318 & n43336;
  assign n43890 = n43311 & n43639;
  assign n43891 = ~n43889 & ~n43890;
  assign n43892 = ~n43849 & n43891;
  assign n43893 = n43305 & ~n43892;
  assign n43894 = n43888 & ~n43893;
  assign n43895 = n43354 & ~n43894;
  assign n43896 = ~n43882 & ~n43895;
  assign n43897 = n43311 & n43334;
  assign n43898 = ~n43634 & ~n43897;
  assign n43899 = n43305 & ~n43898;
  assign n43900 = ~n43338 & ~n43899;
  assign n43901 = ~n43333 & ~n43392;
  assign n43902 = ~n43311 & n43396;
  assign n43903 = ~n43639 & ~n43902;
  assign n43904 = ~n43889 & n43903;
  assign n43905 = ~n43305 & ~n43904;
  assign n43906 = n43311 & n43377;
  assign n43907 = ~n43905 & ~n43906;
  assign n43908 = n43901 & n43907;
  assign n43909 = n43900 & n43908;
  assign n43910 = ~n43354 & ~n43909;
  assign n43911 = ~n43369 & ~n43845;
  assign n43912 = ~n43305 & ~n43911;
  assign n43913 = ~n43910 & ~n43912;
  assign n43914 = n43896 & n43913;
  assign n43915 = pi1068 & n43914;
  assign n43916 = ~pi1068 & ~n43914;
  assign po1057 = n43915 | n43916;
  assign n43918 = pi3974 & pi9040;
  assign n43919 = pi4005 & ~pi9040;
  assign n43920 = ~n43918 & ~n43919;
  assign n43921 = pi1104 & n43920;
  assign n43922 = ~pi1104 & ~n43920;
  assign n43923 = ~n43921 & ~n43922;
  assign n43924 = pi3996 & pi9040;
  assign n43925 = pi4012 & ~pi9040;
  assign n43926 = ~n43924 & ~n43925;
  assign n43927 = ~pi1133 & n43926;
  assign n43928 = pi1133 & ~n43926;
  assign n43929 = ~n43927 & ~n43928;
  assign n43930 = pi3977 & pi9040;
  assign n43931 = pi3992 & ~pi9040;
  assign n43932 = ~n43930 & ~n43931;
  assign n43933 = pi1073 & n43932;
  assign n43934 = ~pi1073 & ~n43932;
  assign n43935 = ~n43933 & ~n43934;
  assign n43936 = pi4009 & pi9040;
  assign n43937 = pi3991 & ~pi9040;
  assign n43938 = ~n43936 & ~n43937;
  assign n43939 = ~pi1116 & ~n43938;
  assign n43940 = pi1116 & ~n43936;
  assign n43941 = ~n43937 & n43940;
  assign n43942 = ~n43939 & ~n43941;
  assign n43943 = pi4006 & pi9040;
  assign n43944 = pi3999 & ~pi9040;
  assign n43945 = ~n43943 & ~n43944;
  assign n43946 = ~pi1083 & n43945;
  assign n43947 = pi1083 & ~n43945;
  assign n43948 = ~n43946 & ~n43947;
  assign n43949 = ~n43942 & n43948;
  assign n43950 = n43935 & n43949;
  assign n43951 = ~n43929 & n43950;
  assign n43952 = n43942 & n43948;
  assign n43953 = ~n43935 & n43952;
  assign n43954 = ~n43929 & n43953;
  assign n43955 = ~n43951 & ~n43954;
  assign n43956 = n43942 & ~n43948;
  assign n43957 = ~n43935 & n43956;
  assign n43958 = n43929 & n43957;
  assign n43959 = ~n43935 & n43949;
  assign n43960 = n43929 & n43959;
  assign n43961 = ~n43958 & ~n43960;
  assign n43962 = n43955 & n43961;
  assign n43963 = n43923 & ~n43962;
  assign n43964 = ~n43929 & ~n43935;
  assign n43965 = ~n43948 & n43964;
  assign n43966 = ~n43942 & n43965;
  assign n43967 = ~n43953 & ~n43966;
  assign n43968 = n43923 & ~n43967;
  assign n43969 = n43929 & ~n43948;
  assign n43970 = ~n43923 & n43969;
  assign n43971 = n43935 & n43942;
  assign n43972 = ~n43929 & n43949;
  assign n43973 = ~n43971 & ~n43972;
  assign n43974 = ~n43923 & ~n43973;
  assign n43975 = ~n43970 & ~n43974;
  assign n43976 = ~n43942 & ~n43948;
  assign n43977 = n43935 & n43976;
  assign n43978 = n43929 & n43977;
  assign n43979 = n43975 & ~n43978;
  assign n43980 = ~n43948 & n43971;
  assign n43981 = ~n43929 & n43980;
  assign n43982 = n43979 & ~n43981;
  assign n43983 = ~n43968 & n43982;
  assign n43984 = ~pi3988 & ~pi9040;
  assign n43985 = ~pi3973 & pi9040;
  assign n43986 = ~n43984 & ~n43985;
  assign n43987 = ~pi1102 & n43986;
  assign n43988 = pi1102 & ~n43986;
  assign n43989 = ~n43987 & ~n43988;
  assign n43990 = ~n43983 & ~n43989;
  assign n43991 = ~n43935 & ~n43948;
  assign n43992 = ~n43923 & ~n43929;
  assign n43993 = n43989 & n43992;
  assign n43994 = n43991 & n43993;
  assign n43995 = n43929 & ~n43935;
  assign n43996 = n43948 & n43995;
  assign n43997 = ~n43923 & ~n43996;
  assign n43998 = ~n43929 & n43935;
  assign n43999 = ~n43942 & n43998;
  assign n44000 = ~n43956 & ~n43991;
  assign n44001 = n43929 & ~n44000;
  assign n44002 = n43923 & ~n43950;
  assign n44003 = ~n44001 & n44002;
  assign n44004 = ~n43999 & n44003;
  assign n44005 = ~n43997 & ~n44004;
  assign n44006 = n43935 & n43952;
  assign n44007 = ~n43929 & n44006;
  assign n44008 = ~n44005 & ~n44007;
  assign n44009 = n43989 & ~n44008;
  assign n44010 = ~n43994 & ~n44009;
  assign n44011 = ~n43990 & n44010;
  assign n44012 = ~n43963 & n44011;
  assign n44013 = ~n43923 & n43978;
  assign n44014 = n44012 & ~n44013;
  assign n44015 = pi0994 & ~n44014;
  assign n44016 = n44011 & ~n44013;
  assign n44017 = ~pi0994 & n44016;
  assign n44018 = ~n43963 & n44017;
  assign po1075 = n44015 | n44018;
  assign n44020 = pi4019 & pi9040;
  assign n44021 = pi3973 & ~pi9040;
  assign n44022 = ~n44020 & ~n44021;
  assign n44023 = ~pi1109 & n44022;
  assign n44024 = pi1109 & ~n44022;
  assign n44025 = ~n44023 & ~n44024;
  assign n44026 = pi4033 & pi9040;
  assign n44027 = pi3984 & ~pi9040;
  assign n44028 = ~n44026 & ~n44027;
  assign n44029 = pi1117 & n44028;
  assign n44030 = ~pi1117 & ~n44028;
  assign n44031 = ~n44029 & ~n44030;
  assign n44032 = pi4034 & pi9040;
  assign n44033 = pi3996 & ~pi9040;
  assign n44034 = ~n44032 & ~n44033;
  assign n44035 = ~pi1092 & ~n44034;
  assign n44036 = pi1092 & ~n44032;
  assign n44037 = ~n44033 & n44036;
  assign n44038 = ~n44035 & ~n44037;
  assign n44039 = pi3982 & pi9040;
  assign n44040 = pi3981 & ~pi9040;
  assign n44041 = ~n44039 & ~n44040;
  assign n44042 = ~pi1073 & n44041;
  assign n44043 = pi1073 & ~n44041;
  assign n44044 = ~n44042 & ~n44043;
  assign n44045 = pi3994 & pi9040;
  assign n44046 = pi3993 & ~pi9040;
  assign n44047 = ~n44045 & ~n44046;
  assign n44048 = ~pi1103 & n44047;
  assign n44049 = pi1103 & ~n44047;
  assign n44050 = ~n44048 & ~n44049;
  assign n44051 = ~n44044 & n44050;
  assign n44052 = ~n44038 & n44051;
  assign n44053 = n44031 & n44052;
  assign n44054 = n44044 & ~n44050;
  assign n44055 = ~n44038 & n44054;
  assign n44056 = n44044 & n44050;
  assign n44057 = n44038 & n44056;
  assign n44058 = n44031 & n44057;
  assign n44059 = ~n44055 & ~n44058;
  assign n44060 = ~n44053 & n44059;
  assign n44061 = ~n44025 & ~n44060;
  assign n44062 = ~n44038 & n44044;
  assign n44063 = ~n44025 & n44062;
  assign n44064 = ~n44031 & n44063;
  assign n44065 = n44038 & n44050;
  assign n44066 = ~n44031 & n44065;
  assign n44067 = n44038 & ~n44050;
  assign n44068 = n44031 & n44067;
  assign n44069 = ~n44066 & ~n44068;
  assign n44070 = n44025 & ~n44069;
  assign n44071 = ~n44064 & ~n44070;
  assign n44072 = ~n44038 & ~n44044;
  assign n44073 = ~n44031 & n44072;
  assign n44074 = ~n44050 & n44073;
  assign n44075 = n44038 & n44051;
  assign n44076 = ~n44074 & ~n44075;
  assign n44077 = n44025 & ~n44076;
  assign n44078 = ~n44031 & ~n44038;
  assign n44079 = n44044 & n44078;
  assign n44080 = n44050 & n44079;
  assign n44081 = ~n44053 & ~n44080;
  assign n44082 = n44031 & ~n44038;
  assign n44083 = ~n44050 & n44082;
  assign n44084 = ~n44044 & ~n44050;
  assign n44085 = n44038 & n44084;
  assign n44086 = ~n44031 & n44085;
  assign n44087 = ~n44083 & ~n44086;
  assign n44088 = ~n44025 & ~n44087;
  assign n44089 = n44081 & ~n44088;
  assign n44090 = ~n44077 & n44089;
  assign n44091 = pi4020 & pi9040;
  assign n44092 = pi3978 & ~pi9040;
  assign n44093 = ~n44091 & ~n44092;
  assign n44094 = pi1083 & n44093;
  assign n44095 = ~pi1083 & ~n44093;
  assign n44096 = ~n44094 & ~n44095;
  assign n44097 = ~n44090 & n44096;
  assign n44098 = n44025 & ~n44031;
  assign n44099 = n44051 & n44098;
  assign n44100 = n44038 & n44054;
  assign n44101 = n44044 & n44082;
  assign n44102 = n44050 & n44101;
  assign n44103 = ~n44100 & ~n44102;
  assign n44104 = n44031 & n44084;
  assign n44105 = n44103 & ~n44104;
  assign n44106 = n44025 & ~n44105;
  assign n44107 = ~n44099 & ~n44106;
  assign n44108 = n44031 & n44085;
  assign n44109 = ~n44031 & n44075;
  assign n44110 = ~n44038 & ~n44050;
  assign n44111 = ~n44025 & ~n44031;
  assign n44112 = n44110 & n44111;
  assign n44113 = ~n44031 & n44055;
  assign n44114 = ~n44112 & ~n44113;
  assign n44115 = ~n44109 & n44114;
  assign n44116 = ~n44108 & n44115;
  assign n44117 = n44107 & n44116;
  assign n44118 = ~n44096 & ~n44117;
  assign n44119 = ~n44097 & ~n44118;
  assign n44120 = n44071 & n44119;
  assign n44121 = ~n44061 & n44120;
  assign n44122 = ~pi0993 & ~n44121;
  assign n44123 = pi0993 & n44121;
  assign po1083 = n44122 | n44123;
  assign n44125 = pi3998 & pi9040;
  assign n44126 = pi4030 & ~pi9040;
  assign n44127 = ~n44125 & ~n44126;
  assign n44128 = pi1089 & n44127;
  assign n44129 = ~pi1089 & ~n44127;
  assign n44130 = ~n44128 & ~n44129;
  assign n44131 = pi4007 & pi9040;
  assign n44132 = pi4013 & ~pi9040;
  assign n44133 = ~n44131 & ~n44132;
  assign n44134 = ~pi1116 & n44133;
  assign n44135 = pi1116 & ~n44133;
  assign n44136 = ~n44134 & ~n44135;
  assign n44137 = pi4027 & pi9040;
  assign n44138 = pi3983 & ~pi9040;
  assign n44139 = ~n44137 & ~n44138;
  assign n44140 = ~pi1102 & n44139;
  assign n44141 = pi1102 & ~n44139;
  assign n44142 = ~n44140 & ~n44141;
  assign n44143 = pi4008 & pi9040;
  assign n44144 = pi4028 & ~pi9040;
  assign n44145 = ~n44143 & ~n44144;
  assign n44146 = ~pi1074 & n44145;
  assign n44147 = pi1074 & ~n44145;
  assign n44148 = ~n44146 & ~n44147;
  assign n44149 = n44142 & ~n44148;
  assign n44150 = pi4017 & pi9040;
  assign n44151 = pi3985 & ~pi9040;
  assign n44152 = ~n44150 & ~n44151;
  assign n44153 = pi1105 & n44152;
  assign n44154 = ~pi1105 & ~n44152;
  assign n44155 = ~n44153 & ~n44154;
  assign n44156 = pi4014 & pi9040;
  assign n44157 = pi3995 & ~pi9040;
  assign n44158 = ~n44156 & ~n44157;
  assign n44159 = ~pi1150 & n44158;
  assign n44160 = pi1150 & ~n44158;
  assign n44161 = ~n44159 & ~n44160;
  assign n44162 = n44155 & ~n44161;
  assign n44163 = n44149 & n44162;
  assign n44164 = ~n44136 & n44163;
  assign n44165 = ~n44155 & ~n44161;
  assign n44166 = ~n44142 & ~n44148;
  assign n44167 = n44165 & n44166;
  assign n44168 = n44142 & n44148;
  assign n44169 = ~n44136 & n44168;
  assign n44170 = ~n44155 & n44169;
  assign n44171 = ~n44142 & n44148;
  assign n44172 = ~n44136 & n44171;
  assign n44173 = ~n44161 & n44172;
  assign n44174 = n44155 & n44173;
  assign n44175 = ~n44170 & ~n44174;
  assign n44176 = ~n44167 & n44175;
  assign n44177 = ~n44164 & n44176;
  assign n44178 = n44136 & ~n44155;
  assign n44179 = ~n44148 & n44178;
  assign n44180 = ~n44142 & n44179;
  assign n44181 = n44177 & ~n44180;
  assign n44182 = ~n44130 & ~n44181;
  assign n44183 = ~n44136 & ~n44155;
  assign n44184 = n44148 & n44183;
  assign n44185 = ~n44136 & ~n44142;
  assign n44186 = ~n44148 & n44185;
  assign n44187 = n44155 & n44186;
  assign n44188 = ~n44184 & ~n44187;
  assign n44189 = n44136 & n44149;
  assign n44190 = n44155 & n44189;
  assign n44191 = n44188 & ~n44190;
  assign n44192 = n44161 & ~n44191;
  assign n44193 = n44136 & n44148;
  assign n44194 = ~n44142 & n44193;
  assign n44195 = n44161 & n44194;
  assign n44196 = n44155 & n44195;
  assign n44197 = n44142 & n44183;
  assign n44198 = ~n44155 & n44168;
  assign n44199 = ~n44197 & ~n44198;
  assign n44200 = n44161 & ~n44199;
  assign n44201 = ~n44196 & ~n44200;
  assign n44202 = ~n44130 & ~n44201;
  assign n44203 = ~n44192 & ~n44202;
  assign n44204 = ~n44182 & n44203;
  assign n44205 = n44136 & n44155;
  assign n44206 = ~n44161 & n44205;
  assign n44207 = n44168 & n44206;
  assign n44208 = n44136 & ~n44142;
  assign n44209 = n44165 & n44208;
  assign n44210 = n44161 & n44185;
  assign n44211 = n44142 & n44155;
  assign n44212 = n44136 & n44211;
  assign n44213 = ~n44189 & ~n44212;
  assign n44214 = ~n44210 & n44213;
  assign n44215 = ~n44155 & n44194;
  assign n44216 = n44214 & ~n44215;
  assign n44217 = n44136 & ~n44148;
  assign n44218 = n44155 & n44168;
  assign n44219 = ~n44217 & ~n44218;
  assign n44220 = ~n44161 & ~n44219;
  assign n44221 = n44149 & ~n44161;
  assign n44222 = ~n44155 & n44221;
  assign n44223 = ~n44220 & ~n44222;
  assign n44224 = n44216 & n44223;
  assign n44225 = n44130 & ~n44224;
  assign n44226 = ~n44209 & ~n44225;
  assign n44227 = ~n44207 & n44226;
  assign n44228 = n44204 & n44227;
  assign n44229 = pi0992 & n44228;
  assign n44230 = ~pi0992 & ~n44228;
  assign po1084 = n44229 | n44230;
  assign n44232 = pi4027 & ~pi9040;
  assign n44233 = pi3975 & pi9040;
  assign n44234 = ~n44232 & ~n44233;
  assign n44235 = ~pi1110 & ~n44234;
  assign n44236 = pi1110 & n44234;
  assign n44237 = ~n44235 & ~n44236;
  assign n44238 = pi4015 & pi9040;
  assign n44239 = pi3997 & ~pi9040;
  assign n44240 = ~n44238 & ~n44239;
  assign n44241 = ~pi1114 & n44240;
  assign n44242 = pi1114 & ~n44240;
  assign n44243 = ~n44241 & ~n44242;
  assign n44244 = pi4004 & pi9040;
  assign n44245 = pi4035 & ~pi9040;
  assign n44246 = ~n44244 & ~n44245;
  assign n44247 = ~pi1128 & ~n44246;
  assign n44248 = pi1128 & ~n44244;
  assign n44249 = ~n44245 & n44248;
  assign n44250 = ~n44247 & ~n44249;
  assign n44251 = pi3986 & pi9040;
  assign n44252 = pi4007 & ~pi9040;
  assign n44253 = ~n44251 & ~n44252;
  assign n44254 = ~pi1082 & ~n44253;
  assign n44255 = pi1082 & n44253;
  assign n44256 = ~n44254 & ~n44255;
  assign n44257 = pi4030 & pi9040;
  assign n44258 = pi4026 & ~pi9040;
  assign n44259 = ~n44257 & ~n44258;
  assign n44260 = ~pi1095 & n44259;
  assign n44261 = pi1095 & ~n44259;
  assign n44262 = ~n44260 & ~n44261;
  assign n44263 = ~n44256 & ~n44262;
  assign n44264 = n44250 & n44263;
  assign n44265 = ~n44243 & n44264;
  assign n44266 = pi3979 & pi9040;
  assign n44267 = pi4010 & ~pi9040;
  assign n44268 = ~n44266 & ~n44267;
  assign n44269 = ~pi1129 & n44268;
  assign n44270 = pi1129 & ~n44268;
  assign n44271 = ~n44269 & ~n44270;
  assign n44272 = n44256 & ~n44262;
  assign n44273 = ~n44243 & n44272;
  assign n44274 = ~n44250 & n44263;
  assign n44275 = n44243 & n44274;
  assign n44276 = ~n44273 & ~n44275;
  assign n44277 = n44271 & ~n44276;
  assign n44278 = ~n44265 & ~n44277;
  assign n44279 = ~pi1095 & ~n44259;
  assign n44280 = pi1095 & n44259;
  assign n44281 = ~n44279 & ~n44280;
  assign n44282 = ~n44256 & ~n44281;
  assign n44283 = ~n44250 & n44282;
  assign n44284 = ~n44271 & n44283;
  assign n44285 = n44263 & ~n44271;
  assign n44286 = ~n44243 & n44285;
  assign n44287 = ~n44284 & ~n44286;
  assign n44288 = n44278 & n44287;
  assign n44289 = n44256 & ~n44281;
  assign n44290 = n44250 & n44289;
  assign n44291 = ~n44243 & n44290;
  assign n44292 = n44250 & n44282;
  assign n44293 = n44243 & n44292;
  assign n44294 = ~n44291 & ~n44293;
  assign n44295 = n44288 & n44294;
  assign n44296 = n44237 & ~n44295;
  assign n44297 = ~n44237 & n44271;
  assign n44298 = ~n44243 & ~n44250;
  assign n44299 = ~n44256 & n44298;
  assign n44300 = ~n44250 & ~n44281;
  assign n44301 = ~n44299 & ~n44300;
  assign n44302 = n44297 & ~n44301;
  assign n44303 = ~n44250 & n44289;
  assign n44304 = n44271 & n44303;
  assign n44305 = n44243 & n44304;
  assign n44306 = n44250 & n44272;
  assign n44307 = n44243 & n44306;
  assign n44308 = ~n44293 & ~n44307;
  assign n44309 = n44271 & ~n44308;
  assign n44310 = ~n44305 & ~n44309;
  assign n44311 = n44243 & n44256;
  assign n44312 = ~n44250 & n44311;
  assign n44313 = n44243 & n44250;
  assign n44314 = ~n44262 & n44313;
  assign n44315 = ~n44256 & n44314;
  assign n44316 = ~n44312 & ~n44315;
  assign n44317 = ~n44243 & ~n44271;
  assign n44318 = n44250 & n44317;
  assign n44319 = ~n44263 & n44318;
  assign n44320 = ~n44271 & n44290;
  assign n44321 = ~n44319 & ~n44320;
  assign n44322 = n44316 & n44321;
  assign n44323 = ~n44237 & ~n44322;
  assign n44324 = ~n44271 & n44315;
  assign n44325 = ~n44323 & ~n44324;
  assign n44326 = n44310 & n44325;
  assign n44327 = ~n44302 & n44326;
  assign n44328 = ~n44296 & n44327;
  assign n44329 = ~n44250 & n44272;
  assign n44330 = n44243 & ~n44271;
  assign n44331 = n44329 & n44330;
  assign n44332 = n44328 & ~n44331;
  assign n44333 = ~pi1027 & ~n44332;
  assign n44334 = pi1027 & ~n44331;
  assign n44335 = n44327 & n44334;
  assign n44336 = ~n44296 & n44335;
  assign po1088 = n44333 | n44336;
  assign n44338 = n44243 & n44283;
  assign n44339 = ~n44243 & n44303;
  assign n44340 = ~n44338 & ~n44339;
  assign n44341 = ~n44271 & ~n44340;
  assign n44342 = n44271 & n44315;
  assign n44343 = ~n44315 & ~n44320;
  assign n44344 = ~n44256 & n44313;
  assign n44345 = ~n44312 & ~n44344;
  assign n44346 = n44271 & ~n44345;
  assign n44347 = ~n44243 & n44271;
  assign n44348 = n44282 & n44347;
  assign n44349 = ~n44250 & n44348;
  assign n44350 = ~n44243 & n44250;
  assign n44351 = ~n44262 & n44350;
  assign n44352 = n44256 & n44351;
  assign n44353 = ~n44271 & n44274;
  assign n44354 = ~n44352 & ~n44353;
  assign n44355 = ~n44349 & n44354;
  assign n44356 = ~n44346 & n44355;
  assign n44357 = n44343 & n44356;
  assign n44358 = n44237 & ~n44357;
  assign n44359 = n44243 & n44320;
  assign n44360 = ~n44358 & ~n44359;
  assign n44361 = ~n44342 & n44360;
  assign n44362 = ~n44341 & n44361;
  assign n44363 = n44250 & ~n44256;
  assign n44364 = n44317 & n44363;
  assign n44365 = ~n44284 & ~n44364;
  assign n44366 = ~n44271 & n44306;
  assign n44367 = n44243 & n44329;
  assign n44368 = ~n44366 & ~n44367;
  assign n44369 = ~n44243 & n44292;
  assign n44370 = ~n44338 & ~n44369;
  assign n44371 = ~n44243 & n44289;
  assign n44372 = ~n44250 & n44281;
  assign n44373 = ~n44371 & ~n44372;
  assign n44374 = n44271 & ~n44373;
  assign n44375 = n44370 & ~n44374;
  assign n44376 = n44368 & n44375;
  assign n44377 = n44365 & n44376;
  assign n44378 = ~n44237 & ~n44377;
  assign n44379 = n44362 & ~n44378;
  assign n44380 = ~pi1004 & ~n44379;
  assign n44381 = pi1004 & n44362;
  assign n44382 = ~n44378 & n44381;
  assign po1091 = n44380 | n44382;
  assign n44384 = ~n44359 & ~n44364;
  assign n44385 = ~n44303 & ~n44315;
  assign n44386 = ~n44371 & n44385;
  assign n44387 = n44271 & ~n44386;
  assign n44388 = ~n44262 & n44298;
  assign n44389 = ~n44256 & n44388;
  assign n44390 = ~n44352 & ~n44389;
  assign n44391 = ~n44331 & n44390;
  assign n44392 = ~n44271 & n44292;
  assign n44393 = n44391 & ~n44392;
  assign n44394 = ~n44387 & n44393;
  assign n44395 = n44237 & ~n44394;
  assign n44396 = n44243 & n44285;
  assign n44397 = n44256 & n44298;
  assign n44398 = ~n44303 & ~n44397;
  assign n44399 = ~n44271 & ~n44398;
  assign n44400 = ~n44396 & ~n44399;
  assign n44401 = n44243 & n44271;
  assign n44402 = n44272 & n44401;
  assign n44403 = n44271 & n44283;
  assign n44404 = ~n44402 & ~n44403;
  assign n44405 = n44400 & n44404;
  assign n44406 = n44256 & n44313;
  assign n44407 = ~n44338 & ~n44406;
  assign n44408 = ~n44369 & n44407;
  assign n44409 = n44405 & n44408;
  assign n44410 = ~n44237 & ~n44409;
  assign n44411 = ~n44338 & n44390;
  assign n44412 = n44271 & ~n44411;
  assign n44413 = ~n44410 & ~n44412;
  assign n44414 = ~n44395 & n44413;
  assign n44415 = n44384 & n44414;
  assign n44416 = pi1017 & ~n44415;
  assign n44417 = ~pi1017 & n44415;
  assign po1092 = n44416 | n44417;
  assign n44419 = ~n44136 & n44142;
  assign n44420 = ~n44180 & ~n44419;
  assign n44421 = ~n44211 & n44420;
  assign n44422 = ~n44161 & ~n44421;
  assign n44423 = n44155 & n44161;
  assign n44424 = ~n44142 & n44423;
  assign n44425 = ~n44136 & n44155;
  assign n44426 = ~n44148 & n44425;
  assign n44427 = ~n44155 & n44172;
  assign n44428 = ~n44426 & ~n44427;
  assign n44429 = n44136 & n44142;
  assign n44430 = ~n44155 & n44161;
  assign n44431 = n44429 & n44430;
  assign n44432 = n44428 & ~n44431;
  assign n44433 = ~n44424 & n44432;
  assign n44434 = ~n44422 & n44433;
  assign n44435 = n44130 & ~n44434;
  assign n44436 = ~n44136 & n44149;
  assign n44437 = ~n44155 & n44436;
  assign n44438 = n44155 & n44169;
  assign n44439 = ~n44437 & ~n44438;
  assign n44440 = ~n44161 & ~n44439;
  assign n44441 = ~n44435 & ~n44440;
  assign n44442 = n44155 & n44172;
  assign n44443 = ~n44186 & ~n44194;
  assign n44444 = ~n44161 & ~n44443;
  assign n44445 = ~n44442 & ~n44444;
  assign n44446 = ~n44190 & n44445;
  assign n44447 = ~n44130 & ~n44446;
  assign n44448 = ~n44166 & ~n44168;
  assign n44449 = n44136 & ~n44448;
  assign n44450 = ~n44198 & ~n44449;
  assign n44451 = n44161 & ~n44450;
  assign n44452 = ~n44130 & n44451;
  assign n44453 = ~n44447 & ~n44452;
  assign n44454 = n44441 & n44453;
  assign n44455 = pi0996 & ~n44454;
  assign n44456 = ~pi0996 & n44441;
  assign n44457 = n44453 & n44456;
  assign po1093 = n44455 | n44457;
  assign n44459 = ~n44155 & n44189;
  assign n44460 = ~n44427 & ~n44459;
  assign n44461 = n44161 & ~n44460;
  assign n44462 = n44186 & n44423;
  assign n44463 = ~n44461 & ~n44462;
  assign n44464 = ~n44209 & n44463;
  assign n44465 = ~n44136 & ~n44161;
  assign n44466 = n44148 & n44465;
  assign n44467 = n44142 & n44466;
  assign n44468 = ~n44155 & n44467;
  assign n44469 = ~n44161 & n44436;
  assign n44470 = ~n44180 & ~n44207;
  assign n44471 = ~n44174 & n44470;
  assign n44472 = ~n44469 & n44471;
  assign n44473 = n44130 & ~n44472;
  assign n44474 = ~n44142 & n44155;
  assign n44475 = n44136 & n44474;
  assign n44476 = n44148 & n44475;
  assign n44477 = ~n44169 & ~n44476;
  assign n44478 = ~n44189 & n44477;
  assign n44479 = n44161 & ~n44478;
  assign n44480 = n44130 & n44479;
  assign n44481 = n44155 & n44221;
  assign n44482 = ~n44467 & ~n44481;
  assign n44483 = ~n44426 & n44482;
  assign n44484 = n44148 & n44178;
  assign n44485 = n44155 & n44166;
  assign n44486 = ~n44185 & ~n44485;
  assign n44487 = n44161 & ~n44486;
  assign n44488 = ~n44484 & ~n44487;
  assign n44489 = n44483 & n44488;
  assign n44490 = ~n44130 & ~n44489;
  assign n44491 = ~n44480 & ~n44490;
  assign n44492 = ~n44473 & n44491;
  assign n44493 = ~n44468 & n44492;
  assign n44494 = n44464 & n44493;
  assign n44495 = pi0997 & ~n44494;
  assign n44496 = ~pi0997 & n44464;
  assign n44497 = n44493 & n44496;
  assign po1094 = n44495 | n44497;
  assign n44499 = n44155 & ~n44448;
  assign n44500 = n44136 & n44499;
  assign n44501 = n44148 & n44425;
  assign n44502 = ~n44217 & ~n44501;
  assign n44503 = ~n44169 & n44502;
  assign n44504 = ~n44161 & ~n44503;
  assign n44505 = ~n44193 & ~n44436;
  assign n44506 = n44161 & ~n44505;
  assign n44507 = ~n44504 & ~n44506;
  assign n44508 = ~n44500 & n44507;
  assign n44509 = ~n44155 & n44186;
  assign n44510 = n44508 & ~n44509;
  assign n44511 = ~n44130 & ~n44510;
  assign n44512 = n44165 & ~n44505;
  assign n44513 = ~n44189 & ~n44194;
  assign n44514 = ~n44169 & ~n44186;
  assign n44515 = n44513 & n44514;
  assign n44516 = n44155 & ~n44515;
  assign n44517 = ~n44512 & ~n44516;
  assign n44518 = ~n44427 & n44517;
  assign n44519 = n44130 & ~n44518;
  assign n44520 = ~n44511 & ~n44519;
  assign n44521 = n44155 & n44436;
  assign n44522 = ~n44509 & ~n44521;
  assign n44523 = n44161 & ~n44522;
  assign n44524 = n44520 & ~n44523;
  assign n44525 = pi0998 & ~n44524;
  assign n44526 = ~pi0998 & ~n44523;
  assign n44527 = ~n44519 & n44526;
  assign n44528 = ~n44511 & n44527;
  assign po1097 = n44525 | n44528;
  assign n44530 = ~n44050 & n44101;
  assign n44531 = ~n44067 & ~n44080;
  assign n44532 = ~n44025 & ~n44531;
  assign n44533 = ~n44530 & ~n44532;
  assign n44534 = ~n44074 & n44533;
  assign n44535 = n44025 & n44031;
  assign n44536 = n44052 & n44535;
  assign n44537 = ~n44109 & ~n44536;
  assign n44538 = ~n44058 & n44537;
  assign n44539 = n44534 & n44538;
  assign n44540 = n44096 & ~n44539;
  assign n44541 = ~n44038 & n44084;
  assign n44542 = n44031 & n44541;
  assign n44543 = ~n44102 & ~n44542;
  assign n44544 = ~n44025 & n44052;
  assign n44545 = n44031 & n44075;
  assign n44546 = ~n44544 & ~n44545;
  assign n44547 = n44038 & ~n44044;
  assign n44548 = n44031 & ~n44050;
  assign n44549 = ~n44547 & ~n44548;
  assign n44550 = ~n44062 & n44549;
  assign n44551 = n44025 & ~n44550;
  assign n44552 = ~n44031 & n44057;
  assign n44553 = ~n44113 & ~n44552;
  assign n44554 = ~n44551 & n44553;
  assign n44555 = n44546 & n44554;
  assign n44556 = n44543 & n44555;
  assign n44557 = ~n44096 & ~n44556;
  assign n44558 = ~n44540 & ~n44557;
  assign n44559 = pi1005 & ~n44558;
  assign n44560 = ~pi1005 & ~n44540;
  assign n44561 = ~n44557 & n44560;
  assign po1098 = n44559 | n44561;
  assign n44563 = ~n43935 & n43942;
  assign n44564 = ~n43923 & n44563;
  assign n44565 = ~n43929 & n44564;
  assign n44566 = n43942 & n43965;
  assign n44567 = n43935 & ~n43948;
  assign n44568 = n43929 & n44567;
  assign n44569 = ~n43951 & ~n44568;
  assign n44570 = ~n44566 & n44569;
  assign n44571 = ~n44565 & n44570;
  assign n44572 = n43923 & n43959;
  assign n44573 = n44571 & ~n44572;
  assign n44574 = n43989 & ~n44573;
  assign n44575 = n43929 & n43953;
  assign n44576 = ~n44007 & ~n44575;
  assign n44577 = n43923 & ~n44576;
  assign n44578 = ~n43989 & n43991;
  assign n44579 = ~n43923 & n44578;
  assign n44580 = n43929 & n43935;
  assign n44581 = ~n43942 & n44580;
  assign n44582 = ~n44567 & ~n44581;
  assign n44583 = ~n43953 & n44582;
  assign n44584 = n43923 & ~n44583;
  assign n44585 = ~n43935 & n43976;
  assign n44586 = n43929 & n44585;
  assign n44587 = ~n44584 & ~n44586;
  assign n44588 = ~n43989 & ~n44587;
  assign n44589 = ~n44579 & ~n44588;
  assign n44590 = ~n44577 & n44589;
  assign n44591 = ~n43951 & ~n43960;
  assign n44592 = ~n43929 & ~n43948;
  assign n44593 = ~n43935 & n44592;
  assign n44594 = n43929 & n44006;
  assign n44595 = ~n44593 & ~n44594;
  assign n44596 = n44591 & n44595;
  assign n44597 = ~n43923 & ~n44596;
  assign n44598 = n44590 & ~n44597;
  assign n44599 = ~n44574 & n44598;
  assign n44600 = ~pi1001 & ~n44599;
  assign n44601 = pi1001 & n44590;
  assign n44602 = ~n44574 & n44601;
  assign n44603 = ~n44597 & n44602;
  assign po1099 = n44600 | n44603;
  assign n44605 = pi4020 & ~pi9040;
  assign n44606 = pi3991 & pi9040;
  assign n44607 = ~n44605 & ~n44606;
  assign n44608 = ~pi1103 & ~n44607;
  assign n44609 = pi1103 & n44607;
  assign n44610 = ~n44608 & ~n44609;
  assign n44611 = pi3993 & pi9040;
  assign n44612 = pi4006 & ~pi9040;
  assign n44613 = ~n44611 & ~n44612;
  assign n44614 = ~pi1136 & n44613;
  assign n44615 = pi1136 & ~n44613;
  assign n44616 = ~n44614 & ~n44615;
  assign n44617 = pi3984 & pi9040;
  assign n44618 = pi4032 & ~pi9040;
  assign n44619 = ~n44617 & ~n44618;
  assign n44620 = pi1098 & n44619;
  assign n44621 = ~pi1098 & ~n44619;
  assign n44622 = ~n44620 & ~n44621;
  assign n44623 = pi3990 & pi9040;
  assign n44624 = pi4034 & ~pi9040;
  assign n44625 = ~n44623 & ~n44624;
  assign n44626 = ~pi1092 & ~n44625;
  assign n44627 = pi1092 & ~n44623;
  assign n44628 = ~n44624 & n44627;
  assign n44629 = ~n44626 & ~n44628;
  assign n44630 = pi3988 & pi9040;
  assign n44631 = pi4031 & ~pi9040;
  assign n44632 = ~n44630 & ~n44631;
  assign n44633 = pi1080 & n44632;
  assign n44634 = ~pi1080 & ~n44632;
  assign n44635 = ~n44633 & ~n44634;
  assign n44636 = n44629 & ~n44635;
  assign n44637 = n44622 & n44636;
  assign n44638 = ~n44629 & ~n44635;
  assign n44639 = ~n44622 & n44638;
  assign n44640 = ~n44637 & ~n44639;
  assign n44641 = n44616 & ~n44640;
  assign n44642 = pi4012 & pi9040;
  assign n44643 = pi4002 & ~pi9040;
  assign n44644 = ~n44642 & ~n44643;
  assign n44645 = ~pi1111 & n44644;
  assign n44646 = pi1111 & ~n44644;
  assign n44647 = ~n44645 & ~n44646;
  assign n44648 = n44629 & n44635;
  assign n44649 = n44622 & n44648;
  assign n44650 = ~n44647 & n44649;
  assign n44651 = ~n44641 & ~n44650;
  assign n44652 = ~n44622 & n44635;
  assign n44653 = n44635 & ~n44647;
  assign n44654 = ~n44652 & ~n44653;
  assign n44655 = n44622 & n44638;
  assign n44656 = n44654 & ~n44655;
  assign n44657 = ~n44616 & ~n44656;
  assign n44658 = n44651 & ~n44657;
  assign n44659 = ~n44610 & ~n44658;
  assign n44660 = n44629 & n44652;
  assign n44661 = n44647 & n44660;
  assign n44662 = n44616 & n44661;
  assign n44663 = ~n44629 & n44635;
  assign n44664 = n44616 & n44647;
  assign n44665 = n44663 & n44664;
  assign n44666 = n44622 & n44665;
  assign n44667 = ~n44662 & ~n44666;
  assign n44668 = ~n44622 & n44647;
  assign n44669 = n44629 & n44668;
  assign n44670 = ~n44635 & n44669;
  assign n44671 = ~n44616 & n44670;
  assign n44672 = n44667 & ~n44671;
  assign n44673 = ~n44622 & n44636;
  assign n44674 = ~n44616 & n44673;
  assign n44675 = n44622 & n44647;
  assign n44676 = ~n44629 & n44675;
  assign n44677 = ~n44670 & ~n44676;
  assign n44678 = ~n44616 & n44635;
  assign n44679 = n44675 & n44678;
  assign n44680 = n44637 & ~n44647;
  assign n44681 = n44616 & n44652;
  assign n44682 = ~n44680 & ~n44681;
  assign n44683 = n44639 & ~n44647;
  assign n44684 = n44682 & ~n44683;
  assign n44685 = ~n44679 & n44684;
  assign n44686 = n44677 & n44685;
  assign n44687 = ~n44674 & n44686;
  assign n44688 = n44610 & ~n44687;
  assign n44689 = n44672 & ~n44688;
  assign n44690 = ~n44659 & n44689;
  assign n44691 = ~pi1006 & ~n44690;
  assign n44692 = pi1006 & n44672;
  assign n44693 = ~n44659 & n44692;
  assign n44694 = ~n44688 & n44693;
  assign po1100 = n44691 | n44694;
  assign n44696 = n43929 & n43980;
  assign n44697 = ~n43977 & ~n44593;
  assign n44698 = n43923 & ~n44697;
  assign n44699 = ~n44696 & ~n44698;
  assign n44700 = ~n43923 & n43950;
  assign n44701 = ~n43923 & n43929;
  assign n44702 = ~n43948 & n44701;
  assign n44703 = n43942 & n44702;
  assign n44704 = n43952 & n43992;
  assign n44705 = ~n44703 & ~n44704;
  assign n44706 = ~n44700 & n44705;
  assign n44707 = ~n43960 & ~n43966;
  assign n44708 = n43948 & n43998;
  assign n44709 = n44707 & ~n44708;
  assign n44710 = n44706 & n44709;
  assign n44711 = n44699 & n44710;
  assign n44712 = ~n43989 & ~n44711;
  assign n44713 = ~n43959 & ~n43977;
  assign n44714 = ~n43929 & ~n44713;
  assign n44715 = ~n43929 & n44567;
  assign n44716 = n43942 & n43995;
  assign n44717 = ~n44006 & ~n44716;
  assign n44718 = ~n44715 & n44717;
  assign n44719 = n43923 & ~n44718;
  assign n44720 = n43929 & n43976;
  assign n44721 = ~n44566 & ~n44720;
  assign n44722 = ~n43923 & ~n44721;
  assign n44723 = ~n44575 & ~n44722;
  assign n44724 = ~n44719 & n44723;
  assign n44725 = ~n44714 & n44724;
  assign n44726 = n43989 & ~n44725;
  assign n44727 = n43923 & n43996;
  assign n44728 = ~n44726 & ~n44727;
  assign n44729 = n43971 & n44701;
  assign n44730 = ~n43948 & n44729;
  assign n44731 = n44728 & ~n44730;
  assign n44732 = ~n44712 & n44731;
  assign n44733 = ~pi1002 & ~n44732;
  assign n44734 = pi1002 & n44728;
  assign n44735 = ~n44712 & n44734;
  assign n44736 = ~n44730 & n44735;
  assign po1101 = n44733 | n44736;
  assign n44738 = pi4028 & pi9040;
  assign n44739 = pi4004 & ~pi9040;
  assign n44740 = ~n44738 & ~n44739;
  assign n44741 = pi1121 & n44740;
  assign n44742 = ~pi1121 & ~n44740;
  assign n44743 = ~n44741 & ~n44742;
  assign n44744 = pi4026 & pi9040;
  assign n44745 = pi4000 & ~pi9040;
  assign n44746 = ~n44744 & ~n44745;
  assign n44747 = pi1089 & n44746;
  assign n44748 = ~pi1089 & ~n44746;
  assign n44749 = ~n44747 & ~n44748;
  assign n44750 = pi3976 & pi9040;
  assign n44751 = pi4017 & ~pi9040;
  assign n44752 = ~n44750 & ~n44751;
  assign n44753 = pi1122 & n44752;
  assign n44754 = ~pi1122 & ~n44752;
  assign n44755 = ~n44753 & ~n44754;
  assign n44756 = n44749 & ~n44755;
  assign n44757 = pi3983 & pi9040;
  assign n44758 = pi3986 & ~pi9040;
  assign n44759 = ~n44757 & ~n44758;
  assign n44760 = ~pi1120 & n44759;
  assign n44761 = pi1120 & ~n44759;
  assign n44762 = ~n44760 & ~n44761;
  assign n44763 = pi3997 & pi9040;
  assign n44764 = pi3998 & ~pi9040;
  assign n44765 = ~n44763 & ~n44764;
  assign n44766 = pi1074 & n44765;
  assign n44767 = ~pi1074 & ~n44765;
  assign n44768 = ~n44766 & ~n44767;
  assign n44769 = ~n44762 & n44768;
  assign n44770 = n44756 & n44769;
  assign n44771 = ~n44762 & ~n44768;
  assign n44772 = ~n44749 & n44771;
  assign n44773 = ~n44770 & ~n44772;
  assign n44774 = ~n44743 & ~n44773;
  assign n44775 = pi4010 & pi9040;
  assign n44776 = pi4011 & ~pi9040;
  assign n44777 = ~n44775 & ~n44776;
  assign n44778 = ~pi1099 & ~n44777;
  assign n44779 = pi1099 & n44777;
  assign n44780 = ~n44778 & ~n44779;
  assign n44781 = n44743 & n44762;
  assign n44782 = n44749 & n44781;
  assign n44783 = n44756 & ~n44768;
  assign n44784 = n44749 & n44755;
  assign n44785 = n44768 & n44784;
  assign n44786 = ~n44783 & ~n44785;
  assign n44787 = ~n44749 & ~n44755;
  assign n44788 = n44768 & n44787;
  assign n44789 = ~n44762 & n44788;
  assign n44790 = n44786 & ~n44789;
  assign n44791 = n44743 & ~n44790;
  assign n44792 = ~n44782 & ~n44791;
  assign n44793 = ~n44749 & n44755;
  assign n44794 = ~n44768 & n44793;
  assign n44795 = ~n44762 & n44794;
  assign n44796 = n44792 & ~n44795;
  assign n44797 = n44762 & n44787;
  assign n44798 = ~n44749 & n44768;
  assign n44799 = n44755 & n44798;
  assign n44800 = ~n44797 & ~n44799;
  assign n44801 = ~n44743 & ~n44800;
  assign n44802 = ~n44768 & n44784;
  assign n44803 = n44762 & n44802;
  assign n44804 = ~n44801 & ~n44803;
  assign n44805 = n44796 & n44804;
  assign n44806 = n44780 & ~n44805;
  assign n44807 = ~n44774 & ~n44806;
  assign n44808 = n44743 & ~n44780;
  assign n44809 = ~n44800 & n44808;
  assign n44810 = ~n44768 & n44787;
  assign n44811 = ~n44802 & ~n44810;
  assign n44812 = ~n44762 & ~n44811;
  assign n44813 = ~n44770 & ~n44812;
  assign n44814 = ~n44780 & ~n44813;
  assign n44815 = ~n44809 & ~n44814;
  assign n44816 = ~n44743 & ~n44780;
  assign n44817 = n44756 & n44762;
  assign n44818 = ~n44794 & ~n44817;
  assign n44819 = n44749 & n44768;
  assign n44820 = n44818 & ~n44819;
  assign n44821 = n44816 & ~n44820;
  assign n44822 = n44815 & ~n44821;
  assign n44823 = n44807 & n44822;
  assign n44824 = ~pi1007 & ~n44823;
  assign n44825 = pi1007 & n44815;
  assign n44826 = n44807 & n44825;
  assign n44827 = ~n44821 & n44826;
  assign po1102 = n44824 | n44827;
  assign n44829 = ~n44610 & n44616;
  assign n44830 = n44622 & ~n44635;
  assign n44831 = n44647 & n44830;
  assign n44832 = n44622 & n44663;
  assign n44833 = ~n44647 & n44832;
  assign n44834 = n44647 & n44648;
  assign n44835 = ~n44833 & ~n44834;
  assign n44836 = ~n44831 & n44835;
  assign n44837 = n44829 & ~n44836;
  assign n44838 = ~n44629 & n44668;
  assign n44839 = ~n44647 & n44655;
  assign n44840 = ~n44838 & ~n44839;
  assign n44841 = ~n44622 & n44663;
  assign n44842 = ~n44649 & ~n44841;
  assign n44843 = n44840 & n44842;
  assign n44844 = ~n44616 & ~n44843;
  assign n44845 = ~n44647 & n44673;
  assign n44846 = ~n44844 & ~n44845;
  assign n44847 = ~n44610 & ~n44846;
  assign n44848 = ~n44837 & ~n44847;
  assign n44849 = ~n44616 & n44647;
  assign n44850 = n44622 & n44849;
  assign n44851 = n44629 & n44850;
  assign n44852 = n44647 & n44841;
  assign n44853 = ~n44851 & ~n44852;
  assign n44854 = ~n44638 & ~n44648;
  assign n44855 = ~n44647 & ~n44854;
  assign n44856 = ~n44639 & ~n44855;
  assign n44857 = n44616 & ~n44856;
  assign n44858 = ~n44637 & ~n44831;
  assign n44859 = ~n44833 & n44858;
  assign n44860 = ~n44616 & ~n44859;
  assign n44861 = ~n44857 & ~n44860;
  assign n44862 = ~n44647 & n44660;
  assign n44863 = ~n44683 & ~n44862;
  assign n44864 = ~n44670 & n44863;
  assign n44865 = ~n44665 & n44864;
  assign n44866 = n44861 & n44865;
  assign n44867 = n44610 & ~n44866;
  assign n44868 = n44853 & ~n44867;
  assign n44869 = n44848 & n44868;
  assign n44870 = pi1008 & ~n44869;
  assign n44871 = ~pi1008 & n44853;
  assign n44872 = n44848 & n44871;
  assign n44873 = ~n44867 & n44872;
  assign po1103 = n44870 | n44873;
  assign n44875 = ~n44647 & n44830;
  assign n44876 = ~n44649 & ~n44875;
  assign n44877 = ~n44852 & n44876;
  assign n44878 = ~n44616 & ~n44877;
  assign n44879 = n44629 & n44647;
  assign n44880 = n44652 & n44879;
  assign n44881 = n44637 & n44647;
  assign n44882 = ~n44622 & ~n44635;
  assign n44883 = ~n44663 & ~n44882;
  assign n44884 = ~n44647 & ~n44883;
  assign n44885 = ~n44881 & ~n44884;
  assign n44886 = ~n44880 & n44885;
  assign n44887 = n44616 & ~n44886;
  assign n44888 = ~n44878 & ~n44887;
  assign n44889 = n44610 & ~n44888;
  assign n44890 = n44616 & n44639;
  assign n44891 = n44647 & n44890;
  assign n44892 = ~n44666 & ~n44891;
  assign n44893 = ~n44671 & n44892;
  assign n44894 = ~n44635 & n44849;
  assign n44895 = n44635 & n44675;
  assign n44896 = ~n44875 & ~n44895;
  assign n44897 = n44616 & ~n44896;
  assign n44898 = ~n44665 & ~n44897;
  assign n44899 = n44647 & n44832;
  assign n44900 = ~n44862 & ~n44899;
  assign n44901 = ~n44616 & n44652;
  assign n44902 = ~n44647 & n44901;
  assign n44903 = ~n44674 & ~n44902;
  assign n44904 = n44900 & n44903;
  assign n44905 = n44898 & n44904;
  assign n44906 = ~n44894 & n44905;
  assign n44907 = ~n44610 & ~n44906;
  assign n44908 = n44647 & n44655;
  assign n44909 = ~n44647 & n44648;
  assign n44910 = ~n44908 & ~n44909;
  assign n44911 = ~n44616 & ~n44910;
  assign n44912 = ~n44907 & ~n44911;
  assign n44913 = n44893 & n44912;
  assign n44914 = ~n44889 & n44913;
  assign n44915 = ~pi1000 & n44914;
  assign n44916 = pi1000 & ~n44914;
  assign po1104 = n44915 | n44916;
  assign n44918 = ~n44291 & ~n44299;
  assign n44919 = n44237 & ~n44918;
  assign n44920 = n44281 & n44313;
  assign n44921 = ~n44344 & ~n44920;
  assign n44922 = n44271 & ~n44921;
  assign n44923 = n44264 & n44271;
  assign n44924 = ~n44922 & ~n44923;
  assign n44925 = n44237 & ~n44924;
  assign n44926 = ~n44919 & ~n44925;
  assign n44927 = n44290 & n44347;
  assign n44928 = ~n44349 & ~n44927;
  assign n44929 = ~n44312 & ~n44372;
  assign n44930 = ~n44271 & ~n44929;
  assign n44931 = n44237 & n44930;
  assign n44932 = n44928 & ~n44931;
  assign n44933 = ~n44281 & n44313;
  assign n44934 = n44256 & n44933;
  assign n44935 = n44243 & n44282;
  assign n44936 = ~n44339 & ~n44935;
  assign n44937 = ~n44271 & ~n44936;
  assign n44938 = ~n44315 & ~n44352;
  assign n44939 = n44243 & n44289;
  assign n44940 = ~n44329 & ~n44939;
  assign n44941 = n44271 & ~n44940;
  assign n44942 = n44938 & ~n44941;
  assign n44943 = ~n44937 & n44942;
  assign n44944 = ~n44934 & n44943;
  assign n44945 = ~n44237 & ~n44944;
  assign n44946 = ~n44369 & n44390;
  assign n44947 = ~n44271 & ~n44946;
  assign n44948 = ~n44945 & ~n44947;
  assign n44949 = n44932 & n44948;
  assign n44950 = n44926 & n44949;
  assign n44951 = ~pi1040 & ~n44950;
  assign n44952 = pi1040 & n44932;
  assign n44953 = n44926 & n44952;
  assign n44954 = n44948 & n44953;
  assign po1105 = n44951 | n44954;
  assign n44956 = ~n44743 & ~n44762;
  assign n44957 = ~n44787 & ~n44802;
  assign n44958 = n44956 & ~n44957;
  assign n44959 = ~n44743 & ~n44768;
  assign n44960 = n44787 & n44959;
  assign n44961 = ~n44958 & ~n44960;
  assign n44962 = n44780 & ~n44961;
  assign n44963 = n44762 & n44768;
  assign n44964 = n44755 & n44963;
  assign n44965 = n44749 & n44964;
  assign n44966 = ~n44819 & ~n44963;
  assign n44967 = n44743 & ~n44966;
  assign n44968 = n44762 & ~n44768;
  assign n44969 = ~n44755 & n44968;
  assign n44970 = n44749 & n44969;
  assign n44971 = ~n44967 & ~n44970;
  assign n44972 = ~n44965 & n44971;
  assign n44973 = n44780 & ~n44972;
  assign n44974 = ~n44962 & ~n44973;
  assign n44975 = n44755 & n44769;
  assign n44976 = ~n44749 & n44975;
  assign n44977 = n44762 & n44794;
  assign n44978 = ~n44976 & ~n44977;
  assign n44979 = ~n44743 & ~n44978;
  assign n44980 = ~n44762 & n44810;
  assign n44981 = n44762 & n44819;
  assign n44982 = ~n44980 & ~n44981;
  assign n44983 = n44743 & ~n44982;
  assign n44984 = ~n44756 & ~n44819;
  assign n44985 = ~n44762 & ~n44984;
  assign n44986 = ~n44794 & ~n44985;
  assign n44987 = ~n44743 & ~n44986;
  assign n44988 = n44755 & n44762;
  assign n44989 = ~n44743 & n44988;
  assign n44990 = ~n44768 & n44989;
  assign n44991 = ~n44755 & n44768;
  assign n44992 = ~n44794 & ~n44991;
  assign n44993 = n44762 & ~n44992;
  assign n44994 = n44743 & ~n44762;
  assign n44995 = n44784 & n44994;
  assign n44996 = ~n44768 & n44995;
  assign n44997 = ~n44993 & ~n44996;
  assign n44998 = ~n44990 & n44997;
  assign n44999 = ~n44987 & n44998;
  assign n45000 = ~n44976 & n44999;
  assign n45001 = ~n44780 & ~n45000;
  assign n45002 = ~n44983 & ~n45001;
  assign n45003 = ~n44979 & n45002;
  assign n45004 = n44974 & n45003;
  assign n45005 = pi1020 & n45004;
  assign n45006 = ~pi1020 & ~n45004;
  assign po1106 = n45005 | n45006;
  assign n45008 = ~n44635 & n44647;
  assign n45009 = ~n44676 & ~n45008;
  assign n45010 = n44616 & ~n45009;
  assign n45011 = n44622 & ~n44647;
  assign n45012 = n44629 & n45011;
  assign n45013 = ~n45010 & ~n45012;
  assign n45014 = ~n44616 & n44648;
  assign n45015 = n44647 & n45014;
  assign n45016 = ~n44908 & ~n45015;
  assign n45017 = n45013 & n45016;
  assign n45018 = n44610 & ~n45017;
  assign n45019 = ~n44832 & ~n44862;
  assign n45020 = n44636 & n44647;
  assign n45021 = n45019 & ~n45020;
  assign n45022 = ~n44616 & ~n45021;
  assign n45023 = n44648 & n44664;
  assign n45024 = ~n44852 & ~n45023;
  assign n45025 = ~n45022 & n45024;
  assign n45026 = ~n44655 & ~n44845;
  assign n45027 = n44616 & ~n45026;
  assign n45028 = n45025 & ~n45027;
  assign n45029 = ~n44610 & ~n45028;
  assign n45030 = ~n45018 & ~n45029;
  assign n45031 = ~n44647 & n44842;
  assign n45032 = ~n44638 & n44647;
  assign n45033 = ~n45031 & ~n45032;
  assign n45034 = n44616 & n45033;
  assign n45035 = ~n44616 & ~n44647;
  assign n45036 = n44640 & ~n44832;
  assign n45037 = n45035 & ~n45036;
  assign n45038 = ~n45034 & ~n45037;
  assign n45039 = n45030 & n45038;
  assign n45040 = ~pi1021 & ~n45039;
  assign n45041 = pi1021 & n45038;
  assign n45042 = ~n45029 & n45041;
  assign n45043 = ~n45018 & n45042;
  assign po1107 = n45040 | n45043;
  assign n45045 = ~n44031 & n44084;
  assign n45046 = ~n44552 & ~n45045;
  assign n45047 = ~n44025 & n45046;
  assign n45048 = n44031 & n44065;
  assign n45049 = ~n44051 & ~n44054;
  assign n45050 = n44038 & ~n45049;
  assign n45051 = n44050 & n44078;
  assign n45052 = n44031 & n44054;
  assign n45053 = ~n45051 & ~n45052;
  assign n45054 = ~n45050 & n45053;
  assign n45055 = n44025 & n45054;
  assign n45056 = ~n45048 & n45055;
  assign n45057 = ~n45047 & ~n45056;
  assign n45058 = n44031 & n45050;
  assign n45059 = ~n44542 & ~n45058;
  assign n45060 = ~n45057 & n45059;
  assign n45061 = n44096 & ~n45060;
  assign n45062 = ~n44025 & ~n45049;
  assign n45063 = ~n44031 & n45062;
  assign n45064 = n44031 & n44056;
  assign n45065 = ~n44108 & ~n45064;
  assign n45066 = ~n44025 & ~n45065;
  assign n45067 = ~n44038 & n45062;
  assign n45068 = ~n45066 & ~n45067;
  assign n45069 = ~n45063 & n45068;
  assign n45070 = ~n44096 & ~n45069;
  assign n45071 = ~n45061 & ~n45070;
  assign n45072 = n44025 & ~n45046;
  assign n45073 = ~n44102 & ~n45072;
  assign n45074 = ~n44096 & ~n45073;
  assign n45075 = ~n44025 & n44102;
  assign n45076 = n44025 & ~n45059;
  assign n45077 = ~n45075 & ~n45076;
  assign n45078 = ~n45074 & n45077;
  assign n45079 = n45071 & n45078;
  assign n45080 = pi1012 & ~n45079;
  assign n45081 = ~pi1012 & n45078;
  assign n45082 = ~n45070 & n45081;
  assign n45083 = ~n45061 & n45082;
  assign po1108 = n45080 | n45083;
  assign n45085 = pi3999 & pi9040;
  assign n45086 = pi3990 & ~pi9040;
  assign n45087 = ~n45085 & ~n45086;
  assign n45088 = ~pi1080 & ~n45087;
  assign n45089 = pi1080 & n45087;
  assign n45090 = ~n45088 & ~n45089;
  assign n45091 = pi4031 & pi9040;
  assign n45092 = pi4009 & ~pi9040;
  assign n45093 = ~n45091 & ~n45092;
  assign n45094 = pi1162 & n45093;
  assign n45095 = ~pi1162 & ~n45093;
  assign n45096 = ~n45094 & ~n45095;
  assign n45097 = pi4005 & pi9040;
  assign n45098 = pi4001 & ~pi9040;
  assign n45099 = ~n45097 & ~n45098;
  assign n45100 = ~pi1115 & n45099;
  assign n45101 = pi1115 & ~n45099;
  assign n45102 = ~n45100 & ~n45101;
  assign n45103 = ~n45096 & n45102;
  assign n45104 = pi4032 & pi9040;
  assign n45105 = pi3977 & ~pi9040;
  assign n45106 = ~n45104 & ~n45105;
  assign n45107 = ~pi1110 & ~n45106;
  assign n45108 = pi1110 & ~n45104;
  assign n45109 = ~n45105 & n45108;
  assign n45110 = ~n45107 & ~n45109;
  assign n45111 = n45103 & n45110;
  assign n45112 = pi4002 & pi9040;
  assign n45113 = pi3982 & ~pi9040;
  assign n45114 = ~n45112 & ~n45113;
  assign n45115 = ~pi1095 & n45114;
  assign n45116 = pi1095 & ~n45114;
  assign n45117 = ~n45115 & ~n45116;
  assign n45118 = pi4003 & pi9040;
  assign n45119 = pi4019 & ~pi9040;
  assign n45120 = ~n45118 & ~n45119;
  assign n45121 = pi1098 & n45120;
  assign n45122 = ~pi1098 & ~n45120;
  assign n45123 = ~n45121 & ~n45122;
  assign n45124 = ~n45110 & ~n45123;
  assign n45125 = ~n45117 & n45124;
  assign n45126 = n45096 & n45125;
  assign n45127 = ~n45110 & n45123;
  assign n45128 = n45117 & n45127;
  assign n45129 = n45096 & n45128;
  assign n45130 = ~n45126 & ~n45129;
  assign n45131 = n45110 & n45123;
  assign n45132 = n45117 & n45131;
  assign n45133 = n45117 & n45124;
  assign n45134 = ~n45096 & n45133;
  assign n45135 = ~n45132 & ~n45134;
  assign n45136 = ~n45102 & ~n45135;
  assign n45137 = n45130 & ~n45136;
  assign n45138 = ~n45111 & n45137;
  assign n45139 = n45090 & ~n45138;
  assign n45140 = n45096 & n45110;
  assign n45141 = n45117 & n45140;
  assign n45142 = ~n45123 & n45141;
  assign n45143 = n45102 & n45142;
  assign n45144 = ~n45096 & ~n45102;
  assign n45145 = n45110 & ~n45123;
  assign n45146 = n45117 & n45145;
  assign n45147 = n45144 & n45146;
  assign n45148 = ~n45096 & ~n45117;
  assign n45149 = ~n45110 & n45148;
  assign n45150 = ~n45147 & ~n45149;
  assign n45151 = ~n45117 & n45127;
  assign n45152 = ~n45132 & ~n45151;
  assign n45153 = ~n45096 & n45127;
  assign n45154 = n45152 & ~n45153;
  assign n45155 = n45102 & ~n45154;
  assign n45156 = n45096 & n45133;
  assign n45157 = ~n45117 & ~n45123;
  assign n45158 = n45110 & n45157;
  assign n45159 = n45096 & n45158;
  assign n45160 = ~n45156 & ~n45159;
  assign n45161 = ~n45117 & n45131;
  assign n45162 = ~n45102 & n45161;
  assign n45163 = n45160 & ~n45162;
  assign n45164 = ~n45155 & n45163;
  assign n45165 = n45150 & n45164;
  assign n45166 = ~n45090 & ~n45165;
  assign n45167 = ~n45143 & ~n45166;
  assign n45168 = ~n45139 & n45167;
  assign n45169 = n45144 & n45151;
  assign n45170 = ~n45102 & n45157;
  assign n45171 = n45096 & n45170;
  assign n45172 = ~n45169 & ~n45171;
  assign n45173 = ~n45102 & n45129;
  assign n45174 = n45172 & ~n45173;
  assign n45175 = n45168 & n45174;
  assign n45176 = ~pi1046 & ~n45175;
  assign n45177 = pi1046 & n45174;
  assign n45178 = n45167 & n45177;
  assign n45179 = ~n45139 & n45178;
  assign po1109 = n45176 | n45179;
  assign n45181 = ~n43951 & ~n43958;
  assign n45182 = ~n43923 & ~n45181;
  assign n45183 = ~n44013 & ~n45182;
  assign n45184 = ~n43935 & ~n43942;
  assign n45185 = n43923 & n45184;
  assign n45186 = ~n43929 & n45185;
  assign n45187 = ~n43923 & n43956;
  assign n45188 = ~n43929 & n45187;
  assign n45189 = ~n44700 & ~n45188;
  assign n45190 = n43942 & n44580;
  assign n45191 = ~n43929 & n43976;
  assign n45192 = ~n45190 & ~n45191;
  assign n45193 = ~n45184 & n45192;
  assign n45194 = n43923 & ~n45193;
  assign n45195 = ~n43954 & ~n45194;
  assign n45196 = n45189 & n45195;
  assign n45197 = ~n43989 & ~n45196;
  assign n45198 = ~n45186 & ~n45197;
  assign n45199 = ~n43977 & ~n43996;
  assign n45200 = ~n44006 & n45199;
  assign n45201 = ~n43923 & ~n45200;
  assign n45202 = n43929 & n43950;
  assign n45203 = ~n43980 & ~n45202;
  assign n45204 = n43923 & ~n45203;
  assign n45205 = ~n45201 & ~n45204;
  assign n45206 = ~n44716 & n45205;
  assign n45207 = ~n43966 & ~n44007;
  assign n45208 = n45206 & n45207;
  assign n45209 = n43989 & ~n45208;
  assign n45210 = n45198 & ~n45209;
  assign n45211 = n45183 & n45210;
  assign n45212 = ~pi1014 & ~n45211;
  assign n45213 = pi1014 & n45198;
  assign n45214 = n45183 & n45213;
  assign n45215 = ~n45209 & n45214;
  assign po1111 = n45212 | n45215;
  assign n45217 = ~n45096 & n45157;
  assign n45218 = ~n45110 & n45217;
  assign n45219 = ~n45096 & n45161;
  assign n45220 = ~n45128 & ~n45219;
  assign n45221 = n45096 & n45157;
  assign n45222 = ~n45096 & n45146;
  assign n45223 = ~n45221 & ~n45222;
  assign n45224 = n45220 & n45223;
  assign n45225 = n45102 & ~n45224;
  assign n45226 = n45096 & n45131;
  assign n45227 = ~n45149 & ~n45226;
  assign n45228 = ~n45133 & n45227;
  assign n45229 = ~n45102 & ~n45228;
  assign n45230 = n45096 & n45117;
  assign n45231 = n45123 & n45230;
  assign n45232 = n45110 & n45231;
  assign n45233 = ~n45229 & ~n45232;
  assign n45234 = ~n45225 & n45233;
  assign n45235 = ~n45218 & n45234;
  assign n45236 = ~n45090 & ~n45235;
  assign n45237 = n45096 & n45102;
  assign n45238 = n45161 & n45237;
  assign n45239 = n45102 & n45133;
  assign n45240 = n45102 & n45151;
  assign n45241 = ~n45239 & ~n45240;
  assign n45242 = ~n45096 & ~n45241;
  assign n45243 = ~n45238 & ~n45242;
  assign n45244 = n45096 & n45127;
  assign n45245 = ~n45096 & n45131;
  assign n45246 = ~n45244 & ~n45245;
  assign n45247 = ~n45158 & n45246;
  assign n45248 = ~n45128 & n45247;
  assign n45249 = ~n45102 & ~n45248;
  assign n45250 = ~n45096 & n45132;
  assign n45251 = ~n45249 & ~n45250;
  assign n45252 = ~n45096 & n45158;
  assign n45253 = ~n45142 & ~n45252;
  assign n45254 = n45251 & n45253;
  assign n45255 = n45243 & n45254;
  assign n45256 = n45090 & ~n45255;
  assign n45257 = n45102 & ~n45130;
  assign n45258 = ~n45256 & ~n45257;
  assign n45259 = ~n45156 & ~n45252;
  assign n45260 = ~n45102 & ~n45259;
  assign n45261 = n45258 & ~n45260;
  assign n45262 = ~n45236 & n45261;
  assign n45263 = pi1018 & ~n45262;
  assign n45264 = ~pi1018 & n45262;
  assign po1112 = n45263 | n45264;
  assign n45266 = n45123 & n45148;
  assign n45267 = ~n45132 & ~n45149;
  assign n45268 = n45102 & ~n45267;
  assign n45269 = ~n45266 & ~n45268;
  assign n45270 = ~n45110 & n45117;
  assign n45271 = n45117 & ~n45123;
  assign n45272 = ~n45096 & n45271;
  assign n45273 = n45096 & n45124;
  assign n45274 = ~n45272 & ~n45273;
  assign n45275 = ~n45270 & n45274;
  assign n45276 = ~n45161 & n45275;
  assign n45277 = ~n45102 & ~n45276;
  assign n45278 = n45269 & ~n45277;
  assign n45279 = ~n45159 & n45278;
  assign n45280 = n45090 & ~n45279;
  assign n45281 = ~n45096 & n45128;
  assign n45282 = n45160 & ~n45281;
  assign n45283 = ~n45102 & ~n45282;
  assign n45284 = ~n45280 & ~n45283;
  assign n45285 = n45110 & n45117;
  assign n45286 = n45102 & n45285;
  assign n45287 = n45096 & n45286;
  assign n45288 = n45144 & n45157;
  assign n45289 = n45096 & n45151;
  assign n45290 = ~n45288 & ~n45289;
  assign n45291 = ~n45110 & ~n45117;
  assign n45292 = n45096 & n45291;
  assign n45293 = ~n45146 & ~n45292;
  assign n45294 = n45102 & ~n45293;
  assign n45295 = n45102 & n45270;
  assign n45296 = ~n45096 & n45295;
  assign n45297 = ~n45294 & ~n45296;
  assign n45298 = n45290 & n45297;
  assign n45299 = ~n45090 & ~n45298;
  assign n45300 = ~n45287 & ~n45299;
  assign n45301 = ~n45219 & n45300;
  assign n45302 = n45284 & n45301;
  assign n45303 = ~pi1019 & ~n45302;
  assign n45304 = ~n45219 & ~n45280;
  assign n45305 = ~n45283 & n45304;
  assign n45306 = n45300 & n45305;
  assign n45307 = pi1019 & n45306;
  assign po1113 = n45303 | n45307;
  assign n45309 = ~n44755 & n44771;
  assign n45310 = ~n44802 & ~n45309;
  assign n45311 = ~n44743 & ~n45310;
  assign n45312 = ~n44762 & n44793;
  assign n45313 = ~n44969 & ~n45312;
  assign n45314 = n44743 & ~n45313;
  assign n45315 = n44762 & n44788;
  assign n45316 = ~n44990 & ~n45315;
  assign n45317 = ~n44770 & n45316;
  assign n45318 = ~n45314 & n45317;
  assign n45319 = ~n45311 & n45318;
  assign n45320 = ~n44965 & ~n44976;
  assign n45321 = n45319 & n45320;
  assign n45322 = n44780 & ~n45321;
  assign n45323 = n44756 & n44963;
  assign n45324 = n44811 & ~n45323;
  assign n45325 = n44743 & ~n45324;
  assign n45326 = n44762 & n44799;
  assign n45327 = ~n45325 & ~n45326;
  assign n45328 = n44749 & n44771;
  assign n45329 = ~n44762 & n44784;
  assign n45330 = ~n45328 & ~n45329;
  assign n45331 = n44743 & ~n45330;
  assign n45332 = n44743 & n44793;
  assign n45333 = n44762 & n45332;
  assign n45334 = ~n45331 & ~n45333;
  assign n45335 = n45327 & n45334;
  assign n45336 = ~n44780 & ~n45335;
  assign n45337 = ~n44788 & ~n44795;
  assign n45338 = ~n44970 & n45337;
  assign n45339 = n44816 & ~n45338;
  assign n45340 = ~n45336 & ~n45339;
  assign n45341 = ~n44770 & ~n44965;
  assign n45342 = ~n44743 & ~n45341;
  assign n45343 = n45340 & ~n45342;
  assign n45344 = ~n45322 & n45343;
  assign n45345 = ~pi1010 & n45344;
  assign n45346 = pi1010 & ~n45344;
  assign po1114 = n45345 | n45346;
  assign n45348 = ~n44025 & n44053;
  assign n45349 = n44078 & ~n45049;
  assign n45350 = ~n44057 & ~n45349;
  assign n45351 = ~n44542 & n45350;
  assign n45352 = n44025 & ~n45351;
  assign n45353 = n44031 & n44100;
  assign n45354 = ~n45352 & ~n45353;
  assign n45355 = ~n44038 & n44056;
  assign n45356 = ~n44031 & n44547;
  assign n45357 = ~n45355 & ~n45356;
  assign n45358 = ~n45052 & n45357;
  assign n45359 = ~n44025 & ~n45358;
  assign n45360 = n45354 & ~n45359;
  assign n45361 = n44096 & ~n45360;
  assign n45362 = ~n45348 & ~n45361;
  assign n45363 = ~n44031 & n44054;
  assign n45364 = ~n44541 & ~n45363;
  assign n45365 = ~n44025 & ~n45364;
  assign n45366 = ~n44058 & ~n45365;
  assign n45367 = ~n44053 & ~n44108;
  assign n45368 = n44031 & n44062;
  assign n45369 = ~n44547 & ~n45368;
  assign n45370 = ~n45355 & n45369;
  assign n45371 = n44025 & ~n45370;
  assign n45372 = ~n44031 & n44100;
  assign n45373 = ~n45371 & ~n45372;
  assign n45374 = n45367 & n45373;
  assign n45375 = n45366 & n45374;
  assign n45376 = ~n44096 & ~n45375;
  assign n45377 = ~n44086 & ~n45048;
  assign n45378 = n44025 & ~n45377;
  assign n45379 = ~n45376 & ~n45378;
  assign n45380 = n45362 & n45379;
  assign n45381 = pi1011 & n45380;
  assign n45382 = ~pi1011 & ~n45380;
  assign po1115 = n45381 | n45382;
  assign n45384 = pi3987 & pi9040;
  assign n45385 = pi3979 & ~pi9040;
  assign n45386 = ~n45384 & ~n45385;
  assign n45387 = pi1122 & n45386;
  assign n45388 = ~pi1122 & ~n45386;
  assign n45389 = ~n45387 & ~n45388;
  assign n45390 = pi4035 & pi9040;
  assign n45391 = pi4018 & ~pi9040;
  assign n45392 = ~n45390 & ~n45391;
  assign n45393 = pi1128 & n45392;
  assign n45394 = ~pi1128 & ~n45392;
  assign n45395 = ~n45393 & ~n45394;
  assign n45396 = pi3980 & pi9040;
  assign n45397 = pi4014 & ~pi9040;
  assign n45398 = ~n45396 & ~n45397;
  assign n45399 = ~pi1099 & n45398;
  assign n45400 = pi1099 & ~n45398;
  assign n45401 = ~n45399 & ~n45400;
  assign n45402 = ~n45395 & ~n45401;
  assign n45403 = ~n45389 & n45402;
  assign n45404 = n45395 & ~n45401;
  assign n45405 = n45389 & n45404;
  assign n45406 = ~n45403 & ~n45405;
  assign n45407 = pi3985 & pi9040;
  assign n45408 = pi3975 & ~pi9040;
  assign n45409 = ~n45407 & ~n45408;
  assign n45410 = pi1127 & n45409;
  assign n45411 = ~pi1127 & ~n45409;
  assign n45412 = ~n45410 & ~n45411;
  assign n45413 = n45389 & ~n45412;
  assign n45414 = n45395 & n45413;
  assign n45415 = n45406 & ~n45414;
  assign n45416 = pi4000 & pi9040;
  assign n45417 = pi4008 & ~pi9040;
  assign n45418 = ~n45416 & ~n45417;
  assign n45419 = ~pi1094 & n45418;
  assign n45420 = pi1094 & ~n45418;
  assign n45421 = ~n45419 & ~n45420;
  assign n45422 = pi4016 & pi9040;
  assign n45423 = pi4015 & ~pi9040;
  assign n45424 = ~n45422 & ~n45423;
  assign n45425 = ~pi1082 & n45424;
  assign n45426 = pi1082 & ~n45424;
  assign n45427 = ~n45425 & ~n45426;
  assign n45428 = n45421 & ~n45427;
  assign n45429 = ~n45415 & n45428;
  assign n45430 = ~n45395 & n45401;
  assign n45431 = n45389 & n45430;
  assign n45432 = ~n45427 & n45431;
  assign n45433 = n45412 & n45432;
  assign n45434 = n45389 & n45402;
  assign n45435 = ~n45421 & n45434;
  assign n45436 = ~n45389 & n45395;
  assign n45437 = n45395 & n45401;
  assign n45438 = n45412 & n45437;
  assign n45439 = ~n45436 & ~n45438;
  assign n45440 = ~n45421 & ~n45439;
  assign n45441 = ~n45435 & ~n45440;
  assign n45442 = ~n45427 & ~n45441;
  assign n45443 = ~n45433 & ~n45442;
  assign n45444 = ~n45389 & n45412;
  assign n45445 = n45395 & n45444;
  assign n45446 = ~n45389 & ~n45412;
  assign n45447 = ~n45395 & n45446;
  assign n45448 = n45401 & n45447;
  assign n45449 = ~n45445 & ~n45448;
  assign n45450 = ~n45421 & ~n45449;
  assign n45451 = n45443 & ~n45450;
  assign n45452 = n45412 & n45421;
  assign n45453 = n45437 & n45452;
  assign n45454 = n45389 & n45453;
  assign n45455 = ~n45404 & ~n45430;
  assign n45456 = n45413 & ~n45455;
  assign n45457 = n45403 & ~n45412;
  assign n45458 = ~n45456 & ~n45457;
  assign n45459 = ~n45389 & n45437;
  assign n45460 = n45421 & n45459;
  assign n45461 = ~n45412 & n45460;
  assign n45462 = n45444 & ~n45455;
  assign n45463 = n45412 & n45434;
  assign n45464 = ~n45462 & ~n45463;
  assign n45465 = ~n45461 & n45464;
  assign n45466 = n45458 & n45465;
  assign n45467 = ~n45454 & n45466;
  assign n45468 = ~n45412 & ~n45421;
  assign n45469 = n45389 & n45468;
  assign n45470 = n45401 & n45469;
  assign n45471 = n45467 & ~n45470;
  assign n45472 = n45427 & ~n45471;
  assign n45473 = n45451 & ~n45472;
  assign n45474 = ~n45429 & n45473;
  assign n45475 = ~pi1024 & ~n45474;
  assign n45476 = pi1024 & n45451;
  assign n45477 = ~n45429 & n45476;
  assign n45478 = ~n45472 & n45477;
  assign po1116 = n45475 | n45478;
  assign n45480 = ~n45134 & ~n45252;
  assign n45481 = ~n45232 & n45480;
  assign n45482 = n45102 & ~n45481;
  assign n45483 = ~n45147 & ~n45173;
  assign n45484 = ~n45142 & ~n45240;
  assign n45485 = ~n45125 & ~n45245;
  assign n45486 = ~n45102 & ~n45485;
  assign n45487 = ~n45219 & ~n45486;
  assign n45488 = n45484 & n45487;
  assign n45489 = n45090 & ~n45488;
  assign n45490 = n45117 & n45123;
  assign n45491 = ~n45270 & ~n45490;
  assign n45492 = n45096 & ~n45491;
  assign n45493 = ~n45153 & ~n45158;
  assign n45494 = ~n45102 & ~n45493;
  assign n45495 = n45096 & n45123;
  assign n45496 = ~n45132 & ~n45495;
  assign n45497 = ~n45124 & n45496;
  assign n45498 = n45102 & ~n45497;
  assign n45499 = ~n45494 & ~n45498;
  assign n45500 = ~n45492 & n45499;
  assign n45501 = ~n45090 & ~n45500;
  assign n45502 = ~n45489 & ~n45501;
  assign n45503 = n45483 & n45502;
  assign n45504 = ~n45482 & n45503;
  assign n45505 = ~pi1025 & ~n45504;
  assign n45506 = pi1025 & n45483;
  assign n45507 = ~n45482 & n45506;
  assign n45508 = n45502 & n45507;
  assign po1117 = n45505 | n45508;
  assign n45510 = n45412 & n45430;
  assign n45511 = ~n45389 & n45510;
  assign n45512 = ~n45463 & ~n45511;
  assign n45513 = ~n45421 & ~n45512;
  assign n45514 = ~n45389 & n45404;
  assign n45515 = n45389 & n45437;
  assign n45516 = ~n45514 & ~n45515;
  assign n45517 = ~n45421 & ~n45516;
  assign n45518 = ~n45412 & n45430;
  assign n45519 = ~n45405 & ~n45518;
  assign n45520 = ~n45459 & n45519;
  assign n45521 = n45421 & ~n45520;
  assign n45522 = ~n45517 & ~n45521;
  assign n45523 = ~n45435 & ~n45448;
  assign n45524 = n45522 & n45523;
  assign n45525 = n45427 & ~n45524;
  assign n45526 = n45412 & n45515;
  assign n45527 = n45402 & ~n45412;
  assign n45528 = ~n45510 & ~n45527;
  assign n45529 = n45421 & ~n45528;
  assign n45530 = ~n45526 & ~n45529;
  assign n45531 = n45389 & ~n45421;
  assign n45532 = ~n45395 & n45531;
  assign n45533 = n45401 & n45532;
  assign n45534 = n45406 & ~n45533;
  assign n45535 = ~n45459 & n45534;
  assign n45536 = ~n45412 & ~n45535;
  assign n45537 = n45530 & ~n45536;
  assign n45538 = ~n45427 & ~n45537;
  assign n45539 = ~n45525 & ~n45538;
  assign n45540 = ~n45389 & ~n45401;
  assign n45541 = n45452 & n45540;
  assign n45542 = n45539 & ~n45541;
  assign n45543 = ~n45513 & n45542;
  assign n45544 = ~pi1035 & ~n45543;
  assign n45545 = pi1035 & ~n45513;
  assign n45546 = n45539 & n45545;
  assign n45547 = ~n45541 & n45546;
  assign po1118 = n45544 | n45547;
  assign n45549 = ~n45421 & n45515;
  assign n45550 = ~n45412 & n45549;
  assign n45551 = n45402 & n45468;
  assign n45552 = ~n45389 & n45551;
  assign n45553 = ~n45550 & ~n45552;
  assign n45554 = ~n45457 & ~n45461;
  assign n45555 = ~n45401 & n45412;
  assign n45556 = n45389 & n45555;
  assign n45557 = ~n45438 & ~n45556;
  assign n45558 = ~n45421 & ~n45557;
  assign n45559 = n45421 & ~n45446;
  assign n45560 = ~n45455 & n45559;
  assign n45561 = ~n45389 & ~n45437;
  assign n45562 = ~n45421 & n45561;
  assign n45563 = ~n45412 & n45562;
  assign n45564 = ~n45560 & ~n45563;
  assign n45565 = ~n45558 & n45564;
  assign n45566 = n45554 & n45565;
  assign n45567 = ~n45427 & ~n45566;
  assign n45568 = n45553 & ~n45567;
  assign n45569 = n45405 & n45421;
  assign n45570 = n45412 & n45569;
  assign n45571 = n45421 & n45427;
  assign n45572 = n45446 & ~n45455;
  assign n45573 = ~n45438 & ~n45572;
  assign n45574 = ~n45434 & n45573;
  assign n45575 = n45571 & ~n45574;
  assign n45576 = n45403 & n45412;
  assign n45577 = ~n45389 & n45555;
  assign n45578 = ~n45510 & ~n45577;
  assign n45579 = ~n45412 & n45437;
  assign n45580 = ~n45431 & ~n45579;
  assign n45581 = n45578 & n45580;
  assign n45582 = ~n45421 & ~n45581;
  assign n45583 = ~n45576 & ~n45582;
  assign n45584 = n45427 & ~n45583;
  assign n45585 = ~n45575 & ~n45584;
  assign n45586 = ~n45570 & n45585;
  assign n45587 = n45568 & n45586;
  assign n45588 = pi1036 & ~n45587;
  assign n45589 = ~pi1036 & n45568;
  assign n45590 = n45586 & n45589;
  assign po1119 = n45588 | n45590;
  assign n45592 = ~n45431 & ~n45555;
  assign n45593 = n45428 & ~n45592;
  assign n45594 = n45389 & n45412;
  assign n45595 = ~n45404 & n45594;
  assign n45596 = ~n45427 & n45595;
  assign n45597 = ~n45421 & n45444;
  assign n45598 = n45404 & n45597;
  assign n45599 = n45389 & n45452;
  assign n45600 = ~n45395 & n45599;
  assign n45601 = ~n45598 & ~n45600;
  assign n45602 = ~n45596 & n45601;
  assign n45603 = ~n45510 & ~n45579;
  assign n45604 = ~n45421 & ~n45603;
  assign n45605 = ~n45552 & ~n45604;
  assign n45606 = ~n45427 & ~n45605;
  assign n45607 = ~n45404 & ~n45540;
  assign n45608 = ~n45412 & ~n45607;
  assign n45609 = ~n45515 & ~n45608;
  assign n45610 = n45421 & ~n45609;
  assign n45611 = ~n45572 & ~n45610;
  assign n45612 = n45412 & n45459;
  assign n45613 = ~n45395 & n45413;
  assign n45614 = n45412 & ~n45607;
  assign n45615 = ~n45613 & ~n45614;
  assign n45616 = ~n45421 & ~n45615;
  assign n45617 = ~n45612 & ~n45616;
  assign n45618 = n45611 & n45617;
  assign n45619 = n45427 & ~n45618;
  assign n45620 = ~n45606 & ~n45619;
  assign n45621 = n45602 & n45620;
  assign n45622 = ~n45593 & n45621;
  assign n45623 = pi1037 & ~n45622;
  assign n45624 = ~pi1037 & n45602;
  assign n45625 = ~n45593 & n45624;
  assign n45626 = n45620 & n45625;
  assign po1120 = n45623 | n45626;
  assign n45628 = ~n44743 & n44799;
  assign n45629 = n44762 & n44784;
  assign n45630 = ~n44783 & ~n45629;
  assign n45631 = ~n44743 & ~n45630;
  assign n45632 = n44743 & ~n44992;
  assign n45633 = ~n45631 & ~n45632;
  assign n45634 = ~n44980 & n45633;
  assign n45635 = n44780 & ~n45634;
  assign n45636 = ~n45628 & ~n45635;
  assign n45637 = n44768 & n44956;
  assign n45638 = ~n44968 & ~n45637;
  assign n45639 = ~n44749 & ~n45638;
  assign n45640 = ~n44770 & ~n45639;
  assign n45641 = ~n44969 & n45640;
  assign n45642 = ~n44762 & n44802;
  assign n45643 = n44743 & n44785;
  assign n45644 = ~n45642 & ~n45643;
  assign n45645 = n45641 & n45644;
  assign n45646 = ~n44780 & ~n45645;
  assign n45647 = ~n45315 & ~n45329;
  assign n45648 = n44743 & ~n45647;
  assign n45649 = ~n45646 & ~n45648;
  assign n45650 = n45636 & n45649;
  assign n45651 = ~pi1039 & ~n45650;
  assign n45652 = ~n45635 & n45649;
  assign n45653 = pi1039 & n45652;
  assign n45654 = ~n45628 & n45653;
  assign po1121 = n45651 | n45654;
  assign n45656 = pi3937 & pi9040;
  assign n45657 = pi4277 & ~pi9040;
  assign n45658 = ~n45656 & ~n45657;
  assign n45659 = ~pi1146 & ~n45658;
  assign n45660 = pi1146 & n45658;
  assign n45661 = ~n45659 & ~n45660;
  assign n45662 = pi3932 & pi9040;
  assign n45663 = pi3953 & ~pi9040;
  assign n45664 = ~n45662 & ~n45663;
  assign n45665 = ~pi1177 & ~n45664;
  assign n45666 = pi1177 & n45664;
  assign n45667 = ~n45665 & ~n45666;
  assign n45668 = pi4025 & pi9040;
  assign n45669 = pi3954 & ~pi9040;
  assign n45670 = ~n45668 & ~n45669;
  assign n45671 = ~pi1175 & n45670;
  assign n45672 = pi1175 & ~n45670;
  assign n45673 = ~n45671 & ~n45672;
  assign n45674 = pi3934 & pi9040;
  assign n45675 = pi3971 & ~pi9040;
  assign n45676 = ~n45674 & ~n45675;
  assign n45677 = ~pi1131 & ~n45676;
  assign n45678 = pi1131 & n45676;
  assign n45679 = ~n45677 & ~n45678;
  assign n45680 = n45673 & ~n45679;
  assign n45681 = n45667 & n45680;
  assign n45682 = pi4119 & ~pi9040;
  assign n45683 = pi3933 & pi9040;
  assign n45684 = ~n45682 & ~n45683;
  assign n45685 = ~pi1167 & n45684;
  assign n45686 = pi1167 & ~n45684;
  assign n45687 = ~n45685 & ~n45686;
  assign n45688 = pi4210 & pi9040;
  assign n45689 = pi3947 & ~pi9040;
  assign n45690 = ~n45688 & ~n45689;
  assign n45691 = pi1182 & n45690;
  assign n45692 = ~pi1182 & ~n45690;
  assign n45693 = ~n45691 & ~n45692;
  assign n45694 = ~n45687 & ~n45693;
  assign n45695 = n45681 & n45694;
  assign n45696 = ~n45673 & n45687;
  assign n45697 = ~n45667 & n45696;
  assign n45698 = ~n45667 & n45687;
  assign n45699 = ~n45679 & n45698;
  assign n45700 = ~n45697 & ~n45699;
  assign n45701 = ~n45693 & ~n45700;
  assign n45702 = ~n45695 & ~n45701;
  assign n45703 = ~n45661 & ~n45702;
  assign n45704 = ~n45667 & n45679;
  assign n45705 = ~n45687 & n45693;
  assign n45706 = n45704 & n45705;
  assign n45707 = ~n45673 & n45706;
  assign n45708 = n45687 & n45693;
  assign n45709 = n45667 & n45679;
  assign n45710 = n45708 & n45709;
  assign n45711 = ~n45679 & n45696;
  assign n45712 = ~n45667 & n45711;
  assign n45713 = n45667 & ~n45679;
  assign n45714 = ~n45673 & n45713;
  assign n45715 = n45693 & n45714;
  assign n45716 = ~n45687 & n45715;
  assign n45717 = ~n45712 & ~n45716;
  assign n45718 = ~n45710 & n45717;
  assign n45719 = ~n45707 & n45718;
  assign n45720 = n45673 & n45687;
  assign n45721 = n45709 & n45720;
  assign n45722 = n45719 & ~n45721;
  assign n45723 = ~n45661 & ~n45722;
  assign n45724 = ~n45667 & ~n45679;
  assign n45725 = n45673 & ~n45687;
  assign n45726 = n45693 & n45725;
  assign n45727 = n45724 & n45726;
  assign n45728 = n45673 & n45704;
  assign n45729 = ~n45687 & n45728;
  assign n45730 = n45667 & ~n45673;
  assign n45731 = n45679 & n45730;
  assign n45732 = ~n45687 & n45731;
  assign n45733 = ~n45729 & ~n45732;
  assign n45734 = ~n45711 & n45733;
  assign n45735 = ~n45693 & ~n45734;
  assign n45736 = ~n45727 & ~n45735;
  assign n45737 = ~n45723 & n45736;
  assign n45738 = ~n45703 & n45737;
  assign n45739 = n45673 & n45708;
  assign n45740 = n45667 & n45739;
  assign n45741 = ~n45667 & ~n45687;
  assign n45742 = n45673 & n45741;
  assign n45743 = ~n45673 & ~n45693;
  assign n45744 = n45667 & n45743;
  assign n45745 = ~n45742 & ~n45744;
  assign n45746 = ~n45728 & n45745;
  assign n45747 = n45681 & n45687;
  assign n45748 = n45746 & ~n45747;
  assign n45749 = ~n45687 & n45724;
  assign n45750 = n45673 & n45679;
  assign n45751 = ~n45749 & ~n45750;
  assign n45752 = n45693 & ~n45751;
  assign n45753 = n45693 & n45704;
  assign n45754 = n45687 & n45753;
  assign n45755 = ~n45752 & ~n45754;
  assign n45756 = n45748 & n45755;
  assign n45757 = n45661 & ~n45756;
  assign n45758 = ~n45740 & ~n45757;
  assign po1127 = n45738 & n45758;
  assign n45760 = pi3951 & pi9040;
  assign n45761 = pi3966 & ~pi9040;
  assign n45762 = ~n45760 & ~n45761;
  assign n45763 = ~pi1160 & ~n45762;
  assign n45764 = pi1160 & n45762;
  assign n45765 = ~n45763 & ~n45764;
  assign n45766 = pi3955 & pi9040;
  assign n45767 = pi4117 & ~pi9040;
  assign n45768 = ~n45766 & ~n45767;
  assign n45769 = ~pi1166 & ~n45768;
  assign n45770 = pi1166 & n45768;
  assign n45771 = ~n45769 & ~n45770;
  assign n45772 = pi4266 & pi9040;
  assign n45773 = pi4138 & ~pi9040;
  assign n45774 = ~n45772 & ~n45773;
  assign n45775 = ~pi1151 & ~n45774;
  assign n45776 = pi1151 & n45774;
  assign n45777 = ~n45775 & ~n45776;
  assign n45778 = n45771 & n45777;
  assign n45779 = n45765 & n45778;
  assign n45780 = ~n45771 & n45777;
  assign n45781 = ~n45765 & n45780;
  assign n45782 = ~n45779 & ~n45781;
  assign n45783 = pi4132 & pi9040;
  assign n45784 = ~pi4039 & ~pi9040;
  assign n45785 = ~n45783 & ~n45784;
  assign n45786 = pi1163 & n45785;
  assign n45787 = ~pi1163 & ~n45785;
  assign n45788 = ~n45786 & ~n45787;
  assign n45789 = ~n45782 & n45788;
  assign n45790 = pi4043 & pi9040;
  assign n45791 = pi3967 & ~pi9040;
  assign n45792 = ~n45790 & ~n45791;
  assign n45793 = ~pi1130 & ~n45792;
  assign n45794 = pi1130 & n45792;
  assign n45795 = ~n45793 & ~n45794;
  assign n45796 = ~n45771 & n45795;
  assign n45797 = ~n45777 & n45796;
  assign n45798 = n45765 & n45797;
  assign n45799 = n45771 & ~n45795;
  assign n45800 = ~n45777 & n45799;
  assign n45801 = ~n45771 & ~n45795;
  assign n45802 = n45777 & n45801;
  assign n45803 = n45765 & n45802;
  assign n45804 = ~n45800 & ~n45803;
  assign n45805 = ~n45798 & n45804;
  assign n45806 = ~n45788 & ~n45805;
  assign n45807 = ~n45789 & ~n45806;
  assign n45808 = ~n45777 & ~n45795;
  assign n45809 = ~n45788 & n45808;
  assign n45810 = ~n45765 & n45809;
  assign n45811 = n45765 & ~n45777;
  assign n45812 = n45771 & n45811;
  assign n45813 = n45771 & n45795;
  assign n45814 = n45777 & n45813;
  assign n45815 = ~n45765 & n45814;
  assign n45816 = ~n45812 & ~n45815;
  assign n45817 = ~n45788 & ~n45816;
  assign n45818 = ~n45777 & n45813;
  assign n45819 = ~n45765 & n45818;
  assign n45820 = n45777 & n45796;
  assign n45821 = ~n45819 & ~n45820;
  assign n45822 = n45788 & ~n45821;
  assign n45823 = ~n45817 & ~n45822;
  assign n45824 = ~n45765 & ~n45777;
  assign n45825 = ~n45795 & n45824;
  assign n45826 = ~n45771 & n45825;
  assign n45827 = ~n45798 & ~n45826;
  assign n45828 = n45823 & n45827;
  assign n45829 = pi4107 & pi9040;
  assign n45830 = ~pi4022 & ~pi9040;
  assign n45831 = ~n45829 & ~n45830;
  assign n45832 = pi1161 & n45831;
  assign n45833 = ~pi1161 & ~n45831;
  assign n45834 = ~n45832 & ~n45833;
  assign n45835 = ~n45828 & n45834;
  assign n45836 = n45788 & n45796;
  assign n45837 = ~n45765 & n45836;
  assign n45838 = ~n45777 & n45801;
  assign n45839 = n45765 & n45838;
  assign n45840 = n45777 & n45799;
  assign n45841 = ~n45839 & ~n45840;
  assign n45842 = n45765 & n45813;
  assign n45843 = n45841 & ~n45842;
  assign n45844 = n45788 & ~n45843;
  assign n45845 = n45771 & ~n45777;
  assign n45846 = ~n45765 & ~n45788;
  assign n45847 = n45845 & n45846;
  assign n45848 = ~n45765 & n45800;
  assign n45849 = ~n45847 & ~n45848;
  assign n45850 = ~n45844 & n45849;
  assign n45851 = ~n45837 & n45850;
  assign n45852 = ~n45765 & n45820;
  assign n45853 = n45765 & n45814;
  assign n45854 = ~n45852 & ~n45853;
  assign n45855 = n45851 & n45854;
  assign n45856 = ~n45834 & ~n45855;
  assign n45857 = ~n45835 & ~n45856;
  assign n45858 = ~n45810 & n45857;
  assign po1132 = n45807 & n45858;
  assign n45860 = pi3963 & ~pi9040;
  assign n45861 = pi3970 & pi9040;
  assign n45862 = ~n45860 & ~n45861;
  assign n45863 = pi1161 & n45862;
  assign n45864 = ~pi1161 & ~n45862;
  assign n45865 = ~n45863 & ~n45864;
  assign n45866 = pi3949 & pi9040;
  assign n45867 = pi3950 & ~pi9040;
  assign n45868 = ~n45866 & ~n45867;
  assign n45869 = pi1130 & n45868;
  assign n45870 = ~pi1130 & ~n45868;
  assign n45871 = ~n45869 & ~n45870;
  assign n45872 = n45865 & ~n45871;
  assign n45873 = ~pi4130 & ~pi9040;
  assign n45874 = pi4039 & pi9040;
  assign n45875 = ~n45873 & ~n45874;
  assign n45876 = ~pi1177 & n45875;
  assign n45877 = pi1177 & ~n45875;
  assign n45878 = ~n45876 & ~n45877;
  assign n45879 = pi4138 & pi9040;
  assign n45880 = pi4041 & ~pi9040;
  assign n45881 = ~n45879 & ~n45880;
  assign n45882 = pi1172 & n45881;
  assign n45883 = ~pi1172 & ~n45881;
  assign n45884 = ~n45882 & ~n45883;
  assign n45885 = pi4118 & ~pi9040;
  assign n45886 = pi3946 & pi9040;
  assign n45887 = ~n45885 & ~n45886;
  assign n45888 = pi1153 & n45887;
  assign n45889 = ~pi1153 & ~n45887;
  assign n45890 = ~n45888 & ~n45889;
  assign n45891 = n45884 & n45890;
  assign n45892 = n45878 & n45891;
  assign n45893 = n45872 & n45892;
  assign n45894 = pi3968 & pi9040;
  assign n45895 = pi3969 & ~pi9040;
  assign n45896 = ~n45894 & ~n45895;
  assign n45897 = ~pi1175 & n45896;
  assign n45898 = pi1175 & ~n45896;
  assign n45899 = ~n45897 & ~n45898;
  assign n45900 = ~n45865 & n45899;
  assign n45901 = n45871 & n45900;
  assign n45902 = n45865 & ~n45899;
  assign n45903 = ~n45872 & ~n45902;
  assign n45904 = ~n45884 & ~n45903;
  assign n45905 = n45871 & n45884;
  assign n45906 = n45899 & n45905;
  assign n45907 = ~n45904 & ~n45906;
  assign n45908 = ~n45901 & n45907;
  assign n45909 = ~n45890 & n45908;
  assign n45910 = ~n45871 & ~n45884;
  assign n45911 = ~n45865 & n45910;
  assign n45912 = n45890 & ~n45911;
  assign n45913 = ~n45909 & ~n45912;
  assign n45914 = ~n45865 & ~n45899;
  assign n45915 = n45871 & n45914;
  assign n45916 = n45884 & n45915;
  assign n45917 = ~n45913 & ~n45916;
  assign n45918 = n45878 & ~n45917;
  assign n45919 = ~n45871 & n45914;
  assign n45920 = n45884 & n45919;
  assign n45921 = n45884 & n45901;
  assign n45922 = ~n45871 & n45900;
  assign n45923 = ~n45884 & n45922;
  assign n45924 = ~n45921 & ~n45923;
  assign n45925 = ~n45920 & n45924;
  assign n45926 = ~n45871 & n45902;
  assign n45927 = ~n45884 & n45926;
  assign n45928 = n45925 & ~n45927;
  assign n45929 = ~n45890 & ~n45928;
  assign n45930 = n45865 & ~n45884;
  assign n45931 = n45890 & n45930;
  assign n45932 = n45884 & n45900;
  assign n45933 = n45871 & ~n45899;
  assign n45934 = ~n45932 & ~n45933;
  assign n45935 = n45890 & ~n45934;
  assign n45936 = n45865 & n45899;
  assign n45937 = ~n45871 & n45936;
  assign n45938 = n45884 & n45937;
  assign n45939 = ~n45919 & ~n45938;
  assign n45940 = ~n45890 & ~n45939;
  assign n45941 = n45871 & n45902;
  assign n45942 = n45884 & n45941;
  assign n45943 = ~n45940 & ~n45942;
  assign n45944 = n45871 & n45936;
  assign n45945 = ~n45884 & n45944;
  assign n45946 = n45943 & ~n45945;
  assign n45947 = ~n45935 & n45946;
  assign n45948 = ~n45931 & n45947;
  assign n45949 = ~n45878 & ~n45948;
  assign n45950 = ~n45929 & ~n45949;
  assign n45951 = n45890 & n45945;
  assign n45952 = n45950 & ~n45951;
  assign n45953 = ~n45918 & n45952;
  assign po1138 = n45893 | ~n45953;
  assign n45955 = ~n45667 & n45673;
  assign n45956 = ~n45693 & n45955;
  assign n45957 = n45687 & n45956;
  assign n45958 = ~n45673 & ~n45687;
  assign n45959 = n45679 & n45958;
  assign n45960 = n45687 & n45714;
  assign n45961 = ~n45959 & ~n45960;
  assign n45962 = n45667 & n45694;
  assign n45963 = ~n45667 & ~n45673;
  assign n45964 = ~n45741 & ~n45963;
  assign n45965 = ~n45721 & n45964;
  assign n45966 = n45693 & ~n45965;
  assign n45967 = ~n45962 & ~n45966;
  assign n45968 = n45961 & n45967;
  assign n45969 = ~n45957 & n45968;
  assign n45970 = n45661 & ~n45969;
  assign n45971 = ~n45673 & n45704;
  assign n45972 = n45687 & n45971;
  assign n45973 = ~n45673 & n45724;
  assign n45974 = ~n45687 & n45973;
  assign n45975 = ~n45972 & ~n45974;
  assign n45976 = n45693 & ~n45975;
  assign n45977 = ~n45970 & ~n45976;
  assign n45978 = ~n45681 & ~n45731;
  assign n45979 = n45693 & ~n45978;
  assign n45980 = ~n45729 & ~n45979;
  assign n45981 = ~n45687 & n45714;
  assign n45982 = n45980 & ~n45981;
  assign n45983 = ~n45661 & ~n45982;
  assign n45984 = ~n45709 & ~n45724;
  assign n45985 = n45673 & ~n45984;
  assign n45986 = ~n45699 & ~n45985;
  assign n45987 = ~n45693 & ~n45986;
  assign n45988 = ~n45661 & n45987;
  assign n45989 = ~n45983 & ~n45988;
  assign po1146 = ~n45977 | ~n45989;
  assign n45991 = n45680 & n45687;
  assign n45992 = ~n45687 & n45709;
  assign n45993 = ~n45730 & ~n45992;
  assign n45994 = ~n45693 & ~n45993;
  assign n45995 = n45693 & n45973;
  assign n45996 = ~n45687 & n45753;
  assign n45997 = ~n45959 & ~n45996;
  assign n45998 = ~n45995 & n45997;
  assign n45999 = ~n45994 & n45998;
  assign n46000 = ~n45991 & n45999;
  assign n46001 = ~n45661 & ~n46000;
  assign n46002 = n45694 & n45731;
  assign n46003 = n45687 & n45728;
  assign n46004 = ~n45960 & ~n46003;
  assign n46005 = ~n45693 & ~n46004;
  assign n46006 = ~n46002 & ~n46005;
  assign n46007 = ~n45740 & n46006;
  assign n46008 = n45661 & ~n45693;
  assign n46009 = n45681 & ~n45687;
  assign n46010 = ~n45728 & ~n46009;
  assign n46011 = ~n45973 & n46010;
  assign n46012 = n46008 & ~n46011;
  assign n46013 = ~n45721 & ~n45727;
  assign n46014 = n45693 & n45971;
  assign n46015 = ~n45716 & ~n46014;
  assign n46016 = n46013 & n46015;
  assign n46017 = n45661 & ~n46016;
  assign n46018 = ~n46012 & ~n46017;
  assign n46019 = n45687 & n45995;
  assign n46020 = n46018 & ~n46019;
  assign n46021 = n46007 & n46020;
  assign n46022 = ~n46001 & n46021;
  assign n46023 = ~pi1227 & n46022;
  assign n46024 = pi1227 & ~n46022;
  assign po1151 = n46023 | n46024;
  assign n46026 = ~n45728 & ~n45973;
  assign n46027 = ~n45681 & n46026;
  assign n46028 = ~n45731 & n46027;
  assign n46029 = ~n45687 & ~n46028;
  assign n46030 = ~n45960 & ~n46029;
  assign n46031 = ~n45680 & ~n45971;
  assign n46032 = n45708 & ~n46031;
  assign n46033 = n46030 & ~n46032;
  assign n46034 = n45661 & ~n46033;
  assign n46035 = ~n45687 & n45985;
  assign n46036 = ~n45693 & ~n46031;
  assign n46037 = ~n46035 & ~n46036;
  assign n46038 = n45687 & n45731;
  assign n46039 = ~n45679 & n45958;
  assign n46040 = ~n45750 & ~n46039;
  assign n46041 = ~n45973 & n46040;
  assign n46042 = n45693 & ~n46041;
  assign n46043 = ~n46038 & ~n46042;
  assign n46044 = n46037 & n46043;
  assign n46045 = ~n45661 & ~n46044;
  assign n46046 = ~n46034 & ~n46045;
  assign n46047 = ~n45687 & n45971;
  assign n46048 = ~n46038 & ~n46047;
  assign n46049 = ~n45693 & ~n46048;
  assign po1154 = ~n46046 | n46049;
  assign n46051 = pi3969 & pi9040;
  assign n46052 = pi4107 & ~pi9040;
  assign n46053 = ~n46051 & ~n46052;
  assign n46054 = ~pi1166 & ~n46053;
  assign n46055 = pi1166 & n46053;
  assign n46056 = ~n46054 & ~n46055;
  assign n46057 = pi4117 & pi9040;
  assign n46058 = pi3970 & ~pi9040;
  assign n46059 = ~n46057 & ~n46058;
  assign n46060 = pi1181 & n46059;
  assign n46061 = ~pi1181 & ~n46059;
  assign n46062 = ~n46060 & ~n46061;
  assign n46063 = pi3957 & ~pi9040;
  assign n46064 = pi4041 & pi9040;
  assign n46065 = ~n46063 & ~n46064;
  assign n46066 = pi1154 & n46065;
  assign n46067 = ~pi1154 & ~n46065;
  assign n46068 = ~n46066 & ~n46067;
  assign n46069 = pi4023 & ~pi9040;
  assign n46070 = pi4130 & pi9040;
  assign n46071 = ~n46069 & ~n46070;
  assign n46072 = ~pi1155 & n46071;
  assign n46073 = pi1155 & ~n46071;
  assign n46074 = ~n46072 & ~n46073;
  assign n46075 = pi3966 & pi9040;
  assign n46076 = pi3948 & ~pi9040;
  assign n46077 = ~n46075 & ~n46076;
  assign n46078 = pi1169 & n46077;
  assign n46079 = ~pi1169 & ~n46077;
  assign n46080 = ~n46078 & ~n46079;
  assign n46081 = n46074 & n46080;
  assign n46082 = n46068 & n46081;
  assign n46083 = pi4131 & pi9040;
  assign n46084 = pi4266 & ~pi9040;
  assign n46085 = ~n46083 & ~n46084;
  assign n46086 = pi1151 & n46085;
  assign n46087 = ~pi1151 & ~n46085;
  assign n46088 = ~n46086 & ~n46087;
  assign n46089 = ~n46074 & n46088;
  assign n46090 = ~pi1169 & n46077;
  assign n46091 = pi1169 & ~n46077;
  assign n46092 = ~n46090 & ~n46091;
  assign n46093 = n46089 & ~n46092;
  assign n46094 = ~n46082 & ~n46093;
  assign n46095 = ~n46074 & ~n46088;
  assign n46096 = ~n46080 & n46095;
  assign n46097 = ~n46068 & n46096;
  assign n46098 = n46094 & ~n46097;
  assign n46099 = ~n46062 & ~n46098;
  assign n46100 = ~n46074 & ~n46080;
  assign n46101 = n46088 & n46100;
  assign n46102 = ~n46068 & n46101;
  assign n46103 = n46074 & ~n46080;
  assign n46104 = ~n46095 & ~n46103;
  assign n46105 = n46068 & n46104;
  assign n46106 = n46074 & n46088;
  assign n46107 = n46080 & n46106;
  assign n46108 = ~n46068 & ~n46107;
  assign n46109 = ~n46105 & ~n46108;
  assign n46110 = ~n46102 & ~n46109;
  assign n46111 = n46062 & ~n46110;
  assign n46112 = ~n46099 & ~n46111;
  assign n46113 = n46056 & ~n46112;
  assign n46114 = ~n46092 & n46095;
  assign n46115 = ~n46068 & n46114;
  assign n46116 = n46062 & n46115;
  assign n46117 = n46092 & n46106;
  assign n46118 = ~n46068 & n46117;
  assign n46119 = ~n46062 & n46118;
  assign n46120 = n46068 & n46089;
  assign n46121 = n46074 & ~n46088;
  assign n46122 = n46080 & n46121;
  assign n46123 = ~n46068 & n46122;
  assign n46124 = ~n46120 & ~n46123;
  assign n46125 = ~n46062 & ~n46124;
  assign n46126 = ~n46119 & ~n46125;
  assign n46127 = ~n46062 & n46068;
  assign n46128 = n46100 & n46127;
  assign n46129 = ~n46062 & n46117;
  assign n46130 = ~n46128 & ~n46129;
  assign n46131 = n46068 & n46088;
  assign n46132 = ~n46080 & n46131;
  assign n46133 = ~n46074 & n46132;
  assign n46134 = ~n46115 & ~n46133;
  assign n46135 = ~n46068 & ~n46092;
  assign n46136 = ~n46074 & n46135;
  assign n46137 = ~n46082 & ~n46136;
  assign n46138 = n46062 & ~n46137;
  assign n46139 = n46062 & ~n46068;
  assign n46140 = n46095 & n46139;
  assign n46141 = ~n46138 & ~n46140;
  assign n46142 = ~n46062 & ~n46068;
  assign n46143 = n46074 & n46142;
  assign n46144 = n46141 & ~n46143;
  assign n46145 = n46134 & n46144;
  assign n46146 = n46130 & n46145;
  assign n46147 = ~n46056 & ~n46146;
  assign n46148 = n46092 & n46121;
  assign n46149 = n46062 & n46148;
  assign n46150 = ~n46068 & n46149;
  assign n46151 = ~n46147 & ~n46150;
  assign n46152 = n46126 & n46151;
  assign n46153 = ~n46116 & n46152;
  assign po1157 = n46113 | ~n46153;
  assign n46155 = ~n45890 & n45911;
  assign n46156 = ~n45884 & n45919;
  assign n46157 = n45884 & n45926;
  assign n46158 = ~n45884 & n45936;
  assign n46159 = ~n46157 & ~n46158;
  assign n46160 = n45890 & ~n46159;
  assign n46161 = ~n45922 & ~n45944;
  assign n46162 = n45884 & ~n46161;
  assign n46163 = n45865 & n45871;
  assign n46164 = n45884 & n46163;
  assign n46165 = ~n45899 & n45910;
  assign n46166 = ~n46164 & ~n46165;
  assign n46167 = ~n45915 & n46166;
  assign n46168 = ~n45890 & ~n46167;
  assign n46169 = ~n46162 & ~n46168;
  assign n46170 = ~n46160 & n46169;
  assign n46171 = ~n46156 & n46170;
  assign n46172 = n45878 & ~n46171;
  assign n46173 = ~n46155 & ~n46172;
  assign n46174 = n45872 & n45884;
  assign n46175 = ~n45944 & ~n46174;
  assign n46176 = ~n45890 & ~n46175;
  assign n46177 = ~n45884 & n45941;
  assign n46178 = ~n46176 & ~n46177;
  assign n46179 = ~n45923 & ~n45938;
  assign n46180 = n45891 & n45914;
  assign n46181 = n45890 & n45902;
  assign n46182 = ~n45884 & n46181;
  assign n46183 = ~n46180 & ~n46182;
  assign n46184 = n45890 & n45901;
  assign n46185 = n46183 & ~n46184;
  assign n46186 = ~n45865 & n45905;
  assign n46187 = n46185 & ~n46186;
  assign n46188 = n46179 & n46187;
  assign n46189 = n46178 & n46188;
  assign n46190 = ~n45878 & ~n46189;
  assign n46191 = ~n45884 & n45890;
  assign n46192 = n45941 & n46191;
  assign n46193 = ~n46190 & ~n46192;
  assign po1164 = n46173 & n46193;
  assign n46195 = ~n45871 & ~n45899;
  assign n46196 = n45891 & n46195;
  assign n46197 = ~n45921 & ~n46196;
  assign n46198 = ~n46157 & n46197;
  assign n46199 = ~n45884 & n46163;
  assign n46200 = n46198 & ~n46199;
  assign n46201 = ~n45890 & n45922;
  assign n46202 = n46200 & ~n46201;
  assign n46203 = n45878 & ~n46202;
  assign n46204 = ~n45884 & n45915;
  assign n46205 = n45924 & ~n46204;
  assign n46206 = ~n46174 & n46205;
  assign n46207 = n45890 & ~n46206;
  assign n46208 = ~n46203 & ~n46207;
  assign n46209 = ~n45916 & ~n46156;
  assign n46210 = ~n45890 & ~n46209;
  assign n46211 = ~n45878 & n45890;
  assign n46212 = n45872 & n46211;
  assign n46213 = n45871 & ~n45884;
  assign n46214 = n45899 & n46213;
  assign n46215 = ~n46163 & ~n46214;
  assign n46216 = ~n45919 & n46215;
  assign n46217 = ~n45890 & ~n46216;
  assign n46218 = ~n45884 & n45937;
  assign n46219 = ~n46217 & ~n46218;
  assign n46220 = ~n45878 & ~n46219;
  assign n46221 = ~n46212 & ~n46220;
  assign n46222 = ~n46210 & n46221;
  assign n46223 = n46208 & n46222;
  assign n46224 = pi1232 & n46223;
  assign n46225 = ~pi1232 & ~n46223;
  assign po1167 = n46224 | n46225;
  assign n46227 = pi4040 & pi9040;
  assign n46228 = pi4021 & ~pi9040;
  assign n46229 = ~n46227 & ~n46228;
  assign n46230 = pi1174 & n46229;
  assign n46231 = ~pi1174 & ~n46229;
  assign n46232 = ~n46230 & ~n46231;
  assign n46233 = pi4133 & ~pi9040;
  assign n46234 = pi3964 & pi9040;
  assign n46235 = ~n46233 & ~n46234;
  assign n46236 = ~pi1176 & ~n46235;
  assign n46237 = pi1176 & n46235;
  assign n46238 = ~n46236 & ~n46237;
  assign n46239 = pi3956 & pi9040;
  assign n46240 = pi4024 & ~pi9040;
  assign n46241 = ~n46239 & ~n46240;
  assign n46242 = ~pi1180 & n46241;
  assign n46243 = pi1180 & ~n46241;
  assign n46244 = ~n46242 & ~n46243;
  assign n46245 = pi3945 & pi9040;
  assign n46246 = pi4025 & ~pi9040;
  assign n46247 = ~n46245 & ~n46246;
  assign n46248 = pi1159 & n46247;
  assign n46249 = ~pi1159 & ~n46247;
  assign n46250 = ~n46248 & ~n46249;
  assign n46251 = pi4277 & pi9040;
  assign n46252 = pi3952 & ~pi9040;
  assign n46253 = ~n46251 & ~n46252;
  assign n46254 = pi1173 & n46253;
  assign n46255 = ~pi1173 & ~n46253;
  assign n46256 = ~n46254 & ~n46255;
  assign n46257 = ~n46250 & ~n46256;
  assign n46258 = n46244 & n46257;
  assign n46259 = ~n46238 & n46258;
  assign n46260 = n46250 & ~n46256;
  assign n46261 = n46244 & n46260;
  assign n46262 = n46238 & n46261;
  assign n46263 = ~n46259 & ~n46262;
  assign n46264 = ~n46232 & ~n46263;
  assign n46265 = pi3932 & ~pi9040;
  assign n46266 = pi3962 & pi9040;
  assign n46267 = ~n46265 & ~n46266;
  assign n46268 = ~pi1171 & ~n46267;
  assign n46269 = pi1171 & n46267;
  assign n46270 = ~n46268 & ~n46269;
  assign n46271 = ~n46250 & n46256;
  assign n46272 = ~n46244 & n46271;
  assign n46273 = ~n46238 & n46272;
  assign n46274 = ~n46244 & n46260;
  assign n46275 = ~n46232 & n46274;
  assign n46276 = ~n46273 & ~n46275;
  assign n46277 = n46238 & ~n46244;
  assign n46278 = n46256 & n46277;
  assign n46279 = n46250 & n46278;
  assign n46280 = n46232 & n46238;
  assign n46281 = n46257 & n46280;
  assign n46282 = n46244 & n46281;
  assign n46283 = ~n46238 & n46250;
  assign n46284 = n46244 & n46283;
  assign n46285 = ~n46238 & ~n46250;
  assign n46286 = ~n46244 & n46285;
  assign n46287 = ~n46284 & ~n46286;
  assign n46288 = n46232 & ~n46287;
  assign n46289 = n46244 & n46271;
  assign n46290 = ~n46232 & n46289;
  assign n46291 = ~n46288 & ~n46290;
  assign n46292 = ~n46282 & n46291;
  assign n46293 = ~n46279 & n46292;
  assign n46294 = n46276 & n46293;
  assign n46295 = n46270 & ~n46294;
  assign n46296 = n46232 & n46273;
  assign n46297 = ~n46238 & n46275;
  assign n46298 = ~n46296 & ~n46297;
  assign n46299 = ~n46295 & n46298;
  assign n46300 = ~n46264 & n46299;
  assign n46301 = ~n46244 & n46257;
  assign n46302 = n46238 & n46301;
  assign n46303 = ~n46259 & ~n46302;
  assign n46304 = ~n46232 & n46238;
  assign n46305 = ~n46244 & ~n46250;
  assign n46306 = n46304 & n46305;
  assign n46307 = ~n46232 & n46258;
  assign n46308 = n46238 & n46260;
  assign n46309 = n46244 & n46256;
  assign n46310 = ~n46308 & ~n46309;
  assign n46311 = n46232 & ~n46310;
  assign n46312 = n46250 & n46256;
  assign n46313 = ~n46244 & n46312;
  assign n46314 = ~n46232 & n46313;
  assign n46315 = n46244 & n46312;
  assign n46316 = ~n46238 & n46315;
  assign n46317 = ~n46314 & ~n46316;
  assign n46318 = ~n46311 & n46317;
  assign n46319 = ~n46307 & n46318;
  assign n46320 = ~n46306 & n46319;
  assign n46321 = n46303 & n46320;
  assign n46322 = ~n46270 & ~n46321;
  assign po1171 = n46300 & ~n46322;
  assign n46324 = n46068 & n46093;
  assign n46325 = n46062 & n46107;
  assign n46326 = ~n46324 & ~n46325;
  assign n46327 = n46068 & ~n46074;
  assign n46328 = ~n46100 & ~n46327;
  assign n46329 = ~n46122 & n46328;
  assign n46330 = ~n46062 & ~n46329;
  assign n46331 = n46326 & ~n46330;
  assign n46332 = ~n46149 & n46331;
  assign n46333 = ~n46056 & ~n46332;
  assign n46334 = ~n46088 & n46135;
  assign n46335 = ~n46118 & ~n46334;
  assign n46336 = n46068 & n46107;
  assign n46337 = n46062 & n46100;
  assign n46338 = ~n46336 & ~n46337;
  assign n46339 = n46068 & n46148;
  assign n46340 = n46338 & ~n46339;
  assign n46341 = ~n46062 & n46136;
  assign n46342 = n46340 & ~n46341;
  assign n46343 = n46335 & n46342;
  assign n46344 = ~n46129 & n46343;
  assign n46345 = n46056 & ~n46344;
  assign n46346 = ~n46116 & ~n46119;
  assign n46347 = n46062 & n46102;
  assign n46348 = n46346 & ~n46347;
  assign n46349 = ~n46345 & n46348;
  assign po1175 = n46333 | ~n46349;
  assign n46351 = pi4192 & ~pi9040;
  assign n46352 = pi4021 & pi9040;
  assign n46353 = ~n46351 & ~n46352;
  assign n46354 = ~pi1158 & ~n46353;
  assign n46355 = pi1158 & n46353;
  assign n46356 = ~n46354 & ~n46355;
  assign n46357 = pi3945 & ~pi9040;
  assign n46358 = pi3953 & pi9040;
  assign n46359 = ~n46357 & ~n46358;
  assign n46360 = ~pi1164 & ~n46359;
  assign n46361 = pi1164 & n46359;
  assign n46362 = ~n46360 & ~n46361;
  assign n46363 = pi4133 & pi9040;
  assign n46364 = pi3937 & ~pi9040;
  assign n46365 = ~n46363 & ~n46364;
  assign n46366 = ~pi1131 & ~n46365;
  assign n46367 = pi1131 & n46365;
  assign n46368 = ~n46366 & ~n46367;
  assign n46369 = pi3952 & pi9040;
  assign n46370 = pi4126 & ~pi9040;
  assign n46371 = ~n46369 & ~n46370;
  assign n46372 = ~pi1146 & n46371;
  assign n46373 = pi1146 & ~n46371;
  assign n46374 = ~n46372 & ~n46373;
  assign n46375 = pi3933 & ~pi9040;
  assign n46376 = pi4029 & pi9040;
  assign n46377 = ~n46375 & ~n46376;
  assign n46378 = ~pi1178 & ~n46377;
  assign n46379 = pi1178 & n46377;
  assign n46380 = ~n46378 & ~n46379;
  assign n46381 = n46374 & n46380;
  assign n46382 = ~n46368 & n46381;
  assign n46383 = n46362 & n46382;
  assign n46384 = pi3956 & ~pi9040;
  assign n46385 = pi3971 & pi9040;
  assign n46386 = ~n46384 & ~n46385;
  assign n46387 = pi1165 & n46386;
  assign n46388 = ~pi1165 & ~n46386;
  assign n46389 = ~n46387 & ~n46388;
  assign n46390 = ~n46374 & n46380;
  assign n46391 = n46368 & n46390;
  assign n46392 = n46374 & ~n46380;
  assign n46393 = n46368 & n46392;
  assign n46394 = n46362 & n46393;
  assign n46395 = ~n46391 & ~n46394;
  assign n46396 = ~n46374 & ~n46380;
  assign n46397 = ~n46368 & n46396;
  assign n46398 = n46395 & ~n46397;
  assign n46399 = n46389 & ~n46398;
  assign n46400 = ~n46362 & n46389;
  assign n46401 = ~n46374 & n46400;
  assign n46402 = ~n46399 & ~n46401;
  assign n46403 = ~n46362 & n46392;
  assign n46404 = n46368 & n46381;
  assign n46405 = ~n46403 & ~n46404;
  assign n46406 = ~n46389 & ~n46405;
  assign n46407 = ~n46368 & ~n46374;
  assign n46408 = n46380 & n46407;
  assign n46409 = ~n46362 & n46408;
  assign n46410 = ~n46406 & ~n46409;
  assign n46411 = n46402 & n46410;
  assign n46412 = ~n46383 & n46411;
  assign n46413 = n46356 & ~n46412;
  assign n46414 = n46362 & n46368;
  assign n46415 = n46396 & n46414;
  assign n46416 = n46362 & ~n46368;
  assign n46417 = n46374 & n46416;
  assign n46418 = ~n46415 & ~n46417;
  assign n46419 = ~n46389 & ~n46418;
  assign n46420 = ~n46356 & ~n46389;
  assign n46421 = n46368 & ~n46374;
  assign n46422 = ~n46362 & n46396;
  assign n46423 = ~n46421 & ~n46422;
  assign n46424 = ~n46382 & n46423;
  assign n46425 = n46420 & ~n46424;
  assign n46426 = ~n46368 & n46392;
  assign n46427 = ~n46408 & ~n46426;
  assign n46428 = n46362 & ~n46427;
  assign n46429 = ~n46415 & ~n46428;
  assign n46430 = ~n46356 & ~n46429;
  assign n46431 = ~n46356 & n46389;
  assign n46432 = ~n46405 & n46431;
  assign n46433 = ~n46430 & ~n46432;
  assign n46434 = ~n46425 & n46433;
  assign n46435 = ~n46419 & n46434;
  assign po1178 = n46413 | ~n46435;
  assign n46437 = n46088 & ~n46092;
  assign n46438 = n46142 & n46437;
  assign n46439 = ~n46089 & ~n46121;
  assign n46440 = n46068 & ~n46439;
  assign n46441 = ~n46148 & ~n46440;
  assign n46442 = n46062 & ~n46441;
  assign n46443 = ~n46068 & n46081;
  assign n46444 = ~n46107 & ~n46443;
  assign n46445 = n46068 & n46114;
  assign n46446 = n46444 & ~n46445;
  assign n46447 = ~n46062 & ~n46446;
  assign n46448 = ~n46442 & ~n46447;
  assign n46449 = ~n46133 & ~n46339;
  assign n46450 = ~n46118 & n46449;
  assign n46451 = ~n46140 & n46450;
  assign n46452 = n46448 & n46451;
  assign n46453 = n46056 & ~n46452;
  assign n46454 = ~n46088 & n46092;
  assign n46455 = ~n46068 & n46454;
  assign n46456 = n46068 & n46122;
  assign n46457 = ~n46455 & ~n46456;
  assign n46458 = ~n46093 & ~n46096;
  assign n46459 = n46457 & n46458;
  assign n46460 = ~n46062 & ~n46459;
  assign n46461 = n46068 & n46117;
  assign n46462 = ~n46460 & ~n46461;
  assign n46463 = ~n46056 & ~n46462;
  assign n46464 = ~n46056 & n46062;
  assign n46465 = ~n46068 & n46089;
  assign n46466 = ~n46445 & ~n46465;
  assign n46467 = ~n46443 & n46466;
  assign n46468 = n46464 & ~n46467;
  assign n46469 = ~n46463 & ~n46468;
  assign n46470 = ~n46453 & n46469;
  assign n46471 = ~n46097 & n46470;
  assign po1181 = n46438 | ~n46471;
  assign n46473 = ~n45765 & n45802;
  assign n46474 = ~n45848 & ~n46473;
  assign n46475 = n45795 & n45811;
  assign n46476 = n45771 & n46475;
  assign n46477 = n45765 & n45820;
  assign n46478 = ~n45788 & n45797;
  assign n46479 = ~n46477 & ~n46478;
  assign n46480 = ~n45839 & n46479;
  assign n46481 = ~n46476 & n46480;
  assign n46482 = n45777 & n45795;
  assign n46483 = n45765 & n45771;
  assign n46484 = ~n45808 & ~n46483;
  assign n46485 = ~n46482 & n46484;
  assign n46486 = n45788 & ~n46485;
  assign n46487 = n46481 & ~n46486;
  assign n46488 = n46474 & n46487;
  assign n46489 = ~n45834 & ~n46488;
  assign n46490 = n45765 & n45800;
  assign n46491 = ~n45778 & ~n45826;
  assign n46492 = ~n45788 & ~n46491;
  assign n46493 = ~n45819 & ~n46492;
  assign n46494 = ~n46490 & n46493;
  assign n46495 = n45788 & n45798;
  assign n46496 = ~n45852 & ~n46495;
  assign n46497 = ~n45803 & n46496;
  assign n46498 = n46494 & n46497;
  assign n46499 = n45834 & ~n46498;
  assign po1184 = ~n46489 & ~n46499;
  assign n46501 = n46389 & ~n46427;
  assign n46502 = n46362 & n46390;
  assign n46503 = ~n46374 & n46416;
  assign n46504 = ~n46502 & ~n46503;
  assign n46505 = n46389 & ~n46504;
  assign n46506 = n46381 & n46389;
  assign n46507 = ~n46362 & n46506;
  assign n46508 = ~n46505 & ~n46507;
  assign n46509 = ~n46362 & n46368;
  assign n46510 = n46396 & n46509;
  assign n46511 = n46389 & n46510;
  assign n46512 = ~n46362 & n46404;
  assign n46513 = ~n46511 & ~n46512;
  assign n46514 = n46508 & n46513;
  assign n46515 = ~n46501 & n46514;
  assign n46516 = ~n46356 & ~n46515;
  assign n46517 = ~n46362 & n46397;
  assign n46518 = ~n46383 & ~n46517;
  assign n46519 = ~n46393 & n46518;
  assign n46520 = n46420 & ~n46519;
  assign n46521 = ~n46516 & ~n46520;
  assign n46522 = ~n46380 & n46416;
  assign n46523 = ~n46408 & ~n46522;
  assign n46524 = ~n46389 & n46523;
  assign n46525 = ~n46362 & ~n46368;
  assign n46526 = ~n46380 & n46525;
  assign n46527 = n46362 & n46381;
  assign n46528 = ~n46526 & ~n46527;
  assign n46529 = n46389 & n46528;
  assign n46530 = ~n46524 & ~n46529;
  assign n46531 = ~n46362 & n46380;
  assign n46532 = ~n46389 & n46531;
  assign n46533 = ~n46368 & n46532;
  assign n46534 = ~n46362 & n46393;
  assign n46535 = ~n46533 & ~n46534;
  assign n46536 = ~n46362 & n46391;
  assign n46537 = ~n46415 & ~n46536;
  assign n46538 = n46362 & n46404;
  assign n46539 = n46537 & ~n46538;
  assign n46540 = n46535 & n46539;
  assign n46541 = ~n46530 & n46540;
  assign n46542 = n46356 & ~n46541;
  assign n46543 = ~n46389 & ~n46537;
  assign n46544 = ~n46542 & ~n46543;
  assign po1187 = ~n46521 | ~n46544;
  assign n46546 = ~n45796 & ~n45799;
  assign n46547 = n45777 & ~n46546;
  assign n46548 = n45765 & n46547;
  assign n46549 = ~n46476 & ~n46548;
  assign n46550 = n45788 & ~n46549;
  assign n46551 = ~n45788 & n45839;
  assign n46552 = ~n46550 & ~n46551;
  assign n46553 = ~n45765 & n45813;
  assign n46554 = ~n46473 & ~n46553;
  assign n46555 = ~n45788 & n46554;
  assign n46556 = ~n45771 & ~n45777;
  assign n46557 = ~n45765 & n46556;
  assign n46558 = n45765 & n45799;
  assign n46559 = n45765 & n45780;
  assign n46560 = ~n46558 & ~n46559;
  assign n46561 = n45788 & n46560;
  assign n46562 = ~n46547 & n46561;
  assign n46563 = ~n46557 & n46562;
  assign n46564 = ~n46555 & ~n46563;
  assign n46565 = n46549 & ~n46564;
  assign n46566 = n45834 & ~n46565;
  assign n46567 = ~n45788 & ~n46546;
  assign n46568 = ~n45777 & n46567;
  assign n46569 = n45765 & n45801;
  assign n46570 = ~n45853 & ~n46569;
  assign n46571 = ~n45788 & ~n46570;
  assign n46572 = ~n46568 & ~n46571;
  assign n46573 = ~n45765 & n46567;
  assign n46574 = n46572 & ~n46573;
  assign n46575 = ~n45834 & ~n46574;
  assign n46576 = ~n46566 & ~n46575;
  assign n46577 = n45788 & ~n46554;
  assign n46578 = ~n45839 & ~n46577;
  assign n46579 = ~n45834 & ~n46578;
  assign n46580 = n46576 & ~n46579;
  assign po1190 = ~n46552 | ~n46580;
  assign n46582 = n45824 & ~n46546;
  assign n46583 = ~n46476 & ~n46582;
  assign n46584 = ~n45802 & n46583;
  assign n46585 = n45788 & ~n46584;
  assign n46586 = n45765 & n45840;
  assign n46587 = ~n46585 & ~n46586;
  assign n46588 = ~n45765 & n46482;
  assign n46589 = ~n46558 & ~n46588;
  assign n46590 = ~n45838 & n46589;
  assign n46591 = ~n45788 & ~n46590;
  assign n46592 = n46587 & ~n46591;
  assign n46593 = n45834 & ~n46592;
  assign n46594 = ~n45788 & n45798;
  assign n46595 = ~n46593 & ~n46594;
  assign n46596 = ~n45815 & ~n46559;
  assign n46597 = n45788 & ~n46596;
  assign n46598 = ~n45765 & n45799;
  assign n46599 = ~n45818 & ~n46598;
  assign n46600 = ~n45788 & ~n46599;
  assign n46601 = ~n45803 & ~n46600;
  assign n46602 = ~n45798 & ~n45853;
  assign n46603 = n45765 & n45808;
  assign n46604 = ~n46482 & ~n46603;
  assign n46605 = ~n45838 & n46604;
  assign n46606 = n45788 & ~n46605;
  assign n46607 = ~n45765 & n45840;
  assign n46608 = ~n46606 & ~n46607;
  assign n46609 = n46602 & n46608;
  assign n46610 = n46601 & n46609;
  assign n46611 = ~n45834 & ~n46610;
  assign n46612 = ~n46597 & ~n46611;
  assign po1193 = ~n46595 | ~n46612;
  assign n46614 = ~n45921 & ~n45927;
  assign n46615 = n45890 & ~n46614;
  assign n46616 = ~n45871 & n45899;
  assign n46617 = n45884 & n45936;
  assign n46618 = ~n46616 & ~n46617;
  assign n46619 = ~n45899 & n46213;
  assign n46620 = n46618 & ~n46619;
  assign n46621 = ~n45890 & ~n46620;
  assign n46622 = ~n45920 & ~n46621;
  assign n46623 = n45884 & n46181;
  assign n46624 = ~n46184 & ~n46623;
  assign n46625 = n46622 & n46624;
  assign n46626 = ~n45878 & ~n46625;
  assign n46627 = ~n45890 & n46616;
  assign n46628 = n45884 & n46627;
  assign n46629 = ~n46626 & ~n46628;
  assign n46630 = ~n45884 & n45901;
  assign n46631 = ~n45941 & ~n46630;
  assign n46632 = ~n45890 & ~n46631;
  assign n46633 = ~n45911 & ~n45944;
  assign n46634 = ~n45915 & n46633;
  assign n46635 = n45890 & ~n46634;
  assign n46636 = ~n45916 & ~n45938;
  assign n46637 = ~n46165 & n46636;
  assign n46638 = ~n46635 & n46637;
  assign n46639 = ~n46632 & n46638;
  assign n46640 = n45878 & ~n46639;
  assign n46641 = n46629 & ~n46640;
  assign n46642 = ~n45951 & n46641;
  assign po1199 = n46615 | ~n46642;
  assign n46644 = pi4131 & ~pi9040;
  assign n46645 = pi3963 & pi9040;
  assign n46646 = ~n46644 & ~n46645;
  assign n46647 = ~pi1155 & ~n46646;
  assign n46648 = pi1155 & n46646;
  assign n46649 = ~n46647 & ~n46648;
  assign n46650 = pi4193 & pi9040;
  assign n46651 = pi4132 & ~pi9040;
  assign n46652 = ~n46650 & ~n46651;
  assign n46653 = ~pi1169 & n46652;
  assign n46654 = pi1169 & ~n46652;
  assign n46655 = ~n46653 & ~n46654;
  assign n46656 = pi3957 & pi9040;
  assign n46657 = pi4043 & ~pi9040;
  assign n46658 = ~n46656 & ~n46657;
  assign n46659 = ~pi1173 & ~n46658;
  assign n46660 = pi1173 & n46658;
  assign n46661 = ~n46659 & ~n46660;
  assign n46662 = pi4023 & pi9040;
  assign n46663 = pi3968 & ~pi9040;
  assign n46664 = ~n46662 & ~n46663;
  assign n46665 = ~pi1183 & ~n46664;
  assign n46666 = pi1183 & n46664;
  assign n46667 = ~n46665 & ~n46666;
  assign n46668 = n46661 & ~n46667;
  assign n46669 = ~n46655 & n46668;
  assign n46670 = pi3965 & ~pi9040;
  assign n46671 = pi4118 & pi9040;
  assign n46672 = ~n46670 & ~n46671;
  assign n46673 = pi1157 & ~n46672;
  assign n46674 = ~pi1157 & n46672;
  assign n46675 = ~n46673 & ~n46674;
  assign n46676 = pi3948 & pi9040;
  assign n46677 = pi3949 & ~pi9040;
  assign n46678 = ~n46676 & ~n46677;
  assign n46679 = ~pi1171 & ~n46678;
  assign n46680 = pi1171 & n46678;
  assign n46681 = ~n46679 & ~n46680;
  assign n46682 = n46668 & ~n46681;
  assign n46683 = ~n46655 & n46681;
  assign n46684 = ~n46661 & n46683;
  assign n46685 = ~n46682 & ~n46684;
  assign n46686 = n46675 & ~n46685;
  assign n46687 = ~n46669 & ~n46686;
  assign n46688 = n46661 & n46681;
  assign n46689 = n46655 & n46688;
  assign n46690 = n46667 & n46689;
  assign n46691 = n46655 & ~n46681;
  assign n46692 = n46667 & n46691;
  assign n46693 = n46655 & ~n46661;
  assign n46694 = ~n46667 & n46693;
  assign n46695 = ~n46692 & ~n46694;
  assign n46696 = ~n46661 & ~n46681;
  assign n46697 = n46661 & n46683;
  assign n46698 = ~n46696 & ~n46697;
  assign n46699 = n46695 & n46698;
  assign n46700 = ~n46675 & ~n46699;
  assign n46701 = ~n46690 & ~n46700;
  assign n46702 = n46687 & n46701;
  assign n46703 = n46649 & ~n46702;
  assign n46704 = ~n46655 & ~n46681;
  assign n46705 = ~n46661 & n46704;
  assign n46706 = ~n46667 & n46705;
  assign n46707 = ~n46661 & n46691;
  assign n46708 = n46667 & n46707;
  assign n46709 = ~n46690 & ~n46708;
  assign n46710 = ~n46706 & n46709;
  assign n46711 = ~n46675 & ~n46710;
  assign n46712 = ~n46703 & ~n46711;
  assign n46713 = n46669 & n46681;
  assign n46714 = ~n46661 & n46681;
  assign n46715 = n46675 & n46714;
  assign n46716 = n46667 & n46715;
  assign n46717 = n46661 & n46704;
  assign n46718 = n46667 & n46717;
  assign n46719 = n46655 & n46661;
  assign n46720 = ~n46675 & n46719;
  assign n46721 = ~n46667 & n46720;
  assign n46722 = ~n46718 & ~n46721;
  assign n46723 = n46661 & n46667;
  assign n46724 = ~n46681 & n46723;
  assign n46725 = n46655 & n46681;
  assign n46726 = ~n46661 & n46725;
  assign n46727 = ~n46724 & ~n46726;
  assign n46728 = n46675 & ~n46727;
  assign n46729 = n46675 & n46696;
  assign n46730 = ~n46667 & n46729;
  assign n46731 = ~n46728 & ~n46730;
  assign n46732 = n46722 & n46731;
  assign n46733 = ~n46649 & ~n46732;
  assign n46734 = ~n46716 & ~n46733;
  assign n46735 = ~n46713 & n46734;
  assign po1204 = ~n46712 | ~n46735;
  assign n46737 = ~n46362 & n46382;
  assign n46738 = ~n46538 & ~n46737;
  assign n46739 = ~n46389 & ~n46738;
  assign n46740 = n46362 & ~n46389;
  assign n46741 = ~n46392 & ~n46408;
  assign n46742 = n46740 & ~n46741;
  assign n46743 = ~n46389 & n46392;
  assign n46744 = ~n46368 & n46743;
  assign n46745 = ~n46742 & ~n46744;
  assign n46746 = n46389 & n46421;
  assign n46747 = n46368 & n46400;
  assign n46748 = ~n46746 & ~n46747;
  assign n46749 = n46745 & n46748;
  assign n46750 = ~n46517 & n46749;
  assign n46751 = ~n46536 & n46750;
  assign n46752 = n46356 & ~n46751;
  assign n46753 = ~n46739 & ~n46752;
  assign n46754 = n46362 & n46426;
  assign n46755 = n46389 & n46754;
  assign n46756 = ~n46362 & n46746;
  assign n46757 = ~n46755 & ~n46756;
  assign n46758 = n46368 & ~n46380;
  assign n46759 = ~n46382 & ~n46758;
  assign n46760 = ~n46362 & ~n46759;
  assign n46761 = n46362 & n46396;
  assign n46762 = n46362 & n46421;
  assign n46763 = ~n46761 & ~n46762;
  assign n46764 = ~n46382 & n46763;
  assign n46765 = ~n46389 & ~n46764;
  assign n46766 = n46362 & n46389;
  assign n46767 = n46408 & n46766;
  assign n46768 = ~n46765 & ~n46767;
  assign n46769 = ~n46533 & n46768;
  assign n46770 = ~n46760 & n46769;
  assign n46771 = ~n46538 & n46770;
  assign n46772 = ~n46356 & ~n46771;
  assign n46773 = n46757 & ~n46772;
  assign po1207 = ~n46753 | ~n46773;
  assign n46775 = ~n46238 & ~n46244;
  assign n46776 = n46250 & n46775;
  assign n46777 = ~n46259 & ~n46776;
  assign n46778 = n46238 & n46244;
  assign n46779 = n46250 & n46778;
  assign n46780 = ~n46261 & ~n46779;
  assign n46781 = ~n46232 & ~n46780;
  assign n46782 = ~n46232 & n46271;
  assign n46783 = ~n46238 & n46782;
  assign n46784 = ~n46781 & ~n46783;
  assign n46785 = n46232 & n46258;
  assign n46786 = n46232 & n46312;
  assign n46787 = ~n46238 & n46786;
  assign n46788 = ~n46785 & ~n46787;
  assign n46789 = n46784 & n46788;
  assign n46790 = ~n46302 & n46789;
  assign n46791 = n46777 & n46790;
  assign n46792 = ~n46270 & ~n46791;
  assign n46793 = n46238 & n46289;
  assign n46794 = ~n46279 & ~n46793;
  assign n46795 = ~n46232 & ~n46238;
  assign n46796 = n46315 & n46795;
  assign n46797 = n46794 & ~n46796;
  assign n46798 = ~n46273 & ~n46308;
  assign n46799 = ~n46261 & n46798;
  assign n46800 = n46232 & ~n46799;
  assign n46801 = ~n46232 & n46301;
  assign n46802 = ~n46800 & ~n46801;
  assign n46803 = n46797 & n46802;
  assign n46804 = n46270 & ~n46803;
  assign n46805 = ~n46297 & ~n46306;
  assign n46806 = ~n46259 & n46794;
  assign n46807 = n46232 & ~n46806;
  assign n46808 = n46805 & ~n46807;
  assign n46809 = ~n46804 & n46808;
  assign po1210 = n46792 | ~n46809;
  assign n46811 = ~n46062 & n46089;
  assign n46812 = ~n46068 & n46811;
  assign n46813 = ~n46123 & ~n46812;
  assign n46814 = n46068 & n46437;
  assign n46815 = ~n46068 & n46074;
  assign n46816 = ~n46334 & ~n46815;
  assign n46817 = n46062 & ~n46816;
  assign n46818 = ~n46814 & ~n46817;
  assign n46819 = n46813 & n46818;
  assign n46820 = n46056 & ~n46819;
  assign n46821 = n46089 & n46139;
  assign n46822 = ~n46122 & ~n46461;
  assign n46823 = n46062 & ~n46822;
  assign n46824 = ~n46068 & n46106;
  assign n46825 = ~n46133 & ~n46824;
  assign n46826 = ~n46114 & n46825;
  assign n46827 = ~n46062 & ~n46826;
  assign n46828 = ~n46097 & ~n46827;
  assign n46829 = ~n46823 & n46828;
  assign n46830 = ~n46821 & n46829;
  assign n46831 = ~n46056 & ~n46830;
  assign n46832 = ~n46820 & ~n46831;
  assign n46833 = n46068 & n46458;
  assign n46834 = ~n46068 & ~n46121;
  assign n46835 = ~n46833 & ~n46834;
  assign n46836 = n46062 & n46835;
  assign n46837 = ~n46114 & ~n46148;
  assign n46838 = ~n46107 & n46837;
  assign n46839 = n46127 & ~n46838;
  assign n46840 = ~n46836 & ~n46839;
  assign po1213 = n46832 & n46840;
  assign n46842 = ~n46667 & n46689;
  assign n46843 = ~n46708 & ~n46842;
  assign n46844 = ~n46675 & ~n46843;
  assign n46845 = n46667 & n46705;
  assign n46846 = n46661 & n46691;
  assign n46847 = n46667 & n46846;
  assign n46848 = ~n46845 & ~n46847;
  assign n46849 = n46675 & ~n46848;
  assign n46850 = ~n46667 & n46846;
  assign n46851 = ~n46667 & n46726;
  assign n46852 = n46667 & n46719;
  assign n46853 = ~n46851 & ~n46852;
  assign n46854 = ~n46705 & ~n46713;
  assign n46855 = n46853 & n46854;
  assign n46856 = n46675 & ~n46855;
  assign n46857 = n46667 & n46683;
  assign n46858 = ~n46682 & ~n46857;
  assign n46859 = ~n46707 & n46858;
  assign n46860 = ~n46675 & ~n46859;
  assign n46861 = n46667 & n46684;
  assign n46862 = ~n46860 & ~n46861;
  assign n46863 = ~n46856 & n46862;
  assign n46864 = ~n46850 & n46863;
  assign n46865 = ~n46649 & ~n46864;
  assign n46866 = n46667 & n46675;
  assign n46867 = n46697 & n46866;
  assign n46868 = n46675 & n46707;
  assign n46869 = n46675 & n46717;
  assign n46870 = ~n46868 & ~n46869;
  assign n46871 = ~n46667 & ~n46870;
  assign n46872 = n46667 & n46726;
  assign n46873 = ~n46842 & ~n46872;
  assign n46874 = ~n46667 & n46683;
  assign n46875 = n46667 & n46704;
  assign n46876 = ~n46874 & ~n46875;
  assign n46877 = ~n46689 & n46876;
  assign n46878 = ~n46705 & n46877;
  assign n46879 = ~n46675 & ~n46878;
  assign n46880 = ~n46667 & n46684;
  assign n46881 = ~n46879 & ~n46880;
  assign n46882 = n46873 & n46881;
  assign n46883 = ~n46871 & n46882;
  assign n46884 = ~n46867 & n46883;
  assign n46885 = n46649 & ~n46884;
  assign n46886 = ~n46865 & ~n46885;
  assign n46887 = ~n46849 & n46886;
  assign po1216 = n46844 | ~n46887;
  assign n46889 = pi4134 & pi9040;
  assign n46890 = pi3964 & ~pi9040;
  assign n46891 = ~n46889 & ~n46890;
  assign n46892 = ~pi1159 & n46891;
  assign n46893 = pi1159 & ~n46891;
  assign n46894 = ~n46892 & ~n46893;
  assign n46895 = pi4126 & pi9040;
  assign n46896 = pi3934 & ~pi9040;
  assign n46897 = ~n46895 & ~n46896;
  assign n46898 = pi1145 & n46897;
  assign n46899 = ~pi1145 & ~n46897;
  assign n46900 = ~n46898 & ~n46899;
  assign n46901 = pi4040 & ~pi9040;
  assign n46902 = pi3961 & pi9040;
  assign n46903 = ~n46901 & ~n46902;
  assign n46904 = ~pi1178 & n46903;
  assign n46905 = pi1178 & ~n46903;
  assign n46906 = ~n46904 & ~n46905;
  assign n46907 = pi3959 & pi9040;
  assign n46908 = pi4210 & ~pi9040;
  assign n46909 = ~n46907 & ~n46908;
  assign n46910 = pi1158 & n46909;
  assign n46911 = ~pi1158 & ~n46909;
  assign n46912 = ~n46910 & ~n46911;
  assign n46913 = pi4024 & pi9040;
  assign n46914 = pi3938 & ~pi9040;
  assign n46915 = ~n46913 & ~n46914;
  assign n46916 = ~pi1180 & ~n46915;
  assign n46917 = pi1180 & n46915;
  assign n46918 = ~n46916 & ~n46917;
  assign n46919 = n46912 & ~n46918;
  assign n46920 = ~n46906 & n46919;
  assign n46921 = ~n46900 & n46920;
  assign n46922 = n46906 & n46918;
  assign n46923 = pi3962 & ~pi9040;
  assign n46924 = pi4119 & pi9040;
  assign n46925 = ~n46923 & ~n46924;
  assign n46926 = ~pi1168 & ~n46925;
  assign n46927 = pi1168 & n46925;
  assign n46928 = ~n46926 & ~n46927;
  assign n46929 = ~n46912 & n46918;
  assign n46930 = n46928 & n46929;
  assign n46931 = ~n46922 & ~n46930;
  assign n46932 = ~n46900 & ~n46931;
  assign n46933 = ~n46921 & ~n46932;
  assign n46934 = ~n46894 & ~n46933;
  assign n46935 = ~n46912 & ~n46918;
  assign n46936 = ~n46906 & n46935;
  assign n46937 = ~n46894 & n46936;
  assign n46938 = n46928 & n46937;
  assign n46939 = ~n46934 & ~n46938;
  assign n46940 = ~n46928 & n46935;
  assign n46941 = n46906 & n46940;
  assign n46942 = n46906 & n46928;
  assign n46943 = n46918 & n46942;
  assign n46944 = ~n46941 & ~n46943;
  assign n46945 = ~n46900 & ~n46944;
  assign n46946 = n46912 & n46918;
  assign n46947 = ~n46935 & ~n46946;
  assign n46948 = ~n46906 & ~n46928;
  assign n46949 = ~n46947 & n46948;
  assign n46950 = n46906 & ~n46928;
  assign n46951 = ~n46918 & n46950;
  assign n46952 = n46912 & n46951;
  assign n46953 = ~n46949 & ~n46952;
  assign n46954 = ~n46906 & n46929;
  assign n46955 = n46928 & n46954;
  assign n46956 = n46900 & n46955;
  assign n46957 = n46953 & ~n46956;
  assign n46958 = n46920 & n46928;
  assign n46959 = n46906 & ~n46947;
  assign n46960 = n46928 & n46959;
  assign n46961 = ~n46958 & ~n46960;
  assign n46962 = ~n46900 & ~n46928;
  assign n46963 = ~n46906 & ~n46912;
  assign n46964 = n46962 & n46963;
  assign n46965 = n46906 & n46929;
  assign n46966 = n46900 & ~n46928;
  assign n46967 = n46965 & n46966;
  assign n46968 = ~n46964 & ~n46967;
  assign n46969 = n46961 & n46968;
  assign n46970 = n46957 & n46969;
  assign n46971 = n46894 & ~n46970;
  assign n46972 = ~n46906 & n46946;
  assign n46973 = n46906 & n46919;
  assign n46974 = ~n46972 & ~n46973;
  assign n46975 = n46918 & n46948;
  assign n46976 = n46974 & ~n46975;
  assign n46977 = ~n46894 & n46900;
  assign n46978 = ~n46976 & n46977;
  assign n46979 = ~n46971 & ~n46978;
  assign n46980 = ~n46945 & n46979;
  assign po1220 = ~n46939 | ~n46980;
  assign n46982 = ~n46667 & n46704;
  assign n46983 = ~n46689 & ~n46982;
  assign n46984 = ~n46675 & ~n46983;
  assign n46985 = ~n46655 & ~n46661;
  assign n46986 = ~n46696 & ~n46985;
  assign n46987 = n46667 & ~n46986;
  assign n46988 = ~n46655 & n46667;
  assign n46989 = ~n46684 & ~n46988;
  assign n46990 = ~n46691 & n46989;
  assign n46991 = n46675 & ~n46990;
  assign n46992 = ~n46987 & ~n46991;
  assign n46993 = ~n46984 & n46992;
  assign n46994 = ~n46649 & ~n46993;
  assign n46995 = ~n46713 & ~n46872;
  assign n46996 = ~n46846 & ~n46874;
  assign n46997 = ~n46675 & ~n46996;
  assign n46998 = n46995 & ~n46997;
  assign n46999 = ~n46869 & n46998;
  assign n47000 = n46649 & ~n46999;
  assign n47001 = ~n46994 & ~n47000;
  assign n47002 = ~n46667 & n46707;
  assign n47003 = ~n46842 & ~n46861;
  assign n47004 = ~n47002 & n47003;
  assign n47005 = n46675 & ~n47004;
  assign n47006 = ~n46675 & n46851;
  assign n47007 = ~n46675 & n46845;
  assign n47008 = ~n47006 & ~n47007;
  assign n47009 = ~n47005 & n47008;
  assign po1223 = ~n47001 | ~n47009;
  assign n47011 = ~n46250 & n46778;
  assign n47012 = n46244 & ~n46256;
  assign n47013 = ~n47011 & ~n47012;
  assign n47014 = n46232 & ~n47013;
  assign n47015 = ~n46270 & n47014;
  assign n47016 = ~n46273 & ~n46284;
  assign n47017 = ~n46244 & n46304;
  assign n47018 = ~n46271 & n47017;
  assign n47019 = ~n46275 & ~n47018;
  assign n47020 = n47016 & n47019;
  assign n47021 = ~n46270 & ~n47020;
  assign n47022 = ~n46238 & n46301;
  assign n47023 = ~n46238 & n46313;
  assign n47024 = ~n47022 & ~n47023;
  assign n47025 = n46232 & ~n47024;
  assign n47026 = n46232 & n46261;
  assign n47027 = ~n46238 & n47026;
  assign n47028 = ~n47025 & ~n47027;
  assign n47029 = ~n46232 & n46273;
  assign n47030 = n47028 & ~n47029;
  assign n47031 = ~n47021 & n47030;
  assign n47032 = ~n47015 & n47031;
  assign n47033 = n46238 & n46782;
  assign n47034 = n46238 & n46272;
  assign n47035 = n46238 & n46312;
  assign n47036 = ~n46238 & n46289;
  assign n47037 = ~n47035 & ~n47036;
  assign n47038 = n46232 & ~n47037;
  assign n47039 = ~n47034 & ~n47038;
  assign n47040 = n46238 & n46274;
  assign n47041 = ~n47022 & ~n47040;
  assign n47042 = ~n46307 & n47041;
  assign n47043 = n47039 & n47042;
  assign n47044 = ~n47033 & n47043;
  assign n47045 = n46270 & ~n47044;
  assign n47046 = n47032 & ~n47045;
  assign po1226 = ~n46796 & n47046;
  assign n47048 = ~n46928 & n46929;
  assign n47049 = n46928 & n46935;
  assign n47050 = ~n47048 & ~n47049;
  assign n47051 = ~n46900 & ~n47050;
  assign n47052 = ~n46900 & n46952;
  assign n47053 = ~n47051 & ~n47052;
  assign n47054 = ~n46894 & ~n47053;
  assign n47055 = ~n46947 & n46950;
  assign n47056 = n46906 & n46912;
  assign n47057 = ~n46946 & ~n47056;
  assign n47058 = ~n46928 & ~n47057;
  assign n47059 = ~n46954 & ~n47058;
  assign n47060 = n46900 & ~n47059;
  assign n47061 = ~n47055 & ~n47060;
  assign n47062 = n46928 & n46965;
  assign n47063 = ~n46918 & n46948;
  assign n47064 = n46928 & ~n47057;
  assign n47065 = ~n47063 & ~n47064;
  assign n47066 = ~n46900 & ~n47065;
  assign n47067 = ~n47062 & ~n47066;
  assign n47068 = n47061 & n47067;
  assign n47069 = n46894 & ~n47068;
  assign n47070 = ~n46900 & n46942;
  assign n47071 = n46946 & n47070;
  assign n47072 = n46900 & n46928;
  assign n47073 = ~n46906 & n47072;
  assign n47074 = ~n46918 & n47073;
  assign n47075 = ~n47071 & ~n47074;
  assign n47076 = ~n46906 & n46928;
  assign n47077 = ~n46894 & ~n46946;
  assign n47078 = n47076 & n47077;
  assign n47079 = n47075 & ~n47078;
  assign n47080 = n46912 & n46928;
  assign n47081 = ~n46936 & ~n47080;
  assign n47082 = n46977 & ~n47081;
  assign n47083 = n47079 & ~n47082;
  assign n47084 = ~n47069 & n47083;
  assign n47085 = ~n47054 & n47084;
  assign n47086 = ~pi1221 & n47085;
  assign n47087 = pi1221 & ~n47085;
  assign po1228 = n47086 | n47087;
  assign n47089 = ~n46930 & ~n47055;
  assign n47090 = ~n46920 & n47089;
  assign n47091 = n46900 & ~n47090;
  assign n47092 = n46894 & n47091;
  assign n47093 = n46906 & n47080;
  assign n47094 = ~n47048 & ~n47093;
  assign n47095 = ~n46936 & n47094;
  assign n47096 = ~n47049 & n47095;
  assign n47097 = ~n46900 & ~n47096;
  assign n47098 = n46928 & n46973;
  assign n47099 = ~n47097 & ~n47098;
  assign n47100 = n46894 & ~n47099;
  assign n47101 = n46954 & n46962;
  assign n47102 = ~n47052 & ~n47101;
  assign n47103 = n46900 & ~n46950;
  assign n47104 = ~n46947 & n47103;
  assign n47105 = ~n46906 & n47080;
  assign n47106 = ~n46930 & ~n47105;
  assign n47107 = ~n46900 & ~n47106;
  assign n47108 = ~n46929 & n46962;
  assign n47109 = n46906 & n47108;
  assign n47110 = ~n47107 & ~n47109;
  assign n47111 = ~n46952 & ~n46967;
  assign n47112 = n47110 & n47111;
  assign n47113 = ~n47104 & n47112;
  assign n47114 = ~n46894 & ~n47113;
  assign n47115 = n47102 & ~n47114;
  assign n47116 = n46972 & n47072;
  assign n47117 = n47115 & ~n47116;
  assign n47118 = ~n47100 & n47117;
  assign po1230 = n47092 | ~n47118;
  assign n47120 = ~n46965 & ~n46972;
  assign n47121 = ~n46940 & n47120;
  assign n47122 = n46900 & ~n47121;
  assign n47123 = n46906 & n46946;
  assign n47124 = ~n46954 & ~n47123;
  assign n47125 = ~n46900 & ~n47124;
  assign n47126 = ~n47122 & ~n47125;
  assign n47127 = ~n46921 & n47126;
  assign n47128 = ~n46941 & n47127;
  assign n47129 = n46894 & ~n47128;
  assign n47130 = n46919 & ~n46928;
  assign n47131 = ~n47049 & ~n47130;
  assign n47132 = n46900 & ~n47131;
  assign n47133 = ~n46955 & ~n47132;
  assign n47134 = ~n46900 & n46936;
  assign n47135 = ~n46965 & ~n47134;
  assign n47136 = n46974 & n47135;
  assign n47137 = ~n46928 & ~n47136;
  assign n47138 = n47133 & ~n47137;
  assign n47139 = ~n46894 & ~n47138;
  assign n47140 = n46906 & n47049;
  assign n47141 = ~n46958 & ~n47140;
  assign n47142 = ~n46900 & ~n47141;
  assign n47143 = n47056 & n47072;
  assign n47144 = ~n47142 & ~n47143;
  assign n47145 = ~n47139 & n47144;
  assign po1233 = n47129 | ~n47145;
  assign n47147 = ~n46502 & ~n46534;
  assign n47148 = n46389 & ~n47147;
  assign n47149 = n46368 & n46740;
  assign n47150 = ~n46525 & ~n47149;
  assign n47151 = n46374 & ~n47150;
  assign n47152 = n46389 & n46391;
  assign n47153 = n46362 & n46408;
  assign n47154 = ~n47152 & ~n47153;
  assign n47155 = ~n46415 & n47154;
  assign n47156 = ~n46526 & n47155;
  assign n47157 = ~n47151 & n47156;
  assign n47158 = ~n46356 & ~n47157;
  assign n47159 = ~n47148 & ~n47158;
  assign n47160 = n46389 & n46759;
  assign n47161 = ~n46362 & n46390;
  assign n47162 = ~n46397 & ~n47161;
  assign n47163 = ~n46389 & n47162;
  assign n47164 = ~n47160 & ~n47163;
  assign n47165 = ~n46754 & ~n47164;
  assign n47166 = n46356 & ~n47165;
  assign n47167 = ~n46389 & n46404;
  assign n47168 = ~n47166 & ~n47167;
  assign n47169 = n47159 & n47168;
  assign n47170 = pi1213 & n47169;
  assign n47171 = ~pi1213 & ~n47169;
  assign po1235 = n47170 | n47171;
  assign n47173 = n46274 & n46280;
  assign n47174 = ~n46282 & ~n47173;
  assign n47175 = ~n46284 & ~n46309;
  assign n47176 = ~n46232 & ~n47175;
  assign n47177 = n46270 & n47176;
  assign n47178 = ~n46238 & n46260;
  assign n47179 = ~n46315 & ~n47178;
  assign n47180 = n46232 & ~n47179;
  assign n47181 = ~n46273 & ~n46279;
  assign n47182 = ~n46238 & n46257;
  assign n47183 = ~n46262 & ~n47182;
  assign n47184 = ~n46232 & ~n47183;
  assign n47185 = ~n46238 & n46274;
  assign n47186 = ~n47184 & ~n47185;
  assign n47187 = n47181 & n47186;
  assign n47188 = ~n47180 & n47187;
  assign n47189 = ~n46270 & ~n47188;
  assign n47190 = ~n46279 & ~n46302;
  assign n47191 = ~n46793 & n47190;
  assign n47192 = ~n46232 & ~n47191;
  assign n47193 = ~n47189 & ~n47192;
  assign n47194 = ~n47011 & ~n47040;
  assign n47195 = n46270 & ~n47194;
  assign n47196 = n46256 & n46775;
  assign n47197 = ~n46286 & ~n47196;
  assign n47198 = ~n46272 & n47197;
  assign n47199 = n46232 & ~n47198;
  assign n47200 = n46270 & n47199;
  assign n47201 = ~n47195 & ~n47200;
  assign n47202 = n47193 & n47201;
  assign n47203 = ~n47177 & n47202;
  assign po1237 = ~n47174 | ~n47203;
  assign n47205 = n46667 & n46720;
  assign n47206 = ~n46675 & n46717;
  assign n47207 = ~n46667 & n47206;
  assign n47208 = ~n47205 & ~n47207;
  assign n47209 = ~n46667 & n46681;
  assign n47210 = n46675 & n47209;
  assign n47211 = ~n46684 & ~n47002;
  assign n47212 = ~n46675 & ~n47211;
  assign n47213 = ~n47210 & ~n47212;
  assign n47214 = n46848 & n47213;
  assign n47215 = n46649 & ~n47214;
  assign n47216 = ~n46682 & ~n47006;
  assign n47217 = ~n46717 & ~n46982;
  assign n47218 = ~n46684 & n47217;
  assign n47219 = n46675 & ~n47218;
  assign n47220 = ~n46675 & n46697;
  assign n47221 = ~n47219 & ~n47220;
  assign n47222 = n47216 & n47221;
  assign n47223 = n46709 & n47222;
  assign n47224 = ~n46649 & ~n47223;
  assign n47225 = n46675 & n46872;
  assign n47226 = ~n47224 & ~n47225;
  assign n47227 = ~n47215 & n47226;
  assign n47228 = ~n47007 & n47227;
  assign po1240 = ~n47208 | ~n47228;
  assign n47230 = pi4110 & pi9040;
  assign n47231 = pi4125 & ~pi9040;
  assign n47232 = ~n47230 & ~n47231;
  assign n47233 = ~pi1240 & ~n47232;
  assign n47234 = pi1240 & n47232;
  assign n47235 = ~n47233 & ~n47234;
  assign n47236 = pi4069 & pi9040;
  assign n47237 = pi4203 & ~pi9040;
  assign n47238 = ~n47236 & ~n47237;
  assign n47239 = ~pi1236 & ~n47238;
  assign n47240 = pi1236 & n47238;
  assign n47241 = ~n47239 & ~n47240;
  assign n47242 = ~n47235 & ~n47241;
  assign n47243 = pi4307 & pi9040;
  assign n47244 = pi4212 & ~pi9040;
  assign n47245 = ~n47243 & ~n47244;
  assign n47246 = pi1222 & n47245;
  assign n47247 = ~pi1222 & ~n47245;
  assign n47248 = ~n47246 & ~n47247;
  assign n47249 = pi4075 & ~pi9040;
  assign n47250 = pi4100 & pi9040;
  assign n47251 = ~n47249 & ~n47250;
  assign n47252 = ~pi1245 & ~n47251;
  assign n47253 = pi1245 & n47251;
  assign n47254 = ~n47252 & ~n47253;
  assign n47255 = pi4069 & ~pi9040;
  assign n47256 = pi4209 & pi9040;
  assign n47257 = ~n47255 & ~n47256;
  assign n47258 = pi1206 & n47257;
  assign n47259 = ~pi1206 & ~n47257;
  assign n47260 = ~n47258 & ~n47259;
  assign n47261 = n47254 & ~n47260;
  assign n47262 = ~n47248 & n47261;
  assign n47263 = pi4307 & ~pi9040;
  assign n47264 = pi4125 & pi9040;
  assign n47265 = ~n47263 & ~n47264;
  assign n47266 = ~pi1239 & ~n47265;
  assign n47267 = pi1239 & n47265;
  assign n47268 = ~n47266 & ~n47267;
  assign n47269 = n47260 & ~n47268;
  assign n47270 = n47254 & n47269;
  assign n47271 = n47248 & n47270;
  assign n47272 = n47260 & n47268;
  assign n47273 = ~n47248 & n47272;
  assign n47274 = ~n47271 & ~n47273;
  assign n47275 = ~n47262 & n47274;
  assign n47276 = n47242 & ~n47275;
  assign n47277 = ~n47248 & ~n47254;
  assign n47278 = ~n47268 & n47277;
  assign n47279 = ~n47260 & ~n47268;
  assign n47280 = n47254 & n47279;
  assign n47281 = n47248 & n47280;
  assign n47282 = ~n47278 & ~n47281;
  assign n47283 = ~n47254 & n47269;
  assign n47284 = n47254 & n47260;
  assign n47285 = n47268 & n47284;
  assign n47286 = ~n47283 & ~n47285;
  assign n47287 = n47282 & n47286;
  assign n47288 = n47235 & ~n47287;
  assign n47289 = ~n47260 & n47268;
  assign n47290 = ~n47254 & n47289;
  assign n47291 = n47248 & n47290;
  assign n47292 = ~n47288 & ~n47291;
  assign n47293 = ~n47241 & ~n47292;
  assign n47294 = ~n47276 & ~n47293;
  assign n47295 = ~n47272 & ~n47279;
  assign n47296 = n47248 & ~n47295;
  assign n47297 = ~n47254 & n47279;
  assign n47298 = ~n47296 & ~n47297;
  assign n47299 = ~n47235 & ~n47298;
  assign n47300 = n47254 & n47289;
  assign n47301 = ~n47262 & ~n47300;
  assign n47302 = ~n47271 & n47301;
  assign n47303 = n47235 & ~n47302;
  assign n47304 = ~n47299 & ~n47303;
  assign n47305 = ~n47235 & ~n47248;
  assign n47306 = n47269 & n47305;
  assign n47307 = n47248 & ~n47254;
  assign n47308 = ~n47268 & n47307;
  assign n47309 = ~n47260 & n47308;
  assign n47310 = ~n47254 & n47260;
  assign n47311 = n47268 & n47310;
  assign n47312 = n47248 & n47311;
  assign n47313 = ~n47309 & ~n47312;
  assign n47314 = n47268 & n47277;
  assign n47315 = ~n47260 & n47314;
  assign n47316 = n47313 & ~n47315;
  assign n47317 = ~n47306 & n47316;
  assign n47318 = n47304 & n47317;
  assign n47319 = n47241 & ~n47318;
  assign n47320 = n47235 & ~n47248;
  assign n47321 = n47254 & n47320;
  assign n47322 = n47268 & n47321;
  assign n47323 = ~n47248 & n47283;
  assign n47324 = ~n47322 & ~n47323;
  assign n47325 = ~n47319 & n47324;
  assign n47326 = n47294 & n47325;
  assign n47327 = pi1254 & ~n47326;
  assign n47328 = ~pi1254 & n47324;
  assign n47329 = n47294 & n47328;
  assign n47330 = ~n47319 & n47329;
  assign po1316 = n47327 | n47330;
  assign n47332 = pi4123 & ~pi9040;
  assign n47333 = pi4203 & pi9040;
  assign n47334 = ~n47332 & ~n47333;
  assign n47335 = pi1214 & n47334;
  assign n47336 = ~pi1214 & ~n47334;
  assign n47337 = ~n47335 & ~n47336;
  assign n47338 = pi4088 & ~pi9040;
  assign n47339 = pi4383 & pi9040;
  assign n47340 = ~n47338 & ~n47339;
  assign n47341 = pi1237 & n47340;
  assign n47342 = ~pi1237 & ~n47340;
  assign n47343 = ~n47341 & ~n47342;
  assign n47344 = pi4110 & ~pi9040;
  assign n47345 = pi4111 & pi9040;
  assign n47346 = ~n47344 & ~n47345;
  assign n47347 = ~pi1210 & n47346;
  assign n47348 = pi1210 & ~n47346;
  assign n47349 = ~n47347 & ~n47348;
  assign n47350 = pi4184 & ~pi9040;
  assign n47351 = pi4136 & pi9040;
  assign n47352 = ~n47350 & ~n47351;
  assign n47353 = ~pi1226 & n47352;
  assign n47354 = pi1226 & ~n47352;
  assign n47355 = ~n47353 & ~n47354;
  assign n47356 = pi4279 & pi9040;
  assign n47357 = pi4299 & ~pi9040;
  assign n47358 = ~n47356 & ~n47357;
  assign n47359 = ~pi1209 & n47358;
  assign n47360 = pi1209 & ~n47358;
  assign n47361 = ~n47359 & ~n47360;
  assign n47362 = n47355 & n47361;
  assign n47363 = ~n47349 & n47362;
  assign n47364 = n47343 & n47363;
  assign n47365 = ~n47355 & n47361;
  assign n47366 = n47349 & n47365;
  assign n47367 = n47343 & n47366;
  assign n47368 = ~n47364 & ~n47367;
  assign n47369 = ~n47355 & ~n47361;
  assign n47370 = n47349 & n47369;
  assign n47371 = ~n47343 & n47370;
  assign n47372 = n47349 & n47362;
  assign n47373 = ~n47343 & n47372;
  assign n47374 = ~n47371 & ~n47373;
  assign n47375 = n47368 & n47374;
  assign n47376 = n47337 & ~n47375;
  assign n47377 = n47355 & ~n47361;
  assign n47378 = n47349 & n47377;
  assign n47379 = n47343 & n47378;
  assign n47380 = ~n47366 & ~n47379;
  assign n47381 = n47337 & ~n47380;
  assign n47382 = ~n47343 & ~n47361;
  assign n47383 = ~n47337 & n47382;
  assign n47384 = ~n47349 & ~n47355;
  assign n47385 = n47343 & n47362;
  assign n47386 = ~n47384 & ~n47385;
  assign n47387 = ~n47337 & ~n47386;
  assign n47388 = ~n47383 & ~n47387;
  assign n47389 = ~n47349 & n47377;
  assign n47390 = ~n47343 & n47389;
  assign n47391 = n47388 & ~n47390;
  assign n47392 = n47343 & ~n47361;
  assign n47393 = ~n47349 & n47392;
  assign n47394 = ~n47355 & n47393;
  assign n47395 = n47391 & ~n47394;
  assign n47396 = ~n47381 & n47395;
  assign n47397 = pi4136 & ~pi9040;
  assign n47398 = pi4216 & pi9040;
  assign n47399 = ~n47397 & ~n47398;
  assign n47400 = ~pi1246 & ~n47399;
  assign n47401 = pi1246 & n47399;
  assign n47402 = ~n47400 & ~n47401;
  assign n47403 = ~n47396 & ~n47402;
  assign n47404 = n47349 & ~n47361;
  assign n47405 = ~n47337 & n47343;
  assign n47406 = n47402 & n47405;
  assign n47407 = n47404 & n47406;
  assign n47408 = ~n47343 & n47349;
  assign n47409 = n47361 & n47408;
  assign n47410 = ~n47337 & ~n47409;
  assign n47411 = n47343 & ~n47349;
  assign n47412 = n47355 & n47411;
  assign n47413 = ~n47369 & ~n47404;
  assign n47414 = ~n47343 & ~n47413;
  assign n47415 = ~n47363 & ~n47414;
  assign n47416 = n47337 & n47415;
  assign n47417 = ~n47412 & n47416;
  assign n47418 = ~n47410 & ~n47417;
  assign n47419 = ~n47349 & n47365;
  assign n47420 = n47343 & n47419;
  assign n47421 = ~n47418 & ~n47420;
  assign n47422 = n47402 & ~n47421;
  assign n47423 = ~n47407 & ~n47422;
  assign n47424 = ~n47403 & n47423;
  assign n47425 = ~n47376 & n47424;
  assign n47426 = ~n47337 & ~n47343;
  assign n47427 = n47377 & n47426;
  assign n47428 = ~n47349 & n47427;
  assign n47429 = n47425 & ~n47428;
  assign n47430 = pi1248 & ~n47429;
  assign n47431 = ~pi1248 & ~n47428;
  assign n47432 = n47424 & n47431;
  assign n47433 = ~n47376 & n47432;
  assign po1317 = n47430 | n47433;
  assign n47435 = n47248 & n47261;
  assign n47436 = ~n47285 & ~n47435;
  assign n47437 = ~n47323 & n47436;
  assign n47438 = n47235 & ~n47437;
  assign n47439 = ~n47248 & n47311;
  assign n47440 = ~n47248 & n47300;
  assign n47441 = ~n47254 & ~n47260;
  assign n47442 = ~n47269 & ~n47441;
  assign n47443 = n47248 & ~n47442;
  assign n47444 = ~n47440 & ~n47443;
  assign n47445 = ~n47439 & n47444;
  assign n47446 = ~n47235 & ~n47445;
  assign n47447 = ~n47438 & ~n47446;
  assign n47448 = n47241 & ~n47447;
  assign n47449 = ~n47260 & n47320;
  assign n47450 = ~n47248 & n47260;
  assign n47451 = n47254 & n47450;
  assign n47452 = ~n47435 & ~n47451;
  assign n47453 = ~n47235 & ~n47452;
  assign n47454 = ~n47306 & ~n47453;
  assign n47455 = ~n47248 & n47270;
  assign n47456 = ~n47312 & ~n47455;
  assign n47457 = n47235 & n47310;
  assign n47458 = n47248 & n47457;
  assign n47459 = n47235 & n47290;
  assign n47460 = ~n47458 & ~n47459;
  assign n47461 = n47456 & n47460;
  assign n47462 = n47454 & n47461;
  assign n47463 = ~n47449 & n47462;
  assign n47464 = ~n47241 & ~n47463;
  assign n47465 = ~n47235 & n47455;
  assign n47466 = ~n47235 & n47297;
  assign n47467 = ~n47248 & n47466;
  assign n47468 = ~n47465 & ~n47467;
  assign n47469 = n47235 & n47315;
  assign n47470 = n47468 & ~n47469;
  assign n47471 = ~n47248 & n47280;
  assign n47472 = n47248 & n47272;
  assign n47473 = ~n47471 & ~n47472;
  assign n47474 = n47235 & ~n47473;
  assign n47475 = n47470 & ~n47474;
  assign n47476 = ~n47464 & n47475;
  assign n47477 = ~n47448 & n47476;
  assign n47478 = ~pi1261 & n47477;
  assign n47479 = pi1261 & ~n47477;
  assign po1331 = n47478 | n47479;
  assign n47481 = n47235 & n47272;
  assign n47482 = ~n47248 & n47481;
  assign n47483 = ~n47471 & ~n47482;
  assign n47484 = ~n47248 & n47254;
  assign n47485 = ~n47268 & n47484;
  assign n47486 = ~n47248 & ~n47260;
  assign n47487 = ~n47485 & ~n47486;
  assign n47488 = ~n47235 & ~n47487;
  assign n47489 = n47248 & n47254;
  assign n47490 = n47268 & n47489;
  assign n47491 = ~n47488 & ~n47490;
  assign n47492 = n47483 & n47491;
  assign n47493 = n47241 & ~n47492;
  assign n47494 = ~n47270 & ~n47312;
  assign n47495 = ~n47248 & n47289;
  assign n47496 = n47494 & ~n47495;
  assign n47497 = n47235 & ~n47496;
  assign n47498 = n47272 & n47305;
  assign n47499 = ~n47323 & ~n47498;
  assign n47500 = ~n47497 & n47499;
  assign n47501 = ~n47280 & ~n47291;
  assign n47502 = ~n47235 & ~n47501;
  assign n47503 = n47500 & ~n47502;
  assign n47504 = ~n47241 & ~n47503;
  assign n47505 = ~n47493 & ~n47504;
  assign n47506 = n47248 & n47286;
  assign n47507 = ~n47248 & ~n47279;
  assign n47508 = ~n47506 & ~n47507;
  assign n47509 = ~n47235 & n47508;
  assign n47510 = n47235 & n47248;
  assign n47511 = ~n47297 & ~n47300;
  assign n47512 = ~n47270 & n47511;
  assign n47513 = n47510 & ~n47512;
  assign n47514 = ~n47509 & ~n47513;
  assign n47515 = n47505 & n47514;
  assign n47516 = ~pi1263 & ~n47515;
  assign n47517 = pi1263 & n47514;
  assign n47518 = ~n47504 & n47517;
  assign n47519 = ~n47493 & n47518;
  assign po1332 = n47516 | n47519;
  assign n47521 = pi4383 & ~pi9040;
  assign n47522 = pi4098 & pi9040;
  assign n47523 = ~n47521 & ~n47522;
  assign n47524 = ~pi1206 & ~n47523;
  assign n47525 = pi1206 & n47523;
  assign n47526 = ~n47524 & ~n47525;
  assign n47527 = pi4298 & pi9040;
  assign n47528 = pi4104 & ~pi9040;
  assign n47529 = ~n47527 & ~n47528;
  assign n47530 = pi1231 & n47529;
  assign n47531 = ~pi1231 & ~n47529;
  assign n47532 = ~n47530 & ~n47531;
  assign n47533 = pi4114 & ~pi9040;
  assign n47534 = pi4127 & pi9040;
  assign n47535 = ~n47533 & ~n47534;
  assign n47536 = pi1235 & n47535;
  assign n47537 = ~pi1235 & ~n47535;
  assign n47538 = ~n47536 & ~n47537;
  assign n47539 = pi4207 & pi9040;
  assign n47540 = pi4135 & ~pi9040;
  assign n47541 = ~n47539 & ~n47540;
  assign n47542 = ~pi1225 & ~n47541;
  assign n47543 = pi1225 & n47541;
  assign n47544 = ~n47542 & ~n47543;
  assign n47545 = pi4135 & pi9040;
  assign n47546 = pi4209 & ~pi9040;
  assign n47547 = ~n47545 & ~n47546;
  assign n47548 = pi1245 & n47547;
  assign n47549 = ~pi1245 & ~n47547;
  assign n47550 = ~n47548 & ~n47549;
  assign n47551 = n47544 & ~n47550;
  assign n47552 = n47538 & n47551;
  assign n47553 = n47532 & n47552;
  assign n47554 = pi4038 & pi9040;
  assign n47555 = pi4100 & ~pi9040;
  assign n47556 = ~n47554 & ~n47555;
  assign n47557 = ~pi1220 & n47556;
  assign n47558 = pi1220 & ~n47556;
  assign n47559 = ~n47557 & ~n47558;
  assign n47560 = n47538 & n47550;
  assign n47561 = n47544 & n47560;
  assign n47562 = ~n47538 & ~n47544;
  assign n47563 = ~n47544 & ~n47550;
  assign n47564 = ~n47532 & n47563;
  assign n47565 = ~n47538 & ~n47550;
  assign n47566 = n47532 & n47565;
  assign n47567 = ~n47564 & ~n47566;
  assign n47568 = ~n47562 & n47567;
  assign n47569 = ~n47561 & n47568;
  assign n47570 = ~n47559 & ~n47569;
  assign n47571 = ~n47532 & n47544;
  assign n47572 = n47550 & n47571;
  assign n47573 = ~n47538 & n47571;
  assign n47574 = ~n47544 & n47560;
  assign n47575 = ~n47573 & ~n47574;
  assign n47576 = n47559 & ~n47575;
  assign n47577 = ~n47572 & ~n47576;
  assign n47578 = ~n47570 & n47577;
  assign n47579 = ~n47553 & n47578;
  assign n47580 = n47526 & ~n47579;
  assign n47581 = ~n47538 & n47550;
  assign n47582 = ~n47544 & n47581;
  assign n47583 = ~n47532 & n47582;
  assign n47584 = ~n47544 & n47565;
  assign n47585 = n47532 & n47584;
  assign n47586 = ~n47553 & ~n47585;
  assign n47587 = ~n47583 & n47586;
  assign n47588 = ~n47559 & ~n47587;
  assign n47589 = ~n47580 & ~n47588;
  assign n47590 = ~n47532 & n47561;
  assign n47591 = n47532 & ~n47544;
  assign n47592 = n47559 & n47591;
  assign n47593 = n47538 & n47592;
  assign n47594 = n47532 & n47544;
  assign n47595 = n47550 & n47594;
  assign n47596 = ~n47538 & n47595;
  assign n47597 = n47551 & ~n47559;
  assign n47598 = ~n47532 & n47597;
  assign n47599 = ~n47596 & ~n47598;
  assign n47600 = ~n47538 & n47544;
  assign n47601 = n47532 & n47600;
  assign n47602 = n47538 & ~n47550;
  assign n47603 = ~n47544 & n47602;
  assign n47604 = ~n47601 & ~n47603;
  assign n47605 = n47559 & ~n47604;
  assign n47606 = n47559 & n47562;
  assign n47607 = ~n47532 & n47606;
  assign n47608 = ~n47605 & ~n47607;
  assign n47609 = n47599 & n47608;
  assign n47610 = ~n47526 & ~n47609;
  assign n47611 = ~n47593 & ~n47610;
  assign n47612 = ~n47590 & n47611;
  assign n47613 = n47589 & n47612;
  assign n47614 = ~pi1256 & ~n47613;
  assign n47615 = ~n47580 & ~n47590;
  assign n47616 = ~n47588 & n47615;
  assign n47617 = n47611 & n47616;
  assign n47618 = pi1256 & n47617;
  assign po1337 = n47614 | n47618;
  assign n47620 = pi4300 & pi9040;
  assign n47621 = pi4099 & ~pi9040;
  assign n47622 = ~n47620 & ~n47621;
  assign n47623 = ~pi1229 & n47622;
  assign n47624 = pi1229 & ~n47622;
  assign n47625 = ~n47623 & ~n47624;
  assign n47626 = pi4106 & pi9040;
  assign n47627 = pi4122 & ~pi9040;
  assign n47628 = ~n47626 & ~n47627;
  assign n47629 = ~pi1226 & n47628;
  assign n47630 = pi1226 & ~n47628;
  assign n47631 = ~n47629 & ~n47630;
  assign n47632 = pi4106 & ~pi9040;
  assign n47633 = pi4124 & pi9040;
  assign n47634 = ~n47632 & ~n47633;
  assign n47635 = ~pi1246 & ~n47634;
  assign n47636 = pi1246 & n47634;
  assign n47637 = ~n47635 & ~n47636;
  assign n47638 = pi4105 & ~pi9040;
  assign n47639 = pi4301 & pi9040;
  assign n47640 = ~n47638 & ~n47639;
  assign n47641 = ~pi1216 & ~n47640;
  assign n47642 = pi1216 & n47640;
  assign n47643 = ~n47641 & ~n47642;
  assign n47644 = ~n47637 & n47643;
  assign n47645 = pi4169 & pi9040;
  assign n47646 = pi4124 & ~pi9040;
  assign n47647 = ~n47645 & ~n47646;
  assign n47648 = ~pi1217 & ~n47647;
  assign n47649 = pi1217 & n47647;
  assign n47650 = ~n47648 & ~n47649;
  assign n47651 = pi4121 & pi9040;
  assign n47652 = pi4295 & ~pi9040;
  assign n47653 = ~n47651 & ~n47652;
  assign n47654 = pi1247 & n47653;
  assign n47655 = ~pi1247 & ~n47653;
  assign n47656 = ~n47654 & ~n47655;
  assign n47657 = n47650 & n47656;
  assign n47658 = n47644 & n47657;
  assign n47659 = ~n47631 & n47658;
  assign n47660 = ~n47631 & ~n47650;
  assign n47661 = ~n47643 & n47660;
  assign n47662 = ~n47637 & n47661;
  assign n47663 = ~n47650 & n47656;
  assign n47664 = n47637 & n47643;
  assign n47665 = n47663 & n47664;
  assign n47666 = n47637 & ~n47643;
  assign n47667 = ~n47631 & n47666;
  assign n47668 = n47656 & n47667;
  assign n47669 = n47650 & n47668;
  assign n47670 = ~n47665 & ~n47669;
  assign n47671 = ~n47662 & n47670;
  assign n47672 = ~n47659 & n47671;
  assign n47673 = n47631 & ~n47650;
  assign n47674 = n47643 & n47673;
  assign n47675 = n47637 & n47674;
  assign n47676 = n47672 & ~n47675;
  assign n47677 = n47625 & ~n47676;
  assign n47678 = ~n47631 & n47637;
  assign n47679 = n47643 & n47678;
  assign n47680 = n47650 & n47679;
  assign n47681 = ~n47661 & ~n47680;
  assign n47682 = n47631 & n47644;
  assign n47683 = n47650 & n47682;
  assign n47684 = n47681 & ~n47683;
  assign n47685 = ~n47656 & ~n47684;
  assign n47686 = n47631 & ~n47643;
  assign n47687 = n47637 & n47686;
  assign n47688 = ~n47656 & n47687;
  assign n47689 = n47650 & n47688;
  assign n47690 = ~n47637 & n47660;
  assign n47691 = ~n47637 & ~n47643;
  assign n47692 = ~n47650 & n47691;
  assign n47693 = ~n47690 & ~n47692;
  assign n47694 = ~n47656 & ~n47693;
  assign n47695 = ~n47689 & ~n47694;
  assign n47696 = n47625 & ~n47695;
  assign n47697 = ~n47685 & ~n47696;
  assign n47698 = ~n47677 & n47697;
  assign n47699 = n47631 & n47650;
  assign n47700 = n47691 & n47699;
  assign n47701 = n47656 & n47700;
  assign n47702 = n47631 & n47663;
  assign n47703 = n47637 & n47702;
  assign n47704 = ~n47656 & n47678;
  assign n47705 = ~n47637 & n47650;
  assign n47706 = n47631 & n47705;
  assign n47707 = ~n47682 & ~n47706;
  assign n47708 = ~n47704 & n47707;
  assign n47709 = ~n47650 & n47687;
  assign n47710 = n47708 & ~n47709;
  assign n47711 = n47644 & n47656;
  assign n47712 = ~n47650 & n47711;
  assign n47713 = n47631 & n47643;
  assign n47714 = n47650 & n47691;
  assign n47715 = ~n47713 & ~n47714;
  assign n47716 = n47656 & ~n47715;
  assign n47717 = ~n47712 & ~n47716;
  assign n47718 = n47710 & n47717;
  assign n47719 = ~n47625 & ~n47718;
  assign n47720 = ~n47703 & ~n47719;
  assign n47721 = ~n47701 & n47720;
  assign n47722 = n47698 & n47721;
  assign n47723 = pi1253 & n47722;
  assign n47724 = ~pi1253 & ~n47722;
  assign po1339 = n47723 | n47724;
  assign n47726 = pi4104 & pi9040;
  assign n47727 = pi4038 & ~pi9040;
  assign n47728 = ~n47726 & ~n47727;
  assign n47729 = ~pi1209 & ~n47728;
  assign n47730 = pi1209 & n47728;
  assign n47731 = ~n47729 & ~n47730;
  assign n47732 = pi4123 & pi9040;
  assign n47733 = pi4111 & ~pi9040;
  assign n47734 = ~n47732 & ~n47733;
  assign n47735 = ~pi1200 & ~n47734;
  assign n47736 = pi1200 & n47734;
  assign n47737 = ~n47735 & ~n47736;
  assign n47738 = pi4298 & ~pi9040;
  assign n47739 = pi4375 & pi9040;
  assign n47740 = ~n47738 & ~n47739;
  assign n47741 = ~pi1241 & ~n47740;
  assign n47742 = pi1241 & n47740;
  assign n47743 = ~n47741 & ~n47742;
  assign n47744 = pi4098 & ~pi9040;
  assign n47745 = pi4114 & pi9040;
  assign n47746 = ~n47744 & ~n47745;
  assign n47747 = ~pi1236 & ~n47746;
  assign n47748 = pi1236 & n47746;
  assign n47749 = ~n47747 & ~n47748;
  assign n47750 = pi4088 & pi9040;
  assign n47751 = pi4375 & ~pi9040;
  assign n47752 = ~n47750 & ~n47751;
  assign n47753 = ~pi1210 & n47752;
  assign n47754 = pi1210 & ~n47752;
  assign n47755 = ~n47753 & ~n47754;
  assign n47756 = ~n47749 & ~n47755;
  assign n47757 = ~n47743 & n47756;
  assign n47758 = ~n47737 & n47757;
  assign n47759 = pi4207 & ~pi9040;
  assign n47760 = pi4299 & pi9040;
  assign n47761 = ~n47759 & ~n47760;
  assign n47762 = ~pi1239 & ~n47761;
  assign n47763 = pi1239 & n47761;
  assign n47764 = ~n47762 & ~n47763;
  assign n47765 = n47749 & n47755;
  assign n47766 = n47764 & n47765;
  assign n47767 = n47737 & ~n47764;
  assign n47768 = n47755 & n47767;
  assign n47769 = ~n47749 & n47768;
  assign n47770 = ~n47766 & ~n47769;
  assign n47771 = n47749 & ~n47755;
  assign n47772 = n47737 & n47771;
  assign n47773 = n47770 & ~n47772;
  assign n47774 = ~n47743 & ~n47773;
  assign n47775 = n47749 & ~n47764;
  assign n47776 = ~n47737 & n47743;
  assign n47777 = n47775 & n47776;
  assign n47778 = ~n47764 & n47765;
  assign n47779 = ~n47737 & n47778;
  assign n47780 = ~n47777 & ~n47779;
  assign n47781 = ~n47774 & n47780;
  assign n47782 = ~n47758 & n47781;
  assign n47783 = n47756 & n47764;
  assign n47784 = ~n47737 & n47783;
  assign n47785 = n47764 & n47771;
  assign n47786 = n47737 & n47785;
  assign n47787 = ~n47784 & ~n47786;
  assign n47788 = n47782 & n47787;
  assign n47789 = ~n47731 & ~n47788;
  assign n47790 = ~n47737 & ~n47764;
  assign n47791 = ~n47755 & n47790;
  assign n47792 = n47749 & n47791;
  assign n47793 = ~n47783 & ~n47792;
  assign n47794 = ~n47743 & ~n47793;
  assign n47795 = n47756 & ~n47764;
  assign n47796 = n47737 & n47795;
  assign n47797 = n47755 & n47790;
  assign n47798 = ~n47749 & n47797;
  assign n47799 = ~n47796 & ~n47798;
  assign n47800 = n47749 & n47767;
  assign n47801 = ~n47737 & n47785;
  assign n47802 = ~n47800 & ~n47801;
  assign n47803 = n47743 & ~n47802;
  assign n47804 = n47799 & ~n47803;
  assign n47805 = ~n47794 & n47804;
  assign n47806 = n47731 & ~n47805;
  assign n47807 = ~n47749 & n47764;
  assign n47808 = ~n47737 & n47807;
  assign n47809 = n47749 & n47764;
  assign n47810 = n47737 & n47809;
  assign n47811 = ~n47808 & ~n47810;
  assign n47812 = ~n47743 & ~n47811;
  assign n47813 = ~n47749 & n47755;
  assign n47814 = n47764 & n47813;
  assign n47815 = n47737 & n47814;
  assign n47816 = ~n47778 & ~n47815;
  assign n47817 = ~n47796 & n47816;
  assign n47818 = n47743 & ~n47817;
  assign n47819 = ~n47812 & ~n47818;
  assign n47820 = n47755 & ~n47764;
  assign n47821 = n47743 & n47820;
  assign n47822 = ~n47737 & n47821;
  assign n47823 = n47819 & ~n47822;
  assign n47824 = ~n47806 & n47823;
  assign n47825 = ~n47789 & n47824;
  assign n47826 = pi1250 & n47825;
  assign n47827 = ~pi1250 & ~n47825;
  assign po1340 = n47826 | n47827;
  assign n47829 = pi4045 & ~pi9040;
  assign n47830 = pi4295 & pi9040;
  assign n47831 = ~n47829 & ~n47830;
  assign n47832 = ~pi1238 & n47831;
  assign n47833 = pi1238 & ~n47831;
  assign n47834 = ~n47832 & ~n47833;
  assign n47835 = pi4317 & ~pi9040;
  assign n47836 = pi4122 & pi9040;
  assign n47837 = ~n47835 & ~n47836;
  assign n47838 = ~pi1244 & n47837;
  assign n47839 = pi1244 & ~n47837;
  assign n47840 = ~n47838 & ~n47839;
  assign n47841 = pi4036 & ~pi9040;
  assign n47842 = pi4129 & pi9040;
  assign n47843 = ~n47841 & ~n47842;
  assign n47844 = ~pi1219 & n47843;
  assign n47845 = pi1219 & ~n47843;
  assign n47846 = ~n47844 & ~n47845;
  assign n47847 = pi4045 & pi9040;
  assign n47848 = pi4301 & ~pi9040;
  assign n47849 = ~n47847 & ~n47848;
  assign n47850 = ~pi1225 & n47849;
  assign n47851 = pi1225 & ~n47849;
  assign n47852 = ~n47850 & ~n47851;
  assign n47853 = pi4120 & pi9040;
  assign n47854 = pi4101 & ~pi9040;
  assign n47855 = ~n47853 & ~n47854;
  assign n47856 = ~pi1224 & n47855;
  assign n47857 = pi1224 & ~n47855;
  assign n47858 = ~n47856 & ~n47857;
  assign n47859 = n47852 & ~n47858;
  assign n47860 = ~n47846 & n47859;
  assign n47861 = ~n47840 & n47860;
  assign n47862 = n47834 & n47861;
  assign n47863 = n47834 & ~n47846;
  assign n47864 = ~n47852 & n47863;
  assign n47865 = n47858 & n47864;
  assign n47866 = n47840 & n47865;
  assign n47867 = ~n47862 & ~n47866;
  assign n47868 = ~n47834 & n47846;
  assign n47869 = n47852 & n47868;
  assign n47870 = ~n47858 & n47869;
  assign n47871 = n47852 & n47858;
  assign n47872 = n47846 & n47871;
  assign n47873 = n47834 & n47872;
  assign n47874 = ~n47870 & ~n47873;
  assign n47875 = ~n47840 & ~n47874;
  assign n47876 = n47867 & ~n47875;
  assign n47877 = ~pi4252 & pi9040;
  assign n47878 = ~pi4120 & ~pi9040;
  assign n47879 = ~n47877 & ~n47878;
  assign n47880 = ~pi1235 & n47879;
  assign n47881 = pi1235 & ~n47879;
  assign n47882 = ~n47880 & ~n47881;
  assign n47883 = ~n47861 & ~n47865;
  assign n47884 = n47834 & ~n47858;
  assign n47885 = n47846 & n47884;
  assign n47886 = n47858 & n47863;
  assign n47887 = ~n47885 & ~n47886;
  assign n47888 = n47840 & ~n47887;
  assign n47889 = ~n47834 & n47840;
  assign n47890 = n47871 & n47889;
  assign n47891 = n47846 & n47890;
  assign n47892 = ~n47852 & ~n47858;
  assign n47893 = ~n47846 & n47892;
  assign n47894 = ~n47834 & n47893;
  assign n47895 = ~n47840 & n47846;
  assign n47896 = ~n47852 & n47895;
  assign n47897 = n47858 & n47896;
  assign n47898 = ~n47894 & ~n47897;
  assign n47899 = ~n47891 & n47898;
  assign n47900 = ~n47888 & n47899;
  assign n47901 = n47883 & n47900;
  assign n47902 = n47882 & ~n47901;
  assign n47903 = n47876 & ~n47902;
  assign n47904 = ~n47834 & ~n47840;
  assign n47905 = ~n47846 & n47858;
  assign n47906 = n47904 & n47905;
  assign n47907 = ~n47840 & n47872;
  assign n47908 = ~n47906 & ~n47907;
  assign n47909 = ~n47840 & n47893;
  assign n47910 = n47846 & n47892;
  assign n47911 = n47834 & n47910;
  assign n47912 = ~n47909 & ~n47911;
  assign n47913 = ~n47846 & n47871;
  assign n47914 = ~n47834 & n47913;
  assign n47915 = ~n47873 & ~n47914;
  assign n47916 = ~n47834 & n47859;
  assign n47917 = n47846 & ~n47852;
  assign n47918 = ~n47916 & ~n47917;
  assign n47919 = n47840 & ~n47918;
  assign n47920 = n47915 & ~n47919;
  assign n47921 = n47912 & n47920;
  assign n47922 = n47908 & n47921;
  assign n47923 = ~n47882 & ~n47922;
  assign n47924 = n47903 & ~n47923;
  assign n47925 = ~pi1251 & ~n47924;
  assign n47926 = pi1251 & n47903;
  assign n47927 = ~n47923 & n47926;
  assign po1341 = n47925 | n47927;
  assign n47929 = n47305 & n47311;
  assign n47930 = ~n47465 & ~n47929;
  assign n47931 = ~n47315 & ~n47485;
  assign n47932 = n47235 & n47451;
  assign n47933 = n47248 & n47300;
  assign n47934 = ~n47235 & n47310;
  assign n47935 = ~n47933 & ~n47934;
  assign n47936 = ~n47309 & n47935;
  assign n47937 = ~n47932 & n47936;
  assign n47938 = n47931 & n47937;
  assign n47939 = ~n47459 & n47938;
  assign n47940 = n47241 & ~n47939;
  assign n47941 = n47248 & n47260;
  assign n47942 = ~n47310 & ~n47941;
  assign n47943 = ~n47280 & n47942;
  assign n47944 = n47235 & ~n47943;
  assign n47945 = ~n47235 & ~n47511;
  assign n47946 = n47248 & n47285;
  assign n47947 = ~n47945 & ~n47946;
  assign n47948 = ~n47944 & n47947;
  assign n47949 = ~n47241 & ~n47948;
  assign n47950 = ~n47940 & ~n47949;
  assign n47951 = ~n47469 & n47950;
  assign n47952 = n47930 & n47951;
  assign n47953 = pi1285 & n47952;
  assign n47954 = ~pi1285 & ~n47952;
  assign po1343 = n47953 | n47954;
  assign n47956 = ~n47532 & n47559;
  assign n47957 = n47538 & n47956;
  assign n47958 = n47544 & n47565;
  assign n47959 = n47532 & n47958;
  assign n47960 = n47532 & n47582;
  assign n47961 = ~n47959 & ~n47960;
  assign n47962 = ~n47532 & ~n47544;
  assign n47963 = ~n47550 & n47962;
  assign n47964 = ~n47538 & n47963;
  assign n47965 = ~n47574 & ~n47964;
  assign n47966 = ~n47559 & ~n47965;
  assign n47967 = n47961 & ~n47966;
  assign n47968 = ~n47957 & n47967;
  assign n47969 = n47526 & ~n47968;
  assign n47970 = n47532 & n47603;
  assign n47971 = n47559 & n47970;
  assign n47972 = ~n47532 & ~n47559;
  assign n47973 = n47603 & n47972;
  assign n47974 = ~n47573 & ~n47973;
  assign n47975 = n47544 & n47581;
  assign n47976 = ~n47574 & ~n47975;
  assign n47977 = ~n47532 & n47581;
  assign n47978 = n47976 & ~n47977;
  assign n47979 = n47559 & ~n47978;
  assign n47980 = ~n47559 & n47561;
  assign n47981 = n47586 & ~n47980;
  assign n47982 = ~n47979 & n47981;
  assign n47983 = n47974 & n47982;
  assign n47984 = ~n47526 & ~n47983;
  assign n47985 = ~n47971 & ~n47984;
  assign n47986 = ~n47969 & n47985;
  assign n47987 = n47972 & n47975;
  assign n47988 = n47532 & n47597;
  assign n47989 = ~n47987 & ~n47988;
  assign n47990 = ~n47559 & n47960;
  assign n47991 = n47989 & ~n47990;
  assign n47992 = n47986 & n47991;
  assign n47993 = ~pi1252 & ~n47992;
  assign n47994 = pi1252 & n47991;
  assign n47995 = n47985 & n47994;
  assign n47996 = ~n47969 & n47995;
  assign po1344 = n47993 | n47996;
  assign n47998 = n47737 & n47778;
  assign n47999 = ~n47798 & ~n47809;
  assign n48000 = n47743 & ~n47999;
  assign n48001 = ~n47998 & ~n48000;
  assign n48002 = ~n47792 & n48001;
  assign n48003 = n47737 & ~n47743;
  assign n48004 = n47795 & n48003;
  assign n48005 = ~n47784 & ~n48004;
  assign n48006 = ~n47815 & n48005;
  assign n48007 = n48002 & n48006;
  assign n48008 = n47731 & ~n48007;
  assign n48009 = ~n47755 & n47767;
  assign n48010 = n47749 & n48009;
  assign n48011 = ~n47769 & ~n48010;
  assign n48012 = n47743 & n47795;
  assign n48013 = n47737 & n47783;
  assign n48014 = ~n48012 & ~n48013;
  assign n48015 = ~n47737 & n47814;
  assign n48016 = ~n47779 & ~n48015;
  assign n48017 = ~n47755 & n47764;
  assign n48018 = n47737 & n47749;
  assign n48019 = ~n48017 & ~n48018;
  assign n48020 = ~n47820 & n48019;
  assign n48021 = ~n47743 & ~n48020;
  assign n48022 = n48016 & ~n48021;
  assign n48023 = n48014 & n48022;
  assign n48024 = n48011 & n48023;
  assign n48025 = ~n47731 & ~n48024;
  assign n48026 = ~n48008 & ~n48025;
  assign n48027 = pi1249 & ~n48026;
  assign n48028 = ~pi1249 & ~n48008;
  assign n48029 = ~n48025 & n48028;
  assign po1345 = n48027 | n48029;
  assign n48031 = ~n47834 & n47860;
  assign n48032 = n47834 & n47913;
  assign n48033 = ~n48031 & ~n48032;
  assign n48034 = ~n47852 & n47858;
  assign n48035 = ~n47846 & n48034;
  assign n48036 = ~n47834 & n48035;
  assign n48037 = ~n47834 & n47892;
  assign n48038 = n47846 & n48034;
  assign n48039 = n47834 & n48038;
  assign n48040 = ~n48037 & ~n48039;
  assign n48041 = n47840 & ~n48040;
  assign n48042 = ~n48036 & ~n48041;
  assign n48043 = ~n47840 & n48034;
  assign n48044 = ~n47834 & n48043;
  assign n48045 = ~n47907 & ~n48044;
  assign n48046 = n48042 & n48045;
  assign n48047 = n48033 & n48046;
  assign n48048 = n47882 & ~n48047;
  assign n48049 = n47840 & ~n47882;
  assign n48050 = n47858 & n47868;
  assign n48051 = n47846 & n47852;
  assign n48052 = ~n48050 & ~n48051;
  assign n48053 = n48049 & ~n48052;
  assign n48054 = ~n47865 & ~n47885;
  assign n48055 = ~n47846 & n47904;
  assign n48056 = ~n48034 & n48055;
  assign n48057 = ~n47861 & ~n48056;
  assign n48058 = n48054 & n48057;
  assign n48059 = ~n47882 & ~n48058;
  assign n48060 = n47846 & n47859;
  assign n48061 = n47834 & n47840;
  assign n48062 = n48060 & n48061;
  assign n48063 = n47834 & n47893;
  assign n48064 = ~n48032 & ~n48063;
  assign n48065 = n47840 & ~n48064;
  assign n48066 = ~n48062 & ~n48065;
  assign n48067 = ~n47840 & n47865;
  assign n48068 = n48066 & ~n48067;
  assign n48069 = ~n48059 & n48068;
  assign n48070 = ~n48053 & n48069;
  assign n48071 = ~n48048 & n48070;
  assign n48072 = n47834 & ~n47840;
  assign n48073 = n47910 & n48072;
  assign n48074 = n48071 & ~n48073;
  assign n48075 = ~pi1255 & ~n48074;
  assign n48076 = ~n48048 & ~n48073;
  assign n48077 = n48070 & n48076;
  assign n48078 = pi1255 & n48077;
  assign po1346 = n48075 | n48078;
  assign n48080 = pi4200 & ~pi9040;
  assign n48081 = pi4042 & pi9040;
  assign n48082 = ~n48080 & ~n48081;
  assign n48083 = ~pi1242 & n48082;
  assign n48084 = pi1242 & ~n48082;
  assign n48085 = ~n48083 & ~n48084;
  assign n48086 = pi4042 & ~pi9040;
  assign n48087 = pi4446 & pi9040;
  assign n48088 = ~n48086 & ~n48087;
  assign n48089 = ~pi1229 & ~n48088;
  assign n48090 = pi1229 & n48088;
  assign n48091 = ~n48089 & ~n48090;
  assign n48092 = pi4036 & pi9040;
  assign n48093 = pi4252 & ~pi9040;
  assign n48094 = ~n48092 & ~n48093;
  assign n48095 = ~pi1230 & n48094;
  assign n48096 = pi1230 & ~n48094;
  assign n48097 = ~n48095 & ~n48096;
  assign n48098 = n48091 & n48097;
  assign n48099 = pi4159 & ~pi9040;
  assign n48100 = pi4037 & pi9040;
  assign n48101 = ~n48099 & ~n48100;
  assign n48102 = ~pi1234 & n48101;
  assign n48103 = pi1234 & ~n48101;
  assign n48104 = ~n48102 & ~n48103;
  assign n48105 = pi4137 & pi9040;
  assign n48106 = pi4446 & ~pi9040;
  assign n48107 = ~n48105 & ~n48106;
  assign n48108 = ~pi1216 & n48107;
  assign n48109 = pi1216 & ~n48107;
  assign n48110 = ~n48108 & ~n48109;
  assign n48111 = ~n48104 & ~n48110;
  assign n48112 = n48098 & n48111;
  assign n48113 = ~n48104 & n48110;
  assign n48114 = ~n48091 & n48113;
  assign n48115 = ~n48112 & ~n48114;
  assign n48116 = n48085 & ~n48115;
  assign n48117 = pi4128 & pi9040;
  assign n48118 = pi4121 & ~pi9040;
  assign n48119 = ~n48117 & ~n48118;
  assign n48120 = ~pi1243 & ~n48119;
  assign n48121 = pi1243 & n48119;
  assign n48122 = ~n48120 & ~n48121;
  assign n48123 = ~n48085 & n48104;
  assign n48124 = n48091 & n48123;
  assign n48125 = n48098 & n48110;
  assign n48126 = n48091 & ~n48097;
  assign n48127 = ~n48110 & n48126;
  assign n48128 = ~n48125 & ~n48127;
  assign n48129 = ~n48091 & n48097;
  assign n48130 = ~n48110 & n48129;
  assign n48131 = ~n48104 & n48130;
  assign n48132 = n48128 & ~n48131;
  assign n48133 = ~n48085 & ~n48132;
  assign n48134 = ~n48124 & ~n48133;
  assign n48135 = ~n48091 & ~n48097;
  assign n48136 = n48110 & n48135;
  assign n48137 = ~n48104 & n48136;
  assign n48138 = n48134 & ~n48137;
  assign n48139 = n48104 & n48129;
  assign n48140 = ~n48091 & ~n48110;
  assign n48141 = ~n48097 & n48140;
  assign n48142 = ~n48139 & ~n48141;
  assign n48143 = n48085 & ~n48142;
  assign n48144 = n48110 & n48126;
  assign n48145 = n48104 & n48144;
  assign n48146 = ~n48143 & ~n48145;
  assign n48147 = n48138 & n48146;
  assign n48148 = n48122 & ~n48147;
  assign n48149 = ~n48116 & ~n48148;
  assign n48150 = ~n48085 & ~n48122;
  assign n48151 = ~n48142 & n48150;
  assign n48152 = n48110 & n48129;
  assign n48153 = ~n48144 & ~n48152;
  assign n48154 = ~n48104 & ~n48153;
  assign n48155 = ~n48112 & ~n48154;
  assign n48156 = ~n48122 & ~n48155;
  assign n48157 = ~n48151 & ~n48156;
  assign n48158 = n48085 & ~n48122;
  assign n48159 = n48098 & n48104;
  assign n48160 = ~n48136 & ~n48159;
  assign n48161 = n48091 & ~n48110;
  assign n48162 = n48160 & ~n48161;
  assign n48163 = n48158 & ~n48162;
  assign n48164 = n48157 & ~n48163;
  assign n48165 = n48149 & n48164;
  assign n48166 = ~pi1266 & ~n48165;
  assign n48167 = n48149 & n48157;
  assign n48168 = pi1266 & n48167;
  assign n48169 = ~n48163 & n48168;
  assign po1347 = n48166 | n48169;
  assign n48171 = n47349 & n47355;
  assign n48172 = n47337 & n48171;
  assign n48173 = n47343 & n48172;
  assign n48174 = ~n47337 & n47363;
  assign n48175 = ~n47337 & n47369;
  assign n48176 = n47343 & n48175;
  assign n48177 = ~n48174 & ~n48176;
  assign n48178 = n47343 & n47377;
  assign n48179 = ~n48171 & ~n48178;
  assign n48180 = ~n47343 & ~n47349;
  assign n48181 = ~n47355 & n48180;
  assign n48182 = n48179 & ~n48181;
  assign n48183 = n47337 & ~n48182;
  assign n48184 = ~n47367 & ~n48183;
  assign n48185 = n48177 & n48184;
  assign n48186 = ~n47402 & ~n48185;
  assign n48187 = ~n47389 & ~n47409;
  assign n48188 = ~n47419 & n48187;
  assign n48189 = ~n47337 & ~n48188;
  assign n48190 = ~n47355 & n47408;
  assign n48191 = ~n47343 & n47363;
  assign n48192 = ~n47361 & n47384;
  assign n48193 = ~n48191 & ~n48192;
  assign n48194 = n47337 & ~n48193;
  assign n48195 = ~n48190 & ~n48194;
  assign n48196 = ~n48189 & n48195;
  assign n48197 = ~n47379 & ~n47420;
  assign n48198 = n48196 & n48197;
  assign n48199 = n47402 & ~n48198;
  assign n48200 = ~n47364 & ~n47371;
  assign n48201 = ~n47337 & ~n48200;
  assign n48202 = ~n47428 & ~n48201;
  assign n48203 = ~n48199 & n48202;
  assign n48204 = ~n48186 & n48203;
  assign n48205 = ~n48173 & n48204;
  assign n48206 = pi1272 & n48205;
  assign n48207 = ~pi1272 & ~n48205;
  assign po1349 = n48206 | n48207;
  assign n48209 = pi4190 & ~pi9040;
  assign n48210 = pi4101 & pi9040;
  assign n48211 = ~n48209 & ~n48210;
  assign n48212 = ~pi1230 & n48211;
  assign n48213 = pi1230 & ~n48211;
  assign n48214 = ~n48212 & ~n48213;
  assign n48215 = pi4105 & pi9040;
  assign n48216 = pi4169 & ~pi9040;
  assign n48217 = ~n48215 & ~n48216;
  assign n48218 = ~pi1219 & ~n48217;
  assign n48219 = pi1219 & n48217;
  assign n48220 = ~n48218 & ~n48219;
  assign n48221 = pi4097 & ~pi9040;
  assign n48222 = pi4317 & pi9040;
  assign n48223 = ~n48221 & ~n48222;
  assign n48224 = ~pi1243 & n48223;
  assign n48225 = pi1243 & ~n48223;
  assign n48226 = ~n48224 & ~n48225;
  assign n48227 = ~n48220 & ~n48226;
  assign n48228 = n48214 & n48227;
  assign n48229 = n48220 & ~n48226;
  assign n48230 = ~n48214 & n48229;
  assign n48231 = ~n48228 & ~n48230;
  assign n48232 = pi4037 & ~pi9040;
  assign n48233 = pi4044 & pi9040;
  assign n48234 = ~n48232 & ~n48233;
  assign n48235 = ~pi1208 & ~n48234;
  assign n48236 = pi1208 & n48234;
  assign n48237 = ~n48235 & ~n48236;
  assign n48238 = ~n48214 & ~n48237;
  assign n48239 = n48220 & n48238;
  assign n48240 = n48231 & ~n48239;
  assign n48241 = pi4129 & ~pi9040;
  assign n48242 = pi4099 & pi9040;
  assign n48243 = ~n48241 & ~n48242;
  assign n48244 = pi1223 & n48243;
  assign n48245 = ~pi1223 & ~n48243;
  assign n48246 = ~n48244 & ~n48245;
  assign n48247 = ~pi4300 & ~pi9040;
  assign n48248 = ~pi4097 & pi9040;
  assign n48249 = ~n48247 & ~n48248;
  assign n48250 = ~pi1224 & n48249;
  assign n48251 = pi1224 & ~n48249;
  assign n48252 = ~n48250 & ~n48251;
  assign n48253 = ~n48246 & n48252;
  assign n48254 = ~n48240 & n48253;
  assign n48255 = ~n48220 & n48226;
  assign n48256 = ~n48214 & n48255;
  assign n48257 = n48237 & n48252;
  assign n48258 = n48256 & n48257;
  assign n48259 = ~n48214 & n48227;
  assign n48260 = n48246 & n48259;
  assign n48261 = n48220 & n48226;
  assign n48262 = n48237 & n48261;
  assign n48263 = n48214 & n48220;
  assign n48264 = ~n48262 & ~n48263;
  assign n48265 = n48246 & ~n48264;
  assign n48266 = ~n48260 & ~n48265;
  assign n48267 = n48252 & ~n48266;
  assign n48268 = ~n48258 & ~n48267;
  assign n48269 = n48214 & n48237;
  assign n48270 = n48220 & n48269;
  assign n48271 = n48214 & ~n48237;
  assign n48272 = ~n48220 & n48271;
  assign n48273 = n48226 & n48272;
  assign n48274 = ~n48270 & ~n48273;
  assign n48275 = n48246 & ~n48274;
  assign n48276 = n48268 & ~n48275;
  assign n48277 = n48237 & ~n48246;
  assign n48278 = n48261 & n48277;
  assign n48279 = ~n48214 & n48278;
  assign n48280 = ~n48229 & ~n48255;
  assign n48281 = n48238 & ~n48280;
  assign n48282 = n48228 & ~n48237;
  assign n48283 = ~n48281 & ~n48282;
  assign n48284 = n48214 & n48261;
  assign n48285 = ~n48237 & ~n48246;
  assign n48286 = n48284 & n48285;
  assign n48287 = n48269 & ~n48280;
  assign n48288 = ~n48214 & n48237;
  assign n48289 = ~n48220 & n48288;
  assign n48290 = ~n48226 & n48289;
  assign n48291 = ~n48287 & ~n48290;
  assign n48292 = ~n48286 & n48291;
  assign n48293 = n48283 & n48292;
  assign n48294 = ~n48279 & n48293;
  assign n48295 = ~n48237 & n48246;
  assign n48296 = ~n48214 & n48295;
  assign n48297 = n48226 & n48296;
  assign n48298 = n48294 & ~n48297;
  assign n48299 = ~n48252 & ~n48298;
  assign n48300 = n48276 & ~n48299;
  assign n48301 = ~n48254 & n48300;
  assign n48302 = ~pi1273 & ~n48301;
  assign n48303 = pi1273 & n48276;
  assign n48304 = ~n48254 & n48303;
  assign n48305 = ~n48299 & n48304;
  assign po1350 = n48302 | n48305;
  assign n48307 = ~n47756 & ~n47765;
  assign n48308 = n47743 & ~n48307;
  assign n48309 = ~n47737 & n48308;
  assign n48310 = n47737 & n47813;
  assign n48311 = ~n47786 & ~n48310;
  assign n48312 = n47743 & ~n48311;
  assign n48313 = ~n47764 & n48308;
  assign n48314 = ~n48312 & ~n48313;
  assign n48315 = ~n48309 & n48314;
  assign n48316 = ~n47731 & ~n48315;
  assign n48317 = n47764 & ~n48307;
  assign n48318 = n47737 & n48317;
  assign n48319 = ~n48010 & ~n48318;
  assign n48320 = ~n47737 & n47771;
  assign n48321 = ~n48015 & ~n48320;
  assign n48322 = n47743 & n48321;
  assign n48323 = n47737 & n47807;
  assign n48324 = ~n47749 & n47790;
  assign n48325 = n47737 & n47765;
  assign n48326 = ~n48324 & ~n48325;
  assign n48327 = ~n47743 & n48326;
  assign n48328 = ~n48317 & n48327;
  assign n48329 = ~n48323 & n48328;
  assign n48330 = ~n48322 & ~n48329;
  assign n48331 = n48319 & ~n48330;
  assign n48332 = n47731 & ~n48331;
  assign n48333 = ~n48316 & ~n48332;
  assign n48334 = ~n47743 & ~n48321;
  assign n48335 = ~n47769 & ~n48334;
  assign n48336 = ~n47731 & ~n48335;
  assign n48337 = n47743 & n47769;
  assign n48338 = ~n47743 & ~n48319;
  assign n48339 = ~n48337 & ~n48338;
  assign n48340 = ~n48336 & n48339;
  assign n48341 = n48333 & n48340;
  assign n48342 = pi1260 & n48341;
  assign n48343 = ~pi1260 & ~n48341;
  assign po1351 = n48342 | n48343;
  assign n48345 = ~n48214 & n48261;
  assign n48346 = n48246 & n48345;
  assign n48347 = ~n48237 & n48346;
  assign n48348 = n48227 & n48295;
  assign n48349 = n48214 & n48348;
  assign n48350 = ~n48347 & ~n48349;
  assign n48351 = ~n48282 & ~n48286;
  assign n48352 = ~n48226 & n48237;
  assign n48353 = ~n48214 & n48352;
  assign n48354 = ~n48262 & ~n48353;
  assign n48355 = n48246 & ~n48354;
  assign n48356 = ~n48246 & ~n48271;
  assign n48357 = ~n48280 & n48356;
  assign n48358 = n48214 & ~n48261;
  assign n48359 = n48246 & n48358;
  assign n48360 = ~n48237 & n48359;
  assign n48361 = ~n48357 & ~n48360;
  assign n48362 = ~n48355 & n48361;
  assign n48363 = n48351 & n48362;
  assign n48364 = n48252 & ~n48363;
  assign n48365 = n48350 & ~n48364;
  assign n48366 = n48230 & ~n48246;
  assign n48367 = n48237 & n48366;
  assign n48368 = ~n48246 & ~n48252;
  assign n48369 = n48271 & ~n48280;
  assign n48370 = ~n48262 & ~n48369;
  assign n48371 = ~n48259 & n48370;
  assign n48372 = n48368 & ~n48371;
  assign n48373 = n48228 & n48237;
  assign n48374 = n48214 & n48352;
  assign n48375 = n48237 & n48255;
  assign n48376 = ~n48374 & ~n48375;
  assign n48377 = ~n48237 & n48261;
  assign n48378 = ~n48256 & ~n48377;
  assign n48379 = n48376 & n48378;
  assign n48380 = n48246 & ~n48379;
  assign n48381 = ~n48373 & ~n48380;
  assign n48382 = ~n48252 & ~n48381;
  assign n48383 = ~n48372 & ~n48382;
  assign n48384 = ~n48367 & n48383;
  assign n48385 = n48365 & n48384;
  assign n48386 = pi1267 & ~n48385;
  assign n48387 = ~pi1267 & n48365;
  assign n48388 = n48384 & n48387;
  assign po1352 = n48386 | n48388;
  assign n48390 = n48085 & ~n48104;
  assign n48391 = ~n48129 & ~n48144;
  assign n48392 = n48390 & ~n48391;
  assign n48393 = n48085 & n48110;
  assign n48394 = n48129 & n48393;
  assign n48395 = ~n48392 & ~n48394;
  assign n48396 = n48122 & ~n48395;
  assign n48397 = n48104 & ~n48110;
  assign n48398 = ~n48097 & n48397;
  assign n48399 = n48091 & n48398;
  assign n48400 = ~n48161 & ~n48397;
  assign n48401 = ~n48085 & ~n48400;
  assign n48402 = n48104 & n48110;
  assign n48403 = n48097 & n48402;
  assign n48404 = n48091 & n48403;
  assign n48405 = ~n48401 & ~n48404;
  assign n48406 = ~n48399 & n48405;
  assign n48407 = n48122 & ~n48406;
  assign n48408 = ~n48396 & ~n48407;
  assign n48409 = ~n48097 & n48111;
  assign n48410 = ~n48091 & n48409;
  assign n48411 = n48104 & n48136;
  assign n48412 = ~n48410 & ~n48411;
  assign n48413 = n48085 & ~n48412;
  assign n48414 = ~n48098 & ~n48161;
  assign n48415 = ~n48104 & ~n48414;
  assign n48416 = ~n48136 & ~n48415;
  assign n48417 = n48085 & ~n48416;
  assign n48418 = ~n48097 & n48104;
  assign n48419 = n48085 & n48418;
  assign n48420 = n48110 & n48419;
  assign n48421 = n48097 & ~n48110;
  assign n48422 = ~n48136 & ~n48421;
  assign n48423 = n48104 & ~n48422;
  assign n48424 = ~n48085 & ~n48104;
  assign n48425 = n48126 & n48424;
  assign n48426 = n48110 & n48425;
  assign n48427 = ~n48423 & ~n48426;
  assign n48428 = ~n48420 & n48427;
  assign n48429 = ~n48417 & n48428;
  assign n48430 = ~n48410 & n48429;
  assign n48431 = ~n48122 & ~n48430;
  assign n48432 = ~n48104 & n48152;
  assign n48433 = n48104 & n48161;
  assign n48434 = ~n48432 & ~n48433;
  assign n48435 = ~n48085 & ~n48434;
  assign n48436 = ~n48431 & ~n48435;
  assign n48437 = ~n48413 & n48436;
  assign n48438 = n48408 & n48437;
  assign n48439 = pi1262 & n48438;
  assign n48440 = ~pi1262 & ~n48438;
  assign po1353 = n48439 | n48440;
  assign n48442 = ~n47858 & n47868;
  assign n48443 = ~n48060 & ~n48442;
  assign n48444 = ~n47840 & ~n48443;
  assign n48445 = n47834 & n48043;
  assign n48446 = ~n48444 & ~n48445;
  assign n48447 = n47840 & n47872;
  assign n48448 = n47840 & n47892;
  assign n48449 = n47834 & n48448;
  assign n48450 = ~n48447 & ~n48449;
  assign n48451 = n48446 & n48450;
  assign n48452 = ~n47858 & n47863;
  assign n48453 = ~n47873 & ~n48452;
  assign n48454 = ~n47914 & n48453;
  assign n48455 = n48451 & n48454;
  assign n48456 = ~n47882 & ~n48455;
  assign n48457 = ~n47862 & ~n47906;
  assign n48458 = ~n47865 & ~n48060;
  assign n48459 = ~n47916 & n48458;
  assign n48460 = n47840 & ~n48459;
  assign n48461 = ~n47834 & n48038;
  assign n48462 = ~n47894 & ~n48461;
  assign n48463 = ~n48073 & n48462;
  assign n48464 = ~n47840 & n47913;
  assign n48465 = n48463 & ~n48464;
  assign n48466 = ~n48460 & n48465;
  assign n48467 = n47882 & ~n48466;
  assign n48468 = ~n47873 & n48462;
  assign n48469 = n47840 & ~n48468;
  assign n48470 = ~n48467 & ~n48469;
  assign n48471 = n48457 & n48470;
  assign n48472 = ~n48456 & n48471;
  assign n48473 = pi1265 & n48472;
  assign n48474 = ~pi1265 & ~n48472;
  assign po1354 = n48473 | n48474;
  assign n48476 = ~n47343 & n48192;
  assign n48477 = n47343 & n47404;
  assign n48478 = ~n47389 & ~n48477;
  assign n48479 = n47337 & ~n48478;
  assign n48480 = ~n48476 & ~n48479;
  assign n48481 = ~n47361 & n47426;
  assign n48482 = ~n47355 & n48481;
  assign n48483 = n47365 & n47405;
  assign n48484 = ~n48482 & ~n48483;
  assign n48485 = ~n48174 & n48484;
  assign n48486 = ~n47373 & ~n47379;
  assign n48487 = n47361 & n47411;
  assign n48488 = n48486 & ~n48487;
  assign n48489 = n48485 & n48488;
  assign n48490 = n48480 & n48489;
  assign n48491 = ~n47402 & ~n48490;
  assign n48492 = ~n47372 & ~n47389;
  assign n48493 = n47343 & ~n48492;
  assign n48494 = ~n47419 & ~n48190;
  assign n48495 = ~n47349 & ~n47361;
  assign n48496 = n47343 & n48495;
  assign n48497 = n48494 & ~n48496;
  assign n48498 = n47337 & ~n48497;
  assign n48499 = ~n47343 & n47377;
  assign n48500 = n47343 & n47349;
  assign n48501 = ~n47361 & n48500;
  assign n48502 = ~n47355 & n48501;
  assign n48503 = ~n48499 & ~n48502;
  assign n48504 = ~n47337 & ~n48503;
  assign n48505 = ~n47343 & n47366;
  assign n48506 = ~n48504 & ~n48505;
  assign n48507 = ~n48498 & n48506;
  assign n48508 = ~n48493 & n48507;
  assign n48509 = n47402 & ~n48508;
  assign n48510 = n47337 & n47409;
  assign n48511 = ~n48509 & ~n48510;
  assign n48512 = ~n47337 & n48476;
  assign n48513 = n48511 & ~n48512;
  assign n48514 = ~n48491 & n48513;
  assign n48515 = ~pi1258 & ~n48514;
  assign n48516 = pi1258 & n48511;
  assign n48517 = ~n48491 & n48516;
  assign n48518 = ~n48512 & n48517;
  assign po1355 = n48515 | n48518;
  assign n48520 = n48214 & n48229;
  assign n48521 = ~n48345 & ~n48520;
  assign n48522 = n48246 & ~n48521;
  assign n48523 = ~n48237 & n48255;
  assign n48524 = ~n48230 & ~n48523;
  assign n48525 = ~n48284 & n48524;
  assign n48526 = ~n48246 & ~n48525;
  assign n48527 = ~n48522 & ~n48526;
  assign n48528 = ~n48260 & ~n48273;
  assign n48529 = n48527 & n48528;
  assign n48530 = ~n48252 & ~n48529;
  assign n48531 = n48237 & n48345;
  assign n48532 = n48227 & ~n48237;
  assign n48533 = ~n48375 & ~n48532;
  assign n48534 = ~n48246 & ~n48533;
  assign n48535 = ~n48531 & ~n48534;
  assign n48536 = ~n48214 & n48246;
  assign n48537 = ~n48220 & n48536;
  assign n48538 = n48226 & n48537;
  assign n48539 = n48231 & ~n48538;
  assign n48540 = ~n48284 & n48539;
  assign n48541 = ~n48237 & ~n48540;
  assign n48542 = n48535 & ~n48541;
  assign n48543 = n48252 & ~n48542;
  assign n48544 = ~n48530 & ~n48543;
  assign n48545 = n48214 & n48375;
  assign n48546 = ~n48290 & ~n48545;
  assign n48547 = n48246 & ~n48546;
  assign n48548 = n48214 & ~n48226;
  assign n48549 = n48277 & n48548;
  assign n48550 = ~n48547 & ~n48549;
  assign n48551 = n48544 & n48550;
  assign n48552 = ~pi1284 & ~n48551;
  assign n48553 = pi1284 & ~n48547;
  assign n48554 = n48544 & n48553;
  assign n48555 = ~n48549 & n48554;
  assign po1357 = n48552 | n48555;
  assign n48557 = ~n48256 & ~n48352;
  assign n48558 = n48253 & ~n48557;
  assign n48559 = n48246 & n48269;
  assign n48560 = n48229 & n48559;
  assign n48561 = ~n48214 & ~n48220;
  assign n48562 = n48277 & n48561;
  assign n48563 = ~n48560 & ~n48562;
  assign n48564 = ~n48229 & n48252;
  assign n48565 = n48288 & n48564;
  assign n48566 = n48563 & ~n48565;
  assign n48567 = ~n48375 & ~n48377;
  assign n48568 = n48246 & ~n48567;
  assign n48569 = ~n48349 & ~n48568;
  assign n48570 = n48252 & ~n48569;
  assign n48571 = ~n48229 & ~n48548;
  assign n48572 = ~n48237 & ~n48571;
  assign n48573 = ~n48345 & ~n48572;
  assign n48574 = ~n48246 & ~n48573;
  assign n48575 = ~n48369 & ~n48574;
  assign n48576 = n48237 & n48284;
  assign n48577 = ~n48220 & n48238;
  assign n48578 = n48237 & ~n48571;
  assign n48579 = ~n48577 & ~n48578;
  assign n48580 = n48246 & ~n48579;
  assign n48581 = ~n48576 & ~n48580;
  assign n48582 = n48575 & n48581;
  assign n48583 = ~n48252 & ~n48582;
  assign n48584 = ~n48570 & ~n48583;
  assign n48585 = n48566 & n48584;
  assign n48586 = ~n48558 & n48585;
  assign n48587 = pi1274 & ~n48586;
  assign n48588 = ~pi1274 & n48566;
  assign n48589 = ~n48558 & n48588;
  assign n48590 = n48584 & n48589;
  assign po1358 = n48587 | n48590;
  assign n48592 = ~n47631 & ~n47637;
  assign n48593 = ~n47675 & ~n48592;
  assign n48594 = ~n47705 & n48593;
  assign n48595 = n47656 & ~n48594;
  assign n48596 = n47650 & ~n47656;
  assign n48597 = n47637 & n48596;
  assign n48598 = ~n47631 & n47650;
  assign n48599 = n47643 & n48598;
  assign n48600 = ~n47650 & n47667;
  assign n48601 = ~n48599 & ~n48600;
  assign n48602 = n47631 & ~n47637;
  assign n48603 = ~n47650 & ~n47656;
  assign n48604 = n48602 & n48603;
  assign n48605 = n48601 & ~n48604;
  assign n48606 = ~n48597 & n48605;
  assign n48607 = ~n48595 & n48606;
  assign n48608 = ~n47625 & ~n48607;
  assign n48609 = ~n47631 & n47644;
  assign n48610 = ~n47650 & n48609;
  assign n48611 = ~n47631 & n47691;
  assign n48612 = n47650 & n48611;
  assign n48613 = ~n48610 & ~n48612;
  assign n48614 = n47656 & ~n48613;
  assign n48615 = ~n48608 & ~n48614;
  assign n48616 = n47650 & n47667;
  assign n48617 = ~n47679 & ~n47687;
  assign n48618 = n47656 & ~n48617;
  assign n48619 = ~n48616 & ~n48618;
  assign n48620 = ~n47683 & n48619;
  assign n48621 = n47625 & ~n48620;
  assign n48622 = ~n47664 & ~n47691;
  assign n48623 = n47631 & ~n48622;
  assign n48624 = ~n47692 & ~n48623;
  assign n48625 = ~n47656 & ~n48624;
  assign n48626 = n47625 & n48625;
  assign n48627 = ~n48621 & ~n48626;
  assign n48628 = n48615 & n48627;
  assign n48629 = pi1276 & ~n48628;
  assign n48630 = ~pi1276 & n48615;
  assign n48631 = n48627 & n48630;
  assign po1359 = n48629 | n48631;
  assign n48633 = n47349 & ~n47355;
  assign n48634 = ~n47337 & n48633;
  assign n48635 = n47343 & n48634;
  assign n48636 = ~n47343 & n48495;
  assign n48637 = ~n47364 & ~n48636;
  assign n48638 = ~n48502 & n48637;
  assign n48639 = ~n48635 & n48638;
  assign n48640 = n47337 & n47372;
  assign n48641 = n48639 & ~n48640;
  assign n48642 = n47402 & ~n48641;
  assign n48643 = ~n47420 & ~n48505;
  assign n48644 = n47337 & ~n48643;
  assign n48645 = ~n47337 & ~n47402;
  assign n48646 = n47404 & n48645;
  assign n48647 = n47355 & n48180;
  assign n48648 = ~n48495 & ~n48647;
  assign n48649 = ~n47366 & n48648;
  assign n48650 = n47337 & ~n48649;
  assign n48651 = ~n47343 & n47378;
  assign n48652 = ~n48650 & ~n48651;
  assign n48653 = ~n47402 & ~n48652;
  assign n48654 = ~n48646 & ~n48653;
  assign n48655 = ~n48644 & n48654;
  assign n48656 = ~n47343 & n47419;
  assign n48657 = ~n48477 & ~n48656;
  assign n48658 = ~n47373 & n48657;
  assign n48659 = ~n47364 & n48658;
  assign n48660 = ~n47337 & ~n48659;
  assign n48661 = n48655 & ~n48660;
  assign n48662 = ~n48642 & n48661;
  assign n48663 = ~pi1270 & ~n48662;
  assign n48664 = pi1270 & n48655;
  assign n48665 = ~n48642 & n48664;
  assign n48666 = ~n48660 & n48665;
  assign po1360 = n48663 | n48666;
  assign n48668 = ~n48031 & ~n48050;
  assign n48669 = n47882 & ~n48668;
  assign n48670 = ~n47864 & ~n47886;
  assign n48671 = ~n48035 & n48670;
  assign n48672 = n47840 & ~n48671;
  assign n48673 = n47882 & n48672;
  assign n48674 = ~n48669 & ~n48673;
  assign n48675 = n47860 & n47889;
  assign n48676 = ~n47891 & ~n48675;
  assign n48677 = ~n47885 & ~n47917;
  assign n48678 = ~n47840 & ~n48677;
  assign n48679 = n47882 & n48678;
  assign n48680 = n48676 & ~n48679;
  assign n48681 = ~n47846 & ~n47858;
  assign n48682 = n47852 & n48681;
  assign n48683 = n47834 & n48682;
  assign n48684 = n47834 & n47871;
  assign n48685 = ~n47870 & ~n48684;
  assign n48686 = ~n47840 & ~n48685;
  assign n48687 = ~n47865 & ~n47894;
  assign n48688 = n47834 & n47859;
  assign n48689 = ~n47910 & ~n48688;
  assign n48690 = n47840 & ~n48689;
  assign n48691 = n48687 & ~n48690;
  assign n48692 = ~n48686 & n48691;
  assign n48693 = ~n48683 & n48692;
  assign n48694 = ~n47882 & ~n48693;
  assign n48695 = ~n47914 & n48462;
  assign n48696 = ~n47840 & ~n48695;
  assign n48697 = ~n48694 & ~n48696;
  assign n48698 = n48680 & n48697;
  assign n48699 = n48674 & n48698;
  assign n48700 = ~pi1264 & ~n48699;
  assign n48701 = pi1264 & n48680;
  assign n48702 = n48674 & n48701;
  assign n48703 = n48697 & n48702;
  assign po1361 = n48700 | n48703;
  assign n48705 = ~n47532 & n47958;
  assign n48706 = n47532 & n47560;
  assign n48707 = ~n47573 & ~n48706;
  assign n48708 = ~n47584 & n48707;
  assign n48709 = ~n47559 & ~n48708;
  assign n48710 = ~n47582 & ~n47590;
  assign n48711 = n47532 & n47551;
  assign n48712 = ~n47532 & n47603;
  assign n48713 = ~n48711 & ~n48712;
  assign n48714 = n48710 & n48713;
  assign n48715 = n47559 & ~n48714;
  assign n48716 = n47550 & n47591;
  assign n48717 = n47538 & n48716;
  assign n48718 = ~n48715 & ~n48717;
  assign n48719 = ~n48709 & n48718;
  assign n48720 = ~n48705 & n48719;
  assign n48721 = ~n47526 & ~n48720;
  assign n48722 = ~n47532 & n47552;
  assign n48723 = ~n47585 & ~n48722;
  assign n48724 = ~n47559 & ~n48723;
  assign n48725 = n47559 & ~n47961;
  assign n48726 = ~n48724 & ~n48725;
  assign n48727 = n47532 & n47559;
  assign n48728 = n47561 & n48727;
  assign n48729 = n47559 & n47584;
  assign n48730 = n47559 & n47975;
  assign n48731 = ~n48729 & ~n48730;
  assign n48732 = ~n47532 & ~n48731;
  assign n48733 = ~n48728 & ~n48732;
  assign n48734 = ~n47970 & ~n48722;
  assign n48735 = n47532 & n47581;
  assign n48736 = ~n47532 & n47560;
  assign n48737 = ~n48735 & ~n48736;
  assign n48738 = ~n47552 & ~n47582;
  assign n48739 = n48737 & n48738;
  assign n48740 = ~n47559 & ~n48739;
  assign n48741 = ~n47532 & n47574;
  assign n48742 = ~n48740 & ~n48741;
  assign n48743 = n48734 & n48742;
  assign n48744 = n48733 & n48743;
  assign n48745 = n47526 & ~n48744;
  assign n48746 = n48726 & ~n48745;
  assign n48747 = ~n48721 & n48746;
  assign n48748 = pi1269 & ~n48747;
  assign n48749 = ~pi1269 & n48747;
  assign po1362 = n48748 | n48749;
  assign n48751 = n47743 & n47796;
  assign n48752 = n47790 & ~n48307;
  assign n48753 = ~n47814 & ~n48752;
  assign n48754 = ~n48010 & n48753;
  assign n48755 = ~n47743 & ~n48754;
  assign n48756 = n47737 & n47766;
  assign n48757 = ~n48755 & ~n48756;
  assign n48758 = ~n47764 & n47813;
  assign n48759 = ~n47737 & n48017;
  assign n48760 = ~n48758 & ~n48759;
  assign n48761 = ~n48325 & n48760;
  assign n48762 = n47743 & ~n48761;
  assign n48763 = n48757 & ~n48762;
  assign n48764 = n47731 & ~n48763;
  assign n48765 = ~n48751 & ~n48764;
  assign n48766 = ~n47737 & n47765;
  assign n48767 = ~n47764 & n47771;
  assign n48768 = ~n48766 & ~n48767;
  assign n48769 = n47743 & ~n48768;
  assign n48770 = ~n47815 & ~n48769;
  assign n48771 = ~n47786 & ~n47796;
  assign n48772 = n47737 & n47820;
  assign n48773 = ~n48017 & ~n48772;
  assign n48774 = ~n48758 & n48773;
  assign n48775 = ~n47743 & ~n48774;
  assign n48776 = ~n47737 & n47766;
  assign n48777 = ~n48775 & ~n48776;
  assign n48778 = n48771 & n48777;
  assign n48779 = n48770 & n48778;
  assign n48780 = ~n47731 & ~n48779;
  assign n48781 = ~n47801 & ~n48323;
  assign n48782 = ~n47743 & ~n48781;
  assign n48783 = ~n48780 & ~n48782;
  assign n48784 = n48765 & n48783;
  assign n48785 = pi1257 & n48784;
  assign n48786 = ~pi1257 & ~n48784;
  assign po1363 = n48785 | n48786;
  assign n48788 = n47650 & n48623;
  assign n48789 = ~n47643 & n48598;
  assign n48790 = ~n47713 & ~n48789;
  assign n48791 = ~n48611 & n48790;
  assign n48792 = n47656 & ~n48791;
  assign n48793 = ~n47686 & ~n48609;
  assign n48794 = ~n47656 & ~n48793;
  assign n48795 = ~n48792 & ~n48794;
  assign n48796 = ~n48788 & n48795;
  assign n48797 = ~n47650 & n47679;
  assign n48798 = n48796 & ~n48797;
  assign n48799 = n47625 & ~n48798;
  assign n48800 = ~n47682 & ~n47687;
  assign n48801 = ~n47679 & ~n48611;
  assign n48802 = n48800 & n48801;
  assign n48803 = n47650 & ~n48802;
  assign n48804 = n47663 & ~n48793;
  assign n48805 = ~n48803 & ~n48804;
  assign n48806 = ~n48600 & n48805;
  assign n48807 = ~n47625 & ~n48806;
  assign n48808 = ~n48799 & ~n48807;
  assign n48809 = n47650 & n48609;
  assign n48810 = ~n48797 & ~n48809;
  assign n48811 = ~n47656 & ~n48810;
  assign n48812 = n48808 & ~n48811;
  assign n48813 = pi1283 & ~n48812;
  assign n48814 = ~pi1283 & ~n48811;
  assign n48815 = ~n48807 & n48814;
  assign n48816 = ~n48799 & n48815;
  assign po1364 = n48813 | n48816;
  assign n48818 = n48097 & ~n48104;
  assign n48819 = n48110 & n48818;
  assign n48820 = ~n48144 & ~n48819;
  assign n48821 = n48085 & ~n48820;
  assign n48822 = ~n48104 & n48135;
  assign n48823 = ~n48403 & ~n48822;
  assign n48824 = ~n48085 & ~n48823;
  assign n48825 = n48104 & n48130;
  assign n48826 = ~n48420 & ~n48825;
  assign n48827 = ~n48112 & n48826;
  assign n48828 = ~n48824 & n48827;
  assign n48829 = ~n48821 & n48828;
  assign n48830 = ~n48399 & ~n48410;
  assign n48831 = n48829 & n48830;
  assign n48832 = n48122 & ~n48831;
  assign n48833 = n48098 & n48397;
  assign n48834 = n48153 & ~n48833;
  assign n48835 = ~n48085 & ~n48834;
  assign n48836 = n48104 & n48141;
  assign n48837 = ~n48835 & ~n48836;
  assign n48838 = n48091 & n48113;
  assign n48839 = ~n48104 & n48126;
  assign n48840 = ~n48838 & ~n48839;
  assign n48841 = ~n48085 & ~n48840;
  assign n48842 = ~n48085 & n48135;
  assign n48843 = n48104 & n48842;
  assign n48844 = ~n48841 & ~n48843;
  assign n48845 = n48837 & n48844;
  assign n48846 = ~n48122 & ~n48845;
  assign n48847 = ~n48130 & ~n48137;
  assign n48848 = ~n48404 & n48847;
  assign n48849 = n48158 & ~n48848;
  assign n48850 = ~n48846 & ~n48849;
  assign n48851 = ~n48112 & ~n48399;
  assign n48852 = n48085 & ~n48851;
  assign n48853 = n48850 & ~n48852;
  assign n48854 = ~n48832 & n48853;
  assign n48855 = ~pi1278 & n48854;
  assign n48856 = pi1278 & ~n48854;
  assign po1366 = n48855 | n48856;
  assign n48858 = ~n47650 & n47686;
  assign n48859 = n47650 & n47664;
  assign n48860 = ~n47678 & ~n48859;
  assign n48861 = ~n47656 & ~n48860;
  assign n48862 = n47656 & n48611;
  assign n48863 = n47650 & n47711;
  assign n48864 = ~n48599 & ~n48863;
  assign n48865 = ~n48862 & n48864;
  assign n48866 = ~n48861 & n48865;
  assign n48867 = ~n48858 & n48866;
  assign n48868 = n47625 & ~n48867;
  assign n48869 = ~n47625 & ~n47656;
  assign n48870 = n47650 & n47687;
  assign n48871 = ~n47682 & ~n48870;
  assign n48872 = ~n48611 & n48871;
  assign n48873 = n48869 & ~n48872;
  assign n48874 = ~n47675 & ~n47701;
  assign n48875 = n47656 & n48609;
  assign n48876 = ~n47669 & ~n48875;
  assign n48877 = n48874 & n48876;
  assign n48878 = ~n47625 & ~n48877;
  assign n48879 = ~n48873 & ~n48878;
  assign n48880 = n47679 & n48596;
  assign n48881 = ~n47650 & n47682;
  assign n48882 = ~n48600 & ~n48881;
  assign n48883 = ~n47656 & ~n48882;
  assign n48884 = ~n48880 & ~n48883;
  assign n48885 = ~n47703 & n48884;
  assign n48886 = ~n47650 & n48862;
  assign n48887 = n48885 & ~n48886;
  assign n48888 = n48879 & n48887;
  assign n48889 = ~n48868 & n48888;
  assign n48890 = ~pi1286 & n48889;
  assign n48891 = pi1286 & ~n48889;
  assign po1367 = n48890 | n48891;
  assign n48893 = ~n47964 & ~n48722;
  assign n48894 = ~n48717 & n48893;
  assign n48895 = n47559 & ~n48894;
  assign n48896 = ~n47973 & ~n47990;
  assign n48897 = ~n47970 & ~n48730;
  assign n48898 = ~n47958 & ~n48736;
  assign n48899 = ~n47559 & ~n48898;
  assign n48900 = ~n47590 & ~n48899;
  assign n48901 = n48897 & n48900;
  assign n48902 = n47526 & ~n48901;
  assign n48903 = ~n47544 & n47550;
  assign n48904 = ~n47562 & ~n48903;
  assign n48905 = n47532 & ~n48904;
  assign n48906 = ~n47552 & ~n47977;
  assign n48907 = ~n47559 & ~n48906;
  assign n48908 = n47532 & n47550;
  assign n48909 = ~n47574 & ~n48908;
  assign n48910 = ~n47565 & n48909;
  assign n48911 = n47559 & ~n48910;
  assign n48912 = ~n48907 & ~n48911;
  assign n48913 = ~n48905 & n48912;
  assign n48914 = ~n47526 & ~n48913;
  assign n48915 = ~n48902 & ~n48914;
  assign n48916 = n48896 & n48915;
  assign n48917 = ~n48895 & n48916;
  assign n48918 = ~pi1282 & ~n48917;
  assign n48919 = pi1282 & n48896;
  assign n48920 = ~n48895 & n48919;
  assign n48921 = n48915 & n48920;
  assign po1368 = n48918 | n48921;
  assign n48923 = n48085 & n48141;
  assign n48924 = n48104 & n48126;
  assign n48925 = ~n48125 & ~n48924;
  assign n48926 = n48085 & ~n48925;
  assign n48927 = ~n48085 & ~n48422;
  assign n48928 = ~n48926 & ~n48927;
  assign n48929 = ~n48432 & n48928;
  assign n48930 = n48122 & ~n48929;
  assign n48931 = ~n48923 & ~n48930;
  assign n48932 = ~n48110 & n48390;
  assign n48933 = ~n48402 & ~n48932;
  assign n48934 = ~n48091 & ~n48933;
  assign n48935 = ~n48112 & ~n48934;
  assign n48936 = ~n48403 & n48935;
  assign n48937 = ~n48085 & n48127;
  assign n48938 = ~n48104 & n48144;
  assign n48939 = ~n48937 & ~n48938;
  assign n48940 = n48936 & n48939;
  assign n48941 = ~n48122 & ~n48940;
  assign n48942 = ~n48825 & ~n48839;
  assign n48943 = ~n48085 & ~n48942;
  assign n48944 = ~n48941 & ~n48943;
  assign n48945 = n48931 & n48944;
  assign n48946 = ~pi1292 & ~n48945;
  assign n48947 = pi1292 & n48944;
  assign n48948 = ~n48930 & n48947;
  assign n48949 = ~n48923 & n48948;
  assign po1369 = n48946 | n48949;
  assign n48951 = pi4379 & pi9040;
  assign n48952 = pi4306 & ~pi9040;
  assign n48953 = ~n48951 & ~n48952;
  assign n48954 = ~pi1310 & ~n48953;
  assign n48955 = pi1310 & n48953;
  assign n48956 = ~n48954 & ~n48955;
  assign n48957 = pi4491 & pi9040;
  assign n48958 = pi4292 & ~pi9040;
  assign n48959 = ~n48957 & ~n48958;
  assign n48960 = ~pi1302 & n48959;
  assign n48961 = pi1302 & ~n48959;
  assign n48962 = ~n48960 & ~n48961;
  assign n48963 = pi4505 & pi9040;
  assign n48964 = pi4214 & ~pi9040;
  assign n48965 = ~n48963 & ~n48964;
  assign n48966 = pi1307 & n48965;
  assign n48967 = ~pi1307 & ~n48965;
  assign n48968 = ~n48966 & ~n48967;
  assign n48969 = pi4303 & pi9040;
  assign n48970 = pi4309 & ~pi9040;
  assign n48971 = ~n48969 & ~n48970;
  assign n48972 = ~pi1271 & ~n48971;
  assign n48973 = pi1271 & n48971;
  assign n48974 = ~n48972 & ~n48973;
  assign n48975 = pi4308 & ~pi9040;
  assign n48976 = pi4302 & pi9040;
  assign n48977 = ~n48975 & ~n48976;
  assign n48978 = ~pi1306 & n48977;
  assign n48979 = pi1306 & ~n48977;
  assign n48980 = ~n48978 & ~n48979;
  assign n48981 = ~n48974 & ~n48980;
  assign n48982 = n48968 & n48981;
  assign n48983 = ~n48962 & n48982;
  assign n48984 = pi4491 & ~pi9040;
  assign n48985 = pi4306 & pi9040;
  assign n48986 = ~n48984 & ~n48985;
  assign n48987 = pi1288 & n48986;
  assign n48988 = ~pi1288 & ~n48986;
  assign n48989 = ~n48987 & ~n48988;
  assign n48990 = n48974 & ~n48980;
  assign n48991 = ~n48962 & n48990;
  assign n48992 = ~n48968 & n48981;
  assign n48993 = n48962 & n48992;
  assign n48994 = ~n48991 & ~n48993;
  assign n48995 = ~n48989 & ~n48994;
  assign n48996 = ~n48983 & ~n48995;
  assign n48997 = ~n48974 & n48980;
  assign n48998 = ~n48968 & n48997;
  assign n48999 = n48989 & n48998;
  assign n49000 = n48981 & n48989;
  assign n49001 = ~n48962 & n49000;
  assign n49002 = ~n48999 & ~n49001;
  assign n49003 = n48996 & n49002;
  assign n49004 = n48974 & n48980;
  assign n49005 = n48968 & n49004;
  assign n49006 = ~n48962 & n49005;
  assign n49007 = n48968 & n48997;
  assign n49008 = n48962 & n49007;
  assign n49009 = ~n49006 & ~n49008;
  assign n49010 = n49003 & n49009;
  assign n49011 = n48956 & ~n49010;
  assign n49012 = ~n48956 & ~n48989;
  assign n49013 = ~n48962 & ~n48968;
  assign n49014 = ~n48974 & n49013;
  assign n49015 = ~n48968 & n48980;
  assign n49016 = ~n49014 & ~n49015;
  assign n49017 = n49012 & ~n49016;
  assign n49018 = n48962 & n48968;
  assign n49019 = ~n48980 & n49018;
  assign n49020 = ~n48974 & n49019;
  assign n49021 = n48962 & n48974;
  assign n49022 = ~n48968 & n49021;
  assign n49023 = ~n49020 & ~n49022;
  assign n49024 = ~n48962 & n48989;
  assign n49025 = n48968 & n49024;
  assign n49026 = ~n48981 & n49025;
  assign n49027 = n48989 & n49005;
  assign n49028 = ~n49026 & ~n49027;
  assign n49029 = n49023 & n49028;
  assign n49030 = ~n48956 & ~n49029;
  assign n49031 = ~n48968 & n49004;
  assign n49032 = n48962 & ~n48989;
  assign n49033 = n49031 & n49032;
  assign n49034 = n48968 & n48990;
  assign n49035 = n48962 & n49034;
  assign n49036 = ~n49008 & ~n49035;
  assign n49037 = ~n48989 & ~n49036;
  assign n49038 = ~n49033 & ~n49037;
  assign n49039 = n48989 & n49020;
  assign n49040 = n49038 & ~n49039;
  assign n49041 = ~n49030 & n49040;
  assign n49042 = ~n49017 & n49041;
  assign n49043 = ~n49011 & n49042;
  assign n49044 = ~n48968 & n48990;
  assign n49045 = n48962 & n48989;
  assign n49046 = n49044 & n49045;
  assign n49047 = n49043 & ~n49046;
  assign n49048 = ~pi1318 & ~n49047;
  assign n49049 = ~n49011 & ~n49046;
  assign n49050 = n49042 & n49049;
  assign n49051 = pi1318 & n49050;
  assign po1386 = n49048 | n49051;
  assign n49053 = n48962 & n48998;
  assign n49054 = n48980 & n49013;
  assign n49055 = n48974 & n49054;
  assign n49056 = ~n49053 & ~n49055;
  assign n49057 = n48989 & ~n49056;
  assign n49058 = ~n49020 & ~n49027;
  assign n49059 = ~n48974 & n49018;
  assign n49060 = ~n49022 & ~n49059;
  assign n49061 = ~n48989 & ~n49060;
  assign n49062 = ~n48962 & ~n48989;
  assign n49063 = n48997 & n49062;
  assign n49064 = ~n48968 & n49063;
  assign n49065 = ~n48962 & n48968;
  assign n49066 = ~n48980 & n49065;
  assign n49067 = n48974 & n49066;
  assign n49068 = ~n48968 & n48989;
  assign n49069 = ~n48980 & n49068;
  assign n49070 = ~n48974 & n49069;
  assign n49071 = ~n49067 & ~n49070;
  assign n49072 = ~n49064 & n49071;
  assign n49073 = ~n49061 & n49072;
  assign n49074 = n49058 & n49073;
  assign n49075 = n48956 & ~n49074;
  assign n49076 = ~n48989 & n49020;
  assign n49077 = n48962 & n49027;
  assign n49078 = ~n49076 & ~n49077;
  assign n49079 = ~n49075 & n49078;
  assign n49080 = ~n49057 & n49079;
  assign n49081 = n48968 & ~n48974;
  assign n49082 = n49024 & n49081;
  assign n49083 = ~n48999 & ~n49082;
  assign n49084 = n48989 & n49034;
  assign n49085 = n48962 & n49044;
  assign n49086 = ~n49084 & ~n49085;
  assign n49087 = ~n48962 & n49007;
  assign n49088 = ~n49053 & ~n49087;
  assign n49089 = ~n48962 & n49004;
  assign n49090 = ~n48968 & ~n48980;
  assign n49091 = ~n49089 & ~n49090;
  assign n49092 = ~n48989 & ~n49091;
  assign n49093 = n49088 & ~n49092;
  assign n49094 = n49086 & n49093;
  assign n49095 = n49083 & n49094;
  assign n49096 = ~n48956 & ~n49095;
  assign n49097 = n49080 & ~n49096;
  assign n49098 = ~pi1317 & ~n49097;
  assign n49099 = pi1317 & n49080;
  assign n49100 = ~n49096 & n49099;
  assign po1392 = n49098 | n49100;
  assign n49102 = ~n49077 & ~n49082;
  assign n49103 = ~n48962 & n48992;
  assign n49104 = ~n49067 & ~n49103;
  assign n49105 = ~n49053 & n49104;
  assign n49106 = ~n48989 & ~n49105;
  assign n49107 = n48974 & n49018;
  assign n49108 = ~n49087 & ~n49107;
  assign n49109 = n48990 & n49032;
  assign n49110 = ~n48989 & n48998;
  assign n49111 = ~n49109 & ~n49110;
  assign n49112 = n48962 & n49000;
  assign n49113 = n48974 & n49013;
  assign n49114 = ~n49031 & ~n49113;
  assign n49115 = n48989 & ~n49114;
  assign n49116 = ~n49112 & ~n49115;
  assign n49117 = n49111 & n49116;
  assign n49118 = n49108 & n49117;
  assign n49119 = ~n49053 & n49118;
  assign n49120 = ~n48956 & ~n49119;
  assign n49121 = ~n49020 & ~n49031;
  assign n49122 = ~n49089 & n49121;
  assign n49123 = ~n48989 & ~n49122;
  assign n49124 = ~n49046 & n49104;
  assign n49125 = n48989 & n49007;
  assign n49126 = n49124 & ~n49125;
  assign n49127 = ~n49123 & n49126;
  assign n49128 = n48956 & ~n49127;
  assign n49129 = ~n49120 & ~n49128;
  assign n49130 = ~n49106 & n49129;
  assign n49131 = n49102 & n49130;
  assign n49132 = pi1320 & ~n49131;
  assign n49133 = ~pi1320 & n49131;
  assign po1394 = n49132 | n49133;
  assign n49135 = pi4292 & pi9040;
  assign n49136 = pi4379 & ~pi9040;
  assign n49137 = ~n49135 & ~n49136;
  assign n49138 = ~pi1294 & ~n49137;
  assign n49139 = pi1294 & n49137;
  assign n49140 = ~n49138 & ~n49139;
  assign n49141 = pi4249 & ~pi9040;
  assign n49142 = pi4493 & pi9040;
  assign n49143 = ~n49141 & ~n49142;
  assign n49144 = ~pi1296 & ~n49143;
  assign n49145 = pi1296 & n49143;
  assign n49146 = ~n49144 & ~n49145;
  assign n49147 = pi4249 & pi9040;
  assign n49148 = pi4215 & ~pi9040;
  assign n49149 = ~n49147 & ~n49148;
  assign n49150 = ~pi1309 & ~n49149;
  assign n49151 = pi1309 & n49149;
  assign n49152 = ~n49150 & ~n49151;
  assign n49153 = n49146 & ~n49152;
  assign n49154 = pi4404 & pi9040;
  assign n49155 = pi4297 & ~pi9040;
  assign n49156 = ~n49154 & ~n49155;
  assign n49157 = ~pi1304 & ~n49156;
  assign n49158 = pi1304 & n49156;
  assign n49159 = ~n49157 & ~n49158;
  assign n49160 = pi4246 & pi9040;
  assign n49161 = pi4505 & ~pi9040;
  assign n49162 = ~n49160 & ~n49161;
  assign n49163 = ~pi1259 & ~n49162;
  assign n49164 = pi1259 & n49162;
  assign n49165 = ~n49163 & ~n49164;
  assign n49166 = n49159 & n49165;
  assign n49167 = n49153 & n49166;
  assign n49168 = n49159 & ~n49165;
  assign n49169 = ~n49146 & n49168;
  assign n49170 = ~n49167 & ~n49169;
  assign n49171 = ~n49140 & ~n49170;
  assign n49172 = pi4211 & pi9040;
  assign n49173 = pi4246 & ~pi9040;
  assign n49174 = ~n49172 & ~n49173;
  assign n49175 = ~pi1291 & ~n49174;
  assign n49176 = pi1291 & n49174;
  assign n49177 = ~n49175 & ~n49176;
  assign n49178 = n49140 & ~n49159;
  assign n49179 = n49146 & n49178;
  assign n49180 = n49153 & ~n49165;
  assign n49181 = n49146 & n49152;
  assign n49182 = n49165 & n49181;
  assign n49183 = ~n49180 & ~n49182;
  assign n49184 = ~n49146 & ~n49152;
  assign n49185 = n49165 & n49184;
  assign n49186 = n49159 & n49185;
  assign n49187 = n49183 & ~n49186;
  assign n49188 = n49140 & ~n49187;
  assign n49189 = ~n49179 & ~n49188;
  assign n49190 = ~n49146 & n49152;
  assign n49191 = ~n49165 & n49190;
  assign n49192 = n49159 & n49191;
  assign n49193 = n49189 & ~n49192;
  assign n49194 = ~n49159 & n49184;
  assign n49195 = ~n49146 & n49165;
  assign n49196 = n49152 & n49195;
  assign n49197 = ~n49194 & ~n49196;
  assign n49198 = ~n49140 & ~n49197;
  assign n49199 = ~n49165 & n49181;
  assign n49200 = ~n49159 & n49199;
  assign n49201 = ~n49198 & ~n49200;
  assign n49202 = n49193 & n49201;
  assign n49203 = n49177 & ~n49202;
  assign n49204 = ~n49171 & ~n49203;
  assign n49205 = n49140 & ~n49177;
  assign n49206 = ~n49197 & n49205;
  assign n49207 = ~n49165 & n49184;
  assign n49208 = ~n49199 & ~n49207;
  assign n49209 = n49159 & ~n49208;
  assign n49210 = ~n49167 & ~n49209;
  assign n49211 = ~n49177 & ~n49210;
  assign n49212 = ~n49206 & ~n49211;
  assign n49213 = ~n49140 & ~n49177;
  assign n49214 = n49153 & ~n49159;
  assign n49215 = ~n49191 & ~n49214;
  assign n49216 = n49146 & n49165;
  assign n49217 = n49215 & ~n49216;
  assign n49218 = n49213 & ~n49217;
  assign n49219 = n49212 & ~n49218;
  assign n49220 = n49204 & n49219;
  assign n49221 = ~pi1319 & ~n49220;
  assign n49222 = pi1319 & n49212;
  assign n49223 = n49204 & n49222;
  assign n49224 = ~n49218 & n49223;
  assign po1395 = n49221 | n49224;
  assign n49226 = pi4285 & pi9040;
  assign n49227 = pi4593 & ~pi9040;
  assign n49228 = ~n49226 & ~n49227;
  assign n49229 = ~pi1303 & n49228;
  assign n49230 = pi1303 & ~n49228;
  assign n49231 = ~n49229 & ~n49230;
  assign n49232 = pi4311 & ~pi9040;
  assign n49233 = pi4391 & pi9040;
  assign n49234 = ~n49232 & ~n49233;
  assign n49235 = ~pi1300 & ~n49234;
  assign n49236 = pi1300 & n49234;
  assign n49237 = ~n49235 & ~n49236;
  assign n49238 = n49231 & ~n49237;
  assign n49239 = pi4588 & ~pi9040;
  assign n49240 = pi4497 & pi9040;
  assign n49241 = ~n49239 & ~n49240;
  assign n49242 = pi1268 & n49241;
  assign n49243 = ~pi1268 & ~n49241;
  assign n49244 = ~n49242 & ~n49243;
  assign n49245 = pi4284 & ~pi9040;
  assign n49246 = pi4311 & pi9040;
  assign n49247 = ~n49245 & ~n49246;
  assign n49248 = ~pi1289 & ~n49247;
  assign n49249 = pi1289 & n49247;
  assign n49250 = ~n49248 & ~n49249;
  assign n49251 = pi4588 & pi9040;
  assign n49252 = pi4316 & ~pi9040;
  assign n49253 = ~n49251 & ~n49252;
  assign n49254 = ~pi1279 & n49253;
  assign n49255 = pi1279 & ~n49253;
  assign n49256 = ~n49254 & ~n49255;
  assign n49257 = n49250 & n49256;
  assign n49258 = ~n49244 & n49257;
  assign n49259 = pi4293 & ~pi9040;
  assign n49260 = pi4484 & pi9040;
  assign n49261 = ~n49259 & ~n49260;
  assign n49262 = ~pi1280 & ~n49261;
  assign n49263 = pi1280 & n49261;
  assign n49264 = ~n49262 & ~n49263;
  assign n49265 = ~n49256 & ~n49264;
  assign n49266 = n49244 & n49250;
  assign n49267 = n49265 & n49266;
  assign n49268 = ~n49256 & n49264;
  assign n49269 = ~n49244 & n49268;
  assign n49270 = ~n49267 & ~n49269;
  assign n49271 = ~n49258 & n49270;
  assign n49272 = n49238 & ~n49271;
  assign n49273 = ~n49244 & ~n49250;
  assign n49274 = ~n49264 & n49273;
  assign n49275 = n49256 & ~n49264;
  assign n49276 = n49250 & n49275;
  assign n49277 = n49244 & n49276;
  assign n49278 = ~n49274 & ~n49277;
  assign n49279 = ~n49250 & n49265;
  assign n49280 = n49250 & n49268;
  assign n49281 = ~n49279 & ~n49280;
  assign n49282 = n49278 & n49281;
  assign n49283 = ~n49231 & ~n49282;
  assign n49284 = n49244 & ~n49250;
  assign n49285 = n49264 & n49284;
  assign n49286 = n49256 & n49285;
  assign n49287 = ~n49283 & ~n49286;
  assign n49288 = ~n49237 & ~n49287;
  assign n49289 = ~n49272 & ~n49288;
  assign n49290 = ~n49250 & n49275;
  assign n49291 = ~n49268 & ~n49275;
  assign n49292 = n49244 & ~n49291;
  assign n49293 = ~n49290 & ~n49292;
  assign n49294 = n49231 & ~n49293;
  assign n49295 = n49256 & n49264;
  assign n49296 = n49250 & n49295;
  assign n49297 = ~n49258 & ~n49296;
  assign n49298 = ~n49267 & n49297;
  assign n49299 = ~n49231 & ~n49298;
  assign n49300 = ~n49294 & ~n49299;
  assign n49301 = n49231 & ~n49244;
  assign n49302 = n49265 & n49301;
  assign n49303 = n49244 & n49290;
  assign n49304 = ~n49250 & ~n49256;
  assign n49305 = n49264 & n49304;
  assign n49306 = n49244 & n49305;
  assign n49307 = ~n49303 & ~n49306;
  assign n49308 = n49264 & n49273;
  assign n49309 = n49256 & n49308;
  assign n49310 = n49307 & ~n49309;
  assign n49311 = ~n49302 & n49310;
  assign n49312 = n49300 & n49311;
  assign n49313 = n49237 & ~n49312;
  assign n49314 = ~n49231 & ~n49244;
  assign n49315 = n49250 & n49314;
  assign n49316 = n49264 & n49315;
  assign n49317 = ~n49244 & n49279;
  assign n49318 = ~n49316 & ~n49317;
  assign n49319 = ~n49313 & n49318;
  assign n49320 = n49289 & n49319;
  assign n49321 = pi1316 & ~n49320;
  assign n49322 = ~pi1316 & n49318;
  assign n49323 = n49289 & n49322;
  assign n49324 = ~n49313 & n49323;
  assign po1396 = n49321 | n49324;
  assign n49326 = pi4398 & pi9040;
  assign n49327 = pi4205 & ~pi9040;
  assign n49328 = ~n49326 & ~n49327;
  assign n49329 = ~pi1296 & n49328;
  assign n49330 = pi1296 & ~n49328;
  assign n49331 = ~n49329 & ~n49330;
  assign n49332 = pi4215 & pi9040;
  assign n49333 = pi4373 & ~pi9040;
  assign n49334 = ~n49332 & ~n49333;
  assign n49335 = ~pi1298 & n49334;
  assign n49336 = pi1298 & ~n49334;
  assign n49337 = ~n49335 & ~n49336;
  assign n49338 = pi4214 & pi9040;
  assign n49339 = pi4211 & ~pi9040;
  assign n49340 = ~n49338 & ~n49339;
  assign n49341 = pi1299 & n49340;
  assign n49342 = ~pi1299 & ~n49340;
  assign n49343 = ~n49341 & ~n49342;
  assign n49344 = pi4213 & ~pi9040;
  assign n49345 = pi4698 & pi9040;
  assign n49346 = ~n49344 & ~n49345;
  assign n49347 = ~pi1259 & n49346;
  assign n49348 = pi1259 & ~n49346;
  assign n49349 = ~n49347 & ~n49348;
  assign n49350 = ~n49343 & ~n49349;
  assign n49351 = pi4286 & ~pi9040;
  assign n49352 = pi4310 & pi9040;
  assign n49353 = ~n49351 & ~n49352;
  assign n49354 = pi1295 & ~n49353;
  assign n49355 = ~pi1295 & n49353;
  assign n49356 = ~n49354 & ~n49355;
  assign n49357 = pi4373 & pi9040;
  assign n49358 = pi4493 & ~pi9040;
  assign n49359 = ~n49357 & ~n49358;
  assign n49360 = pi1308 & n49359;
  assign n49361 = ~pi1308 & ~n49359;
  assign n49362 = ~n49360 & ~n49361;
  assign n49363 = ~n49356 & n49362;
  assign n49364 = n49350 & n49363;
  assign n49365 = ~n49337 & n49364;
  assign n49366 = n49356 & n49362;
  assign n49367 = n49343 & ~n49349;
  assign n49368 = n49366 & n49367;
  assign n49369 = ~n49337 & n49356;
  assign n49370 = n49349 & n49369;
  assign n49371 = ~n49343 & n49370;
  assign n49372 = n49343 & n49349;
  assign n49373 = ~n49337 & n49372;
  assign n49374 = n49362 & n49373;
  assign n49375 = ~n49356 & n49374;
  assign n49376 = ~n49371 & ~n49375;
  assign n49377 = ~n49368 & n49376;
  assign n49378 = ~n49365 & n49377;
  assign n49379 = n49337 & n49356;
  assign n49380 = n49367 & n49379;
  assign n49381 = n49378 & ~n49380;
  assign n49382 = n49331 & ~n49381;
  assign n49383 = ~n49337 & n49343;
  assign n49384 = ~n49349 & n49383;
  assign n49385 = ~n49356 & n49384;
  assign n49386 = ~n49370 & ~n49385;
  assign n49387 = n49337 & n49350;
  assign n49388 = ~n49356 & n49387;
  assign n49389 = n49386 & ~n49388;
  assign n49390 = ~n49362 & ~n49389;
  assign n49391 = n49337 & n49349;
  assign n49392 = n49343 & n49391;
  assign n49393 = ~n49362 & n49392;
  assign n49394 = ~n49356 & n49393;
  assign n49395 = ~n49343 & n49369;
  assign n49396 = ~n49343 & n49349;
  assign n49397 = n49356 & n49396;
  assign n49398 = ~n49395 & ~n49397;
  assign n49399 = ~n49362 & ~n49398;
  assign n49400 = ~n49394 & ~n49399;
  assign n49401 = n49331 & ~n49400;
  assign n49402 = ~n49390 & ~n49401;
  assign n49403 = ~n49382 & n49402;
  assign n49404 = n49337 & ~n49356;
  assign n49405 = n49362 & n49404;
  assign n49406 = n49396 & n49405;
  assign n49407 = n49337 & n49366;
  assign n49408 = n49343 & n49407;
  assign n49409 = ~n49362 & n49383;
  assign n49410 = ~n49343 & ~n49356;
  assign n49411 = n49337 & n49410;
  assign n49412 = ~n49387 & ~n49411;
  assign n49413 = ~n49409 & n49412;
  assign n49414 = n49356 & n49392;
  assign n49415 = n49413 & ~n49414;
  assign n49416 = n49337 & ~n49349;
  assign n49417 = ~n49356 & n49396;
  assign n49418 = ~n49416 & ~n49417;
  assign n49419 = n49362 & ~n49418;
  assign n49420 = n49350 & n49362;
  assign n49421 = n49356 & n49420;
  assign n49422 = ~n49419 & ~n49421;
  assign n49423 = n49415 & n49422;
  assign n49424 = ~n49331 & ~n49423;
  assign n49425 = ~n49408 & ~n49424;
  assign n49426 = ~n49406 & n49425;
  assign n49427 = n49403 & n49426;
  assign n49428 = pi1312 & n49427;
  assign n49429 = ~pi1312 & ~n49427;
  assign po1400 = n49428 | n49429;
  assign n49431 = pi4204 & pi9040;
  assign n49432 = pi4296 & ~pi9040;
  assign n49433 = ~n49431 & ~n49432;
  assign n49434 = pi1275 & n49433;
  assign n49435 = ~pi1275 & ~n49433;
  assign n49436 = ~n49434 & ~n49435;
  assign n49437 = pi4280 & ~pi9040;
  assign n49438 = pi4247 & pi9040;
  assign n49439 = ~n49437 & ~n49438;
  assign n49440 = ~pi1287 & n49439;
  assign n49441 = pi1287 & ~n49439;
  assign n49442 = ~n49440 & ~n49441;
  assign n49443 = pi4208 & ~pi9040;
  assign n49444 = pi4380 & pi9040;
  assign n49445 = ~n49443 & ~n49444;
  assign n49446 = ~pi1298 & n49445;
  assign n49447 = pi1298 & ~n49445;
  assign n49448 = ~n49446 & ~n49447;
  assign n49449 = pi4254 & pi9040;
  assign n49450 = pi4495 & ~pi9040;
  assign n49451 = ~n49449 & ~n49450;
  assign n49452 = ~pi1290 & ~n49451;
  assign n49453 = pi1290 & n49451;
  assign n49454 = ~n49452 & ~n49453;
  assign n49455 = ~n49448 & n49454;
  assign n49456 = n49442 & n49455;
  assign n49457 = pi4281 & ~pi9040;
  assign n49458 = pi4294 & pi9040;
  assign n49459 = ~n49457 & ~n49458;
  assign n49460 = pi1305 & n49459;
  assign n49461 = ~pi1305 & ~n49459;
  assign n49462 = ~n49460 & ~n49461;
  assign n49463 = n49456 & ~n49462;
  assign n49464 = n49448 & ~n49454;
  assign n49465 = n49442 & n49464;
  assign n49466 = ~n49462 & n49465;
  assign n49467 = ~n49463 & ~n49466;
  assign n49468 = ~n49442 & n49464;
  assign n49469 = n49462 & n49468;
  assign n49470 = ~n49448 & ~n49454;
  assign n49471 = n49442 & n49470;
  assign n49472 = n49462 & n49471;
  assign n49473 = ~n49469 & ~n49472;
  assign n49474 = n49467 & n49473;
  assign n49475 = n49436 & ~n49474;
  assign n49476 = n49448 & n49454;
  assign n49477 = n49442 & n49476;
  assign n49478 = n49462 & n49477;
  assign n49479 = ~n49471 & ~n49478;
  assign n49480 = n49436 & ~n49479;
  assign n49481 = n49454 & ~n49462;
  assign n49482 = ~n49436 & n49481;
  assign n49483 = ~n49442 & ~n49448;
  assign n49484 = n49462 & n49464;
  assign n49485 = ~n49483 & ~n49484;
  assign n49486 = ~n49436 & ~n49485;
  assign n49487 = ~n49482 & ~n49486;
  assign n49488 = ~n49442 & n49476;
  assign n49489 = ~n49462 & n49488;
  assign n49490 = n49487 & ~n49489;
  assign n49491 = ~n49442 & n49454;
  assign n49492 = n49462 & n49491;
  assign n49493 = ~n49448 & n49492;
  assign n49494 = n49490 & ~n49493;
  assign n49495 = ~n49480 & n49494;
  assign n49496 = pi4204 & ~pi9040;
  assign n49497 = pi4281 & pi9040;
  assign n49498 = ~n49496 & ~n49497;
  assign n49499 = ~pi1299 & ~n49498;
  assign n49500 = pi1299 & n49498;
  assign n49501 = ~n49499 & ~n49500;
  assign n49502 = ~n49495 & ~n49501;
  assign n49503 = n49442 & n49454;
  assign n49504 = ~n49436 & n49462;
  assign n49505 = n49501 & n49504;
  assign n49506 = n49503 & n49505;
  assign n49507 = n49442 & ~n49462;
  assign n49508 = ~n49454 & n49507;
  assign n49509 = ~n49436 & ~n49508;
  assign n49510 = ~n49442 & n49462;
  assign n49511 = n49448 & n49510;
  assign n49512 = ~n49455 & ~n49503;
  assign n49513 = ~n49462 & ~n49512;
  assign n49514 = n49436 & ~n49468;
  assign n49515 = ~n49513 & n49514;
  assign n49516 = ~n49511 & n49515;
  assign n49517 = ~n49509 & ~n49516;
  assign n49518 = ~n49442 & n49470;
  assign n49519 = n49462 & n49518;
  assign n49520 = ~n49517 & ~n49519;
  assign n49521 = n49501 & ~n49520;
  assign n49522 = ~n49506 & ~n49521;
  assign n49523 = ~n49502 & n49522;
  assign n49524 = ~n49475 & n49523;
  assign n49525 = ~n49436 & ~n49462;
  assign n49526 = n49476 & n49525;
  assign n49527 = ~n49442 & n49526;
  assign n49528 = n49524 & ~n49527;
  assign n49529 = pi1314 & ~n49528;
  assign n49530 = ~pi1314 & ~n49527;
  assign n49531 = n49524 & n49530;
  assign po1402 = n49529 | n49531;
  assign n49533 = ~n49140 & n49159;
  assign n49534 = ~n49184 & ~n49199;
  assign n49535 = n49533 & ~n49534;
  assign n49536 = ~n49140 & ~n49165;
  assign n49537 = n49184 & n49536;
  assign n49538 = ~n49535 & ~n49537;
  assign n49539 = n49177 & ~n49538;
  assign n49540 = ~n49159 & n49165;
  assign n49541 = n49152 & n49540;
  assign n49542 = n49146 & n49541;
  assign n49543 = ~n49216 & ~n49540;
  assign n49544 = n49140 & ~n49543;
  assign n49545 = ~n49159 & ~n49165;
  assign n49546 = ~n49152 & n49545;
  assign n49547 = n49146 & n49546;
  assign n49548 = ~n49544 & ~n49547;
  assign n49549 = ~n49542 & n49548;
  assign n49550 = n49177 & ~n49549;
  assign n49551 = ~n49539 & ~n49550;
  assign n49552 = n49152 & n49166;
  assign n49553 = ~n49146 & n49552;
  assign n49554 = ~n49159 & n49191;
  assign n49555 = ~n49553 & ~n49554;
  assign n49556 = ~n49140 & ~n49555;
  assign n49557 = ~n49153 & ~n49216;
  assign n49558 = n49159 & ~n49557;
  assign n49559 = ~n49191 & ~n49558;
  assign n49560 = ~n49140 & ~n49559;
  assign n49561 = ~n49140 & ~n49159;
  assign n49562 = n49152 & n49561;
  assign n49563 = ~n49165 & n49562;
  assign n49564 = ~n49152 & n49165;
  assign n49565 = ~n49191 & ~n49564;
  assign n49566 = ~n49159 & ~n49565;
  assign n49567 = n49140 & n49159;
  assign n49568 = n49181 & n49567;
  assign n49569 = ~n49165 & n49568;
  assign n49570 = ~n49566 & ~n49569;
  assign n49571 = ~n49563 & n49570;
  assign n49572 = ~n49560 & n49571;
  assign n49573 = ~n49553 & n49572;
  assign n49574 = ~n49177 & ~n49573;
  assign n49575 = n49159 & n49207;
  assign n49576 = ~n49159 & n49216;
  assign n49577 = ~n49575 & ~n49576;
  assign n49578 = n49140 & ~n49577;
  assign n49579 = ~n49574 & ~n49578;
  assign n49580 = ~n49556 & n49579;
  assign n49581 = n49551 & n49580;
  assign n49582 = pi1322 & n49581;
  assign n49583 = ~pi1322 & ~n49581;
  assign po1403 = n49582 | n49583;
  assign n49585 = n49159 & n49190;
  assign n49586 = ~n49546 & ~n49585;
  assign n49587 = n49140 & ~n49586;
  assign n49588 = ~n49152 & n49168;
  assign n49589 = ~n49199 & ~n49588;
  assign n49590 = ~n49140 & ~n49589;
  assign n49591 = ~n49159 & n49185;
  assign n49592 = ~n49563 & ~n49591;
  assign n49593 = ~n49590 & n49592;
  assign n49594 = ~n49587 & n49593;
  assign n49595 = ~n49167 & n49594;
  assign n49596 = ~n49542 & ~n49553;
  assign n49597 = n49595 & n49596;
  assign n49598 = n49177 & ~n49597;
  assign n49599 = n49153 & n49540;
  assign n49600 = n49208 & ~n49599;
  assign n49601 = n49140 & ~n49600;
  assign n49602 = ~n49159 & n49196;
  assign n49603 = ~n49601 & ~n49602;
  assign n49604 = n49146 & n49168;
  assign n49605 = n49159 & n49181;
  assign n49606 = ~n49604 & ~n49605;
  assign n49607 = n49140 & ~n49606;
  assign n49608 = n49140 & n49190;
  assign n49609 = ~n49159 & n49608;
  assign n49610 = ~n49607 & ~n49609;
  assign n49611 = n49603 & n49610;
  assign n49612 = ~n49177 & ~n49611;
  assign n49613 = ~n49185 & ~n49192;
  assign n49614 = ~n49547 & n49613;
  assign n49615 = n49213 & ~n49614;
  assign n49616 = ~n49612 & ~n49615;
  assign n49617 = ~n49167 & ~n49542;
  assign n49618 = ~n49140 & ~n49617;
  assign n49619 = n49616 & ~n49618;
  assign n49620 = ~n49598 & n49619;
  assign n49621 = ~pi1340 & n49620;
  assign n49622 = pi1340 & ~n49620;
  assign po1405 = n49621 | n49622;
  assign n49624 = ~n49290 & ~n49296;
  assign n49625 = n49231 & ~n49624;
  assign n49626 = n49244 & n49280;
  assign n49627 = ~n49625 & ~n49626;
  assign n49628 = n49244 & ~n49256;
  assign n49629 = ~n49304 & ~n49628;
  assign n49630 = ~n49276 & n49629;
  assign n49631 = ~n49231 & ~n49630;
  assign n49632 = n49627 & ~n49631;
  assign n49633 = ~n49237 & ~n49632;
  assign n49634 = ~n49231 & n49309;
  assign n49635 = ~n49244 & n49305;
  assign n49636 = n49231 & n49635;
  assign n49637 = n49250 & n49265;
  assign n49638 = ~n49244 & n49637;
  assign n49639 = n49231 & n49638;
  assign n49640 = ~n49636 & ~n49639;
  assign n49641 = ~n49634 & n49640;
  assign n49642 = ~n49250 & n49295;
  assign n49643 = ~n49231 & n49642;
  assign n49644 = ~n49244 & n49250;
  assign n49645 = ~n49264 & n49644;
  assign n49646 = ~n49309 & ~n49645;
  assign n49647 = ~n49244 & ~n49256;
  assign n49648 = n49250 & n49647;
  assign n49649 = ~n49231 & n49648;
  assign n49650 = n49244 & n49296;
  assign n49651 = n49231 & n49304;
  assign n49652 = ~n49650 & ~n49651;
  assign n49653 = ~n49303 & n49652;
  assign n49654 = ~n49649 & n49653;
  assign n49655 = n49646 & n49654;
  assign n49656 = ~n49643 & n49655;
  assign n49657 = n49237 & ~n49656;
  assign n49658 = n49641 & ~n49657;
  assign n49659 = ~n49633 & n49658;
  assign n49660 = ~pi1329 & ~n49659;
  assign n49661 = pi1329 & n49641;
  assign n49662 = ~n49633 & n49661;
  assign n49663 = ~n49657 & n49662;
  assign po1406 = n49660 | n49663;
  assign n49665 = pi4282 & pi9040;
  assign n49666 = pi4221 & ~pi9040;
  assign n49667 = ~n49665 & ~n49666;
  assign n49668 = ~pi1290 & ~n49667;
  assign n49669 = pi1290 & n49667;
  assign n49670 = ~n49668 & ~n49669;
  assign n49671 = pi4495 & pi9040;
  assign n49672 = pi4380 & ~pi9040;
  assign n49673 = ~n49671 & ~n49672;
  assign n49674 = pi1287 & n49673;
  assign n49675 = ~pi1287 & ~n49673;
  assign n49676 = ~n49674 & ~n49675;
  assign n49677 = pi4288 & pi9040;
  assign n49678 = pi4497 & ~pi9040;
  assign n49679 = ~n49677 & ~n49678;
  assign n49680 = ~pi1300 & n49679;
  assign n49681 = pi1300 & ~n49679;
  assign n49682 = ~n49680 & ~n49681;
  assign n49683 = n49676 & n49682;
  assign n49684 = pi4208 & pi9040;
  assign n49685 = pi4254 & ~pi9040;
  assign n49686 = ~n49684 & ~n49685;
  assign n49687 = ~pi1281 & n49686;
  assign n49688 = pi1281 & ~n49686;
  assign n49689 = ~n49687 & ~n49688;
  assign n49690 = pi4382 & pi9040;
  assign n49691 = pi4220 & ~pi9040;
  assign n49692 = ~n49690 & ~n49691;
  assign n49693 = pi1293 & n49692;
  assign n49694 = ~pi1293 & ~n49692;
  assign n49695 = ~n49693 & ~n49694;
  assign n49696 = n49689 & ~n49695;
  assign n49697 = n49683 & n49696;
  assign n49698 = ~n49676 & ~n49682;
  assign n49699 = pi4280 & pi9040;
  assign n49700 = pi4382 & ~pi9040;
  assign n49701 = ~n49699 & ~n49700;
  assign n49702 = pi1280 & n49701;
  assign n49703 = ~pi1280 & ~n49701;
  assign n49704 = ~n49702 & ~n49703;
  assign n49705 = n49698 & n49704;
  assign n49706 = ~n49676 & n49682;
  assign n49707 = ~n49704 & n49706;
  assign n49708 = ~n49689 & n49707;
  assign n49709 = ~n49705 & ~n49708;
  assign n49710 = n49676 & ~n49682;
  assign n49711 = ~n49689 & n49710;
  assign n49712 = n49709 & ~n49711;
  assign n49713 = ~n49695 & ~n49712;
  assign n49714 = ~n49682 & ~n49704;
  assign n49715 = n49689 & n49695;
  assign n49716 = n49714 & n49715;
  assign n49717 = n49698 & ~n49704;
  assign n49718 = n49689 & n49717;
  assign n49719 = ~n49716 & ~n49718;
  assign n49720 = ~n49713 & n49719;
  assign n49721 = ~n49697 & n49720;
  assign n49722 = n49683 & n49704;
  assign n49723 = n49689 & n49722;
  assign n49724 = ~n49689 & n49704;
  assign n49725 = n49676 & n49724;
  assign n49726 = ~n49682 & n49725;
  assign n49727 = ~n49723 & ~n49726;
  assign n49728 = n49721 & n49727;
  assign n49729 = ~n49670 & ~n49728;
  assign n49730 = n49689 & ~n49704;
  assign n49731 = n49676 & n49730;
  assign n49732 = ~n49682 & n49731;
  assign n49733 = ~n49722 & ~n49732;
  assign n49734 = ~n49695 & ~n49733;
  assign n49735 = n49683 & ~n49704;
  assign n49736 = ~n49689 & n49735;
  assign n49737 = ~n49676 & n49730;
  assign n49738 = n49682 & n49737;
  assign n49739 = ~n49736 & ~n49738;
  assign n49740 = ~n49689 & ~n49704;
  assign n49741 = ~n49682 & n49740;
  assign n49742 = n49689 & n49704;
  assign n49743 = n49676 & n49742;
  assign n49744 = ~n49682 & n49743;
  assign n49745 = ~n49741 & ~n49744;
  assign n49746 = n49695 & ~n49745;
  assign n49747 = n49739 & ~n49746;
  assign n49748 = ~n49734 & n49747;
  assign n49749 = n49670 & ~n49748;
  assign n49750 = n49704 & n49706;
  assign n49751 = ~n49689 & n49750;
  assign n49752 = ~n49717 & ~n49751;
  assign n49753 = ~n49736 & n49752;
  assign n49754 = n49695 & ~n49753;
  assign n49755 = n49682 & n49704;
  assign n49756 = n49689 & n49755;
  assign n49757 = ~n49682 & n49704;
  assign n49758 = ~n49689 & n49757;
  assign n49759 = ~n49756 & ~n49758;
  assign n49760 = ~n49695 & ~n49759;
  assign n49761 = ~n49754 & ~n49760;
  assign n49762 = ~n49676 & ~n49704;
  assign n49763 = n49695 & n49762;
  assign n49764 = n49689 & n49763;
  assign n49765 = n49761 & ~n49764;
  assign n49766 = ~n49749 & n49765;
  assign n49767 = ~n49729 & n49766;
  assign n49768 = ~pi1313 & ~n49767;
  assign n49769 = pi1313 & n49767;
  assign po1408 = n49768 | n49769;
  assign n49771 = n49244 & n49257;
  assign n49772 = ~n49280 & ~n49771;
  assign n49773 = ~n49317 & n49772;
  assign n49774 = ~n49231 & ~n49773;
  assign n49775 = ~n49244 & n49296;
  assign n49776 = ~n49250 & n49256;
  assign n49777 = ~n49265 & ~n49776;
  assign n49778 = n49244 & ~n49777;
  assign n49779 = ~n49775 & ~n49778;
  assign n49780 = ~n49635 & n49779;
  assign n49781 = n49231 & ~n49780;
  assign n49782 = ~n49774 & ~n49781;
  assign n49783 = n49237 & ~n49782;
  assign n49784 = n49256 & n49314;
  assign n49785 = ~n49648 & ~n49771;
  assign n49786 = n49231 & ~n49785;
  assign n49787 = ~n49302 & ~n49786;
  assign n49788 = ~n49306 & ~n49638;
  assign n49789 = ~n49231 & n49304;
  assign n49790 = n49244 & n49789;
  assign n49791 = ~n49643 & ~n49790;
  assign n49792 = n49788 & n49791;
  assign n49793 = n49787 & n49792;
  assign n49794 = ~n49784 & n49793;
  assign n49795 = ~n49237 & ~n49794;
  assign n49796 = n49231 & n49290;
  assign n49797 = ~n49244 & n49796;
  assign n49798 = ~n49639 & ~n49797;
  assign n49799 = ~n49634 & n49798;
  assign n49800 = ~n49244 & n49276;
  assign n49801 = n49244 & n49268;
  assign n49802 = ~n49800 & ~n49801;
  assign n49803 = ~n49231 & ~n49802;
  assign n49804 = n49799 & ~n49803;
  assign n49805 = ~n49795 & n49804;
  assign n49806 = ~n49783 & n49805;
  assign n49807 = ~pi1327 & n49806;
  assign n49808 = pi1327 & ~n49806;
  assign po1409 = n49807 | n49808;
  assign n49810 = ~n49689 & n49717;
  assign n49811 = ~n49738 & ~n49757;
  assign n49812 = n49695 & ~n49811;
  assign n49813 = ~n49810 & ~n49812;
  assign n49814 = ~n49732 & n49813;
  assign n49815 = ~n49689 & ~n49695;
  assign n49816 = n49735 & n49815;
  assign n49817 = ~n49723 & ~n49816;
  assign n49818 = ~n49751 & n49817;
  assign n49819 = n49814 & n49818;
  assign n49820 = n49670 & ~n49819;
  assign n49821 = ~n49704 & n49710;
  assign n49822 = ~n49689 & n49821;
  assign n49823 = ~n49708 & ~n49822;
  assign n49824 = n49695 & n49735;
  assign n49825 = ~n49689 & n49722;
  assign n49826 = ~n49824 & ~n49825;
  assign n49827 = n49689 & n49750;
  assign n49828 = ~n49718 & ~n49827;
  assign n49829 = n49676 & n49704;
  assign n49830 = ~n49682 & ~n49689;
  assign n49831 = ~n49829 & ~n49830;
  assign n49832 = ~n49762 & n49831;
  assign n49833 = ~n49695 & ~n49832;
  assign n49834 = n49828 & ~n49833;
  assign n49835 = n49826 & n49834;
  assign n49836 = n49823 & n49835;
  assign n49837 = ~n49670 & ~n49836;
  assign n49838 = ~n49820 & ~n49837;
  assign n49839 = pi1315 & ~n49838;
  assign n49840 = ~pi1315 & ~n49820;
  assign n49841 = ~n49837 & n49840;
  assign po1410 = n49839 | n49841;
  assign n49843 = ~n49337 & ~n49343;
  assign n49844 = ~n49380 & ~n49843;
  assign n49845 = ~n49410 & n49844;
  assign n49846 = n49362 & ~n49845;
  assign n49847 = ~n49356 & ~n49362;
  assign n49848 = n49343 & n49847;
  assign n49849 = n49337 & ~n49343;
  assign n49850 = n49356 & ~n49362;
  assign n49851 = n49849 & n49850;
  assign n49852 = ~n49337 & ~n49356;
  assign n49853 = ~n49349 & n49852;
  assign n49854 = n49356 & n49373;
  assign n49855 = ~n49853 & ~n49854;
  assign n49856 = ~n49851 & n49855;
  assign n49857 = ~n49848 & n49856;
  assign n49858 = ~n49846 & n49857;
  assign n49859 = ~n49331 & ~n49858;
  assign n49860 = ~n49337 & n49350;
  assign n49861 = n49356 & n49860;
  assign n49862 = ~n49337 & n49396;
  assign n49863 = ~n49356 & n49862;
  assign n49864 = ~n49861 & ~n49863;
  assign n49865 = n49362 & ~n49864;
  assign n49866 = ~n49859 & ~n49865;
  assign n49867 = ~n49356 & n49373;
  assign n49868 = ~n49384 & ~n49392;
  assign n49869 = n49362 & ~n49868;
  assign n49870 = ~n49867 & ~n49869;
  assign n49871 = ~n49388 & n49870;
  assign n49872 = n49331 & ~n49871;
  assign n49873 = ~n49367 & ~n49396;
  assign n49874 = n49337 & ~n49873;
  assign n49875 = ~n49397 & ~n49874;
  assign n49876 = ~n49362 & ~n49875;
  assign n49877 = n49331 & n49876;
  assign n49878 = ~n49872 & ~n49877;
  assign n49879 = n49866 & n49878;
  assign n49880 = pi1321 & ~n49879;
  assign n49881 = ~pi1321 & n49866;
  assign n49882 = n49878 & n49881;
  assign po1411 = n49880 | n49882;
  assign n49884 = ~n49006 & ~n49014;
  assign n49885 = n48956 & ~n49884;
  assign n49886 = ~n49019 & ~n49059;
  assign n49887 = ~n48982 & n49886;
  assign n49888 = ~n48989 & ~n49887;
  assign n49889 = n48956 & n49888;
  assign n49890 = ~n49885 & ~n49889;
  assign n49891 = n49005 & n49062;
  assign n49892 = ~n49064 & ~n49891;
  assign n49893 = ~n49022 & ~n49090;
  assign n49894 = n48989 & ~n49893;
  assign n49895 = n48956 & n49894;
  assign n49896 = n49892 & ~n49895;
  assign n49897 = n48980 & n49018;
  assign n49898 = n48974 & n49897;
  assign n49899 = n48962 & n48997;
  assign n49900 = ~n49055 & ~n49899;
  assign n49901 = n48989 & ~n49900;
  assign n49902 = ~n49020 & ~n49067;
  assign n49903 = n48962 & n49004;
  assign n49904 = ~n49044 & ~n49903;
  assign n49905 = ~n48989 & ~n49904;
  assign n49906 = n49902 & ~n49905;
  assign n49907 = ~n49901 & n49906;
  assign n49908 = ~n49898 & n49907;
  assign n49909 = ~n48956 & ~n49908;
  assign n49910 = ~n49087 & n49104;
  assign n49911 = n48989 & ~n49910;
  assign n49912 = ~n49909 & ~n49911;
  assign n49913 = n49896 & n49912;
  assign n49914 = n49890 & n49913;
  assign n49915 = ~pi1337 & ~n49914;
  assign n49916 = pi1337 & n49896;
  assign n49917 = n49890 & n49916;
  assign n49918 = n49912 & n49917;
  assign po1412 = n49915 | n49918;
  assign n49920 = n49268 & n49314;
  assign n49921 = ~n49800 & ~n49920;
  assign n49922 = ~n49244 & n49256;
  assign n49923 = ~n49645 & ~n49922;
  assign n49924 = n49231 & ~n49923;
  assign n49925 = n49264 & n49266;
  assign n49926 = ~n49924 & ~n49925;
  assign n49927 = n49921 & n49926;
  assign n49928 = n49237 & ~n49927;
  assign n49929 = ~n49306 & ~n49637;
  assign n49930 = ~n49244 & n49295;
  assign n49931 = n49929 & ~n49930;
  assign n49932 = ~n49231 & ~n49931;
  assign n49933 = n49268 & n49301;
  assign n49934 = ~n49317 & ~n49933;
  assign n49935 = ~n49932 & n49934;
  assign n49936 = ~n49276 & ~n49286;
  assign n49937 = n49231 & ~n49936;
  assign n49938 = n49935 & ~n49937;
  assign n49939 = ~n49237 & ~n49938;
  assign n49940 = ~n49928 & ~n49939;
  assign n49941 = ~n49244 & n49275;
  assign n49942 = n49244 & ~n49281;
  assign n49943 = ~n49941 & ~n49942;
  assign n49944 = n49231 & ~n49943;
  assign n49945 = ~n49231 & n49244;
  assign n49946 = n49624 & ~n49637;
  assign n49947 = n49945 & ~n49946;
  assign n49948 = ~n49944 & ~n49947;
  assign n49949 = n49940 & n49948;
  assign n49950 = ~pi1323 & ~n49949;
  assign n49951 = pi1323 & n49948;
  assign n49952 = ~n49939 & n49951;
  assign n49953 = ~n49928 & n49952;
  assign po1415 = n49950 | n49953;
  assign n49955 = ~n49356 & n49874;
  assign n49956 = n49349 & n49852;
  assign n49957 = ~n49416 & ~n49956;
  assign n49958 = ~n49862 & n49957;
  assign n49959 = n49362 & ~n49958;
  assign n49960 = ~n49391 & ~n49860;
  assign n49961 = ~n49362 & ~n49960;
  assign n49962 = ~n49959 & ~n49961;
  assign n49963 = ~n49955 & n49962;
  assign n49964 = n49356 & n49384;
  assign n49965 = n49963 & ~n49964;
  assign n49966 = n49331 & ~n49965;
  assign n49967 = n49366 & ~n49960;
  assign n49968 = ~n49387 & ~n49392;
  assign n49969 = ~n49384 & ~n49862;
  assign n49970 = n49968 & n49969;
  assign n49971 = ~n49356 & ~n49970;
  assign n49972 = ~n49967 & ~n49971;
  assign n49973 = ~n49854 & n49972;
  assign n49974 = ~n49331 & ~n49973;
  assign n49975 = ~n49966 & ~n49974;
  assign n49976 = ~n49356 & n49860;
  assign n49977 = ~n49964 & ~n49976;
  assign n49978 = ~n49362 & ~n49977;
  assign n49979 = n49975 & ~n49978;
  assign n49980 = pi1333 & ~n49979;
  assign n49981 = ~pi1333 & ~n49978;
  assign n49982 = ~n49974 & n49981;
  assign n49983 = ~n49966 & n49982;
  assign po1416 = n49980 | n49983;
  assign n49985 = ~n49140 & n49196;
  assign n49986 = ~n49159 & n49181;
  assign n49987 = ~n49180 & ~n49986;
  assign n49988 = ~n49140 & ~n49987;
  assign n49989 = n49140 & ~n49565;
  assign n49990 = ~n49988 & ~n49989;
  assign n49991 = ~n49575 & n49990;
  assign n49992 = n49177 & ~n49991;
  assign n49993 = ~n49985 & ~n49992;
  assign n49994 = n49165 & n49533;
  assign n49995 = ~n49545 & ~n49994;
  assign n49996 = ~n49146 & ~n49995;
  assign n49997 = ~n49167 & ~n49996;
  assign n49998 = ~n49546 & n49997;
  assign n49999 = n49159 & n49199;
  assign n50000 = n49140 & n49182;
  assign n50001 = ~n49999 & ~n50000;
  assign n50002 = n49998 & n50001;
  assign n50003 = ~n49177 & ~n50002;
  assign n50004 = ~n49591 & ~n49605;
  assign n50005 = n49140 & ~n50004;
  assign n50006 = ~n50003 & ~n50005;
  assign n50007 = n49993 & n50006;
  assign n50008 = ~pi1348 & ~n50007;
  assign n50009 = ~n49992 & n50006;
  assign n50010 = pi1348 & n50009;
  assign n50011 = ~n49985 & n50010;
  assign po1417 = n50008 | n50011;
  assign n50013 = pi4287 & pi9040;
  assign n50014 = pi4228 & ~pi9040;
  assign n50015 = ~n50013 & ~n50014;
  assign n50016 = pi1309 & n50015;
  assign n50017 = ~pi1309 & ~n50015;
  assign n50018 = ~n50016 & ~n50017;
  assign n50019 = pi4309 & pi9040;
  assign n50020 = pi4302 & ~pi9040;
  assign n50021 = ~n50019 & ~n50020;
  assign n50022 = pi1291 & n50021;
  assign n50023 = ~pi1291 & ~n50021;
  assign n50024 = ~n50022 & ~n50023;
  assign n50025 = pi4205 & pi9040;
  assign n50026 = pi4404 & ~pi9040;
  assign n50027 = ~n50025 & ~n50026;
  assign n50028 = ~pi1307 & n50027;
  assign n50029 = pi1307 & ~n50027;
  assign n50030 = ~n50028 & ~n50029;
  assign n50031 = n50024 & ~n50030;
  assign n50032 = n50018 & n50031;
  assign n50033 = pi1307 & n50027;
  assign n50034 = ~pi1307 & ~n50027;
  assign n50035 = ~n50033 & ~n50034;
  assign n50036 = n50024 & ~n50035;
  assign n50037 = ~n50018 & n50036;
  assign n50038 = ~n50032 & ~n50037;
  assign n50039 = pi4213 & pi9040;
  assign n50040 = pi4287 & ~pi9040;
  assign n50041 = ~n50039 & ~n50040;
  assign n50042 = pi1297 & n50041;
  assign n50043 = ~pi1297 & ~n50041;
  assign n50044 = ~n50042 & ~n50043;
  assign n50045 = n50018 & ~n50044;
  assign n50046 = n50035 & n50045;
  assign n50047 = n50038 & ~n50046;
  assign n50048 = pi4206 & pi9040;
  assign n50049 = pi4310 & ~pi9040;
  assign n50050 = ~n50048 & ~n50049;
  assign n50051 = ~pi1277 & n50050;
  assign n50052 = pi1277 & ~n50050;
  assign n50053 = ~n50051 & ~n50052;
  assign n50054 = ~pi4698 & ~pi9040;
  assign n50055 = ~pi4228 & pi9040;
  assign n50056 = ~n50054 & ~n50055;
  assign n50057 = ~pi1271 & n50056;
  assign n50058 = pi1271 & ~n50056;
  assign n50059 = ~n50057 & ~n50058;
  assign n50060 = n50053 & n50059;
  assign n50061 = ~n50047 & n50060;
  assign n50062 = ~n50024 & ~n50035;
  assign n50063 = n50018 & n50062;
  assign n50064 = n50044 & n50059;
  assign n50065 = n50063 & n50064;
  assign n50066 = n50018 & n50036;
  assign n50067 = ~n50053 & n50066;
  assign n50068 = ~n50024 & ~n50030;
  assign n50069 = n50044 & n50068;
  assign n50070 = ~n50018 & n50035;
  assign n50071 = ~n50069 & ~n50070;
  assign n50072 = ~n50053 & ~n50071;
  assign n50073 = ~n50067 & ~n50072;
  assign n50074 = n50059 & ~n50073;
  assign n50075 = ~n50065 & ~n50074;
  assign n50076 = ~n50018 & ~n50044;
  assign n50077 = ~n50035 & n50076;
  assign n50078 = ~n50024 & n50077;
  assign n50079 = ~n50018 & n50044;
  assign n50080 = n50035 & n50079;
  assign n50081 = ~n50078 & ~n50080;
  assign n50082 = ~n50053 & ~n50081;
  assign n50083 = n50075 & ~n50082;
  assign n50084 = n50044 & n50053;
  assign n50085 = n50068 & n50084;
  assign n50086 = n50018 & n50085;
  assign n50087 = ~n50031 & ~n50062;
  assign n50088 = n50045 & ~n50087;
  assign n50089 = n50024 & n50077;
  assign n50090 = ~n50088 & ~n50089;
  assign n50091 = ~n50018 & n50068;
  assign n50092 = ~n50044 & n50053;
  assign n50093 = n50091 & n50092;
  assign n50094 = n50079 & ~n50087;
  assign n50095 = n50044 & n50066;
  assign n50096 = ~n50094 & ~n50095;
  assign n50097 = ~n50093 & n50096;
  assign n50098 = n50090 & n50097;
  assign n50099 = ~n50086 & n50098;
  assign n50100 = ~n50044 & ~n50053;
  assign n50101 = n50018 & n50100;
  assign n50102 = ~n50024 & n50101;
  assign n50103 = n50099 & ~n50102;
  assign n50104 = ~n50059 & ~n50103;
  assign n50105 = n50083 & ~n50104;
  assign n50106 = ~n50061 & n50105;
  assign n50107 = ~pi1330 & ~n50106;
  assign n50108 = pi1330 & n50083;
  assign n50109 = ~n50061 & n50108;
  assign n50110 = ~n50104 & n50109;
  assign po1420 = n50107 | n50110;
  assign n50112 = ~n50018 & n50031;
  assign n50113 = n50018 & n50068;
  assign n50114 = ~n50112 & ~n50113;
  assign n50115 = ~n50053 & ~n50114;
  assign n50116 = ~n50044 & n50062;
  assign n50117 = ~n50032 & ~n50116;
  assign n50118 = ~n50091 & n50117;
  assign n50119 = n50053 & ~n50118;
  assign n50120 = ~n50115 & ~n50119;
  assign n50121 = ~n50067 & ~n50078;
  assign n50122 = n50120 & n50121;
  assign n50123 = ~n50059 & ~n50122;
  assign n50124 = n50044 & n50113;
  assign n50125 = n50044 & n50062;
  assign n50126 = n50036 & ~n50044;
  assign n50127 = ~n50125 & ~n50126;
  assign n50128 = n50053 & ~n50127;
  assign n50129 = ~n50124 & ~n50128;
  assign n50130 = n50018 & ~n50053;
  assign n50131 = ~n50035 & n50130;
  assign n50132 = ~n50024 & n50131;
  assign n50133 = n50038 & ~n50132;
  assign n50134 = ~n50091 & n50133;
  assign n50135 = ~n50044 & ~n50134;
  assign n50136 = n50129 & ~n50135;
  assign n50137 = n50059 & ~n50136;
  assign n50138 = ~n50123 & ~n50137;
  assign n50139 = ~n50018 & n50125;
  assign n50140 = ~n50095 & ~n50139;
  assign n50141 = ~n50053 & ~n50140;
  assign n50142 = ~n50018 & n50024;
  assign n50143 = n50084 & n50142;
  assign n50144 = ~n50141 & ~n50143;
  assign n50145 = n50138 & n50144;
  assign n50146 = ~pi1326 & ~n50145;
  assign n50147 = pi1326 & ~n50141;
  assign n50148 = n50138 & n50147;
  assign n50149 = ~n50143 & n50148;
  assign po1421 = n50146 | n50149;
  assign n50151 = ~n50018 & ~n50068;
  assign n50152 = ~n50053 & n50151;
  assign n50153 = ~n50044 & n50152;
  assign n50154 = n50024 & n50044;
  assign n50155 = n50018 & n50154;
  assign n50156 = ~n50069 & ~n50155;
  assign n50157 = ~n50053 & ~n50156;
  assign n50158 = ~n50153 & ~n50157;
  assign n50159 = n50053 & ~n50076;
  assign n50160 = ~n50087 & n50159;
  assign n50161 = ~n50093 & ~n50160;
  assign n50162 = ~n50089 & n50161;
  assign n50163 = n50158 & n50162;
  assign n50164 = n50059 & ~n50163;
  assign n50165 = n50036 & n50100;
  assign n50166 = ~n50018 & n50165;
  assign n50167 = ~n50053 & n50113;
  assign n50168 = ~n50044 & n50167;
  assign n50169 = ~n50166 & ~n50168;
  assign n50170 = ~n50164 & n50169;
  assign n50171 = n50032 & n50053;
  assign n50172 = n50044 & n50171;
  assign n50173 = n50053 & ~n50059;
  assign n50174 = n50076 & ~n50087;
  assign n50175 = ~n50069 & ~n50174;
  assign n50176 = ~n50066 & n50175;
  assign n50177 = n50173 & ~n50176;
  assign n50178 = n50037 & n50044;
  assign n50179 = ~n50018 & n50154;
  assign n50180 = ~n50125 & ~n50179;
  assign n50181 = ~n50044 & n50068;
  assign n50182 = ~n50063 & ~n50181;
  assign n50183 = n50180 & n50182;
  assign n50184 = ~n50053 & ~n50183;
  assign n50185 = ~n50178 & ~n50184;
  assign n50186 = ~n50059 & ~n50185;
  assign n50187 = ~n50177 & ~n50186;
  assign n50188 = ~n50172 & n50187;
  assign n50189 = n50170 & n50188;
  assign n50190 = pi1332 & ~n50189;
  assign n50191 = ~pi1332 & n50170;
  assign n50192 = n50188 & n50191;
  assign po1422 = n50190 | n50192;
  assign n50194 = ~n50063 & ~n50154;
  assign n50195 = n50060 & ~n50194;
  assign n50196 = ~n50053 & n50079;
  assign n50197 = n50031 & n50196;
  assign n50198 = n50018 & n50084;
  assign n50199 = ~n50035 & n50198;
  assign n50200 = ~n50197 & ~n50199;
  assign n50201 = n50018 & n50044;
  assign n50202 = ~n50031 & n50059;
  assign n50203 = n50201 & n50202;
  assign n50204 = n50200 & ~n50203;
  assign n50205 = ~n50125 & ~n50181;
  assign n50206 = ~n50053 & ~n50205;
  assign n50207 = ~n50166 & ~n50206;
  assign n50208 = n50059 & ~n50207;
  assign n50209 = ~n50031 & ~n50142;
  assign n50210 = ~n50044 & ~n50209;
  assign n50211 = ~n50113 & ~n50210;
  assign n50212 = n50053 & ~n50211;
  assign n50213 = ~n50174 & ~n50212;
  assign n50214 = n50044 & n50091;
  assign n50215 = ~n50035 & n50045;
  assign n50216 = n50044 & ~n50209;
  assign n50217 = ~n50215 & ~n50216;
  assign n50218 = ~n50053 & ~n50217;
  assign n50219 = ~n50214 & ~n50218;
  assign n50220 = n50213 & n50219;
  assign n50221 = ~n50059 & ~n50220;
  assign n50222 = ~n50208 & ~n50221;
  assign n50223 = n50204 & n50222;
  assign n50224 = ~n50195 & n50223;
  assign n50225 = pi1342 & ~n50224;
  assign n50226 = ~pi1342 & n50204;
  assign n50227 = ~n50195 & n50226;
  assign n50228 = n50222 & n50227;
  assign po1423 = n50225 | n50228;
  assign n50230 = pi4284 & pi9040;
  assign n50231 = pi4304 & ~pi9040;
  assign n50232 = ~n50230 & ~n50231;
  assign n50233 = pi1279 & n50232;
  assign n50234 = ~pi1279 & ~n50232;
  assign n50235 = ~n50233 & ~n50234;
  assign n50236 = pi4374 & ~pi9040;
  assign n50237 = pi4384 & pi9040;
  assign n50238 = ~n50236 & ~n50237;
  assign n50239 = ~pi1311 & n50238;
  assign n50240 = pi1311 & ~n50238;
  assign n50241 = ~n50239 & ~n50240;
  assign n50242 = pi4384 & ~pi9040;
  assign n50243 = pi4593 & pi9040;
  assign n50244 = ~n50242 & ~n50243;
  assign n50245 = ~pi1306 & n50244;
  assign n50246 = pi1306 & ~n50244;
  assign n50247 = ~n50245 & ~n50246;
  assign n50248 = pi4221 & pi9040;
  assign n50249 = pi4484 & ~pi9040;
  assign n50250 = ~n50248 & ~n50249;
  assign n50251 = ~pi1310 & n50250;
  assign n50252 = pi1310 & ~n50250;
  assign n50253 = ~n50251 & ~n50252;
  assign n50254 = pi4293 & pi9040;
  assign n50255 = pi4282 & ~pi9040;
  assign n50256 = ~n50254 & ~n50255;
  assign n50257 = pi1289 & n50256;
  assign n50258 = ~pi1289 & ~n50256;
  assign n50259 = ~n50257 & ~n50258;
  assign n50260 = n50253 & ~n50259;
  assign n50261 = ~n50247 & n50260;
  assign n50262 = n50241 & n50261;
  assign n50263 = pi4316 & pi9040;
  assign n50264 = pi4288 & ~pi9040;
  assign n50265 = ~n50263 & ~n50264;
  assign n50266 = pi1301 & n50265;
  assign n50267 = ~pi1301 & ~n50265;
  assign n50268 = ~n50266 & ~n50267;
  assign n50269 = ~pi1289 & n50256;
  assign n50270 = pi1289 & ~n50256;
  assign n50271 = ~n50269 & ~n50270;
  assign n50272 = n50253 & ~n50271;
  assign n50273 = n50247 & n50272;
  assign n50274 = ~n50253 & ~n50271;
  assign n50275 = ~n50247 & n50274;
  assign n50276 = n50241 & n50275;
  assign n50277 = ~n50273 & ~n50276;
  assign n50278 = ~n50247 & ~n50259;
  assign n50279 = ~n50241 & n50278;
  assign n50280 = ~n50253 & ~n50259;
  assign n50281 = n50247 & n50280;
  assign n50282 = n50241 & n50281;
  assign n50283 = ~n50279 & ~n50282;
  assign n50284 = n50277 & n50283;
  assign n50285 = ~n50268 & ~n50284;
  assign n50286 = n50247 & n50260;
  assign n50287 = ~n50241 & n50274;
  assign n50288 = n50241 & ~n50247;
  assign n50289 = n50253 & n50288;
  assign n50290 = ~n50287 & ~n50289;
  assign n50291 = ~n50286 & n50290;
  assign n50292 = n50268 & ~n50291;
  assign n50293 = n50247 & n50274;
  assign n50294 = ~n50241 & n50293;
  assign n50295 = ~n50292 & ~n50294;
  assign n50296 = ~n50285 & n50295;
  assign n50297 = ~n50262 & n50296;
  assign n50298 = ~n50235 & ~n50297;
  assign n50299 = ~n50241 & ~n50268;
  assign n50300 = n50275 & n50299;
  assign n50301 = ~n50268 & n50286;
  assign n50302 = ~n50247 & n50272;
  assign n50303 = ~n50268 & n50302;
  assign n50304 = ~n50301 & ~n50303;
  assign n50305 = n50241 & ~n50304;
  assign n50306 = ~n50300 & ~n50305;
  assign n50307 = ~n50241 & n50272;
  assign n50308 = n50241 & n50274;
  assign n50309 = ~n50307 & ~n50308;
  assign n50310 = ~n50253 & n50278;
  assign n50311 = n50309 & ~n50310;
  assign n50312 = ~n50273 & n50311;
  assign n50313 = n50268 & ~n50312;
  assign n50314 = n50241 & n50293;
  assign n50315 = ~n50313 & ~n50314;
  assign n50316 = n50241 & n50310;
  assign n50317 = ~n50241 & ~n50253;
  assign n50318 = n50247 & n50317;
  assign n50319 = ~n50259 & n50318;
  assign n50320 = ~n50316 & ~n50319;
  assign n50321 = n50315 & n50320;
  assign n50322 = n50306 & n50321;
  assign n50323 = n50235 & ~n50322;
  assign n50324 = ~n50241 & n50261;
  assign n50325 = ~n50241 & n50273;
  assign n50326 = ~n50324 & ~n50325;
  assign n50327 = ~n50268 & ~n50326;
  assign n50328 = ~n50323 & ~n50327;
  assign n50329 = ~n50241 & n50286;
  assign n50330 = ~n50316 & ~n50329;
  assign n50331 = n50268 & ~n50330;
  assign n50332 = n50328 & ~n50331;
  assign n50333 = ~n50298 & n50332;
  assign n50334 = pi1336 & ~n50333;
  assign n50335 = ~pi1336 & n50333;
  assign po1424 = n50334 | n50335;
  assign n50337 = ~n50241 & n50310;
  assign n50338 = ~n50271 & n50288;
  assign n50339 = ~n50289 & ~n50293;
  assign n50340 = ~n50268 & ~n50339;
  assign n50341 = ~n50338 & ~n50340;
  assign n50342 = n50247 & ~n50259;
  assign n50343 = n50241 & n50342;
  assign n50344 = ~n50241 & n50260;
  assign n50345 = ~n50343 & ~n50344;
  assign n50346 = n50247 & n50253;
  assign n50347 = n50345 & ~n50346;
  assign n50348 = ~n50275 & n50347;
  assign n50349 = n50268 & ~n50348;
  assign n50350 = n50341 & ~n50349;
  assign n50351 = ~n50337 & n50350;
  assign n50352 = n50235 & ~n50351;
  assign n50353 = n50241 & n50273;
  assign n50354 = ~n50329 & ~n50337;
  assign n50355 = ~n50353 & n50354;
  assign n50356 = n50268 & ~n50355;
  assign n50357 = ~n50352 & ~n50356;
  assign n50358 = n50247 & ~n50253;
  assign n50359 = ~n50268 & n50358;
  assign n50360 = ~n50241 & n50359;
  assign n50361 = n50241 & n50268;
  assign n50362 = n50278 & n50361;
  assign n50363 = ~n50241 & n50302;
  assign n50364 = ~n50362 & ~n50363;
  assign n50365 = ~n50247 & n50253;
  assign n50366 = ~n50241 & n50365;
  assign n50367 = ~n50281 & ~n50366;
  assign n50368 = ~n50268 & ~n50367;
  assign n50369 = n50253 & ~n50268;
  assign n50370 = n50247 & n50369;
  assign n50371 = n50241 & n50370;
  assign n50372 = ~n50368 & ~n50371;
  assign n50373 = n50364 & n50372;
  assign n50374 = ~n50235 & ~n50373;
  assign n50375 = ~n50360 & ~n50374;
  assign n50376 = ~n50276 & n50375;
  assign n50377 = n50357 & n50376;
  assign n50378 = ~pi1328 & ~n50377;
  assign n50379 = ~n50276 & ~n50352;
  assign n50380 = ~n50356 & n50379;
  assign n50381 = n50375 & n50380;
  assign n50382 = pi1328 & n50381;
  assign po1425 = n50378 | n50382;
  assign n50384 = n49384 & n49847;
  assign n50385 = n49356 & n49387;
  assign n50386 = ~n49854 & ~n50385;
  assign n50387 = ~n49362 & ~n50386;
  assign n50388 = ~n50384 & ~n50387;
  assign n50389 = ~n49408 & n50388;
  assign n50390 = ~n49331 & ~n49362;
  assign n50391 = ~n49356 & n49392;
  assign n50392 = ~n49387 & ~n50391;
  assign n50393 = ~n49862 & n50392;
  assign n50394 = n50390 & ~n50393;
  assign n50395 = n49362 & n49860;
  assign n50396 = ~n49380 & ~n49406;
  assign n50397 = ~n49375 & n50396;
  assign n50398 = ~n50395 & n50397;
  assign n50399 = ~n49331 & ~n50398;
  assign n50400 = ~n50394 & ~n50399;
  assign n50401 = n49356 & n49391;
  assign n50402 = ~n49356 & n49367;
  assign n50403 = ~n49383 & ~n50402;
  assign n50404 = ~n49362 & ~n50403;
  assign n50405 = ~n49356 & n49420;
  assign n50406 = ~n49853 & ~n50405;
  assign n50407 = n49362 & n49862;
  assign n50408 = n50406 & ~n50407;
  assign n50409 = ~n50404 & n50408;
  assign n50410 = ~n50401 & n50409;
  assign n50411 = n49331 & ~n50410;
  assign n50412 = n49356 & n50407;
  assign n50413 = ~n50411 & ~n50412;
  assign n50414 = n50400 & n50413;
  assign n50415 = n50389 & n50414;
  assign n50416 = ~pi1344 & n50415;
  assign n50417 = pi1344 & ~n50415;
  assign po1426 = n50416 | n50417;
  assign n50419 = n49442 & n49448;
  assign n50420 = n49436 & n50419;
  assign n50421 = n49462 & n50420;
  assign n50422 = ~n49436 & n49464;
  assign n50423 = ~n49442 & n50422;
  assign n50424 = ~n49436 & n49455;
  assign n50425 = n49462 & n50424;
  assign n50426 = ~n50423 & ~n50425;
  assign n50427 = n49462 & n49476;
  assign n50428 = ~n50419 & ~n50427;
  assign n50429 = ~n49442 & ~n49462;
  assign n50430 = ~n49448 & n50429;
  assign n50431 = n50428 & ~n50430;
  assign n50432 = n49436 & ~n50431;
  assign n50433 = ~n49472 & ~n50432;
  assign n50434 = n50426 & n50433;
  assign n50435 = ~n49501 & ~n50434;
  assign n50436 = ~n49488 & ~n49508;
  assign n50437 = ~n49518 & n50436;
  assign n50438 = ~n49436 & ~n50437;
  assign n50439 = ~n49448 & n49507;
  assign n50440 = ~n49462 & n49468;
  assign n50441 = n49454 & n49483;
  assign n50442 = ~n50440 & ~n50441;
  assign n50443 = n49436 & ~n50442;
  assign n50444 = ~n50439 & ~n50443;
  assign n50445 = ~n50438 & n50444;
  assign n50446 = ~n49478 & ~n49519;
  assign n50447 = n50445 & n50446;
  assign n50448 = n49501 & ~n50447;
  assign n50449 = ~n49463 & ~n49469;
  assign n50450 = ~n49436 & ~n50449;
  assign n50451 = ~n49527 & ~n50450;
  assign n50452 = ~n50448 & n50451;
  assign n50453 = ~n50435 & n50452;
  assign n50454 = ~n50421 & n50453;
  assign n50455 = pi1354 & n50454;
  assign n50456 = ~pi1354 & ~n50454;
  assign po1427 = n50455 | n50456;
  assign n50458 = n49689 & n49710;
  assign n50459 = ~n49827 & ~n50458;
  assign n50460 = n49695 & n50459;
  assign n50461 = ~n49689 & n49755;
  assign n50462 = ~n49683 & ~n49698;
  assign n50463 = n49704 & ~n50462;
  assign n50464 = n49682 & n49730;
  assign n50465 = ~n49689 & n49698;
  assign n50466 = ~n50464 & ~n50465;
  assign n50467 = ~n49695 & n50466;
  assign n50468 = ~n50463 & n50467;
  assign n50469 = ~n50461 & n50468;
  assign n50470 = ~n50460 & ~n50469;
  assign n50471 = ~n49689 & n50463;
  assign n50472 = ~n49822 & ~n50471;
  assign n50473 = ~n50470 & n50472;
  assign n50474 = n49670 & ~n50473;
  assign n50475 = n49695 & ~n50462;
  assign n50476 = n49689 & n50475;
  assign n50477 = ~n49689 & n49706;
  assign n50478 = ~n49726 & ~n50477;
  assign n50479 = n49695 & ~n50478;
  assign n50480 = ~n49704 & n50475;
  assign n50481 = ~n50479 & ~n50480;
  assign n50482 = ~n50476 & n50481;
  assign n50483 = ~n49670 & ~n50482;
  assign n50484 = ~n50474 & ~n50483;
  assign n50485 = ~n49695 & ~n50459;
  assign n50486 = ~n49708 & ~n50485;
  assign n50487 = ~n49670 & ~n50486;
  assign n50488 = n49695 & n49708;
  assign n50489 = ~n49695 & ~n50472;
  assign n50490 = ~n50488 & ~n50489;
  assign n50491 = ~n50487 & n50490;
  assign n50492 = n50484 & n50491;
  assign n50493 = pi1331 & ~n50492;
  assign n50494 = ~pi1331 & n50491;
  assign n50495 = ~n50483 & n50494;
  assign n50496 = ~n50474 & n50495;
  assign po1428 = n50493 | n50496;
  assign n50498 = n50241 & ~n50268;
  assign n50499 = ~n50253 & n50498;
  assign n50500 = n50241 & n50247;
  assign n50501 = ~n50259 & n50500;
  assign n50502 = n50253 & n50501;
  assign n50503 = ~n50293 & ~n50502;
  assign n50504 = n50268 & ~n50503;
  assign n50505 = n50326 & ~n50504;
  assign n50506 = ~n50499 & n50505;
  assign n50507 = n50235 & ~n50506;
  assign n50508 = ~n50268 & n50319;
  assign n50509 = n50281 & n50361;
  assign n50510 = ~n50289 & ~n50509;
  assign n50511 = ~n50293 & ~n50302;
  assign n50512 = n50241 & n50272;
  assign n50513 = n50511 & ~n50512;
  assign n50514 = ~n50268 & ~n50513;
  assign n50515 = n50268 & n50275;
  assign n50516 = n50354 & ~n50515;
  assign n50517 = ~n50514 & n50516;
  assign n50518 = n50510 & n50517;
  assign n50519 = ~n50235 & ~n50518;
  assign n50520 = ~n50508 & ~n50519;
  assign n50521 = ~n50507 & n50520;
  assign n50522 = n50302 & n50361;
  assign n50523 = n50268 & n50278;
  assign n50524 = ~n50241 & n50523;
  assign n50525 = ~n50522 & ~n50524;
  assign n50526 = n50268 & n50325;
  assign n50527 = n50525 & ~n50526;
  assign n50528 = n50521 & n50527;
  assign n50529 = ~pi1325 & ~n50528;
  assign n50530 = pi1325 & n50527;
  assign n50531 = n50520 & n50530;
  assign n50532 = ~n50507 & n50531;
  assign po1429 = n50529 | n50532;
  assign n50534 = n49442 & ~n49448;
  assign n50535 = ~n49436 & n50534;
  assign n50536 = n49462 & n50535;
  assign n50537 = n49442 & n49462;
  assign n50538 = n49454 & n50537;
  assign n50539 = ~n49448 & n50538;
  assign n50540 = ~n49462 & n49491;
  assign n50541 = ~n49469 & ~n50540;
  assign n50542 = ~n50539 & n50541;
  assign n50543 = ~n50536 & n50542;
  assign n50544 = n49436 & n49465;
  assign n50545 = n50543 & ~n50544;
  assign n50546 = n49501 & ~n50545;
  assign n50547 = ~n49462 & n49471;
  assign n50548 = ~n49519 & ~n50547;
  assign n50549 = n49436 & ~n50548;
  assign n50550 = ~n49436 & ~n49501;
  assign n50551 = n49503 & n50550;
  assign n50552 = n49448 & n50429;
  assign n50553 = ~n49491 & ~n50552;
  assign n50554 = ~n49471 & n50553;
  assign n50555 = n49436 & ~n50554;
  assign n50556 = ~n49462 & n49477;
  assign n50557 = ~n50555 & ~n50556;
  assign n50558 = ~n49501 & ~n50557;
  assign n50559 = ~n50551 & ~n50558;
  assign n50560 = ~n50549 & n50559;
  assign n50561 = n49462 & n49503;
  assign n50562 = ~n49462 & n49518;
  assign n50563 = ~n50561 & ~n50562;
  assign n50564 = ~n49466 & n50563;
  assign n50565 = ~n49469 & n50564;
  assign n50566 = ~n49436 & ~n50565;
  assign n50567 = n50560 & ~n50566;
  assign n50568 = ~n50546 & n50567;
  assign n50569 = ~pi1349 & ~n50568;
  assign n50570 = pi1349 & n50560;
  assign n50571 = ~n50546 & n50570;
  assign n50572 = ~n50566 & n50571;
  assign po1430 = n50569 | n50572;
  assign n50574 = ~n49462 & n50441;
  assign n50575 = ~n49488 & ~n50561;
  assign n50576 = n49436 & ~n50575;
  assign n50577 = ~n50574 & ~n50576;
  assign n50578 = n49454 & n49525;
  assign n50579 = ~n49448 & n50578;
  assign n50580 = ~n49454 & n49504;
  assign n50581 = ~n49448 & n50580;
  assign n50582 = ~n50579 & ~n50581;
  assign n50583 = ~n50423 & n50582;
  assign n50584 = ~n49466 & ~n49478;
  assign n50585 = ~n49454 & n49510;
  assign n50586 = n50584 & ~n50585;
  assign n50587 = n50583 & n50586;
  assign n50588 = n50577 & n50587;
  assign n50589 = ~n49501 & ~n50588;
  assign n50590 = ~n49465 & ~n49488;
  assign n50591 = n49462 & ~n50590;
  assign n50592 = ~n49518 & ~n50439;
  assign n50593 = ~n49492 & n50592;
  assign n50594 = n49436 & ~n50593;
  assign n50595 = ~n49462 & n49476;
  assign n50596 = ~n50539 & ~n50595;
  assign n50597 = ~n49436 & ~n50596;
  assign n50598 = ~n50547 & ~n50597;
  assign n50599 = ~n50594 & n50598;
  assign n50600 = ~n50591 & n50599;
  assign n50601 = n49501 & ~n50600;
  assign n50602 = n49436 & n49508;
  assign n50603 = ~n50601 & ~n50602;
  assign n50604 = ~n49436 & n50574;
  assign n50605 = n50603 & ~n50604;
  assign n50606 = ~n50589 & n50605;
  assign n50607 = ~pi1338 & ~n50606;
  assign n50608 = pi1338 & n50603;
  assign n50609 = ~n50589 & n50608;
  assign n50610 = ~n50604 & n50609;
  assign po1431 = n50607 | n50610;
  assign n50612 = n49695 & n49736;
  assign n50613 = n49730 & ~n50462;
  assign n50614 = ~n49750 & ~n50613;
  assign n50615 = ~n49822 & n50614;
  assign n50616 = ~n49695 & ~n50615;
  assign n50617 = ~n49689 & n49705;
  assign n50618 = ~n50616 & ~n50617;
  assign n50619 = n49689 & n49829;
  assign n50620 = ~n49707 & ~n50619;
  assign n50621 = ~n50465 & n50620;
  assign n50622 = n49695 & ~n50621;
  assign n50623 = n50618 & ~n50622;
  assign n50624 = n49670 & ~n50623;
  assign n50625 = ~n50612 & ~n50624;
  assign n50626 = n49689 & n49698;
  assign n50627 = ~n49821 & ~n50626;
  assign n50628 = n49695 & ~n50627;
  assign n50629 = ~n49751 & ~n50628;
  assign n50630 = ~n49726 & ~n49736;
  assign n50631 = ~n49689 & n49762;
  assign n50632 = ~n49829 & ~n50631;
  assign n50633 = ~n49707 & n50632;
  assign n50634 = ~n49695 & ~n50633;
  assign n50635 = n49689 & n49705;
  assign n50636 = ~n50634 & ~n50635;
  assign n50637 = n50630 & n50636;
  assign n50638 = n50629 & n50637;
  assign n50639 = ~n49670 & ~n50638;
  assign n50640 = ~n49744 & ~n50461;
  assign n50641 = ~n49695 & ~n50640;
  assign n50642 = ~n50639 & ~n50641;
  assign n50643 = n50625 & n50642;
  assign n50644 = pi1324 & n50643;
  assign n50645 = ~pi1324 & ~n50643;
  assign po1432 = n50644 | n50645;
  assign n50647 = ~n50316 & ~n50502;
  assign n50648 = ~n50294 & n50647;
  assign n50649 = ~n50268 & ~n50648;
  assign n50650 = ~n50509 & ~n50526;
  assign n50651 = ~n50303 & ~n50319;
  assign n50652 = ~n50261 & ~n50308;
  assign n50653 = n50268 & ~n50652;
  assign n50654 = ~n50276 & ~n50653;
  assign n50655 = n50651 & n50654;
  assign n50656 = n50235 & ~n50655;
  assign n50657 = n50247 & n50259;
  assign n50658 = ~n50346 & ~n50657;
  assign n50659 = ~n50241 & ~n50658;
  assign n50660 = ~n50310 & ~n50512;
  assign n50661 = n50268 & ~n50660;
  assign n50662 = ~n50241 & n50259;
  assign n50663 = ~n50293 & ~n50662;
  assign n50664 = ~n50260 & n50663;
  assign n50665 = ~n50268 & ~n50664;
  assign n50666 = ~n50661 & ~n50665;
  assign n50667 = ~n50659 & n50666;
  assign n50668 = ~n50235 & ~n50667;
  assign n50669 = ~n50656 & ~n50668;
  assign n50670 = n50650 & n50669;
  assign n50671 = ~n50649 & n50670;
  assign n50672 = ~pi1347 & ~n50671;
  assign n50673 = pi1347 & n50650;
  assign n50674 = ~n50649 & n50673;
  assign n50675 = n50669 & n50674;
  assign po1433 = n50672 | n50675;
  assign n50677 = pi4402 & ~pi9040;
  assign n50678 = pi4409 & pi9040;
  assign n50679 = ~n50677 & ~n50678;
  assign n50680 = pi1335 & n50679;
  assign n50681 = ~pi1335 & ~n50679;
  assign n50682 = ~n50680 & ~n50681;
  assign n50683 = pi4735 & ~pi9040;
  assign n50684 = pi4521 & pi9040;
  assign n50685 = ~n50683 & ~n50684;
  assign n50686 = ~pi1341 & ~n50685;
  assign n50687 = pi1341 & n50685;
  assign n50688 = ~n50686 & ~n50687;
  assign n50689 = pi4805 & pi9040;
  assign n50690 = pi4490 & ~pi9040;
  assign n50691 = ~n50689 & ~n50690;
  assign n50692 = ~pi1367 & ~n50691;
  assign n50693 = pi1367 & n50691;
  assign n50694 = ~n50692 & ~n50693;
  assign n50695 = pi4482 & ~pi9040;
  assign n50696 = pi4477 & pi9040;
  assign n50697 = ~n50695 & ~n50696;
  assign n50698 = ~pi1346 & n50697;
  assign n50699 = pi1346 & ~n50697;
  assign n50700 = ~n50698 & ~n50699;
  assign n50701 = n50694 & ~n50700;
  assign n50702 = ~n50688 & n50701;
  assign n50703 = pi4553 & ~pi9040;
  assign n50704 = pi4678 & pi9040;
  assign n50705 = ~n50703 & ~n50704;
  assign n50706 = ~pi1373 & n50705;
  assign n50707 = pi1373 & ~n50705;
  assign n50708 = ~n50706 & ~n50707;
  assign n50709 = n50702 & n50708;
  assign n50710 = ~n50694 & n50700;
  assign n50711 = ~n50688 & n50708;
  assign n50712 = n50710 & n50711;
  assign n50713 = ~n50709 & ~n50712;
  assign n50714 = n50688 & ~n50708;
  assign n50715 = n50710 & n50714;
  assign n50716 = ~n50688 & ~n50708;
  assign n50717 = n50700 & n50716;
  assign n50718 = n50694 & n50717;
  assign n50719 = ~n50715 & ~n50718;
  assign n50720 = n50713 & n50719;
  assign n50721 = n50682 & ~n50720;
  assign n50722 = ~n50694 & ~n50700;
  assign n50723 = ~n50688 & n50722;
  assign n50724 = ~n50708 & n50723;
  assign n50725 = n50694 & n50700;
  assign n50726 = ~n50688 & n50725;
  assign n50727 = ~n50724 & ~n50726;
  assign n50728 = n50682 & ~n50727;
  assign n50729 = ~n50682 & ~n50700;
  assign n50730 = n50708 & n50729;
  assign n50731 = n50688 & n50694;
  assign n50732 = ~n50708 & n50710;
  assign n50733 = ~n50731 & ~n50732;
  assign n50734 = ~n50682 & ~n50733;
  assign n50735 = ~n50730 & ~n50734;
  assign n50736 = n50688 & n50722;
  assign n50737 = n50708 & n50736;
  assign n50738 = n50735 & ~n50737;
  assign n50739 = ~n50700 & n50731;
  assign n50740 = ~n50708 & n50739;
  assign n50741 = n50738 & ~n50740;
  assign n50742 = ~n50728 & n50741;
  assign n50743 = ~pi4578 & ~pi9040;
  assign n50744 = ~pi4482 & pi9040;
  assign n50745 = ~n50743 & ~n50744;
  assign n50746 = ~pi1371 & n50745;
  assign n50747 = pi1371 & ~n50745;
  assign n50748 = ~n50746 & ~n50747;
  assign n50749 = ~n50742 & ~n50748;
  assign n50750 = ~n50682 & ~n50708;
  assign n50751 = ~n50688 & ~n50700;
  assign n50752 = n50748 & n50751;
  assign n50753 = n50750 & n50752;
  assign n50754 = n50700 & n50711;
  assign n50755 = ~n50682 & ~n50754;
  assign n50756 = ~n50694 & n50714;
  assign n50757 = ~n50701 & ~n50751;
  assign n50758 = n50708 & ~n50757;
  assign n50759 = n50688 & n50710;
  assign n50760 = ~n50758 & ~n50759;
  assign n50761 = n50682 & n50760;
  assign n50762 = ~n50756 & n50761;
  assign n50763 = ~n50755 & ~n50762;
  assign n50764 = n50688 & n50725;
  assign n50765 = ~n50708 & n50764;
  assign n50766 = ~n50763 & ~n50765;
  assign n50767 = n50748 & ~n50766;
  assign n50768 = ~n50753 & ~n50767;
  assign n50769 = ~n50749 & n50768;
  assign n50770 = ~n50721 & n50769;
  assign n50771 = ~n50682 & n50737;
  assign n50772 = n50770 & ~n50771;
  assign n50773 = pi1384 & ~n50772;
  assign n50774 = n50769 & ~n50771;
  assign n50775 = ~pi1384 & n50774;
  assign n50776 = ~n50721 & n50775;
  assign po1445 = n50773 | n50776;
  assign n50778 = pi4603 & pi9040;
  assign n50779 = pi4479 & ~pi9040;
  assign n50780 = ~n50778 & ~n50779;
  assign n50781 = ~pi1346 & ~n50780;
  assign n50782 = pi1346 & n50780;
  assign n50783 = ~n50781 & ~n50782;
  assign n50784 = pi4730 & ~pi9040;
  assign n50785 = pi4401 & pi9040;
  assign n50786 = ~n50784 & ~n50785;
  assign n50787 = ~pi1363 & ~n50786;
  assign n50788 = pi1363 & n50786;
  assign n50789 = ~n50787 & ~n50788;
  assign n50790 = pi4735 & pi9040;
  assign n50791 = pi4409 & ~pi9040;
  assign n50792 = ~n50790 & ~n50791;
  assign n50793 = ~pi1341 & ~n50792;
  assign n50794 = pi1341 & n50792;
  assign n50795 = ~n50793 & ~n50794;
  assign n50796 = ~n50789 & n50795;
  assign n50797 = pi4561 & pi9040;
  assign n50798 = pi4678 & ~pi9040;
  assign n50799 = ~n50797 & ~n50798;
  assign n50800 = ~pi1345 & n50799;
  assign n50801 = pi1345 & ~n50799;
  assign n50802 = ~n50800 & ~n50801;
  assign n50803 = pi4507 & pi9040;
  assign n50804 = pi4561 & ~pi9040;
  assign n50805 = ~n50803 & ~n50804;
  assign n50806 = pi1370 & n50805;
  assign n50807 = ~pi1370 & ~n50805;
  assign n50808 = ~n50806 & ~n50807;
  assign n50809 = n50802 & ~n50808;
  assign n50810 = n50796 & n50809;
  assign n50811 = pi4483 & pi9040;
  assign n50812 = pi4805 & ~pi9040;
  assign n50813 = ~n50811 & ~n50812;
  assign n50814 = ~pi1358 & n50813;
  assign n50815 = pi1358 & ~n50813;
  assign n50816 = ~n50814 & ~n50815;
  assign n50817 = n50789 & ~n50795;
  assign n50818 = ~n50816 & n50817;
  assign n50819 = ~n50802 & n50816;
  assign n50820 = ~n50795 & n50819;
  assign n50821 = ~n50789 & n50820;
  assign n50822 = ~n50818 & ~n50821;
  assign n50823 = n50789 & n50795;
  assign n50824 = ~n50802 & n50823;
  assign n50825 = n50822 & ~n50824;
  assign n50826 = ~n50808 & ~n50825;
  assign n50827 = n50789 & n50816;
  assign n50828 = n50802 & n50808;
  assign n50829 = n50827 & n50828;
  assign n50830 = n50816 & n50817;
  assign n50831 = n50802 & n50830;
  assign n50832 = ~n50829 & ~n50831;
  assign n50833 = ~n50826 & n50832;
  assign n50834 = ~n50810 & n50833;
  assign n50835 = n50796 & ~n50816;
  assign n50836 = n50802 & n50835;
  assign n50837 = ~n50816 & n50823;
  assign n50838 = ~n50802 & n50837;
  assign n50839 = ~n50836 & ~n50838;
  assign n50840 = n50834 & n50839;
  assign n50841 = ~n50783 & ~n50840;
  assign n50842 = n50795 & n50816;
  assign n50843 = n50802 & n50842;
  assign n50844 = n50789 & n50843;
  assign n50845 = ~n50835 & ~n50844;
  assign n50846 = ~n50808 & ~n50845;
  assign n50847 = n50796 & n50816;
  assign n50848 = ~n50802 & n50847;
  assign n50849 = n50802 & n50816;
  assign n50850 = ~n50795 & n50849;
  assign n50851 = ~n50789 & n50850;
  assign n50852 = ~n50848 & ~n50851;
  assign n50853 = n50789 & n50819;
  assign n50854 = n50802 & n50837;
  assign n50855 = ~n50853 & ~n50854;
  assign n50856 = n50808 & ~n50855;
  assign n50857 = n50852 & ~n50856;
  assign n50858 = ~n50846 & n50857;
  assign n50859 = n50783 & ~n50858;
  assign n50860 = n50789 & ~n50816;
  assign n50861 = ~n50802 & n50860;
  assign n50862 = ~n50789 & ~n50816;
  assign n50863 = n50802 & n50862;
  assign n50864 = ~n50861 & ~n50863;
  assign n50865 = ~n50808 & ~n50864;
  assign n50866 = ~n50789 & ~n50795;
  assign n50867 = ~n50816 & n50866;
  assign n50868 = ~n50802 & n50867;
  assign n50869 = ~n50848 & ~n50868;
  assign n50870 = ~n50830 & n50869;
  assign n50871 = n50808 & ~n50870;
  assign n50872 = ~n50865 & ~n50871;
  assign n50873 = ~n50795 & n50816;
  assign n50874 = n50808 & n50873;
  assign n50875 = n50802 & n50874;
  assign n50876 = n50872 & ~n50875;
  assign n50877 = ~n50859 & n50876;
  assign n50878 = ~n50841 & n50877;
  assign n50879 = pi1377 & n50878;
  assign n50880 = ~pi1377 & ~n50878;
  assign po1454 = n50879 | n50880;
  assign n50882 = ~n50851 & ~n50860;
  assign n50883 = n50808 & ~n50882;
  assign n50884 = ~n50802 & n50830;
  assign n50885 = ~n50883 & ~n50884;
  assign n50886 = ~n50844 & n50885;
  assign n50887 = ~n50808 & n50848;
  assign n50888 = ~n50836 & ~n50887;
  assign n50889 = ~n50868 & n50888;
  assign n50890 = n50886 & n50889;
  assign n50891 = n50783 & ~n50890;
  assign n50892 = n50795 & n50819;
  assign n50893 = n50789 & n50892;
  assign n50894 = ~n50821 & ~n50893;
  assign n50895 = n50808 & n50847;
  assign n50896 = ~n50802 & n50835;
  assign n50897 = ~n50895 & ~n50896;
  assign n50898 = n50795 & ~n50816;
  assign n50899 = n50789 & ~n50802;
  assign n50900 = ~n50898 & ~n50899;
  assign n50901 = ~n50873 & n50900;
  assign n50902 = ~n50808 & ~n50901;
  assign n50903 = n50802 & n50867;
  assign n50904 = ~n50831 & ~n50903;
  assign n50905 = ~n50902 & n50904;
  assign n50906 = n50897 & n50905;
  assign n50907 = n50894 & n50906;
  assign n50908 = ~n50783 & ~n50907;
  assign n50909 = ~n50891 & ~n50908;
  assign n50910 = pi1380 & ~n50909;
  assign n50911 = ~pi1380 & ~n50891;
  assign n50912 = ~n50908 & n50911;
  assign po1457 = n50910 | n50912;
  assign n50914 = pi4393 & pi9040;
  assign n50915 = pi4509 & ~pi9040;
  assign n50916 = ~n50914 & ~n50915;
  assign n50917 = pi1371 & n50916;
  assign n50918 = ~pi1371 & ~n50916;
  assign n50919 = ~n50917 & ~n50918;
  assign n50920 = pi4403 & ~pi9040;
  assign n50921 = pi4650 & pi9040;
  assign n50922 = ~n50920 & ~n50921;
  assign n50923 = ~pi1367 & ~n50922;
  assign n50924 = pi1367 & n50922;
  assign n50925 = ~n50923 & ~n50924;
  assign n50926 = pi4485 & pi9040;
  assign n50927 = pi4852 & ~pi9040;
  assign n50928 = ~n50926 & ~n50927;
  assign n50929 = ~pi1374 & ~n50928;
  assign n50930 = pi1374 & n50928;
  assign n50931 = ~n50929 & ~n50930;
  assign n50932 = n50925 & ~n50931;
  assign n50933 = n50919 & n50932;
  assign n50934 = pi4510 & ~pi9040;
  assign n50935 = pi4492 & pi9040;
  assign n50936 = ~n50934 & ~n50935;
  assign n50937 = pi1355 & n50936;
  assign n50938 = ~pi1355 & ~n50936;
  assign n50939 = ~n50937 & ~n50938;
  assign n50940 = ~n50919 & n50939;
  assign n50941 = ~n50925 & n50940;
  assign n50942 = ~n50933 & ~n50941;
  assign n50943 = pi4718 & pi9040;
  assign n50944 = pi4394 & ~pi9040;
  assign n50945 = ~n50943 & ~n50944;
  assign n50946 = ~pi1339 & n50945;
  assign n50947 = pi1339 & ~n50945;
  assign n50948 = ~n50946 & ~n50947;
  assign n50949 = ~n50919 & ~n50948;
  assign n50950 = ~n50925 & n50949;
  assign n50951 = n50942 & ~n50950;
  assign n50952 = ~pi1339 & ~n50945;
  assign n50953 = pi1339 & n50945;
  assign n50954 = ~n50952 & ~n50953;
  assign n50955 = ~n50925 & ~n50954;
  assign n50956 = n50919 & n50955;
  assign n50957 = ~n50939 & n50956;
  assign n50958 = n50951 & ~n50957;
  assign n50959 = ~n50919 & ~n50954;
  assign n50960 = n50939 & n50959;
  assign n50961 = ~n50925 & ~n50948;
  assign n50962 = ~n50960 & ~n50961;
  assign n50963 = n50931 & ~n50962;
  assign n50964 = n50931 & n50949;
  assign n50965 = ~n50939 & n50964;
  assign n50966 = ~n50963 & ~n50965;
  assign n50967 = n50958 & n50966;
  assign n50968 = pi4396 & ~pi9040;
  assign n50969 = pi4591 & pi9040;
  assign n50970 = ~n50968 & ~n50969;
  assign n50971 = ~pi1356 & ~n50970;
  assign n50972 = pi1356 & n50970;
  assign n50973 = ~n50971 & ~n50972;
  assign n50974 = ~n50967 & n50973;
  assign n50975 = n50919 & ~n50954;
  assign n50976 = ~n50925 & n50975;
  assign n50977 = ~n50931 & n50939;
  assign n50978 = n50976 & n50977;
  assign n50979 = n50925 & ~n50939;
  assign n50980 = ~n50919 & n50979;
  assign n50981 = ~n50939 & n50959;
  assign n50982 = ~n50980 & ~n50981;
  assign n50983 = ~n50931 & ~n50982;
  assign n50984 = ~n50978 & ~n50983;
  assign n50985 = ~n50973 & ~n50984;
  assign n50986 = ~n50925 & n50939;
  assign n50987 = n50931 & n50986;
  assign n50988 = n50959 & n50987;
  assign n50989 = n50948 & n50979;
  assign n50990 = n50919 & n50925;
  assign n50991 = ~n50948 & n50990;
  assign n50992 = n50939 & n50991;
  assign n50993 = ~n50989 & ~n50992;
  assign n50994 = n50939 & n50950;
  assign n50995 = n50993 & ~n50994;
  assign n50996 = ~n50931 & ~n50995;
  assign n50997 = n50931 & n50939;
  assign n50998 = n50949 & n50997;
  assign n50999 = n50925 & n50998;
  assign n51000 = n50919 & ~n50948;
  assign n51001 = n50931 & ~n50939;
  assign n51002 = n51000 & n51001;
  assign n51003 = ~n50954 & n50979;
  assign n51004 = ~n50919 & n51003;
  assign n51005 = n50925 & n50975;
  assign n51006 = n50931 & n51005;
  assign n51007 = n50939 & n51006;
  assign n51008 = ~n51004 & ~n51007;
  assign n51009 = ~n51002 & n51008;
  assign n51010 = ~n50999 & n51009;
  assign n51011 = ~n50925 & ~n50939;
  assign n51012 = ~n50948 & n51011;
  assign n51013 = n50919 & n51012;
  assign n51014 = n51010 & ~n51013;
  assign n51015 = ~n50973 & ~n51014;
  assign n51016 = ~n50996 & ~n51015;
  assign n51017 = ~n50988 & n51016;
  assign n51018 = ~n50985 & n51017;
  assign n51019 = ~n50974 & n51018;
  assign n51020 = n50919 & ~n50925;
  assign n51021 = n51001 & n51020;
  assign n51022 = n51019 & ~n51021;
  assign n51023 = ~pi1382 & ~n51022;
  assign n51024 = pi1382 & ~n51021;
  assign n51025 = n51018 & n51024;
  assign n51026 = ~n50974 & n51025;
  assign po1461 = n51023 | n51026;
  assign n51028 = pi4401 & ~pi9040;
  assign n51029 = pi4553 & pi9040;
  assign n51030 = ~n51028 & ~n51029;
  assign n51031 = ~pi1363 & ~n51030;
  assign n51032 = pi1363 & n51030;
  assign n51033 = ~n51031 & ~n51032;
  assign n51034 = pi4507 & ~pi9040;
  assign n51035 = pi4479 & pi9040;
  assign n51036 = ~n51034 & ~n51035;
  assign n51037 = ~pi1361 & ~n51036;
  assign n51038 = pi1361 & n51036;
  assign n51039 = ~n51037 & ~n51038;
  assign n51040 = pi4475 & pi9040;
  assign n51041 = pi4603 & ~pi9040;
  assign n51042 = ~n51040 & ~n51041;
  assign n51043 = ~pi1334 & ~n51042;
  assign n51044 = pi1334 & n51042;
  assign n51045 = ~n51043 & ~n51044;
  assign n51046 = pi4400 & ~pi9040;
  assign n51047 = pi4615 & pi9040;
  assign n51048 = ~n51046 & ~n51047;
  assign n51049 = ~pi1350 & n51048;
  assign n51050 = pi1350 & ~n51048;
  assign n51051 = ~n51049 & ~n51050;
  assign n51052 = pi4475 & ~pi9040;
  assign n51053 = pi4578 & pi9040;
  assign n51054 = ~n51052 & ~n51053;
  assign n51055 = ~pi1368 & n51054;
  assign n51056 = pi1368 & ~n51054;
  assign n51057 = ~n51055 & ~n51056;
  assign n51058 = n51051 & ~n51057;
  assign n51059 = n51045 & n51058;
  assign n51060 = pi4473 & pi9040;
  assign n51061 = pi4413 & ~pi9040;
  assign n51062 = ~n51060 & ~n51061;
  assign n51063 = ~pi1358 & n51062;
  assign n51064 = pi1358 & ~n51062;
  assign n51065 = ~n51063 & ~n51064;
  assign n51066 = ~n51051 & ~n51065;
  assign n51067 = ~n51057 & n51066;
  assign n51068 = ~n51059 & ~n51067;
  assign n51069 = ~n51045 & n51057;
  assign n51070 = n51065 & n51069;
  assign n51071 = ~n51051 & n51070;
  assign n51072 = n51068 & ~n51071;
  assign n51073 = n51039 & ~n51072;
  assign n51074 = ~n51051 & n51057;
  assign n51075 = ~n51065 & n51074;
  assign n51076 = ~n51045 & n51075;
  assign n51077 = n51051 & ~n51065;
  assign n51078 = ~n51057 & n51077;
  assign n51079 = ~n51045 & n51078;
  assign n51080 = ~n51051 & n51065;
  assign n51081 = n51051 & n51057;
  assign n51082 = ~n51080 & ~n51081;
  assign n51083 = n51045 & ~n51082;
  assign n51084 = ~n51079 & ~n51083;
  assign n51085 = ~n51076 & n51084;
  assign n51086 = ~n51039 & ~n51085;
  assign n51087 = ~n51073 & ~n51086;
  assign n51088 = n51033 & ~n51087;
  assign n51089 = n51039 & ~n51045;
  assign n51090 = n51051 & n51089;
  assign n51091 = ~n51039 & ~n51045;
  assign n51092 = n51080 & n51091;
  assign n51093 = ~n51045 & ~n51051;
  assign n51094 = ~n51057 & n51093;
  assign n51095 = ~n51059 & ~n51094;
  assign n51096 = ~n51039 & ~n51095;
  assign n51097 = ~n51092 & ~n51096;
  assign n51098 = ~n51057 & n51080;
  assign n51099 = ~n51045 & n51098;
  assign n51100 = n51045 & n51075;
  assign n51101 = ~n51099 & ~n51100;
  assign n51102 = n51039 & n51045;
  assign n51103 = n51074 & n51102;
  assign n51104 = n51057 & n51077;
  assign n51105 = n51039 & n51104;
  assign n51106 = ~n51103 & ~n51105;
  assign n51107 = n51101 & n51106;
  assign n51108 = n51097 & n51107;
  assign n51109 = ~n51090 & n51108;
  assign n51110 = ~n51033 & ~n51109;
  assign n51111 = n51051 & n51065;
  assign n51112 = n51057 & n51111;
  assign n51113 = ~n51039 & n51112;
  assign n51114 = ~n51045 & n51113;
  assign n51115 = ~n51039 & n51099;
  assign n51116 = ~n51114 & ~n51115;
  assign n51117 = ~n51065 & n51069;
  assign n51118 = n51051 & n51117;
  assign n51119 = n51039 & n51118;
  assign n51120 = n51116 & ~n51119;
  assign n51121 = ~n51045 & ~n51057;
  assign n51122 = n51065 & n51121;
  assign n51123 = n51051 & n51122;
  assign n51124 = n51045 & n51066;
  assign n51125 = ~n51123 & ~n51124;
  assign n51126 = n51039 & ~n51125;
  assign n51127 = n51120 & ~n51126;
  assign n51128 = ~n51110 & n51127;
  assign n51129 = ~n51088 & n51128;
  assign n51130 = ~pi1376 & ~n51129;
  assign n51131 = pi1376 & n51129;
  assign po1463 = n51130 | n51131;
  assign n51133 = pi4480 & pi9040;
  assign n51134 = pi4602 & ~pi9040;
  assign n51135 = ~n51133 & ~n51134;
  assign n51136 = ~pi1366 & n51135;
  assign n51137 = pi1366 & ~n51135;
  assign n51138 = ~n51136 & ~n51137;
  assign n51139 = pi4711 & ~pi9040;
  assign n51140 = pi4394 & pi9040;
  assign n51141 = ~n51139 & ~n51140;
  assign n51142 = ~pi1352 & ~n51141;
  assign n51143 = pi1352 & n51141;
  assign n51144 = ~n51142 & ~n51143;
  assign n51145 = pi4579 & ~pi9040;
  assign n51146 = pi4481 & pi9040;
  assign n51147 = ~n51145 & ~n51146;
  assign n51148 = ~pi1353 & ~n51147;
  assign n51149 = pi1353 & n51147;
  assign n51150 = ~n51148 & ~n51149;
  assign n51151 = pi4511 & ~pi9040;
  assign n51152 = pi4852 & pi9040;
  assign n51153 = ~n51151 & ~n51152;
  assign n51154 = ~pi1369 & n51153;
  assign n51155 = pi1369 & ~n51153;
  assign n51156 = ~n51154 & ~n51155;
  assign n51157 = pi4711 & pi9040;
  assign n51158 = pi4397 & ~pi9040;
  assign n51159 = ~n51157 & ~n51158;
  assign n51160 = ~pi1365 & n51159;
  assign n51161 = pi1365 & ~n51159;
  assign n51162 = ~n51160 & ~n51161;
  assign n51163 = n51156 & n51162;
  assign n51164 = ~n51150 & n51163;
  assign n51165 = ~n51144 & n51164;
  assign n51166 = n51156 & ~n51162;
  assign n51167 = ~n51150 & n51166;
  assign n51168 = n51144 & n51167;
  assign n51169 = ~n51165 & ~n51168;
  assign n51170 = ~n51138 & ~n51169;
  assign n51171 = ~n51156 & n51162;
  assign n51172 = n51150 & n51171;
  assign n51173 = ~n51144 & n51172;
  assign n51174 = n51138 & n51173;
  assign n51175 = pi4485 & ~pi9040;
  assign n51176 = pi4579 & pi9040;
  assign n51177 = ~n51175 & ~n51176;
  assign n51178 = ~pi1372 & ~n51177;
  assign n51179 = pi1372 & n51177;
  assign n51180 = ~n51178 & ~n51179;
  assign n51181 = n51144 & ~n51150;
  assign n51182 = ~n51156 & n51181;
  assign n51183 = ~n51138 & n51182;
  assign n51184 = ~n51173 & ~n51183;
  assign n51185 = n51144 & n51162;
  assign n51186 = n51156 & n51185;
  assign n51187 = ~n51144 & n51171;
  assign n51188 = ~n51186 & ~n51187;
  assign n51189 = n51138 & ~n51188;
  assign n51190 = ~n51144 & ~n51150;
  assign n51191 = n51138 & ~n51162;
  assign n51192 = n51190 & n51191;
  assign n51193 = n51156 & n51192;
  assign n51194 = ~n51156 & ~n51162;
  assign n51195 = n51150 & n51194;
  assign n51196 = n51144 & n51195;
  assign n51197 = ~n51144 & n51150;
  assign n51198 = n51156 & n51197;
  assign n51199 = ~n51138 & n51198;
  assign n51200 = ~n51196 & ~n51199;
  assign n51201 = ~n51193 & n51200;
  assign n51202 = ~n51189 & n51201;
  assign n51203 = n51184 & n51202;
  assign n51204 = n51180 & ~n51203;
  assign n51205 = n51162 & n51183;
  assign n51206 = ~n51204 & ~n51205;
  assign n51207 = ~n51174 & n51206;
  assign n51208 = ~n51170 & n51207;
  assign n51209 = ~n51138 & ~n51162;
  assign n51210 = ~n51144 & ~n51156;
  assign n51211 = n51209 & n51210;
  assign n51212 = n51156 & n51190;
  assign n51213 = ~n51138 & n51212;
  assign n51214 = ~n51211 & ~n51213;
  assign n51215 = n51144 & n51150;
  assign n51216 = ~n51156 & n51215;
  assign n51217 = ~n51138 & n51216;
  assign n51218 = n51156 & n51215;
  assign n51219 = n51162 & n51218;
  assign n51220 = ~n51217 & ~n51219;
  assign n51221 = ~n51162 & n51181;
  assign n51222 = n51150 & n51156;
  assign n51223 = ~n51221 & ~n51222;
  assign n51224 = n51138 & ~n51223;
  assign n51225 = ~n51156 & n51190;
  assign n51226 = ~n51162 & n51225;
  assign n51227 = ~n51165 & ~n51226;
  assign n51228 = ~n51224 & n51227;
  assign n51229 = n51220 & n51228;
  assign n51230 = n51214 & n51229;
  assign n51231 = ~n51180 & ~n51230;
  assign n51232 = n51208 & ~n51231;
  assign n51233 = ~pi1383 & ~n51232;
  assign n51234 = pi1383 & n51208;
  assign n51235 = ~n51231 & n51234;
  assign po1465 = n51233 | n51235;
  assign n51237 = pi4402 & pi9040;
  assign n51238 = pi4615 & ~pi9040;
  assign n51239 = ~n51237 & ~n51238;
  assign n51240 = ~pi1350 & ~n51239;
  assign n51241 = pi1350 & n51239;
  assign n51242 = ~n51240 & ~n51241;
  assign n51243 = pi4413 & pi9040;
  assign n51244 = pi4521 & ~pi9040;
  assign n51245 = ~n51243 & ~n51244;
  assign n51246 = pi1375 & n51245;
  assign n51247 = ~pi1375 & ~n51245;
  assign n51248 = ~n51246 & ~n51247;
  assign n51249 = pi4400 & pi9040;
  assign n51250 = pi4506 & ~pi9040;
  assign n51251 = ~n51249 & ~n51250;
  assign n51252 = pi1372 & n51251;
  assign n51253 = ~pi1372 & ~n51251;
  assign n51254 = ~n51252 & ~n51253;
  assign n51255 = pi4512 & ~pi9040;
  assign n51256 = pi4506 & pi9040;
  assign n51257 = ~n51255 & ~n51256;
  assign n51258 = ~pi1353 & ~n51257;
  assign n51259 = pi1353 & n51257;
  assign n51260 = ~n51258 & ~n51259;
  assign n51261 = pi4730 & pi9040;
  assign n51262 = pi4381 & ~pi9040;
  assign n51263 = ~n51261 & ~n51262;
  assign n51264 = ~pi1368 & ~n51263;
  assign n51265 = pi1368 & n51263;
  assign n51266 = ~n51264 & ~n51265;
  assign n51267 = n51260 & ~n51266;
  assign n51268 = n51254 & n51267;
  assign n51269 = n51248 & n51268;
  assign n51270 = pi4473 & ~pi9040;
  assign n51271 = pi4408 & pi9040;
  assign n51272 = ~n51270 & ~n51271;
  assign n51273 = ~pi1360 & n51272;
  assign n51274 = pi1360 & ~n51272;
  assign n51275 = ~n51273 & ~n51274;
  assign n51276 = n51254 & n51266;
  assign n51277 = n51260 & n51276;
  assign n51278 = ~n51254 & ~n51260;
  assign n51279 = ~n51260 & ~n51266;
  assign n51280 = ~n51248 & n51279;
  assign n51281 = ~n51254 & ~n51266;
  assign n51282 = n51248 & n51281;
  assign n51283 = ~n51280 & ~n51282;
  assign n51284 = ~n51278 & n51283;
  assign n51285 = ~n51277 & n51284;
  assign n51286 = ~n51275 & ~n51285;
  assign n51287 = ~n51248 & n51260;
  assign n51288 = n51266 & n51287;
  assign n51289 = ~n51254 & n51287;
  assign n51290 = ~n51260 & n51276;
  assign n51291 = ~n51289 & ~n51290;
  assign n51292 = n51275 & ~n51291;
  assign n51293 = ~n51288 & ~n51292;
  assign n51294 = ~n51286 & n51293;
  assign n51295 = ~n51269 & n51294;
  assign n51296 = n51242 & ~n51295;
  assign n51297 = ~n51254 & n51266;
  assign n51298 = ~n51260 & n51297;
  assign n51299 = ~n51248 & n51298;
  assign n51300 = ~n51260 & n51281;
  assign n51301 = n51248 & n51300;
  assign n51302 = ~n51269 & ~n51301;
  assign n51303 = ~n51299 & n51302;
  assign n51304 = ~n51275 & ~n51303;
  assign n51305 = ~n51296 & ~n51304;
  assign n51306 = n51254 & n51288;
  assign n51307 = n51254 & ~n51260;
  assign n51308 = n51275 & n51307;
  assign n51309 = n51248 & n51308;
  assign n51310 = n51248 & n51260;
  assign n51311 = n51266 & n51310;
  assign n51312 = ~n51254 & n51311;
  assign n51313 = n51267 & ~n51275;
  assign n51314 = ~n51248 & n51313;
  assign n51315 = ~n51312 & ~n51314;
  assign n51316 = ~n51254 & n51260;
  assign n51317 = n51248 & n51316;
  assign n51318 = n51254 & ~n51266;
  assign n51319 = ~n51260 & n51318;
  assign n51320 = ~n51317 & ~n51319;
  assign n51321 = n51275 & ~n51320;
  assign n51322 = n51275 & n51278;
  assign n51323 = ~n51248 & n51322;
  assign n51324 = ~n51321 & ~n51323;
  assign n51325 = n51315 & n51324;
  assign n51326 = ~n51242 & ~n51325;
  assign n51327 = ~n51309 & ~n51326;
  assign n51328 = ~n51306 & n51327;
  assign n51329 = n51305 & n51328;
  assign n51330 = ~pi1381 & ~n51329;
  assign n51331 = ~n51296 & ~n51306;
  assign n51332 = ~n51304 & n51331;
  assign n51333 = n51327 & n51332;
  assign n51334 = pi1381 & n51333;
  assign po1466 = n51330 | n51334;
  assign n51336 = ~n51156 & n51197;
  assign n51337 = ~n51162 & n51336;
  assign n51338 = ~n51162 & n51215;
  assign n51339 = n51162 & n51198;
  assign n51340 = ~n51338 & ~n51339;
  assign n51341 = n51138 & ~n51340;
  assign n51342 = ~n51337 & ~n51341;
  assign n51343 = ~n51138 & n51197;
  assign n51344 = ~n51162 & n51343;
  assign n51345 = ~n51213 & ~n51344;
  assign n51346 = n51342 & n51345;
  assign n51347 = ~n51162 & n51182;
  assign n51348 = n51162 & n51225;
  assign n51349 = ~n51347 & ~n51348;
  assign n51350 = n51346 & n51349;
  assign n51351 = n51180 & ~n51350;
  assign n51352 = n51138 & ~n51180;
  assign n51353 = ~n51144 & n51166;
  assign n51354 = ~n51150 & n51156;
  assign n51355 = ~n51353 & ~n51354;
  assign n51356 = n51352 & ~n51355;
  assign n51357 = ~n51173 & ~n51186;
  assign n51358 = ~n51156 & n51209;
  assign n51359 = ~n51197 & n51358;
  assign n51360 = ~n51183 & ~n51359;
  assign n51361 = n51357 & n51360;
  assign n51362 = ~n51180 & ~n51361;
  assign n51363 = n51156 & n51181;
  assign n51364 = n51138 & n51363;
  assign n51365 = n51162 & n51364;
  assign n51366 = n51162 & n51216;
  assign n51367 = ~n51348 & ~n51366;
  assign n51368 = n51138 & ~n51367;
  assign n51369 = ~n51365 & ~n51368;
  assign n51370 = ~n51138 & n51173;
  assign n51371 = n51369 & ~n51370;
  assign n51372 = ~n51362 & n51371;
  assign n51373 = ~n51356 & n51372;
  assign n51374 = ~n51351 & n51373;
  assign n51375 = ~n51138 & n51162;
  assign n51376 = n51218 & n51375;
  assign n51377 = n51374 & ~n51376;
  assign n51378 = ~pi1386 & ~n51377;
  assign n51379 = n51373 & ~n51376;
  assign n51380 = pi1386 & n51379;
  assign n51381 = ~n51351 & n51380;
  assign po1467 = n51378 | n51381;
  assign n51383 = ~n51033 & ~n51039;
  assign n51384 = ~n51045 & n51058;
  assign n51385 = n51045 & n51098;
  assign n51386 = ~n51045 & n51066;
  assign n51387 = ~n51385 & ~n51386;
  assign n51388 = ~n51384 & n51387;
  assign n51389 = n51383 & ~n51388;
  assign n51390 = ~n51057 & n51111;
  assign n51391 = n51045 & n51390;
  assign n51392 = ~n51070 & ~n51391;
  assign n51393 = n51057 & n51080;
  assign n51394 = ~n51067 & ~n51393;
  assign n51395 = n51392 & n51394;
  assign n51396 = n51039 & ~n51395;
  assign n51397 = n51045 & n51104;
  assign n51398 = ~n51396 & ~n51397;
  assign n51399 = ~n51033 & ~n51398;
  assign n51400 = ~n51389 & ~n51399;
  assign n51401 = ~n51057 & n51089;
  assign n51402 = ~n51065 & n51401;
  assign n51403 = ~n51071 & ~n51402;
  assign n51404 = ~n51066 & ~n51111;
  assign n51405 = n51045 & ~n51404;
  assign n51406 = ~n51112 & ~n51405;
  assign n51407 = ~n51039 & ~n51406;
  assign n51408 = ~n51078 & ~n51384;
  assign n51409 = ~n51385 & n51408;
  assign n51410 = n51039 & ~n51409;
  assign n51411 = ~n51407 & ~n51410;
  assign n51412 = n51045 & n51112;
  assign n51413 = ~n51100 & ~n51412;
  assign n51414 = ~n51118 & n51413;
  assign n51415 = ~n51092 & n51414;
  assign n51416 = n51411 & n51415;
  assign n51417 = n51033 & ~n51416;
  assign n51418 = n51403 & ~n51417;
  assign n51419 = n51400 & n51418;
  assign n51420 = pi1378 & ~n51419;
  assign n51421 = ~pi1378 & n51403;
  assign n51422 = n51400 & n51421;
  assign n51423 = ~n51417 & n51422;
  assign po1473 = n51420 | n51423;
  assign n51425 = ~n50688 & n50694;
  assign n51426 = ~n50682 & n51425;
  assign n51427 = ~n50708 & n51426;
  assign n51428 = ~n50700 & n50716;
  assign n51429 = n50694 & n51428;
  assign n51430 = n50688 & ~n50700;
  assign n51431 = n50708 & n51430;
  assign n51432 = ~n50715 & ~n51431;
  assign n51433 = ~n51429 & n51432;
  assign n51434 = ~n51427 & n51433;
  assign n51435 = ~n50688 & n50710;
  assign n51436 = n50682 & n51435;
  assign n51437 = n51434 & ~n51436;
  assign n51438 = n50748 & ~n51437;
  assign n51439 = n50694 & n50711;
  assign n51440 = n50700 & n51439;
  assign n51441 = ~n50765 & ~n51440;
  assign n51442 = n50682 & ~n51441;
  assign n51443 = ~n50682 & ~n50748;
  assign n51444 = n50751 & n51443;
  assign n51445 = n50688 & n50708;
  assign n51446 = ~n50694 & n51445;
  assign n51447 = ~n51430 & ~n51446;
  assign n51448 = ~n50726 & n51447;
  assign n51449 = n50682 & ~n51448;
  assign n51450 = n50708 & n50723;
  assign n51451 = ~n51449 & ~n51450;
  assign n51452 = ~n50748 & ~n51451;
  assign n51453 = ~n51444 & ~n51452;
  assign n51454 = ~n51442 & n51453;
  assign n51455 = ~n50708 & n50751;
  assign n51456 = n50708 & n50764;
  assign n51457 = ~n51455 & ~n51456;
  assign n51458 = ~n50712 & n51457;
  assign n51459 = ~n50715 & n51458;
  assign n51460 = ~n50682 & ~n51459;
  assign n51461 = n51454 & ~n51460;
  assign n51462 = ~n51438 & n51461;
  assign n51463 = ~pi1417 & ~n51462;
  assign n51464 = pi1417 & n51454;
  assign n51465 = ~n51438 & n51464;
  assign n51466 = ~n51460 & n51465;
  assign po1474 = n51463 | n51466;
  assign n51468 = n50708 & n50739;
  assign n51469 = ~n50736 & ~n51455;
  assign n51470 = n50682 & ~n51469;
  assign n51471 = ~n51468 & ~n51470;
  assign n51472 = ~n50682 & n50759;
  assign n51473 = ~n50682 & n50708;
  assign n51474 = ~n50700 & n51473;
  assign n51475 = n50694 & n51474;
  assign n51476 = n50725 & n50750;
  assign n51477 = ~n51475 & ~n51476;
  assign n51478 = ~n51472 & n51477;
  assign n51479 = n50708 & n51435;
  assign n51480 = ~n50724 & ~n51479;
  assign n51481 = n50700 & n50714;
  assign n51482 = n51480 & ~n51481;
  assign n51483 = n51478 & n51482;
  assign n51484 = n51471 & n51483;
  assign n51485 = ~n50748 & ~n51484;
  assign n51486 = ~n50736 & ~n51435;
  assign n51487 = ~n50708 & ~n51486;
  assign n51488 = n50682 & n50754;
  assign n51489 = ~n50708 & n51430;
  assign n51490 = ~n50764 & ~n51439;
  assign n51491 = ~n51489 & n51490;
  assign n51492 = n50682 & ~n51491;
  assign n51493 = ~n51488 & ~n51492;
  assign n51494 = n50708 & n50722;
  assign n51495 = ~n51429 & ~n51494;
  assign n51496 = ~n50682 & ~n51495;
  assign n51497 = n51493 & ~n51496;
  assign n51498 = ~n51487 & n51497;
  assign n51499 = ~n51440 & n51498;
  assign n51500 = ~n50748 & ~n51488;
  assign n51501 = ~n51499 & ~n51500;
  assign n51502 = ~n50682 & n51468;
  assign n51503 = ~n51501 & ~n51502;
  assign n51504 = ~n51485 & n51503;
  assign n51505 = ~pi1403 & ~n51504;
  assign n51506 = pi1403 & ~n51501;
  assign n51507 = ~n51485 & n51506;
  assign n51508 = ~n51502 & n51507;
  assign po1475 = n51505 | n51508;
  assign n51510 = pi4494 & ~pi9040;
  assign n51511 = pi4425 & pi9040;
  assign n51512 = ~n51510 & ~n51511;
  assign n51513 = ~pi1357 & ~n51512;
  assign n51514 = pi1357 & n51512;
  assign n51515 = ~n51513 & ~n51514;
  assign n51516 = pi4508 & ~pi9040;
  assign n51517 = pi4583 & pi9040;
  assign n51518 = ~n51516 & ~n51517;
  assign n51519 = pi1359 & n51518;
  assign n51520 = ~pi1359 & ~n51518;
  assign n51521 = ~n51519 & ~n51520;
  assign n51522 = pi4403 & pi9040;
  assign n51523 = pi4492 & ~pi9040;
  assign n51524 = ~n51522 & ~n51523;
  assign n51525 = ~pi1339 & n51524;
  assign n51526 = pi1339 & ~n51524;
  assign n51527 = ~n51525 & ~n51526;
  assign n51528 = pi4393 & ~pi9040;
  assign n51529 = pi4602 & pi9040;
  assign n51530 = ~n51528 & ~n51529;
  assign n51531 = ~pi1356 & ~n51530;
  assign n51532 = pi1356 & n51530;
  assign n51533 = ~n51531 & ~n51532;
  assign n51534 = pi4425 & ~pi9040;
  assign n51535 = pi4397 & pi9040;
  assign n51536 = ~n51534 & ~n51535;
  assign n51537 = ~pi1364 & ~n51536;
  assign n51538 = pi1364 & n51536;
  assign n51539 = ~n51537 & ~n51538;
  assign n51540 = ~n51533 & n51539;
  assign n51541 = n51527 & n51540;
  assign n51542 = n51521 & n51541;
  assign n51543 = pi4385 & pi9040;
  assign n51544 = pi4650 & ~pi9040;
  assign n51545 = ~n51543 & ~n51544;
  assign n51546 = ~pi1362 & ~n51545;
  assign n51547 = pi1362 & n51545;
  assign n51548 = ~n51546 & ~n51547;
  assign n51549 = ~n51521 & n51548;
  assign n51550 = n51533 & n51549;
  assign n51551 = n51533 & ~n51539;
  assign n51552 = n51527 & n51551;
  assign n51553 = n51533 & n51539;
  assign n51554 = ~n51527 & n51553;
  assign n51555 = ~n51552 & ~n51554;
  assign n51556 = ~n51533 & ~n51539;
  assign n51557 = ~n51527 & n51556;
  assign n51558 = n51521 & n51557;
  assign n51559 = n51555 & ~n51558;
  assign n51560 = n51548 & ~n51559;
  assign n51561 = ~n51550 & ~n51560;
  assign n51562 = ~n51542 & n51561;
  assign n51563 = ~n51521 & n51556;
  assign n51564 = ~n51527 & n51540;
  assign n51565 = ~n51563 & ~n51564;
  assign n51566 = ~n51548 & ~n51565;
  assign n51567 = n51527 & n51553;
  assign n51568 = ~n51521 & n51567;
  assign n51569 = ~n51566 & ~n51568;
  assign n51570 = n51562 & n51569;
  assign n51571 = n51515 & ~n51570;
  assign n51572 = ~n51515 & n51548;
  assign n51573 = ~n51565 & n51572;
  assign n51574 = ~n51527 & n51533;
  assign n51575 = ~n51521 & n51551;
  assign n51576 = ~n51541 & ~n51575;
  assign n51577 = ~n51574 & n51576;
  assign n51578 = ~n51515 & ~n51548;
  assign n51579 = ~n51577 & n51578;
  assign n51580 = ~n51573 & ~n51579;
  assign n51581 = n51521 & n51527;
  assign n51582 = ~n51533 & n51581;
  assign n51583 = n51521 & ~n51527;
  assign n51584 = n51551 & n51583;
  assign n51585 = ~n51582 & ~n51584;
  assign n51586 = ~n51548 & ~n51585;
  assign n51587 = n51527 & n51556;
  assign n51588 = ~n51567 & ~n51587;
  assign n51589 = n51521 & ~n51588;
  assign n51590 = ~n51584 & ~n51589;
  assign n51591 = ~n51515 & ~n51590;
  assign n51592 = ~n51586 & ~n51591;
  assign n51593 = n51580 & n51592;
  assign n51594 = ~n51571 & n51593;
  assign n51595 = ~pi1394 & ~n51594;
  assign n51596 = ~n51571 & ~n51586;
  assign n51597 = ~n51573 & ~n51591;
  assign n51598 = pi1394 & n51597;
  assign n51599 = n51596 & n51598;
  assign n51600 = ~n51579 & n51599;
  assign po1476 = n51595 | n51600;
  assign n51602 = n51260 & n51281;
  assign n51603 = n51248 & n51602;
  assign n51604 = n51248 & n51298;
  assign n51605 = ~n51603 & ~n51604;
  assign n51606 = ~n51248 & n51300;
  assign n51607 = ~n51290 & ~n51606;
  assign n51608 = ~n51275 & ~n51607;
  assign n51609 = n51605 & ~n51608;
  assign n51610 = ~n51248 & n51275;
  assign n51611 = n51254 & n51610;
  assign n51612 = n51609 & ~n51611;
  assign n51613 = n51242 & ~n51612;
  assign n51614 = n51248 & n51319;
  assign n51615 = n51275 & n51614;
  assign n51616 = ~n51248 & ~n51275;
  assign n51617 = n51319 & n51616;
  assign n51618 = ~n51289 & ~n51617;
  assign n51619 = n51260 & n51297;
  assign n51620 = ~n51290 & ~n51619;
  assign n51621 = ~n51248 & n51297;
  assign n51622 = n51620 & ~n51621;
  assign n51623 = n51275 & ~n51622;
  assign n51624 = ~n51275 & n51277;
  assign n51625 = n51302 & ~n51624;
  assign n51626 = ~n51623 & n51625;
  assign n51627 = n51618 & n51626;
  assign n51628 = ~n51242 & ~n51627;
  assign n51629 = ~n51615 & ~n51628;
  assign n51630 = ~n51613 & n51629;
  assign n51631 = n51616 & n51619;
  assign n51632 = n51248 & n51313;
  assign n51633 = ~n51631 & ~n51632;
  assign n51634 = ~n51275 & n51604;
  assign n51635 = n51633 & ~n51634;
  assign n51636 = n51630 & n51635;
  assign n51637 = ~pi1379 & ~n51636;
  assign n51638 = pi1379 & n51635;
  assign n51639 = n51629 & n51638;
  assign n51640 = ~n51613 & n51639;
  assign po1477 = n51637 | n51640;
  assign n51642 = ~n50709 & ~n50715;
  assign n51643 = ~n50682 & ~n51642;
  assign n51644 = ~n50771 & ~n51643;
  assign n51645 = ~n50688 & ~n50694;
  assign n51646 = n50682 & n51645;
  assign n51647 = ~n50708 & n51646;
  assign n51648 = ~n50708 & n50722;
  assign n51649 = ~n51645 & ~n51648;
  assign n51650 = n50694 & n51445;
  assign n51651 = n51649 & ~n51650;
  assign n51652 = n50682 & ~n51651;
  assign n51653 = ~n50718 & ~n51652;
  assign n51654 = ~n50748 & ~n51653;
  assign n51655 = ~n50682 & n50701;
  assign n51656 = ~n50708 & n51655;
  assign n51657 = ~n51472 & ~n51656;
  assign n51658 = ~n50748 & ~n51657;
  assign n51659 = ~n51654 & ~n51658;
  assign n51660 = ~n51647 & n51659;
  assign n51661 = ~n50736 & ~n50754;
  assign n51662 = ~n50764 & n51661;
  assign n51663 = ~n50682 & ~n51662;
  assign n51664 = n50708 & n50759;
  assign n51665 = ~n50739 & ~n51664;
  assign n51666 = n50682 & ~n51665;
  assign n51667 = ~n51663 & ~n51666;
  assign n51668 = ~n51439 & n51667;
  assign n51669 = ~n50724 & ~n50765;
  assign n51670 = n51668 & n51669;
  assign n51671 = n50748 & ~n51670;
  assign n51672 = n51660 & ~n51671;
  assign n51673 = n51644 & n51672;
  assign n51674 = ~pi1425 & ~n51673;
  assign n51675 = pi1425 & n51660;
  assign n51676 = n51644 & n51675;
  assign n51677 = ~n51671 & n51676;
  assign po1479 = n51674 | n51677;
  assign n51679 = n50802 & n50823;
  assign n51680 = ~n50903 & ~n51679;
  assign n51681 = n50808 & n51680;
  assign n51682 = ~n50796 & ~n50817;
  assign n51683 = ~n50816 & ~n51682;
  assign n51684 = ~n50802 & n50862;
  assign n51685 = ~n50789 & n50849;
  assign n51686 = ~n50802 & n50817;
  assign n51687 = ~n51685 & ~n51686;
  assign n51688 = ~n51684 & n51687;
  assign n51689 = ~n51683 & n51688;
  assign n51690 = ~n50808 & n51689;
  assign n51691 = ~n51681 & ~n51690;
  assign n51692 = ~n50802 & n51683;
  assign n51693 = ~n50893 & ~n51692;
  assign n51694 = ~n51691 & n51693;
  assign n51695 = n50783 & ~n51694;
  assign n51696 = n50808 & ~n51682;
  assign n51697 = n50802 & n51696;
  assign n51698 = ~n50837 & ~n50866;
  assign n51699 = ~n50802 & ~n51698;
  assign n51700 = n50808 & n51699;
  assign n51701 = n50816 & n51696;
  assign n51702 = ~n51700 & ~n51701;
  assign n51703 = ~n51697 & n51702;
  assign n51704 = ~n50783 & ~n51703;
  assign n51705 = ~n51695 & ~n51704;
  assign n51706 = n50808 & n50821;
  assign n51707 = ~n50808 & ~n51693;
  assign n51708 = ~n51706 & ~n51707;
  assign n51709 = ~n50808 & ~n51680;
  assign n51710 = ~n50821 & ~n51709;
  assign n51711 = ~n50783 & ~n51710;
  assign n51712 = n51708 & ~n51711;
  assign n51713 = n51705 & n51712;
  assign n51714 = pi1387 & ~n51713;
  assign n51715 = ~pi1387 & n51712;
  assign n51716 = ~n51704 & n51715;
  assign n51717 = ~n51695 & n51716;
  assign po1480 = n51714 | n51717;
  assign n51719 = n51521 & ~n51548;
  assign n51720 = ~n51556 & ~n51567;
  assign n51721 = n51719 & ~n51720;
  assign n51722 = n51527 & ~n51548;
  assign n51723 = n51556 & n51722;
  assign n51724 = ~n51721 & ~n51723;
  assign n51725 = n51515 & ~n51724;
  assign n51726 = ~n51521 & ~n51527;
  assign n51727 = n51539 & n51726;
  assign n51728 = n51533 & n51727;
  assign n51729 = ~n51574 & ~n51726;
  assign n51730 = n51548 & ~n51729;
  assign n51731 = ~n51521 & n51527;
  assign n51732 = ~n51539 & n51731;
  assign n51733 = n51533 & n51732;
  assign n51734 = ~n51730 & ~n51733;
  assign n51735 = ~n51728 & n51734;
  assign n51736 = n51515 & ~n51735;
  assign n51737 = ~n51725 & ~n51736;
  assign n51738 = n51539 & n51583;
  assign n51739 = ~n51533 & n51738;
  assign n51740 = ~n51521 & n51541;
  assign n51741 = ~n51739 & ~n51740;
  assign n51742 = ~n51548 & ~n51741;
  assign n51743 = ~n51527 & ~n51539;
  assign n51744 = ~n51541 & ~n51743;
  assign n51745 = ~n51521 & ~n51744;
  assign n51746 = ~n51521 & n51539;
  assign n51747 = n51722 & n51746;
  assign n51748 = ~n51551 & ~n51574;
  assign n51749 = n51521 & ~n51748;
  assign n51750 = ~n51541 & ~n51749;
  assign n51751 = ~n51548 & ~n51750;
  assign n51752 = n51521 & n51548;
  assign n51753 = n51553 & n51752;
  assign n51754 = n51527 & n51753;
  assign n51755 = ~n51751 & ~n51754;
  assign n51756 = ~n51747 & n51755;
  assign n51757 = ~n51745 & n51756;
  assign n51758 = ~n51739 & n51757;
  assign n51759 = ~n51515 & ~n51758;
  assign n51760 = n51521 & n51587;
  assign n51761 = ~n51521 & n51574;
  assign n51762 = ~n51760 & ~n51761;
  assign n51763 = n51548 & ~n51762;
  assign n51764 = ~n51759 & ~n51763;
  assign n51765 = ~n51742 & n51764;
  assign n51766 = n51737 & n51765;
  assign n51767 = pi1390 & n51766;
  assign n51768 = ~pi1390 & ~n51766;
  assign po1481 = n51767 | n51768;
  assign n51770 = n51039 & n51066;
  assign n51771 = ~n51045 & n51770;
  assign n51772 = ~n51123 & ~n51771;
  assign n51773 = n51045 & ~n51065;
  assign n51774 = ~n51057 & n51773;
  assign n51775 = ~n51045 & n51051;
  assign n51776 = ~n51122 & ~n51775;
  assign n51777 = ~n51039 & ~n51776;
  assign n51778 = ~n51774 & ~n51777;
  assign n51779 = n51772 & n51778;
  assign n51780 = n51033 & ~n51779;
  assign n51781 = ~n51098 & ~n51100;
  assign n51782 = ~n51045 & n51077;
  assign n51783 = n51781 & ~n51782;
  assign n51784 = n51039 & ~n51783;
  assign n51785 = n51066 & n51091;
  assign n51786 = ~n51071 & ~n51785;
  assign n51787 = ~n51784 & n51786;
  assign n51788 = ~n51390 & ~n51397;
  assign n51789 = ~n51039 & ~n51788;
  assign n51790 = n51787 & ~n51789;
  assign n51791 = ~n51033 & ~n51790;
  assign n51792 = ~n51780 & ~n51791;
  assign n51793 = ~n51045 & n51111;
  assign n51794 = n51045 & ~n51394;
  assign n51795 = ~n51793 & ~n51794;
  assign n51796 = ~n51039 & ~n51795;
  assign n51797 = ~n51078 & ~n51112;
  assign n51798 = ~n51098 & n51797;
  assign n51799 = n51102 & ~n51798;
  assign n51800 = ~n51796 & ~n51799;
  assign n51801 = n51792 & n51800;
  assign n51802 = ~pi1385 & ~n51801;
  assign n51803 = ~n51791 & n51800;
  assign n51804 = pi1385 & n51803;
  assign n51805 = ~n51780 & n51804;
  assign po1482 = n51802 | n51805;
  assign n51807 = n51162 & n51343;
  assign n51808 = n51144 & n51166;
  assign n51809 = ~n51363 & ~n51808;
  assign n51810 = ~n51138 & ~n51809;
  assign n51811 = ~n51807 & ~n51810;
  assign n51812 = n51138 & n51162;
  assign n51813 = n51215 & n51812;
  assign n51814 = n51138 & n51212;
  assign n51815 = ~n51813 & ~n51814;
  assign n51816 = n51811 & n51815;
  assign n51817 = n51144 & n51171;
  assign n51818 = ~n51165 & ~n51817;
  assign n51819 = ~n51226 & n51818;
  assign n51820 = n51816 & n51819;
  assign n51821 = ~n51180 & ~n51820;
  assign n51822 = ~n51205 & ~n51211;
  assign n51823 = ~n51173 & ~n51363;
  assign n51824 = ~n51221 & n51823;
  assign n51825 = n51138 & ~n51824;
  assign n51826 = ~n51162 & n51198;
  assign n51827 = ~n51196 & ~n51826;
  assign n51828 = ~n51376 & n51827;
  assign n51829 = ~n51138 & n51225;
  assign n51830 = n51828 & ~n51829;
  assign n51831 = ~n51825 & n51830;
  assign n51832 = n51180 & ~n51831;
  assign n51833 = ~n51165 & n51827;
  assign n51834 = n51138 & ~n51833;
  assign n51835 = ~n51832 & ~n51834;
  assign n51836 = n51822 & n51835;
  assign n51837 = ~n51821 & n51836;
  assign n51838 = pi1393 & ~n51837;
  assign n51839 = ~pi1393 & n51837;
  assign po1483 = n51838 | n51839;
  assign n51841 = ~n51347 & ~n51353;
  assign n51842 = n51180 & ~n51841;
  assign n51843 = ~n51172 & ~n51187;
  assign n51844 = ~n51336 & n51843;
  assign n51845 = n51138 & ~n51844;
  assign n51846 = n51180 & n51845;
  assign n51847 = ~n51842 & ~n51846;
  assign n51848 = n51182 & n51191;
  assign n51849 = ~n51193 & ~n51848;
  assign n51850 = ~n51186 & ~n51222;
  assign n51851 = ~n51138 & ~n51850;
  assign n51852 = n51180 & n51851;
  assign n51853 = n51849 & ~n51852;
  assign n51854 = n51162 & n51182;
  assign n51855 = n51162 & n51190;
  assign n51856 = ~n51168 & ~n51855;
  assign n51857 = ~n51138 & ~n51856;
  assign n51858 = ~n51173 & ~n51196;
  assign n51859 = n51162 & n51181;
  assign n51860 = ~n51218 & ~n51859;
  assign n51861 = n51138 & ~n51860;
  assign n51862 = n51858 & ~n51861;
  assign n51863 = ~n51857 & n51862;
  assign n51864 = ~n51854 & n51863;
  assign n51865 = ~n51180 & ~n51864;
  assign n51866 = ~n51226 & n51827;
  assign n51867 = ~n51138 & ~n51866;
  assign n51868 = ~n51865 & ~n51867;
  assign n51869 = n51853 & n51868;
  assign n51870 = n51847 & n51869;
  assign n51871 = ~pi1402 & ~n51870;
  assign n51872 = pi1402 & n51853;
  assign n51873 = n51847 & n51872;
  assign n51874 = n51868 & n51873;
  assign po1484 = n51871 | n51874;
  assign n51876 = n50808 & n50848;
  assign n51877 = n50849 & ~n51682;
  assign n51878 = ~n50867 & ~n51877;
  assign n51879 = ~n50893 & n51878;
  assign n51880 = ~n50808 & ~n51879;
  assign n51881 = ~n50802 & n50818;
  assign n51882 = ~n51880 & ~n51881;
  assign n51883 = n50816 & n50866;
  assign n51884 = n50802 & n50898;
  assign n51885 = ~n51883 & ~n51884;
  assign n51886 = ~n51686 & n51885;
  assign n51887 = n50808 & ~n51886;
  assign n51888 = n51882 & ~n51887;
  assign n51889 = n50783 & ~n51888;
  assign n51890 = ~n51876 & ~n51889;
  assign n51891 = n50802 & n50817;
  assign n51892 = n50816 & n50823;
  assign n51893 = ~n51891 & ~n51892;
  assign n51894 = n50808 & ~n51893;
  assign n51895 = ~n50868 & ~n51894;
  assign n51896 = ~n50838 & ~n50848;
  assign n51897 = ~n50802 & n50873;
  assign n51898 = ~n50898 & ~n51897;
  assign n51899 = ~n51883 & n51898;
  assign n51900 = ~n50808 & ~n51899;
  assign n51901 = n50802 & n50818;
  assign n51902 = ~n51900 & ~n51901;
  assign n51903 = n51896 & n51902;
  assign n51904 = n51895 & n51903;
  assign n51905 = ~n50783 & ~n51904;
  assign n51906 = ~n50854 & ~n51684;
  assign n51907 = ~n50808 & ~n51906;
  assign n51908 = ~n51905 & ~n51907;
  assign n51909 = n51890 & n51908;
  assign n51910 = pi1397 & n51909;
  assign n51911 = ~pi1397 & ~n51909;
  assign po1485 = n51910 | n51911;
  assign n51913 = pi4396 & pi9040;
  assign n51914 = pi4399 & ~pi9040;
  assign n51915 = ~n51913 & ~n51914;
  assign n51916 = ~pi1351 & n51915;
  assign n51917 = pi1351 & ~n51915;
  assign n51918 = ~n51916 & ~n51917;
  assign n51919 = pi4494 & pi9040;
  assign n51920 = pi4583 & ~pi9040;
  assign n51921 = ~n51919 & ~n51920;
  assign n51922 = ~pi1343 & ~n51921;
  assign n51923 = pi1343 & n51921;
  assign n51924 = ~n51922 & ~n51923;
  assign n51925 = pi4392 & pi9040;
  assign n51926 = pi4481 & ~pi9040;
  assign n51927 = ~n51925 & ~n51926;
  assign n51928 = ~pi1364 & n51927;
  assign n51929 = pi1364 & ~n51927;
  assign n51930 = ~n51928 & ~n51929;
  assign n51931 = pi4385 & ~pi9040;
  assign n51932 = pi4399 & pi9040;
  assign n51933 = ~n51931 & ~n51932;
  assign n51934 = ~pi1357 & n51933;
  assign n51935 = pi1357 & ~n51933;
  assign n51936 = ~n51934 & ~n51935;
  assign n51937 = pi4392 & ~pi9040;
  assign n51938 = pi4419 & pi9040;
  assign n51939 = ~n51937 & ~n51938;
  assign n51940 = ~pi1369 & ~n51939;
  assign n51941 = pi1369 & n51939;
  assign n51942 = ~n51940 & ~n51941;
  assign n51943 = n51936 & n51942;
  assign n51944 = ~n51930 & n51943;
  assign n51945 = n51924 & n51944;
  assign n51946 = n51918 & n51945;
  assign n51947 = n51918 & n51930;
  assign n51948 = ~n51942 & n51947;
  assign n51949 = ~n51936 & n51948;
  assign n51950 = n51924 & n51949;
  assign n51951 = ~n51946 & ~n51950;
  assign n51952 = n51930 & n51943;
  assign n51953 = n51918 & ~n51924;
  assign n51954 = n51952 & n51953;
  assign n51955 = ~n51949 & ~n51954;
  assign n51956 = ~n51930 & ~n51936;
  assign n51957 = ~n51918 & n51956;
  assign n51958 = ~n51918 & n51943;
  assign n51959 = ~n51957 & ~n51958;
  assign n51960 = n51924 & ~n51959;
  assign n51961 = ~n51936 & n51942;
  assign n51962 = n51936 & ~n51942;
  assign n51963 = ~n51961 & ~n51962;
  assign n51964 = ~n51924 & ~n51947;
  assign n51965 = ~n51963 & n51964;
  assign n51966 = n51918 & ~n51943;
  assign n51967 = n51924 & n51966;
  assign n51968 = n51930 & n51967;
  assign n51969 = ~n51965 & ~n51968;
  assign n51970 = ~n51960 & n51969;
  assign n51971 = n51955 & n51970;
  assign n51972 = pi4609 & ~pi9040;
  assign n51973 = pi4508 & pi9040;
  assign n51974 = ~n51972 & ~n51973;
  assign n51975 = ~pi1352 & ~n51974;
  assign n51976 = pi1352 & n51974;
  assign n51977 = ~n51975 & ~n51976;
  assign n51978 = ~n51971 & n51977;
  assign n51979 = n51951 & ~n51978;
  assign n51980 = ~n51930 & n51961;
  assign n51981 = ~n51924 & n51980;
  assign n51982 = ~n51918 & n51981;
  assign n51983 = ~n51924 & ~n51977;
  assign n51984 = ~n51936 & ~n51942;
  assign n51985 = ~n51930 & n51984;
  assign n51986 = ~n51958 & ~n51985;
  assign n51987 = n51947 & ~n51963;
  assign n51988 = n51986 & ~n51987;
  assign n51989 = n51983 & ~n51988;
  assign n51990 = n51930 & n51984;
  assign n51991 = ~n51918 & n51990;
  assign n51992 = ~n51918 & ~n51936;
  assign n51993 = n51930 & n51992;
  assign n51994 = ~n51918 & n51962;
  assign n51995 = ~n51993 & ~n51994;
  assign n51996 = n51918 & n51943;
  assign n51997 = ~n51930 & n51962;
  assign n51998 = ~n51996 & ~n51997;
  assign n51999 = n51995 & n51998;
  assign n52000 = n51924 & ~n51999;
  assign n52001 = ~n51991 & ~n52000;
  assign n52002 = ~n51977 & ~n52001;
  assign n52003 = ~n51989 & ~n52002;
  assign n52004 = ~n51982 & n52003;
  assign n52005 = n51979 & n52004;
  assign n52006 = pi1398 & ~n52005;
  assign n52007 = ~pi1398 & n51979;
  assign n52008 = n52004 & n52007;
  assign po1486 = n52006 | n52008;
  assign n52010 = ~n51039 & ~n51797;
  assign n52011 = n51045 & n51067;
  assign n52012 = ~n52010 & ~n52011;
  assign n52013 = n51045 & ~n51051;
  assign n52014 = ~n51074 & ~n52013;
  assign n52015 = ~n51390 & n52014;
  assign n52016 = n51039 & ~n52015;
  assign n52017 = n52012 & ~n52016;
  assign n52018 = ~n51033 & ~n52017;
  assign n52019 = ~n51039 & n51076;
  assign n52020 = ~n51115 & ~n52019;
  assign n52021 = ~n51119 & n52020;
  assign n52022 = ~n51118 & ~n51122;
  assign n52023 = n51039 & n51094;
  assign n52024 = n51045 & n51078;
  assign n52025 = ~n51039 & n51074;
  assign n52026 = ~n52024 & ~n52025;
  assign n52027 = ~n51412 & n52026;
  assign n52028 = ~n52023 & n52027;
  assign n52029 = n52022 & n52028;
  assign n52030 = ~n51105 & n52029;
  assign n52031 = n51033 & ~n52030;
  assign n52032 = n52021 & ~n52031;
  assign n52033 = ~n52018 & n52032;
  assign n52034 = ~pi1392 & ~n52033;
  assign n52035 = pi1392 & n52021;
  assign n52036 = ~n52018 & n52035;
  assign n52037 = ~n52031 & n52036;
  assign po1487 = n52034 | n52037;
  assign n52039 = ~n51248 & n51602;
  assign n52040 = ~n51298 & ~n51306;
  assign n52041 = n51248 & n51267;
  assign n52042 = ~n51248 & n51319;
  assign n52043 = ~n52041 & ~n52042;
  assign n52044 = n52040 & n52043;
  assign n52045 = n51275 & ~n52044;
  assign n52046 = n51248 & n51276;
  assign n52047 = ~n51289 & ~n52046;
  assign n52048 = ~n51300 & n52047;
  assign n52049 = ~n51275 & ~n52048;
  assign n52050 = n51248 & ~n51260;
  assign n52051 = n51266 & n52050;
  assign n52052 = n51254 & n52051;
  assign n52053 = ~n52049 & ~n52052;
  assign n52054 = ~n52045 & n52053;
  assign n52055 = ~n52039 & n52054;
  assign n52056 = ~n51242 & ~n52055;
  assign n52057 = n51248 & n51275;
  assign n52058 = n51277 & n52057;
  assign n52059 = n51275 & n51300;
  assign n52060 = n51275 & n51619;
  assign n52061 = ~n52059 & ~n52060;
  assign n52062 = ~n51248 & ~n52061;
  assign n52063 = ~n52058 & ~n52062;
  assign n52064 = n51248 & n51297;
  assign n52065 = ~n51248 & n51276;
  assign n52066 = ~n52064 & ~n52065;
  assign n52067 = ~n51268 & n52066;
  assign n52068 = ~n51298 & n52067;
  assign n52069 = ~n51275 & ~n52068;
  assign n52070 = ~n51248 & n51290;
  assign n52071 = ~n52069 & ~n52070;
  assign n52072 = ~n51248 & n51268;
  assign n52073 = ~n51614 & ~n52072;
  assign n52074 = n52071 & n52073;
  assign n52075 = n52063 & n52074;
  assign n52076 = n51242 & ~n52075;
  assign n52077 = n51275 & ~n51605;
  assign n52078 = ~n52076 & ~n52077;
  assign n52079 = ~n51301 & ~n52072;
  assign n52080 = ~n51275 & ~n52079;
  assign n52081 = n52078 & ~n52080;
  assign n52082 = ~n52056 & n52081;
  assign n52083 = pi1391 & ~n52082;
  assign n52084 = ~pi1391 & n52082;
  assign po1488 = n52083 | n52084;
  assign n52086 = ~n50939 & n51005;
  assign n52087 = ~n50939 & n50950;
  assign n52088 = ~n52086 & ~n52087;
  assign n52089 = ~n50931 & ~n52088;
  assign n52090 = n50977 & n50991;
  assign n52091 = ~n52089 & ~n52090;
  assign n52092 = ~n51021 & n52091;
  assign n52093 = n50939 & n50956;
  assign n52094 = ~n50950 & ~n52093;
  assign n52095 = n50925 & n50959;
  assign n52096 = n52094 & ~n52095;
  assign n52097 = ~n50931 & ~n52096;
  assign n52098 = n50973 & n52097;
  assign n52099 = n50925 & n50949;
  assign n52100 = n50931 & n52099;
  assign n52101 = ~n50988 & ~n51013;
  assign n52102 = ~n51007 & n52101;
  assign n52103 = ~n52100 & n52102;
  assign n52104 = n50973 & ~n52103;
  assign n52105 = n50925 & n50931;
  assign n52106 = ~n50954 & n52105;
  assign n52107 = ~n50919 & n52106;
  assign n52108 = ~n50939 & n52107;
  assign n52109 = n50925 & n50939;
  assign n52110 = ~n50948 & n52109;
  assign n52111 = n50939 & n50964;
  assign n52112 = ~n52107 & ~n52111;
  assign n52113 = ~n52110 & n52112;
  assign n52114 = n50948 & n51011;
  assign n52115 = n50939 & n51000;
  assign n52116 = ~n50990 & ~n52115;
  assign n52117 = ~n50931 & ~n52116;
  assign n52118 = ~n52114 & ~n52117;
  assign n52119 = n52113 & n52118;
  assign n52120 = ~n50973 & ~n52119;
  assign n52121 = ~n52108 & ~n52120;
  assign n52122 = ~n52104 & n52121;
  assign n52123 = ~n52098 & n52122;
  assign n52124 = n52092 & n52123;
  assign n52125 = pi1396 & ~n52124;
  assign n52126 = ~pi1396 & n52092;
  assign n52127 = n52123 & n52126;
  assign po1489 = n52125 | n52127;
  assign n52129 = n51918 & ~n51930;
  assign n52130 = n51942 & n52129;
  assign n52131 = ~n51980 & ~n51990;
  assign n52132 = ~n52130 & n52131;
  assign n52133 = ~n51924 & n51977;
  assign n52134 = ~n52132 & n52133;
  assign n52135 = ~n51918 & n51977;
  assign n52136 = n51997 & n52135;
  assign n52137 = n51924 & n51985;
  assign n52138 = n51930 & n51942;
  assign n52139 = ~n51958 & ~n52138;
  assign n52140 = n51924 & ~n52139;
  assign n52141 = ~n52137 & ~n52140;
  assign n52142 = n51977 & ~n52141;
  assign n52143 = ~n52136 & ~n52142;
  assign n52144 = ~n51918 & n51930;
  assign n52145 = n51942 & n52144;
  assign n52146 = n51936 & n51948;
  assign n52147 = ~n52145 & ~n52146;
  assign n52148 = n51924 & ~n52147;
  assign n52149 = n52143 & ~n52148;
  assign n52150 = ~n51918 & ~n51924;
  assign n52151 = n51943 & n52150;
  assign n52152 = ~n51930 & n52151;
  assign n52153 = ~n51963 & n52129;
  assign n52154 = ~n51949 & ~n52153;
  assign n52155 = ~n51963 & n52144;
  assign n52156 = ~n51918 & ~n51930;
  assign n52157 = ~n51942 & n52156;
  assign n52158 = ~n51936 & n52157;
  assign n52159 = ~n52155 & ~n52158;
  assign n52160 = ~n51954 & n52159;
  assign n52161 = n52154 & n52160;
  assign n52162 = ~n52152 & n52161;
  assign n52163 = n51918 & n51924;
  assign n52164 = ~n51930 & n52163;
  assign n52165 = n51936 & n52164;
  assign n52166 = n52162 & ~n52165;
  assign n52167 = ~n51977 & ~n52166;
  assign n52168 = n52149 & ~n52167;
  assign n52169 = ~n52134 & n52168;
  assign n52170 = ~pi1408 & ~n52169;
  assign n52171 = pi1408 & n52149;
  assign n52172 = ~n52134 & n52171;
  assign n52173 = ~n52167 & n52172;
  assign po1490 = n52170 | n52173;
  assign n52175 = ~n51994 & ~n51996;
  assign n52176 = n51924 & ~n52175;
  assign n52177 = ~n51950 & ~n52176;
  assign n52178 = n51977 & ~n52177;
  assign n52179 = ~n51918 & n51952;
  assign n52180 = ~n51942 & n52129;
  assign n52181 = n51930 & ~n51936;
  assign n52182 = ~n51961 & ~n52181;
  assign n52183 = ~n51918 & ~n52182;
  assign n52184 = ~n52180 & ~n52183;
  assign n52185 = n51924 & ~n52184;
  assign n52186 = ~n52179 & ~n52185;
  assign n52187 = n51918 & ~n52182;
  assign n52188 = ~n51944 & ~n52187;
  assign n52189 = ~n51924 & ~n52188;
  assign n52190 = ~n51987 & ~n52189;
  assign n52191 = n52186 & n52190;
  assign n52192 = ~n51977 & ~n52191;
  assign n52193 = ~n51961 & n52156;
  assign n52194 = n51977 & n52193;
  assign n52195 = n51961 & n52144;
  assign n52196 = n51924 & n52195;
  assign n52197 = ~n51930 & n52150;
  assign n52198 = ~n51942 & n52197;
  assign n52199 = ~n52196 & ~n52198;
  assign n52200 = ~n52194 & n52199;
  assign n52201 = ~n51992 & ~n51997;
  assign n52202 = n52133 & ~n52201;
  assign n52203 = n52200 & ~n52202;
  assign n52204 = ~n52192 & n52203;
  assign n52205 = ~n52178 & n52204;
  assign n52206 = pi1399 & ~n52205;
  assign n52207 = ~pi1399 & n52205;
  assign po1491 = n52206 | n52207;
  assign n52209 = n50939 & n52095;
  assign n52210 = ~n50939 & n52099;
  assign n52211 = ~n52209 & ~n52210;
  assign n52212 = n50931 & ~n52211;
  assign n52213 = ~n50919 & n50925;
  assign n52214 = ~n51013 & ~n52213;
  assign n52215 = ~n50940 & n52214;
  assign n52216 = n50931 & ~n52215;
  assign n52217 = n50919 & n50977;
  assign n52218 = ~n52086 & ~n52110;
  assign n52219 = ~n50919 & ~n50925;
  assign n52220 = ~n50931 & ~n50939;
  assign n52221 = n52219 & n52220;
  assign n52222 = n52218 & ~n52221;
  assign n52223 = ~n52217 & n52222;
  assign n52224 = ~n52216 & n52223;
  assign n52225 = n50973 & ~n52224;
  assign n52226 = ~n52212 & ~n52225;
  assign n52227 = n50939 & n51005;
  assign n52228 = ~n50956 & ~n50991;
  assign n52229 = n50931 & ~n52228;
  assign n52230 = ~n52227 & ~n52229;
  assign n52231 = ~n50994 & n52230;
  assign n52232 = ~n50973 & ~n52231;
  assign n52233 = ~n50959 & ~n51000;
  assign n52234 = ~n50925 & ~n52233;
  assign n52235 = ~n50981 & ~n52234;
  assign n52236 = ~n50931 & ~n52235;
  assign n52237 = ~n50973 & n52236;
  assign n52238 = ~n52232 & ~n52237;
  assign n52239 = n52226 & n52238;
  assign n52240 = pi1389 & ~n52239;
  assign n52241 = ~pi1389 & n52226;
  assign n52242 = n52238 & n52241;
  assign po1492 = n52240 | n52242;
  assign n52244 = ~n51539 & n51581;
  assign n52245 = ~n51567 & ~n52244;
  assign n52246 = ~n51548 & ~n52245;
  assign n52247 = n51521 & n51540;
  assign n52248 = ~n51521 & ~n51539;
  assign n52249 = n51527 & n52248;
  assign n52250 = ~n52247 & ~n52249;
  assign n52251 = n51548 & ~n52250;
  assign n52252 = ~n51521 & n51557;
  assign n52253 = ~n51747 & ~n52252;
  assign n52254 = ~n51584 & n52253;
  assign n52255 = ~n52251 & n52254;
  assign n52256 = ~n52246 & n52255;
  assign n52257 = ~n51728 & ~n51739;
  assign n52258 = n52256 & n52257;
  assign n52259 = n51515 & ~n52258;
  assign n52260 = n51533 & n51581;
  assign n52261 = n51521 & n51553;
  assign n52262 = ~n52260 & ~n52261;
  assign n52263 = n51548 & ~n52262;
  assign n52264 = n51540 & n51548;
  assign n52265 = ~n51521 & n52264;
  assign n52266 = ~n52263 & ~n52265;
  assign n52267 = n51551 & n51726;
  assign n52268 = n51588 & ~n52267;
  assign n52269 = n51548 & ~n52268;
  assign n52270 = ~n51521 & n51564;
  assign n52271 = ~n52269 & ~n52270;
  assign n52272 = n52266 & n52271;
  assign n52273 = ~n51515 & ~n52272;
  assign n52274 = ~n51542 & ~n51557;
  assign n52275 = ~n51733 & n52274;
  assign n52276 = n51578 & ~n52275;
  assign n52277 = ~n52273 & ~n52276;
  assign n52278 = ~n51584 & ~n51728;
  assign n52279 = ~n51548 & ~n52278;
  assign n52280 = n52277 & ~n52279;
  assign n52281 = ~n52259 & n52280;
  assign n52282 = ~pi1401 & n52281;
  assign n52283 = pi1401 & ~n52281;
  assign po1493 = n52282 | n52283;
  assign n52285 = ~n51606 & ~n52072;
  assign n52286 = ~n52052 & n52285;
  assign n52287 = n51275 & ~n52286;
  assign n52288 = ~n51614 & ~n52060;
  assign n52289 = ~n51602 & ~n52065;
  assign n52290 = ~n51275 & ~n52289;
  assign n52291 = ~n51306 & ~n52290;
  assign n52292 = n52288 & n52291;
  assign n52293 = n51242 & ~n52292;
  assign n52294 = ~n51260 & n51266;
  assign n52295 = ~n51278 & ~n52294;
  assign n52296 = n51248 & ~n52295;
  assign n52297 = ~n51268 & ~n51621;
  assign n52298 = ~n51275 & ~n52297;
  assign n52299 = n51248 & n51266;
  assign n52300 = ~n51290 & ~n52299;
  assign n52301 = ~n51281 & n52300;
  assign n52302 = n51275 & ~n52301;
  assign n52303 = ~n52298 & ~n52302;
  assign n52304 = ~n52296 & n52303;
  assign n52305 = ~n51242 & ~n52304;
  assign n52306 = ~n52293 & ~n52305;
  assign n52307 = ~n51617 & ~n51634;
  assign n52308 = n52306 & n52307;
  assign n52309 = ~n52287 & n52308;
  assign n52310 = ~pi1407 & ~n52309;
  assign n52311 = pi1407 & n52307;
  assign n52312 = ~n52287 & n52311;
  assign n52313 = n52306 & n52312;
  assign po1494 = n52310 | n52313;
  assign n52315 = ~n50955 & ~n52099;
  assign n52316 = n51001 & ~n52315;
  assign n52317 = ~n50950 & ~n50976;
  assign n52318 = ~n50991 & ~n52095;
  assign n52319 = n52317 & n52318;
  assign n52320 = n50939 & ~n52319;
  assign n52321 = ~n52316 & ~n52320;
  assign n52322 = ~n52086 & n52321;
  assign n52323 = n50973 & ~n52322;
  assign n52324 = ~n50939 & n50991;
  assign n52325 = n50939 & n52099;
  assign n52326 = ~n52324 & ~n52325;
  assign n52327 = ~n50931 & ~n52326;
  assign n52328 = n50939 & ~n52233;
  assign n52329 = ~n50925 & n52328;
  assign n52330 = ~n50931 & ~n52315;
  assign n52331 = n50948 & n52109;
  assign n52332 = ~n50961 & ~n52331;
  assign n52333 = ~n52095 & n52332;
  assign n52334 = n50931 & ~n52333;
  assign n52335 = ~n52330 & ~n52334;
  assign n52336 = ~n52329 & n52335;
  assign n52337 = ~n52324 & n52336;
  assign n52338 = ~n50973 & ~n52337;
  assign n52339 = ~n52327 & ~n52338;
  assign n52340 = ~n52323 & n52339;
  assign n52341 = ~pi1388 & ~n52340;
  assign n52342 = pi1388 & ~n52327;
  assign n52343 = ~n52323 & n52342;
  assign n52344 = ~n52338 & n52343;
  assign po1495 = n52341 | n52344;
  assign n52346 = n51930 & n51961;
  assign n52347 = ~n51944 & ~n52346;
  assign n52348 = n51924 & ~n52347;
  assign n52349 = n51918 & n51962;
  assign n52350 = ~n51980 & ~n52349;
  assign n52351 = ~n51952 & n52350;
  assign n52352 = ~n51924 & ~n52351;
  assign n52353 = ~n52348 & ~n52352;
  assign n52354 = ~n51977 & ~n52146;
  assign n52355 = n52353 & n52354;
  assign n52356 = ~n52137 & n52355;
  assign n52357 = ~n51918 & n51944;
  assign n52358 = n51918 & n51984;
  assign n52359 = ~n51994 & ~n52358;
  assign n52360 = ~n51924 & ~n52359;
  assign n52361 = ~n52357 & ~n52360;
  assign n52362 = n51924 & n51997;
  assign n52363 = n52131 & ~n52362;
  assign n52364 = ~n51952 & n52363;
  assign n52365 = n51918 & ~n52364;
  assign n52366 = n52361 & ~n52365;
  assign n52367 = n51977 & n52366;
  assign n52368 = ~n52356 & ~n52367;
  assign n52369 = n51930 & n51994;
  assign n52370 = ~n52158 & ~n52369;
  assign n52371 = n51924 & ~n52370;
  assign n52372 = ~n51924 & n52181;
  assign n52373 = ~n51918 & n52372;
  assign n52374 = ~n52371 & ~n52373;
  assign n52375 = ~n52368 & n52374;
  assign n52376 = ~pi1409 & ~n52375;
  assign n52377 = pi1409 & ~n52371;
  assign n52378 = ~n52368 & n52377;
  assign n52379 = ~n52373 & n52378;
  assign po1496 = n52376 | n52379;
  assign n52381 = ~n51521 & n51553;
  assign n52382 = ~n51552 & ~n52381;
  assign n52383 = ~n51548 & ~n52382;
  assign n52384 = n51548 & ~n51744;
  assign n52385 = ~n52383 & ~n52384;
  assign n52386 = ~n51760 & n52385;
  assign n52387 = n51515 & ~n52386;
  assign n52388 = ~n51548 & n51564;
  assign n52389 = ~n52387 & ~n52388;
  assign n52390 = ~n52252 & ~n52261;
  assign n52391 = n51548 & ~n52390;
  assign n52392 = n51548 & n51554;
  assign n52393 = n51521 & n51567;
  assign n52394 = ~n52392 & ~n52393;
  assign n52395 = ~n51527 & n51719;
  assign n52396 = ~n51731 & ~n52395;
  assign n52397 = ~n51533 & ~n52396;
  assign n52398 = ~n51584 & ~n52397;
  assign n52399 = ~n52249 & n52398;
  assign n52400 = n52394 & n52399;
  assign n52401 = ~n51515 & ~n52400;
  assign n52402 = ~n52391 & ~n52401;
  assign n52403 = n52389 & n52402;
  assign n52404 = pi1437 & n52403;
  assign n52405 = ~pi1437 & ~n52403;
  assign po1497 = n52404 | n52405;
  assign n52407 = pi4604 & ~pi9040;
  assign n52408 = pi4937 & pi9040;
  assign n52409 = ~n52407 & ~n52408;
  assign n52410 = ~pi1423 & ~n52409;
  assign n52411 = pi1423 & n52409;
  assign n52412 = ~n52410 & ~n52411;
  assign n52413 = pi4710 & ~pi9040;
  assign n52414 = pi4754 & pi9040;
  assign n52415 = ~n52413 & ~n52414;
  assign n52416 = ~pi1427 & n52415;
  assign n52417 = pi1427 & ~n52415;
  assign n52418 = ~n52416 & ~n52417;
  assign n52419 = pi4689 & pi9040;
  assign n52420 = pi4590 & ~pi9040;
  assign n52421 = ~n52419 & ~n52420;
  assign n52422 = pi1404 & n52421;
  assign n52423 = ~pi1404 & ~n52421;
  assign n52424 = ~n52422 & ~n52423;
  assign n52425 = n52418 & n52424;
  assign n52426 = pi4715 & ~pi9040;
  assign n52427 = pi4695 & pi9040;
  assign n52428 = ~n52426 & ~n52427;
  assign n52429 = pi1414 & n52428;
  assign n52430 = ~pi1414 & ~n52428;
  assign n52431 = ~n52429 & ~n52430;
  assign n52432 = pi4616 & ~pi9040;
  assign n52433 = pi4958 & pi9040;
  assign n52434 = ~n52432 & ~n52433;
  assign n52435 = pi1438 & n52434;
  assign n52436 = ~pi1438 & ~n52434;
  assign n52437 = ~n52435 & ~n52436;
  assign n52438 = ~n52431 & ~n52437;
  assign n52439 = n52425 & n52438;
  assign n52440 = pi4604 & pi9040;
  assign n52441 = pi4816 & ~pi9040;
  assign n52442 = ~n52440 & ~n52441;
  assign n52443 = ~pi1406 & n52442;
  assign n52444 = pi1406 & ~n52442;
  assign n52445 = ~n52443 & ~n52444;
  assign n52446 = ~n52418 & ~n52424;
  assign n52447 = ~n52445 & n52446;
  assign n52448 = n52431 & n52445;
  assign n52449 = ~n52424 & n52448;
  assign n52450 = n52418 & n52449;
  assign n52451 = ~n52447 & ~n52450;
  assign n52452 = ~n52418 & n52424;
  assign n52453 = n52431 & n52452;
  assign n52454 = n52451 & ~n52453;
  assign n52455 = ~n52437 & ~n52454;
  assign n52456 = ~n52418 & n52445;
  assign n52457 = ~n52431 & n52437;
  assign n52458 = n52456 & n52457;
  assign n52459 = n52445 & n52446;
  assign n52460 = ~n52431 & n52459;
  assign n52461 = ~n52458 & ~n52460;
  assign n52462 = ~n52455 & n52461;
  assign n52463 = ~n52439 & n52462;
  assign n52464 = n52425 & ~n52445;
  assign n52465 = ~n52431 & n52464;
  assign n52466 = ~n52445 & n52452;
  assign n52467 = n52431 & n52466;
  assign n52468 = ~n52465 & ~n52467;
  assign n52469 = n52463 & n52468;
  assign n52470 = ~n52412 & ~n52469;
  assign n52471 = ~n52418 & ~n52431;
  assign n52472 = n52445 & n52471;
  assign n52473 = n52424 & n52472;
  assign n52474 = ~n52464 & ~n52473;
  assign n52475 = ~n52437 & ~n52474;
  assign n52476 = n52425 & n52448;
  assign n52477 = ~n52431 & n52445;
  assign n52478 = ~n52424 & n52477;
  assign n52479 = n52418 & n52478;
  assign n52480 = ~n52476 & ~n52479;
  assign n52481 = ~n52418 & n52448;
  assign n52482 = ~n52431 & n52466;
  assign n52483 = ~n52481 & ~n52482;
  assign n52484 = n52437 & ~n52483;
  assign n52485 = n52480 & ~n52484;
  assign n52486 = ~n52475 & n52485;
  assign n52487 = n52412 & ~n52486;
  assign n52488 = ~n52418 & ~n52445;
  assign n52489 = n52431 & n52488;
  assign n52490 = n52418 & ~n52445;
  assign n52491 = ~n52431 & n52490;
  assign n52492 = ~n52489 & ~n52491;
  assign n52493 = ~n52437 & ~n52492;
  assign n52494 = n52418 & ~n52424;
  assign n52495 = ~n52445 & n52494;
  assign n52496 = n52431 & n52495;
  assign n52497 = ~n52476 & ~n52496;
  assign n52498 = ~n52459 & n52497;
  assign n52499 = n52437 & ~n52498;
  assign n52500 = ~n52493 & ~n52499;
  assign n52501 = ~n52424 & n52445;
  assign n52502 = n52437 & n52501;
  assign n52503 = ~n52431 & n52502;
  assign n52504 = n52500 & ~n52503;
  assign n52505 = ~n52487 & n52504;
  assign n52506 = ~n52470 & n52505;
  assign n52507 = ~pi1442 & ~n52506;
  assign n52508 = pi1442 & n52506;
  assign po1520 = n52507 | n52508;
  assign n52510 = pi4617 & pi9040;
  assign n52511 = pi4850 & ~pi9040;
  assign n52512 = ~n52510 & ~n52511;
  assign n52513 = ~pi1433 & ~n52512;
  assign n52514 = pi1433 & n52512;
  assign n52515 = ~n52513 & ~n52514;
  assign n52516 = pi4623 & ~pi9040;
  assign n52517 = pi4772 & pi9040;
  assign n52518 = ~n52516 & ~n52517;
  assign n52519 = ~pi1431 & ~n52518;
  assign n52520 = pi1431 & n52518;
  assign n52521 = ~n52519 & ~n52520;
  assign n52522 = pi4738 & pi9040;
  assign n52523 = pi4817 & ~pi9040;
  assign n52524 = ~n52522 & ~n52523;
  assign n52525 = ~pi1434 & n52524;
  assign n52526 = pi1434 & ~n52524;
  assign n52527 = ~n52525 & ~n52526;
  assign n52528 = n52521 & n52527;
  assign n52529 = n52515 & n52528;
  assign n52530 = pi4817 & pi9040;
  assign n52531 = pi4618 & ~pi9040;
  assign n52532 = ~n52530 & ~n52531;
  assign n52533 = ~pi1419 & n52532;
  assign n52534 = pi1419 & ~n52532;
  assign n52535 = ~n52533 & ~n52534;
  assign n52536 = ~n52515 & ~n52535;
  assign n52537 = ~n52521 & n52536;
  assign n52538 = ~n52529 & ~n52537;
  assign n52539 = pi4737 & ~pi9040;
  assign n52540 = pi4815 & pi9040;
  assign n52541 = ~n52539 & ~n52540;
  assign n52542 = ~pi1413 & ~n52541;
  assign n52543 = pi1413 & n52541;
  assign n52544 = ~n52542 & ~n52543;
  assign n52545 = ~n52515 & n52544;
  assign n52546 = ~n52521 & n52545;
  assign n52547 = n52538 & ~n52546;
  assign n52548 = ~n52521 & ~n52544;
  assign n52549 = n52515 & n52548;
  assign n52550 = n52535 & n52549;
  assign n52551 = n52547 & ~n52550;
  assign n52552 = ~n52515 & ~n52544;
  assign n52553 = ~n52535 & n52552;
  assign n52554 = ~n52521 & n52544;
  assign n52555 = ~n52553 & ~n52554;
  assign n52556 = ~n52527 & ~n52555;
  assign n52557 = ~n52527 & n52545;
  assign n52558 = n52535 & n52557;
  assign n52559 = ~n52556 & ~n52558;
  assign n52560 = n52551 & n52559;
  assign n52561 = pi4850 & pi9040;
  assign n52562 = pi4619 & ~pi9040;
  assign n52563 = ~n52561 & ~n52562;
  assign n52564 = ~pi1412 & ~n52563;
  assign n52565 = pi1412 & n52563;
  assign n52566 = ~n52564 & ~n52565;
  assign n52567 = ~n52560 & n52566;
  assign n52568 = n52527 & ~n52535;
  assign n52569 = n52549 & n52568;
  assign n52570 = n52521 & n52535;
  assign n52571 = ~n52515 & n52570;
  assign n52572 = n52535 & n52552;
  assign n52573 = ~n52571 & ~n52572;
  assign n52574 = n52527 & ~n52573;
  assign n52575 = ~n52569 & ~n52574;
  assign n52576 = ~n52566 & ~n52575;
  assign n52577 = ~n52527 & ~n52535;
  assign n52578 = n52545 & n52577;
  assign n52579 = n52521 & n52578;
  assign n52580 = n52515 & n52544;
  assign n52581 = ~n52527 & n52535;
  assign n52582 = n52580 & n52581;
  assign n52583 = ~n52544 & n52570;
  assign n52584 = ~n52515 & n52583;
  assign n52585 = n52515 & ~n52544;
  assign n52586 = n52521 & n52585;
  assign n52587 = ~n52527 & n52586;
  assign n52588 = ~n52535 & n52587;
  assign n52589 = ~n52584 & ~n52588;
  assign n52590 = ~n52582 & n52589;
  assign n52591 = ~n52579 & n52590;
  assign n52592 = ~n52521 & n52535;
  assign n52593 = n52544 & n52592;
  assign n52594 = n52515 & n52593;
  assign n52595 = n52591 & ~n52594;
  assign n52596 = ~n52566 & ~n52595;
  assign n52597 = n52515 & n52521;
  assign n52598 = n52544 & n52597;
  assign n52599 = ~n52535 & n52598;
  assign n52600 = ~n52583 & ~n52599;
  assign n52601 = ~n52535 & n52546;
  assign n52602 = n52600 & ~n52601;
  assign n52603 = n52527 & ~n52602;
  assign n52604 = ~n52521 & ~n52535;
  assign n52605 = ~n52527 & n52604;
  assign n52606 = n52552 & n52605;
  assign n52607 = ~n52603 & ~n52606;
  assign n52608 = ~n52596 & n52607;
  assign n52609 = ~n52576 & n52608;
  assign n52610 = ~n52567 & n52609;
  assign n52611 = n52515 & ~n52521;
  assign n52612 = n52581 & n52611;
  assign n52613 = n52610 & ~n52612;
  assign n52614 = ~pi1441 & ~n52613;
  assign n52615 = pi1441 & ~n52612;
  assign n52616 = n52609 & n52615;
  assign n52617 = ~n52567 & n52616;
  assign po1521 = n52614 | n52617;
  assign n52619 = pi4709 & ~pi9040;
  assign n52620 = pi4816 & pi9040;
  assign n52621 = ~n52619 & ~n52620;
  assign n52622 = ~pi1410 & ~n52621;
  assign n52623 = pi1410 & n52621;
  assign n52624 = ~n52622 & ~n52623;
  assign n52625 = pi4774 & pi9040;
  assign n52626 = pi4959 & ~pi9040;
  assign n52627 = ~n52625 & ~n52626;
  assign n52628 = ~pi1404 & n52627;
  assign n52629 = pi1404 & ~n52627;
  assign n52630 = ~n52628 & ~n52629;
  assign n52631 = pi4831 & pi9040;
  assign n52632 = pi4608 & ~pi9040;
  assign n52633 = ~n52631 & ~n52632;
  assign n52634 = ~pi1431 & n52633;
  assign n52635 = pi1431 & ~n52633;
  assign n52636 = ~n52634 & ~n52635;
  assign n52637 = pi4612 & ~pi9040;
  assign n52638 = pi4692 & pi9040;
  assign n52639 = ~n52637 & ~n52638;
  assign n52640 = ~pi1423 & n52639;
  assign n52641 = pi1423 & ~n52639;
  assign n52642 = ~n52640 & ~n52641;
  assign n52643 = ~n52636 & ~n52642;
  assign n52644 = n52630 & n52643;
  assign n52645 = pi4736 & ~pi9040;
  assign n52646 = pi4654 & pi9040;
  assign n52647 = ~n52645 & ~n52646;
  assign n52648 = pi1428 & n52647;
  assign n52649 = ~pi1428 & ~n52647;
  assign n52650 = ~n52648 & ~n52649;
  assign n52651 = n52644 & ~n52650;
  assign n52652 = n52636 & n52642;
  assign n52653 = n52630 & n52652;
  assign n52654 = ~n52650 & n52653;
  assign n52655 = ~n52651 & ~n52654;
  assign n52656 = ~n52630 & n52652;
  assign n52657 = n52650 & n52656;
  assign n52658 = ~n52636 & n52642;
  assign n52659 = n52630 & n52658;
  assign n52660 = n52650 & n52659;
  assign n52661 = ~n52657 & ~n52660;
  assign n52662 = n52655 & n52661;
  assign n52663 = n52624 & ~n52662;
  assign n52664 = n52630 & n52650;
  assign n52665 = ~n52642 & n52664;
  assign n52666 = n52636 & n52665;
  assign n52667 = ~n52659 & ~n52666;
  assign n52668 = n52624 & ~n52667;
  assign n52669 = ~n52624 & ~n52642;
  assign n52670 = ~n52650 & n52669;
  assign n52671 = ~n52630 & ~n52636;
  assign n52672 = n52650 & n52652;
  assign n52673 = ~n52671 & ~n52672;
  assign n52674 = ~n52624 & ~n52673;
  assign n52675 = ~n52670 & ~n52674;
  assign n52676 = n52636 & ~n52642;
  assign n52677 = ~n52630 & n52676;
  assign n52678 = ~n52650 & n52677;
  assign n52679 = n52675 & ~n52678;
  assign n52680 = ~n52642 & n52671;
  assign n52681 = n52650 & n52680;
  assign n52682 = n52679 & ~n52681;
  assign n52683 = ~n52668 & n52682;
  assign n52684 = pi4959 & pi9040;
  assign n52685 = pi4754 & ~pi9040;
  assign n52686 = ~n52684 & ~n52685;
  assign n52687 = pi1433 & n52686;
  assign n52688 = ~pi1433 & ~n52686;
  assign n52689 = ~n52687 & ~n52688;
  assign n52690 = ~n52683 & ~n52689;
  assign n52691 = n52630 & ~n52642;
  assign n52692 = ~n52624 & n52650;
  assign n52693 = n52689 & n52692;
  assign n52694 = n52691 & n52693;
  assign n52695 = n52630 & ~n52650;
  assign n52696 = n52642 & n52695;
  assign n52697 = ~n52624 & ~n52696;
  assign n52698 = ~n52630 & n52650;
  assign n52699 = n52636 & n52698;
  assign n52700 = ~n52643 & ~n52691;
  assign n52701 = ~n52650 & ~n52700;
  assign n52702 = n52624 & ~n52656;
  assign n52703 = ~n52701 & n52702;
  assign n52704 = ~n52699 & n52703;
  assign n52705 = ~n52697 & ~n52704;
  assign n52706 = ~n52630 & n52658;
  assign n52707 = n52650 & n52706;
  assign n52708 = ~n52705 & ~n52707;
  assign n52709 = n52689 & ~n52708;
  assign n52710 = ~n52694 & ~n52709;
  assign n52711 = ~n52690 & n52710;
  assign n52712 = ~n52663 & n52711;
  assign n52713 = ~n52624 & n52678;
  assign n52714 = n52712 & ~n52713;
  assign n52715 = pi1443 & ~n52714;
  assign n52716 = ~pi1443 & ~n52713;
  assign n52717 = n52711 & n52716;
  assign n52718 = ~n52663 & n52717;
  assign po1525 = n52715 | n52718;
  assign n52720 = pi4780 & ~pi9040;
  assign n52721 = pi4606 & pi9040;
  assign n52722 = ~n52720 & ~n52721;
  assign n52723 = ~pi1406 & n52722;
  assign n52724 = pi1406 & ~n52722;
  assign n52725 = ~n52723 & ~n52724;
  assign n52726 = pi4590 & pi9040;
  assign n52727 = pi4949 & ~pi9040;
  assign n52728 = ~n52726 & ~n52727;
  assign n52729 = ~pi1432 & ~n52728;
  assign n52730 = pi1432 & n52728;
  assign n52731 = ~n52729 & ~n52730;
  assign n52732 = pi4709 & pi9040;
  assign n52733 = pi4691 & ~pi9040;
  assign n52734 = ~n52732 & ~n52733;
  assign n52735 = ~pi1400 & ~n52734;
  assign n52736 = pi1400 & n52734;
  assign n52737 = ~n52735 & ~n52736;
  assign n52738 = pi4675 & pi9040;
  assign n52739 = pi4831 & ~pi9040;
  assign n52740 = ~n52738 & ~n52739;
  assign n52741 = pi1424 & n52740;
  assign n52742 = ~pi1424 & ~n52740;
  assign n52743 = ~n52741 & ~n52742;
  assign n52744 = ~n52737 & n52743;
  assign n52745 = n52731 & n52744;
  assign n52746 = ~n52725 & n52745;
  assign n52747 = pi4675 & ~pi9040;
  assign n52748 = pi4733 & pi9040;
  assign n52749 = ~n52747 & ~n52748;
  assign n52750 = ~pi1411 & n52749;
  assign n52751 = pi1411 & ~n52749;
  assign n52752 = ~n52750 & ~n52751;
  assign n52753 = n52725 & ~n52752;
  assign n52754 = ~n52731 & n52753;
  assign n52755 = ~n52737 & n52754;
  assign n52756 = ~n52746 & ~n52755;
  assign n52757 = pi4606 & ~pi9040;
  assign n52758 = pi4612 & pi9040;
  assign n52759 = ~n52757 & ~n52758;
  assign n52760 = ~pi1427 & ~n52759;
  assign n52761 = pi1427 & n52759;
  assign n52762 = ~n52760 & ~n52761;
  assign n52763 = ~n52743 & ~n52762;
  assign n52764 = ~n52725 & ~n52752;
  assign n52765 = ~n52737 & n52764;
  assign n52766 = n52731 & n52753;
  assign n52767 = n52737 & n52766;
  assign n52768 = ~n52765 & ~n52767;
  assign n52769 = n52731 & n52752;
  assign n52770 = ~n52737 & n52769;
  assign n52771 = n52768 & ~n52770;
  assign n52772 = n52763 & ~n52771;
  assign n52773 = ~n52731 & ~n52737;
  assign n52774 = n52725 & n52773;
  assign n52775 = n52725 & n52752;
  assign n52776 = n52731 & n52775;
  assign n52777 = n52737 & n52776;
  assign n52778 = ~n52774 & ~n52777;
  assign n52779 = n52731 & n52764;
  assign n52780 = ~n52754 & ~n52779;
  assign n52781 = n52778 & n52780;
  assign n52782 = n52743 & ~n52781;
  assign n52783 = ~n52731 & n52737;
  assign n52784 = ~n52725 & n52783;
  assign n52785 = n52752 & n52784;
  assign n52786 = ~n52782 & ~n52785;
  assign n52787 = ~n52762 & ~n52786;
  assign n52788 = ~n52772 & ~n52787;
  assign n52789 = ~n52731 & n52775;
  assign n52790 = ~n52764 & ~n52775;
  assign n52791 = n52737 & ~n52790;
  assign n52792 = ~n52789 & ~n52791;
  assign n52793 = ~n52743 & ~n52792;
  assign n52794 = ~n52725 & n52752;
  assign n52795 = n52731 & n52794;
  assign n52796 = ~n52770 & ~n52795;
  assign n52797 = ~n52767 & n52796;
  assign n52798 = n52743 & ~n52797;
  assign n52799 = ~n52793 & ~n52798;
  assign n52800 = ~n52737 & ~n52743;
  assign n52801 = n52753 & n52800;
  assign n52802 = n52737 & n52789;
  assign n52803 = ~n52731 & ~n52752;
  assign n52804 = ~n52725 & n52803;
  assign n52805 = n52737 & n52804;
  assign n52806 = ~n52802 & ~n52805;
  assign n52807 = ~n52725 & n52773;
  assign n52808 = n52752 & n52807;
  assign n52809 = n52806 & ~n52808;
  assign n52810 = ~n52801 & n52809;
  assign n52811 = n52799 & n52810;
  assign n52812 = n52762 & ~n52811;
  assign n52813 = n52788 & ~n52812;
  assign n52814 = n52756 & n52813;
  assign n52815 = pi1452 & ~n52814;
  assign n52816 = ~pi1452 & n52756;
  assign n52817 = n52788 & n52816;
  assign n52818 = ~n52812 & n52817;
  assign po1527 = n52815 | n52818;
  assign n52820 = n52737 & n52769;
  assign n52821 = ~n52779 & ~n52820;
  assign n52822 = ~n52755 & n52821;
  assign n52823 = n52743 & ~n52822;
  assign n52824 = ~n52737 & n52804;
  assign n52825 = ~n52737 & n52795;
  assign n52826 = ~n52731 & n52752;
  assign n52827 = ~n52753 & ~n52826;
  assign n52828 = n52737 & ~n52827;
  assign n52829 = ~n52825 & ~n52828;
  assign n52830 = ~n52824 & n52829;
  assign n52831 = ~n52743 & ~n52830;
  assign n52832 = ~n52823 & ~n52831;
  assign n52833 = n52762 & ~n52832;
  assign n52834 = ~n52743 & n52789;
  assign n52835 = ~n52737 & n52834;
  assign n52836 = n52731 & ~n52737;
  assign n52837 = n52753 & n52836;
  assign n52838 = ~n52743 & n52837;
  assign n52839 = ~n52835 & ~n52838;
  assign n52840 = n52743 & n52808;
  assign n52841 = n52839 & ~n52840;
  assign n52842 = n52744 & n52752;
  assign n52843 = ~n52752 & n52836;
  assign n52844 = ~n52820 & ~n52843;
  assign n52845 = ~n52743 & ~n52844;
  assign n52846 = ~n52801 & ~n52845;
  assign n52847 = ~n52805 & ~n52837;
  assign n52848 = n52737 & n52743;
  assign n52849 = n52803 & n52848;
  assign n52850 = ~n52725 & n52826;
  assign n52851 = n52743 & n52850;
  assign n52852 = ~n52849 & ~n52851;
  assign n52853 = n52847 & n52852;
  assign n52854 = n52846 & n52853;
  assign n52855 = ~n52842 & n52854;
  assign n52856 = ~n52762 & ~n52855;
  assign n52857 = ~n52737 & n52776;
  assign n52858 = n52737 & n52764;
  assign n52859 = ~n52857 & ~n52858;
  assign n52860 = n52743 & ~n52859;
  assign n52861 = ~n52856 & ~n52860;
  assign n52862 = n52841 & n52861;
  assign n52863 = ~n52833 & n52862;
  assign n52864 = ~pi1449 & ~n52863;
  assign n52865 = pi1449 & n52863;
  assign po1529 = n52864 | n52865;
  assign n52867 = pi4707 & ~pi9040;
  assign n52868 = pi4610 & pi9040;
  assign n52869 = ~n52867 & ~n52868;
  assign n52870 = ~pi1436 & ~n52869;
  assign n52871 = pi1436 & n52869;
  assign n52872 = ~n52870 & ~n52871;
  assign n52873 = pi4737 & pi9040;
  assign n52874 = pi4947 & ~pi9040;
  assign n52875 = ~n52873 & ~n52874;
  assign n52876 = ~pi1430 & n52875;
  assign n52877 = pi1430 & ~n52875;
  assign n52878 = ~n52876 & ~n52877;
  assign n52879 = pi4617 & ~pi9040;
  assign n52880 = pi4734 & pi9040;
  assign n52881 = ~n52879 & ~n52880;
  assign n52882 = ~pi1421 & n52881;
  assign n52883 = pi1421 & ~n52881;
  assign n52884 = ~n52882 & ~n52883;
  assign n52885 = pi4619 & pi9040;
  assign n52886 = pi4839 & ~pi9040;
  assign n52887 = ~n52885 & ~n52886;
  assign n52888 = ~pi1420 & ~n52887;
  assign n52889 = pi1420 & n52887;
  assign n52890 = ~n52888 & ~n52889;
  assign n52891 = pi4690 & pi9040;
  assign n52892 = pi4772 & ~pi9040;
  assign n52893 = ~n52891 & ~n52892;
  assign n52894 = ~pi1418 & n52893;
  assign n52895 = pi1418 & ~n52893;
  assign n52896 = ~n52894 & ~n52895;
  assign n52897 = n52890 & ~n52896;
  assign n52898 = ~n52884 & n52897;
  assign n52899 = pi4652 & ~pi9040;
  assign n52900 = pi4947 & pi9040;
  assign n52901 = ~n52899 & ~n52900;
  assign n52902 = pi1429 & n52901;
  assign n52903 = ~pi1429 & ~n52901;
  assign n52904 = ~n52902 & ~n52903;
  assign n52905 = ~n52890 & ~n52896;
  assign n52906 = ~n52904 & n52905;
  assign n52907 = n52884 & n52906;
  assign n52908 = ~n52898 & ~n52907;
  assign n52909 = n52878 & ~n52908;
  assign n52910 = n52904 & n52905;
  assign n52911 = ~n52884 & n52910;
  assign n52912 = ~n52890 & n52896;
  assign n52913 = n52904 & n52912;
  assign n52914 = n52884 & n52913;
  assign n52915 = ~n52911 & ~n52914;
  assign n52916 = ~n52909 & n52915;
  assign n52917 = n52890 & n52896;
  assign n52918 = n52904 & n52917;
  assign n52919 = ~n52884 & n52918;
  assign n52920 = ~n52904 & n52912;
  assign n52921 = ~n52878 & n52920;
  assign n52922 = ~n52878 & n52905;
  assign n52923 = ~n52884 & n52922;
  assign n52924 = ~n52921 & ~n52923;
  assign n52925 = ~n52919 & n52924;
  assign n52926 = n52916 & n52925;
  assign n52927 = n52872 & ~n52926;
  assign n52928 = ~n52872 & n52878;
  assign n52929 = ~n52884 & ~n52904;
  assign n52930 = ~n52890 & n52929;
  assign n52931 = n52896 & ~n52904;
  assign n52932 = ~n52930 & ~n52931;
  assign n52933 = n52928 & ~n52932;
  assign n52934 = n52884 & n52904;
  assign n52935 = ~n52896 & n52934;
  assign n52936 = ~n52890 & n52935;
  assign n52937 = n52884 & n52890;
  assign n52938 = ~n52904 & n52937;
  assign n52939 = ~n52936 & ~n52938;
  assign n52940 = ~n52878 & ~n52884;
  assign n52941 = n52904 & n52940;
  assign n52942 = ~n52905 & n52941;
  assign n52943 = ~n52878 & n52918;
  assign n52944 = ~n52942 & ~n52943;
  assign n52945 = n52939 & n52944;
  assign n52946 = ~n52872 & ~n52945;
  assign n52947 = ~n52904 & n52917;
  assign n52948 = n52878 & n52947;
  assign n52949 = n52884 & n52948;
  assign n52950 = n52897 & n52904;
  assign n52951 = n52884 & n52950;
  assign n52952 = ~n52914 & ~n52951;
  assign n52953 = n52878 & ~n52952;
  assign n52954 = ~n52949 & ~n52953;
  assign n52955 = ~n52878 & n52936;
  assign n52956 = n52954 & ~n52955;
  assign n52957 = ~n52946 & n52956;
  assign n52958 = ~n52933 & n52957;
  assign n52959 = ~n52927 & n52958;
  assign n52960 = n52897 & ~n52904;
  assign n52961 = ~n52878 & n52884;
  assign n52962 = n52960 & n52961;
  assign n52963 = n52959 & ~n52962;
  assign n52964 = ~pi1444 & ~n52963;
  assign n52965 = pi1444 & ~n52962;
  assign n52966 = n52958 & n52965;
  assign n52967 = ~n52927 & n52966;
  assign po1531 = n52964 | n52967;
  assign n52969 = pi4794 & pi9040;
  assign n52970 = pi4690 & ~pi9040;
  assign n52971 = ~n52969 & ~n52970;
  assign n52972 = ~pi1435 & n52971;
  assign n52973 = pi1435 & ~n52971;
  assign n52974 = ~n52972 & ~n52973;
  assign n52975 = pi4839 & pi9040;
  assign n52976 = pi4605 & ~pi9040;
  assign n52977 = ~n52975 & ~n52976;
  assign n52978 = ~pi1412 & ~n52977;
  assign n52979 = pi1412 & n52977;
  assign n52980 = ~n52978 & ~n52979;
  assign n52981 = pi4699 & pi9040;
  assign n52982 = pi4620 & ~pi9040;
  assign n52983 = ~n52981 & ~n52982;
  assign n52984 = pi1426 & n52983;
  assign n52985 = ~pi1426 & ~n52983;
  assign n52986 = ~n52984 & ~n52985;
  assign n52987 = ~n52980 & ~n52986;
  assign n52988 = n52974 & n52987;
  assign n52989 = pi4794 & ~pi9040;
  assign n52990 = pi4707 & pi9040;
  assign n52991 = ~n52989 & ~n52990;
  assign n52992 = ~pi1413 & n52991;
  assign n52993 = pi1413 & ~n52991;
  assign n52994 = ~n52992 & ~n52993;
  assign n52995 = ~n52980 & ~n52994;
  assign n52996 = n52986 & n52995;
  assign n52997 = ~n52988 & ~n52996;
  assign n52998 = pi4613 & ~pi9040;
  assign n52999 = pi4716 & pi9040;
  assign n53000 = ~n52998 & ~n52999;
  assign n53001 = ~pi1416 & ~n53000;
  assign n53002 = pi1416 & n53000;
  assign n53003 = ~n53001 & ~n53002;
  assign n53004 = pi4613 & pi9040;
  assign n53005 = pi4607 & ~pi9040;
  assign n53006 = ~n53004 & ~n53005;
  assign n53007 = pi1415 & n53006;
  assign n53008 = ~pi1415 & ~n53006;
  assign n53009 = ~n53007 & ~n53008;
  assign n53010 = n53003 & ~n53009;
  assign n53011 = ~n52997 & n53010;
  assign n53012 = n52980 & ~n52986;
  assign n53013 = ~n52974 & ~n52994;
  assign n53014 = n53012 & n53013;
  assign n53015 = n52980 & n52986;
  assign n53016 = n52994 & n53015;
  assign n53017 = n52987 & n52994;
  assign n53018 = ~n53016 & ~n53017;
  assign n53019 = ~n52974 & ~n53018;
  assign n53020 = ~n53014 & ~n53019;
  assign n53021 = ~n53009 & ~n53020;
  assign n53022 = ~n53011 & ~n53021;
  assign n53023 = ~n52974 & n52994;
  assign n53024 = ~n52980 & n53023;
  assign n53025 = ~n53014 & ~n53024;
  assign n53026 = ~n53003 & ~n53025;
  assign n53027 = n52974 & n53003;
  assign n53028 = n52980 & n53027;
  assign n53029 = n52994 & n53012;
  assign n53030 = ~n52994 & n53015;
  assign n53031 = ~n53029 & ~n53030;
  assign n53032 = n52987 & ~n52994;
  assign n53033 = ~n52974 & n53032;
  assign n53034 = n53031 & ~n53033;
  assign n53035 = n53003 & ~n53034;
  assign n53036 = ~n53028 & ~n53035;
  assign n53037 = ~n52980 & n52986;
  assign n53038 = n52994 & n53037;
  assign n53039 = ~n52974 & n53038;
  assign n53040 = n53036 & ~n53039;
  assign n53041 = ~n52997 & ~n53003;
  assign n53042 = n52974 & n53016;
  assign n53043 = ~n53041 & ~n53042;
  assign n53044 = n53040 & n53043;
  assign n53045 = n53009 & ~n53044;
  assign n53046 = ~n53026 & ~n53045;
  assign n53047 = ~n53003 & ~n53009;
  assign n53048 = n52974 & n53012;
  assign n53049 = ~n53038 & ~n53048;
  assign n53050 = n52980 & ~n52994;
  assign n53051 = n53049 & ~n53050;
  assign n53052 = n53047 & ~n53051;
  assign n53053 = n53046 & ~n53052;
  assign n53054 = n53022 & n53053;
  assign n53055 = ~pi1447 & ~n53054;
  assign n53056 = pi1447 & n53022;
  assign n53057 = n53046 & n53056;
  assign n53058 = ~n53052 & n53057;
  assign po1532 = n53055 | n53058;
  assign n53060 = n52884 & n52920;
  assign n53061 = n52896 & n52929;
  assign n53062 = n52890 & n53061;
  assign n53063 = ~n53060 & ~n53062;
  assign n53064 = ~n52878 & ~n53063;
  assign n53065 = n52878 & n52936;
  assign n53066 = ~n52936 & ~n52943;
  assign n53067 = ~n52890 & n52934;
  assign n53068 = ~n52938 & ~n53067;
  assign n53069 = n52878 & ~n53068;
  assign n53070 = n52878 & ~n52884;
  assign n53071 = n52912 & n53070;
  assign n53072 = ~n52904 & n53071;
  assign n53073 = ~n52884 & n52904;
  assign n53074 = ~n52896 & n53073;
  assign n53075 = n52890 & n53074;
  assign n53076 = ~n52878 & n52906;
  assign n53077 = ~n53075 & ~n53076;
  assign n53078 = ~n53072 & n53077;
  assign n53079 = ~n53069 & n53078;
  assign n53080 = n53066 & n53079;
  assign n53081 = n52872 & ~n53080;
  assign n53082 = n52884 & n52943;
  assign n53083 = ~n53081 & ~n53082;
  assign n53084 = ~n53065 & n53083;
  assign n53085 = ~n53064 & n53084;
  assign n53086 = ~n52890 & n52904;
  assign n53087 = n52940 & n53086;
  assign n53088 = ~n52921 & ~n53087;
  assign n53089 = ~n52878 & n52950;
  assign n53090 = n52884 & n52960;
  assign n53091 = ~n53089 & ~n53090;
  assign n53092 = ~n52884 & n52913;
  assign n53093 = ~n53060 & ~n53092;
  assign n53094 = ~n52884 & n52917;
  assign n53095 = ~n52896 & ~n52904;
  assign n53096 = ~n53094 & ~n53095;
  assign n53097 = n52878 & ~n53096;
  assign n53098 = n53093 & ~n53097;
  assign n53099 = n53091 & n53098;
  assign n53100 = n53088 & n53099;
  assign n53101 = ~n52872 & ~n53100;
  assign n53102 = n53085 & ~n53101;
  assign n53103 = ~pi1446 & ~n53102;
  assign n53104 = pi1446 & n53085;
  assign n53105 = ~n53101 & n53104;
  assign po1536 = n53103 | n53105;
  assign n53107 = ~n53082 & ~n53087;
  assign n53108 = ~n52936 & ~n52947;
  assign n53109 = ~n53094 & n53108;
  assign n53110 = n52878 & ~n53109;
  assign n53111 = ~n52896 & n52929;
  assign n53112 = ~n52890 & n53111;
  assign n53113 = ~n53075 & ~n53112;
  assign n53114 = ~n52962 & n53113;
  assign n53115 = ~n52878 & n52913;
  assign n53116 = n53114 & ~n53115;
  assign n53117 = ~n53110 & n53116;
  assign n53118 = n52872 & ~n53117;
  assign n53119 = n52884 & n52922;
  assign n53120 = n52890 & n52929;
  assign n53121 = ~n52947 & ~n53120;
  assign n53122 = ~n52878 & ~n53121;
  assign n53123 = ~n53119 & ~n53122;
  assign n53124 = n52878 & n52884;
  assign n53125 = n52897 & n53124;
  assign n53126 = n52878 & n52920;
  assign n53127 = ~n53125 & ~n53126;
  assign n53128 = n53123 & n53127;
  assign n53129 = n52890 & n52934;
  assign n53130 = ~n53060 & ~n53129;
  assign n53131 = ~n53092 & n53130;
  assign n53132 = n53128 & n53131;
  assign n53133 = ~n52872 & ~n53132;
  assign n53134 = ~n53060 & n53113;
  assign n53135 = n52878 & ~n53134;
  assign n53136 = ~n53133 & ~n53135;
  assign n53137 = ~n53118 & n53136;
  assign n53138 = n53107 & n53137;
  assign n53139 = pi1450 & ~n53138;
  assign n53140 = ~pi1450 & n53138;
  assign po1537 = n53139 | n53140;
  assign n53142 = n52431 & n52459;
  assign n53143 = ~n52479 & ~n52488;
  assign n53144 = n52437 & ~n53143;
  assign n53145 = ~n52473 & ~n53144;
  assign n53146 = ~n53142 & n53145;
  assign n53147 = ~n52437 & n52476;
  assign n53148 = ~n52465 & ~n53147;
  assign n53149 = ~n52496 & n53148;
  assign n53150 = n53146 & n53149;
  assign n53151 = n52412 & ~n53150;
  assign n53152 = n52445 & n52452;
  assign n53153 = n52431 & n53152;
  assign n53154 = ~n52450 & ~n53153;
  assign n53155 = ~n52431 & n52495;
  assign n53156 = ~n52460 & ~n53155;
  assign n53157 = n52425 & n52445;
  assign n53158 = n52437 & n53157;
  assign n53159 = n52431 & n52464;
  assign n53160 = ~n53158 & ~n53159;
  assign n53161 = n52424 & ~n52445;
  assign n53162 = ~n52418 & n52431;
  assign n53163 = ~n53161 & ~n53162;
  assign n53164 = ~n52501 & n53163;
  assign n53165 = ~n52437 & ~n53164;
  assign n53166 = n53160 & ~n53165;
  assign n53167 = n53156 & n53166;
  assign n53168 = n53154 & n53167;
  assign n53169 = ~n52412 & ~n53168;
  assign n53170 = ~n53151 & ~n53169;
  assign n53171 = pi1440 & ~n53170;
  assign n53172 = ~pi1440 & ~n53151;
  assign n53173 = ~n53169 & n53172;
  assign po1538 = n53171 | n53173;
  assign n53175 = ~n52515 & n52521;
  assign n53176 = ~n52594 & ~n53175;
  assign n53177 = ~n52536 & n53176;
  assign n53178 = ~n52527 & ~n53177;
  assign n53179 = n52515 & n52568;
  assign n53180 = n52521 & ~n52535;
  assign n53181 = n52544 & n53180;
  assign n53182 = n52535 & n52586;
  assign n53183 = ~n53181 & ~n53182;
  assign n53184 = ~n52515 & ~n52521;
  assign n53185 = n52527 & n52535;
  assign n53186 = n53184 & n53185;
  assign n53187 = n53183 & ~n53186;
  assign n53188 = ~n53179 & n53187;
  assign n53189 = ~n53178 & n53188;
  assign n53190 = n52566 & ~n53189;
  assign n53191 = n52521 & n52552;
  assign n53192 = ~n52535 & n53191;
  assign n53193 = n52521 & n52545;
  assign n53194 = n52535 & n53193;
  assign n53195 = ~n53192 & ~n53194;
  assign n53196 = ~n52527 & ~n53195;
  assign n53197 = ~n53190 & ~n53196;
  assign n53198 = ~n52535 & n52586;
  assign n53199 = ~n52549 & ~n52598;
  assign n53200 = ~n52527 & ~n53199;
  assign n53201 = ~n53198 & ~n53200;
  assign n53202 = ~n52601 & n53201;
  assign n53203 = ~n52566 & ~n53202;
  assign n53204 = ~n52552 & ~n52580;
  assign n53205 = ~n52521 & ~n53204;
  assign n53206 = ~n52572 & ~n53205;
  assign n53207 = n52527 & ~n53206;
  assign n53208 = ~n52566 & n53207;
  assign n53209 = ~n53203 & ~n53208;
  assign n53210 = n53197 & n53209;
  assign n53211 = pi1451 & ~n53210;
  assign n53212 = ~pi1451 & n53197;
  assign n53213 = n53209 & n53212;
  assign po1539 = n53211 | n53213;
  assign n53215 = ~n52974 & n53017;
  assign n53216 = n52974 & n53050;
  assign n53217 = ~n53215 & ~n53216;
  assign n53218 = n53003 & ~n53217;
  assign n53219 = n52986 & n53013;
  assign n53220 = ~n52980 & n53219;
  assign n53221 = n52974 & n53038;
  assign n53222 = ~n53220 & ~n53221;
  assign n53223 = ~n53003 & ~n53222;
  assign n53224 = ~n52974 & ~n53003;
  assign n53225 = ~n52987 & ~n53016;
  assign n53226 = n53224 & ~n53225;
  assign n53227 = n52994 & ~n53003;
  assign n53228 = n52987 & n53227;
  assign n53229 = ~n53226 & ~n53228;
  assign n53230 = n53009 & ~n53229;
  assign n53231 = n52974 & n53030;
  assign n53232 = n52974 & ~n52994;
  assign n53233 = ~n53050 & ~n53232;
  assign n53234 = n53003 & ~n53233;
  assign n53235 = n52974 & n52994;
  assign n53236 = ~n52986 & n53235;
  assign n53237 = n52980 & n53236;
  assign n53238 = ~n53234 & ~n53237;
  assign n53239 = ~n53231 & n53238;
  assign n53240 = n53009 & ~n53239;
  assign n53241 = ~n53230 & ~n53240;
  assign n53242 = ~n53012 & ~n53050;
  assign n53243 = ~n52974 & ~n53242;
  assign n53244 = ~n53038 & ~n53243;
  assign n53245 = ~n53003 & ~n53244;
  assign n53246 = n52974 & n52986;
  assign n53247 = n53227 & n53246;
  assign n53248 = ~n52986 & ~n52994;
  assign n53249 = ~n53038 & ~n53248;
  assign n53250 = n52974 & ~n53249;
  assign n53251 = ~n52974 & n53003;
  assign n53252 = n53015 & n53251;
  assign n53253 = n52994 & n53252;
  assign n53254 = ~n53250 & ~n53253;
  assign n53255 = ~n53247 & n53254;
  assign n53256 = ~n53245 & n53255;
  assign n53257 = ~n53220 & n53256;
  assign n53258 = ~n53009 & ~n53257;
  assign n53259 = n53241 & ~n53258;
  assign n53260 = ~n53223 & n53259;
  assign n53261 = ~n53218 & n53260;
  assign n53262 = pi1458 & n53261;
  assign n53263 = ~pi1458 & ~n53261;
  assign po1541 = n53262 | n53263;
  assign n53265 = n52743 & n52764;
  assign n53266 = ~n52737 & n53265;
  assign n53267 = ~n52857 & ~n53266;
  assign n53268 = n52731 & n52737;
  assign n53269 = ~n52725 & n53268;
  assign n53270 = n52725 & n52836;
  assign n53271 = ~n52737 & n52752;
  assign n53272 = ~n53270 & ~n53271;
  assign n53273 = ~n52743 & ~n53272;
  assign n53274 = ~n53269 & ~n53273;
  assign n53275 = n53267 & n53274;
  assign n53276 = n52762 & ~n53275;
  assign n53277 = ~n52766 & ~n52805;
  assign n53278 = ~n52737 & n52794;
  assign n53279 = n53277 & ~n53278;
  assign n53280 = n52743 & ~n53279;
  assign n53281 = n52764 & n52800;
  assign n53282 = ~n52755 & ~n53281;
  assign n53283 = ~n53280 & n53282;
  assign n53284 = ~n52776 & ~n52785;
  assign n53285 = ~n52743 & ~n53284;
  assign n53286 = n53283 & ~n53285;
  assign n53287 = ~n52762 & ~n53286;
  assign n53288 = ~n53276 & ~n53287;
  assign n53289 = ~n52737 & n52775;
  assign n53290 = n52737 & ~n52780;
  assign n53291 = ~n53289 & ~n53290;
  assign n53292 = ~n52743 & ~n53291;
  assign n53293 = ~n52789 & ~n52795;
  assign n53294 = ~n52766 & n53293;
  assign n53295 = n52848 & ~n53294;
  assign n53296 = ~n53292 & ~n53295;
  assign n53297 = n53288 & n53296;
  assign n53298 = ~pi1466 & ~n53297;
  assign n53299 = pi1466 & n53296;
  assign n53300 = ~n53287 & n53299;
  assign n53301 = ~n53276 & n53300;
  assign po1542 = n53298 | n53301;
  assign n53303 = pi4608 & pi9040;
  assign n53304 = pi4937 & ~pi9040;
  assign n53305 = ~n53303 & ~n53304;
  assign n53306 = ~pi1411 & ~n53305;
  assign n53307 = pi1411 & n53305;
  assign n53308 = ~n53306 & ~n53307;
  assign n53309 = pi4710 & pi9040;
  assign n53310 = pi4692 & ~pi9040;
  assign n53311 = ~n53309 & ~n53310;
  assign n53312 = pi1439 & n53311;
  assign n53313 = ~pi1439 & ~n53311;
  assign n53314 = ~n53312 & ~n53313;
  assign n53315 = pi4736 & pi9040;
  assign n53316 = pi4883 & ~pi9040;
  assign n53317 = ~n53315 & ~n53316;
  assign n53318 = pi1405 & n53317;
  assign n53319 = ~pi1405 & ~n53317;
  assign n53320 = ~n53318 & ~n53319;
  assign n53321 = ~n53314 & ~n53320;
  assign n53322 = pi4781 & pi9040;
  assign n53323 = pi4958 & ~pi9040;
  assign n53324 = ~n53322 & ~n53323;
  assign n53325 = ~pi1436 & n53324;
  assign n53326 = pi1436 & ~n53324;
  assign n53327 = ~n53325 & ~n53326;
  assign n53328 = n53321 & ~n53327;
  assign n53329 = pi4883 & pi9040;
  assign n53330 = pi4695 & ~pi9040;
  assign n53331 = ~n53329 & ~n53330;
  assign n53332 = pi1418 & n53331;
  assign n53333 = ~pi1418 & ~n53331;
  assign n53334 = ~n53332 & ~n53333;
  assign n53335 = pi4774 & ~pi9040;
  assign n53336 = pi4949 & pi9040;
  assign n53337 = ~n53335 & ~n53336;
  assign n53338 = pi1432 & n53337;
  assign n53339 = ~pi1432 & ~n53337;
  assign n53340 = ~n53338 & ~n53339;
  assign n53341 = n53327 & ~n53340;
  assign n53342 = n53334 & n53341;
  assign n53343 = n53314 & n53342;
  assign n53344 = n53327 & n53340;
  assign n53345 = ~n53334 & n53344;
  assign n53346 = n53314 & n53345;
  assign n53347 = ~n53343 & ~n53346;
  assign n53348 = ~n53327 & n53340;
  assign n53349 = ~n53334 & n53348;
  assign n53350 = ~n53314 & ~n53334;
  assign n53351 = ~n53340 & n53350;
  assign n53352 = n53327 & n53351;
  assign n53353 = ~n53349 & ~n53352;
  assign n53354 = n53320 & ~n53353;
  assign n53355 = n53347 & ~n53354;
  assign n53356 = ~n53328 & n53355;
  assign n53357 = n53308 & ~n53356;
  assign n53358 = ~n53327 & ~n53340;
  assign n53359 = ~n53334 & n53358;
  assign n53360 = n53314 & n53359;
  assign n53361 = ~n53320 & n53360;
  assign n53362 = ~n53314 & n53320;
  assign n53363 = n53359 & n53362;
  assign n53364 = ~n53314 & n53334;
  assign n53365 = n53327 & n53364;
  assign n53366 = ~n53363 & ~n53365;
  assign n53367 = n53334 & n53344;
  assign n53368 = ~n53349 & ~n53367;
  assign n53369 = ~n53314 & n53344;
  assign n53370 = n53368 & ~n53369;
  assign n53371 = ~n53320 & ~n53370;
  assign n53372 = n53334 & ~n53340;
  assign n53373 = ~n53327 & n53372;
  assign n53374 = n53314 & n53373;
  assign n53375 = ~n53334 & n53341;
  assign n53376 = n53314 & n53375;
  assign n53377 = ~n53374 & ~n53376;
  assign n53378 = n53334 & n53348;
  assign n53379 = n53320 & n53378;
  assign n53380 = n53377 & ~n53379;
  assign n53381 = ~n53371 & n53380;
  assign n53382 = n53366 & n53381;
  assign n53383 = ~n53308 & ~n53382;
  assign n53384 = ~n53361 & ~n53383;
  assign n53385 = ~n53357 & n53384;
  assign n53386 = n53362 & n53367;
  assign n53387 = n53320 & n53372;
  assign n53388 = n53314 & n53387;
  assign n53389 = ~n53386 & ~n53388;
  assign n53390 = n53320 & n53346;
  assign n53391 = n53389 & ~n53390;
  assign n53392 = n53385 & n53391;
  assign n53393 = ~pi1448 & ~n53392;
  assign n53394 = pi1448 & n53391;
  assign n53395 = n53384 & n53394;
  assign n53396 = ~n53357 & n53395;
  assign po1543 = n53393 | n53396;
  assign n53398 = ~n53334 & ~n53340;
  assign n53399 = ~n53314 & n53398;
  assign n53400 = n53314 & n53341;
  assign n53401 = ~n53399 & ~n53400;
  assign n53402 = n53327 & ~n53334;
  assign n53403 = n53401 & ~n53402;
  assign n53404 = ~n53378 & n53403;
  assign n53405 = n53320 & ~n53404;
  assign n53406 = n53340 & n53364;
  assign n53407 = ~n53349 & ~n53365;
  assign n53408 = ~n53320 & ~n53407;
  assign n53409 = ~n53406 & ~n53408;
  assign n53410 = ~n53405 & n53409;
  assign n53411 = ~n53374 & n53410;
  assign n53412 = n53308 & ~n53411;
  assign n53413 = ~n53314 & n53345;
  assign n53414 = n53377 & ~n53413;
  assign n53415 = n53320 & ~n53414;
  assign n53416 = ~n53412 & ~n53415;
  assign n53417 = ~n53314 & n53378;
  assign n53418 = ~n53327 & ~n53334;
  assign n53419 = ~n53320 & n53418;
  assign n53420 = n53314 & n53419;
  assign n53421 = n53334 & n53362;
  assign n53422 = ~n53340 & n53421;
  assign n53423 = n53314 & n53367;
  assign n53424 = ~n53422 & ~n53423;
  assign n53425 = n53327 & n53334;
  assign n53426 = n53314 & n53425;
  assign n53427 = ~n53359 & ~n53426;
  assign n53428 = ~n53320 & ~n53427;
  assign n53429 = ~n53320 & n53327;
  assign n53430 = ~n53334 & n53429;
  assign n53431 = ~n53314 & n53430;
  assign n53432 = ~n53428 & ~n53431;
  assign n53433 = n53424 & n53432;
  assign n53434 = ~n53308 & ~n53433;
  assign n53435 = ~n53420 & ~n53434;
  assign n53436 = ~n53417 & n53435;
  assign n53437 = n53416 & n53436;
  assign n53438 = ~pi1445 & ~n53437;
  assign n53439 = ~n53412 & ~n53417;
  assign n53440 = ~n53415 & n53439;
  assign n53441 = n53435 & n53440;
  assign n53442 = pi1445 & n53441;
  assign po1544 = n53438 | n53442;
  assign n53444 = pi4891 & pi9040;
  assign n53445 = pi4716 & ~pi9040;
  assign n53446 = ~n53444 & ~n53445;
  assign n53447 = pi1426 & n53446;
  assign n53448 = ~pi1426 & ~n53446;
  assign n53449 = ~n53447 & ~n53448;
  assign n53450 = pi4607 & pi9040;
  assign n53451 = pi4685 & ~pi9040;
  assign n53452 = ~n53450 & ~n53451;
  assign n53453 = pi1429 & n53452;
  assign n53454 = ~pi1429 & ~n53452;
  assign n53455 = ~n53453 & ~n53454;
  assign n53456 = pi4685 & pi9040;
  assign n53457 = pi4699 & ~pi9040;
  assign n53458 = ~n53456 & ~n53457;
  assign n53459 = ~pi1415 & n53458;
  assign n53460 = pi1415 & ~n53458;
  assign n53461 = ~n53459 & ~n53460;
  assign n53462 = n53455 & ~n53461;
  assign n53463 = n53449 & n53462;
  assign n53464 = ~n53455 & ~n53461;
  assign n53465 = ~n53449 & n53464;
  assign n53466 = ~n53463 & ~n53465;
  assign n53467 = pi4611 & pi9040;
  assign n53468 = pi4734 & ~pi9040;
  assign n53469 = ~n53467 & ~n53468;
  assign n53470 = pi1422 & n53469;
  assign n53471 = ~pi1422 & ~n53469;
  assign n53472 = ~n53470 & ~n53471;
  assign n53473 = n53449 & ~n53472;
  assign n53474 = n53455 & n53473;
  assign n53475 = n53466 & ~n53474;
  assign n53476 = pi4623 & pi9040;
  assign n53477 = pi4891 & ~pi9040;
  assign n53478 = ~n53476 & ~n53477;
  assign n53479 = ~pi1395 & n53478;
  assign n53480 = pi1395 & ~n53478;
  assign n53481 = ~n53479 & ~n53480;
  assign n53482 = pi4618 & pi9040;
  assign n53483 = pi4610 & ~pi9040;
  assign n53484 = ~n53482 & ~n53483;
  assign n53485 = ~pi1420 & ~n53484;
  assign n53486 = pi1420 & n53484;
  assign n53487 = ~n53485 & ~n53486;
  assign n53488 = n53481 & n53487;
  assign n53489 = ~n53475 & n53488;
  assign n53490 = ~n53455 & n53461;
  assign n53491 = n53449 & n53490;
  assign n53492 = n53472 & n53487;
  assign n53493 = n53491 & n53492;
  assign n53494 = n53449 & n53464;
  assign n53495 = ~n53481 & n53494;
  assign n53496 = n53455 & n53461;
  assign n53497 = n53472 & n53496;
  assign n53498 = ~n53449 & n53455;
  assign n53499 = ~n53497 & ~n53498;
  assign n53500 = ~n53481 & ~n53499;
  assign n53501 = ~n53495 & ~n53500;
  assign n53502 = n53487 & ~n53501;
  assign n53503 = ~n53493 & ~n53502;
  assign n53504 = ~n53449 & ~n53472;
  assign n53505 = ~n53455 & n53504;
  assign n53506 = n53461 & n53505;
  assign n53507 = ~n53449 & n53472;
  assign n53508 = n53455 & n53507;
  assign n53509 = ~n53506 & ~n53508;
  assign n53510 = ~n53481 & ~n53509;
  assign n53511 = n53503 & ~n53510;
  assign n53512 = n53472 & n53481;
  assign n53513 = n53496 & n53512;
  assign n53514 = n53449 & n53513;
  assign n53515 = ~n53462 & ~n53490;
  assign n53516 = n53473 & ~n53515;
  assign n53517 = ~n53461 & n53505;
  assign n53518 = ~n53516 & ~n53517;
  assign n53519 = n53507 & ~n53515;
  assign n53520 = n53472 & n53494;
  assign n53521 = ~n53519 & ~n53520;
  assign n53522 = ~n53449 & n53496;
  assign n53523 = ~n53472 & n53481;
  assign n53524 = n53522 & n53523;
  assign n53525 = n53521 & ~n53524;
  assign n53526 = n53518 & n53525;
  assign n53527 = ~n53514 & n53526;
  assign n53528 = ~n53472 & ~n53481;
  assign n53529 = n53449 & n53528;
  assign n53530 = n53461 & n53529;
  assign n53531 = n53527 & ~n53530;
  assign n53532 = ~n53487 & ~n53531;
  assign n53533 = n53511 & ~n53532;
  assign n53534 = ~n53489 & n53533;
  assign n53535 = ~pi1461 & ~n53534;
  assign n53536 = pi1461 & n53511;
  assign n53537 = ~n53489 & n53536;
  assign n53538 = ~n53532 & n53537;
  assign po1545 = n53535 | n53538;
  assign n53540 = ~n52743 & ~n53293;
  assign n53541 = n52737 & n52779;
  assign n53542 = ~n53540 & ~n53541;
  assign n53543 = n52737 & ~n52752;
  assign n53544 = ~n52803 & ~n53543;
  assign n53545 = ~n52776 & n53544;
  assign n53546 = n52743 & ~n53545;
  assign n53547 = n53542 & ~n53546;
  assign n53548 = ~n52762 & ~n53547;
  assign n53549 = ~n52743 & n52824;
  assign n53550 = ~n52838 & ~n53549;
  assign n53551 = ~n52840 & n53550;
  assign n53552 = ~n52808 & ~n53270;
  assign n53553 = n52743 & n52843;
  assign n53554 = n52737 & n52795;
  assign n53555 = ~n52743 & n52803;
  assign n53556 = ~n53554 & ~n53555;
  assign n53557 = ~n52802 & n53556;
  assign n53558 = ~n53553 & n53557;
  assign n53559 = n53552 & n53558;
  assign n53560 = ~n52851 & n53559;
  assign n53561 = n52762 & ~n53560;
  assign n53562 = n53551 & ~n53561;
  assign n53563 = ~n53548 & n53562;
  assign n53564 = ~pi1468 & ~n53563;
  assign n53565 = pi1468 & n53551;
  assign n53566 = ~n53548 & n53565;
  assign n53567 = ~n53561 & n53566;
  assign po1546 = n53564 | n53567;
  assign n53569 = n52535 & n52546;
  assign n53570 = ~n53182 & ~n53569;
  assign n53571 = n52527 & ~n53570;
  assign n53572 = n52568 & n52598;
  assign n53573 = ~n53571 & ~n53572;
  assign n53574 = ~n52612 & n53573;
  assign n53575 = ~n52535 & n52549;
  assign n53576 = ~n52546 & ~n53575;
  assign n53577 = ~n53191 & n53576;
  assign n53578 = n52527 & ~n53577;
  assign n53579 = n52566 & n53578;
  assign n53580 = ~n52527 & n53193;
  assign n53581 = ~n52594 & ~n52606;
  assign n53582 = ~n52588 & n53581;
  assign n53583 = ~n53580 & n53582;
  assign n53584 = n52566 & ~n53583;
  assign n53585 = n52521 & ~n52527;
  assign n53586 = ~n52544 & n53585;
  assign n53587 = ~n52515 & n53586;
  assign n53588 = ~n52535 & n52557;
  assign n53589 = ~n53587 & ~n53588;
  assign n53590 = ~n53181 & n53589;
  assign n53591 = ~n52544 & n52592;
  assign n53592 = ~n52535 & n52580;
  assign n53593 = ~n52597 & ~n53592;
  assign n53594 = n52527 & ~n53593;
  assign n53595 = ~n53591 & ~n53594;
  assign n53596 = n53590 & n53595;
  assign n53597 = ~n52566 & ~n53596;
  assign n53598 = n52535 & n53587;
  assign n53599 = ~n53597 & ~n53598;
  assign n53600 = ~n53584 & n53599;
  assign n53601 = ~n53579 & n53600;
  assign n53602 = n53574 & n53601;
  assign n53603 = pi1459 & ~n53602;
  assign n53604 = ~pi1459 & n53574;
  assign n53605 = n53601 & n53604;
  assign po1547 = n53603 | n53605;
  assign n53607 = ~n52431 & n52452;
  assign n53608 = ~n53155 & ~n53607;
  assign n53609 = n52437 & n53608;
  assign n53610 = ~n52425 & ~n52446;
  assign n53611 = ~n52445 & ~n53610;
  assign n53612 = n52418 & n52477;
  assign n53613 = n52431 & n52446;
  assign n53614 = ~n53612 & ~n53613;
  assign n53615 = n52431 & n52490;
  assign n53616 = n53614 & ~n53615;
  assign n53617 = ~n53611 & n53616;
  assign n53618 = ~n52437 & n53617;
  assign n53619 = ~n53609 & ~n53618;
  assign n53620 = n52431 & n53611;
  assign n53621 = ~n53153 & ~n53620;
  assign n53622 = ~n53619 & n53621;
  assign n53623 = n52412 & ~n53622;
  assign n53624 = n52437 & ~n53610;
  assign n53625 = ~n52431 & n53624;
  assign n53626 = ~n52466 & ~n52494;
  assign n53627 = n52431 & ~n53626;
  assign n53628 = n52437 & n53627;
  assign n53629 = n52445 & n53624;
  assign n53630 = ~n53628 & ~n53629;
  assign n53631 = ~n53625 & n53630;
  assign n53632 = ~n52412 & ~n53631;
  assign n53633 = ~n53623 & ~n53632;
  assign n53634 = ~n52437 & ~n53608;
  assign n53635 = ~n52450 & ~n53634;
  assign n53636 = ~n52412 & ~n53635;
  assign n53637 = n52437 & n52450;
  assign n53638 = ~n52437 & ~n53621;
  assign n53639 = ~n53637 & ~n53638;
  assign n53640 = ~n53636 & n53639;
  assign n53641 = n53633 & n53640;
  assign n53642 = pi1462 & ~n53641;
  assign n53643 = ~n53623 & n53640;
  assign n53644 = ~n53632 & n53643;
  assign n53645 = ~pi1462 & n53644;
  assign po1548 = n53642 | n53645;
  assign n53647 = n53463 & n53481;
  assign n53648 = n53472 & n53647;
  assign n53649 = n53481 & ~n53487;
  assign n53650 = ~n53494 & ~n53497;
  assign n53651 = n53504 & ~n53515;
  assign n53652 = n53650 & ~n53651;
  assign n53653 = n53649 & ~n53652;
  assign n53654 = n53465 & n53472;
  assign n53655 = ~n53461 & n53472;
  assign n53656 = ~n53449 & n53655;
  assign n53657 = n53472 & n53490;
  assign n53658 = ~n53656 & ~n53657;
  assign n53659 = ~n53472 & n53496;
  assign n53660 = ~n53491 & ~n53659;
  assign n53661 = n53658 & n53660;
  assign n53662 = ~n53481 & ~n53661;
  assign n53663 = ~n53654 & ~n53662;
  assign n53664 = ~n53487 & ~n53663;
  assign n53665 = ~n53653 & ~n53664;
  assign n53666 = ~n53648 & n53665;
  assign n53667 = n53449 & n53496;
  assign n53668 = ~n53481 & n53667;
  assign n53669 = ~n53472 & n53668;
  assign n53670 = n53464 & n53528;
  assign n53671 = ~n53449 & n53670;
  assign n53672 = ~n53669 & ~n53671;
  assign n53673 = ~n53517 & ~n53524;
  assign n53674 = n53449 & ~n53461;
  assign n53675 = n53472 & n53674;
  assign n53676 = ~n53497 & ~n53675;
  assign n53677 = ~n53481 & ~n53676;
  assign n53678 = n53481 & ~n53504;
  assign n53679 = ~n53515 & n53678;
  assign n53680 = ~n53496 & n53528;
  assign n53681 = ~n53449 & n53680;
  assign n53682 = ~n53679 & ~n53681;
  assign n53683 = ~n53677 & n53682;
  assign n53684 = n53673 & n53683;
  assign n53685 = n53487 & ~n53684;
  assign n53686 = n53672 & ~n53685;
  assign n53687 = ~pi1454 & n53686;
  assign n53688 = n53666 & n53687;
  assign n53689 = n53666 & n53686;
  assign n53690 = pi1454 & ~n53689;
  assign po1549 = n53688 | n53690;
  assign n53692 = ~n52535 & n53205;
  assign n53693 = ~n52548 & ~n53193;
  assign n53694 = n52527 & ~n53693;
  assign n53695 = ~n53692 & ~n53694;
  assign n53696 = ~n52544 & n53180;
  assign n53697 = ~n52554 & ~n53696;
  assign n53698 = ~n53191 & n53697;
  assign n53699 = ~n52527 & ~n53698;
  assign n53700 = n53695 & ~n53699;
  assign n53701 = n52535 & n52598;
  assign n53702 = n53700 & ~n53701;
  assign n53703 = ~n52566 & ~n53702;
  assign n53704 = n52581 & ~n53693;
  assign n53705 = ~n52546 & ~n52549;
  assign n53706 = ~n52598 & ~n53191;
  assign n53707 = n53705 & n53706;
  assign n53708 = ~n52535 & ~n53707;
  assign n53709 = ~n53704 & ~n53708;
  assign n53710 = ~n53182 & n53709;
  assign n53711 = n52566 & ~n53710;
  assign n53712 = ~n53703 & ~n53711;
  assign n53713 = ~n52535 & n53193;
  assign n53714 = ~n53701 & ~n53713;
  assign n53715 = n52527 & ~n53714;
  assign n53716 = n53712 & ~n53715;
  assign n53717 = pi1471 & ~n53716;
  assign n53718 = ~pi1471 & ~n53715;
  assign n53719 = ~n53711 & n53718;
  assign n53720 = ~n53703 & n53719;
  assign po1550 = n53717 | n53720;
  assign n53722 = ~n53314 & n53342;
  assign n53723 = ~n53345 & ~n53417;
  assign n53724 = n53314 & n53372;
  assign n53725 = ~n53314 & n53359;
  assign n53726 = ~n53724 & ~n53725;
  assign n53727 = n53723 & n53726;
  assign n53728 = ~n53320 & ~n53727;
  assign n53729 = n53314 & n53348;
  assign n53730 = ~n53365 & ~n53729;
  assign n53731 = ~n53375 & n53730;
  assign n53732 = n53320 & ~n53731;
  assign n53733 = n53314 & ~n53334;
  assign n53734 = n53340 & n53733;
  assign n53735 = ~n53327 & n53734;
  assign n53736 = ~n53732 & ~n53735;
  assign n53737 = ~n53728 & n53736;
  assign n53738 = ~n53722 & n53737;
  assign n53739 = ~n53308 & ~n53738;
  assign n53740 = n53314 & ~n53320;
  assign n53741 = n53378 & n53740;
  assign n53742 = ~n53320 & n53375;
  assign n53743 = ~n53320 & n53367;
  assign n53744 = ~n53742 & ~n53743;
  assign n53745 = ~n53314 & ~n53744;
  assign n53746 = ~n53741 & ~n53745;
  assign n53747 = n53314 & n53344;
  assign n53748 = ~n53314 & n53348;
  assign n53749 = ~n53747 & ~n53748;
  assign n53750 = ~n53373 & n53749;
  assign n53751 = ~n53345 & n53750;
  assign n53752 = n53320 & ~n53751;
  assign n53753 = ~n53314 & n53349;
  assign n53754 = ~n53752 & ~n53753;
  assign n53755 = ~n53314 & n53373;
  assign n53756 = ~n53360 & ~n53755;
  assign n53757 = n53754 & n53756;
  assign n53758 = n53746 & n53757;
  assign n53759 = n53308 & ~n53758;
  assign n53760 = ~n53320 & ~n53347;
  assign n53761 = ~n53759 & ~n53760;
  assign n53762 = ~n53376 & ~n53755;
  assign n53763 = n53320 & ~n53762;
  assign n53764 = n53761 & ~n53763;
  assign n53765 = ~n53739 & n53764;
  assign n53766 = pi1456 & ~n53765;
  assign n53767 = ~pi1456 & n53765;
  assign po1551 = n53766 | n53767;
  assign n53769 = n52630 & ~n52636;
  assign n53770 = ~n52624 & n53769;
  assign n53771 = n52650 & n53770;
  assign n53772 = n52644 & n52650;
  assign n53773 = ~n52630 & ~n52642;
  assign n53774 = ~n52650 & n53773;
  assign n53775 = ~n52657 & ~n53774;
  assign n53776 = ~n53772 & n53775;
  assign n53777 = ~n53771 & n53776;
  assign n53778 = n52624 & n52653;
  assign n53779 = n53777 & ~n53778;
  assign n53780 = n52689 & ~n53779;
  assign n53781 = n52630 & n52676;
  assign n53782 = ~n52650 & n53781;
  assign n53783 = ~n52630 & ~n52650;
  assign n53784 = n52636 & n53783;
  assign n53785 = ~n53773 & ~n53784;
  assign n53786 = ~n52659 & n53785;
  assign n53787 = n52624 & ~n53786;
  assign n53788 = ~n53782 & ~n53787;
  assign n53789 = ~n52689 & ~n53788;
  assign n53790 = ~n52650 & n52659;
  assign n53791 = ~n52707 & ~n53790;
  assign n53792 = n52624 & ~n53791;
  assign n53793 = ~n52624 & ~n52689;
  assign n53794 = n52691 & n53793;
  assign n53795 = ~n53792 & ~n53794;
  assign n53796 = ~n53789 & n53795;
  assign n53797 = ~n52642 & n52650;
  assign n53798 = n52630 & n53797;
  assign n53799 = ~n52650 & n52706;
  assign n53800 = ~n53798 & ~n53799;
  assign n53801 = ~n52654 & n53800;
  assign n53802 = ~n52657 & n53801;
  assign n53803 = ~n52624 & ~n53802;
  assign n53804 = n53796 & ~n53803;
  assign n53805 = ~n53780 & n53804;
  assign n53806 = ~pi1492 & ~n53805;
  assign n53807 = pi1492 & n53796;
  assign n53808 = ~n53780 & n53807;
  assign n53809 = ~n53803 & n53808;
  assign po1552 = n53806 | n53809;
  assign n53811 = ~n52919 & ~n52930;
  assign n53812 = n52872 & ~n53811;
  assign n53813 = ~n52935 & ~n53067;
  assign n53814 = ~n52910 & n53813;
  assign n53815 = n52878 & ~n53814;
  assign n53816 = n52872 & n53815;
  assign n53817 = ~n53812 & ~n53816;
  assign n53818 = n52918 & n53070;
  assign n53819 = ~n53072 & ~n53818;
  assign n53820 = ~n52938 & ~n53095;
  assign n53821 = ~n52878 & ~n53820;
  assign n53822 = n52872 & n53821;
  assign n53823 = n53819 & ~n53822;
  assign n53824 = n52884 & n52918;
  assign n53825 = n52884 & n52912;
  assign n53826 = ~n53062 & ~n53825;
  assign n53827 = ~n52878 & ~n53826;
  assign n53828 = ~n52936 & ~n53075;
  assign n53829 = n52884 & n52917;
  assign n53830 = ~n52960 & ~n53829;
  assign n53831 = n52878 & ~n53830;
  assign n53832 = n53828 & ~n53831;
  assign n53833 = ~n53827 & n53832;
  assign n53834 = ~n53824 & n53833;
  assign n53835 = ~n52872 & ~n53834;
  assign n53836 = ~n53092 & n53113;
  assign n53837 = ~n52878 & ~n53836;
  assign n53838 = ~n53835 & ~n53837;
  assign n53839 = n53823 & n53838;
  assign n53840 = n53817 & n53839;
  assign n53841 = ~pi1457 & ~n53840;
  assign n53842 = pi1457 & n53823;
  assign n53843 = n53817 & n53842;
  assign n53844 = n53838 & n53843;
  assign po1553 = n53841 | n53844;
  assign n53846 = n52642 & n52698;
  assign n53847 = ~n52666 & ~n53846;
  assign n53848 = ~n52677 & ~n53798;
  assign n53849 = n52624 & ~n53848;
  assign n53850 = ~n52624 & ~n52630;
  assign n53851 = n52652 & n53850;
  assign n53852 = ~n53849 & ~n53851;
  assign n53853 = ~n52650 & n52680;
  assign n53854 = ~n52654 & ~n53853;
  assign n53855 = ~n52624 & ~n52650;
  assign n53856 = ~n52642 & n53855;
  assign n53857 = ~n52636 & n53856;
  assign n53858 = n52658 & n52692;
  assign n53859 = ~n53857 & ~n53858;
  assign n53860 = n53854 & n53859;
  assign n53861 = n53852 & n53860;
  assign n53862 = n53847 & n53861;
  assign n53863 = ~n52689 & ~n53862;
  assign n53864 = ~n52653 & ~n52677;
  assign n53865 = n52650 & ~n53864;
  assign n53866 = ~n52636 & n52695;
  assign n53867 = ~n52706 & ~n53866;
  assign n53868 = n52650 & n53773;
  assign n53869 = n53867 & ~n53868;
  assign n53870 = n52624 & ~n53869;
  assign n53871 = ~n52650 & n52676;
  assign n53872 = ~n53772 & ~n53871;
  assign n53873 = ~n52624 & ~n53872;
  assign n53874 = ~n53790 & ~n53873;
  assign n53875 = ~n53870 & n53874;
  assign n53876 = ~n53865 & n53875;
  assign n53877 = n52689 & ~n53876;
  assign n53878 = n52624 & n52696;
  assign n53879 = ~n53877 & ~n53878;
  assign n53880 = n52671 & n53855;
  assign n53881 = ~n52642 & n53880;
  assign n53882 = n53879 & ~n53881;
  assign n53883 = ~n53863 & n53882;
  assign n53884 = ~pi1465 & ~n53883;
  assign n53885 = pi1465 & n53879;
  assign n53886 = ~n53863 & n53885;
  assign n53887 = ~n53881 & n53886;
  assign po1554 = n53884 | n53887;
  assign n53889 = ~n52986 & n53023;
  assign n53890 = ~n53016 & ~n53889;
  assign n53891 = ~n53003 & ~n53890;
  assign n53892 = ~n52974 & n53037;
  assign n53893 = ~n53236 & ~n53892;
  assign n53894 = n53003 & ~n53893;
  assign n53895 = n52974 & n53032;
  assign n53896 = ~n53247 & ~n53895;
  assign n53897 = ~n53014 & n53896;
  assign n53898 = ~n53894 & n53897;
  assign n53899 = ~n53891 & n53898;
  assign n53900 = ~n53220 & ~n53231;
  assign n53901 = n53899 & n53900;
  assign n53902 = n53009 & ~n53901;
  assign n53903 = n53012 & n53232;
  assign n53904 = n53018 & ~n53903;
  assign n53905 = n53003 & ~n53904;
  assign n53906 = n52974 & n52996;
  assign n53907 = ~n53905 & ~n53906;
  assign n53908 = n52980 & n53023;
  assign n53909 = ~n52974 & n53015;
  assign n53910 = ~n53908 & ~n53909;
  assign n53911 = n53003 & ~n53910;
  assign n53912 = n53003 & n53037;
  assign n53913 = n52974 & n53912;
  assign n53914 = ~n53911 & ~n53913;
  assign n53915 = n53907 & n53914;
  assign n53916 = ~n53009 & ~n53915;
  assign n53917 = ~n53032 & ~n53039;
  assign n53918 = ~n53237 & n53917;
  assign n53919 = n53047 & ~n53918;
  assign n53920 = ~n53916 & ~n53919;
  assign n53921 = ~n53014 & ~n53231;
  assign n53922 = ~n53003 & ~n53921;
  assign n53923 = n53920 & ~n53922;
  assign n53924 = ~n53902 & n53923;
  assign n53925 = ~pi1472 & n53924;
  assign n53926 = pi1472 & ~n53924;
  assign po1555 = n53925 | n53926;
  assign n53928 = ~n52651 & ~n52657;
  assign n53929 = ~n52624 & ~n53928;
  assign n53930 = ~n52713 & ~n53929;
  assign n53931 = n52630 & n52636;
  assign n53932 = n52624 & n53931;
  assign n53933 = n52650 & n53932;
  assign n53934 = n52650 & n52676;
  assign n53935 = ~n53931 & ~n53934;
  assign n53936 = ~n52636 & n53783;
  assign n53937 = n53935 & ~n53936;
  assign n53938 = n52624 & ~n53937;
  assign n53939 = ~n52660 & ~n53938;
  assign n53940 = ~n52689 & ~n53939;
  assign n53941 = ~n52624 & n52643;
  assign n53942 = n52650 & n53941;
  assign n53943 = ~n53851 & ~n53942;
  assign n53944 = ~n52689 & ~n53943;
  assign n53945 = ~n53940 & ~n53944;
  assign n53946 = ~n53933 & n53945;
  assign n53947 = ~n52677 & ~n52696;
  assign n53948 = ~n52706 & n53947;
  assign n53949 = ~n52624 & ~n53948;
  assign n53950 = ~n52650 & n52656;
  assign n53951 = ~n52680 & ~n53950;
  assign n53952 = n52624 & ~n53951;
  assign n53953 = ~n53949 & ~n53952;
  assign n53954 = ~n53866 & n53953;
  assign n53955 = ~n52666 & ~n52707;
  assign n53956 = n53954 & n53955;
  assign n53957 = n52689 & ~n53956;
  assign n53958 = n53946 & ~n53957;
  assign n53959 = n53930 & n53958;
  assign n53960 = ~pi1479 & ~n53959;
  assign n53961 = pi1479 & n53946;
  assign n53962 = n53930 & n53961;
  assign n53963 = ~n53957 & n53962;
  assign po1556 = n53960 | n53963;
  assign n53965 = n52431 & n53157;
  assign n53966 = n52437 & n53965;
  assign n53967 = n52477 & ~n53610;
  assign n53968 = ~n52495 & ~n53967;
  assign n53969 = ~n53153 & n53968;
  assign n53970 = ~n52437 & ~n53969;
  assign n53971 = n52431 & n52447;
  assign n53972 = ~n53970 & ~n53971;
  assign n53973 = n52445 & n52494;
  assign n53974 = ~n52431 & n53161;
  assign n53975 = ~n53973 & ~n53974;
  assign n53976 = ~n53613 & n53975;
  assign n53977 = n52437 & ~n53976;
  assign n53978 = n53972 & ~n53977;
  assign n53979 = n52412 & ~n53978;
  assign n53980 = ~n53966 & ~n53979;
  assign n53981 = ~n52431 & n52446;
  assign n53982 = ~n53152 & ~n53981;
  assign n53983 = n52437 & ~n53982;
  assign n53984 = ~n52496 & ~n53983;
  assign n53985 = ~n52467 & ~n53965;
  assign n53986 = n52431 & n52501;
  assign n53987 = ~n53161 & ~n53986;
  assign n53988 = ~n53973 & n53987;
  assign n53989 = ~n52437 & ~n53988;
  assign n53990 = ~n52431 & n52447;
  assign n53991 = ~n53989 & ~n53990;
  assign n53992 = n53985 & n53991;
  assign n53993 = n53984 & n53992;
  assign n53994 = ~n52412 & ~n53993;
  assign n53995 = ~n52482 & ~n53615;
  assign n53996 = ~n52437 & ~n53995;
  assign n53997 = ~n53994 & ~n53996;
  assign n53998 = n53980 & n53997;
  assign n53999 = pi1460 & n53998;
  assign n54000 = ~pi1460 & ~n53998;
  assign po1557 = n53999 | n54000;
  assign n54002 = ~n53449 & n53462;
  assign n54003 = ~n53667 & ~n54002;
  assign n54004 = ~n53481 & ~n54003;
  assign n54005 = ~n53472 & n53490;
  assign n54006 = ~n53463 & ~n54005;
  assign n54007 = ~n53522 & n54006;
  assign n54008 = n53481 & ~n54007;
  assign n54009 = ~n54004 & ~n54008;
  assign n54010 = ~n53495 & ~n53506;
  assign n54011 = n54009 & n54010;
  assign n54012 = ~n53487 & ~n54011;
  assign n54013 = n53472 & n53667;
  assign n54014 = n53464 & ~n53472;
  assign n54015 = ~n53657 & ~n54014;
  assign n54016 = n53481 & ~n54015;
  assign n54017 = ~n54013 & ~n54016;
  assign n54018 = n53449 & ~n53481;
  assign n54019 = ~n53455 & n54018;
  assign n54020 = n53461 & n54019;
  assign n54021 = n53466 & ~n54020;
  assign n54022 = ~n53522 & n54021;
  assign n54023 = ~n53472 & ~n54022;
  assign n54024 = n54017 & ~n54023;
  assign n54025 = n53487 & ~n54024;
  assign n54026 = ~n54012 & ~n54025;
  assign n54027 = ~n53449 & n53657;
  assign n54028 = ~n53520 & ~n54027;
  assign n54029 = ~n53481 & ~n54028;
  assign n54030 = ~n53449 & ~n53461;
  assign n54031 = n53512 & n54030;
  assign n54032 = ~n54029 & ~n54031;
  assign n54033 = n54026 & n54032;
  assign n54034 = ~pi1453 & ~n54033;
  assign n54035 = pi1453 & ~n54029;
  assign n54036 = n54026 & n54035;
  assign n54037 = ~n54031 & n54036;
  assign po1558 = n54034 | n54037;
  assign n54039 = n53462 & n53507;
  assign n54040 = ~n53481 & n54039;
  assign n54041 = n53449 & ~n53455;
  assign n54042 = n53512 & n54041;
  assign n54043 = ~n54040 & ~n54042;
  assign n54044 = ~n53657 & ~n53659;
  assign n54045 = ~n53481 & ~n54044;
  assign n54046 = ~n53671 & ~n54045;
  assign n54047 = n53487 & ~n54046;
  assign n54048 = n53472 & n53522;
  assign n54049 = ~n53455 & n53473;
  assign n54050 = ~n53462 & ~n54030;
  assign n54051 = n53472 & ~n54050;
  assign n54052 = ~n54049 & ~n54051;
  assign n54053 = ~n53481 & ~n54052;
  assign n54054 = ~n54048 & ~n54053;
  assign n54055 = ~n53472 & ~n54050;
  assign n54056 = ~n53667 & ~n54055;
  assign n54057 = n53481 & ~n54056;
  assign n54058 = ~n53651 & ~n54057;
  assign n54059 = n54054 & n54058;
  assign n54060 = ~n53487 & ~n54059;
  assign n54061 = n53449 & n53472;
  assign n54062 = ~n53462 & n54061;
  assign n54063 = n53487 & n54062;
  assign n54064 = ~n53491 & ~n53655;
  assign n54065 = n53488 & ~n54064;
  assign n54066 = ~n54063 & ~n54065;
  assign n54067 = ~n54060 & n54066;
  assign n54068 = ~n54047 & n54067;
  assign n54069 = n54043 & n54068;
  assign n54070 = ~pi1455 & n54069;
  assign n54071 = pi1455 & ~n54069;
  assign po1559 = n54070 | n54071;
  assign n54073 = ~n53352 & ~n53755;
  assign n54074 = ~n53735 & n54073;
  assign n54075 = ~n53320 & ~n54074;
  assign n54076 = ~n53363 & ~n53390;
  assign n54077 = ~n53360 & ~n53743;
  assign n54078 = ~n53342 & ~n53748;
  assign n54079 = n53320 & ~n54078;
  assign n54080 = ~n53417 & ~n54079;
  assign n54081 = n54077 & n54080;
  assign n54082 = n53308 & ~n54081;
  assign n54083 = ~n53334 & n53340;
  assign n54084 = ~n53402 & ~n54083;
  assign n54085 = n53314 & ~n54084;
  assign n54086 = ~n53369 & ~n53373;
  assign n54087 = n53320 & ~n54086;
  assign n54088 = n53314 & n53340;
  assign n54089 = ~n53349 & ~n54088;
  assign n54090 = ~n53341 & n54089;
  assign n54091 = ~n53320 & ~n54090;
  assign n54092 = ~n54087 & ~n54091;
  assign n54093 = ~n54085 & n54092;
  assign n54094 = ~n53308 & ~n54093;
  assign n54095 = ~n54082 & ~n54094;
  assign n54096 = n54076 & n54095;
  assign n54097 = ~n54075 & n54096;
  assign n54098 = ~pi1474 & ~n54097;
  assign n54099 = pi1474 & n54076;
  assign n54100 = ~n54075 & n54099;
  assign n54101 = n54095 & n54100;
  assign po1560 = n54098 | n54101;
  assign n54103 = n52974 & n53015;
  assign n54104 = ~n53029 & ~n54103;
  assign n54105 = ~n53003 & ~n54104;
  assign n54106 = n53003 & ~n53249;
  assign n54107 = ~n54105 & ~n54106;
  assign n54108 = ~n53215 & n54107;
  assign n54109 = n53009 & ~n54108;
  assign n54110 = n52996 & ~n53003;
  assign n54111 = ~n54109 & ~n54110;
  assign n54112 = ~n53895 & ~n53909;
  assign n54113 = n53003 & ~n54112;
  assign n54114 = ~n52994 & n53224;
  assign n54115 = ~n53235 & ~n54114;
  assign n54116 = ~n52980 & ~n54115;
  assign n54117 = n53003 & n53030;
  assign n54118 = ~n52974 & n53016;
  assign n54119 = ~n54117 & ~n54118;
  assign n54120 = ~n53014 & n54119;
  assign n54121 = ~n53236 & n54120;
  assign n54122 = ~n54116 & n54121;
  assign n54123 = ~n53009 & ~n54122;
  assign n54124 = ~n54113 & ~n54123;
  assign n54125 = n54111 & n54124;
  assign n54126 = pi1498 & n54125;
  assign n54127 = ~pi1498 & ~n54125;
  assign po1561 = n54126 | n54127;
  assign n54129 = pi4836 & ~pi9040;
  assign n54130 = pi4832 & pi9040;
  assign n54131 = ~n54129 & ~n54130;
  assign n54132 = ~pi1484 & ~n54131;
  assign n54133 = pi1484 & n54131;
  assign n54134 = ~n54132 & ~n54133;
  assign n54135 = pi4845 & pi9040;
  assign n54136 = pi5150 & ~pi9040;
  assign n54137 = ~n54135 & ~n54136;
  assign n54138 = ~pi1489 & ~n54137;
  assign n54139 = pi1489 & n54137;
  assign n54140 = ~n54138 & ~n54139;
  assign n54141 = pi4841 & pi9040;
  assign n54142 = pi4821 & ~pi9040;
  assign n54143 = ~n54141 & ~n54142;
  assign n54144 = ~pi1463 & ~n54143;
  assign n54145 = pi1463 & n54143;
  assign n54146 = ~n54144 & ~n54145;
  assign n54147 = pi5184 & ~pi9040;
  assign n54148 = pi4874 & pi9040;
  assign n54149 = ~n54147 & ~n54148;
  assign n54150 = ~pi1493 & n54149;
  assign n54151 = pi1493 & ~n54149;
  assign n54152 = ~n54150 & ~n54151;
  assign n54153 = pi5187 & pi9040;
  assign n54154 = pi4843 & ~pi9040;
  assign n54155 = ~n54153 & ~n54154;
  assign n54156 = ~pi1476 & n54155;
  assign n54157 = pi1476 & ~n54155;
  assign n54158 = ~n54156 & ~n54157;
  assign n54159 = ~n54152 & n54158;
  assign n54160 = n54146 & n54159;
  assign n54161 = pi4967 & ~pi9040;
  assign n54162 = pi4906 & pi9040;
  assign n54163 = ~n54161 & ~n54162;
  assign n54164 = ~pi1469 & n54163;
  assign n54165 = pi1469 & ~n54163;
  assign n54166 = ~n54164 & ~n54165;
  assign n54167 = ~n54158 & ~n54166;
  assign n54168 = ~n54152 & n54167;
  assign n54169 = ~n54160 & ~n54168;
  assign n54170 = ~n54158 & n54166;
  assign n54171 = n54152 & n54170;
  assign n54172 = ~n54146 & n54171;
  assign n54173 = n54169 & ~n54172;
  assign n54174 = n54140 & ~n54173;
  assign n54175 = n54152 & ~n54158;
  assign n54176 = ~n54146 & ~n54166;
  assign n54177 = n54175 & n54176;
  assign n54178 = n54158 & ~n54166;
  assign n54179 = ~n54152 & n54178;
  assign n54180 = ~n54146 & n54179;
  assign n54181 = n54152 & n54158;
  assign n54182 = ~n54170 & ~n54181;
  assign n54183 = n54146 & ~n54182;
  assign n54184 = ~n54180 & ~n54183;
  assign n54185 = ~n54177 & n54184;
  assign n54186 = ~n54140 & ~n54185;
  assign n54187 = ~n54174 & ~n54186;
  assign n54188 = n54134 & ~n54187;
  assign n54189 = n54158 & n54166;
  assign n54190 = n54152 & n54189;
  assign n54191 = ~n54140 & n54190;
  assign n54192 = ~n54146 & n54191;
  assign n54193 = ~n54152 & n54170;
  assign n54194 = ~n54146 & n54193;
  assign n54195 = ~n54140 & n54194;
  assign n54196 = ~n54192 & ~n54195;
  assign n54197 = ~n54146 & n54152;
  assign n54198 = ~n54166 & n54197;
  assign n54199 = n54158 & n54198;
  assign n54200 = n54140 & n54199;
  assign n54201 = n54196 & ~n54200;
  assign n54202 = n54140 & ~n54146;
  assign n54203 = n54158 & n54202;
  assign n54204 = ~n54140 & ~n54146;
  assign n54205 = n54170 & n54204;
  assign n54206 = ~n54146 & ~n54158;
  assign n54207 = ~n54152 & n54206;
  assign n54208 = ~n54160 & ~n54207;
  assign n54209 = ~n54140 & ~n54208;
  assign n54210 = ~n54205 & ~n54209;
  assign n54211 = ~n54166 & n54175;
  assign n54212 = n54146 & n54211;
  assign n54213 = ~n54194 & ~n54212;
  assign n54214 = n54140 & n54146;
  assign n54215 = n54175 & n54214;
  assign n54216 = n54152 & n54178;
  assign n54217 = n54140 & n54216;
  assign n54218 = ~n54215 & ~n54217;
  assign n54219 = n54213 & n54218;
  assign n54220 = n54210 & n54219;
  assign n54221 = ~n54203 & n54220;
  assign n54222 = ~n54134 & ~n54221;
  assign n54223 = ~n54146 & ~n54152;
  assign n54224 = n54166 & n54223;
  assign n54225 = n54158 & n54224;
  assign n54226 = n54146 & n54167;
  assign n54227 = ~n54225 & ~n54226;
  assign n54228 = n54140 & ~n54227;
  assign n54229 = ~n54222 & ~n54228;
  assign n54230 = n54201 & n54229;
  assign n54231 = ~n54188 & n54230;
  assign n54232 = ~pi1504 & ~n54231;
  assign n54233 = pi1504 & n54231;
  assign po1581 = n54232 | n54233;
  assign n54235 = pi4965 & pi9040;
  assign n54236 = pi4876 & ~pi9040;
  assign n54237 = ~n54235 & ~n54236;
  assign n54238 = ~pi1480 & ~n54237;
  assign n54239 = pi1480 & n54237;
  assign n54240 = ~n54238 & ~n54239;
  assign n54241 = pi4987 & pi9040;
  assign n54242 = pi4842 & ~pi9040;
  assign n54243 = ~n54241 & ~n54242;
  assign n54244 = ~pi1484 & n54243;
  assign n54245 = pi1484 & ~n54243;
  assign n54246 = ~n54244 & ~n54245;
  assign n54247 = pi4876 & pi9040;
  assign n54248 = pi4987 & ~pi9040;
  assign n54249 = ~n54247 & ~n54248;
  assign n54250 = pi1481 & n54249;
  assign n54251 = ~pi1481 & ~n54249;
  assign n54252 = ~n54250 & ~n54251;
  assign n54253 = n54246 & n54252;
  assign n54254 = pi5187 & ~pi9040;
  assign n54255 = pi4967 & pi9040;
  assign n54256 = ~n54254 & ~n54255;
  assign n54257 = ~pi1470 & ~n54256;
  assign n54258 = pi1470 & n54256;
  assign n54259 = ~n54257 & ~n54258;
  assign n54260 = pi4890 & ~pi9040;
  assign n54261 = pi4964 & pi9040;
  assign n54262 = ~n54260 & ~n54261;
  assign n54263 = pi1496 & n54262;
  assign n54264 = ~pi1496 & ~n54262;
  assign n54265 = ~n54263 & ~n54264;
  assign n54266 = ~n54259 & ~n54265;
  assign n54267 = n54253 & n54266;
  assign n54268 = pi4843 & pi9040;
  assign n54269 = pi4874 & ~pi9040;
  assign n54270 = ~n54268 & ~n54269;
  assign n54271 = ~pi1469 & n54270;
  assign n54272 = pi1469 & ~n54270;
  assign n54273 = ~n54271 & ~n54272;
  assign n54274 = ~n54246 & ~n54252;
  assign n54275 = ~n54273 & n54274;
  assign n54276 = n54259 & n54273;
  assign n54277 = ~n54252 & n54276;
  assign n54278 = n54246 & n54277;
  assign n54279 = ~n54275 & ~n54278;
  assign n54280 = ~n54246 & n54252;
  assign n54281 = n54259 & n54280;
  assign n54282 = n54279 & ~n54281;
  assign n54283 = ~n54265 & ~n54282;
  assign n54284 = ~n54246 & n54273;
  assign n54285 = ~n54259 & n54265;
  assign n54286 = n54284 & n54285;
  assign n54287 = n54273 & n54274;
  assign n54288 = ~n54259 & n54287;
  assign n54289 = ~n54286 & ~n54288;
  assign n54290 = ~n54283 & n54289;
  assign n54291 = ~n54267 & n54290;
  assign n54292 = n54253 & ~n54273;
  assign n54293 = ~n54259 & n54292;
  assign n54294 = ~n54273 & n54280;
  assign n54295 = n54259 & n54294;
  assign n54296 = ~n54293 & ~n54295;
  assign n54297 = n54291 & n54296;
  assign n54298 = ~n54240 & ~n54297;
  assign n54299 = ~n54259 & n54273;
  assign n54300 = n54252 & n54299;
  assign n54301 = ~n54246 & n54300;
  assign n54302 = ~n54292 & ~n54301;
  assign n54303 = ~n54265 & ~n54302;
  assign n54304 = n54253 & n54276;
  assign n54305 = ~n54252 & n54299;
  assign n54306 = n54246 & n54305;
  assign n54307 = ~n54304 & ~n54306;
  assign n54308 = ~n54246 & n54276;
  assign n54309 = ~n54259 & n54294;
  assign n54310 = ~n54308 & ~n54309;
  assign n54311 = n54265 & ~n54310;
  assign n54312 = n54307 & ~n54311;
  assign n54313 = ~n54303 & n54312;
  assign n54314 = n54240 & ~n54313;
  assign n54315 = ~n54246 & ~n54273;
  assign n54316 = n54259 & n54315;
  assign n54317 = n54246 & ~n54273;
  assign n54318 = ~n54259 & n54317;
  assign n54319 = ~n54316 & ~n54318;
  assign n54320 = ~n54265 & ~n54319;
  assign n54321 = n54246 & ~n54252;
  assign n54322 = ~n54273 & n54321;
  assign n54323 = n54259 & n54322;
  assign n54324 = ~n54304 & ~n54323;
  assign n54325 = ~n54287 & n54324;
  assign n54326 = n54265 & ~n54325;
  assign n54327 = ~n54320 & ~n54326;
  assign n54328 = ~n54252 & n54273;
  assign n54329 = n54265 & n54328;
  assign n54330 = ~n54259 & n54329;
  assign n54331 = n54327 & ~n54330;
  assign n54332 = ~n54314 & n54331;
  assign n54333 = ~n54298 & n54332;
  assign n54334 = ~pi1509 & ~n54333;
  assign n54335 = pi1509 & n54333;
  assign po1586 = n54334 | n54335;
  assign n54337 = ~n54134 & ~n54140;
  assign n54338 = ~n54146 & n54159;
  assign n54339 = n54146 & n54193;
  assign n54340 = ~n54146 & n54167;
  assign n54341 = ~n54339 & ~n54340;
  assign n54342 = ~n54338 & n54341;
  assign n54343 = n54337 & ~n54342;
  assign n54344 = ~n54168 & ~n54171;
  assign n54345 = n54166 & n54197;
  assign n54346 = ~n54152 & n54189;
  assign n54347 = n54146 & n54346;
  assign n54348 = ~n54345 & ~n54347;
  assign n54349 = n54344 & n54348;
  assign n54350 = n54140 & ~n54349;
  assign n54351 = n54146 & n54216;
  assign n54352 = ~n54350 & ~n54351;
  assign n54353 = ~n54134 & ~n54352;
  assign n54354 = ~n54343 & ~n54353;
  assign n54355 = ~n54152 & n54202;
  assign n54356 = ~n54166 & n54355;
  assign n54357 = ~n54172 & ~n54356;
  assign n54358 = ~n54167 & ~n54189;
  assign n54359 = n54146 & ~n54358;
  assign n54360 = ~n54190 & ~n54359;
  assign n54361 = ~n54140 & ~n54360;
  assign n54362 = ~n54179 & ~n54338;
  assign n54363 = ~n54339 & n54362;
  assign n54364 = n54140 & ~n54363;
  assign n54365 = ~n54361 & ~n54364;
  assign n54366 = n54146 & n54190;
  assign n54367 = ~n54212 & ~n54366;
  assign n54368 = ~n54199 & n54367;
  assign n54369 = ~n54205 & n54368;
  assign n54370 = n54365 & n54369;
  assign n54371 = n54134 & ~n54370;
  assign n54372 = n54357 & ~n54371;
  assign n54373 = n54354 & n54372;
  assign n54374 = pi1505 & ~n54373;
  assign n54375 = ~pi1505 & n54357;
  assign n54376 = n54354 & n54375;
  assign n54377 = ~n54371 & n54376;
  assign po1590 = n54374 | n54377;
  assign n54379 = ~n54179 & ~n54190;
  assign n54380 = ~n54140 & ~n54379;
  assign n54381 = n54146 & n54168;
  assign n54382 = ~n54380 & ~n54381;
  assign n54383 = n54146 & ~n54158;
  assign n54384 = ~n54175 & ~n54383;
  assign n54385 = ~n54346 & n54384;
  assign n54386 = n54140 & ~n54385;
  assign n54387 = n54382 & ~n54386;
  assign n54388 = ~n54134 & ~n54387;
  assign n54389 = ~n54146 & n54211;
  assign n54390 = ~n54140 & n54389;
  assign n54391 = ~n54195 & ~n54390;
  assign n54392 = ~n54200 & n54391;
  assign n54393 = n54140 & n54207;
  assign n54394 = n54146 & n54179;
  assign n54395 = ~n54140 & n54175;
  assign n54396 = ~n54394 & ~n54395;
  assign n54397 = ~n54366 & n54396;
  assign n54398 = ~n54393 & n54397;
  assign n54399 = ~n54199 & ~n54224;
  assign n54400 = n54398 & n54399;
  assign n54401 = ~n54217 & n54400;
  assign n54402 = n54134 & ~n54401;
  assign n54403 = n54392 & ~n54402;
  assign n54404 = ~n54388 & n54403;
  assign n54405 = ~pi1511 & ~n54404;
  assign n54406 = pi1511 & n54392;
  assign n54407 = ~n54388 & n54406;
  assign n54408 = ~n54402 & n54407;
  assign po1591 = n54405 | n54408;
  assign n54410 = pi4890 & pi9040;
  assign n54411 = pi4960 & ~pi9040;
  assign n54412 = ~n54410 & ~n54411;
  assign n54413 = pi1476 & n54412;
  assign n54414 = ~pi1476 & ~n54412;
  assign n54415 = ~n54413 & ~n54414;
  assign n54416 = pi5184 & pi9040;
  assign n54417 = pi4818 & ~pi9040;
  assign n54418 = ~n54416 & ~n54417;
  assign n54419 = pi1503 & n54418;
  assign n54420 = ~pi1503 & ~n54418;
  assign n54421 = ~n54419 & ~n54420;
  assign n54422 = pi4957 & ~pi9040;
  assign n54423 = pi4911 & pi9040;
  assign n54424 = ~n54422 & ~n54423;
  assign n54425 = ~pi1483 & n54424;
  assign n54426 = pi1483 & ~n54424;
  assign n54427 = ~n54425 & ~n54426;
  assign n54428 = pi4836 & pi9040;
  assign n54429 = pi4988 & ~pi9040;
  assign n54430 = ~n54428 & ~n54429;
  assign n54431 = pi1478 & n54430;
  assign n54432 = ~pi1478 & ~n54430;
  assign n54433 = ~n54431 & ~n54432;
  assign n54434 = pi4881 & pi9040;
  assign n54435 = pi5038 & ~pi9040;
  assign n54436 = ~n54434 & ~n54435;
  assign n54437 = ~pi1493 & ~n54436;
  assign n54438 = pi1493 & n54436;
  assign n54439 = ~n54437 & ~n54438;
  assign n54440 = n54433 & ~n54439;
  assign n54441 = ~n54427 & n54440;
  assign n54442 = n54421 & n54441;
  assign n54443 = ~n54421 & n54433;
  assign n54444 = n54439 & n54443;
  assign n54445 = pi4990 & pi9040;
  assign n54446 = pi4964 & ~pi9040;
  assign n54447 = ~n54445 & ~n54446;
  assign n54448 = ~pi1495 & n54447;
  assign n54449 = pi1495 & ~n54447;
  assign n54450 = ~n54448 & ~n54449;
  assign n54451 = n54427 & n54443;
  assign n54452 = ~n54427 & n54439;
  assign n54453 = ~n54433 & n54452;
  assign n54454 = ~n54451 & ~n54453;
  assign n54455 = n54450 & ~n54454;
  assign n54456 = ~n54444 & ~n54455;
  assign n54457 = n54433 & n54452;
  assign n54458 = n54427 & ~n54433;
  assign n54459 = ~n54433 & ~n54439;
  assign n54460 = ~n54421 & n54459;
  assign n54461 = n54427 & ~n54439;
  assign n54462 = n54421 & n54461;
  assign n54463 = ~n54460 & ~n54462;
  assign n54464 = ~n54458 & n54463;
  assign n54465 = ~n54457 & n54464;
  assign n54466 = ~n54450 & ~n54465;
  assign n54467 = n54456 & ~n54466;
  assign n54468 = ~n54442 & n54467;
  assign n54469 = n54415 & ~n54468;
  assign n54470 = n54427 & n54439;
  assign n54471 = ~n54433 & n54470;
  assign n54472 = ~n54421 & n54471;
  assign n54473 = n54421 & ~n54433;
  assign n54474 = ~n54439 & n54473;
  assign n54475 = n54427 & n54474;
  assign n54476 = ~n54442 & ~n54475;
  assign n54477 = ~n54472 & n54476;
  assign n54478 = ~n54450 & ~n54477;
  assign n54479 = ~n54469 & ~n54478;
  assign n54480 = ~n54427 & n54444;
  assign n54481 = n54450 & n54473;
  assign n54482 = ~n54427 & n54481;
  assign n54483 = n54433 & n54470;
  assign n54484 = n54421 & n54483;
  assign n54485 = n54440 & ~n54450;
  assign n54486 = ~n54421 & n54485;
  assign n54487 = ~n54484 & ~n54486;
  assign n54488 = n54427 & n54433;
  assign n54489 = n54421 & n54488;
  assign n54490 = ~n54427 & ~n54439;
  assign n54491 = ~n54433 & n54490;
  assign n54492 = ~n54489 & ~n54491;
  assign n54493 = n54450 & ~n54492;
  assign n54494 = n54450 & n54458;
  assign n54495 = ~n54421 & n54494;
  assign n54496 = ~n54493 & ~n54495;
  assign n54497 = n54487 & n54496;
  assign n54498 = ~n54415 & ~n54497;
  assign n54499 = ~n54482 & ~n54498;
  assign n54500 = ~n54480 & n54499;
  assign n54501 = n54479 & n54500;
  assign n54502 = ~pi1512 & ~n54501;
  assign n54503 = ~n54469 & ~n54480;
  assign n54504 = ~n54478 & n54503;
  assign n54505 = n54499 & n54504;
  assign n54506 = pi1512 & n54505;
  assign po1592 = n54502 | n54506;
  assign n54508 = pi4962 & pi9040;
  assign n54509 = pi4844 & ~pi9040;
  assign n54510 = ~n54508 & ~n54509;
  assign n54511 = ~pi1494 & ~n54510;
  assign n54512 = pi1494 & n54510;
  assign n54513 = ~n54511 & ~n54512;
  assign n54514 = pi5039 & pi9040;
  assign n54515 = pi4961 & ~pi9040;
  assign n54516 = ~n54514 & ~n54515;
  assign n54517 = ~pi1487 & ~n54516;
  assign n54518 = pi1487 & n54516;
  assign n54519 = ~n54517 & ~n54518;
  assign n54520 = pi5063 & ~pi9040;
  assign n54521 = pi4833 & pi9040;
  assign n54522 = ~n54520 & ~n54521;
  assign n54523 = ~pi1497 & ~n54522;
  assign n54524 = pi1497 & n54522;
  assign n54525 = ~n54523 & ~n54524;
  assign n54526 = pi5063 & pi9040;
  assign n54527 = pi4854 & ~pi9040;
  assign n54528 = ~n54526 & ~n54527;
  assign n54529 = ~pi1467 & n54528;
  assign n54530 = pi1467 & ~n54528;
  assign n54531 = ~n54529 & ~n54530;
  assign n54532 = ~n54525 & ~n54531;
  assign n54533 = pi4898 & ~pi9040;
  assign n54534 = pi5278 & pi9040;
  assign n54535 = ~n54533 & ~n54534;
  assign n54536 = pi1488 & n54535;
  assign n54537 = ~pi1488 & ~n54535;
  assign n54538 = ~n54536 & ~n54537;
  assign n54539 = pi4854 & pi9040;
  assign n54540 = pi4840 & ~pi9040;
  assign n54541 = ~n54539 & ~n54540;
  assign n54542 = ~pi1501 & ~n54541;
  assign n54543 = pi1501 & n54541;
  assign n54544 = ~n54542 & ~n54543;
  assign n54545 = n54538 & n54544;
  assign n54546 = n54532 & n54545;
  assign n54547 = n54519 & n54546;
  assign n54548 = ~n54538 & n54544;
  assign n54549 = n54525 & ~n54531;
  assign n54550 = n54548 & n54549;
  assign n54551 = n54525 & n54531;
  assign n54552 = n54519 & n54551;
  assign n54553 = n54544 & n54552;
  assign n54554 = n54538 & n54553;
  assign n54555 = n54519 & ~n54538;
  assign n54556 = n54531 & n54555;
  assign n54557 = ~n54525 & n54556;
  assign n54558 = ~n54554 & ~n54557;
  assign n54559 = ~n54550 & n54558;
  assign n54560 = ~n54547 & n54559;
  assign n54561 = ~n54519 & ~n54538;
  assign n54562 = ~n54531 & n54561;
  assign n54563 = n54525 & n54562;
  assign n54564 = n54560 & ~n54563;
  assign n54565 = ~n54513 & ~n54564;
  assign n54566 = n54519 & n54525;
  assign n54567 = ~n54531 & n54566;
  assign n54568 = n54538 & n54567;
  assign n54569 = ~n54556 & ~n54568;
  assign n54570 = ~n54519 & n54532;
  assign n54571 = n54538 & n54570;
  assign n54572 = n54569 & ~n54571;
  assign n54573 = ~n54544 & ~n54572;
  assign n54574 = ~n54519 & n54531;
  assign n54575 = n54525 & n54574;
  assign n54576 = ~n54544 & n54575;
  assign n54577 = n54538 & n54576;
  assign n54578 = ~n54525 & n54555;
  assign n54579 = ~n54525 & n54531;
  assign n54580 = ~n54538 & n54579;
  assign n54581 = ~n54578 & ~n54580;
  assign n54582 = ~n54544 & ~n54581;
  assign n54583 = ~n54577 & ~n54582;
  assign n54584 = ~n54513 & ~n54583;
  assign n54585 = ~n54573 & ~n54584;
  assign n54586 = ~n54565 & n54585;
  assign n54587 = ~n54519 & n54538;
  assign n54588 = n54544 & n54587;
  assign n54589 = n54579 & n54588;
  assign n54590 = ~n54519 & n54525;
  assign n54591 = n54548 & n54590;
  assign n54592 = n54519 & ~n54544;
  assign n54593 = n54525 & n54592;
  assign n54594 = ~n54525 & n54538;
  assign n54595 = ~n54519 & n54594;
  assign n54596 = ~n54593 & ~n54595;
  assign n54597 = ~n54538 & n54575;
  assign n54598 = n54596 & ~n54597;
  assign n54599 = ~n54570 & n54598;
  assign n54600 = n54532 & n54544;
  assign n54601 = ~n54538 & n54600;
  assign n54602 = n54538 & n54579;
  assign n54603 = ~n54519 & ~n54531;
  assign n54604 = ~n54602 & ~n54603;
  assign n54605 = n54544 & ~n54604;
  assign n54606 = ~n54601 & ~n54605;
  assign n54607 = n54599 & n54606;
  assign n54608 = n54513 & ~n54607;
  assign n54609 = ~n54591 & ~n54608;
  assign n54610 = ~n54589 & n54609;
  assign n54611 = n54586 & n54610;
  assign n54612 = pi1508 & n54611;
  assign n54613 = ~pi1508 & ~n54611;
  assign po1596 = n54612 | n54613;
  assign n54615 = pi4844 & pi9040;
  assign n54616 = pi5278 & ~pi9040;
  assign n54617 = ~n54615 & ~n54616;
  assign n54618 = ~pi1502 & n54617;
  assign n54619 = pi1502 & ~n54617;
  assign n54620 = ~n54618 & ~n54619;
  assign n54621 = pi4847 & ~pi9040;
  assign n54622 = pi4835 & pi9040;
  assign n54623 = ~n54621 & ~n54622;
  assign n54624 = ~pi1486 & n54623;
  assign n54625 = pi1486 & ~n54623;
  assign n54626 = ~n54624 & ~n54625;
  assign n54627 = pi4909 & ~pi9040;
  assign n54628 = pi5060 & pi9040;
  assign n54629 = ~n54627 & ~n54628;
  assign n54630 = pi1500 & n54629;
  assign n54631 = ~pi1500 & ~n54629;
  assign n54632 = ~n54630 & ~n54631;
  assign n54633 = pi4898 & pi9040;
  assign n54634 = pi5116 & ~pi9040;
  assign n54635 = ~n54633 & ~n54634;
  assign n54636 = ~pi1478 & n54635;
  assign n54637 = pi1478 & ~n54635;
  assign n54638 = ~n54636 & ~n54637;
  assign n54639 = pi4849 & pi9040;
  assign n54640 = pi5060 & ~pi9040;
  assign n54641 = ~n54639 & ~n54640;
  assign n54642 = pi1473 & n54641;
  assign n54643 = ~pi1473 & ~n54641;
  assign n54644 = ~n54642 & ~n54643;
  assign n54645 = n54638 & ~n54644;
  assign n54646 = ~n54632 & n54645;
  assign n54647 = n54626 & n54646;
  assign n54648 = ~pi1473 & n54641;
  assign n54649 = pi1473 & ~n54641;
  assign n54650 = ~n54648 & ~n54649;
  assign n54651 = ~n54626 & ~n54632;
  assign n54652 = n54638 & n54651;
  assign n54653 = ~n54650 & n54652;
  assign n54654 = ~n54647 & ~n54653;
  assign n54655 = ~n54620 & ~n54654;
  assign n54656 = n54626 & n54632;
  assign n54657 = ~n54638 & n54656;
  assign n54658 = ~n54644 & n54657;
  assign n54659 = n54620 & n54658;
  assign n54660 = pi4966 & pi9040;
  assign n54661 = pi4837 & ~pi9040;
  assign n54662 = ~n54660 & ~n54661;
  assign n54663 = ~pi1483 & ~n54662;
  assign n54664 = pi1483 & n54662;
  assign n54665 = ~n54663 & ~n54664;
  assign n54666 = n54638 & ~n54650;
  assign n54667 = n54632 & n54666;
  assign n54668 = ~n54620 & n54667;
  assign n54669 = ~n54658 & ~n54668;
  assign n54670 = n54626 & ~n54650;
  assign n54671 = ~n54632 & n54670;
  assign n54672 = ~n54644 & n54656;
  assign n54673 = ~n54671 & ~n54672;
  assign n54674 = n54620 & ~n54673;
  assign n54675 = n54620 & ~n54626;
  assign n54676 = n54645 & n54675;
  assign n54677 = ~n54632 & n54676;
  assign n54678 = ~n54626 & n54632;
  assign n54679 = ~n54638 & n54678;
  assign n54680 = ~n54650 & n54679;
  assign n54681 = ~n54620 & ~n54632;
  assign n54682 = ~n54638 & n54681;
  assign n54683 = ~n54644 & n54682;
  assign n54684 = ~n54680 & ~n54683;
  assign n54685 = ~n54677 & n54684;
  assign n54686 = ~n54674 & n54685;
  assign n54687 = n54669 & n54686;
  assign n54688 = n54665 & ~n54687;
  assign n54689 = n54626 & n54668;
  assign n54690 = ~n54688 & ~n54689;
  assign n54691 = ~n54659 & n54690;
  assign n54692 = ~n54655 & n54691;
  assign n54693 = ~n54620 & ~n54626;
  assign n54694 = n54632 & ~n54644;
  assign n54695 = n54693 & n54694;
  assign n54696 = ~n54620 & n54646;
  assign n54697 = ~n54695 & ~n54696;
  assign n54698 = ~n54638 & ~n54650;
  assign n54699 = n54632 & n54698;
  assign n54700 = ~n54620 & n54699;
  assign n54701 = ~n54632 & n54698;
  assign n54702 = n54626 & n54701;
  assign n54703 = ~n54700 & ~n54702;
  assign n54704 = n54632 & n54645;
  assign n54705 = ~n54626 & n54704;
  assign n54706 = ~n54647 & ~n54705;
  assign n54707 = ~n54626 & n54666;
  assign n54708 = ~n54632 & ~n54638;
  assign n54709 = ~n54707 & ~n54708;
  assign n54710 = n54620 & ~n54709;
  assign n54711 = n54706 & ~n54710;
  assign n54712 = n54703 & n54711;
  assign n54713 = n54697 & n54712;
  assign n54714 = ~n54665 & ~n54713;
  assign n54715 = n54692 & ~n54714;
  assign n54716 = ~pi1514 & ~n54715;
  assign n54717 = pi1514 & n54692;
  assign n54718 = ~n54714 & n54717;
  assign po1597 = n54716 | n54718;
  assign n54720 = n54140 & n54167;
  assign n54721 = ~n54146 & n54720;
  assign n54722 = ~n54225 & ~n54721;
  assign n54723 = n54146 & ~n54166;
  assign n54724 = ~n54152 & n54723;
  assign n54725 = ~n54146 & n54158;
  assign n54726 = ~n54224 & ~n54725;
  assign n54727 = ~n54140 & ~n54726;
  assign n54728 = ~n54724 & ~n54727;
  assign n54729 = n54722 & n54728;
  assign n54730 = n54134 & ~n54729;
  assign n54731 = ~n54193 & ~n54212;
  assign n54732 = ~n54146 & n54178;
  assign n54733 = n54731 & ~n54732;
  assign n54734 = n54140 & ~n54733;
  assign n54735 = n54167 & n54204;
  assign n54736 = ~n54172 & ~n54735;
  assign n54737 = ~n54734 & n54736;
  assign n54738 = ~n54346 & ~n54351;
  assign n54739 = ~n54140 & ~n54738;
  assign n54740 = n54737 & ~n54739;
  assign n54741 = ~n54134 & ~n54740;
  assign n54742 = ~n54730 & ~n54741;
  assign n54743 = ~n54146 & n54189;
  assign n54744 = n54146 & ~n54344;
  assign n54745 = ~n54743 & ~n54744;
  assign n54746 = ~n54140 & ~n54745;
  assign n54747 = ~n54193 & n54379;
  assign n54748 = n54214 & ~n54747;
  assign n54749 = ~n54746 & ~n54748;
  assign n54750 = n54742 & n54749;
  assign n54751 = ~pi1515 & ~n54750;
  assign n54752 = ~n54741 & n54749;
  assign n54753 = pi1515 & n54752;
  assign n54754 = ~n54730 & n54753;
  assign po1598 = n54751 | n54754;
  assign n54756 = pi4881 & ~pi9040;
  assign n54757 = pi5150 & pi9040;
  assign n54758 = ~n54756 & ~n54757;
  assign n54759 = pi1464 & n54758;
  assign n54760 = ~pi1464 & ~n54758;
  assign n54761 = ~n54759 & ~n54760;
  assign n54762 = pi4832 & ~pi9040;
  assign n54763 = pi4821 & pi9040;
  assign n54764 = ~n54762 & ~n54763;
  assign n54765 = ~pi1481 & n54764;
  assign n54766 = pi1481 & ~n54764;
  assign n54767 = ~n54765 & ~n54766;
  assign n54768 = pi4957 & pi9040;
  assign n54769 = pi4841 & ~pi9040;
  assign n54770 = ~n54768 & ~n54769;
  assign n54771 = ~pi1487 & n54770;
  assign n54772 = pi1487 & ~n54770;
  assign n54773 = ~n54771 & ~n54772;
  assign n54774 = pi4990 & ~pi9040;
  assign n54775 = pi5038 & pi9040;
  assign n54776 = ~n54774 & ~n54775;
  assign n54777 = ~pi1480 & n54776;
  assign n54778 = pi1480 & ~n54776;
  assign n54779 = ~n54777 & ~n54778;
  assign n54780 = ~n54773 & ~n54779;
  assign n54781 = n54767 & n54780;
  assign n54782 = pi4818 & pi9040;
  assign n54783 = pi4911 & ~pi9040;
  assign n54784 = ~n54782 & ~n54783;
  assign n54785 = pi1485 & n54784;
  assign n54786 = ~pi1485 & ~n54784;
  assign n54787 = ~n54785 & ~n54786;
  assign n54788 = n54781 & ~n54787;
  assign n54789 = pi1480 & n54776;
  assign n54790 = ~pi1480 & ~n54776;
  assign n54791 = ~n54789 & ~n54790;
  assign n54792 = n54773 & ~n54791;
  assign n54793 = n54767 & n54792;
  assign n54794 = ~n54787 & n54793;
  assign n54795 = ~n54788 & ~n54794;
  assign n54796 = ~n54767 & n54787;
  assign n54797 = n54792 & n54796;
  assign n54798 = ~n54773 & ~n54791;
  assign n54799 = n54767 & n54798;
  assign n54800 = n54787 & n54799;
  assign n54801 = ~n54797 & ~n54800;
  assign n54802 = n54795 & n54801;
  assign n54803 = n54761 & ~n54802;
  assign n54804 = n54767 & n54787;
  assign n54805 = ~n54779 & n54804;
  assign n54806 = n54773 & n54805;
  assign n54807 = ~n54799 & ~n54806;
  assign n54808 = n54761 & ~n54807;
  assign n54809 = ~n54761 & ~n54779;
  assign n54810 = ~n54787 & n54809;
  assign n54811 = ~n54767 & ~n54773;
  assign n54812 = n54787 & n54792;
  assign n54813 = ~n54811 & ~n54812;
  assign n54814 = ~n54761 & ~n54813;
  assign n54815 = ~n54810 & ~n54814;
  assign n54816 = n54773 & ~n54779;
  assign n54817 = ~n54767 & n54816;
  assign n54818 = ~n54787 & n54817;
  assign n54819 = n54815 & ~n54818;
  assign n54820 = ~n54779 & n54811;
  assign n54821 = n54787 & n54820;
  assign n54822 = n54819 & ~n54821;
  assign n54823 = ~n54808 & n54822;
  assign n54824 = pi5185 & pi9040;
  assign n54825 = pi4906 & ~pi9040;
  assign n54826 = ~n54824 & ~n54825;
  assign n54827 = ~pi1497 & ~n54826;
  assign n54828 = pi1497 & n54826;
  assign n54829 = ~n54827 & ~n54828;
  assign n54830 = ~n54823 & ~n54829;
  assign n54831 = n54767 & ~n54779;
  assign n54832 = ~n54761 & n54787;
  assign n54833 = n54829 & n54832;
  assign n54834 = n54831 & n54833;
  assign n54835 = n54767 & ~n54787;
  assign n54836 = ~n54791 & n54835;
  assign n54837 = ~n54761 & ~n54836;
  assign n54838 = n54773 & n54796;
  assign n54839 = ~n54780 & ~n54831;
  assign n54840 = ~n54787 & ~n54839;
  assign n54841 = ~n54767 & n54792;
  assign n54842 = n54761 & ~n54841;
  assign n54843 = ~n54840 & n54842;
  assign n54844 = ~n54838 & n54843;
  assign n54845 = ~n54837 & ~n54844;
  assign n54846 = ~n54767 & n54798;
  assign n54847 = n54787 & n54846;
  assign n54848 = ~n54845 & ~n54847;
  assign n54849 = n54829 & ~n54848;
  assign n54850 = ~n54834 & ~n54849;
  assign n54851 = ~n54830 & n54850;
  assign n54852 = ~n54803 & n54851;
  assign n54853 = ~n54761 & n54818;
  assign n54854 = n54852 & ~n54853;
  assign n54855 = pi1506 & ~n54854;
  assign n54856 = ~pi1506 & ~n54853;
  assign n54857 = n54851 & n54856;
  assign n54858 = ~n54803 & n54857;
  assign po1599 = n54855 | n54858;
  assign n54860 = ~n54638 & ~n54644;
  assign n54861 = n54632 & n54860;
  assign n54862 = ~n54626 & n54861;
  assign n54863 = ~n54626 & n54698;
  assign n54864 = ~n54632 & n54860;
  assign n54865 = n54626 & n54864;
  assign n54866 = ~n54863 & ~n54865;
  assign n54867 = n54620 & ~n54866;
  assign n54868 = ~n54862 & ~n54867;
  assign n54869 = ~n54620 & n54860;
  assign n54870 = ~n54626 & n54869;
  assign n54871 = ~n54696 & ~n54870;
  assign n54872 = n54868 & n54871;
  assign n54873 = ~n54626 & n54667;
  assign n54874 = n54626 & n54704;
  assign n54875 = ~n54873 & ~n54874;
  assign n54876 = n54872 & n54875;
  assign n54877 = n54665 & ~n54876;
  assign n54878 = n54620 & ~n54665;
  assign n54879 = n54650 & n54651;
  assign n54880 = ~n54632 & n54638;
  assign n54881 = ~n54879 & ~n54880;
  assign n54882 = n54878 & ~n54881;
  assign n54883 = ~n54658 & ~n54671;
  assign n54884 = n54632 & n54693;
  assign n54885 = ~n54860 & n54884;
  assign n54886 = ~n54668 & ~n54885;
  assign n54887 = n54883 & n54886;
  assign n54888 = ~n54665 & ~n54887;
  assign n54889 = ~n54632 & n54666;
  assign n54890 = n54620 & n54889;
  assign n54891 = n54626 & n54890;
  assign n54892 = n54626 & n54699;
  assign n54893 = ~n54874 & ~n54892;
  assign n54894 = n54620 & ~n54893;
  assign n54895 = ~n54891 & ~n54894;
  assign n54896 = ~n54620 & n54658;
  assign n54897 = n54895 & ~n54896;
  assign n54898 = ~n54888 & n54897;
  assign n54899 = ~n54882 & n54898;
  assign n54900 = ~n54877 & n54899;
  assign n54901 = ~n54620 & n54626;
  assign n54902 = n54701 & n54901;
  assign n54903 = n54900 & ~n54902;
  assign n54904 = ~pi1518 & ~n54903;
  assign n54905 = ~n54877 & ~n54902;
  assign n54906 = n54899 & n54905;
  assign n54907 = pi1518 & n54906;
  assign po1600 = n54904 | n54907;
  assign n54909 = ~n54421 & n54450;
  assign n54910 = ~n54427 & n54909;
  assign n54911 = n54433 & n54461;
  assign n54912 = n54421 & n54911;
  assign n54913 = n54470 & n54473;
  assign n54914 = ~n54912 & ~n54913;
  assign n54915 = ~n54433 & n54461;
  assign n54916 = ~n54421 & n54915;
  assign n54917 = ~n54453 & ~n54916;
  assign n54918 = ~n54450 & ~n54917;
  assign n54919 = n54914 & ~n54918;
  assign n54920 = ~n54910 & n54919;
  assign n54921 = n54415 & ~n54920;
  assign n54922 = n54421 & n54491;
  assign n54923 = n54450 & n54922;
  assign n54924 = ~n54421 & ~n54450;
  assign n54925 = n54491 & n54924;
  assign n54926 = ~n54453 & ~n54483;
  assign n54927 = ~n54421 & n54470;
  assign n54928 = n54926 & ~n54927;
  assign n54929 = n54450 & ~n54928;
  assign n54930 = ~n54925 & ~n54929;
  assign n54931 = ~n54450 & n54457;
  assign n54932 = ~n54451 & n54476;
  assign n54933 = ~n54931 & n54932;
  assign n54934 = n54930 & n54933;
  assign n54935 = ~n54415 & ~n54934;
  assign n54936 = ~n54923 & ~n54935;
  assign n54937 = ~n54921 & n54936;
  assign n54938 = n54483 & n54924;
  assign n54939 = n54421 & n54485;
  assign n54940 = ~n54938 & ~n54939;
  assign n54941 = ~n54450 & n54913;
  assign n54942 = n54940 & ~n54941;
  assign n54943 = n54937 & n54942;
  assign n54944 = ~pi1513 & ~n54943;
  assign n54945 = pi1513 & n54942;
  assign n54946 = n54936 & n54945;
  assign n54947 = ~n54921 & n54946;
  assign po1601 = n54944 | n54947;
  assign n54949 = ~n54259 & n54280;
  assign n54950 = ~n54259 & n54322;
  assign n54951 = ~n54949 & ~n54950;
  assign n54952 = n54265 & n54951;
  assign n54953 = ~n54253 & ~n54274;
  assign n54954 = ~n54273 & ~n54953;
  assign n54955 = n54246 & n54299;
  assign n54956 = n54259 & n54274;
  assign n54957 = ~n54955 & ~n54956;
  assign n54958 = n54259 & n54317;
  assign n54959 = n54957 & ~n54958;
  assign n54960 = ~n54954 & n54959;
  assign n54961 = ~n54265 & n54960;
  assign n54962 = ~n54952 & ~n54961;
  assign n54963 = n54273 & n54280;
  assign n54964 = n54259 & n54963;
  assign n54965 = n54259 & n54954;
  assign n54966 = ~n54964 & ~n54965;
  assign n54967 = ~n54962 & n54966;
  assign n54968 = n54240 & ~n54967;
  assign n54969 = n54265 & ~n54953;
  assign n54970 = ~n54259 & n54969;
  assign n54971 = ~n54294 & ~n54321;
  assign n54972 = n54259 & ~n54971;
  assign n54973 = n54265 & n54972;
  assign n54974 = n54273 & n54969;
  assign n54975 = ~n54973 & ~n54974;
  assign n54976 = ~n54970 & n54975;
  assign n54977 = ~n54240 & ~n54976;
  assign n54978 = ~n54968 & ~n54977;
  assign n54979 = ~n54265 & ~n54951;
  assign n54980 = ~n54278 & ~n54979;
  assign n54981 = ~n54240 & ~n54980;
  assign n54982 = n54265 & n54278;
  assign n54983 = ~n54265 & ~n54966;
  assign n54984 = ~n54982 & ~n54983;
  assign n54985 = ~n54981 & n54984;
  assign n54986 = n54978 & n54985;
  assign n54987 = pi1522 & ~n54986;
  assign n54988 = ~n54968 & n54985;
  assign n54989 = ~n54977 & n54988;
  assign n54990 = ~pi1522 & n54989;
  assign po1602 = n54987 | n54990;
  assign n54992 = n54519 & ~n54525;
  assign n54993 = ~n54563 & ~n54992;
  assign n54994 = ~n54594 & n54993;
  assign n54995 = n54544 & ~n54994;
  assign n54996 = n54538 & ~n54544;
  assign n54997 = n54525 & n54996;
  assign n54998 = n54519 & n54538;
  assign n54999 = ~n54531 & n54998;
  assign n55000 = ~n54538 & n54552;
  assign n55001 = ~n54999 & ~n55000;
  assign n55002 = ~n54519 & ~n54525;
  assign n55003 = ~n54538 & ~n54544;
  assign n55004 = n55002 & n55003;
  assign n55005 = n55001 & ~n55004;
  assign n55006 = ~n54997 & n55005;
  assign n55007 = ~n54995 & n55006;
  assign n55008 = n54513 & ~n55007;
  assign n55009 = n54519 & n54579;
  assign n55010 = n54538 & n55009;
  assign n55011 = n54519 & n54532;
  assign n55012 = ~n54538 & n55011;
  assign n55013 = ~n55010 & ~n55012;
  assign n55014 = n54544 & ~n55013;
  assign n55015 = ~n55008 & ~n55014;
  assign n55016 = n54538 & n54552;
  assign n55017 = ~n54567 & ~n54575;
  assign n55018 = n54544 & ~n55017;
  assign n55019 = ~n55016 & ~n55018;
  assign n55020 = ~n54571 & n55019;
  assign n55021 = ~n54513 & ~n55020;
  assign n55022 = ~n54549 & ~n54579;
  assign n55023 = ~n54519 & ~n55022;
  assign n55024 = ~n54580 & ~n55023;
  assign n55025 = ~n54544 & ~n55024;
  assign n55026 = ~n54513 & n55025;
  assign n55027 = ~n55021 & ~n55026;
  assign n55028 = n55015 & n55027;
  assign n55029 = ~pi1510 & n55028;
  assign n55030 = pi1510 & ~n55028;
  assign po1604 = n55029 | n55030;
  assign n55032 = pi5116 & pi9040;
  assign n55033 = pi4882 & ~pi9040;
  assign n55034 = ~n55032 & ~n55033;
  assign n55035 = ~pi1482 & ~n55034;
  assign n55036 = pi1482 & n55034;
  assign n55037 = ~n55035 & ~n55036;
  assign n55038 = pi4840 & pi9040;
  assign n55039 = pi4923 & ~pi9040;
  assign n55040 = ~n55038 & ~n55039;
  assign n55041 = ~pi1490 & ~n55040;
  assign n55042 = pi1490 & n55040;
  assign n55043 = ~n55041 & ~n55042;
  assign n55044 = pi4943 & ~pi9040;
  assign n55045 = pi4923 & pi9040;
  assign n55046 = ~n55044 & ~n55045;
  assign n55047 = ~pi1491 & ~n55046;
  assign n55048 = pi1491 & n55046;
  assign n55049 = ~n55047 & ~n55048;
  assign n55050 = n55043 & ~n55049;
  assign n55051 = pi5059 & pi9040;
  assign n55052 = pi4963 & ~pi9040;
  assign n55053 = ~n55051 & ~n55052;
  assign n55054 = ~pi1494 & ~n55053;
  assign n55055 = pi1494 & n55053;
  assign n55056 = ~n55054 & ~n55055;
  assign n55057 = pi4846 & pi9040;
  assign n55058 = pi4962 & ~pi9040;
  assign n55059 = ~n55057 & ~n55058;
  assign n55060 = ~pi1499 & n55059;
  assign n55061 = pi1499 & ~n55059;
  assign n55062 = ~n55060 & ~n55061;
  assign n55063 = ~n55056 & n55062;
  assign n55064 = pi4838 & pi9040;
  assign n55065 = pi4984 & ~pi9040;
  assign n55066 = ~n55064 & ~n55065;
  assign n55067 = ~pi1467 & n55066;
  assign n55068 = pi1467 & ~n55066;
  assign n55069 = ~n55067 & ~n55068;
  assign n55070 = n55056 & ~n55062;
  assign n55071 = n55069 & n55070;
  assign n55072 = ~n55063 & ~n55071;
  assign n55073 = n55050 & ~n55072;
  assign n55074 = ~n55049 & n55069;
  assign n55075 = n55063 & n55074;
  assign n55076 = ~n55073 & ~n55075;
  assign n55077 = n55037 & ~n55076;
  assign n55078 = ~n55043 & ~n55069;
  assign n55079 = ~n55062 & n55078;
  assign n55080 = n55056 & n55079;
  assign n55081 = n55056 & ~n55069;
  assign n55082 = ~n55078 & ~n55081;
  assign n55083 = n55049 & ~n55082;
  assign n55084 = ~n55043 & n55069;
  assign n55085 = n55062 & n55084;
  assign n55086 = n55056 & n55085;
  assign n55087 = ~n55083 & ~n55086;
  assign n55088 = ~n55080 & n55087;
  assign n55089 = n55037 & ~n55088;
  assign n55090 = ~n55077 & ~n55089;
  assign n55091 = n55043 & ~n55069;
  assign n55092 = ~n55062 & n55091;
  assign n55093 = ~n55056 & n55092;
  assign n55094 = ~n55056 & ~n55062;
  assign n55095 = n55069 & n55094;
  assign n55096 = ~n55043 & n55095;
  assign n55097 = ~n55093 & ~n55096;
  assign n55098 = ~n55049 & ~n55097;
  assign n55099 = n55062 & ~n55069;
  assign n55100 = ~n55095 & ~n55099;
  assign n55101 = ~n55043 & ~n55100;
  assign n55102 = ~n55043 & ~n55062;
  assign n55103 = n55074 & n55102;
  assign n55104 = n55056 & n55062;
  assign n55105 = ~n55081 & ~n55104;
  assign n55106 = n55043 & ~n55105;
  assign n55107 = ~n55095 & ~n55106;
  assign n55108 = ~n55049 & ~n55107;
  assign n55109 = n55043 & n55049;
  assign n55110 = n55070 & n55109;
  assign n55111 = n55069 & n55110;
  assign n55112 = ~n55108 & ~n55111;
  assign n55113 = ~n55103 & n55112;
  assign n55114 = ~n55101 & n55113;
  assign n55115 = ~n55093 & n55114;
  assign n55116 = ~n55037 & ~n55115;
  assign n55117 = n55063 & n55069;
  assign n55118 = n55043 & n55117;
  assign n55119 = ~n55043 & n55081;
  assign n55120 = ~n55118 & ~n55119;
  assign n55121 = n55049 & ~n55120;
  assign n55122 = ~n55116 & ~n55121;
  assign n55123 = ~n55098 & n55122;
  assign n55124 = n55090 & n55123;
  assign n55125 = pi1519 & n55124;
  assign n55126 = ~pi1519 & ~n55124;
  assign po1605 = n55125 | n55126;
  assign n55128 = n54259 & n54287;
  assign n55129 = ~n54306 & ~n54315;
  assign n55130 = n54265 & ~n55129;
  assign n55131 = ~n55128 & ~n55130;
  assign n55132 = ~n54301 & n55131;
  assign n55133 = ~n54265 & n54304;
  assign n55134 = ~n54293 & ~n55133;
  assign n55135 = ~n54323 & n55134;
  assign n55136 = n55132 & n55135;
  assign n55137 = n54240 & ~n55136;
  assign n55138 = ~n54278 & ~n54964;
  assign n55139 = ~n54288 & ~n54950;
  assign n55140 = n54253 & n54273;
  assign n55141 = n54265 & n55140;
  assign n55142 = n54259 & n54292;
  assign n55143 = ~n55141 & ~n55142;
  assign n55144 = n54252 & ~n54273;
  assign n55145 = ~n54246 & n54259;
  assign n55146 = ~n55144 & ~n55145;
  assign n55147 = ~n54328 & n55146;
  assign n55148 = ~n54265 & ~n55147;
  assign n55149 = n55143 & ~n55148;
  assign n55150 = n55139 & n55149;
  assign n55151 = n55138 & n55150;
  assign n55152 = ~n54240 & ~n55151;
  assign n55153 = ~n55137 & ~n55152;
  assign n55154 = pi1521 & ~n55153;
  assign n55155 = ~pi1521 & ~n55137;
  assign n55156 = ~n55152 & n55155;
  assign po1606 = n55154 | n55156;
  assign n55158 = ~n54421 & n54911;
  assign n55159 = ~n54471 & ~n54480;
  assign n55160 = n54421 & n54440;
  assign n55161 = ~n54421 & n54491;
  assign n55162 = ~n55160 & ~n55161;
  assign n55163 = n55159 & n55162;
  assign n55164 = n54450 & ~n55163;
  assign n55165 = n54421 & n54452;
  assign n55166 = ~n54451 & ~n55165;
  assign n55167 = ~n54915 & n55166;
  assign n55168 = ~n54450 & ~n55167;
  assign n55169 = n54439 & n54473;
  assign n55170 = ~n54427 & n55169;
  assign n55171 = ~n55168 & ~n55170;
  assign n55172 = ~n55164 & n55171;
  assign n55173 = ~n55158 & n55172;
  assign n55174 = ~n54415 & ~n55173;
  assign n55175 = n54421 & n54450;
  assign n55176 = n54457 & n55175;
  assign n55177 = n54450 & n54915;
  assign n55178 = n54450 & n54483;
  assign n55179 = ~n55177 & ~n55178;
  assign n55180 = ~n54421 & ~n55179;
  assign n55181 = ~n55176 & ~n55180;
  assign n55182 = n54421 & n54470;
  assign n55183 = ~n54421 & n54452;
  assign n55184 = ~n55182 & ~n55183;
  assign n55185 = ~n54441 & n55184;
  assign n55186 = ~n54471 & n55185;
  assign n55187 = ~n54450 & ~n55186;
  assign n55188 = ~n54421 & n54453;
  assign n55189 = ~n55187 & ~n55188;
  assign n55190 = ~n54421 & n54441;
  assign n55191 = ~n54922 & ~n55190;
  assign n55192 = n55189 & n55191;
  assign n55193 = n55181 & n55192;
  assign n55194 = n54415 & ~n55193;
  assign n55195 = n54450 & ~n54914;
  assign n55196 = ~n55194 & ~n55195;
  assign n55197 = ~n54475 & ~n55190;
  assign n55198 = ~n54450 & ~n55197;
  assign n55199 = n55196 & ~n55198;
  assign n55200 = ~n55174 & n55199;
  assign n55201 = pi1520 & ~n55200;
  assign n55202 = ~pi1520 & n55200;
  assign po1607 = n55201 | n55202;
  assign n55204 = n54626 & n54869;
  assign n55205 = n54644 & n54651;
  assign n55206 = ~n54889 & ~n55205;
  assign n55207 = ~n54620 & ~n55206;
  assign n55208 = ~n55204 & ~n55207;
  assign n55209 = n54620 & n54626;
  assign n55210 = n54698 & n55209;
  assign n55211 = n54620 & n54646;
  assign n55212 = ~n55210 & ~n55211;
  assign n55213 = n55208 & n55212;
  assign n55214 = n54644 & n54656;
  assign n55215 = ~n54647 & ~n55214;
  assign n55216 = ~n54705 & n55215;
  assign n55217 = n55213 & n55216;
  assign n55218 = ~n54665 & ~n55217;
  assign n55219 = ~n54689 & ~n54695;
  assign n55220 = ~n54658 & ~n54889;
  assign n55221 = ~n54707 & n55220;
  assign n55222 = n54620 & ~n55221;
  assign n55223 = ~n54626 & n54864;
  assign n55224 = ~n54680 & ~n55223;
  assign n55225 = ~n54902 & n55224;
  assign n55226 = ~n54620 & n54704;
  assign n55227 = n55225 & ~n55226;
  assign n55228 = ~n55222 & n55227;
  assign n55229 = n54665 & ~n55228;
  assign n55230 = ~n54647 & n55224;
  assign n55231 = n54620 & ~n55230;
  assign n55232 = ~n55229 & ~n55231;
  assign n55233 = n55219 & n55232;
  assign n55234 = ~n55218 & n55233;
  assign n55235 = pi1526 & ~n55234;
  assign n55236 = ~pi1526 & n55234;
  assign po1608 = n55235 | n55236;
  assign n55238 = n55091 & n55104;
  assign n55239 = n55043 & n55069;
  assign n55240 = ~n55056 & n55239;
  assign n55241 = ~n55238 & ~n55240;
  assign n55242 = ~n55049 & ~n55241;
  assign n55243 = ~n55043 & n55049;
  assign n55244 = n55056 & n55243;
  assign n55245 = n55069 & n55104;
  assign n55246 = ~n55069 & n55070;
  assign n55247 = ~n55245 & ~n55246;
  assign n55248 = n55063 & ~n55069;
  assign n55249 = n55043 & n55248;
  assign n55250 = n55247 & ~n55249;
  assign n55251 = n55049 & ~n55250;
  assign n55252 = ~n55244 & ~n55251;
  assign n55253 = n55043 & n55095;
  assign n55254 = n55252 & ~n55253;
  assign n55255 = ~n55043 & n55063;
  assign n55256 = ~n55069 & n55094;
  assign n55257 = ~n55255 & ~n55256;
  assign n55258 = ~n55049 & ~n55257;
  assign n55259 = ~n55043 & n55071;
  assign n55260 = ~n55258 & ~n55259;
  assign n55261 = n55254 & n55260;
  assign n55262 = n55037 & ~n55261;
  assign n55263 = ~n55242 & ~n55262;
  assign n55264 = ~n55037 & n55049;
  assign n55265 = ~n55257 & n55264;
  assign n55266 = ~n55071 & ~n55117;
  assign n55267 = n55043 & ~n55266;
  assign n55268 = ~n55238 & ~n55267;
  assign n55269 = ~n55037 & ~n55268;
  assign n55270 = ~n55265 & ~n55269;
  assign n55271 = ~n55037 & ~n55049;
  assign n55272 = ~n55043 & n55104;
  assign n55273 = ~n55095 & ~n55272;
  assign n55274 = ~n55081 & n55273;
  assign n55275 = n55271 & ~n55274;
  assign n55276 = n55270 & ~n55275;
  assign n55277 = n55263 & n55276;
  assign n55278 = ~pi1517 & ~n55277;
  assign n55279 = pi1517 & n55270;
  assign n55280 = n55263 & n55279;
  assign n55281 = ~n55275 & n55280;
  assign po1609 = n55278 | n55281;
  assign n55283 = ~n54538 & n54570;
  assign n55284 = ~n55000 & ~n55283;
  assign n55285 = ~n54544 & ~n55284;
  assign n55286 = n54567 & n54996;
  assign n55287 = ~n55285 & ~n55286;
  assign n55288 = ~n54591 & n55287;
  assign n55289 = n54519 & n54544;
  assign n55290 = n54531 & n55289;
  assign n55291 = ~n54525 & n55290;
  assign n55292 = ~n54538 & n55291;
  assign n55293 = n54538 & n54575;
  assign n55294 = ~n54570 & ~n55293;
  assign n55295 = ~n55009 & n55294;
  assign n55296 = ~n54544 & ~n55295;
  assign n55297 = n54513 & n55296;
  assign n55298 = n54544 & n55011;
  assign n55299 = ~n54563 & ~n54589;
  assign n55300 = ~n54554 & n55299;
  assign n55301 = ~n55298 & n55300;
  assign n55302 = n54513 & ~n55301;
  assign n55303 = n54538 & n54600;
  assign n55304 = ~n55291 & ~n55303;
  assign n55305 = ~n54999 & n55304;
  assign n55306 = n54531 & n54561;
  assign n55307 = n54538 & n54549;
  assign n55308 = ~n54566 & ~n55307;
  assign n55309 = ~n54544 & ~n55308;
  assign n55310 = ~n55306 & ~n55309;
  assign n55311 = n55305 & n55310;
  assign n55312 = ~n54513 & ~n55311;
  assign n55313 = ~n55302 & ~n55312;
  assign n55314 = ~n55297 & n55313;
  assign n55315 = ~n55292 & n55314;
  assign n55316 = n55288 & n55315;
  assign n55317 = pi1516 & ~n55316;
  assign n55318 = ~pi1516 & n55288;
  assign n55319 = n55315 & n55318;
  assign po1610 = n55317 | n55319;
  assign n55321 = ~n54574 & ~n55011;
  assign n55322 = n54548 & ~n55321;
  assign n55323 = ~n54570 & ~n54575;
  assign n55324 = ~n54567 & ~n55009;
  assign n55325 = n55323 & n55324;
  assign n55326 = n54538 & ~n55325;
  assign n55327 = ~n55322 & ~n55326;
  assign n55328 = ~n55000 & n55327;
  assign n55329 = n54513 & ~n55328;
  assign n55330 = ~n54538 & n54567;
  assign n55331 = n54538 & n55011;
  assign n55332 = ~n55330 & ~n55331;
  assign n55333 = ~n54544 & ~n55332;
  assign n55334 = n54538 & ~n55022;
  assign n55335 = ~n54519 & n55334;
  assign n55336 = ~n54544 & ~n55321;
  assign n55337 = n54531 & n54998;
  assign n55338 = ~n54603 & ~n55337;
  assign n55339 = ~n55009 & n55338;
  assign n55340 = n54544 & ~n55339;
  assign n55341 = ~n55336 & ~n55340;
  assign n55342 = ~n55335 & n55341;
  assign n55343 = ~n55330 & n55342;
  assign n55344 = ~n54513 & ~n55343;
  assign n55345 = ~n55333 & ~n55344;
  assign n55346 = ~n55329 & n55345;
  assign n55347 = ~pi1507 & ~n55346;
  assign n55348 = pi1507 & ~n55333;
  assign n55349 = ~n55329 & n55348;
  assign n55350 = ~n55344 & n55349;
  assign po1612 = n55347 | n55350;
  assign n55352 = pi5059 & ~pi9040;
  assign n55353 = pi4882 & pi9040;
  assign n55354 = ~n55352 & ~n55353;
  assign n55355 = pi1477 & n55354;
  assign n55356 = ~pi1477 & ~n55354;
  assign n55357 = ~n55355 & ~n55356;
  assign n55358 = pi4837 & pi9040;
  assign n55359 = pi4834 & ~pi9040;
  assign n55360 = ~n55358 & ~n55359;
  assign n55361 = ~pi1475 & n55360;
  assign n55362 = pi1475 & ~n55360;
  assign n55363 = ~n55361 & ~n55362;
  assign n55364 = pi4846 & ~pi9040;
  assign n55365 = pi4984 & pi9040;
  assign n55366 = ~n55364 & ~n55365;
  assign n55367 = ~pi1499 & ~n55366;
  assign n55368 = pi1499 & n55366;
  assign n55369 = ~n55367 & ~n55368;
  assign n55370 = pi4834 & pi9040;
  assign n55371 = pi4833 & ~pi9040;
  assign n55372 = ~n55370 & ~n55371;
  assign n55373 = ~pi1482 & n55372;
  assign n55374 = pi1482 & ~n55372;
  assign n55375 = ~n55373 & ~n55374;
  assign n55376 = pi4961 & pi9040;
  assign n55377 = pi4835 & ~pi9040;
  assign n55378 = ~n55376 & ~n55377;
  assign n55379 = ~pi1500 & ~n55378;
  assign n55380 = pi1500 & n55378;
  assign n55381 = ~n55379 & ~n55380;
  assign n55382 = n55375 & n55381;
  assign n55383 = n55369 & n55382;
  assign n55384 = ~n55363 & n55383;
  assign n55385 = ~n55357 & n55384;
  assign n55386 = ~n55375 & ~n55381;
  assign n55387 = ~n55357 & ~n55363;
  assign n55388 = n55386 & n55387;
  assign n55389 = ~n55369 & n55388;
  assign n55390 = ~n55385 & ~n55389;
  assign n55391 = ~n55369 & n55382;
  assign n55392 = ~n55357 & n55363;
  assign n55393 = n55391 & n55392;
  assign n55394 = ~n55369 & n55386;
  assign n55395 = ~n55357 & n55394;
  assign n55396 = ~n55393 & ~n55395;
  assign n55397 = ~n55375 & n55381;
  assign n55398 = n55375 & ~n55381;
  assign n55399 = ~n55397 & ~n55398;
  assign n55400 = ~n55357 & ~n55369;
  assign n55401 = n55363 & ~n55400;
  assign n55402 = ~n55399 & n55401;
  assign n55403 = n55369 & ~n55375;
  assign n55404 = n55357 & n55403;
  assign n55405 = n55357 & n55382;
  assign n55406 = ~n55404 & ~n55405;
  assign n55407 = ~n55363 & ~n55406;
  assign n55408 = ~n55357 & ~n55382;
  assign n55409 = ~n55363 & n55408;
  assign n55410 = ~n55369 & n55409;
  assign n55411 = ~n55407 & ~n55410;
  assign n55412 = ~n55402 & n55411;
  assign n55413 = n55396 & n55412;
  assign n55414 = pi4909 & pi9040;
  assign n55415 = pi5039 & ~pi9040;
  assign n55416 = ~n55414 & ~n55415;
  assign n55417 = ~pi1473 & ~n55416;
  assign n55418 = pi1473 & n55416;
  assign n55419 = ~n55417 & ~n55418;
  assign n55420 = ~n55413 & n55419;
  assign n55421 = n55390 & ~n55420;
  assign n55422 = n55369 & n55397;
  assign n55423 = n55363 & n55422;
  assign n55424 = n55357 & n55423;
  assign n55425 = n55363 & ~n55419;
  assign n55426 = n55369 & n55386;
  assign n55427 = ~n55405 & ~n55426;
  assign n55428 = ~n55399 & n55400;
  assign n55429 = n55427 & ~n55428;
  assign n55430 = n55425 & ~n55429;
  assign n55431 = n55357 & n55394;
  assign n55432 = n55357 & ~n55375;
  assign n55433 = ~n55369 & n55432;
  assign n55434 = n55357 & n55398;
  assign n55435 = ~n55433 & ~n55434;
  assign n55436 = ~n55357 & n55382;
  assign n55437 = n55369 & n55398;
  assign n55438 = ~n55436 & ~n55437;
  assign n55439 = n55435 & n55438;
  assign n55440 = ~n55363 & ~n55439;
  assign n55441 = ~n55431 & ~n55440;
  assign n55442 = ~n55419 & ~n55441;
  assign n55443 = ~n55430 & ~n55442;
  assign n55444 = ~n55424 & n55443;
  assign n55445 = n55421 & n55444;
  assign n55446 = pi1533 & ~n55445;
  assign n55447 = ~pi1533 & n55421;
  assign n55448 = n55444 & n55447;
  assign po1613 = n55446 | n55448;
  assign n55450 = ~n55434 & ~n55436;
  assign n55451 = ~n55363 & ~n55450;
  assign n55452 = ~n55389 & ~n55451;
  assign n55453 = n55419 & ~n55452;
  assign n55454 = ~n55369 & ~n55375;
  assign n55455 = ~n55397 & ~n55454;
  assign n55456 = ~n55357 & ~n55455;
  assign n55457 = ~n55383 & ~n55456;
  assign n55458 = n55363 & ~n55457;
  assign n55459 = ~n55428 & ~n55458;
  assign n55460 = n55357 & n55391;
  assign n55461 = ~n55357 & n55369;
  assign n55462 = ~n55381 & n55461;
  assign n55463 = n55357 & ~n55455;
  assign n55464 = ~n55462 & ~n55463;
  assign n55465 = ~n55363 & ~n55464;
  assign n55466 = ~n55460 & ~n55465;
  assign n55467 = n55459 & n55466;
  assign n55468 = ~n55419 & ~n55467;
  assign n55469 = n55357 & n55369;
  assign n55470 = ~n55397 & n55469;
  assign n55471 = n55419 & n55470;
  assign n55472 = n55357 & ~n55369;
  assign n55473 = n55397 & n55472;
  assign n55474 = ~n55363 & n55473;
  assign n55475 = n55357 & n55363;
  assign n55476 = n55369 & n55475;
  assign n55477 = ~n55381 & n55476;
  assign n55478 = ~n55474 & ~n55477;
  assign n55479 = ~n55471 & n55478;
  assign n55480 = ~n55432 & ~n55437;
  assign n55481 = n55363 & n55419;
  assign n55482 = ~n55480 & n55481;
  assign n55483 = n55479 & ~n55482;
  assign n55484 = ~n55468 & n55483;
  assign n55485 = ~n55453 & n55484;
  assign n55486 = pi1532 & ~n55485;
  assign n55487 = ~pi1532 & n55485;
  assign po1614 = n55486 | n55487;
  assign n55489 = n55062 & n55239;
  assign n55490 = ~n55071 & ~n55489;
  assign n55491 = ~n55049 & ~n55490;
  assign n55492 = n55043 & n55094;
  assign n55493 = ~n55085 & ~n55492;
  assign n55494 = n55049 & ~n55493;
  assign n55495 = ~n55043 & n55248;
  assign n55496 = ~n55103 & ~n55495;
  assign n55497 = ~n55238 & n55496;
  assign n55498 = ~n55494 & n55497;
  assign n55499 = ~n55491 & n55498;
  assign n55500 = ~n55080 & ~n55093;
  assign n55501 = n55499 & n55500;
  assign n55502 = n55037 & ~n55501;
  assign n55503 = n55078 & n55104;
  assign n55504 = n55266 & ~n55503;
  assign n55505 = n55049 & ~n55504;
  assign n55506 = ~n55043 & n55256;
  assign n55507 = ~n55505 & ~n55506;
  assign n55508 = n55056 & n55239;
  assign n55509 = n55043 & n55070;
  assign n55510 = ~n55508 & ~n55509;
  assign n55511 = n55049 & ~n55510;
  assign n55512 = n55049 & n55094;
  assign n55513 = ~n55043 & n55512;
  assign n55514 = ~n55511 & ~n55513;
  assign n55515 = n55507 & n55514;
  assign n55516 = ~n55037 & ~n55515;
  assign n55517 = ~n55248 & ~n55253;
  assign n55518 = ~n55086 & n55517;
  assign n55519 = n55271 & ~n55518;
  assign n55520 = ~n55516 & ~n55519;
  assign n55521 = ~n55080 & ~n55238;
  assign n55522 = ~n55049 & ~n55521;
  assign n55523 = n55520 & ~n55522;
  assign n55524 = ~n55502 & n55523;
  assign n55525 = ~pi1525 & n55524;
  assign n55526 = pi1525 & ~n55524;
  assign po1615 = n55525 | n55526;
  assign n55528 = n54767 & ~n54773;
  assign n55529 = ~n54761 & n55528;
  assign n55530 = n54787 & n55529;
  assign n55531 = ~n54773 & n54805;
  assign n55532 = ~n54767 & ~n54779;
  assign n55533 = ~n54787 & n55532;
  assign n55534 = ~n54797 & ~n55533;
  assign n55535 = ~n55531 & n55534;
  assign n55536 = ~n55530 & n55535;
  assign n55537 = n54761 & n54793;
  assign n55538 = n55536 & ~n55537;
  assign n55539 = n54829 & ~n55538;
  assign n55540 = ~n54787 & n54799;
  assign n55541 = ~n54847 & ~n55540;
  assign n55542 = n54761 & ~n55541;
  assign n55543 = ~n54761 & ~n54829;
  assign n55544 = n54831 & n55543;
  assign n55545 = ~n54767 & ~n54787;
  assign n55546 = n54773 & n55545;
  assign n55547 = ~n55532 & ~n55546;
  assign n55548 = ~n54799 & n55547;
  assign n55549 = n54761 & ~n55548;
  assign n55550 = n54767 & n54816;
  assign n55551 = ~n54787 & n55550;
  assign n55552 = ~n55549 & ~n55551;
  assign n55553 = ~n54829 & ~n55552;
  assign n55554 = ~n55544 & ~n55553;
  assign n55555 = ~n55542 & n55554;
  assign n55556 = n54787 & n54831;
  assign n55557 = ~n54787 & n54846;
  assign n55558 = ~n55556 & ~n55557;
  assign n55559 = ~n54794 & n55558;
  assign n55560 = ~n54797 & n55559;
  assign n55561 = ~n54761 & ~n55560;
  assign n55562 = n55555 & ~n55561;
  assign n55563 = ~n55539 & n55562;
  assign n55564 = ~pi1553 & ~n55563;
  assign n55565 = pi1553 & n55555;
  assign n55566 = ~n55539 & n55565;
  assign n55567 = ~n55561 & n55566;
  assign po1616 = n55564 | n55567;
  assign n55569 = ~n54873 & ~n54879;
  assign n55570 = n54665 & ~n55569;
  assign n55571 = ~n54657 & ~n54672;
  assign n55572 = ~n54861 & n55571;
  assign n55573 = n54620 & ~n55572;
  assign n55574 = n54665 & n55573;
  assign n55575 = ~n55570 & ~n55574;
  assign n55576 = n54667 & n54675;
  assign n55577 = ~n54677 & ~n55576;
  assign n55578 = ~n54671 & ~n54708;
  assign n55579 = ~n54620 & ~n55578;
  assign n55580 = n54665 & n55579;
  assign n55581 = n55577 & ~n55580;
  assign n55582 = n54626 & n54667;
  assign n55583 = n54626 & n54645;
  assign n55584 = ~n54653 & ~n55583;
  assign n55585 = ~n54620 & ~n55584;
  assign n55586 = ~n54658 & ~n54680;
  assign n55587 = n54626 & n54666;
  assign n55588 = ~n54701 & ~n55587;
  assign n55589 = n54620 & ~n55588;
  assign n55590 = n55586 & ~n55589;
  assign n55591 = ~n55585 & n55590;
  assign n55592 = ~n55582 & n55591;
  assign n55593 = ~n54665 & ~n55592;
  assign n55594 = ~n54705 & n55224;
  assign n55595 = ~n54620 & ~n55594;
  assign n55596 = ~n55593 & ~n55595;
  assign n55597 = n55581 & n55596;
  assign n55598 = n55575 & n55597;
  assign n55599 = ~pi1537 & ~n55598;
  assign n55600 = pi1537 & n55581;
  assign n55601 = n55575 & n55600;
  assign n55602 = n55596 & n55601;
  assign po1617 = n55599 | n55602;
  assign n55604 = ~n54794 & ~n54806;
  assign n55605 = ~n54761 & ~n54787;
  assign n55606 = ~n54779 & n55605;
  assign n55607 = ~n54773 & n55606;
  assign n55608 = n54798 & n54832;
  assign n55609 = ~n55607 & ~n55608;
  assign n55610 = ~n54761 & n54841;
  assign n55611 = n55609 & ~n55610;
  assign n55612 = ~n54787 & n54820;
  assign n55613 = ~n54817 & ~n55556;
  assign n55614 = n54761 & ~n55613;
  assign n55615 = ~n55612 & ~n55614;
  assign n55616 = n54779 & n54796;
  assign n55617 = n55615 & ~n55616;
  assign n55618 = n55611 & n55617;
  assign n55619 = n55604 & n55618;
  assign n55620 = ~n54829 & ~n55619;
  assign n55621 = ~n54793 & ~n54817;
  assign n55622 = n54787 & ~n55621;
  assign n55623 = ~n54787 & n54816;
  assign n55624 = ~n55531 & ~n55623;
  assign n55625 = ~n54761 & ~n55624;
  assign n55626 = ~n54773 & n54835;
  assign n55627 = ~n54846 & ~n55626;
  assign n55628 = n54787 & n55532;
  assign n55629 = n55627 & ~n55628;
  assign n55630 = n54761 & ~n55629;
  assign n55631 = ~n55540 & ~n55630;
  assign n55632 = ~n55625 & n55631;
  assign n55633 = ~n55622 & n55632;
  assign n55634 = n54829 & ~n55633;
  assign n55635 = n54761 & n54836;
  assign n55636 = ~n55634 & ~n55635;
  assign n55637 = n54811 & n55605;
  assign n55638 = ~n54779 & n55637;
  assign n55639 = n55636 & ~n55638;
  assign n55640 = ~n55620 & n55639;
  assign n55641 = ~pi1527 & ~n55640;
  assign n55642 = pi1527 & n55636;
  assign n55643 = ~n55620 & n55642;
  assign n55644 = ~n55638 & n55643;
  assign po1618 = n55641 | n55644;
  assign n55646 = n54259 & n55140;
  assign n55647 = n54265 & n55646;
  assign n55648 = n54299 & ~n54953;
  assign n55649 = ~n54322 & ~n55648;
  assign n55650 = ~n54964 & n55649;
  assign n55651 = ~n54265 & ~n55650;
  assign n55652 = n54259 & n54275;
  assign n55653 = ~n55651 & ~n55652;
  assign n55654 = n54273 & n54321;
  assign n55655 = ~n54259 & n55144;
  assign n55656 = ~n55654 & ~n55655;
  assign n55657 = ~n54956 & n55656;
  assign n55658 = n54265 & ~n55657;
  assign n55659 = n55653 & ~n55658;
  assign n55660 = n54240 & ~n55659;
  assign n55661 = ~n55647 & ~n55660;
  assign n55662 = ~n54259 & n54274;
  assign n55663 = ~n54963 & ~n55662;
  assign n55664 = n54265 & ~n55663;
  assign n55665 = ~n54323 & ~n55664;
  assign n55666 = ~n54295 & ~n55646;
  assign n55667 = n54259 & n54328;
  assign n55668 = ~n55144 & ~n55667;
  assign n55669 = ~n55654 & n55668;
  assign n55670 = ~n54265 & ~n55669;
  assign n55671 = ~n54259 & n54275;
  assign n55672 = ~n55670 & ~n55671;
  assign n55673 = n55666 & n55672;
  assign n55674 = n55665 & n55673;
  assign n55675 = ~n54240 & ~n55674;
  assign n55676 = ~n54309 & ~n54958;
  assign n55677 = ~n54265 & ~n55676;
  assign n55678 = ~n55675 & ~n55677;
  assign n55679 = n55661 & n55678;
  assign n55680 = pi1530 & n55679;
  assign n55681 = ~pi1530 & ~n55679;
  assign po1619 = n55680 | n55681;
  assign n55683 = ~n54916 & ~n55190;
  assign n55684 = ~n55170 & n55683;
  assign n55685 = n54450 & ~n55684;
  assign n55686 = ~n54925 & ~n54941;
  assign n55687 = ~n54922 & ~n55178;
  assign n55688 = ~n54911 & ~n55183;
  assign n55689 = ~n54450 & ~n55688;
  assign n55690 = ~n54480 & ~n55689;
  assign n55691 = n55687 & n55690;
  assign n55692 = n54415 & ~n55691;
  assign n55693 = ~n54433 & n54439;
  assign n55694 = ~n54458 & ~n55693;
  assign n55695 = n54421 & ~n55694;
  assign n55696 = ~n54441 & ~n54927;
  assign n55697 = ~n54450 & ~n55696;
  assign n55698 = n54421 & n54439;
  assign n55699 = ~n54453 & ~n55698;
  assign n55700 = ~n54461 & n55699;
  assign n55701 = n54450 & ~n55700;
  assign n55702 = ~n55697 & ~n55701;
  assign n55703 = ~n55695 & n55702;
  assign n55704 = ~n54415 & ~n55703;
  assign n55705 = ~n55692 & ~n55704;
  assign n55706 = n55686 & n55705;
  assign n55707 = ~n55685 & n55706;
  assign n55708 = ~pi1540 & ~n55707;
  assign n55709 = pi1540 & n55686;
  assign n55710 = ~n55685 & n55709;
  assign n55711 = n55705 & n55710;
  assign po1620 = n55708 | n55711;
  assign n55713 = n55381 & n55461;
  assign n55714 = ~n55394 & ~n55422;
  assign n55715 = ~n55713 & n55714;
  assign n55716 = n55481 & ~n55715;
  assign n55717 = n55357 & n55419;
  assign n55718 = n55437 & n55717;
  assign n55719 = ~n55363 & n55426;
  assign n55720 = ~n55369 & n55381;
  assign n55721 = ~n55405 & ~n55720;
  assign n55722 = ~n55363 & ~n55721;
  assign n55723 = ~n55719 & ~n55722;
  assign n55724 = n55419 & ~n55723;
  assign n55725 = ~n55718 & ~n55724;
  assign n55726 = n55381 & n55472;
  assign n55727 = ~n55357 & n55398;
  assign n55728 = ~n55369 & n55727;
  assign n55729 = ~n55726 & ~n55728;
  assign n55730 = ~n55363 & ~n55729;
  assign n55731 = n55725 & ~n55730;
  assign n55732 = n55382 & n55475;
  assign n55733 = n55369 & n55732;
  assign n55734 = ~n55399 & n55461;
  assign n55735 = ~n55395 & ~n55734;
  assign n55736 = ~n55399 & n55472;
  assign n55737 = n55357 & n55426;
  assign n55738 = ~n55736 & ~n55737;
  assign n55739 = ~n55393 & n55738;
  assign n55740 = n55735 & n55739;
  assign n55741 = ~n55733 & n55740;
  assign n55742 = n55369 & n55387;
  assign n55743 = n55375 & n55742;
  assign n55744 = n55741 & ~n55743;
  assign n55745 = ~n55419 & ~n55744;
  assign n55746 = n55731 & ~n55745;
  assign n55747 = ~n55716 & n55746;
  assign n55748 = ~pi1531 & ~n55747;
  assign n55749 = pi1531 & n55731;
  assign n55750 = ~n55716 & n55749;
  assign n55751 = ~n55745 & n55750;
  assign po1621 = n55748 | n55751;
  assign n55753 = ~n55369 & n55397;
  assign n55754 = ~n55383 & ~n55753;
  assign n55755 = ~n55363 & ~n55754;
  assign n55756 = ~n55422 & ~n55727;
  assign n55757 = ~n55391 & n55756;
  assign n55758 = n55363 & ~n55757;
  assign n55759 = ~n55755 & ~n55758;
  assign n55760 = ~n55719 & ~n55728;
  assign n55761 = n55759 & n55760;
  assign n55762 = ~n55419 & ~n55761;
  assign n55763 = ~n55357 & n55386;
  assign n55764 = ~n55434 & ~n55763;
  assign n55765 = n55363 & ~n55764;
  assign n55766 = n55357 & n55383;
  assign n55767 = ~n55765 & ~n55766;
  assign n55768 = ~n55363 & n55369;
  assign n55769 = ~n55381 & n55768;
  assign n55770 = n55375 & n55769;
  assign n55771 = n55714 & ~n55770;
  assign n55772 = ~n55391 & n55771;
  assign n55773 = ~n55357 & ~n55772;
  assign n55774 = n55767 & ~n55773;
  assign n55775 = n55419 & ~n55774;
  assign n55776 = ~n55762 & ~n55775;
  assign n55777 = ~n55369 & n55434;
  assign n55778 = ~n55737 & ~n55777;
  assign n55779 = ~n55363 & ~n55778;
  assign n55780 = n55363 & n55454;
  assign n55781 = n55357 & n55780;
  assign n55782 = ~n55779 & ~n55781;
  assign n55783 = n55776 & n55782;
  assign n55784 = ~pi1523 & ~n55783;
  assign n55785 = pi1523 & ~n55779;
  assign n55786 = n55776 & n55785;
  assign n55787 = ~n55781 & n55786;
  assign po1622 = n55784 | n55787;
  assign n55789 = ~n54788 & ~n54797;
  assign n55790 = ~n54761 & ~n55789;
  assign n55791 = ~n54853 & ~n55790;
  assign n55792 = n54767 & n54773;
  assign n55793 = n54761 & n55792;
  assign n55794 = n54787 & n55793;
  assign n55795 = n54787 & n54816;
  assign n55796 = ~n55792 & ~n55795;
  assign n55797 = ~n54773 & n55545;
  assign n55798 = n55796 & ~n55797;
  assign n55799 = n54761 & ~n55798;
  assign n55800 = ~n54800 & ~n55799;
  assign n55801 = ~n54829 & ~n55800;
  assign n55802 = ~n54761 & n54780;
  assign n55803 = n54787 & n55802;
  assign n55804 = ~n55610 & ~n55803;
  assign n55805 = ~n54829 & ~n55804;
  assign n55806 = ~n55801 & ~n55805;
  assign n55807 = ~n55794 & n55806;
  assign n55808 = ~n54817 & ~n54836;
  assign n55809 = ~n54846 & n55808;
  assign n55810 = ~n54761 & ~n55809;
  assign n55811 = ~n54787 & n54841;
  assign n55812 = ~n54820 & ~n55811;
  assign n55813 = n54761 & ~n55812;
  assign n55814 = ~n55810 & ~n55813;
  assign n55815 = ~n55626 & n55814;
  assign n55816 = ~n54806 & ~n54847;
  assign n55817 = n55815 & n55816;
  assign n55818 = n54829 & ~n55817;
  assign n55819 = n55807 & ~n55818;
  assign n55820 = n55791 & n55819;
  assign n55821 = ~pi1543 & ~n55820;
  assign n55822 = pi1543 & n55807;
  assign n55823 = n55791 & n55822;
  assign n55824 = ~n55818 & n55823;
  assign po1624 = n55821 | n55824;
  assign n55826 = ~n55043 & n55070;
  assign n55827 = ~n55245 & ~n55826;
  assign n55828 = ~n55049 & ~n55827;
  assign n55829 = n55049 & ~n55100;
  assign n55830 = ~n55828 & ~n55829;
  assign n55831 = ~n55118 & n55830;
  assign n55832 = n55037 & ~n55831;
  assign n55833 = ~n55049 & n55256;
  assign n55834 = ~n55832 & ~n55833;
  assign n55835 = ~n55495 & ~n55509;
  assign n55836 = n55049 & ~n55835;
  assign n55837 = n55050 & ~n55069;
  assign n55838 = ~n55084 & ~n55837;
  assign n55839 = ~n55056 & ~n55838;
  assign n55840 = n55049 & n55246;
  assign n55841 = n55043 & n55071;
  assign n55842 = ~n55840 & ~n55841;
  assign n55843 = ~n55238 & n55842;
  assign n55844 = ~n55085 & n55843;
  assign n55845 = ~n55839 & n55844;
  assign n55846 = ~n55037 & ~n55845;
  assign n55847 = ~n55836 & ~n55846;
  assign n55848 = n55834 & n55847;
  assign n55849 = pi1557 & n55848;
  assign n55850 = ~pi1557 & ~n55848;
  assign po1625 = n55849 | n55850;
  assign n55852 = pi5194 & pi9040;
  assign n55853 = pi5112 & ~pi9040;
  assign n55854 = ~n55852 & ~n55853;
  assign n55855 = ~pi1551 & ~n55854;
  assign n55856 = pi1551 & n55854;
  assign n55857 = ~n55855 & ~n55856;
  assign n55858 = pi5262 & ~pi9040;
  assign n55859 = pi5065 & pi9040;
  assign n55860 = ~n55858 & ~n55859;
  assign n55861 = ~pi1560 & n55860;
  assign n55862 = pi1560 & ~n55860;
  assign n55863 = ~n55861 & ~n55862;
  assign n55864 = pi5075 & pi9040;
  assign n55865 = pi5245 & ~pi9040;
  assign n55866 = ~n55864 & ~n55865;
  assign n55867 = ~pi1528 & n55866;
  assign n55868 = pi1528 & ~n55866;
  assign n55869 = ~n55867 & ~n55868;
  assign n55870 = pi5262 & pi9040;
  assign n55871 = pi5194 & ~pi9040;
  assign n55872 = ~n55870 & ~n55871;
  assign n55873 = ~pi1542 & n55872;
  assign n55874 = pi1542 & ~n55872;
  assign n55875 = ~n55873 & ~n55874;
  assign n55876 = pi5255 & pi9040;
  assign n55877 = pi5067 & ~pi9040;
  assign n55878 = ~n55876 & ~n55877;
  assign n55879 = pi1558 & n55878;
  assign n55880 = ~pi1558 & ~n55878;
  assign n55881 = ~n55879 & ~n55880;
  assign n55882 = n55875 & ~n55881;
  assign n55883 = ~n55869 & n55882;
  assign n55884 = n55863 & n55883;
  assign n55885 = pi5151 & pi9040;
  assign n55886 = pi5065 & ~pi9040;
  assign n55887 = ~n55885 & ~n55886;
  assign n55888 = ~pi1539 & n55887;
  assign n55889 = pi1539 & ~n55887;
  assign n55890 = ~n55888 & ~n55889;
  assign n55891 = ~n55863 & n55869;
  assign n55892 = ~n55890 & n55891;
  assign n55893 = ~n55875 & n55890;
  assign n55894 = n55869 & n55893;
  assign n55895 = n55863 & n55894;
  assign n55896 = ~n55892 & ~n55895;
  assign n55897 = ~n55863 & ~n55869;
  assign n55898 = ~n55875 & n55897;
  assign n55899 = n55896 & ~n55898;
  assign n55900 = ~n55881 & ~n55899;
  assign n55901 = ~n55863 & n55890;
  assign n55902 = n55875 & n55881;
  assign n55903 = n55901 & n55902;
  assign n55904 = n55875 & n55890;
  assign n55905 = n55891 & n55904;
  assign n55906 = ~n55903 & ~n55905;
  assign n55907 = ~n55900 & n55906;
  assign n55908 = ~n55884 & n55907;
  assign n55909 = n55863 & ~n55869;
  assign n55910 = ~n55890 & n55909;
  assign n55911 = n55875 & n55910;
  assign n55912 = ~n55890 & n55897;
  assign n55913 = ~n55875 & n55912;
  assign n55914 = ~n55911 & ~n55913;
  assign n55915 = n55908 & n55914;
  assign n55916 = ~n55857 & ~n55915;
  assign n55917 = n55890 & n55897;
  assign n55918 = n55875 & n55917;
  assign n55919 = ~n55910 & ~n55918;
  assign n55920 = ~n55881 & ~n55919;
  assign n55921 = n55893 & n55909;
  assign n55922 = n55869 & n55904;
  assign n55923 = n55863 & n55922;
  assign n55924 = ~n55921 & ~n55923;
  assign n55925 = ~n55863 & n55893;
  assign n55926 = n55875 & n55912;
  assign n55927 = ~n55925 & ~n55926;
  assign n55928 = n55881 & ~n55927;
  assign n55929 = n55924 & ~n55928;
  assign n55930 = ~n55920 & n55929;
  assign n55931 = n55857 & ~n55930;
  assign n55932 = ~n55863 & ~n55890;
  assign n55933 = ~n55875 & n55932;
  assign n55934 = n55863 & ~n55890;
  assign n55935 = n55875 & n55934;
  assign n55936 = ~n55933 & ~n55935;
  assign n55937 = ~n55881 & ~n55936;
  assign n55938 = n55863 & n55869;
  assign n55939 = ~n55890 & n55938;
  assign n55940 = ~n55875 & n55939;
  assign n55941 = ~n55921 & ~n55940;
  assign n55942 = n55890 & n55891;
  assign n55943 = n55941 & ~n55942;
  assign n55944 = n55881 & ~n55943;
  assign n55945 = ~n55937 & ~n55944;
  assign n55946 = n55869 & n55890;
  assign n55947 = n55881 & n55946;
  assign n55948 = n55875 & n55947;
  assign n55949 = n55945 & ~n55948;
  assign n55950 = ~n55931 & n55949;
  assign n55951 = ~n55916 & n55950;
  assign n55952 = ~pi1571 & ~n55951;
  assign n55953 = pi1571 & n55951;
  assign po1649 = n55952 | n55953;
  assign n55955 = pi5144 & pi9040;
  assign n55956 = pi5302 & ~pi9040;
  assign n55957 = ~n55955 & ~n55956;
  assign n55958 = ~pi1564 & ~n55957;
  assign n55959 = pi1564 & n55957;
  assign n55960 = ~n55958 & ~n55959;
  assign n55961 = pi5069 & ~pi9040;
  assign n55962 = pi5064 & pi9040;
  assign n55963 = ~n55961 & ~n55962;
  assign n55964 = ~pi1562 & ~n55963;
  assign n55965 = pi1562 & n55963;
  assign n55966 = ~n55964 & ~n55965;
  assign n55967 = pi5267 & ~pi9040;
  assign n55968 = pi5193 & pi9040;
  assign n55969 = ~n55967 & ~n55968;
  assign n55970 = ~pi1563 & n55969;
  assign n55971 = pi1563 & ~n55969;
  assign n55972 = ~n55970 & ~n55971;
  assign n55973 = n55966 & n55972;
  assign n55974 = n55960 & n55973;
  assign n55975 = pi5078 & ~pi9040;
  assign n55976 = pi5312 & pi9040;
  assign n55977 = ~n55975 & ~n55976;
  assign n55978 = pi1547 & n55977;
  assign n55979 = ~pi1547 & ~n55977;
  assign n55980 = ~n55978 & ~n55979;
  assign n55981 = ~n55960 & n55980;
  assign n55982 = ~n55966 & n55981;
  assign n55983 = ~n55974 & ~n55982;
  assign n55984 = pi5117 & ~pi9040;
  assign n55985 = pi5314 & pi9040;
  assign n55986 = ~n55984 & ~n55985;
  assign n55987 = ~pi1529 & n55986;
  assign n55988 = pi1529 & ~n55986;
  assign n55989 = ~n55987 & ~n55988;
  assign n55990 = ~n55960 & ~n55989;
  assign n55991 = ~n55966 & n55990;
  assign n55992 = n55983 & ~n55991;
  assign n55993 = ~n55966 & n55989;
  assign n55994 = n55960 & n55993;
  assign n55995 = ~n55980 & n55994;
  assign n55996 = n55992 & ~n55995;
  assign n55997 = ~n55960 & n55989;
  assign n55998 = n55980 & n55997;
  assign n55999 = ~n55966 & ~n55989;
  assign n56000 = ~n55998 & ~n55999;
  assign n56001 = ~n55972 & ~n56000;
  assign n56002 = ~n55972 & n55990;
  assign n56003 = ~n55980 & n56002;
  assign n56004 = ~n56001 & ~n56003;
  assign n56005 = n55996 & n56004;
  assign n56006 = pi5066 & pi9040;
  assign n56007 = pi5193 & ~pi9040;
  assign n56008 = ~n56006 & ~n56007;
  assign n56009 = ~pi1548 & ~n56008;
  assign n56010 = pi1548 & n56008;
  assign n56011 = ~n56009 & ~n56010;
  assign n56012 = ~n56005 & n56011;
  assign n56013 = n55972 & n55980;
  assign n56014 = n55994 & n56013;
  assign n56015 = n55966 & ~n55980;
  assign n56016 = ~n55960 & n56015;
  assign n56017 = ~n55980 & n55997;
  assign n56018 = ~n56016 & ~n56017;
  assign n56019 = n55972 & ~n56018;
  assign n56020 = ~n56014 & ~n56019;
  assign n56021 = ~n56011 & ~n56020;
  assign n56022 = n55960 & n55989;
  assign n56023 = n55966 & n56022;
  assign n56024 = ~n55972 & n56023;
  assign n56025 = n55980 & n56024;
  assign n56026 = n55980 & n55990;
  assign n56027 = ~n55972 & n56026;
  assign n56028 = n55966 & n56027;
  assign n56029 = ~n55980 & n55989;
  assign n56030 = n55966 & n56029;
  assign n56031 = ~n55960 & n56030;
  assign n56032 = n55960 & ~n55989;
  assign n56033 = ~n55972 & n56032;
  assign n56034 = ~n55980 & n56033;
  assign n56035 = ~n56031 & ~n56034;
  assign n56036 = ~n56028 & n56035;
  assign n56037 = ~n56025 & n56036;
  assign n56038 = ~n55966 & ~n55980;
  assign n56039 = ~n55989 & n56038;
  assign n56040 = n55960 & n56039;
  assign n56041 = n56037 & ~n56040;
  assign n56042 = ~n56011 & ~n56041;
  assign n56043 = n55989 & n56015;
  assign n56044 = n55960 & n55966;
  assign n56045 = ~n55989 & n56044;
  assign n56046 = n55980 & n56045;
  assign n56047 = ~n56043 & ~n56046;
  assign n56048 = n55980 & n55991;
  assign n56049 = n56047 & ~n56048;
  assign n56050 = n55972 & ~n56049;
  assign n56051 = ~n55966 & n55980;
  assign n56052 = ~n55972 & n56051;
  assign n56053 = n55997 & n56052;
  assign n56054 = ~n56050 & ~n56053;
  assign n56055 = ~n56042 & n56054;
  assign n56056 = ~n56021 & n56055;
  assign n56057 = ~n56012 & n56056;
  assign n56058 = ~n55972 & ~n55980;
  assign n56059 = n55960 & ~n55966;
  assign n56060 = n56058 & n56059;
  assign n56061 = n56057 & ~n56060;
  assign n56062 = ~pi1575 & ~n56061;
  assign n56063 = pi1575 & ~n56060;
  assign n56064 = n56057 & n56063;
  assign po1650 = n56062 | n56064;
  assign n56066 = pi5182 & pi9040;
  assign n56067 = pi5439 & ~pi9040;
  assign n56068 = ~n56066 & ~n56067;
  assign n56069 = ~pi1534 & ~n56068;
  assign n56070 = pi1534 & n56068;
  assign n56071 = ~n56069 & ~n56070;
  assign n56072 = pi5076 & ~pi9040;
  assign n56073 = pi5156 & pi9040;
  assign n56074 = ~n56072 & ~n56073;
  assign n56075 = ~pi1528 & n56074;
  assign n56076 = pi1528 & ~n56074;
  assign n56077 = ~n56075 & ~n56076;
  assign n56078 = pi5164 & ~pi9040;
  assign n56079 = pi5440 & pi9040;
  assign n56080 = ~n56078 & ~n56079;
  assign n56081 = ~pi1562 & n56080;
  assign n56082 = pi1562 & ~n56080;
  assign n56083 = ~n56081 & ~n56082;
  assign n56084 = pi5192 & ~pi9040;
  assign n56085 = pi5253 & pi9040;
  assign n56086 = ~n56084 & ~n56085;
  assign n56087 = ~pi1551 & n56086;
  assign n56088 = pi1551 & ~n56086;
  assign n56089 = ~n56087 & ~n56088;
  assign n56090 = ~n56083 & ~n56089;
  assign n56091 = n56077 & n56090;
  assign n56092 = pi5250 & ~pi9040;
  assign n56093 = pi5155 & pi9040;
  assign n56094 = ~n56092 & ~n56093;
  assign n56095 = pi1561 & n56094;
  assign n56096 = ~pi1561 & ~n56094;
  assign n56097 = ~n56095 & ~n56096;
  assign n56098 = n56091 & ~n56097;
  assign n56099 = n56083 & n56089;
  assign n56100 = n56077 & n56099;
  assign n56101 = ~n56097 & n56100;
  assign n56102 = ~n56098 & ~n56101;
  assign n56103 = ~n56077 & n56099;
  assign n56104 = n56097 & n56103;
  assign n56105 = ~n56083 & n56089;
  assign n56106 = n56077 & n56105;
  assign n56107 = n56097 & n56106;
  assign n56108 = ~n56104 & ~n56107;
  assign n56109 = n56102 & n56108;
  assign n56110 = n56071 & ~n56109;
  assign n56111 = n56083 & ~n56089;
  assign n56112 = n56077 & n56111;
  assign n56113 = n56097 & n56112;
  assign n56114 = ~n56106 & ~n56113;
  assign n56115 = n56071 & ~n56114;
  assign n56116 = ~n56071 & ~n56089;
  assign n56117 = ~n56097 & n56116;
  assign n56118 = ~n56077 & ~n56083;
  assign n56119 = n56097 & n56099;
  assign n56120 = ~n56118 & ~n56119;
  assign n56121 = ~n56071 & ~n56120;
  assign n56122 = ~n56117 & ~n56121;
  assign n56123 = ~n56077 & n56111;
  assign n56124 = ~n56097 & n56123;
  assign n56125 = n56122 & ~n56124;
  assign n56126 = ~n56089 & n56118;
  assign n56127 = n56097 & n56126;
  assign n56128 = n56125 & ~n56127;
  assign n56129 = ~n56115 & n56128;
  assign n56130 = pi5112 & pi9040;
  assign n56131 = pi5058 & ~pi9040;
  assign n56132 = ~n56130 & ~n56131;
  assign n56133 = ~pi1564 & ~n56132;
  assign n56134 = pi1564 & n56132;
  assign n56135 = ~n56133 & ~n56134;
  assign n56136 = ~n56129 & ~n56135;
  assign n56137 = n56077 & ~n56089;
  assign n56138 = ~n56071 & n56097;
  assign n56139 = n56135 & n56138;
  assign n56140 = n56137 & n56139;
  assign n56141 = n56077 & ~n56097;
  assign n56142 = n56089 & n56141;
  assign n56143 = ~n56071 & ~n56142;
  assign n56144 = ~n56077 & n56097;
  assign n56145 = n56083 & n56144;
  assign n56146 = ~n56090 & ~n56137;
  assign n56147 = ~n56097 & ~n56146;
  assign n56148 = ~n56103 & ~n56147;
  assign n56149 = n56071 & n56148;
  assign n56150 = ~n56145 & n56149;
  assign n56151 = ~n56143 & ~n56150;
  assign n56152 = ~n56077 & n56105;
  assign n56153 = n56097 & n56152;
  assign n56154 = ~n56151 & ~n56153;
  assign n56155 = n56135 & ~n56154;
  assign n56156 = ~n56140 & ~n56155;
  assign n56157 = ~n56136 & n56156;
  assign n56158 = ~n56110 & n56157;
  assign n56159 = ~n56071 & n56124;
  assign n56160 = n56158 & ~n56159;
  assign n56161 = pi1568 & ~n56160;
  assign n56162 = ~pi1568 & ~n56159;
  assign n56163 = n56157 & n56162;
  assign n56164 = ~n56110 & n56163;
  assign po1653 = n56161 | n56164;
  assign n56166 = pi5083 & pi9040;
  assign n56167 = pi5156 & ~pi9040;
  assign n56168 = ~n56166 & ~n56167;
  assign n56169 = ~pi1546 & ~n56168;
  assign n56170 = pi1546 & n56168;
  assign n56171 = ~n56169 & ~n56170;
  assign n56172 = pi5072 & ~pi9040;
  assign n56173 = pi5439 & pi9040;
  assign n56174 = ~n56172 & ~n56173;
  assign n56175 = pi1567 & n56174;
  assign n56176 = ~pi1567 & ~n56174;
  assign n56177 = ~n56175 & ~n56176;
  assign n56178 = pi5192 & pi9040;
  assign n56179 = pi5182 & ~pi9040;
  assign n56180 = ~n56178 & ~n56179;
  assign n56181 = pi1565 & n56180;
  assign n56182 = ~pi1565 & ~n56180;
  assign n56183 = ~n56181 & ~n56182;
  assign n56184 = pi5083 & ~pi9040;
  assign n56185 = pi5058 & pi9040;
  assign n56186 = ~n56184 & ~n56185;
  assign n56187 = ~pi1536 & n56186;
  assign n56188 = pi1536 & ~n56186;
  assign n56189 = ~n56187 & ~n56188;
  assign n56190 = pi5164 & pi9040;
  assign n56191 = pi5155 & ~pi9040;
  assign n56192 = ~n56190 & ~n56191;
  assign n56193 = pi1556 & n56192;
  assign n56194 = ~pi1556 & ~n56192;
  assign n56195 = ~n56193 & ~n56194;
  assign n56196 = ~n56189 & ~n56195;
  assign n56197 = n56183 & n56196;
  assign n56198 = n56177 & n56197;
  assign n56199 = ~n56177 & ~n56189;
  assign n56200 = n56195 & n56199;
  assign n56201 = pi5076 & pi9040;
  assign n56202 = pi5440 & ~pi9040;
  assign n56203 = ~n56201 & ~n56202;
  assign n56204 = pi1538 & n56203;
  assign n56205 = ~pi1538 & ~n56203;
  assign n56206 = ~n56204 & ~n56205;
  assign n56207 = ~n56183 & n56199;
  assign n56208 = n56183 & n56195;
  assign n56209 = n56189 & n56208;
  assign n56210 = ~n56207 & ~n56209;
  assign n56211 = ~n56206 & ~n56210;
  assign n56212 = ~n56200 & ~n56211;
  assign n56213 = ~n56189 & n56208;
  assign n56214 = ~n56183 & n56189;
  assign n56215 = ~n56213 & ~n56214;
  assign n56216 = n56189 & ~n56195;
  assign n56217 = ~n56177 & n56216;
  assign n56218 = ~n56183 & ~n56195;
  assign n56219 = n56177 & n56218;
  assign n56220 = ~n56217 & ~n56219;
  assign n56221 = n56215 & n56220;
  assign n56222 = n56206 & ~n56221;
  assign n56223 = n56212 & ~n56222;
  assign n56224 = ~n56198 & n56223;
  assign n56225 = n56171 & ~n56224;
  assign n56226 = ~n56183 & n56195;
  assign n56227 = n56189 & n56226;
  assign n56228 = ~n56177 & n56227;
  assign n56229 = n56189 & n56218;
  assign n56230 = n56177 & n56229;
  assign n56231 = ~n56198 & ~n56230;
  assign n56232 = ~n56228 & n56231;
  assign n56233 = n56206 & ~n56232;
  assign n56234 = ~n56225 & ~n56233;
  assign n56235 = n56183 & n56200;
  assign n56236 = n56183 & n56189;
  assign n56237 = ~n56206 & n56236;
  assign n56238 = n56177 & n56237;
  assign n56239 = ~n56177 & n56206;
  assign n56240 = ~n56189 & n56239;
  assign n56241 = ~n56195 & n56240;
  assign n56242 = ~n56189 & n56226;
  assign n56243 = n56177 & n56242;
  assign n56244 = ~n56241 & ~n56243;
  assign n56245 = ~n56183 & ~n56189;
  assign n56246 = n56177 & n56245;
  assign n56247 = n56183 & ~n56195;
  assign n56248 = n56189 & n56247;
  assign n56249 = ~n56246 & ~n56248;
  assign n56250 = ~n56206 & ~n56249;
  assign n56251 = ~n56183 & ~n56206;
  assign n56252 = n56189 & n56251;
  assign n56253 = ~n56177 & n56252;
  assign n56254 = ~n56250 & ~n56253;
  assign n56255 = n56244 & n56254;
  assign n56256 = ~n56171 & ~n56255;
  assign n56257 = ~n56238 & ~n56256;
  assign n56258 = ~n56235 & n56257;
  assign n56259 = n56234 & n56258;
  assign n56260 = ~pi1570 & ~n56259;
  assign n56261 = ~n56225 & ~n56235;
  assign n56262 = ~n56233 & n56261;
  assign n56263 = n56257 & n56262;
  assign n56264 = pi1570 & n56263;
  assign po1655 = n56260 | n56264;
  assign n56266 = pi5355 & pi9040;
  assign n56267 = pi5073 & ~pi9040;
  assign n56268 = ~n56266 & ~n56267;
  assign n56269 = ~pi1565 & ~n56268;
  assign n56270 = pi1565 & n56268;
  assign n56271 = ~n56269 & ~n56270;
  assign n56272 = pi5089 & pi9040;
  assign n56273 = pi5074 & ~pi9040;
  assign n56274 = ~n56272 & ~n56273;
  assign n56275 = ~pi1550 & n56274;
  assign n56276 = pi1550 & ~n56274;
  assign n56277 = ~n56275 & ~n56276;
  assign n56278 = pi5315 & pi9040;
  assign n56279 = pi5061 & ~pi9040;
  assign n56280 = ~n56278 & ~n56279;
  assign n56281 = pi1554 & n56280;
  assign n56282 = ~pi1554 & ~n56280;
  assign n56283 = ~n56281 & ~n56282;
  assign n56284 = pi5068 & pi9040;
  assign n56285 = pi5312 & ~pi9040;
  assign n56286 = ~n56284 & ~n56285;
  assign n56287 = ~pi1549 & n56286;
  assign n56288 = pi1549 & ~n56286;
  assign n56289 = ~n56287 & ~n56288;
  assign n56290 = pi5062 & ~pi9040;
  assign n56291 = pi5061 & pi9040;
  assign n56292 = ~n56290 & ~n56291;
  assign n56293 = ~pi1536 & ~n56292;
  assign n56294 = pi1536 & n56292;
  assign n56295 = ~n56293 & ~n56294;
  assign n56296 = n56289 & n56295;
  assign n56297 = n56283 & n56296;
  assign n56298 = ~n56277 & n56297;
  assign n56299 = pi5070 & pi9040;
  assign n56300 = pi5195 & ~pi9040;
  assign n56301 = ~n56299 & ~n56300;
  assign n56302 = ~pi1566 & n56301;
  assign n56303 = pi1566 & ~n56301;
  assign n56304 = ~n56302 & ~n56303;
  assign n56305 = ~n56289 & n56295;
  assign n56306 = ~n56277 & n56305;
  assign n56307 = ~n56283 & n56296;
  assign n56308 = n56277 & n56307;
  assign n56309 = ~n56306 & ~n56308;
  assign n56310 = n56304 & ~n56309;
  assign n56311 = ~n56298 & ~n56310;
  assign n56312 = n56289 & ~n56295;
  assign n56313 = ~n56283 & n56312;
  assign n56314 = ~n56304 & n56313;
  assign n56315 = n56296 & ~n56304;
  assign n56316 = ~n56277 & n56315;
  assign n56317 = ~n56314 & ~n56316;
  assign n56318 = n56311 & n56317;
  assign n56319 = ~n56289 & ~n56295;
  assign n56320 = n56283 & n56319;
  assign n56321 = ~n56277 & n56320;
  assign n56322 = n56283 & n56312;
  assign n56323 = n56277 & n56322;
  assign n56324 = ~n56321 & ~n56323;
  assign n56325 = n56318 & n56324;
  assign n56326 = n56271 & ~n56325;
  assign n56327 = ~n56271 & n56304;
  assign n56328 = ~n56277 & ~n56283;
  assign n56329 = n56289 & n56328;
  assign n56330 = ~n56283 & ~n56295;
  assign n56331 = ~n56329 & ~n56330;
  assign n56332 = n56327 & ~n56331;
  assign n56333 = n56277 & n56283;
  assign n56334 = n56295 & n56333;
  assign n56335 = n56289 & n56334;
  assign n56336 = n56277 & ~n56289;
  assign n56337 = ~n56283 & n56336;
  assign n56338 = ~n56335 & ~n56337;
  assign n56339 = ~n56277 & ~n56304;
  assign n56340 = n56283 & n56339;
  assign n56341 = ~n56296 & n56340;
  assign n56342 = ~n56304 & n56320;
  assign n56343 = ~n56341 & ~n56342;
  assign n56344 = n56338 & n56343;
  assign n56345 = ~n56271 & ~n56344;
  assign n56346 = ~n56283 & n56319;
  assign n56347 = n56304 & n56346;
  assign n56348 = n56277 & n56347;
  assign n56349 = n56283 & n56305;
  assign n56350 = n56277 & n56349;
  assign n56351 = ~n56323 & ~n56350;
  assign n56352 = n56304 & ~n56351;
  assign n56353 = ~n56348 & ~n56352;
  assign n56354 = ~n56304 & n56335;
  assign n56355 = n56353 & ~n56354;
  assign n56356 = ~n56345 & n56355;
  assign n56357 = ~n56332 & n56356;
  assign n56358 = ~n56326 & n56357;
  assign n56359 = ~n56283 & n56305;
  assign n56360 = n56277 & ~n56304;
  assign n56361 = n56359 & n56360;
  assign n56362 = n56358 & ~n56361;
  assign n56363 = ~pi1573 & ~n56362;
  assign n56364 = pi1573 & ~n56361;
  assign n56365 = n56357 & n56364;
  assign n56366 = ~n56326 & n56365;
  assign po1656 = n56363 | n56366;
  assign n56368 = ~n55875 & n55942;
  assign n56369 = ~n55923 & ~n55932;
  assign n56370 = n55881 & ~n56369;
  assign n56371 = ~n56368 & ~n56370;
  assign n56372 = ~n55918 & n56371;
  assign n56373 = ~n55881 & n55921;
  assign n56374 = ~n55911 & ~n56373;
  assign n56375 = ~n55940 & n56374;
  assign n56376 = n56372 & n56375;
  assign n56377 = n55857 & ~n56376;
  assign n56378 = ~n55875 & n55917;
  assign n56379 = ~n55895 & ~n56378;
  assign n56380 = n55890 & n55909;
  assign n56381 = n55881 & n56380;
  assign n56382 = ~n55875 & n55910;
  assign n56383 = ~n56381 & ~n56382;
  assign n56384 = ~n55869 & ~n55890;
  assign n56385 = ~n55863 & ~n55875;
  assign n56386 = ~n56384 & ~n56385;
  assign n56387 = ~n55946 & n56386;
  assign n56388 = ~n55881 & ~n56387;
  assign n56389 = n55875 & n55939;
  assign n56390 = ~n55905 & ~n56389;
  assign n56391 = ~n56388 & n56390;
  assign n56392 = n56383 & n56391;
  assign n56393 = n56379 & n56392;
  assign n56394 = ~n55857 & ~n56393;
  assign n56395 = ~n56377 & ~n56394;
  assign n56396 = pi1572 & ~n56395;
  assign n56397 = ~pi1572 & ~n56377;
  assign n56398 = ~n56394 & n56397;
  assign po1659 = n56396 | n56398;
  assign n56400 = pi5255 & ~pi9040;
  assign n56401 = pi5326 & pi9040;
  assign n56402 = ~n56400 & ~n56401;
  assign n56403 = ~pi1560 & ~n56402;
  assign n56404 = pi1560 & n56402;
  assign n56405 = ~n56403 & ~n56404;
  assign n56406 = pi5250 & pi9040;
  assign n56407 = pi5189 & ~pi9040;
  assign n56408 = ~n56406 & ~n56407;
  assign n56409 = ~pi1541 & ~n56408;
  assign n56410 = pi1541 & n56408;
  assign n56411 = ~n56409 & ~n56410;
  assign n56412 = pi5253 & ~pi9040;
  assign n56413 = pi5067 & pi9040;
  assign n56414 = ~n56412 & ~n56413;
  assign n56415 = pi1535 & n56414;
  assign n56416 = ~pi1535 & ~n56414;
  assign n56417 = ~n56415 & ~n56416;
  assign n56418 = pi5075 & ~pi9040;
  assign n56419 = pi5188 & pi9040;
  assign n56420 = ~n56418 & ~n56419;
  assign n56421 = ~pi1546 & n56420;
  assign n56422 = pi1546 & ~n56420;
  assign n56423 = ~n56421 & ~n56422;
  assign n56424 = pi5079 & ~pi9040;
  assign n56425 = pi5189 & pi9040;
  assign n56426 = ~n56424 & ~n56425;
  assign n56427 = ~pi1556 & n56426;
  assign n56428 = pi1556 & ~n56426;
  assign n56429 = ~n56427 & ~n56428;
  assign n56430 = n56423 & ~n56429;
  assign n56431 = n56417 & n56430;
  assign n56432 = pi5143 & ~pi9040;
  assign n56433 = pi5245 & pi9040;
  assign n56434 = ~n56432 & ~n56433;
  assign n56435 = ~pi1539 & n56434;
  assign n56436 = pi1539 & ~n56434;
  assign n56437 = ~n56435 & ~n56436;
  assign n56438 = ~n56423 & ~n56437;
  assign n56439 = ~n56429 & n56438;
  assign n56440 = ~n56431 & ~n56439;
  assign n56441 = ~n56417 & n56429;
  assign n56442 = n56437 & n56441;
  assign n56443 = ~n56423 & n56442;
  assign n56444 = n56440 & ~n56443;
  assign n56445 = n56411 & ~n56444;
  assign n56446 = ~n56423 & n56429;
  assign n56447 = ~n56437 & n56446;
  assign n56448 = ~n56417 & n56447;
  assign n56449 = n56423 & ~n56437;
  assign n56450 = ~n56429 & n56449;
  assign n56451 = ~n56417 & n56450;
  assign n56452 = ~n56423 & n56437;
  assign n56453 = n56423 & n56429;
  assign n56454 = ~n56452 & ~n56453;
  assign n56455 = n56417 & ~n56454;
  assign n56456 = ~n56451 & ~n56455;
  assign n56457 = ~n56448 & n56456;
  assign n56458 = ~n56411 & ~n56457;
  assign n56459 = ~n56445 & ~n56458;
  assign n56460 = n56405 & ~n56459;
  assign n56461 = n56423 & n56437;
  assign n56462 = n56429 & n56461;
  assign n56463 = ~n56411 & n56462;
  assign n56464 = ~n56417 & n56463;
  assign n56465 = ~n56429 & n56452;
  assign n56466 = ~n56417 & n56465;
  assign n56467 = ~n56411 & n56466;
  assign n56468 = ~n56464 & ~n56467;
  assign n56469 = n56429 & n56449;
  assign n56470 = ~n56417 & n56469;
  assign n56471 = n56411 & n56470;
  assign n56472 = n56468 & ~n56471;
  assign n56473 = n56411 & ~n56417;
  assign n56474 = n56423 & n56473;
  assign n56475 = n56417 & n56447;
  assign n56476 = ~n56466 & ~n56475;
  assign n56477 = ~n56411 & ~n56417;
  assign n56478 = n56452 & n56477;
  assign n56479 = ~n56417 & ~n56423;
  assign n56480 = ~n56429 & n56479;
  assign n56481 = ~n56431 & ~n56480;
  assign n56482 = ~n56411 & ~n56481;
  assign n56483 = ~n56478 & ~n56482;
  assign n56484 = n56411 & n56417;
  assign n56485 = n56446 & n56484;
  assign n56486 = n56411 & n56429;
  assign n56487 = n56449 & n56486;
  assign n56488 = ~n56485 & ~n56487;
  assign n56489 = n56483 & n56488;
  assign n56490 = n56476 & n56489;
  assign n56491 = ~n56474 & n56490;
  assign n56492 = ~n56405 & ~n56491;
  assign n56493 = ~n56417 & ~n56429;
  assign n56494 = n56437 & n56493;
  assign n56495 = n56423 & n56494;
  assign n56496 = n56417 & n56438;
  assign n56497 = ~n56495 & ~n56496;
  assign n56498 = n56411 & ~n56497;
  assign n56499 = ~n56492 & ~n56498;
  assign n56500 = n56472 & n56499;
  assign n56501 = ~n56460 & n56500;
  assign n56502 = ~pi1588 & ~n56501;
  assign n56503 = pi1588 & n56501;
  assign po1661 = n56502 | n56503;
  assign n56505 = n56277 & n56313;
  assign n56506 = ~n56295 & n56328;
  assign n56507 = ~n56289 & n56506;
  assign n56508 = ~n56505 & ~n56507;
  assign n56509 = ~n56304 & ~n56508;
  assign n56510 = ~n56335 & ~n56342;
  assign n56511 = n56289 & n56333;
  assign n56512 = ~n56337 & ~n56511;
  assign n56513 = n56304 & ~n56512;
  assign n56514 = ~n56277 & n56304;
  assign n56515 = n56312 & n56514;
  assign n56516 = ~n56283 & n56515;
  assign n56517 = ~n56277 & n56283;
  assign n56518 = n56295 & n56517;
  assign n56519 = ~n56289 & n56518;
  assign n56520 = ~n56283 & ~n56304;
  assign n56521 = n56295 & n56520;
  assign n56522 = n56289 & n56521;
  assign n56523 = ~n56519 & ~n56522;
  assign n56524 = ~n56516 & n56523;
  assign n56525 = ~n56513 & n56524;
  assign n56526 = n56510 & n56525;
  assign n56527 = n56271 & ~n56526;
  assign n56528 = n56304 & n56335;
  assign n56529 = n56277 & n56342;
  assign n56530 = ~n56528 & ~n56529;
  assign n56531 = ~n56527 & n56530;
  assign n56532 = ~n56509 & n56531;
  assign n56533 = n56283 & n56289;
  assign n56534 = n56339 & n56533;
  assign n56535 = ~n56314 & ~n56534;
  assign n56536 = ~n56304 & n56349;
  assign n56537 = n56277 & n56359;
  assign n56538 = ~n56536 & ~n56537;
  assign n56539 = ~n56277 & n56322;
  assign n56540 = ~n56505 & ~n56539;
  assign n56541 = ~n56277 & n56319;
  assign n56542 = ~n56283 & n56295;
  assign n56543 = ~n56541 & ~n56542;
  assign n56544 = n56304 & ~n56543;
  assign n56545 = n56540 & ~n56544;
  assign n56546 = n56538 & n56545;
  assign n56547 = n56535 & n56546;
  assign n56548 = ~n56271 & ~n56547;
  assign n56549 = n56532 & ~n56548;
  assign n56550 = ~pi1582 & ~n56549;
  assign n56551 = pi1582 & n56532;
  assign n56552 = ~n56548 & n56551;
  assign po1662 = n56550 | n56552;
  assign n56554 = ~n56529 & ~n56534;
  assign n56555 = ~n56335 & ~n56346;
  assign n56556 = ~n56541 & n56555;
  assign n56557 = n56304 & ~n56556;
  assign n56558 = ~n56277 & n56307;
  assign n56559 = ~n56519 & ~n56558;
  assign n56560 = ~n56361 & n56559;
  assign n56561 = ~n56304 & n56322;
  assign n56562 = n56560 & ~n56561;
  assign n56563 = ~n56557 & n56562;
  assign n56564 = n56271 & ~n56563;
  assign n56565 = n56277 & n56315;
  assign n56566 = ~n56289 & n56328;
  assign n56567 = ~n56346 & ~n56566;
  assign n56568 = ~n56304 & ~n56567;
  assign n56569 = ~n56565 & ~n56568;
  assign n56570 = n56304 & n56305;
  assign n56571 = n56277 & n56570;
  assign n56572 = n56304 & n56313;
  assign n56573 = ~n56571 & ~n56572;
  assign n56574 = n56569 & n56573;
  assign n56575 = ~n56289 & n56333;
  assign n56576 = ~n56505 & ~n56575;
  assign n56577 = ~n56539 & n56576;
  assign n56578 = n56574 & n56577;
  assign n56579 = ~n56271 & ~n56578;
  assign n56580 = ~n56505 & n56559;
  assign n56581 = n56304 & ~n56580;
  assign n56582 = ~n56579 & ~n56581;
  assign n56583 = ~n56564 & n56582;
  assign n56584 = n56554 & n56583;
  assign n56585 = pi1584 & ~n56584;
  assign n56586 = ~pi1584 & n56584;
  assign po1663 = n56585 | n56586;
  assign n56588 = ~n55960 & n55966;
  assign n56589 = ~n56040 & ~n56588;
  assign n56590 = ~n55981 & n56589;
  assign n56591 = ~n55972 & ~n56590;
  assign n56592 = n55960 & n56013;
  assign n56593 = n55966 & n55980;
  assign n56594 = ~n55989 & n56593;
  assign n56595 = ~n55980 & n56023;
  assign n56596 = ~n56594 & ~n56595;
  assign n56597 = ~n55960 & ~n55966;
  assign n56598 = n55972 & ~n55980;
  assign n56599 = n56597 & n56598;
  assign n56600 = n56596 & ~n56599;
  assign n56601 = ~n56592 & n56600;
  assign n56602 = ~n56591 & n56601;
  assign n56603 = n56011 & ~n56602;
  assign n56604 = n55966 & n55997;
  assign n56605 = n55980 & n56604;
  assign n56606 = n55966 & n55990;
  assign n56607 = ~n55980 & n56606;
  assign n56608 = ~n56605 & ~n56607;
  assign n56609 = ~n55972 & ~n56608;
  assign n56610 = ~n56603 & ~n56609;
  assign n56611 = n55980 & n56023;
  assign n56612 = ~n55994 & ~n56045;
  assign n56613 = ~n55972 & ~n56612;
  assign n56614 = ~n56611 & ~n56613;
  assign n56615 = ~n56048 & n56614;
  assign n56616 = ~n56011 & ~n56615;
  assign n56617 = ~n55997 & ~n56032;
  assign n56618 = ~n55966 & ~n56617;
  assign n56619 = ~n56017 & ~n56618;
  assign n56620 = n55972 & ~n56619;
  assign n56621 = ~n56011 & n56620;
  assign n56622 = ~n56616 & ~n56621;
  assign n56623 = n56610 & n56622;
  assign n56624 = pi1576 & ~n56623;
  assign n56625 = ~pi1576 & n56610;
  assign n56626 = n56622 & n56625;
  assign po1664 = n56624 | n56626;
  assign n56628 = pi5078 & pi9040;
  assign n56629 = pi5066 & ~pi9040;
  assign n56630 = ~n56628 & ~n56629;
  assign n56631 = pi1552 & n56630;
  assign n56632 = ~pi1552 & ~n56630;
  assign n56633 = ~n56631 & ~n56632;
  assign n56634 = pi5154 & ~pi9040;
  assign n56635 = pi5196 & pi9040;
  assign n56636 = ~n56634 & ~n56635;
  assign n56637 = ~pi1548 & ~n56636;
  assign n56638 = pi1548 & n56636;
  assign n56639 = ~n56637 & ~n56638;
  assign n56640 = pi5314 & ~pi9040;
  assign n56641 = pi5190 & pi9040;
  assign n56642 = ~n56640 & ~n56641;
  assign n56643 = pi1545 & n56642;
  assign n56644 = ~pi1545 & ~n56642;
  assign n56645 = ~n56643 & ~n56644;
  assign n56646 = n56639 & ~n56645;
  assign n56647 = pi5195 & pi9040;
  assign n56648 = pi5190 & ~pi9040;
  assign n56649 = ~n56647 & ~n56648;
  assign n56650 = pi1559 & n56649;
  assign n56651 = ~pi1559 & ~n56649;
  assign n56652 = ~n56650 & ~n56651;
  assign n56653 = pi5117 & pi9040;
  assign n56654 = pi5416 & ~pi9040;
  assign n56655 = ~n56653 & ~n56654;
  assign n56656 = ~pi1529 & n56655;
  assign n56657 = pi1529 & ~n56655;
  assign n56658 = ~n56656 & ~n56657;
  assign n56659 = n56652 & ~n56658;
  assign n56660 = n56646 & n56659;
  assign n56661 = n56652 & n56658;
  assign n56662 = ~n56639 & n56661;
  assign n56663 = ~n56660 & ~n56662;
  assign n56664 = ~n56633 & ~n56663;
  assign n56665 = pi5252 & pi9040;
  assign n56666 = pi5068 & ~pi9040;
  assign n56667 = ~n56665 & ~n56666;
  assign n56668 = ~pi1544 & ~n56667;
  assign n56669 = pi1544 & n56667;
  assign n56670 = ~n56668 & ~n56669;
  assign n56671 = n56633 & ~n56652;
  assign n56672 = n56639 & n56671;
  assign n56673 = n56646 & n56658;
  assign n56674 = n56639 & n56645;
  assign n56675 = ~n56658 & n56674;
  assign n56676 = ~n56673 & ~n56675;
  assign n56677 = ~n56639 & ~n56645;
  assign n56678 = ~n56658 & n56677;
  assign n56679 = n56652 & n56678;
  assign n56680 = n56676 & ~n56679;
  assign n56681 = n56633 & ~n56680;
  assign n56682 = ~n56672 & ~n56681;
  assign n56683 = ~n56639 & n56645;
  assign n56684 = n56658 & n56683;
  assign n56685 = n56652 & n56684;
  assign n56686 = n56682 & ~n56685;
  assign n56687 = ~n56652 & n56677;
  assign n56688 = ~n56658 & n56683;
  assign n56689 = ~n56687 & ~n56688;
  assign n56690 = ~n56633 & ~n56689;
  assign n56691 = n56658 & n56674;
  assign n56692 = ~n56652 & n56691;
  assign n56693 = ~n56690 & ~n56692;
  assign n56694 = n56686 & n56693;
  assign n56695 = n56670 & ~n56694;
  assign n56696 = ~n56664 & ~n56695;
  assign n56697 = n56633 & ~n56670;
  assign n56698 = ~n56689 & n56697;
  assign n56699 = n56658 & n56677;
  assign n56700 = ~n56691 & ~n56699;
  assign n56701 = n56652 & ~n56700;
  assign n56702 = ~n56660 & ~n56701;
  assign n56703 = ~n56670 & ~n56702;
  assign n56704 = ~n56698 & ~n56703;
  assign n56705 = ~n56633 & ~n56670;
  assign n56706 = n56646 & ~n56652;
  assign n56707 = ~n56684 & ~n56706;
  assign n56708 = n56639 & ~n56658;
  assign n56709 = n56707 & ~n56708;
  assign n56710 = n56705 & ~n56709;
  assign n56711 = n56704 & ~n56710;
  assign n56712 = n56696 & n56711;
  assign n56713 = ~pi1569 & ~n56712;
  assign n56714 = pi1569 & n56704;
  assign n56715 = n56696 & n56714;
  assign n56716 = ~n56710 & n56715;
  assign po1666 = n56713 | n56716;
  assign n56718 = ~n56405 & ~n56411;
  assign n56719 = ~n56417 & n56430;
  assign n56720 = n56417 & n56465;
  assign n56721 = ~n56417 & n56438;
  assign n56722 = ~n56720 & ~n56721;
  assign n56723 = ~n56719 & n56722;
  assign n56724 = n56718 & ~n56723;
  assign n56725 = ~n56429 & n56461;
  assign n56726 = n56417 & n56725;
  assign n56727 = ~n56442 & ~n56726;
  assign n56728 = n56429 & n56452;
  assign n56729 = ~n56439 & ~n56728;
  assign n56730 = n56727 & n56729;
  assign n56731 = n56411 & ~n56730;
  assign n56732 = n56417 & n56469;
  assign n56733 = ~n56731 & ~n56732;
  assign n56734 = ~n56405 & ~n56733;
  assign n56735 = ~n56724 & ~n56734;
  assign n56736 = ~n56429 & n56473;
  assign n56737 = ~n56437 & n56736;
  assign n56738 = ~n56443 & ~n56737;
  assign n56739 = ~n56438 & ~n56461;
  assign n56740 = n56417 & ~n56739;
  assign n56741 = ~n56462 & ~n56740;
  assign n56742 = ~n56411 & ~n56741;
  assign n56743 = ~n56450 & ~n56719;
  assign n56744 = ~n56720 & n56743;
  assign n56745 = n56411 & ~n56744;
  assign n56746 = ~n56742 & ~n56745;
  assign n56747 = n56417 & n56462;
  assign n56748 = ~n56475 & ~n56747;
  assign n56749 = ~n56470 & n56748;
  assign n56750 = ~n56478 & n56749;
  assign n56751 = n56746 & n56750;
  assign n56752 = n56405 & ~n56751;
  assign n56753 = n56738 & ~n56752;
  assign n56754 = n56735 & n56753;
  assign n56755 = pi1577 & ~n56754;
  assign n56756 = ~pi1577 & n56738;
  assign n56757 = n56735 & n56756;
  assign n56758 = ~n56752 & n56757;
  assign po1667 = n56755 | n56758;
  assign n56760 = ~n56177 & ~n56206;
  assign n56761 = n56183 & n56760;
  assign n56762 = ~n56189 & n56218;
  assign n56763 = n56177 & n56762;
  assign n56764 = n56177 & n56227;
  assign n56765 = ~n56763 & ~n56764;
  assign n56766 = ~n56177 & n56189;
  assign n56767 = ~n56195 & n56766;
  assign n56768 = ~n56183 & n56767;
  assign n56769 = ~n56209 & ~n56768;
  assign n56770 = n56206 & ~n56769;
  assign n56771 = n56765 & ~n56770;
  assign n56772 = ~n56761 & n56771;
  assign n56773 = n56171 & ~n56772;
  assign n56774 = n56177 & n56248;
  assign n56775 = ~n56206 & n56774;
  assign n56776 = n56239 & n56248;
  assign n56777 = ~n56207 & ~n56776;
  assign n56778 = ~n56209 & ~n56242;
  assign n56779 = ~n56177 & n56226;
  assign n56780 = n56778 & ~n56779;
  assign n56781 = ~n56206 & ~n56780;
  assign n56782 = n56206 & n56213;
  assign n56783 = n56231 & ~n56782;
  assign n56784 = ~n56781 & n56783;
  assign n56785 = n56777 & n56784;
  assign n56786 = ~n56171 & ~n56785;
  assign n56787 = ~n56775 & ~n56786;
  assign n56788 = ~n56773 & n56787;
  assign n56789 = n56239 & n56242;
  assign n56790 = n56196 & n56206;
  assign n56791 = n56177 & n56790;
  assign n56792 = ~n56789 & ~n56791;
  assign n56793 = n56206 & n56764;
  assign n56794 = n56792 & ~n56793;
  assign n56795 = n56788 & n56794;
  assign n56796 = ~pi1580 & ~n56795;
  assign n56797 = pi1580 & n56794;
  assign n56798 = n56787 & n56797;
  assign n56799 = ~n56773 & n56798;
  assign po1668 = n56796 | n56799;
  assign n56801 = pi5069 & pi9040;
  assign n56802 = pi5315 & ~pi9040;
  assign n56803 = ~n56801 & ~n56802;
  assign n56804 = pi1555 & n56803;
  assign n56805 = ~pi1555 & ~n56803;
  assign n56806 = ~n56804 & ~n56805;
  assign n56807 = pi5089 & ~pi9040;
  assign n56808 = pi5152 & pi9040;
  assign n56809 = ~n56807 & ~n56808;
  assign n56810 = pi1524 & n56809;
  assign n56811 = ~pi1524 & ~n56809;
  assign n56812 = ~n56810 & ~n56811;
  assign n56813 = pi5071 & ~pi9040;
  assign n56814 = pi5416 & pi9040;
  assign n56815 = ~n56813 & ~n56814;
  assign n56816 = pi1544 & n56815;
  assign n56817 = ~pi1544 & ~n56815;
  assign n56818 = ~n56816 & ~n56817;
  assign n56819 = pi5267 & pi9040;
  assign n56820 = pi5144 & ~pi9040;
  assign n56821 = ~n56819 & ~n56820;
  assign n56822 = pi1545 & n56821;
  assign n56823 = ~pi1545 & ~n56821;
  assign n56824 = ~n56822 & ~n56823;
  assign n56825 = n56818 & ~n56824;
  assign n56826 = ~n56812 & n56825;
  assign n56827 = n56806 & n56826;
  assign n56828 = pi5154 & pi9040;
  assign n56829 = pi5252 & ~pi9040;
  assign n56830 = ~n56828 & ~n56829;
  assign n56831 = ~pi1549 & n56830;
  assign n56832 = pi1549 & ~n56830;
  assign n56833 = ~n56831 & ~n56832;
  assign n56834 = pi5073 & pi9040;
  assign n56835 = pi5196 & ~pi9040;
  assign n56836 = ~n56834 & ~n56835;
  assign n56837 = ~pi1554 & n56836;
  assign n56838 = pi1554 & ~n56836;
  assign n56839 = ~n56837 & ~n56838;
  assign n56840 = n56818 & ~n56839;
  assign n56841 = n56824 & n56840;
  assign n56842 = ~n56818 & ~n56839;
  assign n56843 = ~n56824 & n56842;
  assign n56844 = ~n56818 & n56839;
  assign n56845 = ~n56806 & n56844;
  assign n56846 = ~n56843 & ~n56845;
  assign n56847 = ~n56841 & n56846;
  assign n56848 = ~n56812 & ~n56847;
  assign n56849 = n56824 & n56842;
  assign n56850 = ~n56824 & n56840;
  assign n56851 = ~n56849 & ~n56850;
  assign n56852 = n56812 & ~n56851;
  assign n56853 = ~n56848 & ~n56852;
  assign n56854 = n56818 & n56839;
  assign n56855 = n56824 & n56854;
  assign n56856 = n56812 & n56855;
  assign n56857 = ~n56824 & n56845;
  assign n56858 = ~n56856 & ~n56857;
  assign n56859 = n56853 & n56858;
  assign n56860 = n56833 & ~n56859;
  assign n56861 = n56806 & n56849;
  assign n56862 = ~n56806 & n56854;
  assign n56863 = n56806 & n56844;
  assign n56864 = ~n56862 & ~n56863;
  assign n56865 = ~n56812 & ~n56864;
  assign n56866 = ~n56861 & ~n56865;
  assign n56867 = n56824 & n56844;
  assign n56868 = n56812 & n56867;
  assign n56869 = ~n56824 & n56854;
  assign n56870 = ~n56841 & ~n56869;
  assign n56871 = ~n56868 & n56870;
  assign n56872 = ~n56843 & n56871;
  assign n56873 = ~n56806 & ~n56872;
  assign n56874 = n56866 & ~n56873;
  assign n56875 = ~n56833 & ~n56874;
  assign n56876 = ~n56860 & ~n56875;
  assign n56877 = ~n56827 & n56876;
  assign n56878 = n56806 & n56824;
  assign n56879 = n56839 & n56878;
  assign n56880 = n56818 & n56879;
  assign n56881 = ~n56824 & n56863;
  assign n56882 = ~n56880 & ~n56881;
  assign n56883 = n56812 & ~n56882;
  assign n56884 = n56877 & ~n56883;
  assign n56885 = ~pi1597 & ~n56884;
  assign n56886 = pi1597 & ~n56883;
  assign n56887 = n56877 & n56886;
  assign po1669 = n56885 | n56887;
  assign n56889 = n56812 & n56849;
  assign n56890 = ~n56806 & n56889;
  assign n56891 = ~n56806 & n56812;
  assign n56892 = n56854 & n56891;
  assign n56893 = ~n56824 & n56892;
  assign n56894 = ~n56890 & ~n56893;
  assign n56895 = ~n56812 & n56843;
  assign n56896 = ~n56806 & n56895;
  assign n56897 = ~n56806 & n56869;
  assign n56898 = ~n56896 & ~n56897;
  assign n56899 = n56818 & n56824;
  assign n56900 = n56806 & n56899;
  assign n56901 = n56806 & n56842;
  assign n56902 = ~n56900 & ~n56901;
  assign n56903 = n56812 & ~n56902;
  assign n56904 = ~n56840 & ~n56844;
  assign n56905 = ~n56806 & ~n56824;
  assign n56906 = ~n56812 & ~n56905;
  assign n56907 = ~n56904 & n56906;
  assign n56908 = ~n56842 & n56891;
  assign n56909 = ~n56824 & n56908;
  assign n56910 = ~n56907 & ~n56909;
  assign n56911 = ~n56903 & n56910;
  assign n56912 = n56898 & n56911;
  assign n56913 = ~n56833 & ~n56912;
  assign n56914 = n56894 & ~n56913;
  assign n56915 = ~n56812 & n56841;
  assign n56916 = n56806 & n56915;
  assign n56917 = ~n56812 & n56833;
  assign n56918 = ~n56855 & ~n56901;
  assign n56919 = ~n56904 & n56905;
  assign n56920 = n56918 & ~n56919;
  assign n56921 = n56917 & ~n56920;
  assign n56922 = n56806 & n56869;
  assign n56923 = n56806 & n56818;
  assign n56924 = ~n56824 & n56923;
  assign n56925 = ~n56863 & ~n56924;
  assign n56926 = ~n56806 & n56842;
  assign n56927 = ~n56867 & ~n56926;
  assign n56928 = n56925 & n56927;
  assign n56929 = n56812 & ~n56928;
  assign n56930 = ~n56922 & ~n56929;
  assign n56931 = n56833 & ~n56930;
  assign n56932 = ~n56921 & ~n56931;
  assign n56933 = ~n56916 & n56932;
  assign n56934 = n56914 & n56933;
  assign n56935 = pi1581 & ~n56934;
  assign n56936 = ~pi1581 & n56914;
  assign n56937 = n56933 & n56936;
  assign po1670 = n56935 | n56937;
  assign n56939 = ~n56863 & ~n56926;
  assign n56940 = n56812 & ~n56939;
  assign n56941 = ~n56893 & ~n56940;
  assign n56942 = ~n56833 & ~n56941;
  assign n56943 = ~n56840 & n56878;
  assign n56944 = ~n56833 & n56943;
  assign n56945 = n56806 & ~n56824;
  assign n56946 = n56812 & n56945;
  assign n56947 = n56840 & n56946;
  assign n56948 = n56806 & ~n56812;
  assign n56949 = n56824 & n56839;
  assign n56950 = n56948 & n56949;
  assign n56951 = ~n56947 & ~n56950;
  assign n56952 = ~n56944 & n56951;
  assign n56953 = ~n56825 & ~n56840;
  assign n56954 = ~n56806 & ~n56953;
  assign n56955 = ~n56849 & ~n56954;
  assign n56956 = ~n56812 & ~n56955;
  assign n56957 = ~n56919 & ~n56956;
  assign n56958 = n56806 & n56843;
  assign n56959 = ~n56806 & n56824;
  assign n56960 = n56839 & n56959;
  assign n56961 = n56806 & ~n56953;
  assign n56962 = ~n56960 & ~n56961;
  assign n56963 = n56812 & ~n56962;
  assign n56964 = ~n56958 & ~n56963;
  assign n56965 = n56957 & n56964;
  assign n56966 = n56833 & ~n56965;
  assign n56967 = ~n56867 & ~n56923;
  assign n56968 = ~n56812 & ~n56833;
  assign n56969 = ~n56967 & n56968;
  assign n56970 = ~n56966 & ~n56969;
  assign n56971 = n56952 & n56970;
  assign n56972 = ~n56942 & n56971;
  assign n56973 = pi1587 & ~n56972;
  assign n56974 = ~pi1587 & n56972;
  assign po1671 = n56973 | n56974;
  assign n56976 = ~n56177 & n56762;
  assign n56977 = ~n56227 & ~n56235;
  assign n56978 = n56177 & n56196;
  assign n56979 = ~n56177 & n56248;
  assign n56980 = ~n56978 & ~n56979;
  assign n56981 = n56977 & n56980;
  assign n56982 = ~n56206 & ~n56981;
  assign n56983 = n56177 & n56208;
  assign n56984 = ~n56207 & ~n56983;
  assign n56985 = ~n56229 & n56984;
  assign n56986 = n56206 & ~n56985;
  assign n56987 = n56177 & n56209;
  assign n56988 = ~n56986 & ~n56987;
  assign n56989 = ~n56982 & n56988;
  assign n56990 = ~n56976 & n56989;
  assign n56991 = ~n56171 & ~n56990;
  assign n56992 = n56177 & ~n56206;
  assign n56993 = n56213 & n56992;
  assign n56994 = ~n56206 & n56229;
  assign n56995 = ~n56206 & n56242;
  assign n56996 = ~n56994 & ~n56995;
  assign n56997 = ~n56177 & ~n56996;
  assign n56998 = ~n56993 & ~n56997;
  assign n56999 = n56177 & n56226;
  assign n57000 = ~n56177 & n56208;
  assign n57001 = ~n56999 & ~n57000;
  assign n57002 = ~n56197 & n57001;
  assign n57003 = ~n56227 & n57002;
  assign n57004 = n56206 & ~n57003;
  assign n57005 = ~n56177 & n56209;
  assign n57006 = ~n57004 & ~n57005;
  assign n57007 = ~n56177 & n56197;
  assign n57008 = ~n56774 & ~n57007;
  assign n57009 = n57006 & n57008;
  assign n57010 = n56998 & n57009;
  assign n57011 = n56171 & ~n57010;
  assign n57012 = ~n56206 & ~n56765;
  assign n57013 = ~n57011 & ~n57012;
  assign n57014 = ~n56230 & ~n57007;
  assign n57015 = n56206 & ~n57014;
  assign n57016 = n57013 & ~n57015;
  assign n57017 = ~n56991 & n57016;
  assign n57018 = pi1583 & ~n57017;
  assign n57019 = ~pi1583 & n57017;
  assign po1672 = n57018 | n57019;
  assign n57021 = ~n56321 & ~n56329;
  assign n57022 = n56271 & ~n57021;
  assign n57023 = ~n56334 & ~n56511;
  assign n57024 = ~n56297 & n57023;
  assign n57025 = n56304 & ~n57024;
  assign n57026 = n56271 & n57025;
  assign n57027 = ~n57022 & ~n57026;
  assign n57028 = n56320 & n56514;
  assign n57029 = ~n56516 & ~n57028;
  assign n57030 = ~n56337 & ~n56542;
  assign n57031 = ~n56304 & ~n57030;
  assign n57032 = n56271 & n57031;
  assign n57033 = n57029 & ~n57032;
  assign n57034 = n56277 & n56320;
  assign n57035 = n56277 & n56312;
  assign n57036 = ~n56507 & ~n57035;
  assign n57037 = ~n56304 & ~n57036;
  assign n57038 = n56277 & n56319;
  assign n57039 = ~n56359 & ~n57038;
  assign n57040 = n56304 & ~n57039;
  assign n57041 = ~n56335 & ~n56519;
  assign n57042 = ~n57040 & n57041;
  assign n57043 = ~n57037 & n57042;
  assign n57044 = ~n57034 & n57043;
  assign n57045 = ~n56271 & ~n57044;
  assign n57046 = ~n56539 & n56559;
  assign n57047 = ~n56304 & ~n57046;
  assign n57048 = ~n57045 & ~n57047;
  assign n57049 = n57033 & n57048;
  assign n57050 = n57027 & n57049;
  assign n57051 = ~pi1589 & ~n57050;
  assign n57052 = pi1589 & n57033;
  assign n57053 = n57027 & n57052;
  assign n57054 = n57048 & n57053;
  assign po1673 = n57051 | n57054;
  assign n57056 = ~n56633 & ~n56651;
  assign n57057 = ~n56650 & n57056;
  assign n57058 = ~n56677 & ~n56691;
  assign n57059 = n57057 & ~n57058;
  assign n57060 = ~n56633 & n56658;
  assign n57061 = n56677 & n57060;
  assign n57062 = ~n57059 & ~n57061;
  assign n57063 = n56670 & ~n57062;
  assign n57064 = ~n56652 & n56675;
  assign n57065 = ~n56652 & ~n56658;
  assign n57066 = ~n56708 & ~n57065;
  assign n57067 = n56633 & ~n57066;
  assign n57068 = ~n56652 & n56658;
  assign n57069 = ~n56645 & n57068;
  assign n57070 = n56639 & n57069;
  assign n57071 = ~n57067 & ~n57070;
  assign n57072 = ~n57064 & n57071;
  assign n57073 = n56670 & ~n57072;
  assign n57074 = ~n57063 & ~n57073;
  assign n57075 = n56645 & n56659;
  assign n57076 = ~n56639 & n57075;
  assign n57077 = ~n56652 & n56684;
  assign n57078 = ~n57076 & ~n57077;
  assign n57079 = ~n56633 & ~n57078;
  assign n57080 = ~n56645 & n56661;
  assign n57081 = ~n56639 & n57080;
  assign n57082 = ~n56652 & n56708;
  assign n57083 = ~n57081 & ~n57082;
  assign n57084 = n56633 & ~n57083;
  assign n57085 = ~n56646 & ~n56708;
  assign n57086 = n56652 & ~n57085;
  assign n57087 = ~n56684 & ~n57086;
  assign n57088 = ~n56633 & ~n57087;
  assign n57089 = n56645 & ~n56652;
  assign n57090 = n57060 & n57089;
  assign n57091 = ~n56645 & ~n56658;
  assign n57092 = ~n56684 & ~n57091;
  assign n57093 = ~n56652 & ~n57092;
  assign n57094 = n56633 & n56652;
  assign n57095 = n56674 & n57094;
  assign n57096 = n56658 & n57095;
  assign n57097 = ~n57093 & ~n57096;
  assign n57098 = ~n57090 & n57097;
  assign n57099 = ~n57088 & n57098;
  assign n57100 = ~n57076 & n57099;
  assign n57101 = ~n56670 & ~n57100;
  assign n57102 = ~n57084 & ~n57101;
  assign n57103 = ~n57079 & n57102;
  assign n57104 = n57074 & n57103;
  assign n57105 = pi1578 & n57104;
  assign n57106 = ~pi1578 & ~n57104;
  assign po1674 = n57105 | n57106;
  assign n57108 = ~n55980 & n55991;
  assign n57109 = ~n56595 & ~n57108;
  assign n57110 = n55972 & ~n57109;
  assign n57111 = n56013 & n56045;
  assign n57112 = ~n57110 & ~n57111;
  assign n57113 = ~n56060 & n57112;
  assign n57114 = n55966 & ~n55972;
  assign n57115 = n55989 & n57114;
  assign n57116 = ~n55960 & n57115;
  assign n57117 = ~n55980 & n57116;
  assign n57118 = ~n55972 & n56606;
  assign n57119 = ~n56040 & ~n56053;
  assign n57120 = ~n56025 & n57119;
  assign n57121 = ~n57118 & n57120;
  assign n57122 = n56011 & ~n57121;
  assign n57123 = n55980 & n56002;
  assign n57124 = ~n57116 & ~n57123;
  assign n57125 = ~n56594 & n57124;
  assign n57126 = n55989 & n56038;
  assign n57127 = n55980 & n56032;
  assign n57128 = ~n56044 & ~n57127;
  assign n57129 = n55972 & ~n57128;
  assign n57130 = ~n57126 & ~n57129;
  assign n57131 = n57125 & n57130;
  assign n57132 = ~n56011 & ~n57131;
  assign n57133 = n55980 & n55994;
  assign n57134 = ~n55991 & ~n57133;
  assign n57135 = ~n56604 & n57134;
  assign n57136 = n55972 & ~n57135;
  assign n57137 = n56011 & n57136;
  assign n57138 = ~n57132 & ~n57137;
  assign n57139 = ~n57122 & n57138;
  assign n57140 = ~n57117 & n57139;
  assign n57141 = n57113 & n57140;
  assign n57142 = pi1596 & ~n57141;
  assign n57143 = ~pi1596 & n57113;
  assign n57144 = n57140 & n57143;
  assign po1675 = n57142 | n57144;
  assign n57146 = ~n56839 & n56959;
  assign n57147 = n56870 & ~n57146;
  assign n57148 = n56968 & ~n57147;
  assign n57149 = ~n56833 & n56867;
  assign n57150 = n56806 & n57149;
  assign n57151 = ~n56824 & ~n56839;
  assign n57152 = ~n56901 & ~n57151;
  assign n57153 = n56812 & ~n57152;
  assign n57154 = ~n56856 & ~n57153;
  assign n57155 = ~n56833 & ~n57154;
  assign n57156 = ~n57150 & ~n57155;
  assign n57157 = ~n56839 & n56945;
  assign n57158 = ~n56857 & ~n57157;
  assign n57159 = n56812 & ~n57158;
  assign n57160 = n57156 & ~n57159;
  assign n57161 = ~n56904 & n56959;
  assign n57162 = n56842 & n56948;
  assign n57163 = n56824 & n57162;
  assign n57164 = ~n56904 & n56945;
  assign n57165 = n56824 & n56891;
  assign n57166 = ~n56818 & n57165;
  assign n57167 = ~n57164 & ~n57166;
  assign n57168 = ~n57163 & n57167;
  assign n57169 = ~n57161 & n57168;
  assign n57170 = ~n56880 & n56898;
  assign n57171 = n57169 & n57170;
  assign n57172 = n56833 & ~n57171;
  assign n57173 = n57160 & ~n57172;
  assign n57174 = ~n57148 & n57173;
  assign n57175 = ~pi1586 & ~n57174;
  assign n57176 = pi1586 & n57160;
  assign n57177 = ~n57148 & n57176;
  assign n57178 = ~n57172 & n57177;
  assign po1676 = n57175 | n57178;
  assign n57180 = n55875 & n55897;
  assign n57181 = ~n56389 & ~n57180;
  assign n57182 = n55881 & n57181;
  assign n57183 = ~n55875 & n55934;
  assign n57184 = ~n55891 & ~n55909;
  assign n57185 = ~n55890 & ~n57184;
  assign n57186 = n55863 & n55904;
  assign n57187 = ~n55875 & n55891;
  assign n57188 = ~n57186 & ~n57187;
  assign n57189 = ~n55881 & n57188;
  assign n57190 = ~n57185 & n57189;
  assign n57191 = ~n57183 & n57190;
  assign n57192 = ~n57182 & ~n57191;
  assign n57193 = ~n55875 & n57185;
  assign n57194 = ~n56378 & ~n57193;
  assign n57195 = ~n57192 & n57194;
  assign n57196 = n55857 & ~n57195;
  assign n57197 = n55881 & ~n57184;
  assign n57198 = n55875 & n57197;
  assign n57199 = ~n55912 & ~n55938;
  assign n57200 = ~n55875 & ~n57199;
  assign n57201 = n55881 & n57200;
  assign n57202 = n55890 & n57197;
  assign n57203 = ~n57201 & ~n57202;
  assign n57204 = ~n57198 & n57203;
  assign n57205 = ~n55857 & ~n57204;
  assign n57206 = ~n57196 & ~n57205;
  assign n57207 = n55881 & n55895;
  assign n57208 = ~n55881 & ~n57194;
  assign n57209 = ~n57207 & ~n57208;
  assign n57210 = ~n55881 & ~n57181;
  assign n57211 = ~n55895 & ~n57210;
  assign n57212 = ~n55857 & ~n57211;
  assign n57213 = n57209 & ~n57212;
  assign n57214 = n57206 & n57213;
  assign n57215 = pi1595 & ~n57214;
  assign n57216 = ~pi1595 & n57213;
  assign n57217 = ~n57205 & n57216;
  assign n57218 = ~n57196 & n57217;
  assign po1677 = n57215 | n57218;
  assign n57220 = ~n56097 & n56126;
  assign n57221 = ~n56089 & n56097;
  assign n57222 = n56077 & n57221;
  assign n57223 = ~n56123 & ~n57222;
  assign n57224 = n56071 & ~n57223;
  assign n57225 = ~n57220 & ~n57224;
  assign n57226 = ~n56071 & ~n56097;
  assign n57227 = ~n56089 & n57226;
  assign n57228 = ~n56083 & n57227;
  assign n57229 = n56105 & n56138;
  assign n57230 = ~n57228 & ~n57229;
  assign n57231 = ~n56071 & ~n56077;
  assign n57232 = n56099 & n57231;
  assign n57233 = n57230 & ~n57232;
  assign n57234 = ~n56101 & ~n56113;
  assign n57235 = n56089 & n56144;
  assign n57236 = n57234 & ~n57235;
  assign n57237 = n57233 & n57236;
  assign n57238 = n57225 & n57237;
  assign n57239 = ~n56135 & ~n57238;
  assign n57240 = ~n56100 & ~n56123;
  assign n57241 = n56097 & ~n57240;
  assign n57242 = ~n56083 & n56141;
  assign n57243 = ~n56152 & ~n57242;
  assign n57244 = ~n56077 & ~n56089;
  assign n57245 = n56097 & n57244;
  assign n57246 = n57243 & ~n57245;
  assign n57247 = n56071 & ~n57246;
  assign n57248 = ~n56097 & n56111;
  assign n57249 = n56077 & n56097;
  assign n57250 = ~n56089 & n57249;
  assign n57251 = ~n56083 & n57250;
  assign n57252 = ~n57248 & ~n57251;
  assign n57253 = ~n56071 & ~n57252;
  assign n57254 = ~n56097 & n56106;
  assign n57255 = ~n57253 & ~n57254;
  assign n57256 = ~n57247 & n57255;
  assign n57257 = ~n57241 & n57256;
  assign n57258 = n56135 & ~n57257;
  assign n57259 = n56071 & n56142;
  assign n57260 = ~n57258 & ~n57259;
  assign n57261 = n56118 & n57226;
  assign n57262 = ~n56089 & n57261;
  assign n57263 = n57260 & ~n57262;
  assign n57264 = ~n57239 & n57263;
  assign n57265 = ~pi1590 & ~n57264;
  assign n57266 = pi1590 & n57260;
  assign n57267 = ~n57239 & n57266;
  assign n57268 = ~n57262 & n57267;
  assign po1679 = n57265 | n57268;
  assign n57270 = n56411 & n56438;
  assign n57271 = ~n56417 & n57270;
  assign n57272 = ~n56495 & ~n57271;
  assign n57273 = n56417 & ~n56437;
  assign n57274 = ~n56429 & n57273;
  assign n57275 = ~n56417 & n56423;
  assign n57276 = ~n56494 & ~n57275;
  assign n57277 = ~n56411 & ~n57276;
  assign n57278 = ~n57274 & ~n57277;
  assign n57279 = n57272 & n57278;
  assign n57280 = n56405 & ~n57279;
  assign n57281 = ~n56417 & n56449;
  assign n57282 = ~n56465 & ~n56475;
  assign n57283 = ~n57281 & n57282;
  assign n57284 = n56411 & ~n57283;
  assign n57285 = n56438 & n56477;
  assign n57286 = ~n56443 & ~n57285;
  assign n57287 = ~n57284 & n57286;
  assign n57288 = ~n56725 & ~n56732;
  assign n57289 = ~n56411 & ~n57288;
  assign n57290 = n57287 & ~n57289;
  assign n57291 = ~n56405 & ~n57290;
  assign n57292 = ~n57280 & ~n57291;
  assign n57293 = ~n56417 & n56461;
  assign n57294 = n56417 & ~n56729;
  assign n57295 = ~n57293 & ~n57294;
  assign n57296 = ~n56411 & ~n57295;
  assign n57297 = ~n56450 & ~n56462;
  assign n57298 = ~n56465 & n57297;
  assign n57299 = n56484 & ~n57298;
  assign n57300 = ~n57296 & ~n57299;
  assign n57301 = n57292 & n57300;
  assign n57302 = ~pi1585 & ~n57301;
  assign n57303 = ~n57291 & n57300;
  assign n57304 = pi1585 & n57303;
  assign n57305 = ~n57280 & n57304;
  assign po1680 = n57302 | n57305;
  assign n57307 = ~n56411 & ~n57297;
  assign n57308 = n56417 & n56439;
  assign n57309 = ~n57307 & ~n57308;
  assign n57310 = n56417 & ~n56423;
  assign n57311 = ~n56446 & ~n57310;
  assign n57312 = ~n56725 & n57311;
  assign n57313 = n56411 & ~n57312;
  assign n57314 = n57309 & ~n57313;
  assign n57315 = ~n56405 & ~n57314;
  assign n57316 = ~n56411 & n56448;
  assign n57317 = ~n56467 & ~n57316;
  assign n57318 = ~n56471 & n57317;
  assign n57319 = ~n56470 & ~n56494;
  assign n57320 = n56411 & n56480;
  assign n57321 = n56417 & n56450;
  assign n57322 = ~n56411 & n56446;
  assign n57323 = ~n57321 & ~n57322;
  assign n57324 = ~n56747 & n57323;
  assign n57325 = ~n57320 & n57324;
  assign n57326 = n57319 & n57325;
  assign n57327 = ~n56487 & n57326;
  assign n57328 = n56405 & ~n57327;
  assign n57329 = n57318 & ~n57328;
  assign n57330 = ~n57315 & n57329;
  assign n57331 = ~pi1592 & ~n57330;
  assign n57332 = pi1592 & n57318;
  assign n57333 = ~n57315 & n57332;
  assign n57334 = ~n57328 & n57333;
  assign po1681 = n57331 | n57334;
  assign n57336 = ~n56098 & ~n56104;
  assign n57337 = ~n56071 & ~n57336;
  assign n57338 = ~n56159 & ~n57337;
  assign n57339 = n56077 & n56083;
  assign n57340 = n56071 & n57339;
  assign n57341 = n56097 & n57340;
  assign n57342 = n56097 & n56111;
  assign n57343 = ~n57339 & ~n57342;
  assign n57344 = ~n56077 & ~n56097;
  assign n57345 = ~n56083 & n57344;
  assign n57346 = n57343 & ~n57345;
  assign n57347 = n56071 & ~n57346;
  assign n57348 = ~n56107 & ~n57347;
  assign n57349 = ~n56135 & ~n57348;
  assign n57350 = ~n56071 & n56090;
  assign n57351 = n56097 & n57350;
  assign n57352 = ~n57232 & ~n57351;
  assign n57353 = ~n56135 & ~n57352;
  assign n57354 = ~n57349 & ~n57353;
  assign n57355 = ~n57341 & n57354;
  assign n57356 = ~n56123 & ~n56142;
  assign n57357 = ~n56152 & n57356;
  assign n57358 = ~n56071 & ~n57357;
  assign n57359 = n56099 & n57344;
  assign n57360 = ~n56126 & ~n57359;
  assign n57361 = n56071 & ~n57360;
  assign n57362 = ~n57358 & ~n57361;
  assign n57363 = ~n57242 & n57362;
  assign n57364 = ~n56113 & ~n56153;
  assign n57365 = n57363 & n57364;
  assign n57366 = n56135 & ~n57365;
  assign n57367 = n57355 & ~n57366;
  assign n57368 = n57338 & n57367;
  assign n57369 = ~pi1606 & ~n57368;
  assign n57370 = pi1606 & n57355;
  assign n57371 = n57338 & n57370;
  assign n57372 = ~n57366 & n57371;
  assign po1682 = n57369 | n57372;
  assign n57374 = ~n55875 & n56380;
  assign n57375 = n55881 & n57374;
  assign n57376 = n55904 & ~n57184;
  assign n57377 = ~n55939 & ~n57376;
  assign n57378 = ~n56378 & n57377;
  assign n57379 = ~n55881 & ~n57378;
  assign n57380 = ~n55875 & n55892;
  assign n57381 = ~n57379 & ~n57380;
  assign n57382 = n55890 & n55938;
  assign n57383 = n55875 & n56384;
  assign n57384 = ~n57382 & ~n57383;
  assign n57385 = ~n57187 & n57384;
  assign n57386 = n55881 & ~n57385;
  assign n57387 = n57381 & ~n57386;
  assign n57388 = n55857 & ~n57387;
  assign n57389 = ~n57375 & ~n57388;
  assign n57390 = n55875 & n55891;
  assign n57391 = ~n55917 & ~n57390;
  assign n57392 = n55881 & ~n57391;
  assign n57393 = ~n55940 & ~n57392;
  assign n57394 = ~n55913 & ~n57374;
  assign n57395 = ~n55875 & n55946;
  assign n57396 = ~n56384 & ~n57395;
  assign n57397 = ~n57382 & n57396;
  assign n57398 = ~n55881 & ~n57397;
  assign n57399 = n55875 & n55892;
  assign n57400 = ~n57398 & ~n57399;
  assign n57401 = n57394 & n57400;
  assign n57402 = n57393 & n57401;
  assign n57403 = ~n55857 & ~n57402;
  assign n57404 = ~n55926 & ~n57183;
  assign n57405 = ~n55881 & ~n57404;
  assign n57406 = ~n57403 & ~n57405;
  assign n57407 = n57389 & n57406;
  assign n57408 = pi1594 & n57407;
  assign n57409 = ~pi1594 & ~n57407;
  assign po1683 = n57408 | n57409;
  assign n57411 = n55980 & n56618;
  assign n57412 = ~n55993 & ~n56606;
  assign n57413 = n55972 & ~n57412;
  assign n57414 = ~n57411 & ~n57413;
  assign n57415 = n55989 & n56593;
  assign n57416 = ~n55999 & ~n57415;
  assign n57417 = ~n56604 & n57416;
  assign n57418 = ~n55972 & ~n57417;
  assign n57419 = n57414 & ~n57418;
  assign n57420 = ~n55980 & n56045;
  assign n57421 = n57419 & ~n57420;
  assign n57422 = ~n56011 & ~n57421;
  assign n57423 = n56058 & ~n57412;
  assign n57424 = ~n55991 & ~n55994;
  assign n57425 = ~n56045 & ~n56604;
  assign n57426 = n57424 & n57425;
  assign n57427 = n55980 & ~n57426;
  assign n57428 = ~n57423 & ~n57427;
  assign n57429 = ~n56595 & n57428;
  assign n57430 = n56011 & ~n57429;
  assign n57431 = ~n57422 & ~n57430;
  assign n57432 = n55980 & n56606;
  assign n57433 = ~n57420 & ~n57432;
  assign n57434 = n55972 & ~n57433;
  assign n57435 = n57431 & ~n57434;
  assign n57436 = pi1574 & ~n57435;
  assign n57437 = ~pi1574 & ~n57434;
  assign n57438 = ~n57430 & n57437;
  assign n57439 = ~n57422 & n57438;
  assign po1685 = n57436 | n57439;
  assign n57441 = n56646 & n57065;
  assign n57442 = n56700 & ~n57441;
  assign n57443 = n56633 & ~n57442;
  assign n57444 = ~n56652 & n56688;
  assign n57445 = ~n57443 & ~n57444;
  assign n57446 = n56639 & n56661;
  assign n57447 = n56652 & n56674;
  assign n57448 = ~n57446 & ~n57447;
  assign n57449 = n56633 & ~n57448;
  assign n57450 = n56633 & n56683;
  assign n57451 = ~n56652 & n57450;
  assign n57452 = ~n57449 & ~n57451;
  assign n57453 = n57445 & n57452;
  assign n57454 = ~n56670 & ~n57453;
  assign n57455 = ~n56678 & ~n56685;
  assign n57456 = ~n57070 & n57455;
  assign n57457 = n56705 & ~n57456;
  assign n57458 = ~n57454 & ~n57457;
  assign n57459 = ~n56652 & n56678;
  assign n57460 = ~n57090 & ~n57459;
  assign n57461 = ~n56691 & ~n57080;
  assign n57462 = ~n56633 & ~n57461;
  assign n57463 = n56652 & n56683;
  assign n57464 = ~n57069 & ~n57463;
  assign n57465 = n56633 & ~n57464;
  assign n57466 = ~n57462 & ~n57465;
  assign n57467 = ~n56660 & n57466;
  assign n57468 = n57460 & n57467;
  assign n57469 = ~n57064 & ~n57076;
  assign n57470 = n57468 & n57469;
  assign n57471 = n56670 & ~n57470;
  assign n57472 = ~n56660 & ~n57064;
  assign n57473 = ~n56633 & ~n57472;
  assign n57474 = ~n57471 & ~n57473;
  assign n57475 = n57458 & n57474;
  assign n57476 = ~pi1579 & n57475;
  assign n57477 = pi1579 & ~n57475;
  assign po1686 = n57476 | n57477;
  assign n57479 = ~n56768 & ~n57007;
  assign n57480 = ~n56987 & n57479;
  assign n57481 = ~n56206 & ~n57480;
  assign n57482 = ~n56776 & ~n56793;
  assign n57483 = ~n56774 & ~n56995;
  assign n57484 = ~n56762 & ~n57000;
  assign n57485 = n56206 & ~n57484;
  assign n57486 = ~n56235 & ~n57485;
  assign n57487 = n57483 & n57486;
  assign n57488 = n56171 & ~n57487;
  assign n57489 = n56189 & n56195;
  assign n57490 = ~n56214 & ~n57489;
  assign n57491 = n56177 & ~n57490;
  assign n57492 = ~n56197 & ~n56779;
  assign n57493 = n56206 & ~n57492;
  assign n57494 = n56177 & n56195;
  assign n57495 = ~n56209 & ~n57494;
  assign n57496 = ~n56218 & n57495;
  assign n57497 = ~n56206 & ~n57496;
  assign n57498 = ~n57493 & ~n57497;
  assign n57499 = ~n57491 & n57498;
  assign n57500 = ~n56171 & ~n57499;
  assign n57501 = ~n57488 & ~n57500;
  assign n57502 = n57482 & n57501;
  assign n57503 = ~n57481 & n57502;
  assign n57504 = ~pi1601 & ~n57503;
  assign n57505 = pi1601 & n57482;
  assign n57506 = ~n57481 & n57505;
  assign n57507 = n57501 & n57506;
  assign po1687 = n57504 | n57507;
  assign n57509 = ~n56153 & ~n57254;
  assign n57510 = n56071 & ~n57509;
  assign n57511 = ~n56135 & n56137;
  assign n57512 = ~n56071 & n57511;
  assign n57513 = n56083 & n57344;
  assign n57514 = ~n57244 & ~n57513;
  assign n57515 = ~n56106 & n57514;
  assign n57516 = n56071 & ~n57515;
  assign n57517 = ~n56097 & n56112;
  assign n57518 = ~n57516 & ~n57517;
  assign n57519 = ~n56135 & ~n57518;
  assign n57520 = ~n57512 & ~n57519;
  assign n57521 = ~n56101 & ~n56104;
  assign n57522 = ~n56097 & n56152;
  assign n57523 = ~n57222 & ~n57522;
  assign n57524 = n57521 & n57523;
  assign n57525 = ~n56071 & ~n57524;
  assign n57526 = n56077 & ~n56083;
  assign n57527 = ~n56071 & n57526;
  assign n57528 = n56097 & n57527;
  assign n57529 = ~n56097 & n57244;
  assign n57530 = ~n56104 & ~n57529;
  assign n57531 = ~n57251 & n57530;
  assign n57532 = ~n57528 & n57531;
  assign n57533 = n56071 & n56100;
  assign n57534 = n57532 & ~n57533;
  assign n57535 = n56135 & ~n57534;
  assign n57536 = ~n57525 & ~n57535;
  assign n57537 = n57520 & n57536;
  assign n57538 = ~n57510 & n57537;
  assign n57539 = pi1619 & n57538;
  assign n57540 = ~pi1619 & ~n57538;
  assign po1688 = n57539 | n57540;
  assign n57542 = ~n56652 & n56674;
  assign n57543 = ~n56673 & ~n57542;
  assign n57544 = ~n56633 & ~n57543;
  assign n57545 = n56633 & ~n57092;
  assign n57546 = ~n57081 & ~n57545;
  assign n57547 = ~n57544 & n57546;
  assign n57548 = n56670 & ~n57547;
  assign n57549 = ~n56633 & n56688;
  assign n57550 = ~n57548 & ~n57549;
  assign n57551 = ~n57447 & ~n57459;
  assign n57552 = n56633 & ~n57551;
  assign n57553 = n56633 & n56675;
  assign n57554 = n56652 & n56691;
  assign n57555 = ~n56658 & n57057;
  assign n57556 = ~n57068 & ~n57555;
  assign n57557 = ~n56639 & ~n57556;
  assign n57558 = ~n57069 & ~n57557;
  assign n57559 = ~n56660 & n57558;
  assign n57560 = ~n57554 & n57559;
  assign n57561 = ~n57553 & n57560;
  assign n57562 = ~n56670 & ~n57561;
  assign n57563 = ~n57552 & ~n57562;
  assign n57564 = n57550 & n57563;
  assign n57565 = pi1602 & ~n57564;
  assign n57566 = ~pi1602 & n57564;
  assign po1689 = n57565 | n57566;
  assign n57568 = pi5402 & ~pi9040;
  assign n57569 = pi5570 & pi9040;
  assign n57570 = ~n57568 & ~n57569;
  assign n57571 = ~pi1611 & ~n57570;
  assign n57572 = pi1611 & n57570;
  assign n57573 = ~n57571 & ~n57572;
  assign n57574 = pi5400 & pi9040;
  assign n57575 = pi5401 & ~pi9040;
  assign n57576 = ~n57574 & ~n57575;
  assign n57577 = pi1624 & n57576;
  assign n57578 = ~pi1624 & ~n57576;
  assign n57579 = ~n57577 & ~n57578;
  assign n57580 = pi5396 & pi9040;
  assign n57581 = pi5510 & ~pi9040;
  assign n57582 = ~n57580 & ~n57581;
  assign n57583 = ~pi1598 & ~n57582;
  assign n57584 = pi1598 & ~n57580;
  assign n57585 = ~n57581 & n57584;
  assign n57586 = ~n57583 & ~n57585;
  assign n57587 = pi5514 & pi9040;
  assign n57588 = pi5317 & ~pi9040;
  assign n57589 = ~n57587 & ~n57588;
  assign n57590 = ~pi1621 & ~n57589;
  assign n57591 = pi1621 & n57589;
  assign n57592 = ~n57590 & ~n57591;
  assign n57593 = pi5407 & ~pi9040;
  assign n57594 = pi5513 & pi9040;
  assign n57595 = ~n57593 & ~n57594;
  assign n57596 = ~pi1612 & n57595;
  assign n57597 = pi1612 & ~n57595;
  assign n57598 = ~n57596 & ~n57597;
  assign n57599 = n57592 & n57598;
  assign n57600 = n57586 & n57599;
  assign n57601 = pi5509 & pi9040;
  assign n57602 = pi5443 & ~pi9040;
  assign n57603 = ~n57601 & ~n57602;
  assign n57604 = ~pi1593 & ~n57603;
  assign n57605 = pi1593 & n57603;
  assign n57606 = ~n57604 & ~n57605;
  assign n57607 = ~n57598 & n57606;
  assign n57608 = n57592 & n57607;
  assign n57609 = ~n57600 & ~n57608;
  assign n57610 = ~n57598 & ~n57606;
  assign n57611 = ~n57592 & n57610;
  assign n57612 = ~n57586 & n57611;
  assign n57613 = n57609 & ~n57612;
  assign n57614 = n57579 & ~n57613;
  assign n57615 = ~n57592 & ~n57598;
  assign n57616 = n57606 & n57615;
  assign n57617 = ~n57586 & n57616;
  assign n57618 = n57598 & n57606;
  assign n57619 = n57592 & n57618;
  assign n57620 = ~n57586 & n57619;
  assign n57621 = ~n57592 & n57598;
  assign n57622 = ~n57610 & ~n57621;
  assign n57623 = n57586 & ~n57622;
  assign n57624 = ~n57620 & ~n57623;
  assign n57625 = ~n57617 & n57624;
  assign n57626 = ~n57579 & ~n57625;
  assign n57627 = ~n57614 & ~n57626;
  assign n57628 = n57573 & ~n57627;
  assign n57629 = n57579 & ~n57586;
  assign n57630 = n57598 & n57629;
  assign n57631 = ~n57579 & ~n57586;
  assign n57632 = n57610 & n57631;
  assign n57633 = ~n57586 & ~n57598;
  assign n57634 = n57592 & n57633;
  assign n57635 = ~n57600 & ~n57634;
  assign n57636 = ~n57579 & ~n57635;
  assign n57637 = ~n57632 & ~n57636;
  assign n57638 = n57592 & n57610;
  assign n57639 = ~n57586 & n57638;
  assign n57640 = n57586 & n57616;
  assign n57641 = ~n57639 & ~n57640;
  assign n57642 = n57579 & n57586;
  assign n57643 = n57615 & n57642;
  assign n57644 = ~n57592 & n57618;
  assign n57645 = n57579 & n57644;
  assign n57646 = ~n57643 & ~n57645;
  assign n57647 = n57641 & n57646;
  assign n57648 = n57637 & n57647;
  assign n57649 = ~n57630 & n57648;
  assign n57650 = ~n57573 & ~n57649;
  assign n57651 = n57598 & ~n57606;
  assign n57652 = ~n57592 & n57651;
  assign n57653 = ~n57579 & n57652;
  assign n57654 = ~n57586 & n57653;
  assign n57655 = ~n57579 & n57639;
  assign n57656 = ~n57654 & ~n57655;
  assign n57657 = ~n57586 & ~n57592;
  assign n57658 = n57606 & n57657;
  assign n57659 = n57598 & n57658;
  assign n57660 = n57579 & n57659;
  assign n57661 = n57656 & ~n57660;
  assign n57662 = n57599 & ~n57606;
  assign n57663 = ~n57586 & n57662;
  assign n57664 = n57586 & n57607;
  assign n57665 = ~n57663 & ~n57664;
  assign n57666 = n57579 & ~n57665;
  assign n57667 = n57661 & ~n57666;
  assign n57668 = ~n57650 & n57667;
  assign n57669 = ~n57628 & n57668;
  assign n57670 = ~pi1656 & ~n57669;
  assign n57671 = pi1656 & n57669;
  assign po1710 = n57670 | n57671;
  assign n57673 = ~n57573 & ~n57579;
  assign n57674 = ~n57586 & n57599;
  assign n57675 = n57586 & n57638;
  assign n57676 = ~n57586 & n57607;
  assign n57677 = ~n57675 & ~n57676;
  assign n57678 = ~n57674 & n57677;
  assign n57679 = n57673 & ~n57678;
  assign n57680 = ~n57606 & n57657;
  assign n57681 = n57586 & n57662;
  assign n57682 = ~n57680 & ~n57681;
  assign n57683 = ~n57608 & ~n57611;
  assign n57684 = n57682 & n57683;
  assign n57685 = n57579 & ~n57684;
  assign n57686 = n57586 & n57644;
  assign n57687 = ~n57685 & ~n57686;
  assign n57688 = ~n57573 & ~n57687;
  assign n57689 = ~n57679 & ~n57688;
  assign n57690 = n57592 & n57629;
  assign n57691 = n57606 & n57690;
  assign n57692 = ~n57612 & ~n57691;
  assign n57693 = ~n57607 & ~n57651;
  assign n57694 = n57586 & ~n57693;
  assign n57695 = ~n57652 & ~n57694;
  assign n57696 = ~n57579 & ~n57695;
  assign n57697 = ~n57619 & ~n57674;
  assign n57698 = ~n57675 & n57697;
  assign n57699 = n57579 & ~n57698;
  assign n57700 = ~n57696 & ~n57699;
  assign n57701 = n57586 & ~n57592;
  assign n57702 = ~n57606 & n57701;
  assign n57703 = n57598 & n57702;
  assign n57704 = ~n57640 & ~n57703;
  assign n57705 = ~n57659 & n57704;
  assign n57706 = ~n57632 & n57705;
  assign n57707 = n57700 & n57706;
  assign n57708 = n57573 & ~n57707;
  assign n57709 = n57692 & ~n57708;
  assign n57710 = n57689 & n57709;
  assign n57711 = pi1646 & ~n57710;
  assign n57712 = ~pi1646 & n57692;
  assign n57713 = n57689 & n57712;
  assign n57714 = ~n57708 & n57713;
  assign po1714 = n57711 | n57714;
  assign n57716 = pi5441 & pi9040;
  assign n57717 = pi5435 & ~pi9040;
  assign n57718 = ~n57716 & ~n57717;
  assign n57719 = ~pi1603 & ~n57718;
  assign n57720 = pi1603 & n57718;
  assign n57721 = ~n57719 & ~n57720;
  assign n57722 = pi5511 & ~pi9040;
  assign n57723 = pi5438 & pi9040;
  assign n57724 = ~n57722 & ~n57723;
  assign n57725 = pi1608 & n57724;
  assign n57726 = ~pi1608 & ~n57724;
  assign n57727 = ~n57725 & ~n57726;
  assign n57728 = pi5392 & ~pi9040;
  assign n57729 = pi5402 & pi9040;
  assign n57730 = ~n57728 & ~n57729;
  assign n57731 = ~pi1620 & n57730;
  assign n57732 = pi1620 & ~n57730;
  assign n57733 = ~n57731 & ~n57732;
  assign n57734 = pi5316 & pi9040;
  assign n57735 = pi5400 & ~pi9040;
  assign n57736 = ~n57734 & ~n57735;
  assign n57737 = ~pi1600 & n57736;
  assign n57738 = pi1600 & ~n57736;
  assign n57739 = ~n57737 & ~n57738;
  assign n57740 = ~n57733 & ~n57739;
  assign n57741 = ~n57727 & n57740;
  assign n57742 = pi5320 & ~pi9040;
  assign n57743 = pi5510 & pi9040;
  assign n57744 = ~n57742 & ~n57743;
  assign n57745 = pi1617 & n57744;
  assign n57746 = ~pi1617 & ~n57744;
  assign n57747 = ~n57745 & ~n57746;
  assign n57748 = n57741 & ~n57747;
  assign n57749 = ~pi1600 & ~n57736;
  assign n57750 = pi1600 & n57736;
  assign n57751 = ~n57749 & ~n57750;
  assign n57752 = n57733 & ~n57751;
  assign n57753 = ~n57727 & n57752;
  assign n57754 = ~n57747 & n57753;
  assign n57755 = ~n57748 & ~n57754;
  assign n57756 = n57727 & n57752;
  assign n57757 = n57747 & n57756;
  assign n57758 = ~n57733 & ~n57751;
  assign n57759 = ~n57727 & n57758;
  assign n57760 = n57747 & n57759;
  assign n57761 = ~n57757 & ~n57760;
  assign n57762 = n57755 & n57761;
  assign n57763 = n57721 & ~n57762;
  assign n57764 = ~n57727 & n57747;
  assign n57765 = ~n57739 & n57764;
  assign n57766 = n57733 & n57765;
  assign n57767 = ~n57759 & ~n57766;
  assign n57768 = n57721 & ~n57767;
  assign n57769 = ~n57721 & ~n57739;
  assign n57770 = ~n57747 & n57769;
  assign n57771 = n57727 & ~n57733;
  assign n57772 = n57747 & n57752;
  assign n57773 = ~n57771 & ~n57772;
  assign n57774 = ~n57721 & ~n57773;
  assign n57775 = ~n57770 & ~n57774;
  assign n57776 = n57733 & ~n57739;
  assign n57777 = n57727 & n57776;
  assign n57778 = ~n57747 & n57777;
  assign n57779 = n57775 & ~n57778;
  assign n57780 = n57751 & n57771;
  assign n57781 = n57747 & n57780;
  assign n57782 = n57779 & ~n57781;
  assign n57783 = ~n57768 & n57782;
  assign n57784 = pi5407 & pi9040;
  assign n57785 = pi5308 & ~pi9040;
  assign n57786 = ~n57784 & ~n57785;
  assign n57787 = pi1628 & n57786;
  assign n57788 = ~pi1628 & ~n57786;
  assign n57789 = ~n57787 & ~n57788;
  assign n57790 = ~n57783 & ~n57789;
  assign n57791 = ~n57727 & ~n57739;
  assign n57792 = ~n57721 & n57747;
  assign n57793 = n57789 & n57792;
  assign n57794 = n57791 & n57793;
  assign n57795 = ~n57727 & ~n57747;
  assign n57796 = ~n57751 & n57795;
  assign n57797 = ~n57721 & ~n57796;
  assign n57798 = ~n57740 & ~n57791;
  assign n57799 = ~n57747 & ~n57798;
  assign n57800 = n57727 & n57747;
  assign n57801 = n57733 & n57800;
  assign n57802 = ~n57756 & ~n57801;
  assign n57803 = ~n57799 & n57802;
  assign n57804 = n57721 & n57803;
  assign n57805 = ~n57797 & ~n57804;
  assign n57806 = n57727 & n57758;
  assign n57807 = n57747 & n57806;
  assign n57808 = ~n57805 & ~n57807;
  assign n57809 = n57789 & ~n57808;
  assign n57810 = ~n57794 & ~n57809;
  assign n57811 = ~n57790 & n57810;
  assign n57812 = ~n57763 & n57811;
  assign n57813 = ~n57721 & n57778;
  assign n57814 = n57812 & ~n57813;
  assign n57815 = pi1635 & ~n57814;
  assign n57816 = ~pi1635 & ~n57813;
  assign n57817 = n57811 & n57816;
  assign n57818 = ~n57763 & n57817;
  assign po1715 = n57815 | n57818;
  assign n57820 = pi5304 & ~pi9040;
  assign n57821 = pi5310 & pi9040;
  assign n57822 = ~n57820 & ~n57821;
  assign n57823 = ~pi1622 & ~n57822;
  assign n57824 = pi1622 & n57822;
  assign n57825 = ~n57823 & ~n57824;
  assign n57826 = pi5505 & ~pi9040;
  assign n57827 = pi5325 & pi9040;
  assign n57828 = ~n57826 & ~n57827;
  assign n57829 = pi1628 & n57828;
  assign n57830 = ~pi1628 & ~n57828;
  assign n57831 = ~n57829 & ~n57830;
  assign n57832 = pi5303 & ~pi9040;
  assign n57833 = pi5436 & pi9040;
  assign n57834 = ~n57832 & ~n57833;
  assign n57835 = pi1591 & n57834;
  assign n57836 = ~pi1591 & ~n57834;
  assign n57837 = ~n57835 & ~n57836;
  assign n57838 = pi5437 & pi9040;
  assign n57839 = pi5408 & ~pi9040;
  assign n57840 = ~n57838 & ~n57839;
  assign n57841 = ~pi1620 & ~n57840;
  assign n57842 = pi1620 & n57840;
  assign n57843 = ~n57841 & ~n57842;
  assign n57844 = pi5299 & ~pi9040;
  assign n57845 = pi5566 & pi9040;
  assign n57846 = ~n57844 & ~n57845;
  assign n57847 = pi1607 & n57846;
  assign n57848 = ~pi1607 & ~n57846;
  assign n57849 = ~n57847 & ~n57848;
  assign n57850 = n57843 & ~n57849;
  assign n57851 = ~n57837 & n57850;
  assign n57852 = ~n57831 & n57851;
  assign n57853 = pi5322 & pi9040;
  assign n57854 = pi5502 & ~pi9040;
  assign n57855 = ~n57853 & ~n57854;
  assign n57856 = pi1629 & n57855;
  assign n57857 = ~pi1629 & ~n57855;
  assign n57858 = ~n57856 & ~n57857;
  assign n57859 = ~n57849 & n57858;
  assign n57860 = n57837 & n57859;
  assign n57861 = n57831 & n57860;
  assign n57862 = n57831 & ~n57837;
  assign n57863 = n57843 & n57862;
  assign n57864 = n57858 & n57863;
  assign n57865 = n57849 & n57864;
  assign n57866 = ~n57831 & n57837;
  assign n57867 = n57849 & n57858;
  assign n57868 = n57866 & n57867;
  assign n57869 = n57843 & n57868;
  assign n57870 = ~n57865 & ~n57869;
  assign n57871 = ~n57861 & n57870;
  assign n57872 = ~n57852 & n57871;
  assign n57873 = n57831 & n57837;
  assign n57874 = ~n57849 & n57873;
  assign n57875 = ~n57843 & n57874;
  assign n57876 = n57872 & ~n57875;
  assign n57877 = ~n57825 & ~n57876;
  assign n57878 = ~n57831 & n57850;
  assign n57879 = ~n57831 & ~n57837;
  assign n57880 = ~n57849 & n57879;
  assign n57881 = ~n57878 & ~n57880;
  assign n57882 = ~n57858 & ~n57881;
  assign n57883 = ~n57837 & ~n57843;
  assign n57884 = n57831 & n57883;
  assign n57885 = ~n57858 & n57884;
  assign n57886 = n57849 & n57885;
  assign n57887 = ~n57882 & ~n57886;
  assign n57888 = ~n57825 & ~n57887;
  assign n57889 = n57831 & n57843;
  assign n57890 = n57837 & n57889;
  assign n57891 = n57849 & n57890;
  assign n57892 = ~n57851 & ~n57891;
  assign n57893 = ~n57843 & n57866;
  assign n57894 = n57849 & n57893;
  assign n57895 = n57892 & ~n57894;
  assign n57896 = ~n57858 & ~n57895;
  assign n57897 = ~n57888 & ~n57896;
  assign n57898 = ~n57877 & n57897;
  assign n57899 = ~n57843 & n57849;
  assign n57900 = n57858 & n57899;
  assign n57901 = n57879 & n57900;
  assign n57902 = n57831 & ~n57843;
  assign n57903 = n57859 & n57902;
  assign n57904 = ~n57849 & n57884;
  assign n57905 = n57843 & ~n57858;
  assign n57906 = n57831 & n57905;
  assign n57907 = ~n57831 & n57849;
  assign n57908 = ~n57843 & n57907;
  assign n57909 = ~n57906 & ~n57908;
  assign n57910 = ~n57904 & n57909;
  assign n57911 = ~n57893 & n57910;
  assign n57912 = n57858 & n57866;
  assign n57913 = ~n57849 & n57912;
  assign n57914 = n57849 & n57879;
  assign n57915 = n57837 & ~n57843;
  assign n57916 = ~n57914 & ~n57915;
  assign n57917 = n57858 & ~n57916;
  assign n57918 = ~n57913 & ~n57917;
  assign n57919 = n57911 & n57918;
  assign n57920 = n57825 & ~n57919;
  assign n57921 = ~n57903 & ~n57920;
  assign n57922 = ~n57901 & n57921;
  assign n57923 = n57898 & n57922;
  assign n57924 = pi1634 & n57923;
  assign n57925 = ~pi1634 & ~n57923;
  assign po1720 = n57924 | n57925;
  assign n57927 = pi5570 & ~pi9040;
  assign n57928 = pi5565 & pi9040;
  assign n57929 = ~n57927 & ~n57928;
  assign n57930 = ~pi1600 & ~n57929;
  assign n57931 = pi1600 & n57929;
  assign n57932 = ~n57930 & ~n57931;
  assign n57933 = pi5442 & ~pi9040;
  assign n57934 = pi5401 & pi9040;
  assign n57935 = ~n57933 & ~n57934;
  assign n57936 = ~pi1611 & n57935;
  assign n57937 = pi1611 & ~n57935;
  assign n57938 = ~n57936 & ~n57937;
  assign n57939 = pi5309 & pi9040;
  assign n57940 = pi5415 & ~pi9040;
  assign n57941 = ~n57939 & ~n57940;
  assign n57942 = pi1608 & n57941;
  assign n57943 = ~pi1608 & ~n57941;
  assign n57944 = ~n57942 & ~n57943;
  assign n57945 = n57938 & n57944;
  assign n57946 = pi5434 & ~pi9040;
  assign n57947 = pi5317 & pi9040;
  assign n57948 = ~n57946 & ~n57947;
  assign n57949 = ~pi1599 & ~n57948;
  assign n57950 = pi1599 & n57948;
  assign n57951 = ~n57949 & ~n57950;
  assign n57952 = pi5308 & pi9040;
  assign n57953 = pi5323 & ~pi9040;
  assign n57954 = ~n57952 & ~n57953;
  assign n57955 = pi1625 & n57954;
  assign n57956 = ~pi1625 & ~n57954;
  assign n57957 = ~n57955 & ~n57956;
  assign n57958 = ~n57951 & ~n57957;
  assign n57959 = n57945 & n57958;
  assign n57960 = pi5320 & pi9040;
  assign n57961 = pi5509 & ~pi9040;
  assign n57962 = ~n57960 & ~n57961;
  assign n57963 = ~pi1593 & n57962;
  assign n57964 = pi1593 & ~n57962;
  assign n57965 = ~n57963 & ~n57964;
  assign n57966 = ~n57938 & ~n57944;
  assign n57967 = ~n57965 & n57966;
  assign n57968 = n57951 & n57965;
  assign n57969 = ~n57944 & n57968;
  assign n57970 = n57938 & n57969;
  assign n57971 = ~n57967 & ~n57970;
  assign n57972 = ~n57938 & n57944;
  assign n57973 = n57951 & n57972;
  assign n57974 = n57971 & ~n57973;
  assign n57975 = ~n57957 & ~n57974;
  assign n57976 = ~n57938 & n57965;
  assign n57977 = ~n57951 & n57957;
  assign n57978 = n57976 & n57977;
  assign n57979 = n57965 & n57966;
  assign n57980 = ~n57951 & n57979;
  assign n57981 = ~n57978 & ~n57980;
  assign n57982 = ~n57975 & n57981;
  assign n57983 = ~n57959 & n57982;
  assign n57984 = ~n57965 & n57972;
  assign n57985 = n57951 & n57984;
  assign n57986 = n57945 & ~n57965;
  assign n57987 = ~n57951 & n57986;
  assign n57988 = ~n57985 & ~n57987;
  assign n57989 = n57983 & n57988;
  assign n57990 = ~n57932 & ~n57989;
  assign n57991 = ~n57951 & n57965;
  assign n57992 = n57944 & n57991;
  assign n57993 = ~n57938 & n57992;
  assign n57994 = ~n57986 & ~n57993;
  assign n57995 = ~n57957 & ~n57994;
  assign n57996 = ~n57938 & n57968;
  assign n57997 = ~n57951 & n57984;
  assign n57998 = ~n57996 & ~n57997;
  assign n57999 = n57957 & ~n57998;
  assign n58000 = n57945 & n57968;
  assign n58001 = ~n57944 & n57991;
  assign n58002 = n57938 & n58001;
  assign n58003 = ~n58000 & ~n58002;
  assign n58004 = ~n57999 & n58003;
  assign n58005 = ~n57995 & n58004;
  assign n58006 = n57932 & ~n58005;
  assign n58007 = ~n57938 & ~n57965;
  assign n58008 = n57951 & n58007;
  assign n58009 = n57938 & ~n57965;
  assign n58010 = ~n57951 & n58009;
  assign n58011 = ~n58008 & ~n58010;
  assign n58012 = ~n57957 & ~n58011;
  assign n58013 = n57938 & ~n57944;
  assign n58014 = ~n57965 & n58013;
  assign n58015 = n57951 & n58014;
  assign n58016 = ~n58000 & ~n58015;
  assign n58017 = ~n57979 & n58016;
  assign n58018 = n57957 & ~n58017;
  assign n58019 = ~n58012 & ~n58018;
  assign n58020 = ~n57944 & n57965;
  assign n58021 = n57957 & n58020;
  assign n58022 = ~n57951 & n58021;
  assign n58023 = n58019 & ~n58022;
  assign n58024 = ~n58006 & n58023;
  assign n58025 = ~n57990 & n58024;
  assign n58026 = ~pi1639 & ~n58025;
  assign n58027 = pi1639 & n58025;
  assign po1721 = n58026 | n58027;
  assign n58029 = ~n57831 & n57843;
  assign n58030 = ~n57875 & ~n58029;
  assign n58031 = ~n57907 & n58030;
  assign n58032 = n57858 & ~n58031;
  assign n58033 = n57849 & ~n57858;
  assign n58034 = n57831 & n58033;
  assign n58035 = n57843 & n57849;
  assign n58036 = n57837 & n58035;
  assign n58037 = ~n57849 & n57863;
  assign n58038 = ~n58036 & ~n58037;
  assign n58039 = ~n57831 & ~n57843;
  assign n58040 = ~n57849 & ~n57858;
  assign n58041 = n58039 & n58040;
  assign n58042 = n58038 & ~n58041;
  assign n58043 = ~n58034 & n58042;
  assign n58044 = ~n58032 & n58043;
  assign n58045 = n57825 & ~n58044;
  assign n58046 = n57843 & n57866;
  assign n58047 = ~n57849 & n58046;
  assign n58048 = n57843 & n57879;
  assign n58049 = n57849 & n58048;
  assign n58050 = ~n58047 & ~n58049;
  assign n58051 = n57858 & ~n58050;
  assign n58052 = ~n58045 & ~n58051;
  assign n58053 = n57849 & n57863;
  assign n58054 = ~n57884 & ~n57890;
  assign n58055 = n57858 & ~n58054;
  assign n58056 = ~n58053 & ~n58055;
  assign n58057 = ~n57894 & n58056;
  assign n58058 = ~n57825 & ~n58057;
  assign n58059 = ~n57873 & ~n57879;
  assign n58060 = ~n57843 & ~n58059;
  assign n58061 = ~n57880 & ~n58060;
  assign n58062 = ~n57858 & ~n58061;
  assign n58063 = ~n57825 & n58062;
  assign n58064 = ~n58058 & ~n58063;
  assign n58065 = n58052 & n58064;
  assign n58066 = pi1640 & ~n58065;
  assign n58067 = ~pi1640 & n58052;
  assign n58068 = n58064 & n58067;
  assign po1722 = n58066 | n58068;
  assign n58070 = ~n57579 & n57617;
  assign n58071 = ~n57655 & ~n58070;
  assign n58072 = ~n57660 & n58071;
  assign n58073 = n57586 & n57608;
  assign n58074 = ~n57619 & ~n57652;
  assign n58075 = ~n57579 & ~n58074;
  assign n58076 = ~n58073 & ~n58075;
  assign n58077 = n57586 & ~n57598;
  assign n58078 = ~n57615 & ~n58077;
  assign n58079 = ~n57662 & n58078;
  assign n58080 = n57579 & ~n58079;
  assign n58081 = n58076 & ~n58080;
  assign n58082 = ~n57573 & ~n58081;
  assign n58083 = ~n57586 & n57592;
  assign n58084 = ~n57606 & n58083;
  assign n58085 = ~n57659 & ~n58084;
  assign n58086 = n57579 & n57634;
  assign n58087 = n57586 & n57619;
  assign n58088 = ~n57579 & n57615;
  assign n58089 = ~n58087 & ~n58088;
  assign n58090 = ~n57703 & n58089;
  assign n58091 = ~n58086 & n58090;
  assign n58092 = n58085 & n58091;
  assign n58093 = ~n57645 & n58092;
  assign n58094 = n57573 & ~n58093;
  assign n58095 = ~n58082 & ~n58094;
  assign n58096 = n58072 & n58095;
  assign n58097 = ~pi1660 & ~n58096;
  assign n58098 = pi1660 & n58072;
  assign n58099 = ~n58082 & n58098;
  assign n58100 = ~n58094 & n58099;
  assign po1724 = n58097 | n58100;
  assign n58102 = pi5316 & ~pi9040;
  assign n58103 = pi5443 & pi9040;
  assign n58104 = ~n58102 & ~n58103;
  assign n58105 = ~pi1612 & ~n58104;
  assign n58106 = pi1612 & n58104;
  assign n58107 = ~n58105 & ~n58106;
  assign n58108 = pi5392 & pi9040;
  assign n58109 = pi5513 & ~pi9040;
  assign n58110 = ~n58108 & ~n58109;
  assign n58111 = pi1630 & n58110;
  assign n58112 = ~pi1630 & ~n58110;
  assign n58113 = ~n58111 & ~n58112;
  assign n58114 = pi5511 & pi9040;
  assign n58115 = pi5514 & ~pi9040;
  assign n58116 = ~n58114 & ~n58115;
  assign n58117 = ~pi1627 & ~n58116;
  assign n58118 = pi1627 & n58116;
  assign n58119 = ~n58117 & ~n58118;
  assign n58120 = pi5396 & ~pi9040;
  assign n58121 = pi5415 & pi9040;
  assign n58122 = ~n58120 & ~n58121;
  assign n58123 = ~pi1605 & ~n58122;
  assign n58124 = pi1605 & n58122;
  assign n58125 = ~n58123 & ~n58124;
  assign n58126 = pi5323 & pi9040;
  assign n58127 = pi5318 & ~pi9040;
  assign n58128 = ~n58126 & ~n58127;
  assign n58129 = ~pi1621 & ~n58128;
  assign n58130 = pi1621 & n58128;
  assign n58131 = ~n58129 & ~n58130;
  assign n58132 = n58125 & ~n58131;
  assign n58133 = n58119 & n58132;
  assign n58134 = n58113 & n58133;
  assign n58135 = pi5311 & pi9040;
  assign n58136 = pi5441 & ~pi9040;
  assign n58137 = ~n58135 & ~n58136;
  assign n58138 = ~pi1623 & n58137;
  assign n58139 = pi1623 & ~n58137;
  assign n58140 = ~n58138 & ~n58139;
  assign n58141 = n58119 & n58131;
  assign n58142 = n58125 & n58141;
  assign n58143 = ~n58119 & ~n58125;
  assign n58144 = ~n58125 & ~n58131;
  assign n58145 = ~n58113 & n58144;
  assign n58146 = ~n58119 & ~n58131;
  assign n58147 = n58113 & n58146;
  assign n58148 = ~n58145 & ~n58147;
  assign n58149 = ~n58143 & n58148;
  assign n58150 = ~n58142 & n58149;
  assign n58151 = ~n58140 & ~n58150;
  assign n58152 = ~n58113 & n58125;
  assign n58153 = n58131 & n58152;
  assign n58154 = ~n58119 & n58152;
  assign n58155 = ~n58125 & n58141;
  assign n58156 = ~n58154 & ~n58155;
  assign n58157 = n58140 & ~n58156;
  assign n58158 = ~n58153 & ~n58157;
  assign n58159 = ~n58151 & n58158;
  assign n58160 = ~n58134 & n58159;
  assign n58161 = n58107 & ~n58160;
  assign n58162 = ~n58119 & n58131;
  assign n58163 = ~n58125 & n58162;
  assign n58164 = ~n58113 & n58163;
  assign n58165 = ~n58125 & n58146;
  assign n58166 = n58113 & n58165;
  assign n58167 = ~n58134 & ~n58166;
  assign n58168 = ~n58164 & n58167;
  assign n58169 = ~n58140 & ~n58168;
  assign n58170 = ~n58161 & ~n58169;
  assign n58171 = n58119 & n58153;
  assign n58172 = n58119 & ~n58125;
  assign n58173 = n58140 & n58172;
  assign n58174 = n58113 & n58173;
  assign n58175 = n58125 & n58162;
  assign n58176 = n58113 & n58175;
  assign n58177 = n58132 & ~n58140;
  assign n58178 = ~n58113 & n58177;
  assign n58179 = ~n58176 & ~n58178;
  assign n58180 = ~n58119 & n58125;
  assign n58181 = n58113 & n58180;
  assign n58182 = n58119 & ~n58131;
  assign n58183 = ~n58125 & n58182;
  assign n58184 = ~n58181 & ~n58183;
  assign n58185 = n58140 & ~n58184;
  assign n58186 = n58140 & n58143;
  assign n58187 = ~n58113 & n58186;
  assign n58188 = ~n58185 & ~n58187;
  assign n58189 = n58179 & n58188;
  assign n58190 = ~n58107 & ~n58189;
  assign n58191 = ~n58174 & ~n58190;
  assign n58192 = ~n58171 & n58191;
  assign n58193 = n58170 & n58192;
  assign n58194 = ~pi1637 & ~n58193;
  assign n58195 = ~n58161 & ~n58171;
  assign n58196 = ~n58169 & n58195;
  assign n58197 = n58191 & n58196;
  assign n58198 = pi1637 & n58197;
  assign po1725 = n58194 | n58198;
  assign n58200 = ~n57849 & n57893;
  assign n58201 = ~n58037 & ~n58200;
  assign n58202 = ~n57858 & ~n58201;
  assign n58203 = n57890 & n58033;
  assign n58204 = ~n58202 & ~n58203;
  assign n58205 = ~n57903 & n58204;
  assign n58206 = n57843 & n57858;
  assign n58207 = ~n57837 & n58206;
  assign n58208 = ~n57831 & n58207;
  assign n58209 = ~n57849 & n58208;
  assign n58210 = n57858 & n58046;
  assign n58211 = ~n57875 & ~n57901;
  assign n58212 = ~n57865 & n58211;
  assign n58213 = ~n58210 & n58212;
  assign n58214 = n57825 & ~n58213;
  assign n58215 = n57849 & n57884;
  assign n58216 = ~n57893 & ~n58215;
  assign n58217 = ~n58048 & n58216;
  assign n58218 = ~n57858 & ~n58217;
  assign n58219 = n57825 & n58218;
  assign n58220 = n57849 & n57912;
  assign n58221 = ~n58208 & ~n58220;
  assign n58222 = ~n58036 & n58221;
  assign n58223 = ~n57843 & ~n57849;
  assign n58224 = ~n57837 & n58223;
  assign n58225 = n57849 & n57873;
  assign n58226 = ~n57889 & ~n58225;
  assign n58227 = ~n57858 & ~n58226;
  assign n58228 = ~n58224 & ~n58227;
  assign n58229 = n58222 & n58228;
  assign n58230 = ~n57825 & ~n58229;
  assign n58231 = ~n58219 & ~n58230;
  assign n58232 = ~n58214 & n58231;
  assign n58233 = ~n58209 & n58232;
  assign n58234 = n58205 & n58233;
  assign n58235 = pi1644 & ~n58234;
  assign n58236 = ~pi1644 & n58205;
  assign n58237 = n58233 & n58236;
  assign po1727 = n58235 | n58237;
  assign n58239 = pi5399 & ~pi9040;
  assign n58240 = pi5505 & pi9040;
  assign n58241 = ~n58239 & ~n58240;
  assign n58242 = ~pi1627 & ~n58241;
  assign n58243 = pi1627 & n58241;
  assign n58244 = ~n58242 & ~n58243;
  assign n58245 = pi5306 & pi9040;
  assign n58246 = pi5328 & ~pi9040;
  assign n58247 = ~n58245 & ~n58246;
  assign n58248 = ~pi1615 & n58247;
  assign n58249 = pi1615 & ~n58247;
  assign n58250 = ~n58248 & ~n58249;
  assign n58251 = pi5576 & pi9040;
  assign n58252 = pi5398 & ~pi9040;
  assign n58253 = ~n58251 & ~n58252;
  assign n58254 = ~pi1609 & n58253;
  assign n58255 = pi1609 & ~n58253;
  assign n58256 = ~n58254 & ~n58255;
  assign n58257 = pi5408 & pi9040;
  assign n58258 = pi5665 & ~pi9040;
  assign n58259 = ~n58257 & ~n58258;
  assign n58260 = ~pi1614 & n58259;
  assign n58261 = pi1614 & ~n58259;
  assign n58262 = ~n58260 & ~n58261;
  assign n58263 = pi5310 & ~pi9040;
  assign n58264 = pi5403 & pi9040;
  assign n58265 = ~n58263 & ~n58264;
  assign n58266 = ~pi1605 & n58265;
  assign n58267 = pi1605 & ~n58265;
  assign n58268 = ~n58266 & ~n58267;
  assign n58269 = ~n58262 & n58268;
  assign n58270 = ~n58256 & n58269;
  assign n58271 = ~n58250 & n58270;
  assign n58272 = ~pi1614 & ~n58259;
  assign n58273 = pi1614 & n58259;
  assign n58274 = ~n58272 & ~n58273;
  assign n58275 = n58268 & ~n58274;
  assign n58276 = ~n58256 & n58275;
  assign n58277 = n58250 & n58276;
  assign n58278 = ~n58271 & ~n58277;
  assign n58279 = ~n58268 & ~n58274;
  assign n58280 = ~n58256 & n58279;
  assign n58281 = ~n58250 & n58280;
  assign n58282 = pi5305 & pi9040;
  assign n58283 = pi5313 & ~pi9040;
  assign n58284 = ~n58282 & ~n58283;
  assign n58285 = ~pi1631 & ~n58284;
  assign n58286 = pi1631 & n58284;
  assign n58287 = ~n58285 & ~n58286;
  assign n58288 = ~n58262 & ~n58268;
  assign n58289 = ~n58250 & n58288;
  assign n58290 = n58256 & n58279;
  assign n58291 = n58250 & n58290;
  assign n58292 = ~n58289 & ~n58291;
  assign n58293 = ~n58287 & ~n58292;
  assign n58294 = ~n58281 & ~n58293;
  assign n58295 = n58256 & n58275;
  assign n58296 = n58287 & n58295;
  assign n58297 = n58279 & n58287;
  assign n58298 = ~n58250 & n58297;
  assign n58299 = ~n58296 & ~n58298;
  assign n58300 = n58294 & n58299;
  assign n58301 = n58278 & n58300;
  assign n58302 = n58244 & ~n58301;
  assign n58303 = ~n58244 & ~n58287;
  assign n58304 = ~n58250 & n58256;
  assign n58305 = n58262 & n58304;
  assign n58306 = n58256 & n58268;
  assign n58307 = ~n58305 & ~n58306;
  assign n58308 = n58303 & ~n58307;
  assign n58309 = n58250 & ~n58256;
  assign n58310 = ~n58268 & n58309;
  assign n58311 = ~n58274 & n58310;
  assign n58312 = n58250 & ~n58262;
  assign n58313 = n58256 & n58312;
  assign n58314 = ~n58311 & ~n58313;
  assign n58315 = ~n58250 & n58287;
  assign n58316 = ~n58256 & n58315;
  assign n58317 = ~n58279 & n58316;
  assign n58318 = n58270 & n58287;
  assign n58319 = ~n58317 & ~n58318;
  assign n58320 = n58314 & n58319;
  assign n58321 = ~n58244 & ~n58320;
  assign n58322 = n58256 & n58269;
  assign n58323 = ~n58287 & n58322;
  assign n58324 = n58250 & n58323;
  assign n58325 = ~n58256 & n58288;
  assign n58326 = n58250 & n58325;
  assign n58327 = ~n58277 & ~n58326;
  assign n58328 = ~n58287 & ~n58327;
  assign n58329 = ~n58324 & ~n58328;
  assign n58330 = n58287 & n58311;
  assign n58331 = n58329 & ~n58330;
  assign n58332 = ~n58321 & n58331;
  assign n58333 = ~n58308 & n58332;
  assign n58334 = ~n58302 & n58333;
  assign n58335 = n58256 & n58288;
  assign n58336 = n58250 & n58287;
  assign n58337 = n58335 & n58336;
  assign n58338 = n58334 & ~n58337;
  assign n58339 = ~pi1642 & ~n58338;
  assign n58340 = pi1642 & ~n58337;
  assign n58341 = n58333 & n58340;
  assign n58342 = ~n58302 & n58341;
  assign po1728 = n58339 | n58342;
  assign n58344 = n58125 & n58146;
  assign n58345 = n58113 & n58344;
  assign n58346 = n58113 & n58163;
  assign n58347 = ~n58345 & ~n58346;
  assign n58348 = ~n58113 & ~n58125;
  assign n58349 = ~n58131 & n58348;
  assign n58350 = ~n58119 & n58349;
  assign n58351 = ~n58155 & ~n58350;
  assign n58352 = ~n58140 & ~n58351;
  assign n58353 = n58347 & ~n58352;
  assign n58354 = ~n58113 & n58140;
  assign n58355 = n58119 & n58354;
  assign n58356 = n58353 & ~n58355;
  assign n58357 = n58107 & ~n58356;
  assign n58358 = n58113 & n58183;
  assign n58359 = n58140 & n58358;
  assign n58360 = ~n58113 & ~n58140;
  assign n58361 = n58183 & n58360;
  assign n58362 = ~n58154 & ~n58361;
  assign n58363 = ~n58155 & ~n58175;
  assign n58364 = ~n58113 & n58162;
  assign n58365 = n58363 & ~n58364;
  assign n58366 = n58140 & ~n58365;
  assign n58367 = ~n58140 & n58142;
  assign n58368 = n58167 & ~n58367;
  assign n58369 = ~n58366 & n58368;
  assign n58370 = n58362 & n58369;
  assign n58371 = ~n58107 & ~n58370;
  assign n58372 = ~n58359 & ~n58371;
  assign n58373 = ~n58357 & n58372;
  assign n58374 = n58175 & n58360;
  assign n58375 = n58113 & n58177;
  assign n58376 = ~n58374 & ~n58375;
  assign n58377 = ~n58140 & n58346;
  assign n58378 = n58376 & ~n58377;
  assign n58379 = n58373 & n58378;
  assign n58380 = ~pi1632 & ~n58379;
  assign n58381 = n58372 & n58378;
  assign n58382 = pi1632 & n58381;
  assign n58383 = ~n58357 & n58382;
  assign po1730 = n58380 | n58383;
  assign n58385 = n57849 & n58060;
  assign n58386 = ~n57883 & ~n58046;
  assign n58387 = ~n57858 & ~n58386;
  assign n58388 = ~n58385 & ~n58387;
  assign n58389 = ~n57837 & n58035;
  assign n58390 = ~n57915 & ~n58389;
  assign n58391 = ~n58048 & n58390;
  assign n58392 = n57858 & ~n58391;
  assign n58393 = n58388 & ~n58392;
  assign n58394 = ~n57849 & n57890;
  assign n58395 = n58393 & ~n58394;
  assign n58396 = ~n57825 & ~n58395;
  assign n58397 = n57859 & ~n58386;
  assign n58398 = ~n57884 & ~n57893;
  assign n58399 = ~n57890 & ~n58048;
  assign n58400 = n58398 & n58399;
  assign n58401 = n57849 & ~n58400;
  assign n58402 = ~n58397 & ~n58401;
  assign n58403 = ~n58037 & n58402;
  assign n58404 = n57825 & ~n58403;
  assign n58405 = ~n58396 & ~n58404;
  assign n58406 = n57849 & n58046;
  assign n58407 = ~n58394 & ~n58406;
  assign n58408 = ~n57858 & ~n58407;
  assign n58409 = n58405 & ~n58408;
  assign n58410 = pi1633 & ~n58409;
  assign n58411 = ~pi1633 & ~n58408;
  assign n58412 = ~n58404 & n58411;
  assign n58413 = ~n58396 & n58412;
  assign po1731 = n58410 | n58413;
  assign n58415 = n58250 & n58295;
  assign n58416 = ~n58250 & n58322;
  assign n58417 = ~n58415 & ~n58416;
  assign n58418 = n58287 & ~n58417;
  assign n58419 = ~n58287 & n58311;
  assign n58420 = ~n58311 & ~n58318;
  assign n58421 = ~n58250 & ~n58256;
  assign n58422 = ~n58268 & n58421;
  assign n58423 = ~n58262 & n58422;
  assign n58424 = ~n58250 & ~n58287;
  assign n58425 = n58275 & n58424;
  assign n58426 = n58256 & n58425;
  assign n58427 = ~n58274 & n58309;
  assign n58428 = ~n58313 & ~n58427;
  assign n58429 = ~n58287 & ~n58428;
  assign n58430 = n58256 & n58287;
  assign n58431 = ~n58268 & n58430;
  assign n58432 = ~n58274 & n58431;
  assign n58433 = ~n58429 & ~n58432;
  assign n58434 = ~n58426 & n58433;
  assign n58435 = ~n58423 & n58434;
  assign n58436 = n58420 & n58435;
  assign n58437 = n58244 & ~n58436;
  assign n58438 = n58250 & n58318;
  assign n58439 = ~n58437 & ~n58438;
  assign n58440 = ~n58419 & n58439;
  assign n58441 = ~n58418 & n58440;
  assign n58442 = ~n58256 & ~n58274;
  assign n58443 = n58315 & n58442;
  assign n58444 = ~n58296 & ~n58443;
  assign n58445 = n58287 & n58325;
  assign n58446 = n58250 & n58335;
  assign n58447 = ~n58445 & ~n58446;
  assign n58448 = ~n58250 & n58276;
  assign n58449 = ~n58415 & ~n58448;
  assign n58450 = ~n58250 & n58269;
  assign n58451 = n58256 & ~n58268;
  assign n58452 = ~n58450 & ~n58451;
  assign n58453 = ~n58287 & ~n58452;
  assign n58454 = n58449 & ~n58453;
  assign n58455 = n58447 & n58454;
  assign n58456 = n58444 & n58455;
  assign n58457 = ~n58244 & ~n58456;
  assign n58458 = n58441 & ~n58457;
  assign n58459 = ~pi1645 & ~n58458;
  assign n58460 = pi1645 & n58441;
  assign n58461 = ~n58457 & n58460;
  assign po1732 = n58459 | n58461;
  assign n58463 = pi5305 & ~pi9040;
  assign n58464 = pi5405 & pi9040;
  assign n58465 = ~n58463 & ~n58464;
  assign n58466 = ~pi1610 & ~n58465;
  assign n58467 = pi1610 & n58465;
  assign n58468 = ~n58466 & ~n58467;
  assign n58469 = pi5325 & ~pi9040;
  assign n58470 = pi5665 & pi9040;
  assign n58471 = ~n58469 & ~n58470;
  assign n58472 = pi1616 & n58471;
  assign n58473 = ~pi1616 & ~n58471;
  assign n58474 = ~n58472 & ~n58473;
  assign n58475 = pi5398 & pi9040;
  assign n58476 = pi5436 & ~pi9040;
  assign n58477 = ~n58475 & ~n58476;
  assign n58478 = pi1626 & n58477;
  assign n58479 = ~pi1626 & ~n58477;
  assign n58480 = ~n58478 & ~n58479;
  assign n58481 = n58474 & ~n58480;
  assign n58482 = pi5403 & ~pi9040;
  assign n58483 = pi5321 & pi9040;
  assign n58484 = ~n58482 & ~n58483;
  assign n58485 = pi1622 & n58484;
  assign n58486 = ~pi1622 & ~n58484;
  assign n58487 = ~n58485 & ~n58486;
  assign n58488 = pi5573 & ~pi9040;
  assign n58489 = pi5299 & pi9040;
  assign n58490 = ~n58488 & ~n58489;
  assign n58491 = ~pi1618 & n58490;
  assign n58492 = pi1618 & ~n58490;
  assign n58493 = ~n58491 & ~n58492;
  assign n58494 = ~n58487 & n58493;
  assign n58495 = pi5304 & pi9040;
  assign n58496 = pi5306 & ~pi9040;
  assign n58497 = ~n58495 & ~n58496;
  assign n58498 = ~pi1591 & n58497;
  assign n58499 = pi1591 & ~n58497;
  assign n58500 = ~n58498 & ~n58499;
  assign n58501 = n58487 & ~n58493;
  assign n58502 = n58500 & n58501;
  assign n58503 = ~n58494 & ~n58502;
  assign n58504 = n58481 & ~n58503;
  assign n58505 = ~n58480 & n58500;
  assign n58506 = n58494 & n58505;
  assign n58507 = ~n58504 & ~n58506;
  assign n58508 = n58468 & ~n58507;
  assign n58509 = ~n58474 & ~n58500;
  assign n58510 = ~n58493 & n58509;
  assign n58511 = n58487 & n58510;
  assign n58512 = n58487 & ~n58500;
  assign n58513 = ~n58509 & ~n58512;
  assign n58514 = n58480 & ~n58513;
  assign n58515 = ~n58474 & n58500;
  assign n58516 = n58493 & n58515;
  assign n58517 = n58487 & n58516;
  assign n58518 = ~n58514 & ~n58517;
  assign n58519 = ~n58511 & n58518;
  assign n58520 = n58468 & ~n58519;
  assign n58521 = ~n58508 & ~n58520;
  assign n58522 = n58474 & ~n58500;
  assign n58523 = ~n58493 & n58522;
  assign n58524 = ~n58487 & n58523;
  assign n58525 = ~n58487 & ~n58493;
  assign n58526 = n58500 & n58525;
  assign n58527 = ~n58474 & n58526;
  assign n58528 = ~n58524 & ~n58527;
  assign n58529 = ~n58480 & ~n58528;
  assign n58530 = n58494 & n58500;
  assign n58531 = n58474 & n58530;
  assign n58532 = ~n58474 & n58512;
  assign n58533 = ~n58531 & ~n58532;
  assign n58534 = n58480 & ~n58533;
  assign n58535 = n58487 & n58493;
  assign n58536 = ~n58512 & ~n58535;
  assign n58537 = n58474 & ~n58536;
  assign n58538 = ~n58526 & ~n58537;
  assign n58539 = ~n58480 & ~n58538;
  assign n58540 = ~n58474 & ~n58493;
  assign n58541 = n58505 & n58540;
  assign n58542 = n58493 & ~n58500;
  assign n58543 = ~n58526 & ~n58542;
  assign n58544 = ~n58474 & ~n58543;
  assign n58545 = n58474 & n58480;
  assign n58546 = n58501 & n58545;
  assign n58547 = n58500 & n58546;
  assign n58548 = ~n58544 & ~n58547;
  assign n58549 = ~n58541 & n58548;
  assign n58550 = ~n58539 & n58549;
  assign n58551 = ~n58524 & n58550;
  assign n58552 = ~n58468 & ~n58551;
  assign n58553 = ~n58534 & ~n58552;
  assign n58554 = ~n58529 & n58553;
  assign n58555 = n58521 & n58554;
  assign n58556 = pi1641 & n58555;
  assign n58557 = ~pi1641 & ~n58555;
  assign po1733 = n58556 | n58557;
  assign n58559 = n57579 & n57607;
  assign n58560 = ~n57586 & n58559;
  assign n58561 = ~n57663 & ~n58560;
  assign n58562 = n57586 & n57592;
  assign n58563 = n57606 & n58562;
  assign n58564 = ~n57586 & n57598;
  assign n58565 = ~n58084 & ~n58564;
  assign n58566 = ~n57579 & ~n58565;
  assign n58567 = ~n58563 & ~n58566;
  assign n58568 = n58561 & n58567;
  assign n58569 = n57573 & ~n58568;
  assign n58570 = ~n57638 & ~n57640;
  assign n58571 = ~n57586 & n57618;
  assign n58572 = n58570 & ~n58571;
  assign n58573 = n57579 & ~n58572;
  assign n58574 = n57607 & n57631;
  assign n58575 = ~n57612 & ~n58574;
  assign n58576 = ~n58573 & n58575;
  assign n58577 = ~n57662 & ~n57686;
  assign n58578 = ~n57579 & ~n58577;
  assign n58579 = n58576 & ~n58578;
  assign n58580 = ~n57573 & ~n58579;
  assign n58581 = ~n58569 & ~n58580;
  assign n58582 = ~n57586 & n57651;
  assign n58583 = n57586 & ~n57683;
  assign n58584 = ~n58582 & ~n58583;
  assign n58585 = ~n57579 & ~n58584;
  assign n58586 = ~n57638 & n58074;
  assign n58587 = n57642 & ~n58586;
  assign n58588 = ~n58585 & ~n58587;
  assign n58589 = n58581 & n58588;
  assign n58590 = ~pi1658 & ~n58589;
  assign n58591 = pi1658 & n58588;
  assign n58592 = ~n58580 & n58591;
  assign n58593 = ~n58569 & n58592;
  assign po1734 = n58590 | n58593;
  assign n58595 = n57951 & n57979;
  assign n58596 = ~n58002 & ~n58007;
  assign n58597 = n57957 & ~n58596;
  assign n58598 = ~n58595 & ~n58597;
  assign n58599 = ~n57993 & n58598;
  assign n58600 = ~n57957 & n58000;
  assign n58601 = ~n57987 & ~n58600;
  assign n58602 = ~n58015 & n58601;
  assign n58603 = n58599 & n58602;
  assign n58604 = n57932 & ~n58603;
  assign n58605 = ~n57951 & n58014;
  assign n58606 = n57944 & ~n57965;
  assign n58607 = ~n57938 & n57951;
  assign n58608 = ~n58606 & ~n58607;
  assign n58609 = ~n58020 & n58608;
  assign n58610 = ~n57957 & ~n58609;
  assign n58611 = ~n58605 & ~n58610;
  assign n58612 = n57951 & n57986;
  assign n58613 = n57965 & n57972;
  assign n58614 = n57951 & n58613;
  assign n58615 = ~n57970 & ~n58614;
  assign n58616 = n57945 & n57965;
  assign n58617 = n57957 & n58616;
  assign n58618 = n58615 & ~n58617;
  assign n58619 = ~n58612 & n58618;
  assign n58620 = ~n57980 & n58619;
  assign n58621 = n58611 & n58620;
  assign n58622 = ~n57932 & ~n58621;
  assign n58623 = ~n58604 & ~n58622;
  assign n58624 = pi1643 & ~n58623;
  assign n58625 = ~pi1643 & ~n58604;
  assign n58626 = ~n58622 & n58625;
  assign po1735 = n58624 | n58626;
  assign n58628 = ~n58113 & n58344;
  assign n58629 = ~n58163 & ~n58171;
  assign n58630 = n58113 & n58132;
  assign n58631 = ~n58113 & n58183;
  assign n58632 = ~n58630 & ~n58631;
  assign n58633 = n58629 & n58632;
  assign n58634 = n58140 & ~n58633;
  assign n58635 = n58113 & n58141;
  assign n58636 = ~n58154 & ~n58635;
  assign n58637 = ~n58165 & n58636;
  assign n58638 = ~n58140 & ~n58637;
  assign n58639 = n58113 & ~n58125;
  assign n58640 = n58131 & n58639;
  assign n58641 = n58119 & n58640;
  assign n58642 = ~n58638 & ~n58641;
  assign n58643 = ~n58634 & n58642;
  assign n58644 = ~n58628 & n58643;
  assign n58645 = ~n58107 & ~n58644;
  assign n58646 = n58113 & n58140;
  assign n58647 = n58142 & n58646;
  assign n58648 = n58140 & n58165;
  assign n58649 = n58140 & n58175;
  assign n58650 = ~n58648 & ~n58649;
  assign n58651 = ~n58113 & ~n58650;
  assign n58652 = ~n58647 & ~n58651;
  assign n58653 = ~n58113 & n58133;
  assign n58654 = ~n58358 & ~n58653;
  assign n58655 = n58113 & n58162;
  assign n58656 = ~n58113 & n58141;
  assign n58657 = ~n58655 & ~n58656;
  assign n58658 = ~n58133 & n58657;
  assign n58659 = ~n58163 & n58658;
  assign n58660 = ~n58140 & ~n58659;
  assign n58661 = ~n58113 & n58155;
  assign n58662 = ~n58660 & ~n58661;
  assign n58663 = n58654 & n58662;
  assign n58664 = n58652 & n58663;
  assign n58665 = n58107 & ~n58664;
  assign n58666 = n58140 & ~n58347;
  assign n58667 = ~n58665 & ~n58666;
  assign n58668 = ~n58166 & ~n58653;
  assign n58669 = ~n58140 & ~n58668;
  assign n58670 = n58667 & ~n58669;
  assign n58671 = ~n58645 & n58670;
  assign n58672 = pi1636 & ~n58671;
  assign n58673 = ~pi1636 & n58671;
  assign po1736 = n58672 | n58673;
  assign n58675 = n58522 & n58535;
  assign n58676 = n58474 & n58500;
  assign n58677 = ~n58487 & n58676;
  assign n58678 = ~n58675 & ~n58677;
  assign n58679 = ~n58480 & ~n58678;
  assign n58680 = ~n58474 & n58480;
  assign n58681 = n58487 & n58680;
  assign n58682 = n58500 & n58535;
  assign n58683 = ~n58500 & n58501;
  assign n58684 = ~n58682 & ~n58683;
  assign n58685 = n58494 & ~n58500;
  assign n58686 = n58474 & n58685;
  assign n58687 = n58684 & ~n58686;
  assign n58688 = n58480 & ~n58687;
  assign n58689 = ~n58681 & ~n58688;
  assign n58690 = n58474 & n58526;
  assign n58691 = n58689 & ~n58690;
  assign n58692 = ~n58474 & n58494;
  assign n58693 = ~n58500 & n58525;
  assign n58694 = ~n58692 & ~n58693;
  assign n58695 = ~n58480 & ~n58694;
  assign n58696 = ~n58474 & n58502;
  assign n58697 = ~n58695 & ~n58696;
  assign n58698 = n58691 & n58697;
  assign n58699 = n58468 & ~n58698;
  assign n58700 = ~n58679 & ~n58699;
  assign n58701 = ~n58468 & n58480;
  assign n58702 = ~n58694 & n58701;
  assign n58703 = ~n58502 & ~n58530;
  assign n58704 = n58474 & ~n58703;
  assign n58705 = ~n58675 & ~n58704;
  assign n58706 = ~n58468 & ~n58705;
  assign n58707 = ~n58702 & ~n58706;
  assign n58708 = ~n58468 & ~n58480;
  assign n58709 = ~n58474 & n58535;
  assign n58710 = ~n58526 & ~n58709;
  assign n58711 = ~n58512 & n58710;
  assign n58712 = n58708 & ~n58711;
  assign n58713 = n58707 & ~n58712;
  assign n58714 = n58700 & n58713;
  assign n58715 = ~pi1638 & ~n58714;
  assign n58716 = pi1638 & n58707;
  assign n58717 = n58700 & n58716;
  assign n58718 = ~n58712 & n58717;
  assign po1737 = n58715 | n58718;
  assign n58720 = ~n57951 & n57972;
  assign n58721 = ~n58605 & ~n58720;
  assign n58722 = n57957 & n58721;
  assign n58723 = ~n57945 & ~n57966;
  assign n58724 = ~n57965 & ~n58723;
  assign n58725 = n57938 & n57991;
  assign n58726 = n57951 & n57966;
  assign n58727 = ~n58725 & ~n58726;
  assign n58728 = n57951 & n58009;
  assign n58729 = n58727 & ~n58728;
  assign n58730 = ~n58724 & n58729;
  assign n58731 = ~n57957 & n58730;
  assign n58732 = ~n58722 & ~n58731;
  assign n58733 = n57951 & n58724;
  assign n58734 = ~n58614 & ~n58733;
  assign n58735 = ~n58732 & n58734;
  assign n58736 = n57932 & ~n58735;
  assign n58737 = n57957 & ~n58723;
  assign n58738 = ~n57951 & n58737;
  assign n58739 = ~n57984 & ~n58013;
  assign n58740 = n57951 & ~n58739;
  assign n58741 = n57957 & n58740;
  assign n58742 = n57965 & n58737;
  assign n58743 = ~n58741 & ~n58742;
  assign n58744 = ~n58738 & n58743;
  assign n58745 = ~n57932 & ~n58744;
  assign n58746 = ~n58736 & ~n58745;
  assign n58747 = n57957 & n57970;
  assign n58748 = ~n57957 & ~n58734;
  assign n58749 = ~n58747 & ~n58748;
  assign n58750 = ~n57957 & ~n58721;
  assign n58751 = ~n57970 & ~n58750;
  assign n58752 = ~n57932 & ~n58751;
  assign n58753 = n58749 & ~n58752;
  assign n58754 = n58746 & n58753;
  assign n58755 = pi1655 & ~n58754;
  assign n58756 = ~n58736 & n58753;
  assign n58757 = ~n58745 & n58756;
  assign n58758 = ~pi1655 & n58757;
  assign po1738 = n58755 | n58758;
  assign n58760 = n58493 & n58676;
  assign n58761 = ~n58502 & ~n58760;
  assign n58762 = ~n58480 & ~n58761;
  assign n58763 = n58474 & n58525;
  assign n58764 = ~n58516 & ~n58763;
  assign n58765 = n58480 & ~n58764;
  assign n58766 = ~n58474 & n58685;
  assign n58767 = ~n58541 & ~n58766;
  assign n58768 = ~n58675 & n58767;
  assign n58769 = ~n58765 & n58768;
  assign n58770 = ~n58762 & n58769;
  assign n58771 = ~n58511 & ~n58524;
  assign n58772 = n58770 & n58771;
  assign n58773 = n58468 & ~n58772;
  assign n58774 = n58509 & n58535;
  assign n58775 = n58703 & ~n58774;
  assign n58776 = n58480 & ~n58775;
  assign n58777 = ~n58474 & n58693;
  assign n58778 = ~n58776 & ~n58777;
  assign n58779 = n58487 & n58676;
  assign n58780 = n58474 & n58501;
  assign n58781 = ~n58779 & ~n58780;
  assign n58782 = n58480 & ~n58781;
  assign n58783 = n58480 & n58525;
  assign n58784 = ~n58474 & n58783;
  assign n58785 = ~n58782 & ~n58784;
  assign n58786 = n58778 & n58785;
  assign n58787 = ~n58468 & ~n58786;
  assign n58788 = ~n58685 & ~n58690;
  assign n58789 = ~n58517 & n58788;
  assign n58790 = n58708 & ~n58789;
  assign n58791 = ~n58787 & ~n58790;
  assign n58792 = ~n58511 & ~n58675;
  assign n58793 = ~n58480 & ~n58792;
  assign n58794 = n58791 & ~n58793;
  assign n58795 = ~n58773 & n58794;
  assign n58796 = ~pi1647 & n58795;
  assign n58797 = pi1647 & ~n58795;
  assign po1740 = n58796 | n58797;
  assign n58799 = ~n58250 & n58290;
  assign n58800 = ~n58423 & ~n58799;
  assign n58801 = ~n58415 & n58800;
  assign n58802 = ~n58287 & ~n58801;
  assign n58803 = ~n58311 & ~n58322;
  assign n58804 = ~n58450 & n58803;
  assign n58805 = ~n58287 & ~n58804;
  assign n58806 = ~n58337 & n58800;
  assign n58807 = n58276 & n58287;
  assign n58808 = n58806 & ~n58807;
  assign n58809 = ~n58805 & n58808;
  assign n58810 = n58244 & ~n58809;
  assign n58811 = ~n58438 & ~n58443;
  assign n58812 = n58250 & n58297;
  assign n58813 = n58274 & n58304;
  assign n58814 = ~n58322 & ~n58813;
  assign n58815 = n58287 & ~n58814;
  assign n58816 = ~n58812 & ~n58815;
  assign n58817 = ~n58287 & n58288;
  assign n58818 = n58250 & n58817;
  assign n58819 = ~n58287 & n58295;
  assign n58820 = ~n58818 & ~n58819;
  assign n58821 = n58816 & n58820;
  assign n58822 = n58274 & n58309;
  assign n58823 = ~n58415 & ~n58822;
  assign n58824 = ~n58448 & n58823;
  assign n58825 = n58821 & n58824;
  assign n58826 = ~n58244 & ~n58825;
  assign n58827 = n58811 & ~n58826;
  assign n58828 = ~n58810 & n58827;
  assign n58829 = ~n58802 & n58828;
  assign n58830 = ~pi1648 & n58829;
  assign n58831 = pi1648 & ~n58829;
  assign po1741 = n58830 | n58831;
  assign n58833 = ~n57747 & n57780;
  assign n58834 = n57747 & n57791;
  assign n58835 = ~n57777 & ~n58834;
  assign n58836 = n57721 & ~n58835;
  assign n58837 = ~n58833 & ~n58836;
  assign n58838 = ~n57721 & ~n57747;
  assign n58839 = ~n57739 & n58838;
  assign n58840 = ~n57733 & n58839;
  assign n58841 = n57758 & n57792;
  assign n58842 = ~n58840 & ~n58841;
  assign n58843 = ~n57721 & n57756;
  assign n58844 = n58842 & ~n58843;
  assign n58845 = ~n57754 & ~n57766;
  assign n58846 = n57739 & n57800;
  assign n58847 = n58845 & ~n58846;
  assign n58848 = n58844 & n58847;
  assign n58849 = n58837 & n58848;
  assign n58850 = ~n57789 & ~n58849;
  assign n58851 = ~n57753 & ~n57777;
  assign n58852 = n57747 & ~n58851;
  assign n58853 = ~n57733 & n57795;
  assign n58854 = ~n57806 & ~n58853;
  assign n58855 = n57727 & ~n57739;
  assign n58856 = n57747 & n58855;
  assign n58857 = n58854 & ~n58856;
  assign n58858 = n57721 & ~n58857;
  assign n58859 = ~n57747 & n57776;
  assign n58860 = ~n57733 & n57765;
  assign n58861 = ~n58859 & ~n58860;
  assign n58862 = ~n57721 & ~n58861;
  assign n58863 = ~n57747 & n57759;
  assign n58864 = ~n58862 & ~n58863;
  assign n58865 = ~n58858 & n58864;
  assign n58866 = ~n58852 & n58865;
  assign n58867 = n57789 & ~n58866;
  assign n58868 = n57721 & n57796;
  assign n58869 = ~n58867 & ~n58868;
  assign n58870 = ~n57721 & n58833;
  assign n58871 = n58869 & ~n58870;
  assign n58872 = ~n58850 & n58871;
  assign n58873 = ~pi1651 & ~n58872;
  assign n58874 = pi1651 & n58869;
  assign n58875 = ~n58850 & n58874;
  assign n58876 = ~n58870 & n58875;
  assign po1742 = n58873 | n58876;
  assign n58878 = ~n57748 & ~n57757;
  assign n58879 = ~n57721 & ~n58878;
  assign n58880 = ~n57813 & ~n58879;
  assign n58881 = ~n57727 & n57733;
  assign n58882 = n57721 & n58881;
  assign n58883 = n57747 & n58882;
  assign n58884 = n57747 & n57776;
  assign n58885 = ~n58881 & ~n58884;
  assign n58886 = n57727 & ~n57747;
  assign n58887 = ~n57733 & n58886;
  assign n58888 = n58885 & ~n58887;
  assign n58889 = n57721 & ~n58888;
  assign n58890 = ~n57760 & ~n58889;
  assign n58891 = ~n57789 & ~n58890;
  assign n58892 = ~n57721 & n57740;
  assign n58893 = n57747 & n58892;
  assign n58894 = ~n58843 & ~n58893;
  assign n58895 = ~n57789 & ~n58894;
  assign n58896 = ~n58891 & ~n58895;
  assign n58897 = ~n58883 & n58896;
  assign n58898 = ~n57777 & ~n57796;
  assign n58899 = ~n57806 & n58898;
  assign n58900 = ~n57721 & ~n58899;
  assign n58901 = ~n57751 & n58886;
  assign n58902 = n57733 & n58901;
  assign n58903 = ~n57780 & ~n58902;
  assign n58904 = n57721 & ~n58903;
  assign n58905 = ~n58853 & ~n58904;
  assign n58906 = ~n58900 & n58905;
  assign n58907 = ~n57766 & ~n57807;
  assign n58908 = n58906 & n58907;
  assign n58909 = n57789 & ~n58908;
  assign n58910 = n58897 & ~n58909;
  assign n58911 = n58880 & n58910;
  assign n58912 = ~pi1671 & ~n58911;
  assign n58913 = pi1671 & n58897;
  assign n58914 = n58880 & n58913;
  assign n58915 = ~n58909 & n58914;
  assign po1744 = n58912 | n58915;
  assign n58917 = pi5293 & pi9040;
  assign n58918 = pi5576 & ~pi9040;
  assign n58919 = ~n58917 & ~n58918;
  assign n58920 = ~pi1609 & n58919;
  assign n58921 = pi1609 & ~n58919;
  assign n58922 = ~n58920 & ~n58921;
  assign n58923 = pi5399 & pi9040;
  assign n58924 = pi5566 & ~pi9040;
  assign n58925 = ~n58923 & ~n58924;
  assign n58926 = ~pi1613 & n58925;
  assign n58927 = pi1613 & ~n58925;
  assign n58928 = ~n58926 & ~n58927;
  assign n58929 = pi5313 & pi9040;
  assign n58930 = pi5319 & ~pi9040;
  assign n58931 = ~n58929 & ~n58930;
  assign n58932 = ~pi1618 & ~n58931;
  assign n58933 = pi1618 & n58931;
  assign n58934 = ~n58932 & ~n58933;
  assign n58935 = n58928 & n58934;
  assign n58936 = ~n58922 & n58935;
  assign n58937 = pi5324 & ~pi9040;
  assign n58938 = pi5502 & pi9040;
  assign n58939 = ~n58937 & ~n58938;
  assign n58940 = ~pi1610 & n58939;
  assign n58941 = pi1610 & ~n58939;
  assign n58942 = ~n58940 & ~n58941;
  assign n58943 = n58922 & ~n58942;
  assign n58944 = ~n58934 & n58943;
  assign n58945 = ~n58922 & ~n58942;
  assign n58946 = n58934 & n58945;
  assign n58947 = ~n58944 & ~n58946;
  assign n58948 = ~n58936 & n58947;
  assign n58949 = pi5303 & pi9040;
  assign n58950 = pi5321 & ~pi9040;
  assign n58951 = ~n58949 & ~n58950;
  assign n58952 = ~pi1604 & n58951;
  assign n58953 = pi1604 & ~n58951;
  assign n58954 = ~n58952 & ~n58953;
  assign n58955 = pi5508 & ~pi9040;
  assign n58956 = pi5328 & pi9040;
  assign n58957 = ~n58955 & ~n58956;
  assign n58958 = ~pi1614 & ~n58957;
  assign n58959 = pi1614 & n58957;
  assign n58960 = ~n58958 & ~n58959;
  assign n58961 = n58954 & n58960;
  assign n58962 = ~n58948 & n58961;
  assign n58963 = n58922 & n58942;
  assign n58964 = n58934 & n58963;
  assign n58965 = ~n58928 & n58960;
  assign n58966 = n58964 & n58965;
  assign n58967 = n58934 & n58943;
  assign n58968 = ~n58954 & n58967;
  assign n58969 = ~n58922 & n58942;
  assign n58970 = ~n58928 & n58969;
  assign n58971 = ~n58922 & ~n58934;
  assign n58972 = ~n58970 & ~n58971;
  assign n58973 = ~n58954 & ~n58972;
  assign n58974 = ~n58968 & ~n58973;
  assign n58975 = n58960 & ~n58974;
  assign n58976 = ~n58966 & ~n58975;
  assign n58977 = ~n58928 & ~n58934;
  assign n58978 = ~n58922 & n58977;
  assign n58979 = n58928 & ~n58934;
  assign n58980 = n58922 & n58979;
  assign n58981 = n58942 & n58980;
  assign n58982 = ~n58978 & ~n58981;
  assign n58983 = ~n58954 & ~n58982;
  assign n58984 = n58976 & ~n58983;
  assign n58985 = ~n58928 & n58954;
  assign n58986 = n58969 & n58985;
  assign n58987 = n58934 & n58986;
  assign n58988 = ~n58945 & ~n58963;
  assign n58989 = n58935 & ~n58988;
  assign n58990 = n58928 & n58944;
  assign n58991 = ~n58989 & ~n58990;
  assign n58992 = ~n58934 & n58969;
  assign n58993 = n58928 & n58954;
  assign n58994 = n58992 & n58993;
  assign n58995 = n58977 & ~n58988;
  assign n58996 = ~n58928 & n58967;
  assign n58997 = ~n58995 & ~n58996;
  assign n58998 = ~n58994 & n58997;
  assign n58999 = n58991 & n58998;
  assign n59000 = ~n58987 & n58999;
  assign n59001 = n58928 & ~n58954;
  assign n59002 = n58934 & n59001;
  assign n59003 = n58942 & n59002;
  assign n59004 = n59000 & ~n59003;
  assign n59005 = ~n58960 & ~n59004;
  assign n59006 = n58984 & ~n59005;
  assign n59007 = ~n58962 & n59006;
  assign n59008 = ~pi1681 & ~n59007;
  assign n59009 = pi1681 & n58984;
  assign n59010 = ~n58962 & n59009;
  assign n59011 = ~n59005 & n59010;
  assign po1745 = n59008 | n59011;
  assign n59013 = n58934 & n58969;
  assign n59014 = ~n58954 & n59013;
  assign n59015 = n58928 & n59014;
  assign n59016 = n58943 & n59001;
  assign n59017 = ~n58934 & n59016;
  assign n59018 = ~n59015 & ~n59017;
  assign n59019 = ~n58990 & ~n58994;
  assign n59020 = n58934 & ~n58942;
  assign n59021 = ~n58928 & n59020;
  assign n59022 = ~n58970 & ~n59021;
  assign n59023 = ~n58954 & ~n59022;
  assign n59024 = n58928 & ~n58969;
  assign n59025 = ~n58954 & n59024;
  assign n59026 = ~n58934 & n59025;
  assign n59027 = n58954 & ~n58979;
  assign n59028 = ~n58988 & n59027;
  assign n59029 = ~n59026 & ~n59028;
  assign n59030 = ~n59023 & n59029;
  assign n59031 = n59019 & n59030;
  assign n59032 = n58960 & ~n59031;
  assign n59033 = n59018 & ~n59032;
  assign n59034 = n58946 & n58954;
  assign n59035 = ~n58928 & n59034;
  assign n59036 = n58954 & ~n58960;
  assign n59037 = ~n58967 & ~n58970;
  assign n59038 = n58979 & ~n58988;
  assign n59039 = n59037 & ~n59038;
  assign n59040 = n59036 & ~n59039;
  assign n59041 = ~n58928 & n58944;
  assign n59042 = ~n58928 & ~n58942;
  assign n59043 = ~n58934 & n59042;
  assign n59044 = ~n58928 & n58963;
  assign n59045 = ~n59043 & ~n59044;
  assign n59046 = n58928 & n58969;
  assign n59047 = ~n58964 & ~n59046;
  assign n59048 = n59045 & n59047;
  assign n59049 = ~n58954 & ~n59048;
  assign n59050 = ~n59041 & ~n59049;
  assign n59051 = ~n58960 & ~n59050;
  assign n59052 = ~n59040 & ~n59051;
  assign n59053 = ~n59035 & n59052;
  assign n59054 = n59033 & n59053;
  assign n59055 = pi1673 & ~n59054;
  assign n59056 = ~pi1673 & n59033;
  assign n59057 = n59053 & n59056;
  assign po1746 = n59055 | n59057;
  assign n59059 = ~n59044 & ~n59046;
  assign n59060 = ~n58954 & ~n59059;
  assign n59061 = ~n59017 & ~n59060;
  assign n59062 = n58960 & ~n59061;
  assign n59063 = n58934 & n58960;
  assign n59064 = ~n58945 & n59063;
  assign n59065 = ~n58928 & n59064;
  assign n59066 = n58945 & n58977;
  assign n59067 = ~n58954 & n59066;
  assign n59068 = n58934 & n58985;
  assign n59069 = n58922 & n59068;
  assign n59070 = ~n59067 & ~n59069;
  assign n59071 = ~n59065 & n59070;
  assign n59072 = ~n58934 & ~n58942;
  assign n59073 = ~n58945 & ~n59072;
  assign n59074 = n58928 & ~n59073;
  assign n59075 = ~n59013 & ~n59074;
  assign n59076 = n58954 & ~n59075;
  assign n59077 = ~n59038 & ~n59076;
  assign n59078 = ~n58928 & n58992;
  assign n59079 = n58922 & n58935;
  assign n59080 = ~n58928 & ~n59073;
  assign n59081 = ~n59079 & ~n59080;
  assign n59082 = ~n58954 & ~n59081;
  assign n59083 = ~n59078 & ~n59082;
  assign n59084 = n59077 & n59083;
  assign n59085 = ~n58960 & ~n59084;
  assign n59086 = ~n58964 & ~n59042;
  assign n59087 = n58961 & ~n59086;
  assign n59088 = ~n59085 & ~n59087;
  assign n59089 = n59071 & n59088;
  assign n59090 = ~n59062 & n59089;
  assign n59091 = pi1674 & ~n59090;
  assign n59092 = ~pi1674 & n59090;
  assign po1747 = n59091 | n59092;
  assign n59094 = ~n58271 & ~n58305;
  assign n59095 = n58244 & ~n59094;
  assign n59096 = ~n58310 & ~n58427;
  assign n59097 = ~n58280 & n59096;
  assign n59098 = ~n58287 & ~n59097;
  assign n59099 = n58244 & n59098;
  assign n59100 = ~n59095 & ~n59099;
  assign n59101 = n58270 & n58424;
  assign n59102 = ~n58426 & ~n59101;
  assign n59103 = ~n58313 & ~n58451;
  assign n59104 = n58287 & ~n59103;
  assign n59105 = n58244 & n59104;
  assign n59106 = n59102 & ~n59105;
  assign n59107 = n58268 & n58309;
  assign n59108 = ~n58262 & n59107;
  assign n59109 = n58250 & n58275;
  assign n59110 = ~n58416 & ~n59109;
  assign n59111 = n58287 & ~n59110;
  assign n59112 = ~n58311 & ~n58423;
  assign n59113 = n58250 & n58269;
  assign n59114 = ~n58335 & ~n59113;
  assign n59115 = ~n58287 & ~n59114;
  assign n59116 = n59112 & ~n59115;
  assign n59117 = ~n59111 & n59116;
  assign n59118 = ~n59108 & n59117;
  assign n59119 = ~n58244 & ~n59118;
  assign n59120 = ~n58448 & n58800;
  assign n59121 = n58287 & ~n59120;
  assign n59122 = ~n59119 & ~n59121;
  assign n59123 = n59106 & n59122;
  assign n59124 = n59100 & n59123;
  assign n59125 = ~pi1650 & ~n59124;
  assign n59126 = pi1650 & n59106;
  assign n59127 = n59100 & n59126;
  assign n59128 = n59122 & n59127;
  assign po1748 = n59125 | n59128;
  assign n59130 = ~n58350 & ~n58653;
  assign n59131 = ~n58641 & n59130;
  assign n59132 = n58140 & ~n59131;
  assign n59133 = ~n58358 & ~n58649;
  assign n59134 = ~n58344 & ~n58656;
  assign n59135 = ~n58140 & ~n59134;
  assign n59136 = ~n58171 & ~n59135;
  assign n59137 = n59133 & n59136;
  assign n59138 = n58107 & ~n59137;
  assign n59139 = ~n58125 & n58131;
  assign n59140 = ~n58143 & ~n59139;
  assign n59141 = n58113 & ~n59140;
  assign n59142 = ~n58133 & ~n58364;
  assign n59143 = ~n58140 & ~n59142;
  assign n59144 = n58113 & n58131;
  assign n59145 = ~n58155 & ~n59144;
  assign n59146 = ~n58146 & n59145;
  assign n59147 = n58140 & ~n59146;
  assign n59148 = ~n59143 & ~n59147;
  assign n59149 = ~n59141 & n59148;
  assign n59150 = ~n58107 & ~n59149;
  assign n59151 = ~n59138 & ~n59150;
  assign n59152 = ~n58361 & ~n58377;
  assign n59153 = n59151 & n59152;
  assign n59154 = ~n59132 & n59153;
  assign n59155 = ~pi1654 & ~n59154;
  assign n59156 = pi1654 & n59152;
  assign n59157 = ~n59132 & n59156;
  assign n59158 = n59151 & n59157;
  assign po1749 = n59155 | n59158;
  assign n59160 = n57951 & n58616;
  assign n59161 = n57957 & n59160;
  assign n59162 = n57991 & ~n58723;
  assign n59163 = ~n58014 & ~n58614;
  assign n59164 = ~n59162 & n59163;
  assign n59165 = ~n57957 & ~n59164;
  assign n59166 = n57951 & n57967;
  assign n59167 = ~n59165 & ~n59166;
  assign n59168 = n57965 & n58013;
  assign n59169 = ~n57951 & n58606;
  assign n59170 = ~n59168 & ~n59169;
  assign n59171 = ~n58726 & n59170;
  assign n59172 = n57957 & ~n59171;
  assign n59173 = n59167 & ~n59172;
  assign n59174 = n57932 & ~n59173;
  assign n59175 = ~n59161 & ~n59174;
  assign n59176 = ~n57951 & n57966;
  assign n59177 = ~n58613 & ~n59176;
  assign n59178 = n57957 & ~n59177;
  assign n59179 = ~n58015 & ~n59178;
  assign n59180 = ~n57985 & ~n59160;
  assign n59181 = ~n57951 & n57967;
  assign n59182 = n57951 & n58020;
  assign n59183 = ~n58606 & ~n59182;
  assign n59184 = ~n59168 & n59183;
  assign n59185 = ~n57957 & ~n59184;
  assign n59186 = ~n59181 & ~n59185;
  assign n59187 = n59180 & n59186;
  assign n59188 = n59179 & n59187;
  assign n59189 = ~n57932 & ~n59188;
  assign n59190 = ~n57997 & ~n58728;
  assign n59191 = ~n57957 & ~n59190;
  assign n59192 = ~n59189 & ~n59191;
  assign n59193 = n59175 & n59192;
  assign n59194 = pi1653 & n59193;
  assign n59195 = ~pi1653 & ~n59193;
  assign po1750 = n59194 | n59195;
  assign n59197 = ~n58934 & n59044;
  assign n59198 = ~n58996 & ~n59197;
  assign n59199 = ~n58954 & ~n59198;
  assign n59200 = ~n58934 & n58945;
  assign n59201 = ~n59013 & ~n59200;
  assign n59202 = ~n58954 & ~n59201;
  assign n59203 = n58928 & n58963;
  assign n59204 = ~n58946 & ~n59203;
  assign n59205 = ~n58992 & n59204;
  assign n59206 = n58954 & ~n59205;
  assign n59207 = ~n59202 & ~n59206;
  assign n59208 = ~n58968 & ~n58981;
  assign n59209 = n59207 & n59208;
  assign n59210 = ~n58960 & ~n59209;
  assign n59211 = ~n58928 & n59013;
  assign n59212 = n58928 & n58943;
  assign n59213 = ~n59044 & ~n59212;
  assign n59214 = n58954 & ~n59213;
  assign n59215 = ~n59211 & ~n59214;
  assign n59216 = n58934 & ~n58954;
  assign n59217 = n58922 & n59216;
  assign n59218 = n58942 & n59217;
  assign n59219 = n58947 & ~n59218;
  assign n59220 = ~n58992 & n59219;
  assign n59221 = n58928 & ~n59220;
  assign n59222 = n59215 & ~n59221;
  assign n59223 = n58960 & ~n59222;
  assign n59224 = ~n59210 & ~n59223;
  assign n59225 = n58985 & n59072;
  assign n59226 = n59224 & ~n59225;
  assign n59227 = ~n59199 & n59226;
  assign n59228 = ~pi1649 & ~n59227;
  assign n59229 = pi1649 & ~n59199;
  assign n59230 = n59224 & n59229;
  assign n59231 = ~n59225 & n59230;
  assign po1751 = n59228 | n59231;
  assign n59233 = ~n57807 & ~n58863;
  assign n59234 = n57721 & ~n59233;
  assign n59235 = ~n57754 & ~n57757;
  assign n59236 = ~n57747 & n57806;
  assign n59237 = ~n58834 & ~n59236;
  assign n59238 = n59235 & n59237;
  assign n59239 = ~n57721 & ~n59238;
  assign n59240 = ~n57789 & n57791;
  assign n59241 = ~n57721 & n59240;
  assign n59242 = n57733 & n58886;
  assign n59243 = ~n58855 & ~n59242;
  assign n59244 = ~n57759 & n59243;
  assign n59245 = n57721 & ~n59244;
  assign n59246 = ~n57727 & n57776;
  assign n59247 = ~n57747 & n59246;
  assign n59248 = ~n59245 & ~n59247;
  assign n59249 = ~n57789 & ~n59248;
  assign n59250 = ~n59241 & ~n59249;
  assign n59251 = ~n57727 & ~n57733;
  assign n59252 = ~n57721 & n59251;
  assign n59253 = n57747 & n59252;
  assign n59254 = ~n57747 & n58855;
  assign n59255 = ~n57757 & ~n59254;
  assign n59256 = ~n58860 & n59255;
  assign n59257 = ~n59253 & n59256;
  assign n59258 = n57721 & n57753;
  assign n59259 = n59257 & ~n59258;
  assign n59260 = n57789 & ~n59259;
  assign n59261 = n59250 & ~n59260;
  assign n59262 = ~n59239 & n59261;
  assign n59263 = ~n59234 & n59262;
  assign n59264 = pi1682 & n59263;
  assign n59265 = ~pi1682 & ~n59263;
  assign po1752 = n59264 | n59265;
  assign n59267 = ~n58474 & n58501;
  assign n59268 = ~n58682 & ~n59267;
  assign n59269 = ~n58480 & ~n59268;
  assign n59270 = n58480 & ~n58543;
  assign n59271 = ~n58531 & ~n59270;
  assign n59272 = ~n59269 & n59271;
  assign n59273 = n58468 & ~n59272;
  assign n59274 = ~n58480 & n58693;
  assign n59275 = ~n59273 & ~n59274;
  assign n59276 = ~n58766 & ~n58780;
  assign n59277 = n58480 & ~n59276;
  assign n59278 = n58480 & n58683;
  assign n59279 = n58474 & n58502;
  assign n59280 = ~n58480 & n58522;
  assign n59281 = ~n58515 & ~n59280;
  assign n59282 = ~n58487 & ~n59281;
  assign n59283 = ~n58516 & ~n59282;
  assign n59284 = ~n58675 & n59283;
  assign n59285 = ~n59279 & n59284;
  assign n59286 = ~n59278 & n59285;
  assign n59287 = ~n58468 & ~n59286;
  assign n59288 = ~n59277 & ~n59287;
  assign n59289 = n59275 & n59288;
  assign n59290 = pi1666 & ~n59289;
  assign n59291 = ~pi1666 & n59289;
  assign po1753 = n59290 | n59291;
  assign n59293 = pi5697 & ~pi9040;
  assign n59294 = pi5704 & pi9040;
  assign n59295 = ~n59293 & ~n59294;
  assign n59296 = ~pi1657 & ~n59295;
  assign n59297 = pi1657 & n59295;
  assign n59298 = ~n59296 & ~n59297;
  assign n59299 = pi5783 & pi9040;
  assign n59300 = pi5695 & ~pi9040;
  assign n59301 = ~n59299 & ~n59300;
  assign n59302 = ~pi1668 & n59301;
  assign n59303 = pi1668 & ~n59301;
  assign n59304 = ~n59302 & ~n59303;
  assign n59305 = pi5666 & pi9040;
  assign n59306 = pi5572 & ~pi9040;
  assign n59307 = ~n59305 & ~n59306;
  assign n59308 = ~pi1684 & n59307;
  assign n59309 = pi1684 & ~n59307;
  assign n59310 = ~n59308 & ~n59309;
  assign n59311 = pi5579 & ~pi9040;
  assign n59312 = pi5669 & pi9040;
  assign n59313 = ~n59311 & ~n59312;
  assign n59314 = ~pi1665 & n59313;
  assign n59315 = pi1665 & ~n59313;
  assign n59316 = ~n59314 & ~n59315;
  assign n59317 = ~n59310 & ~n59316;
  assign n59318 = n59304 & n59317;
  assign n59319 = pi5577 & pi9040;
  assign n59320 = pi5782 & ~pi9040;
  assign n59321 = ~n59319 & ~n59320;
  assign n59322 = pi1694 & n59321;
  assign n59323 = ~pi1694 & ~n59321;
  assign n59324 = ~n59322 & ~n59323;
  assign n59325 = n59318 & ~n59324;
  assign n59326 = n59310 & n59316;
  assign n59327 = n59304 & n59326;
  assign n59328 = ~n59324 & n59327;
  assign n59329 = ~n59325 & ~n59328;
  assign n59330 = ~n59304 & n59324;
  assign n59331 = n59326 & n59330;
  assign n59332 = ~n59310 & n59316;
  assign n59333 = n59304 & n59332;
  assign n59334 = n59324 & n59333;
  assign n59335 = ~n59331 & ~n59334;
  assign n59336 = n59329 & n59335;
  assign n59337 = n59298 & ~n59336;
  assign n59338 = n59304 & n59324;
  assign n59339 = ~n59316 & n59338;
  assign n59340 = n59310 & n59339;
  assign n59341 = ~n59333 & ~n59340;
  assign n59342 = n59298 & ~n59341;
  assign n59343 = ~n59298 & ~n59316;
  assign n59344 = ~n59324 & n59343;
  assign n59345 = ~n59304 & ~n59310;
  assign n59346 = n59324 & n59326;
  assign n59347 = ~n59345 & ~n59346;
  assign n59348 = ~n59298 & ~n59347;
  assign n59349 = ~n59344 & ~n59348;
  assign n59350 = n59310 & ~n59316;
  assign n59351 = ~n59304 & n59350;
  assign n59352 = ~n59324 & n59351;
  assign n59353 = n59349 & ~n59352;
  assign n59354 = ~n59316 & n59345;
  assign n59355 = n59324 & n59354;
  assign n59356 = n59353 & ~n59355;
  assign n59357 = ~n59342 & n59356;
  assign n59358 = pi5555 & pi9040;
  assign n59359 = pi5672 & ~pi9040;
  assign n59360 = ~n59358 & ~n59359;
  assign n59361 = ~pi1689 & ~n59360;
  assign n59362 = pi1689 & n59360;
  assign n59363 = ~n59361 & ~n59362;
  assign n59364 = ~n59357 & ~n59363;
  assign n59365 = n59304 & ~n59316;
  assign n59366 = ~n59298 & n59324;
  assign n59367 = n59363 & n59366;
  assign n59368 = n59365 & n59367;
  assign n59369 = n59304 & ~n59324;
  assign n59370 = n59316 & n59369;
  assign n59371 = ~n59298 & ~n59370;
  assign n59372 = n59310 & n59330;
  assign n59373 = ~n59317 & ~n59365;
  assign n59374 = ~n59324 & ~n59373;
  assign n59375 = ~n59304 & n59326;
  assign n59376 = n59298 & ~n59375;
  assign n59377 = ~n59374 & n59376;
  assign n59378 = ~n59372 & n59377;
  assign n59379 = ~n59371 & ~n59378;
  assign n59380 = ~n59304 & n59332;
  assign n59381 = n59324 & n59380;
  assign n59382 = ~n59379 & ~n59381;
  assign n59383 = n59363 & ~n59382;
  assign n59384 = ~n59368 & ~n59383;
  assign n59385 = ~n59364 & n59384;
  assign n59386 = ~n59337 & n59385;
  assign n59387 = ~n59298 & n59352;
  assign n59388 = n59386 & ~n59387;
  assign n59389 = pi1696 & ~n59388;
  assign n59390 = ~n59337 & ~n59387;
  assign n59391 = n59385 & n59390;
  assign n59392 = ~pi1696 & n59391;
  assign po1777 = n59389 | n59392;
  assign n59394 = pi5579 & pi9040;
  assign n59395 = pi5696 & ~pi9040;
  assign n59396 = ~n59394 & ~n59395;
  assign n59397 = pi1676 & n59396;
  assign n59398 = ~pi1676 & ~n59396;
  assign n59399 = ~n59397 & ~n59398;
  assign n59400 = pi5666 & ~pi9040;
  assign n59401 = pi5780 & pi9040;
  assign n59402 = ~n59400 & ~n59401;
  assign n59403 = pi1691 & n59402;
  assign n59404 = ~pi1691 & ~n59402;
  assign n59405 = ~n59403 & ~n59404;
  assign n59406 = pi5783 & ~pi9040;
  assign n59407 = pi5785 & pi9040;
  assign n59408 = ~n59406 & ~n59407;
  assign n59409 = pi1690 & n59408;
  assign n59410 = ~pi1690 & ~n59408;
  assign n59411 = ~n59409 & ~n59410;
  assign n59412 = pi5664 & pi9040;
  assign n59413 = pi5588 & ~pi9040;
  assign n59414 = ~n59412 & ~n59413;
  assign n59415 = pi1659 & n59414;
  assign n59416 = ~pi1659 & ~n59414;
  assign n59417 = ~n59415 & ~n59416;
  assign n59418 = pi5557 & ~pi9040;
  assign n59419 = pi5571 & pi9040;
  assign n59420 = ~n59418 & ~n59419;
  assign n59421 = pi1685 & n59420;
  assign n59422 = ~pi1685 & ~n59420;
  assign n59423 = ~n59421 & ~n59422;
  assign n59424 = n59417 & ~n59423;
  assign n59425 = n59411 & n59424;
  assign n59426 = n59405 & n59425;
  assign n59427 = ~n59405 & n59417;
  assign n59428 = n59423 & n59427;
  assign n59429 = pi5582 & ~pi9040;
  assign n59430 = pi5697 & pi9040;
  assign n59431 = ~n59429 & ~n59430;
  assign n59432 = ~pi1680 & ~n59431;
  assign n59433 = pi1680 & n59431;
  assign n59434 = ~n59432 & ~n59433;
  assign n59435 = ~n59411 & n59427;
  assign n59436 = n59411 & n59423;
  assign n59437 = ~n59417 & n59436;
  assign n59438 = ~n59435 & ~n59437;
  assign n59439 = ~n59434 & ~n59438;
  assign n59440 = ~n59428 & ~n59439;
  assign n59441 = n59417 & n59436;
  assign n59442 = ~n59417 & ~n59423;
  assign n59443 = ~n59405 & n59442;
  assign n59444 = ~n59411 & ~n59423;
  assign n59445 = n59405 & n59444;
  assign n59446 = ~n59443 & ~n59445;
  assign n59447 = ~n59411 & ~n59417;
  assign n59448 = n59446 & ~n59447;
  assign n59449 = ~n59441 & n59448;
  assign n59450 = n59434 & ~n59449;
  assign n59451 = n59440 & ~n59450;
  assign n59452 = ~n59426 & n59451;
  assign n59453 = n59399 & ~n59452;
  assign n59454 = ~n59411 & n59423;
  assign n59455 = ~n59417 & n59454;
  assign n59456 = ~n59405 & n59455;
  assign n59457 = ~n59417 & n59444;
  assign n59458 = n59405 & n59457;
  assign n59459 = ~n59426 & ~n59458;
  assign n59460 = ~n59456 & n59459;
  assign n59461 = n59434 & ~n59460;
  assign n59462 = ~n59453 & ~n59461;
  assign n59463 = n59411 & n59428;
  assign n59464 = n59411 & ~n59417;
  assign n59465 = ~n59434 & n59464;
  assign n59466 = n59405 & n59465;
  assign n59467 = ~n59405 & n59434;
  assign n59468 = n59417 & n59467;
  assign n59469 = ~n59423 & n59468;
  assign n59470 = n59417 & n59454;
  assign n59471 = n59405 & n59470;
  assign n59472 = ~n59469 & ~n59471;
  assign n59473 = ~n59411 & n59417;
  assign n59474 = n59405 & n59473;
  assign n59475 = n59411 & ~n59423;
  assign n59476 = ~n59417 & n59475;
  assign n59477 = ~n59474 & ~n59476;
  assign n59478 = ~n59434 & ~n59477;
  assign n59479 = ~n59411 & ~n59434;
  assign n59480 = ~n59417 & n59479;
  assign n59481 = ~n59405 & n59480;
  assign n59482 = ~n59478 & ~n59481;
  assign n59483 = n59472 & n59482;
  assign n59484 = ~n59399 & ~n59483;
  assign n59485 = ~n59466 & ~n59484;
  assign n59486 = ~n59463 & n59485;
  assign n59487 = n59462 & n59486;
  assign n59488 = ~pi1703 & ~n59487;
  assign n59489 = ~n59453 & ~n59463;
  assign n59490 = ~n59461 & n59489;
  assign n59491 = n59485 & n59490;
  assign n59492 = pi1703 & n59491;
  assign po1779 = n59488 | n59492;
  assign n59494 = pi5702 & pi9040;
  assign n59495 = pi5705 & ~pi9040;
  assign n59496 = ~n59494 & ~n59495;
  assign n59497 = ~pi1665 & ~n59496;
  assign n59498 = pi1665 & n59496;
  assign n59499 = ~n59497 & ~n59498;
  assign n59500 = pi5701 & pi9040;
  assign n59501 = pi5661 & ~pi9040;
  assign n59502 = ~n59500 & ~n59501;
  assign n59503 = ~pi1693 & n59502;
  assign n59504 = pi1693 & ~n59502;
  assign n59505 = ~n59503 & ~n59504;
  assign n59506 = pi5574 & ~pi9040;
  assign n59507 = pi5588 & pi9040;
  assign n59508 = ~n59506 & ~n59507;
  assign n59509 = pi1668 & n59508;
  assign n59510 = ~pi1668 & ~n59508;
  assign n59511 = ~n59509 & ~n59510;
  assign n59512 = n59505 & n59511;
  assign n59513 = pi5554 & ~pi9040;
  assign n59514 = pi5699 & pi9040;
  assign n59515 = ~n59513 & ~n59514;
  assign n59516 = pi1670 & n59515;
  assign n59517 = ~pi1670 & ~n59515;
  assign n59518 = ~n59516 & ~n59517;
  assign n59519 = pi5555 & ~pi9040;
  assign n59520 = pi5557 & pi9040;
  assign n59521 = ~n59519 & ~n59520;
  assign n59522 = pi1686 & n59521;
  assign n59523 = ~pi1686 & ~n59521;
  assign n59524 = ~n59522 & ~n59523;
  assign n59525 = ~n59518 & ~n59524;
  assign n59526 = n59512 & n59525;
  assign n59527 = pi5577 & ~pi9040;
  assign n59528 = pi5784 & pi9040;
  assign n59529 = ~n59527 & ~n59528;
  assign n59530 = ~pi1664 & n59529;
  assign n59531 = pi1664 & ~n59529;
  assign n59532 = ~n59530 & ~n59531;
  assign n59533 = ~n59505 & ~n59511;
  assign n59534 = ~n59532 & n59533;
  assign n59535 = n59518 & n59532;
  assign n59536 = ~n59511 & n59535;
  assign n59537 = n59505 & n59536;
  assign n59538 = ~n59534 & ~n59537;
  assign n59539 = ~n59505 & n59511;
  assign n59540 = n59518 & n59539;
  assign n59541 = n59538 & ~n59540;
  assign n59542 = ~n59524 & ~n59541;
  assign n59543 = ~n59505 & n59532;
  assign n59544 = ~n59518 & n59524;
  assign n59545 = n59543 & n59544;
  assign n59546 = n59532 & n59533;
  assign n59547 = ~n59518 & n59546;
  assign n59548 = ~n59545 & ~n59547;
  assign n59549 = ~n59542 & n59548;
  assign n59550 = ~n59526 & n59549;
  assign n59551 = n59512 & ~n59532;
  assign n59552 = ~n59518 & n59551;
  assign n59553 = ~n59532 & n59539;
  assign n59554 = n59518 & n59553;
  assign n59555 = ~n59552 & ~n59554;
  assign n59556 = n59550 & n59555;
  assign n59557 = ~n59499 & ~n59556;
  assign n59558 = ~n59518 & n59532;
  assign n59559 = n59511 & n59558;
  assign n59560 = ~n59505 & n59559;
  assign n59561 = ~n59551 & ~n59560;
  assign n59562 = ~n59524 & ~n59561;
  assign n59563 = n59512 & n59535;
  assign n59564 = n59505 & ~n59511;
  assign n59565 = n59558 & n59564;
  assign n59566 = ~n59563 & ~n59565;
  assign n59567 = ~n59505 & n59535;
  assign n59568 = ~n59518 & n59553;
  assign n59569 = ~n59567 & ~n59568;
  assign n59570 = n59524 & ~n59569;
  assign n59571 = n59566 & ~n59570;
  assign n59572 = ~n59562 & n59571;
  assign n59573 = n59499 & ~n59572;
  assign n59574 = ~n59505 & ~n59532;
  assign n59575 = n59518 & n59574;
  assign n59576 = n59505 & ~n59532;
  assign n59577 = ~n59518 & n59576;
  assign n59578 = ~n59575 & ~n59577;
  assign n59579 = ~n59524 & ~n59578;
  assign n59580 = ~n59532 & n59564;
  assign n59581 = n59518 & n59580;
  assign n59582 = ~n59563 & ~n59581;
  assign n59583 = ~n59546 & n59582;
  assign n59584 = n59524 & ~n59583;
  assign n59585 = ~n59579 & ~n59584;
  assign n59586 = ~n59511 & n59532;
  assign n59587 = n59524 & n59586;
  assign n59588 = ~n59518 & n59587;
  assign n59589 = n59585 & ~n59588;
  assign n59590 = ~n59573 & n59589;
  assign n59591 = ~n59557 & n59590;
  assign n59592 = ~pi1697 & ~n59591;
  assign n59593 = pi1697 & n59591;
  assign po1784 = n59592 | n59593;
  assign n59595 = pi5561 & pi9040;
  assign n59596 = pi5700 & ~pi9040;
  assign n59597 = ~n59595 & ~n59596;
  assign n59598 = ~pi1690 & ~n59597;
  assign n59599 = pi1690 & n59597;
  assign n59600 = ~n59598 & ~n59599;
  assign n59601 = pi5578 & ~pi9040;
  assign n59602 = pi5663 & pi9040;
  assign n59603 = ~n59601 & ~n59602;
  assign n59604 = ~pi1663 & n59603;
  assign n59605 = pi1663 & ~n59603;
  assign n59606 = ~n59604 & ~n59605;
  assign n59607 = pi5834 & ~pi9040;
  assign n59608 = pi5671 & pi9040;
  assign n59609 = ~n59607 & ~n59608;
  assign n59610 = ~pi1678 & n59609;
  assign n59611 = pi1678 & ~n59609;
  assign n59612 = ~n59610 & ~n59611;
  assign n59613 = pi5919 & pi9040;
  assign n59614 = pi5667 & ~pi9040;
  assign n59615 = ~n59613 & ~n59614;
  assign n59616 = pi1677 & n59615;
  assign n59617 = ~pi1677 & ~n59615;
  assign n59618 = ~n59616 & ~n59617;
  assign n59619 = pi5575 & pi9040;
  assign n59620 = pi5677 & ~pi9040;
  assign n59621 = ~n59619 & ~n59620;
  assign n59622 = pi1659 & n59621;
  assign n59623 = ~pi1659 & ~n59621;
  assign n59624 = ~n59622 & ~n59623;
  assign n59625 = ~n59618 & n59624;
  assign n59626 = ~n59612 & n59625;
  assign n59627 = ~n59606 & n59626;
  assign n59628 = pi5564 & ~pi9040;
  assign n59629 = pi5553 & pi9040;
  assign n59630 = ~n59628 & ~n59629;
  assign n59631 = ~pi1692 & ~n59630;
  assign n59632 = pi1692 & n59630;
  assign n59633 = ~n59631 & ~n59632;
  assign n59634 = ~pi1677 & n59615;
  assign n59635 = pi1677 & ~n59615;
  assign n59636 = ~n59634 & ~n59635;
  assign n59637 = n59624 & ~n59636;
  assign n59638 = ~n59606 & n59637;
  assign n59639 = n59612 & n59625;
  assign n59640 = n59606 & n59639;
  assign n59641 = ~n59638 & ~n59640;
  assign n59642 = ~n59633 & ~n59641;
  assign n59643 = ~n59627 & ~n59642;
  assign n59644 = ~n59618 & ~n59624;
  assign n59645 = n59612 & n59644;
  assign n59646 = n59633 & n59645;
  assign n59647 = n59625 & n59633;
  assign n59648 = ~n59606 & n59647;
  assign n59649 = ~n59646 & ~n59648;
  assign n59650 = n59643 & n59649;
  assign n59651 = ~n59624 & ~n59636;
  assign n59652 = ~n59612 & n59651;
  assign n59653 = ~n59606 & n59652;
  assign n59654 = ~n59612 & n59644;
  assign n59655 = n59606 & n59654;
  assign n59656 = ~n59653 & ~n59655;
  assign n59657 = n59650 & n59656;
  assign n59658 = n59600 & ~n59657;
  assign n59659 = ~n59600 & ~n59633;
  assign n59660 = ~n59606 & n59612;
  assign n59661 = n59636 & n59660;
  assign n59662 = n59612 & ~n59624;
  assign n59663 = ~n59661 & ~n59662;
  assign n59664 = n59659 & ~n59663;
  assign n59665 = n59606 & ~n59612;
  assign n59666 = n59624 & n59665;
  assign n59667 = ~n59618 & n59666;
  assign n59668 = n59606 & ~n59636;
  assign n59669 = n59612 & n59668;
  assign n59670 = ~n59667 & ~n59669;
  assign n59671 = ~n59606 & n59633;
  assign n59672 = ~n59612 & n59671;
  assign n59673 = ~n59625 & n59672;
  assign n59674 = n59633 & n59652;
  assign n59675 = ~n59673 & ~n59674;
  assign n59676 = n59670 & n59675;
  assign n59677 = ~n59600 & ~n59676;
  assign n59678 = n59612 & n59651;
  assign n59679 = ~n59633 & n59678;
  assign n59680 = n59606 & n59679;
  assign n59681 = ~n59612 & n59637;
  assign n59682 = n59606 & n59681;
  assign n59683 = ~n59655 & ~n59682;
  assign n59684 = ~n59633 & ~n59683;
  assign n59685 = ~n59680 & ~n59684;
  assign n59686 = n59633 & n59667;
  assign n59687 = n59685 & ~n59686;
  assign n59688 = ~n59677 & n59687;
  assign n59689 = ~n59664 & n59688;
  assign n59690 = ~n59658 & n59689;
  assign n59691 = n59612 & n59637;
  assign n59692 = n59606 & n59633;
  assign n59693 = n59691 & n59692;
  assign n59694 = n59690 & ~n59693;
  assign n59695 = ~pi1712 & ~n59694;
  assign n59696 = ~n59658 & ~n59693;
  assign n59697 = n59689 & n59696;
  assign n59698 = pi1712 & n59697;
  assign po1785 = n59695 | n59698;
  assign n59700 = pi5671 & ~pi9040;
  assign n59701 = pi5698 & pi9040;
  assign n59702 = ~n59700 & ~n59701;
  assign n59703 = pi1688 & n59702;
  assign n59704 = ~pi1688 & ~n59702;
  assign n59705 = ~n59703 & ~n59704;
  assign n59706 = pi5677 & pi9040;
  assign n59707 = pi5559 & ~pi9040;
  assign n59708 = ~n59706 & ~n59707;
  assign n59709 = ~pi1683 & ~n59708;
  assign n59710 = pi1683 & n59708;
  assign n59711 = ~n59709 & ~n59710;
  assign n59712 = pi5826 & pi9040;
  assign n59713 = pi5569 & ~pi9040;
  assign n59714 = ~n59712 & ~n59713;
  assign n59715 = pi1672 & n59714;
  assign n59716 = ~pi1672 & ~n59714;
  assign n59717 = ~n59715 & ~n59716;
  assign n59718 = n59711 & ~n59717;
  assign n59719 = pi5568 & pi9040;
  assign n59720 = pi5919 & ~pi9040;
  assign n59721 = ~n59719 & ~n59720;
  assign n59722 = ~pi1695 & ~n59721;
  assign n59723 = pi1695 & n59721;
  assign n59724 = ~n59722 & ~n59723;
  assign n59725 = pi5563 & ~pi9040;
  assign n59726 = pi5578 & pi9040;
  assign n59727 = ~n59725 & ~n59726;
  assign n59728 = ~pi1652 & ~n59727;
  assign n59729 = pi1652 & n59727;
  assign n59730 = ~n59728 & ~n59729;
  assign n59731 = n59724 & n59730;
  assign n59732 = n59718 & n59731;
  assign n59733 = n59724 & ~n59730;
  assign n59734 = ~n59711 & n59733;
  assign n59735 = ~n59732 & ~n59734;
  assign n59736 = ~n59705 & ~n59735;
  assign n59737 = pi5564 & pi9040;
  assign n59738 = ~pi5567 & ~pi9040;
  assign n59739 = ~n59737 & ~n59738;
  assign n59740 = ~pi1662 & ~n59739;
  assign n59741 = pi1662 & n59739;
  assign n59742 = ~n59740 & ~n59741;
  assign n59743 = n59705 & ~n59724;
  assign n59744 = n59711 & n59743;
  assign n59745 = n59718 & ~n59730;
  assign n59746 = n59711 & n59717;
  assign n59747 = n59730 & n59746;
  assign n59748 = ~n59745 & ~n59747;
  assign n59749 = ~n59711 & ~n59717;
  assign n59750 = n59730 & n59749;
  assign n59751 = n59724 & n59750;
  assign n59752 = n59748 & ~n59751;
  assign n59753 = n59705 & ~n59752;
  assign n59754 = ~n59744 & ~n59753;
  assign n59755 = ~n59711 & n59717;
  assign n59756 = ~n59730 & n59755;
  assign n59757 = n59724 & n59756;
  assign n59758 = n59754 & ~n59757;
  assign n59759 = ~n59724 & n59749;
  assign n59760 = n59730 & n59755;
  assign n59761 = ~n59759 & ~n59760;
  assign n59762 = ~n59705 & ~n59761;
  assign n59763 = ~n59730 & n59746;
  assign n59764 = ~n59724 & n59763;
  assign n59765 = ~n59762 & ~n59764;
  assign n59766 = n59758 & n59765;
  assign n59767 = n59742 & ~n59766;
  assign n59768 = ~n59736 & ~n59767;
  assign n59769 = n59705 & ~n59742;
  assign n59770 = ~n59761 & n59769;
  assign n59771 = ~n59730 & n59749;
  assign n59772 = ~n59763 & ~n59771;
  assign n59773 = n59724 & ~n59772;
  assign n59774 = ~n59732 & ~n59773;
  assign n59775 = ~n59742 & ~n59774;
  assign n59776 = ~n59770 & ~n59775;
  assign n59777 = ~n59705 & ~n59742;
  assign n59778 = n59718 & ~n59724;
  assign n59779 = ~n59756 & ~n59778;
  assign n59780 = n59711 & n59730;
  assign n59781 = n59779 & ~n59780;
  assign n59782 = n59777 & ~n59781;
  assign n59783 = n59776 & ~n59782;
  assign n59784 = n59768 & n59783;
  assign n59785 = ~pi1700 & ~n59784;
  assign n59786 = pi1700 & n59776;
  assign n59787 = n59768 & n59786;
  assign n59788 = ~n59782 & n59787;
  assign po1786 = n59785 | n59788;
  assign n59790 = pi5563 & pi9040;
  assign n59791 = pi5575 & ~pi9040;
  assign n59792 = ~n59790 & ~n59791;
  assign n59793 = ~pi1683 & ~n59792;
  assign n59794 = pi1683 & n59792;
  assign n59795 = ~n59793 & ~n59794;
  assign n59796 = pi5706 & ~pi9040;
  assign n59797 = pi5667 & pi9040;
  assign n59798 = ~n59796 & ~n59797;
  assign n59799 = pi1684 & n59798;
  assign n59800 = ~pi1684 & ~n59798;
  assign n59801 = ~n59799 & ~n59800;
  assign n59802 = pi5568 & ~pi9040;
  assign n59803 = pi5700 & pi9040;
  assign n59804 = ~n59802 & ~n59803;
  assign n59805 = ~pi1689 & ~n59804;
  assign n59806 = pi1689 & n59804;
  assign n59807 = ~n59805 & ~n59806;
  assign n59808 = pi5698 & ~pi9040;
  assign n59809 = pi5581 & pi9040;
  assign n59810 = ~n59808 & ~n59809;
  assign n59811 = ~pi1652 & n59810;
  assign n59812 = pi1652 & ~n59810;
  assign n59813 = ~n59811 & ~n59812;
  assign n59814 = ~n59807 & ~n59813;
  assign n59815 = pi5569 & pi9040;
  assign n59816 = pi5830 & ~pi9040;
  assign n59817 = ~n59815 & ~n59816;
  assign n59818 = ~pi1661 & n59817;
  assign n59819 = pi1661 & ~n59817;
  assign n59820 = ~n59818 & ~n59819;
  assign n59821 = pi5558 & ~pi9040;
  assign n59822 = pi5779 & pi9040;
  assign n59823 = ~n59821 & ~n59822;
  assign n59824 = ~pi1687 & ~n59823;
  assign n59825 = pi1687 & n59823;
  assign n59826 = ~n59824 & ~n59825;
  assign n59827 = ~n59820 & n59826;
  assign n59828 = n59814 & n59827;
  assign n59829 = n59801 & n59828;
  assign n59830 = n59820 & n59826;
  assign n59831 = n59807 & ~n59813;
  assign n59832 = n59830 & n59831;
  assign n59833 = n59801 & n59820;
  assign n59834 = n59813 & n59833;
  assign n59835 = ~n59807 & n59834;
  assign n59836 = n59807 & n59813;
  assign n59837 = n59801 & n59836;
  assign n59838 = n59826 & n59837;
  assign n59839 = ~n59820 & n59838;
  assign n59840 = ~n59835 & ~n59839;
  assign n59841 = ~n59832 & n59840;
  assign n59842 = ~n59829 & n59841;
  assign n59843 = ~n59801 & n59820;
  assign n59844 = n59831 & n59843;
  assign n59845 = n59842 & ~n59844;
  assign n59846 = ~n59795 & ~n59845;
  assign n59847 = ~n59801 & n59813;
  assign n59848 = n59807 & n59847;
  assign n59849 = ~n59826 & n59848;
  assign n59850 = ~n59820 & n59849;
  assign n59851 = ~n59807 & n59833;
  assign n59852 = ~n59807 & n59813;
  assign n59853 = n59820 & n59852;
  assign n59854 = ~n59851 & ~n59853;
  assign n59855 = ~n59826 & ~n59854;
  assign n59856 = ~n59850 & ~n59855;
  assign n59857 = ~n59795 & ~n59856;
  assign n59858 = n59801 & n59807;
  assign n59859 = ~n59813 & n59858;
  assign n59860 = ~n59820 & n59859;
  assign n59861 = ~n59834 & ~n59860;
  assign n59862 = ~n59801 & n59814;
  assign n59863 = ~n59820 & n59862;
  assign n59864 = n59861 & ~n59863;
  assign n59865 = ~n59826 & ~n59864;
  assign n59866 = ~n59857 & ~n59865;
  assign n59867 = ~n59846 & n59866;
  assign n59868 = ~n59801 & ~n59820;
  assign n59869 = n59826 & n59868;
  assign n59870 = n59852 & n59869;
  assign n59871 = ~n59801 & n59807;
  assign n59872 = n59830 & n59871;
  assign n59873 = n59801 & ~n59826;
  assign n59874 = n59807 & n59873;
  assign n59875 = ~n59807 & ~n59820;
  assign n59876 = ~n59801 & n59875;
  assign n59877 = ~n59874 & ~n59876;
  assign n59878 = n59820 & n59848;
  assign n59879 = n59877 & ~n59878;
  assign n59880 = ~n59862 & n59879;
  assign n59881 = n59814 & n59826;
  assign n59882 = n59820 & n59881;
  assign n59883 = ~n59820 & n59852;
  assign n59884 = ~n59801 & ~n59813;
  assign n59885 = ~n59883 & ~n59884;
  assign n59886 = n59826 & ~n59885;
  assign n59887 = ~n59882 & ~n59886;
  assign n59888 = n59880 & n59887;
  assign n59889 = n59795 & ~n59888;
  assign n59890 = ~n59872 & ~n59889;
  assign n59891 = ~n59870 & n59890;
  assign n59892 = n59867 & n59891;
  assign n59893 = pi1708 & n59892;
  assign n59894 = ~pi1708 & ~n59892;
  assign po1789 = n59893 | n59894;
  assign n59896 = pi5572 & pi9040;
  assign n59897 = pi5702 & ~pi9040;
  assign n59898 = ~n59896 & ~n59897;
  assign n59899 = ~pi1693 & ~n59898;
  assign n59900 = pi1693 & n59898;
  assign n59901 = ~n59899 & ~n59900;
  assign n59902 = pi5669 & ~pi9040;
  assign n59903 = pi5661 & pi9040;
  assign n59904 = ~n59902 & ~n59903;
  assign n59905 = ~pi1669 & ~n59904;
  assign n59906 = pi1669 & n59904;
  assign n59907 = ~n59905 & ~n59906;
  assign n59908 = pi5664 & ~pi9040;
  assign n59909 = pi5782 & pi9040;
  assign n59910 = ~n59908 & ~n59909;
  assign n59911 = pi1667 & n59910;
  assign n59912 = ~pi1667 & ~n59910;
  assign n59913 = ~n59911 & ~n59912;
  assign n59914 = pi5785 & ~pi9040;
  assign n59915 = pi5554 & pi9040;
  assign n59916 = ~n59914 & ~n59915;
  assign n59917 = ~pi1685 & ~n59916;
  assign n59918 = pi1685 & n59916;
  assign n59919 = ~n59917 & ~n59918;
  assign n59920 = pi5672 & pi9040;
  assign n59921 = pi5780 & ~pi9040;
  assign n59922 = ~n59920 & ~n59921;
  assign n59923 = ~pi1676 & n59922;
  assign n59924 = pi1676 & ~n59922;
  assign n59925 = ~n59923 & ~n59924;
  assign n59926 = n59919 & n59925;
  assign n59927 = n59913 & n59926;
  assign n59928 = pi5784 & ~pi9040;
  assign n59929 = pi5696 & pi9040;
  assign n59930 = ~n59928 & ~n59929;
  assign n59931 = ~pi1664 & n59930;
  assign n59932 = pi1664 & ~n59930;
  assign n59933 = ~n59931 & ~n59932;
  assign n59934 = ~n59925 & ~n59933;
  assign n59935 = n59919 & n59934;
  assign n59936 = ~n59927 & ~n59935;
  assign n59937 = ~n59913 & ~n59919;
  assign n59938 = n59933 & n59937;
  assign n59939 = ~n59925 & n59938;
  assign n59940 = n59936 & ~n59939;
  assign n59941 = n59907 & ~n59940;
  assign n59942 = ~n59919 & ~n59925;
  assign n59943 = ~n59933 & n59942;
  assign n59944 = ~n59913 & n59943;
  assign n59945 = n59925 & ~n59933;
  assign n59946 = n59919 & n59945;
  assign n59947 = ~n59913 & n59946;
  assign n59948 = ~n59925 & n59933;
  assign n59949 = ~n59919 & n59925;
  assign n59950 = ~n59948 & ~n59949;
  assign n59951 = n59913 & ~n59950;
  assign n59952 = ~n59947 & ~n59951;
  assign n59953 = ~n59944 & n59952;
  assign n59954 = ~n59907 & ~n59953;
  assign n59955 = ~n59941 & ~n59954;
  assign n59956 = n59901 & ~n59955;
  assign n59957 = n59907 & ~n59913;
  assign n59958 = n59925 & n59957;
  assign n59959 = ~n59907 & ~n59913;
  assign n59960 = n59948 & n59959;
  assign n59961 = ~n59913 & ~n59925;
  assign n59962 = n59919 & n59961;
  assign n59963 = ~n59927 & ~n59962;
  assign n59964 = ~n59907 & ~n59963;
  assign n59965 = ~n59960 & ~n59964;
  assign n59966 = n59919 & n59948;
  assign n59967 = ~n59913 & n59966;
  assign n59968 = n59913 & n59943;
  assign n59969 = ~n59967 & ~n59968;
  assign n59970 = n59907 & n59913;
  assign n59971 = n59942 & n59970;
  assign n59972 = ~n59919 & n59945;
  assign n59973 = n59907 & n59972;
  assign n59974 = ~n59971 & ~n59973;
  assign n59975 = n59969 & n59974;
  assign n59976 = n59965 & n59975;
  assign n59977 = ~n59958 & n59976;
  assign n59978 = ~n59901 & ~n59977;
  assign n59979 = n59925 & n59933;
  assign n59980 = ~n59919 & n59979;
  assign n59981 = ~n59907 & n59980;
  assign n59982 = ~n59913 & n59981;
  assign n59983 = ~n59907 & n59967;
  assign n59984 = ~n59982 & ~n59983;
  assign n59985 = ~n59933 & n59937;
  assign n59986 = n59925 & n59985;
  assign n59987 = n59907 & n59986;
  assign n59988 = n59984 & ~n59987;
  assign n59989 = ~n59913 & n59919;
  assign n59990 = n59933 & n59989;
  assign n59991 = n59925 & n59990;
  assign n59992 = n59913 & n59934;
  assign n59993 = ~n59991 & ~n59992;
  assign n59994 = n59907 & ~n59993;
  assign n59995 = n59988 & ~n59994;
  assign n59996 = ~n59978 & n59995;
  assign n59997 = ~n59956 & n59996;
  assign n59998 = ~pi1710 & ~n59997;
  assign n59999 = pi1710 & n59997;
  assign po1790 = n59998 | n59999;
  assign n60001 = n59801 & ~n59807;
  assign n60002 = ~n59844 & ~n60001;
  assign n60003 = ~n59875 & n60002;
  assign n60004 = n59826 & ~n60003;
  assign n60005 = ~n59820 & ~n59826;
  assign n60006 = n59807 & n60005;
  assign n60007 = n59801 & ~n59820;
  assign n60008 = ~n59813 & n60007;
  assign n60009 = n59820 & n59837;
  assign n60010 = ~n60008 & ~n60009;
  assign n60011 = ~n59801 & ~n59807;
  assign n60012 = n59820 & ~n59826;
  assign n60013 = n60011 & n60012;
  assign n60014 = n60010 & ~n60013;
  assign n60015 = ~n60006 & n60014;
  assign n60016 = ~n60004 & n60015;
  assign n60017 = n59795 & ~n60016;
  assign n60018 = n59801 & n59814;
  assign n60019 = n59820 & n60018;
  assign n60020 = n59813 & n60001;
  assign n60021 = ~n59820 & n60020;
  assign n60022 = ~n60019 & ~n60021;
  assign n60023 = n59826 & ~n60022;
  assign n60024 = ~n60017 & ~n60023;
  assign n60025 = ~n59820 & n59837;
  assign n60026 = ~n59848 & ~n59859;
  assign n60027 = n59826 & ~n60026;
  assign n60028 = ~n60025 & ~n60027;
  assign n60029 = ~n59863 & n60028;
  assign n60030 = ~n59795 & ~n60029;
  assign n60031 = ~n59831 & ~n59852;
  assign n60032 = ~n59801 & ~n60031;
  assign n60033 = ~n59853 & ~n60032;
  assign n60034 = ~n59826 & ~n60033;
  assign n60035 = ~n59795 & n60034;
  assign n60036 = ~n60030 & ~n60035;
  assign n60037 = n60024 & n60036;
  assign n60038 = pi1715 & ~n60037;
  assign n60039 = ~pi1715 & n60024;
  assign n60040 = n60036 & n60039;
  assign po1791 = n60038 | n60040;
  assign n60042 = ~n59705 & n59724;
  assign n60043 = ~n59749 & ~n59763;
  assign n60044 = n60042 & ~n60043;
  assign n60045 = ~n59705 & ~n59730;
  assign n60046 = n59749 & n60045;
  assign n60047 = ~n60044 & ~n60046;
  assign n60048 = n59742 & ~n60047;
  assign n60049 = ~n59724 & n59747;
  assign n60050 = ~n59724 & n59730;
  assign n60051 = ~n59780 & ~n60050;
  assign n60052 = n59705 & ~n60051;
  assign n60053 = ~n59724 & ~n59730;
  assign n60054 = ~n59717 & n60053;
  assign n60055 = n59711 & n60054;
  assign n60056 = ~n60052 & ~n60055;
  assign n60057 = ~n60049 & n60056;
  assign n60058 = n59742 & ~n60057;
  assign n60059 = ~n60048 & ~n60058;
  assign n60060 = n59717 & n59731;
  assign n60061 = ~n59711 & n60060;
  assign n60062 = ~n59724 & n59756;
  assign n60063 = ~n60061 & ~n60062;
  assign n60064 = ~n59705 & ~n60063;
  assign n60065 = ~n59718 & ~n59780;
  assign n60066 = n59724 & ~n60065;
  assign n60067 = ~n59756 & ~n60066;
  assign n60068 = ~n59705 & ~n60067;
  assign n60069 = n59717 & ~n59724;
  assign n60070 = n60045 & n60069;
  assign n60071 = ~n59717 & n59730;
  assign n60072 = ~n59756 & ~n60071;
  assign n60073 = ~n59724 & ~n60072;
  assign n60074 = n59705 & n59724;
  assign n60075 = n59746 & n60074;
  assign n60076 = ~n59730 & n60075;
  assign n60077 = ~n60073 & ~n60076;
  assign n60078 = ~n60070 & n60077;
  assign n60079 = ~n60068 & n60078;
  assign n60080 = ~n60061 & n60079;
  assign n60081 = ~n59742 & ~n60080;
  assign n60082 = n59724 & n59771;
  assign n60083 = ~n59724 & n59780;
  assign n60084 = ~n60082 & ~n60083;
  assign n60085 = n59705 & ~n60084;
  assign n60086 = ~n60081 & ~n60085;
  assign n60087 = ~n60064 & n60086;
  assign n60088 = n60059 & n60087;
  assign n60089 = pi1716 & n60088;
  assign n60090 = ~pi1716 & ~n60088;
  assign po1793 = n60089 | n60090;
  assign n60092 = ~n59901 & ~n59907;
  assign n60093 = ~n59913 & n59926;
  assign n60094 = n59913 & n59966;
  assign n60095 = ~n59913 & n59934;
  assign n60096 = ~n60094 & ~n60095;
  assign n60097 = ~n60093 & n60096;
  assign n60098 = n60092 & ~n60097;
  assign n60099 = n59919 & n59979;
  assign n60100 = n59913 & n60099;
  assign n60101 = ~n59938 & ~n60100;
  assign n60102 = ~n59919 & n59948;
  assign n60103 = ~n59935 & ~n60102;
  assign n60104 = n60101 & n60103;
  assign n60105 = n59907 & ~n60104;
  assign n60106 = n59913 & n59972;
  assign n60107 = ~n60105 & ~n60106;
  assign n60108 = ~n59901 & ~n60107;
  assign n60109 = ~n60098 & ~n60108;
  assign n60110 = n59919 & n59957;
  assign n60111 = ~n59933 & n60110;
  assign n60112 = ~n59939 & ~n60111;
  assign n60113 = ~n59934 & ~n59979;
  assign n60114 = n59913 & ~n60113;
  assign n60115 = ~n59980 & ~n60114;
  assign n60116 = ~n59907 & ~n60115;
  assign n60117 = ~n59946 & ~n60093;
  assign n60118 = ~n60094 & n60117;
  assign n60119 = n59907 & ~n60118;
  assign n60120 = ~n60116 & ~n60119;
  assign n60121 = n59913 & n59980;
  assign n60122 = ~n59968 & ~n60121;
  assign n60123 = ~n59986 & n60122;
  assign n60124 = ~n59960 & n60123;
  assign n60125 = n60120 & n60124;
  assign n60126 = n59901 & ~n60125;
  assign n60127 = n60112 & ~n60126;
  assign n60128 = n60109 & n60127;
  assign n60129 = pi1701 & ~n60128;
  assign n60130 = ~pi1701 & n60112;
  assign n60131 = n60109 & n60130;
  assign n60132 = ~n60126 & n60131;
  assign po1794 = n60129 | n60132;
  assign n60134 = ~n59732 & ~n60049;
  assign n60135 = ~n59705 & ~n60134;
  assign n60136 = ~n59750 & ~n59757;
  assign n60137 = ~n60055 & n60136;
  assign n60138 = n59777 & ~n60137;
  assign n60139 = n59718 & n60050;
  assign n60140 = n59772 & ~n60139;
  assign n60141 = n59705 & ~n60140;
  assign n60142 = ~n59724 & n59760;
  assign n60143 = ~n60141 & ~n60142;
  assign n60144 = n59711 & n59733;
  assign n60145 = n59724 & n59746;
  assign n60146 = ~n60144 & ~n60145;
  assign n60147 = n59705 & ~n60146;
  assign n60148 = n59705 & n59755;
  assign n60149 = ~n59724 & n60148;
  assign n60150 = ~n60147 & ~n60149;
  assign n60151 = n60143 & n60150;
  assign n60152 = ~n59742 & ~n60151;
  assign n60153 = ~n60138 & ~n60152;
  assign n60154 = ~n59717 & n59733;
  assign n60155 = ~n59763 & ~n60154;
  assign n60156 = ~n59705 & ~n60155;
  assign n60157 = n59724 & n59755;
  assign n60158 = ~n60054 & ~n60157;
  assign n60159 = n59705 & ~n60158;
  assign n60160 = ~n59724 & n59750;
  assign n60161 = ~n60070 & ~n60160;
  assign n60162 = ~n59732 & n60161;
  assign n60163 = ~n60159 & n60162;
  assign n60164 = ~n60156 & n60163;
  assign n60165 = ~n60049 & ~n60061;
  assign n60166 = n60164 & n60165;
  assign n60167 = n59742 & ~n60166;
  assign n60168 = n60153 & ~n60167;
  assign n60169 = ~n60135 & n60168;
  assign n60170 = ~pi1722 & n60169;
  assign n60171 = pi1722 & ~n60169;
  assign po1795 = n60170 | n60171;
  assign n60173 = ~n59405 & ~n59434;
  assign n60174 = n59411 & n60173;
  assign n60175 = n59417 & n59444;
  assign n60176 = n59405 & n60175;
  assign n60177 = n59405 & n59455;
  assign n60178 = ~n60176 & ~n60177;
  assign n60179 = ~n59405 & ~n59417;
  assign n60180 = ~n59423 & n60179;
  assign n60181 = ~n59411 & n60180;
  assign n60182 = ~n59437 & ~n60181;
  assign n60183 = n59434 & ~n60182;
  assign n60184 = n60178 & ~n60183;
  assign n60185 = ~n60174 & n60184;
  assign n60186 = n59399 & ~n60185;
  assign n60187 = n59405 & n59476;
  assign n60188 = ~n59434 & n60187;
  assign n60189 = n59467 & n59476;
  assign n60190 = ~n59435 & ~n60189;
  assign n60191 = ~n59437 & ~n59470;
  assign n60192 = ~n59405 & n59454;
  assign n60193 = n60191 & ~n60192;
  assign n60194 = ~n59434 & ~n60193;
  assign n60195 = n59434 & n59441;
  assign n60196 = ~n60194 & ~n60195;
  assign n60197 = n59459 & n60196;
  assign n60198 = n60190 & n60197;
  assign n60199 = ~n59399 & ~n60198;
  assign n60200 = ~n60188 & ~n60199;
  assign n60201 = ~n60186 & n60200;
  assign n60202 = n59467 & n59470;
  assign n60203 = n59424 & n59434;
  assign n60204 = n59405 & n60203;
  assign n60205 = ~n60202 & ~n60204;
  assign n60206 = n59434 & n60177;
  assign n60207 = n60205 & ~n60206;
  assign n60208 = n60201 & n60207;
  assign n60209 = ~pi1707 & ~n60208;
  assign n60210 = pi1707 & n60207;
  assign n60211 = n60200 & n60210;
  assign n60212 = ~n60186 & n60211;
  assign po1796 = n60209 | n60212;
  assign n60214 = pi5561 & ~pi9040;
  assign n60215 = pi5830 & pi9040;
  assign n60216 = ~n60214 & ~n60215;
  assign n60217 = pi1679 & n60216;
  assign n60218 = ~pi1679 & ~n60216;
  assign n60219 = ~n60217 & ~n60218;
  assign n60220 = pi5581 & ~pi9040;
  assign n60221 = pi5559 & pi9040;
  assign n60222 = ~n60220 & ~n60221;
  assign n60223 = ~pi1675 & n60222;
  assign n60224 = pi1675 & ~n60222;
  assign n60225 = ~n60223 & ~n60224;
  assign n60226 = pi5553 & ~pi9040;
  assign n60227 = pi5580 & pi9040;
  assign n60228 = ~n60226 & ~n60227;
  assign n60229 = ~pi1672 & n60228;
  assign n60230 = pi1672 & ~n60228;
  assign n60231 = ~n60229 & ~n60230;
  assign n60232 = pi5556 & pi9040;
  assign n60233 = pi5779 & ~pi9040;
  assign n60234 = ~n60232 & ~n60233;
  assign n60235 = ~pi1662 & n60234;
  assign n60236 = pi1662 & ~n60234;
  assign n60237 = ~n60235 & ~n60236;
  assign n60238 = pi5560 & ~pi9040;
  assign n60239 = pi5834 & pi9040;
  assign n60240 = ~n60238 & ~n60239;
  assign n60241 = ~pi1678 & ~n60240;
  assign n60242 = pi1678 & n60240;
  assign n60243 = ~n60241 & ~n60242;
  assign n60244 = n60237 & n60243;
  assign n60245 = ~n60231 & n60244;
  assign n60246 = ~n60225 & n60245;
  assign n60247 = ~n60219 & n60246;
  assign n60248 = ~n60219 & n60231;
  assign n60249 = ~n60243 & n60248;
  assign n60250 = ~n60237 & n60249;
  assign n60251 = ~n60225 & n60250;
  assign n60252 = ~n60247 & ~n60251;
  assign n60253 = n60231 & n60244;
  assign n60254 = ~n60219 & n60225;
  assign n60255 = n60253 & n60254;
  assign n60256 = ~n60250 & ~n60255;
  assign n60257 = ~n60231 & ~n60237;
  assign n60258 = n60219 & n60257;
  assign n60259 = n60219 & n60244;
  assign n60260 = ~n60258 & ~n60259;
  assign n60261 = ~n60225 & ~n60260;
  assign n60262 = ~n60237 & n60243;
  assign n60263 = n60237 & ~n60243;
  assign n60264 = ~n60262 & ~n60263;
  assign n60265 = n60225 & ~n60248;
  assign n60266 = ~n60264 & n60265;
  assign n60267 = ~n60219 & ~n60225;
  assign n60268 = ~n60244 & n60267;
  assign n60269 = n60231 & n60268;
  assign n60270 = ~n60266 & ~n60269;
  assign n60271 = ~n60261 & n60270;
  assign n60272 = n60256 & n60271;
  assign n60273 = pi5675 & pi9040;
  assign n60274 = pi5663 & ~pi9040;
  assign n60275 = ~n60273 & ~n60274;
  assign n60276 = pi1677 & n60275;
  assign n60277 = ~pi1677 & ~n60275;
  assign n60278 = ~n60276 & ~n60277;
  assign n60279 = ~n60272 & n60278;
  assign n60280 = n60252 & ~n60279;
  assign n60281 = ~n60231 & n60262;
  assign n60282 = n60225 & n60281;
  assign n60283 = n60219 & n60282;
  assign n60284 = n60225 & ~n60278;
  assign n60285 = ~n60237 & ~n60243;
  assign n60286 = ~n60231 & n60285;
  assign n60287 = ~n60259 & ~n60286;
  assign n60288 = n60248 & ~n60264;
  assign n60289 = n60287 & ~n60288;
  assign n60290 = n60284 & ~n60289;
  assign n60291 = ~n60283 & ~n60290;
  assign n60292 = n60231 & n60285;
  assign n60293 = n60219 & n60292;
  assign n60294 = n60219 & ~n60237;
  assign n60295 = n60231 & n60294;
  assign n60296 = n60219 & n60263;
  assign n60297 = ~n60295 & ~n60296;
  assign n60298 = ~n60219 & n60244;
  assign n60299 = ~n60231 & n60263;
  assign n60300 = ~n60298 & ~n60299;
  assign n60301 = n60297 & n60300;
  assign n60302 = ~n60225 & ~n60301;
  assign n60303 = ~n60293 & ~n60302;
  assign n60304 = ~n60278 & ~n60303;
  assign n60305 = n60291 & ~n60304;
  assign n60306 = n60280 & n60305;
  assign n60307 = pi1727 & ~n60306;
  assign n60308 = ~pi1727 & n60280;
  assign n60309 = n60305 & n60308;
  assign po1797 = n60307 | n60309;
  assign n60311 = n59606 & n59645;
  assign n60312 = ~n59624 & n59660;
  assign n60313 = ~n59636 & n60312;
  assign n60314 = ~n60311 & ~n60313;
  assign n60315 = n59633 & ~n60314;
  assign n60316 = ~n59633 & n59667;
  assign n60317 = ~n59667 & ~n59674;
  assign n60318 = ~n59606 & ~n59612;
  assign n60319 = n59624 & n60318;
  assign n60320 = ~n59636 & n60319;
  assign n60321 = ~n59606 & ~n59633;
  assign n60322 = n59644 & n60321;
  assign n60323 = n59612 & n60322;
  assign n60324 = ~n59618 & n59665;
  assign n60325 = ~n59669 & ~n60324;
  assign n60326 = ~n59633 & ~n60325;
  assign n60327 = n59612 & n59633;
  assign n60328 = n59624 & n60327;
  assign n60329 = ~n59618 & n60328;
  assign n60330 = ~n60326 & ~n60329;
  assign n60331 = ~n60323 & n60330;
  assign n60332 = ~n60320 & n60331;
  assign n60333 = n60317 & n60332;
  assign n60334 = n59600 & ~n60333;
  assign n60335 = n59606 & n59674;
  assign n60336 = ~n60334 & ~n60335;
  assign n60337 = ~n60316 & n60336;
  assign n60338 = ~n60315 & n60337;
  assign n60339 = ~n59612 & ~n59618;
  assign n60340 = n59671 & n60339;
  assign n60341 = ~n59646 & ~n60340;
  assign n60342 = n59633 & n59681;
  assign n60343 = n59606 & n59691;
  assign n60344 = ~n60342 & ~n60343;
  assign n60345 = ~n59606 & n59654;
  assign n60346 = ~n60311 & ~n60345;
  assign n60347 = ~n59606 & n59651;
  assign n60348 = n59612 & n59624;
  assign n60349 = ~n60347 & ~n60348;
  assign n60350 = ~n59633 & ~n60349;
  assign n60351 = n60346 & ~n60350;
  assign n60352 = n60344 & n60351;
  assign n60353 = n60341 & n60352;
  assign n60354 = ~n59600 & ~n60353;
  assign n60355 = n60338 & ~n60354;
  assign n60356 = ~pi1711 & ~n60355;
  assign n60357 = pi1711 & n60338;
  assign n60358 = ~n60354 & n60357;
  assign po1798 = n60356 | n60358;
  assign n60360 = n59606 & n59647;
  assign n60361 = n59618 & n59660;
  assign n60362 = ~n59678 & ~n60361;
  assign n60363 = n59633 & ~n60362;
  assign n60364 = ~n60360 & ~n60363;
  assign n60365 = ~n59633 & n59637;
  assign n60366 = n59606 & n60365;
  assign n60367 = ~n59633 & n59645;
  assign n60368 = ~n60366 & ~n60367;
  assign n60369 = n60364 & n60368;
  assign n60370 = n59618 & n59665;
  assign n60371 = ~n60311 & ~n60370;
  assign n60372 = ~n60345 & n60371;
  assign n60373 = n60369 & n60372;
  assign n60374 = ~n59600 & ~n60373;
  assign n60375 = ~n59667 & ~n59678;
  assign n60376 = ~n60347 & n60375;
  assign n60377 = ~n59633 & ~n60376;
  assign n60378 = ~n59606 & n59639;
  assign n60379 = ~n60320 & ~n60378;
  assign n60380 = ~n59693 & n60379;
  assign n60381 = n59633 & n59654;
  assign n60382 = n60380 & ~n60381;
  assign n60383 = ~n60377 & n60382;
  assign n60384 = n59600 & ~n60383;
  assign n60385 = ~n60335 & ~n60340;
  assign n60386 = ~n60311 & n60379;
  assign n60387 = ~n59633 & ~n60386;
  assign n60388 = n60385 & ~n60387;
  assign n60389 = ~n60384 & n60388;
  assign n60390 = ~n60374 & n60389;
  assign n60391 = pi1721 & ~n60390;
  assign n60392 = ~pi1721 & n60390;
  assign po1799 = n60391 | n60392;
  assign n60394 = n59518 & n59546;
  assign n60395 = ~n59565 & ~n59574;
  assign n60396 = n59524 & ~n60395;
  assign n60397 = ~n60394 & ~n60396;
  assign n60398 = ~n59560 & n60397;
  assign n60399 = ~n59524 & n59563;
  assign n60400 = ~n59552 & ~n60399;
  assign n60401 = ~n59581 & n60400;
  assign n60402 = n60398 & n60401;
  assign n60403 = n59499 & ~n60402;
  assign n60404 = n59532 & n59539;
  assign n60405 = n59518 & n60404;
  assign n60406 = ~n59537 & ~n60405;
  assign n60407 = ~n59518 & n59580;
  assign n60408 = ~n59547 & ~n60407;
  assign n60409 = n59512 & n59532;
  assign n60410 = n59524 & n60409;
  assign n60411 = n59518 & n59551;
  assign n60412 = ~n60410 & ~n60411;
  assign n60413 = n59511 & ~n59532;
  assign n60414 = ~n59505 & n59518;
  assign n60415 = ~n60413 & ~n60414;
  assign n60416 = ~n59586 & n60415;
  assign n60417 = ~n59524 & ~n60416;
  assign n60418 = n60412 & ~n60417;
  assign n60419 = n60408 & n60418;
  assign n60420 = n60406 & n60419;
  assign n60421 = ~n59499 & ~n60420;
  assign n60422 = ~n60403 & ~n60421;
  assign n60423 = pi1698 & ~n60422;
  assign n60424 = ~pi1698 & ~n60403;
  assign n60425 = ~n60421 & n60424;
  assign po1800 = n60423 | n60425;
  assign n60427 = ~n59405 & n60175;
  assign n60428 = ~n59455 & ~n59463;
  assign n60429 = n59405 & n59424;
  assign n60430 = ~n59405 & n59476;
  assign n60431 = ~n60429 & ~n60430;
  assign n60432 = n60428 & n60431;
  assign n60433 = ~n59434 & ~n60432;
  assign n60434 = n59405 & n59436;
  assign n60435 = ~n59435 & ~n60434;
  assign n60436 = ~n59457 & n60435;
  assign n60437 = n59434 & ~n60436;
  assign n60438 = n59405 & n59437;
  assign n60439 = ~n60437 & ~n60438;
  assign n60440 = ~n60433 & n60439;
  assign n60441 = ~n60427 & n60440;
  assign n60442 = ~n59399 & ~n60441;
  assign n60443 = n59405 & n59441;
  assign n60444 = ~n59434 & n60443;
  assign n60445 = ~n59434 & n59457;
  assign n60446 = ~n59434 & n59470;
  assign n60447 = ~n60445 & ~n60446;
  assign n60448 = ~n59405 & ~n60447;
  assign n60449 = ~n60444 & ~n60448;
  assign n60450 = n59405 & n59454;
  assign n60451 = ~n59405 & n59436;
  assign n60452 = ~n60450 & ~n60451;
  assign n60453 = ~n59425 & n60452;
  assign n60454 = ~n59455 & n60453;
  assign n60455 = n59434 & ~n60454;
  assign n60456 = ~n59405 & n59437;
  assign n60457 = ~n60455 & ~n60456;
  assign n60458 = ~n59405 & n59425;
  assign n60459 = ~n60187 & ~n60458;
  assign n60460 = n60457 & n60459;
  assign n60461 = n60449 & n60460;
  assign n60462 = n59399 & ~n60461;
  assign n60463 = ~n59434 & ~n60178;
  assign n60464 = ~n60462 & ~n60463;
  assign n60465 = ~n59458 & ~n60458;
  assign n60466 = n59434 & ~n60465;
  assign n60467 = n60464 & ~n60466;
  assign n60468 = ~n60442 & n60467;
  assign n60469 = pi1714 & ~n60468;
  assign n60470 = ~pi1714 & n60468;
  assign po1801 = n60469 | n60470;
  assign n60472 = ~n60281 & ~n60292;
  assign n60473 = ~n60219 & ~n60231;
  assign n60474 = n60243 & n60473;
  assign n60475 = n60472 & ~n60474;
  assign n60476 = n60225 & n60278;
  assign n60477 = ~n60475 & n60476;
  assign n60478 = n60219 & n60278;
  assign n60479 = n60299 & n60478;
  assign n60480 = ~n60225 & n60286;
  assign n60481 = n60231 & n60243;
  assign n60482 = ~n60259 & ~n60481;
  assign n60483 = ~n60225 & ~n60482;
  assign n60484 = ~n60480 & ~n60483;
  assign n60485 = n60278 & ~n60484;
  assign n60486 = ~n60479 & ~n60485;
  assign n60487 = n60237 & n60249;
  assign n60488 = n60219 & n60231;
  assign n60489 = n60243 & n60488;
  assign n60490 = ~n60487 & ~n60489;
  assign n60491 = ~n60225 & ~n60490;
  assign n60492 = n60486 & ~n60491;
  assign n60493 = n60219 & n60225;
  assign n60494 = n60244 & n60493;
  assign n60495 = ~n60231 & n60494;
  assign n60496 = ~n60264 & n60473;
  assign n60497 = ~n60250 & ~n60496;
  assign n60498 = ~n60264 & n60488;
  assign n60499 = n60219 & ~n60231;
  assign n60500 = ~n60243 & n60499;
  assign n60501 = ~n60237 & n60500;
  assign n60502 = ~n60498 & ~n60501;
  assign n60503 = ~n60255 & n60502;
  assign n60504 = n60497 & n60503;
  assign n60505 = ~n60495 & n60504;
  assign n60506 = ~n60231 & n60267;
  assign n60507 = n60237 & n60506;
  assign n60508 = n60505 & ~n60507;
  assign n60509 = ~n60278 & ~n60508;
  assign n60510 = n60492 & ~n60509;
  assign n60511 = ~n60477 & n60510;
  assign n60512 = ~pi1726 & ~n60511;
  assign n60513 = pi1726 & n60492;
  assign n60514 = ~n60477 & n60513;
  assign n60515 = ~n60509 & n60514;
  assign po1802 = n60512 | n60515;
  assign n60517 = ~n60296 & ~n60298;
  assign n60518 = ~n60225 & ~n60517;
  assign n60519 = ~n60251 & ~n60518;
  assign n60520 = n60278 & ~n60519;
  assign n60521 = n60231 & ~n60237;
  assign n60522 = ~n60262 & ~n60521;
  assign n60523 = ~n60219 & ~n60522;
  assign n60524 = ~n60245 & ~n60523;
  assign n60525 = n60225 & ~n60524;
  assign n60526 = ~n60288 & ~n60525;
  assign n60527 = n60219 & n60253;
  assign n60528 = ~n60243 & n60473;
  assign n60529 = n60219 & ~n60522;
  assign n60530 = ~n60528 & ~n60529;
  assign n60531 = ~n60225 & ~n60530;
  assign n60532 = ~n60527 & ~n60531;
  assign n60533 = n60526 & n60532;
  assign n60534 = ~n60278 & ~n60533;
  assign n60535 = ~n60262 & n60499;
  assign n60536 = n60278 & n60535;
  assign n60537 = n60262 & n60488;
  assign n60538 = ~n60225 & n60537;
  assign n60539 = ~n60231 & ~n60243;
  assign n60540 = n60493 & n60539;
  assign n60541 = ~n60538 & ~n60540;
  assign n60542 = ~n60536 & n60541;
  assign n60543 = ~n60294 & ~n60299;
  assign n60544 = n60476 & ~n60543;
  assign n60545 = n60542 & ~n60544;
  assign n60546 = ~n60534 & n60545;
  assign n60547 = ~n60520 & n60546;
  assign n60548 = pi1729 & ~n60547;
  assign n60549 = ~pi1729 & n60547;
  assign po1803 = n60548 | n60549;
  assign n60551 = ~n59820 & n60032;
  assign n60552 = ~n59847 & ~n60018;
  assign n60553 = ~n59826 & ~n60552;
  assign n60554 = ~n60551 & ~n60553;
  assign n60555 = n59813 & n60007;
  assign n60556 = ~n59884 & ~n60555;
  assign n60557 = ~n60020 & n60556;
  assign n60558 = n59826 & ~n60557;
  assign n60559 = n60554 & ~n60558;
  assign n60560 = n59820 & n59859;
  assign n60561 = n60559 & ~n60560;
  assign n60562 = ~n59795 & ~n60561;
  assign n60563 = n59830 & ~n60552;
  assign n60564 = ~n59848 & ~n59862;
  assign n60565 = ~n59859 & ~n60020;
  assign n60566 = n60564 & n60565;
  assign n60567 = ~n59820 & ~n60566;
  assign n60568 = ~n60563 & ~n60567;
  assign n60569 = ~n60009 & n60568;
  assign n60570 = n59795 & ~n60569;
  assign n60571 = ~n60562 & ~n60570;
  assign n60572 = ~n59820 & n60018;
  assign n60573 = ~n60560 & ~n60572;
  assign n60574 = ~n59826 & ~n60573;
  assign n60575 = n60571 & ~n60574;
  assign n60576 = pi1719 & ~n60575;
  assign n60577 = ~pi1719 & ~n60574;
  assign n60578 = ~n60570 & n60577;
  assign n60579 = ~n60562 & n60578;
  assign po1804 = n60576 | n60579;
  assign n60581 = ~n59653 & ~n59661;
  assign n60582 = n59600 & ~n60581;
  assign n60583 = ~n59666 & ~n60324;
  assign n60584 = ~n59626 & n60583;
  assign n60585 = ~n59633 & ~n60584;
  assign n60586 = n59600 & n60585;
  assign n60587 = ~n60582 & ~n60586;
  assign n60588 = n59652 & n60321;
  assign n60589 = ~n60323 & ~n60588;
  assign n60590 = ~n59669 & ~n60348;
  assign n60591 = n59633 & ~n60590;
  assign n60592 = n59600 & n60591;
  assign n60593 = n60589 & ~n60592;
  assign n60594 = n59606 & n59652;
  assign n60595 = n59606 & n59644;
  assign n60596 = ~n60313 & ~n60595;
  assign n60597 = n59633 & ~n60596;
  assign n60598 = ~n59667 & ~n60320;
  assign n60599 = n59606 & n59651;
  assign n60600 = ~n59691 & ~n60599;
  assign n60601 = ~n59633 & ~n60600;
  assign n60602 = n60598 & ~n60601;
  assign n60603 = ~n60597 & n60602;
  assign n60604 = ~n60594 & n60603;
  assign n60605 = ~n59600 & ~n60604;
  assign n60606 = ~n60345 & n60379;
  assign n60607 = n59633 & ~n60606;
  assign n60608 = ~n60605 & ~n60607;
  assign n60609 = n60593 & n60608;
  assign n60610 = n60587 & n60609;
  assign n60611 = ~pi1730 & ~n60610;
  assign n60612 = pi1730 & n60593;
  assign n60613 = n60587 & n60612;
  assign n60614 = n60608 & n60613;
  assign po1806 = n60611 | n60614;
  assign n60616 = ~n59324 & n59354;
  assign n60617 = n59324 & n59365;
  assign n60618 = ~n59351 & ~n60617;
  assign n60619 = n59298 & ~n60618;
  assign n60620 = ~n60616 & ~n60619;
  assign n60621 = ~n59298 & ~n59324;
  assign n60622 = ~n59316 & n60621;
  assign n60623 = ~n59310 & n60622;
  assign n60624 = n59332 & n59366;
  assign n60625 = ~n60623 & ~n60624;
  assign n60626 = ~n59298 & ~n59304;
  assign n60627 = n59326 & n60626;
  assign n60628 = n60625 & ~n60627;
  assign n60629 = ~n59328 & ~n59340;
  assign n60630 = n59316 & n59330;
  assign n60631 = n60629 & ~n60630;
  assign n60632 = n60628 & n60631;
  assign n60633 = n60620 & n60632;
  assign n60634 = ~n59363 & ~n60633;
  assign n60635 = ~n59327 & ~n59351;
  assign n60636 = n59324 & ~n60635;
  assign n60637 = ~n59324 & n59350;
  assign n60638 = ~n59310 & n59339;
  assign n60639 = ~n60637 & ~n60638;
  assign n60640 = ~n59298 & ~n60639;
  assign n60641 = ~n59310 & n59369;
  assign n60642 = ~n59380 & ~n60641;
  assign n60643 = ~n59304 & ~n59316;
  assign n60644 = n59324 & n60643;
  assign n60645 = n60642 & ~n60644;
  assign n60646 = n59298 & ~n60645;
  assign n60647 = ~n59324 & n59333;
  assign n60648 = ~n60646 & ~n60647;
  assign n60649 = ~n60640 & n60648;
  assign n60650 = ~n60636 & n60649;
  assign n60651 = n59363 & ~n60650;
  assign n60652 = n59298 & n59370;
  assign n60653 = ~n60651 & ~n60652;
  assign n60654 = n59345 & n60621;
  assign n60655 = ~n59316 & n60654;
  assign n60656 = n60653 & ~n60655;
  assign n60657 = ~n60634 & n60656;
  assign n60658 = ~pi1699 & ~n60657;
  assign n60659 = pi1699 & n60653;
  assign n60660 = ~n60634 & n60659;
  assign n60661 = ~n60655 & n60660;
  assign po1807 = n60658 | n60661;
  assign n60663 = n59907 & n59934;
  assign n60664 = ~n59913 & n60663;
  assign n60665 = ~n59991 & ~n60664;
  assign n60666 = n59913 & ~n59933;
  assign n60667 = n59919 & n60666;
  assign n60668 = ~n59913 & n59925;
  assign n60669 = ~n59990 & ~n60668;
  assign n60670 = ~n59907 & ~n60669;
  assign n60671 = ~n60667 & ~n60670;
  assign n60672 = n60665 & n60671;
  assign n60673 = n59901 & ~n60672;
  assign n60674 = ~n59966 & ~n59968;
  assign n60675 = ~n59913 & n59945;
  assign n60676 = n60674 & ~n60675;
  assign n60677 = n59907 & ~n60676;
  assign n60678 = n59934 & n59959;
  assign n60679 = ~n59939 & ~n60678;
  assign n60680 = ~n60677 & n60679;
  assign n60681 = ~n60099 & ~n60106;
  assign n60682 = ~n59907 & ~n60681;
  assign n60683 = n60680 & ~n60682;
  assign n60684 = ~n59901 & ~n60683;
  assign n60685 = ~n60673 & ~n60684;
  assign n60686 = ~n59913 & n59979;
  assign n60687 = n59913 & ~n60103;
  assign n60688 = ~n60686 & ~n60687;
  assign n60689 = ~n59907 & ~n60688;
  assign n60690 = ~n59946 & ~n59980;
  assign n60691 = ~n59966 & n60690;
  assign n60692 = n59970 & ~n60691;
  assign n60693 = ~n60689 & ~n60692;
  assign n60694 = n60685 & n60693;
  assign n60695 = ~pi1717 & ~n60694;
  assign n60696 = ~n60684 & n60693;
  assign n60697 = pi1717 & n60696;
  assign n60698 = ~n60673 & n60697;
  assign po1808 = n60695 | n60698;
  assign n60700 = ~n59907 & ~n60690;
  assign n60701 = n59913 & n59935;
  assign n60702 = ~n60700 & ~n60701;
  assign n60703 = n59913 & ~n59925;
  assign n60704 = ~n59942 & ~n60703;
  assign n60705 = ~n60099 & n60704;
  assign n60706 = n59907 & ~n60705;
  assign n60707 = n60702 & ~n60706;
  assign n60708 = ~n59901 & ~n60707;
  assign n60709 = ~n59907 & n59944;
  assign n60710 = ~n59983 & ~n60709;
  assign n60711 = ~n59987 & n60710;
  assign n60712 = ~n59986 & ~n59990;
  assign n60713 = n59907 & n59962;
  assign n60714 = n59913 & n59946;
  assign n60715 = ~n59907 & n59942;
  assign n60716 = ~n60714 & ~n60715;
  assign n60717 = ~n60121 & n60716;
  assign n60718 = ~n60713 & n60717;
  assign n60719 = n60712 & n60718;
  assign n60720 = ~n59973 & n60719;
  assign n60721 = n59901 & ~n60720;
  assign n60722 = n60711 & ~n60721;
  assign n60723 = ~n60708 & n60722;
  assign n60724 = ~pi1704 & ~n60723;
  assign n60725 = pi1704 & n60711;
  assign n60726 = ~n60708 & n60725;
  assign n60727 = ~n60721 & n60726;
  assign po1809 = n60724 | n60727;
  assign n60729 = n59820 & n59862;
  assign n60730 = ~n60009 & ~n60729;
  assign n60731 = ~n59826 & ~n60730;
  assign n60732 = n59859 & n60005;
  assign n60733 = ~n60731 & ~n60732;
  assign n60734 = ~n59872 & n60733;
  assign n60735 = n59801 & n59826;
  assign n60736 = n59813 & n60735;
  assign n60737 = ~n59807 & n60736;
  assign n60738 = n59820 & n60737;
  assign n60739 = ~n59820 & n59848;
  assign n60740 = ~n59862 & ~n60739;
  assign n60741 = ~n60020 & n60740;
  assign n60742 = ~n59826 & ~n60741;
  assign n60743 = n59795 & n60742;
  assign n60744 = n59826 & n60018;
  assign n60745 = ~n59844 & ~n59870;
  assign n60746 = ~n59839 & n60745;
  assign n60747 = ~n60744 & n60746;
  assign n60748 = n59795 & ~n60747;
  assign n60749 = ~n59820 & n59881;
  assign n60750 = ~n60737 & ~n60749;
  assign n60751 = ~n60008 & n60750;
  assign n60752 = n59813 & n59843;
  assign n60753 = ~n59820 & n59831;
  assign n60754 = ~n59858 & ~n60753;
  assign n60755 = ~n59826 & ~n60754;
  assign n60756 = ~n60752 & ~n60755;
  assign n60757 = n60751 & n60756;
  assign n60758 = ~n59795 & ~n60757;
  assign n60759 = ~n60748 & ~n60758;
  assign n60760 = ~n60743 & n60759;
  assign n60761 = ~n60738 & n60760;
  assign n60762 = n60734 & n60761;
  assign n60763 = pi1718 & ~n60762;
  assign n60764 = ~pi1718 & n60734;
  assign n60765 = n60761 & n60764;
  assign po1810 = n60763 | n60765;
  assign n60767 = ~n59325 & ~n59331;
  assign n60768 = ~n59298 & ~n60767;
  assign n60769 = ~n59387 & ~n60768;
  assign n60770 = n59304 & n59310;
  assign n60771 = n59298 & n60770;
  assign n60772 = n59324 & n60771;
  assign n60773 = n59324 & n59350;
  assign n60774 = ~n60770 & ~n60773;
  assign n60775 = ~n59304 & ~n59324;
  assign n60776 = ~n59310 & n60775;
  assign n60777 = n60774 & ~n60776;
  assign n60778 = n59298 & ~n60777;
  assign n60779 = ~n59334 & ~n60778;
  assign n60780 = ~n59363 & ~n60779;
  assign n60781 = ~n59298 & n59317;
  assign n60782 = n59324 & n60781;
  assign n60783 = ~n60627 & ~n60782;
  assign n60784 = ~n59363 & ~n60783;
  assign n60785 = ~n60780 & ~n60784;
  assign n60786 = ~n60772 & n60785;
  assign n60787 = ~n59351 & ~n59370;
  assign n60788 = ~n59380 & n60787;
  assign n60789 = ~n59298 & ~n60788;
  assign n60790 = ~n59324 & n59375;
  assign n60791 = ~n59354 & ~n60790;
  assign n60792 = n59298 & ~n60791;
  assign n60793 = ~n60641 & ~n60792;
  assign n60794 = ~n60789 & n60793;
  assign n60795 = ~n59340 & ~n59381;
  assign n60796 = n60794 & n60795;
  assign n60797 = n59363 & ~n60796;
  assign n60798 = n60786 & ~n60797;
  assign n60799 = n60769 & n60798;
  assign n60800 = ~pi1713 & ~n60799;
  assign n60801 = pi1713 & n60786;
  assign n60802 = n60769 & n60801;
  assign n60803 = ~n60797 & n60802;
  assign po1811 = n60800 | n60803;
  assign n60805 = ~n59518 & n59539;
  assign n60806 = ~n60407 & ~n60805;
  assign n60807 = n59524 & n60806;
  assign n60808 = n59518 & n59576;
  assign n60809 = ~n59512 & ~n59533;
  assign n60810 = ~n59532 & ~n60809;
  assign n60811 = n59505 & n59558;
  assign n60812 = n59518 & n59533;
  assign n60813 = ~n60811 & ~n60812;
  assign n60814 = ~n60810 & n60813;
  assign n60815 = ~n60808 & n60814;
  assign n60816 = ~n59524 & n60815;
  assign n60817 = ~n60807 & ~n60816;
  assign n60818 = n59518 & n60810;
  assign n60819 = ~n60405 & ~n60818;
  assign n60820 = ~n60817 & n60819;
  assign n60821 = n59499 & ~n60820;
  assign n60822 = n59524 & ~n60809;
  assign n60823 = ~n59518 & n60822;
  assign n60824 = ~n59553 & ~n59564;
  assign n60825 = n59518 & ~n60824;
  assign n60826 = n59524 & n60825;
  assign n60827 = n59532 & n60822;
  assign n60828 = ~n60826 & ~n60827;
  assign n60829 = ~n60823 & n60828;
  assign n60830 = ~n59499 & ~n60829;
  assign n60831 = ~n60821 & ~n60830;
  assign n60832 = ~n59524 & ~n60806;
  assign n60833 = ~n59537 & ~n60832;
  assign n60834 = ~n59499 & ~n60833;
  assign n60835 = n59524 & n59537;
  assign n60836 = ~n59524 & ~n60819;
  assign n60837 = ~n60835 & ~n60836;
  assign n60838 = ~n60834 & n60837;
  assign n60839 = n60831 & n60838;
  assign n60840 = pi1706 & ~n60839;
  assign n60841 = ~n60821 & n60838;
  assign n60842 = ~n60830 & n60841;
  assign n60843 = ~pi1706 & n60842;
  assign po1812 = n60840 | n60843;
  assign n60845 = n60231 & n60296;
  assign n60846 = ~n60501 & ~n60845;
  assign n60847 = ~n60225 & ~n60846;
  assign n60848 = n60231 & n60262;
  assign n60849 = ~n60245 & ~n60848;
  assign n60850 = ~n60225 & ~n60849;
  assign n60851 = ~n60219 & n60263;
  assign n60852 = ~n60281 & ~n60851;
  assign n60853 = ~n60253 & n60852;
  assign n60854 = n60225 & ~n60853;
  assign n60855 = ~n60850 & ~n60854;
  assign n60856 = ~n60480 & ~n60487;
  assign n60857 = n60855 & n60856;
  assign n60858 = ~n60278 & ~n60857;
  assign n60859 = n60219 & n60245;
  assign n60860 = ~n60219 & n60285;
  assign n60861 = ~n60296 & ~n60860;
  assign n60862 = n60225 & ~n60861;
  assign n60863 = ~n60859 & ~n60862;
  assign n60864 = ~n60225 & n60299;
  assign n60865 = n60472 & ~n60864;
  assign n60866 = ~n60253 & n60865;
  assign n60867 = ~n60219 & ~n60866;
  assign n60868 = n60863 & ~n60867;
  assign n60869 = n60278 & ~n60868;
  assign n60870 = ~n60858 & ~n60869;
  assign n60871 = n60225 & n60521;
  assign n60872 = n60219 & n60871;
  assign n60873 = n60870 & ~n60872;
  assign n60874 = ~n60847 & n60873;
  assign n60875 = ~pi1733 & ~n60874;
  assign n60876 = pi1733 & ~n60847;
  assign n60877 = n60870 & n60876;
  assign n60878 = ~n60872 & n60877;
  assign po1813 = n60875 | n60878;
  assign n60880 = n59518 & n60409;
  assign n60881 = n59524 & n60880;
  assign n60882 = n59558 & ~n60809;
  assign n60883 = ~n59580 & ~n60882;
  assign n60884 = ~n60405 & n60883;
  assign n60885 = ~n59524 & ~n60884;
  assign n60886 = n59518 & n59534;
  assign n60887 = ~n60885 & ~n60886;
  assign n60888 = n59532 & n59564;
  assign n60889 = ~n59518 & n60413;
  assign n60890 = ~n60888 & ~n60889;
  assign n60891 = ~n60812 & n60890;
  assign n60892 = n59524 & ~n60891;
  assign n60893 = n60887 & ~n60892;
  assign n60894 = n59499 & ~n60893;
  assign n60895 = ~n60881 & ~n60894;
  assign n60896 = ~n59518 & n59533;
  assign n60897 = ~n60404 & ~n60896;
  assign n60898 = n59524 & ~n60897;
  assign n60899 = ~n59581 & ~n60898;
  assign n60900 = ~n59554 & ~n60880;
  assign n60901 = ~n59518 & n59534;
  assign n60902 = n59518 & n59586;
  assign n60903 = ~n60413 & ~n60902;
  assign n60904 = ~n60888 & n60903;
  assign n60905 = ~n59524 & ~n60904;
  assign n60906 = ~n60901 & ~n60905;
  assign n60907 = n60900 & n60906;
  assign n60908 = n60899 & n60907;
  assign n60909 = ~n59499 & ~n60908;
  assign n60910 = ~n59568 & ~n60808;
  assign n60911 = ~n59524 & ~n60910;
  assign n60912 = ~n60909 & ~n60911;
  assign n60913 = n60895 & n60912;
  assign n60914 = pi1705 & n60913;
  assign n60915 = ~pi1705 & ~n60913;
  assign po1814 = n60914 | n60915;
  assign n60917 = ~n60181 & ~n60458;
  assign n60918 = ~n60438 & n60917;
  assign n60919 = ~n59434 & ~n60918;
  assign n60920 = ~n60189 & ~n60206;
  assign n60921 = ~n60187 & ~n60446;
  assign n60922 = ~n60175 & ~n60451;
  assign n60923 = n59434 & ~n60922;
  assign n60924 = ~n59463 & ~n60923;
  assign n60925 = n60921 & n60924;
  assign n60926 = n59399 & ~n60925;
  assign n60927 = ~n59417 & n59423;
  assign n60928 = ~n59447 & ~n60927;
  assign n60929 = n59405 & ~n60928;
  assign n60930 = ~n59425 & ~n60192;
  assign n60931 = n59434 & ~n60930;
  assign n60932 = n59405 & n59423;
  assign n60933 = ~n59437 & ~n60932;
  assign n60934 = ~n59444 & n60933;
  assign n60935 = ~n59434 & ~n60934;
  assign n60936 = ~n60931 & ~n60935;
  assign n60937 = ~n60929 & n60936;
  assign n60938 = ~n59399 & ~n60937;
  assign n60939 = ~n60926 & ~n60938;
  assign n60940 = n60920 & n60939;
  assign n60941 = ~n60919 & n60940;
  assign n60942 = ~pi1735 & ~n60941;
  assign n60943 = pi1735 & n60920;
  assign n60944 = ~n60919 & n60943;
  assign n60945 = n60939 & n60944;
  assign po1815 = n60942 | n60945;
  assign n60947 = ~n59724 & n59746;
  assign n60948 = ~n59745 & ~n60947;
  assign n60949 = ~n59705 & ~n60948;
  assign n60950 = n59705 & ~n60072;
  assign n60951 = ~n60082 & ~n60950;
  assign n60952 = ~n60949 & n60951;
  assign n60953 = n59742 & ~n60952;
  assign n60954 = ~n59705 & n59760;
  assign n60955 = ~n60953 & ~n60954;
  assign n60956 = ~n60145 & ~n60160;
  assign n60957 = n59705 & ~n60956;
  assign n60958 = n59705 & n59747;
  assign n60959 = n59717 & n59733;
  assign n60960 = n59711 & n60959;
  assign n60961 = ~n59705 & n59731;
  assign n60962 = ~n60053 & ~n60961;
  assign n60963 = ~n59711 & ~n60962;
  assign n60964 = ~n60054 & ~n60963;
  assign n60965 = ~n59732 & n60964;
  assign n60966 = ~n60960 & n60965;
  assign n60967 = ~n60958 & n60966;
  assign n60968 = ~n59742 & ~n60967;
  assign n60969 = ~n60957 & ~n60968;
  assign n60970 = n60955 & n60969;
  assign n60971 = pi1737 & ~n60970;
  assign n60972 = ~pi1737 & n60970;
  assign po1816 = n60971 | n60972;
  assign n60974 = ~n59381 & ~n60647;
  assign n60975 = n59298 & ~n60974;
  assign n60976 = ~n59328 & ~n59331;
  assign n60977 = ~n59324 & n59380;
  assign n60978 = ~n60617 & ~n60977;
  assign n60979 = n60976 & n60978;
  assign n60980 = ~n59298 & ~n60979;
  assign n60981 = ~n59363 & n59365;
  assign n60982 = ~n59298 & n60981;
  assign n60983 = n59310 & n60775;
  assign n60984 = ~n60643 & ~n60983;
  assign n60985 = ~n59333 & n60984;
  assign n60986 = n59298 & ~n60985;
  assign n60987 = n59304 & n59350;
  assign n60988 = ~n59324 & n60987;
  assign n60989 = ~n60986 & ~n60988;
  assign n60990 = ~n59363 & ~n60989;
  assign n60991 = ~n60982 & ~n60990;
  assign n60992 = n59304 & ~n59310;
  assign n60993 = ~n59298 & n60992;
  assign n60994 = n59324 & n60993;
  assign n60995 = ~n59324 & n60643;
  assign n60996 = ~n59331 & ~n60995;
  assign n60997 = ~n60638 & n60996;
  assign n60998 = ~n60994 & n60997;
  assign n60999 = n59298 & n59327;
  assign n61000 = n60998 & ~n60999;
  assign n61001 = n59363 & ~n61000;
  assign n61002 = n60991 & ~n61001;
  assign n61003 = ~n60980 & n61002;
  assign n61004 = ~n60975 & n61003;
  assign n61005 = pi1720 & n61004;
  assign n61006 = ~pi1720 & ~n61004;
  assign po1817 = n61005 | n61006;
  assign n61008 = pi5938 & ~pi9040;
  assign n61009 = pi5941 & pi9040;
  assign n61010 = ~n61008 & ~n61009;
  assign n61011 = ~pi1738 & n61010;
  assign n61012 = pi1738 & ~n61010;
  assign n61013 = ~n61011 & ~n61012;
  assign n61014 = pi5824 & pi9040;
  assign n61015 = pi5929 & ~pi9040;
  assign n61016 = ~n61014 & ~n61015;
  assign n61017 = pi1725 & n61016;
  assign n61018 = ~pi1725 & ~n61016;
  assign n61019 = ~n61017 & ~n61018;
  assign n61020 = pi5913 & pi9040;
  assign n61021 = pi5945 & ~pi9040;
  assign n61022 = ~n61020 & ~n61021;
  assign n61023 = pi1756 & n61022;
  assign n61024 = ~pi1756 & ~n61022;
  assign n61025 = ~n61023 & ~n61024;
  assign n61026 = pi5943 & pi9040;
  assign n61027 = pi6012 & ~pi9040;
  assign n61028 = ~n61026 & ~n61027;
  assign n61029 = ~pi1732 & n61028;
  assign n61030 = pi1732 & ~n61028;
  assign n61031 = ~n61029 & ~n61030;
  assign n61032 = n61025 & ~n61031;
  assign n61033 = ~n61019 & n61032;
  assign n61034 = pi5940 & pi9040;
  assign n61035 = pi5909 & ~pi9040;
  assign n61036 = ~n61034 & ~n61035;
  assign n61037 = pi1754 & n61036;
  assign n61038 = ~pi1754 & ~n61036;
  assign n61039 = ~n61037 & ~n61038;
  assign n61040 = n61033 & ~n61039;
  assign n61041 = ~n61019 & ~n61039;
  assign n61042 = n61031 & n61041;
  assign n61043 = ~n61025 & n61042;
  assign n61044 = ~n61040 & ~n61043;
  assign n61045 = ~n61025 & n61031;
  assign n61046 = n61019 & n61039;
  assign n61047 = n61045 & n61046;
  assign n61048 = n61025 & n61031;
  assign n61049 = ~n61019 & n61048;
  assign n61050 = n61039 & n61049;
  assign n61051 = ~n61047 & ~n61050;
  assign n61052 = n61044 & n61051;
  assign n61053 = ~n61013 & ~n61052;
  assign n61054 = ~n61025 & ~n61031;
  assign n61055 = ~n61019 & n61054;
  assign n61056 = n61039 & n61055;
  assign n61057 = ~n61049 & ~n61056;
  assign n61058 = ~n61013 & ~n61057;
  assign n61059 = n61013 & ~n61031;
  assign n61060 = ~n61039 & n61059;
  assign n61061 = n61019 & n61025;
  assign n61062 = n61039 & n61045;
  assign n61063 = ~n61061 & ~n61062;
  assign n61064 = n61013 & ~n61063;
  assign n61065 = ~n61060 & ~n61064;
  assign n61066 = n61019 & n61054;
  assign n61067 = ~n61039 & n61066;
  assign n61068 = n61065 & ~n61067;
  assign n61069 = ~n61031 & n61061;
  assign n61070 = n61039 & n61069;
  assign n61071 = n61068 & ~n61070;
  assign n61072 = ~n61058 & n61071;
  assign n61073 = pi5843 & pi9040;
  assign n61074 = ~pi5835 & ~pi9040;
  assign n61075 = ~n61073 & ~n61074;
  assign n61076 = ~pi1742 & ~n61075;
  assign n61077 = pi1742 & n61075;
  assign n61078 = ~n61076 & ~n61077;
  assign n61079 = ~n61072 & ~n61078;
  assign n61080 = ~n61019 & ~n61031;
  assign n61081 = n61013 & n61039;
  assign n61082 = n61078 & n61081;
  assign n61083 = n61080 & n61082;
  assign n61084 = n61013 & ~n61042;
  assign n61085 = ~n61025 & n61046;
  assign n61086 = ~n61032 & ~n61080;
  assign n61087 = ~n61039 & ~n61086;
  assign n61088 = n61019 & n61045;
  assign n61089 = ~n61013 & ~n61088;
  assign n61090 = ~n61087 & n61089;
  assign n61091 = ~n61085 & n61090;
  assign n61092 = ~n61084 & ~n61091;
  assign n61093 = n61019 & n61048;
  assign n61094 = n61039 & n61093;
  assign n61095 = ~n61092 & ~n61094;
  assign n61096 = n61078 & ~n61095;
  assign n61097 = ~n61083 & ~n61096;
  assign n61098 = ~n61079 & n61097;
  assign n61099 = ~n61053 & n61098;
  assign n61100 = n61013 & n61067;
  assign n61101 = n61099 & ~n61100;
  assign n61102 = pi1761 & ~n61101;
  assign n61103 = ~pi1761 & ~n61100;
  assign n61104 = n61098 & n61103;
  assign n61105 = ~n61053 & n61104;
  assign po1838 = n61102 | n61105;
  assign n61107 = pi5921 & pi9040;
  assign n61108 = pi5832 & ~pi9040;
  assign n61109 = ~n61107 & ~n61108;
  assign n61110 = ~pi1748 & ~n61109;
  assign n61111 = pi1748 & n61109;
  assign n61112 = ~n61110 & ~n61111;
  assign n61113 = pi5827 & pi9040;
  assign n61114 = pi5840 & ~pi9040;
  assign n61115 = ~n61113 & ~n61114;
  assign n61116 = pi1756 & n61115;
  assign n61117 = ~pi1756 & ~n61115;
  assign n61118 = ~n61116 & ~n61117;
  assign n61119 = pi5918 & ~pi9040;
  assign n61120 = pi6080 & pi9040;
  assign n61121 = ~n61119 & ~n61120;
  assign n61122 = ~pi1742 & ~n61121;
  assign n61123 = pi1742 & n61121;
  assign n61124 = ~n61122 & ~n61123;
  assign n61125 = pi5923 & pi9040;
  assign n61126 = pi6069 & ~pi9040;
  assign n61127 = ~n61125 & ~n61126;
  assign n61128 = ~pi1702 & n61127;
  assign n61129 = pi1702 & ~n61127;
  assign n61130 = ~n61128 & ~n61129;
  assign n61131 = ~n61124 & ~n61130;
  assign n61132 = pi5823 & pi9040;
  assign n61133 = pi5937 & ~pi9040;
  assign n61134 = ~n61132 & ~n61133;
  assign n61135 = ~pi1747 & n61134;
  assign n61136 = pi1747 & ~n61134;
  assign n61137 = ~n61135 & ~n61136;
  assign n61138 = pi5833 & pi9040;
  assign n61139 = pi5921 & ~pi9040;
  assign n61140 = ~n61138 & ~n61139;
  assign n61141 = pi1758 & n61140;
  assign n61142 = ~pi1758 & ~n61140;
  assign n61143 = ~n61141 & ~n61142;
  assign n61144 = ~n61137 & n61143;
  assign n61145 = n61131 & n61144;
  assign n61146 = n61118 & n61145;
  assign n61147 = n61137 & n61143;
  assign n61148 = n61124 & ~n61130;
  assign n61149 = n61147 & n61148;
  assign n61150 = n61118 & n61137;
  assign n61151 = n61130 & n61150;
  assign n61152 = ~n61124 & n61151;
  assign n61153 = n61124 & n61130;
  assign n61154 = n61118 & n61153;
  assign n61155 = n61143 & n61154;
  assign n61156 = ~n61137 & n61155;
  assign n61157 = ~n61152 & ~n61156;
  assign n61158 = ~n61149 & n61157;
  assign n61159 = ~n61146 & n61158;
  assign n61160 = ~n61118 & n61137;
  assign n61161 = ~n61130 & n61160;
  assign n61162 = n61124 & n61161;
  assign n61163 = n61159 & ~n61162;
  assign n61164 = ~n61112 & ~n61163;
  assign n61165 = n61118 & n61124;
  assign n61166 = ~n61130 & n61165;
  assign n61167 = ~n61137 & n61166;
  assign n61168 = ~n61151 & ~n61167;
  assign n61169 = ~n61118 & n61131;
  assign n61170 = ~n61137 & n61169;
  assign n61171 = n61168 & ~n61170;
  assign n61172 = ~n61143 & ~n61171;
  assign n61173 = ~n61118 & n61130;
  assign n61174 = n61124 & n61173;
  assign n61175 = ~n61143 & n61174;
  assign n61176 = ~n61137 & n61175;
  assign n61177 = ~n61124 & n61150;
  assign n61178 = ~n61124 & n61130;
  assign n61179 = n61137 & n61178;
  assign n61180 = ~n61177 & ~n61179;
  assign n61181 = ~n61143 & ~n61180;
  assign n61182 = ~n61176 & ~n61181;
  assign n61183 = ~n61112 & ~n61182;
  assign n61184 = ~n61172 & ~n61183;
  assign n61185 = ~n61164 & n61184;
  assign n61186 = ~n61118 & ~n61137;
  assign n61187 = n61143 & n61186;
  assign n61188 = n61178 & n61187;
  assign n61189 = ~n61118 & n61124;
  assign n61190 = n61147 & n61189;
  assign n61191 = n61137 & n61174;
  assign n61192 = n61118 & ~n61143;
  assign n61193 = n61124 & n61192;
  assign n61194 = ~n61124 & ~n61137;
  assign n61195 = ~n61118 & n61194;
  assign n61196 = ~n61193 & ~n61195;
  assign n61197 = ~n61191 & n61196;
  assign n61198 = ~n61169 & n61197;
  assign n61199 = n61131 & n61143;
  assign n61200 = n61137 & n61199;
  assign n61201 = ~n61137 & n61178;
  assign n61202 = ~n61118 & ~n61130;
  assign n61203 = ~n61201 & ~n61202;
  assign n61204 = n61143 & ~n61203;
  assign n61205 = ~n61200 & ~n61204;
  assign n61206 = n61198 & n61205;
  assign n61207 = n61112 & ~n61206;
  assign n61208 = ~n61190 & ~n61207;
  assign n61209 = ~n61188 & n61208;
  assign n61210 = n61185 & n61209;
  assign n61211 = pi1764 & n61210;
  assign n61212 = ~pi1764 & ~n61210;
  assign po1843 = n61211 | n61212;
  assign n61214 = n61118 & ~n61124;
  assign n61215 = ~n61162 & ~n61214;
  assign n61216 = ~n61194 & n61215;
  assign n61217 = n61143 & ~n61216;
  assign n61218 = ~n61137 & ~n61143;
  assign n61219 = n61124 & n61218;
  assign n61220 = n61118 & ~n61137;
  assign n61221 = ~n61130 & n61220;
  assign n61222 = n61137 & n61154;
  assign n61223 = ~n61221 & ~n61222;
  assign n61224 = ~n61118 & ~n61124;
  assign n61225 = n61137 & ~n61143;
  assign n61226 = n61224 & n61225;
  assign n61227 = n61223 & ~n61226;
  assign n61228 = ~n61219 & n61227;
  assign n61229 = ~n61217 & n61228;
  assign n61230 = n61112 & ~n61229;
  assign n61231 = n61118 & n61131;
  assign n61232 = n61137 & n61231;
  assign n61233 = n61118 & n61178;
  assign n61234 = ~n61137 & n61233;
  assign n61235 = ~n61232 & ~n61234;
  assign n61236 = n61143 & ~n61235;
  assign n61237 = ~n61230 & ~n61236;
  assign n61238 = ~n61137 & n61154;
  assign n61239 = ~n61166 & ~n61174;
  assign n61240 = n61143 & ~n61239;
  assign n61241 = ~n61238 & ~n61240;
  assign n61242 = ~n61170 & n61241;
  assign n61243 = ~n61112 & ~n61242;
  assign n61244 = ~n61148 & ~n61178;
  assign n61245 = ~n61118 & ~n61244;
  assign n61246 = ~n61179 & ~n61245;
  assign n61247 = ~n61143 & ~n61246;
  assign n61248 = ~n61112 & n61247;
  assign n61249 = ~n61243 & ~n61248;
  assign n61250 = n61237 & n61249;
  assign n61251 = pi1770 & ~n61250;
  assign n61252 = ~pi1770 & n61237;
  assign n61253 = n61249 & n61252;
  assign po1845 = n61251 | n61253;
  assign n61255 = pi5917 & ~pi9040;
  assign n61256 = pi5819 & pi9040;
  assign n61257 = ~n61255 & ~n61256;
  assign n61258 = ~pi1743 & ~n61257;
  assign n61259 = pi1743 & n61257;
  assign n61260 = ~n61258 & ~n61259;
  assign n61261 = pi5948 & ~pi9040;
  assign n61262 = pi5818 & pi9040;
  assign n61263 = ~n61261 & ~n61262;
  assign n61264 = pi1752 & n61263;
  assign n61265 = ~pi1752 & ~n61263;
  assign n61266 = pi5823 & ~pi9040;
  assign n61267 = pi5832 & pi9040;
  assign n61268 = ~n61266 & ~n61267;
  assign n61269 = pi1736 & n61268;
  assign n61270 = ~pi1736 & ~n61268;
  assign n61271 = ~n61269 & ~n61270;
  assign n61272 = ~n61265 & ~n61271;
  assign n61273 = ~n61264 & n61272;
  assign n61274 = pi6069 & pi9040;
  assign n61275 = pi5818 & ~pi9040;
  assign n61276 = ~n61274 & ~n61275;
  assign n61277 = pi1755 & n61276;
  assign n61278 = ~pi1755 & ~n61276;
  assign n61279 = ~n61277 & ~n61278;
  assign n61280 = pi5836 & pi9040;
  assign n61281 = pi5946 & ~pi9040;
  assign n61282 = ~n61280 & ~n61281;
  assign n61283 = ~pi1748 & ~n61282;
  assign n61284 = pi1748 & n61282;
  assign n61285 = ~n61283 & ~n61284;
  assign n61286 = ~n61279 & ~n61285;
  assign n61287 = pi5923 & ~pi9040;
  assign n61288 = pi5911 & pi9040;
  assign n61289 = ~n61287 & ~n61288;
  assign n61290 = ~pi1702 & n61289;
  assign n61291 = pi1702 & ~n61289;
  assign n61292 = ~n61290 & ~n61291;
  assign n61293 = n61279 & n61285;
  assign n61294 = n61292 & n61293;
  assign n61295 = ~n61286 & ~n61294;
  assign n61296 = n61273 & ~n61295;
  assign n61297 = ~n61271 & n61292;
  assign n61298 = n61286 & n61297;
  assign n61299 = ~n61296 & ~n61298;
  assign n61300 = n61260 & ~n61299;
  assign n61301 = ~n61264 & ~n61265;
  assign n61302 = ~n61292 & ~n61301;
  assign n61303 = n61279 & n61302;
  assign n61304 = n61285 & n61303;
  assign n61305 = n61285 & ~n61292;
  assign n61306 = ~n61302 & ~n61305;
  assign n61307 = n61271 & ~n61306;
  assign n61308 = n61292 & ~n61301;
  assign n61309 = ~n61279 & n61308;
  assign n61310 = n61285 & n61309;
  assign n61311 = ~n61307 & ~n61310;
  assign n61312 = ~n61304 & n61311;
  assign n61313 = n61260 & ~n61312;
  assign n61314 = ~n61300 & ~n61313;
  assign n61315 = ~n61292 & n61301;
  assign n61316 = n61279 & n61315;
  assign n61317 = ~n61285 & n61316;
  assign n61318 = n61279 & ~n61285;
  assign n61319 = n61292 & n61318;
  assign n61320 = ~n61301 & n61319;
  assign n61321 = ~n61317 & ~n61320;
  assign n61322 = ~n61271 & ~n61321;
  assign n61323 = ~n61279 & n61285;
  assign n61324 = ~n61305 & ~n61323;
  assign n61325 = n61301 & ~n61324;
  assign n61326 = ~n61319 & ~n61325;
  assign n61327 = ~n61271 & ~n61326;
  assign n61328 = n61279 & ~n61301;
  assign n61329 = n61297 & n61328;
  assign n61330 = ~n61279 & ~n61292;
  assign n61331 = ~n61319 & ~n61330;
  assign n61332 = ~n61301 & ~n61331;
  assign n61333 = n61271 & n61301;
  assign n61334 = n61293 & n61333;
  assign n61335 = n61292 & n61334;
  assign n61336 = ~n61332 & ~n61335;
  assign n61337 = ~n61329 & n61336;
  assign n61338 = ~n61327 & n61337;
  assign n61339 = ~n61317 & n61338;
  assign n61340 = ~n61260 & ~n61339;
  assign n61341 = n61286 & n61292;
  assign n61342 = n61301 & n61341;
  assign n61343 = ~n61301 & n61305;
  assign n61344 = ~n61342 & ~n61343;
  assign n61345 = n61271 & ~n61344;
  assign n61346 = ~n61340 & ~n61345;
  assign n61347 = ~n61322 & n61346;
  assign n61348 = n61314 & n61347;
  assign n61349 = pi1771 & n61348;
  assign n61350 = ~pi1771 & ~n61348;
  assign po1847 = n61349 | n61350;
  assign n61352 = pi5929 & pi9040;
  assign n61353 = pi5842 & ~pi9040;
  assign n61354 = ~n61352 & ~n61353;
  assign n61355 = ~pi1744 & ~n61354;
  assign n61356 = pi1744 & n61354;
  assign n61357 = ~n61355 & ~n61356;
  assign n61358 = pi5837 & pi9040;
  assign n61359 = pi5941 & ~pi9040;
  assign n61360 = ~n61358 & ~n61359;
  assign n61361 = ~pi1759 & n61360;
  assign n61362 = pi1759 & ~n61360;
  assign n61363 = ~n61361 & ~n61362;
  assign n61364 = pi5842 & pi9040;
  assign n61365 = pi5843 & ~pi9040;
  assign n61366 = ~n61364 & ~n61365;
  assign n61367 = ~pi1746 & ~n61366;
  assign n61368 = pi1746 & n61366;
  assign n61369 = ~n61367 & ~n61368;
  assign n61370 = pi5943 & ~pi9040;
  assign n61371 = pi5938 & pi9040;
  assign n61372 = ~n61370 & ~n61371;
  assign n61373 = ~pi1757 & ~n61372;
  assign n61374 = pi1757 & n61372;
  assign n61375 = ~n61373 & ~n61374;
  assign n61376 = pi5913 & ~pi9040;
  assign n61377 = pi5909 & pi9040;
  assign n61378 = ~n61376 & ~n61377;
  assign n61379 = ~pi1724 & ~n61378;
  assign n61380 = pi1724 & n61378;
  assign n61381 = ~n61379 & ~n61380;
  assign n61382 = ~n61375 & ~n61381;
  assign n61383 = n61369 & n61382;
  assign n61384 = ~n61363 & n61383;
  assign n61385 = ~n61375 & n61381;
  assign n61386 = ~n61363 & ~n61369;
  assign n61387 = n61385 & n61386;
  assign n61388 = ~n61384 & ~n61387;
  assign n61389 = n61375 & n61381;
  assign n61390 = ~n61369 & n61389;
  assign n61391 = n61363 & ~n61369;
  assign n61392 = ~n61381 & n61391;
  assign n61393 = ~n61375 & n61392;
  assign n61394 = ~n61390 & ~n61393;
  assign n61395 = pi5824 & ~pi9040;
  assign n61396 = pi5945 & pi9040;
  assign n61397 = ~n61395 & ~n61396;
  assign n61398 = ~pi1734 & n61397;
  assign n61399 = pi1734 & ~n61397;
  assign n61400 = ~n61398 & ~n61399;
  assign n61401 = ~n61394 & ~n61400;
  assign n61402 = n61388 & ~n61401;
  assign n61403 = n61363 & n61400;
  assign n61404 = n61375 & n61403;
  assign n61405 = n61402 & ~n61404;
  assign n61406 = n61357 & ~n61405;
  assign n61407 = n61375 & ~n61381;
  assign n61408 = ~n61369 & n61407;
  assign n61409 = ~n61363 & n61408;
  assign n61410 = n61400 & n61409;
  assign n61411 = n61363 & ~n61400;
  assign n61412 = n61408 & n61411;
  assign n61413 = n61363 & n61369;
  assign n61414 = ~n61375 & n61413;
  assign n61415 = ~n61412 & ~n61414;
  assign n61416 = n61369 & n61385;
  assign n61417 = ~n61390 & ~n61416;
  assign n61418 = n61363 & n61385;
  assign n61419 = n61417 & ~n61418;
  assign n61420 = n61400 & ~n61419;
  assign n61421 = n61369 & ~n61381;
  assign n61422 = n61375 & n61421;
  assign n61423 = ~n61363 & n61422;
  assign n61424 = ~n61381 & n61386;
  assign n61425 = ~n61375 & n61424;
  assign n61426 = ~n61423 & ~n61425;
  assign n61427 = n61369 & n61389;
  assign n61428 = ~n61400 & n61427;
  assign n61429 = n61426 & ~n61428;
  assign n61430 = ~n61420 & n61429;
  assign n61431 = n61415 & n61430;
  assign n61432 = ~n61357 & ~n61431;
  assign n61433 = ~n61410 & ~n61432;
  assign n61434 = ~n61406 & n61433;
  assign n61435 = n61411 & n61416;
  assign n61436 = ~n61400 & n61421;
  assign n61437 = ~n61363 & n61436;
  assign n61438 = ~n61435 & ~n61437;
  assign n61439 = n61387 & ~n61400;
  assign n61440 = n61438 & ~n61439;
  assign n61441 = n61434 & n61440;
  assign n61442 = ~pi1768 & ~n61441;
  assign n61443 = pi1768 & n61440;
  assign n61444 = n61433 & n61443;
  assign n61445 = ~n61406 & n61444;
  assign po1848 = n61442 | n61445;
  assign n61447 = n61363 & n61383;
  assign n61448 = ~n61369 & n61385;
  assign n61449 = n61363 & n61427;
  assign n61450 = ~n61448 & ~n61449;
  assign n61451 = ~n61363 & n61421;
  assign n61452 = n61363 & n61408;
  assign n61453 = ~n61451 & ~n61452;
  assign n61454 = n61450 & n61453;
  assign n61455 = n61400 & ~n61454;
  assign n61456 = ~n61369 & n61382;
  assign n61457 = ~n61363 & n61389;
  assign n61458 = ~n61414 & ~n61457;
  assign n61459 = ~n61456 & n61458;
  assign n61460 = ~n61400 & ~n61459;
  assign n61461 = n61381 & n61386;
  assign n61462 = n61375 & n61461;
  assign n61463 = ~n61460 & ~n61462;
  assign n61464 = ~n61455 & n61463;
  assign n61465 = ~n61447 & n61464;
  assign n61466 = ~n61357 & ~n61465;
  assign n61467 = n61400 & n61427;
  assign n61468 = ~n61363 & n61467;
  assign n61469 = n61400 & n61456;
  assign n61470 = n61400 & n61416;
  assign n61471 = ~n61469 & ~n61470;
  assign n61472 = n61363 & ~n61471;
  assign n61473 = ~n61468 & ~n61472;
  assign n61474 = ~n61363 & n61385;
  assign n61475 = n61363 & n61389;
  assign n61476 = ~n61474 & ~n61475;
  assign n61477 = ~n61422 & n61476;
  assign n61478 = ~n61448 & n61477;
  assign n61479 = ~n61400 & ~n61478;
  assign n61480 = n61363 & n61390;
  assign n61481 = ~n61479 & ~n61480;
  assign n61482 = n61363 & n61422;
  assign n61483 = ~n61409 & ~n61482;
  assign n61484 = n61481 & n61483;
  assign n61485 = n61473 & n61484;
  assign n61486 = n61357 & ~n61485;
  assign n61487 = ~n61388 & n61400;
  assign n61488 = ~n61486 & ~n61487;
  assign n61489 = ~n61425 & ~n61482;
  assign n61490 = ~n61400 & ~n61489;
  assign n61491 = n61488 & ~n61490;
  assign n61492 = ~n61466 & n61491;
  assign n61493 = pi1779 & ~n61492;
  assign n61494 = ~pi1779 & n61492;
  assign po1849 = n61493 | n61494;
  assign n61496 = n61381 & n61413;
  assign n61497 = ~n61390 & ~n61414;
  assign n61498 = n61400 & ~n61497;
  assign n61499 = ~n61496 & ~n61498;
  assign n61500 = ~n61369 & ~n61375;
  assign n61501 = ~n61369 & ~n61381;
  assign n61502 = n61363 & n61501;
  assign n61503 = ~n61363 & n61382;
  assign n61504 = ~n61502 & ~n61503;
  assign n61505 = ~n61500 & n61504;
  assign n61506 = ~n61427 & n61505;
  assign n61507 = ~n61400 & ~n61506;
  assign n61508 = n61499 & ~n61507;
  assign n61509 = ~n61423 & n61508;
  assign n61510 = n61357 & ~n61509;
  assign n61511 = n61363 & n61448;
  assign n61512 = n61426 & ~n61511;
  assign n61513 = ~n61400 & ~n61512;
  assign n61514 = ~n61510 & ~n61513;
  assign n61515 = ~n61369 & n61375;
  assign n61516 = n61400 & n61515;
  assign n61517 = ~n61363 & n61516;
  assign n61518 = ~n61363 & n61416;
  assign n61519 = n61363 & n61436;
  assign n61520 = ~n61518 & ~n61519;
  assign n61521 = n61369 & ~n61375;
  assign n61522 = ~n61363 & n61521;
  assign n61523 = ~n61408 & ~n61522;
  assign n61524 = n61400 & ~n61523;
  assign n61525 = n61400 & n61500;
  assign n61526 = n61363 & n61525;
  assign n61527 = ~n61524 & ~n61526;
  assign n61528 = n61520 & n61527;
  assign n61529 = ~n61357 & ~n61528;
  assign n61530 = ~n61517 & ~n61529;
  assign n61531 = ~n61449 & n61530;
  assign n61532 = n61514 & n61531;
  assign n61533 = ~pi1763 & ~n61532;
  assign n61534 = ~n61449 & ~n61510;
  assign n61535 = ~n61513 & n61534;
  assign n61536 = n61530 & n61535;
  assign n61537 = pi1763 & n61536;
  assign po1850 = n61533 | n61537;
  assign n61539 = n61286 & ~n61301;
  assign n61540 = ~n61292 & n61318;
  assign n61541 = ~n61539 & ~n61540;
  assign n61542 = ~n61260 & n61271;
  assign n61543 = ~n61541 & n61542;
  assign n61544 = n61315 & n61323;
  assign n61545 = ~n61294 & ~n61341;
  assign n61546 = n61301 & ~n61545;
  assign n61547 = ~n61544 & ~n61546;
  assign n61548 = ~n61260 & ~n61547;
  assign n61549 = ~n61543 & ~n61548;
  assign n61550 = n61292 & n61301;
  assign n61551 = ~n61285 & n61550;
  assign n61552 = ~n61544 & ~n61551;
  assign n61553 = ~n61271 & ~n61552;
  assign n61554 = n61271 & ~n61301;
  assign n61555 = n61285 & n61554;
  assign n61556 = n61292 & n61323;
  assign n61557 = ~n61292 & n61293;
  assign n61558 = ~n61556 & ~n61557;
  assign n61559 = n61286 & ~n61292;
  assign n61560 = n61301 & n61559;
  assign n61561 = n61558 & ~n61560;
  assign n61562 = n61271 & ~n61561;
  assign n61563 = ~n61555 & ~n61562;
  assign n61564 = n61301 & n61319;
  assign n61565 = n61563 & ~n61564;
  assign n61566 = ~n61271 & ~n61541;
  assign n61567 = n61294 & ~n61301;
  assign n61568 = ~n61566 & ~n61567;
  assign n61569 = n61565 & n61568;
  assign n61570 = n61260 & ~n61569;
  assign n61571 = ~n61553 & ~n61570;
  assign n61572 = ~n61260 & ~n61271;
  assign n61573 = ~n61301 & n61323;
  assign n61574 = ~n61319 & ~n61573;
  assign n61575 = ~n61305 & n61574;
  assign n61576 = n61572 & ~n61575;
  assign n61577 = n61571 & ~n61576;
  assign n61578 = n61549 & n61577;
  assign n61579 = ~pi1776 & ~n61578;
  assign n61580 = pi1776 & n61549;
  assign n61581 = n61571 & n61580;
  assign n61582 = ~n61576 & n61581;
  assign po1851 = n61579 | n61582;
  assign n61584 = ~pi5835 & pi9040;
  assign n61585 = pi5942 & ~pi9040;
  assign n61586 = ~n61584 & ~n61585;
  assign n61587 = ~pi1732 & ~n61586;
  assign n61588 = pi1732 & n61586;
  assign n61589 = ~n61587 & ~n61588;
  assign n61590 = pi6015 & pi9040;
  assign n61591 = pi5796 & ~pi9040;
  assign n61592 = ~n61590 & ~n61591;
  assign n61593 = ~pi1753 & n61592;
  assign n61594 = pi1753 & ~n61592;
  assign n61595 = ~n61593 & ~n61594;
  assign n61596 = pi5792 & ~pi9040;
  assign n61597 = pi6013 & pi9040;
  assign n61598 = ~n61596 & ~n61597;
  assign n61599 = pi1725 & n61598;
  assign n61600 = ~pi1725 & ~n61598;
  assign n61601 = ~n61599 & ~n61600;
  assign n61602 = n61595 & n61601;
  assign n61603 = pi6015 & ~pi9040;
  assign n61604 = pi5942 & pi9040;
  assign n61605 = ~n61603 & ~n61604;
  assign n61606 = pi1741 & n61605;
  assign n61607 = ~pi1741 & ~n61605;
  assign n61608 = ~n61606 & ~n61607;
  assign n61609 = pi5939 & ~pi9040;
  assign n61610 = pi5825 & pi9040;
  assign n61611 = ~n61609 & ~n61610;
  assign n61612 = pi1728 & n61611;
  assign n61613 = ~pi1728 & ~n61611;
  assign n61614 = ~n61612 & ~n61613;
  assign n61615 = ~n61608 & ~n61614;
  assign n61616 = n61602 & n61615;
  assign n61617 = pi5916 & ~pi9040;
  assign n61618 = pi5796 & pi9040;
  assign n61619 = ~n61617 & ~n61618;
  assign n61620 = ~pi1731 & n61619;
  assign n61621 = pi1731 & ~n61619;
  assign n61622 = ~n61620 & ~n61621;
  assign n61623 = ~n61595 & ~n61601;
  assign n61624 = ~n61622 & n61623;
  assign n61625 = n61608 & n61622;
  assign n61626 = ~n61601 & n61625;
  assign n61627 = n61595 & n61626;
  assign n61628 = ~n61624 & ~n61627;
  assign n61629 = ~n61595 & n61601;
  assign n61630 = n61608 & n61629;
  assign n61631 = n61628 & ~n61630;
  assign n61632 = ~n61614 & ~n61631;
  assign n61633 = ~n61595 & n61622;
  assign n61634 = ~n61608 & n61614;
  assign n61635 = n61633 & n61634;
  assign n61636 = n61622 & n61623;
  assign n61637 = ~n61608 & n61636;
  assign n61638 = ~n61635 & ~n61637;
  assign n61639 = ~n61632 & n61638;
  assign n61640 = ~n61616 & n61639;
  assign n61641 = n61602 & ~n61622;
  assign n61642 = ~n61608 & n61641;
  assign n61643 = ~n61622 & n61629;
  assign n61644 = n61608 & n61643;
  assign n61645 = ~n61642 & ~n61644;
  assign n61646 = n61640 & n61645;
  assign n61647 = ~n61589 & ~n61646;
  assign n61648 = ~n61608 & n61622;
  assign n61649 = n61601 & n61648;
  assign n61650 = ~n61595 & n61649;
  assign n61651 = ~n61641 & ~n61650;
  assign n61652 = ~n61614 & ~n61651;
  assign n61653 = n61602 & n61625;
  assign n61654 = ~n61601 & n61648;
  assign n61655 = n61595 & n61654;
  assign n61656 = ~n61653 & ~n61655;
  assign n61657 = ~n61595 & n61625;
  assign n61658 = ~n61608 & n61643;
  assign n61659 = ~n61657 & ~n61658;
  assign n61660 = n61614 & ~n61659;
  assign n61661 = n61656 & ~n61660;
  assign n61662 = ~n61652 & n61661;
  assign n61663 = n61589 & ~n61662;
  assign n61664 = ~n61595 & ~n61622;
  assign n61665 = n61608 & n61664;
  assign n61666 = n61595 & ~n61622;
  assign n61667 = ~n61608 & n61666;
  assign n61668 = ~n61665 & ~n61667;
  assign n61669 = ~n61614 & ~n61668;
  assign n61670 = n61595 & ~n61601;
  assign n61671 = ~n61622 & n61670;
  assign n61672 = n61608 & n61671;
  assign n61673 = ~n61653 & ~n61672;
  assign n61674 = ~n61636 & n61673;
  assign n61675 = n61614 & ~n61674;
  assign n61676 = ~n61669 & ~n61675;
  assign n61677 = ~n61601 & n61622;
  assign n61678 = n61614 & n61677;
  assign n61679 = ~n61608 & n61678;
  assign n61680 = n61676 & ~n61679;
  assign n61681 = ~n61663 & n61680;
  assign n61682 = ~n61647 & n61681;
  assign n61683 = ~pi1765 & ~n61682;
  assign n61684 = pi1765 & n61682;
  assign po1853 = n61683 | n61684;
  assign n61686 = pi5940 & ~pi9040;
  assign n61687 = pi5947 & pi9040;
  assign n61688 = ~n61686 & ~n61687;
  assign n61689 = pi1749 & n61688;
  assign n61690 = ~pi1749 & ~n61688;
  assign n61691 = ~n61689 & ~n61690;
  assign n61692 = pi5939 & pi9040;
  assign n61693 = pi5816 & ~pi9040;
  assign n61694 = ~n61692 & ~n61693;
  assign n61695 = ~pi1753 & ~n61694;
  assign n61696 = pi1753 & n61694;
  assign n61697 = ~n61695 & ~n61696;
  assign n61698 = ~n61691 & ~n61697;
  assign n61699 = pi6012 & pi9040;
  assign n61700 = pi5825 & ~pi9040;
  assign n61701 = ~n61699 & ~n61700;
  assign n61702 = ~pi1709 & ~n61701;
  assign n61703 = pi1709 & n61701;
  assign n61704 = ~n61702 & ~n61703;
  assign n61705 = pi5792 & pi9040;
  assign n61706 = pi5831 & ~pi9040;
  assign n61707 = ~n61705 & ~n61706;
  assign n61708 = pi1744 & n61707;
  assign n61709 = ~pi1744 & ~n61707;
  assign n61710 = ~n61708 & ~n61709;
  assign n61711 = pi5821 & pi9040;
  assign n61712 = pi5947 & ~pi9040;
  assign n61713 = ~n61711 & ~n61712;
  assign n61714 = ~pi1724 & ~n61713;
  assign n61715 = pi1724 & n61713;
  assign n61716 = ~n61714 & ~n61715;
  assign n61717 = ~n61710 & n61716;
  assign n61718 = ~n61704 & n61717;
  assign n61719 = pi5920 & pi9040;
  assign n61720 = pi6013 & ~pi9040;
  assign n61721 = ~n61719 & ~n61720;
  assign n61722 = ~pi1731 & ~n61721;
  assign n61723 = pi1731 & n61721;
  assign n61724 = ~n61722 & ~n61723;
  assign n61725 = n61710 & ~n61724;
  assign n61726 = n61716 & n61725;
  assign n61727 = n61704 & n61726;
  assign n61728 = n61710 & n61724;
  assign n61729 = ~n61704 & n61728;
  assign n61730 = ~n61727 & ~n61729;
  assign n61731 = ~n61718 & n61730;
  assign n61732 = n61698 & ~n61731;
  assign n61733 = ~n61704 & ~n61716;
  assign n61734 = ~n61724 & n61733;
  assign n61735 = n61717 & ~n61724;
  assign n61736 = n61704 & n61735;
  assign n61737 = ~n61734 & ~n61736;
  assign n61738 = ~n61716 & n61725;
  assign n61739 = n61716 & n61728;
  assign n61740 = ~n61738 & ~n61739;
  assign n61741 = n61737 & n61740;
  assign n61742 = n61691 & ~n61741;
  assign n61743 = ~n61710 & n61724;
  assign n61744 = ~n61716 & n61743;
  assign n61745 = n61704 & n61744;
  assign n61746 = ~n61742 & ~n61745;
  assign n61747 = ~n61697 & ~n61746;
  assign n61748 = ~n61732 & ~n61747;
  assign n61749 = ~n61710 & ~n61724;
  assign n61750 = ~n61716 & n61749;
  assign n61751 = ~n61728 & ~n61749;
  assign n61752 = n61704 & ~n61751;
  assign n61753 = ~n61750 & ~n61752;
  assign n61754 = ~n61691 & ~n61753;
  assign n61755 = n61716 & n61743;
  assign n61756 = ~n61718 & ~n61755;
  assign n61757 = ~n61727 & n61756;
  assign n61758 = n61691 & ~n61757;
  assign n61759 = ~n61754 & ~n61758;
  assign n61760 = ~n61691 & ~n61704;
  assign n61761 = n61725 & n61760;
  assign n61762 = n61704 & n61750;
  assign n61763 = n61704 & n61724;
  assign n61764 = ~n61716 & n61763;
  assign n61765 = n61710 & n61764;
  assign n61766 = ~n61762 & ~n61765;
  assign n61767 = n61724 & n61733;
  assign n61768 = ~n61710 & n61767;
  assign n61769 = n61766 & ~n61768;
  assign n61770 = ~n61761 & n61769;
  assign n61771 = n61759 & n61770;
  assign n61772 = n61697 & ~n61771;
  assign n61773 = n61691 & ~n61704;
  assign n61774 = n61716 & n61773;
  assign n61775 = n61724 & n61774;
  assign n61776 = ~n61704 & n61738;
  assign n61777 = ~n61775 & ~n61776;
  assign n61778 = ~n61772 & n61777;
  assign n61779 = n61748 & n61778;
  assign n61780 = pi1760 & ~n61779;
  assign n61781 = ~pi1760 & n61777;
  assign n61782 = n61748 & n61781;
  assign n61783 = ~n61772 & n61782;
  assign po1854 = n61780 | n61783;
  assign n61785 = n61137 & n61169;
  assign n61786 = ~n61222 & ~n61785;
  assign n61787 = ~n61143 & ~n61786;
  assign n61788 = n61166 & n61218;
  assign n61789 = ~n61787 & ~n61788;
  assign n61790 = ~n61190 & n61789;
  assign n61791 = ~n61137 & n61174;
  assign n61792 = ~n61169 & ~n61791;
  assign n61793 = ~n61233 & n61792;
  assign n61794 = ~n61143 & ~n61793;
  assign n61795 = n61112 & n61794;
  assign n61796 = n61143 & n61231;
  assign n61797 = ~n61162 & ~n61188;
  assign n61798 = ~n61156 & n61797;
  assign n61799 = ~n61796 & n61798;
  assign n61800 = n61112 & ~n61799;
  assign n61801 = n61118 & n61143;
  assign n61802 = n61130 & n61801;
  assign n61803 = ~n61124 & n61802;
  assign n61804 = ~n61137 & n61199;
  assign n61805 = ~n61803 & ~n61804;
  assign n61806 = ~n61221 & n61805;
  assign n61807 = n61130 & n61160;
  assign n61808 = ~n61137 & n61148;
  assign n61809 = ~n61165 & ~n61808;
  assign n61810 = ~n61143 & ~n61809;
  assign n61811 = ~n61807 & ~n61810;
  assign n61812 = n61806 & n61811;
  assign n61813 = ~n61112 & ~n61812;
  assign n61814 = n61137 & n61803;
  assign n61815 = ~n61813 & ~n61814;
  assign n61816 = ~n61800 & n61815;
  assign n61817 = ~n61795 & n61816;
  assign n61818 = n61790 & n61817;
  assign n61819 = pi1780 & ~n61818;
  assign n61820 = ~pi1780 & n61790;
  assign n61821 = n61817 & n61820;
  assign po1855 = n61819 | n61821;
  assign n61823 = pi5949 & ~pi9040;
  assign n61824 = pi5822 & pi9040;
  assign n61825 = ~n61823 & ~n61824;
  assign n61826 = ~pi1757 & ~n61825;
  assign n61827 = pi1757 & n61825;
  assign n61828 = ~n61826 & ~n61827;
  assign n61829 = pi5838 & ~pi9040;
  assign n61830 = pi5829 & pi9040;
  assign n61831 = ~n61829 & ~n61830;
  assign n61832 = ~pi1745 & n61831;
  assign n61833 = pi1745 & ~n61831;
  assign n61834 = ~n61832 & ~n61833;
  assign n61835 = pi6076 & ~pi9040;
  assign n61836 = pi5815 & pi9040;
  assign n61837 = ~n61835 & ~n61836;
  assign n61838 = ~pi1751 & n61837;
  assign n61839 = pi1751 & ~n61837;
  assign n61840 = ~n61838 & ~n61839;
  assign n61841 = pi5819 & ~pi9040;
  assign n61842 = pi5937 & pi9040;
  assign n61843 = ~n61841 & ~n61842;
  assign n61844 = ~pi1723 & n61843;
  assign n61845 = pi1723 & ~n61843;
  assign n61846 = ~n61844 & ~n61845;
  assign n61847 = pi5817 & pi9040;
  assign n61848 = pi5815 & ~pi9040;
  assign n61849 = ~n61847 & ~n61848;
  assign n61850 = ~pi1746 & n61849;
  assign n61851 = pi1746 & ~n61849;
  assign n61852 = ~n61850 & ~n61851;
  assign n61853 = ~n61846 & n61852;
  assign n61854 = ~n61840 & n61853;
  assign n61855 = ~n61834 & n61854;
  assign n61856 = n61846 & n61852;
  assign n61857 = ~n61840 & n61856;
  assign n61858 = n61834 & n61857;
  assign n61859 = ~n61855 & ~n61858;
  assign n61860 = n61846 & ~n61852;
  assign n61861 = ~n61840 & n61860;
  assign n61862 = ~n61834 & n61861;
  assign n61863 = pi5820 & ~pi9040;
  assign n61864 = pi5948 & pi9040;
  assign n61865 = ~n61863 & ~n61864;
  assign n61866 = ~pi1740 & ~n61865;
  assign n61867 = pi1740 & n61865;
  assign n61868 = ~n61866 & ~n61867;
  assign n61869 = ~n61846 & ~n61852;
  assign n61870 = ~n61834 & n61869;
  assign n61871 = n61840 & n61860;
  assign n61872 = n61834 & n61871;
  assign n61873 = ~n61870 & ~n61872;
  assign n61874 = ~n61868 & ~n61873;
  assign n61875 = ~n61862 & ~n61874;
  assign n61876 = n61840 & n61856;
  assign n61877 = n61868 & n61876;
  assign n61878 = n61860 & n61868;
  assign n61879 = ~n61834 & n61878;
  assign n61880 = ~n61877 & ~n61879;
  assign n61881 = n61875 & n61880;
  assign n61882 = n61859 & n61881;
  assign n61883 = n61828 & ~n61882;
  assign n61884 = ~n61828 & ~n61868;
  assign n61885 = n61840 & n61852;
  assign n61886 = ~n61834 & n61840;
  assign n61887 = n61846 & n61886;
  assign n61888 = ~n61885 & ~n61887;
  assign n61889 = n61884 & ~n61888;
  assign n61890 = n61834 & ~n61840;
  assign n61891 = ~n61852 & n61890;
  assign n61892 = n61846 & n61891;
  assign n61893 = n61834 & ~n61846;
  assign n61894 = n61840 & n61893;
  assign n61895 = ~n61892 & ~n61894;
  assign n61896 = ~n61834 & n61868;
  assign n61897 = ~n61840 & n61896;
  assign n61898 = ~n61860 & n61897;
  assign n61899 = n61854 & n61868;
  assign n61900 = ~n61898 & ~n61899;
  assign n61901 = n61895 & n61900;
  assign n61902 = ~n61828 & ~n61901;
  assign n61903 = n61840 & n61853;
  assign n61904 = ~n61868 & n61903;
  assign n61905 = n61834 & n61904;
  assign n61906 = ~n61840 & n61869;
  assign n61907 = n61834 & n61906;
  assign n61908 = ~n61858 & ~n61907;
  assign n61909 = ~n61868 & ~n61908;
  assign n61910 = ~n61905 & ~n61909;
  assign n61911 = n61868 & n61892;
  assign n61912 = n61910 & ~n61911;
  assign n61913 = ~n61902 & n61912;
  assign n61914 = ~n61889 & n61913;
  assign n61915 = ~n61883 & n61914;
  assign n61916 = n61840 & n61869;
  assign n61917 = n61834 & n61868;
  assign n61918 = n61916 & n61917;
  assign n61919 = n61915 & ~n61918;
  assign n61920 = ~pi1772 & ~n61919;
  assign n61921 = n61914 & ~n61918;
  assign n61922 = pi1772 & n61921;
  assign n61923 = ~n61883 & n61922;
  assign po1856 = n61920 | n61923;
  assign n61925 = ~n61137 & n61245;
  assign n61926 = ~n61173 & ~n61231;
  assign n61927 = ~n61143 & ~n61926;
  assign n61928 = ~n61925 & ~n61927;
  assign n61929 = n61130 & n61220;
  assign n61930 = ~n61202 & ~n61929;
  assign n61931 = ~n61233 & n61930;
  assign n61932 = n61143 & ~n61931;
  assign n61933 = n61928 & ~n61932;
  assign n61934 = n61137 & n61166;
  assign n61935 = n61933 & ~n61934;
  assign n61936 = ~n61112 & ~n61935;
  assign n61937 = ~n61169 & ~n61174;
  assign n61938 = ~n61166 & ~n61233;
  assign n61939 = n61937 & n61938;
  assign n61940 = ~n61137 & ~n61939;
  assign n61941 = n61147 & ~n61926;
  assign n61942 = ~n61940 & ~n61941;
  assign n61943 = ~n61222 & n61942;
  assign n61944 = n61112 & ~n61943;
  assign n61945 = ~n61936 & ~n61944;
  assign n61946 = ~n61137 & n61231;
  assign n61947 = ~n61934 & ~n61946;
  assign n61948 = ~n61143 & ~n61947;
  assign n61949 = n61945 & ~n61948;
  assign n61950 = pi1769 & ~n61949;
  assign n61951 = ~pi1769 & ~n61948;
  assign n61952 = ~n61944 & n61951;
  assign n61953 = ~n61936 & n61952;
  assign po1858 = n61950 | n61953;
  assign n61955 = ~n61691 & n61750;
  assign n61956 = ~n61704 & n61955;
  assign n61957 = ~n61704 & n61726;
  assign n61958 = ~n61691 & n61957;
  assign n61959 = ~n61956 & ~n61958;
  assign n61960 = n61691 & n61768;
  assign n61961 = n61959 & ~n61960;
  assign n61962 = ~n61710 & n61773;
  assign n61963 = n61704 & n61717;
  assign n61964 = ~n61704 & n61710;
  assign n61965 = n61716 & n61964;
  assign n61966 = ~n61963 & ~n61965;
  assign n61967 = ~n61691 & ~n61966;
  assign n61968 = ~n61761 & ~n61967;
  assign n61969 = ~n61765 & ~n61957;
  assign n61970 = n61710 & ~n61716;
  assign n61971 = n61691 & n61704;
  assign n61972 = n61970 & n61971;
  assign n61973 = n61691 & n61744;
  assign n61974 = ~n61972 & ~n61973;
  assign n61975 = n61969 & n61974;
  assign n61976 = n61968 & n61975;
  assign n61977 = ~n61962 & n61976;
  assign n61978 = ~n61697 & ~n61977;
  assign n61979 = ~n61739 & ~n61963;
  assign n61980 = ~n61776 & n61979;
  assign n61981 = n61691 & ~n61980;
  assign n61982 = n61724 & n61970;
  assign n61983 = ~n61704 & n61982;
  assign n61984 = ~n61704 & n61755;
  assign n61985 = ~n61710 & ~n61716;
  assign n61986 = ~n61725 & ~n61985;
  assign n61987 = n61704 & ~n61986;
  assign n61988 = ~n61984 & ~n61987;
  assign n61989 = ~n61983 & n61988;
  assign n61990 = ~n61691 & ~n61989;
  assign n61991 = ~n61981 & ~n61990;
  assign n61992 = n61697 & ~n61991;
  assign n61993 = ~n61704 & n61735;
  assign n61994 = n61704 & n61728;
  assign n61995 = ~n61993 & ~n61994;
  assign n61996 = n61691 & ~n61995;
  assign n61997 = ~n61992 & ~n61996;
  assign n61998 = ~n61978 & n61997;
  assign n61999 = n61961 & n61998;
  assign n62000 = pi1783 & n61999;
  assign n62001 = ~pi1783 & ~n61999;
  assign po1861 = n62000 | n62001;
  assign n62003 = n61834 & n61876;
  assign n62004 = ~n61834 & n61903;
  assign n62005 = ~n62003 & ~n62004;
  assign n62006 = n61868 & ~n62005;
  assign n62007 = ~n61892 & ~n61899;
  assign n62008 = n61846 & n61890;
  assign n62009 = ~n61894 & ~n62008;
  assign n62010 = ~n61868 & ~n62009;
  assign n62011 = ~n61834 & ~n61868;
  assign n62012 = n61856 & n62011;
  assign n62013 = n61840 & n62012;
  assign n62014 = ~n61834 & ~n61840;
  assign n62015 = ~n61852 & n62014;
  assign n62016 = ~n61846 & n62015;
  assign n62017 = n61840 & n61868;
  assign n62018 = ~n61852 & n62017;
  assign n62019 = n61846 & n62018;
  assign n62020 = ~n62016 & ~n62019;
  assign n62021 = ~n62013 & n62020;
  assign n62022 = ~n62010 & n62021;
  assign n62023 = n62007 & n62022;
  assign n62024 = n61828 & ~n62023;
  assign n62025 = ~n61868 & n61892;
  assign n62026 = n61853 & n61917;
  assign n62027 = ~n61840 & n62026;
  assign n62028 = ~n62025 & ~n62027;
  assign n62029 = ~n62024 & n62028;
  assign n62030 = ~n62006 & n62029;
  assign n62031 = ~n61840 & n61846;
  assign n62032 = n61896 & n62031;
  assign n62033 = ~n61877 & ~n62032;
  assign n62034 = n61868 & n61906;
  assign n62035 = n61834 & n61916;
  assign n62036 = ~n62034 & ~n62035;
  assign n62037 = ~n61834 & n61853;
  assign n62038 = n61840 & ~n61852;
  assign n62039 = ~n62037 & ~n62038;
  assign n62040 = ~n61868 & ~n62039;
  assign n62041 = ~n61834 & n61857;
  assign n62042 = ~n62003 & ~n62041;
  assign n62043 = ~n62040 & n62042;
  assign n62044 = n62036 & n62043;
  assign n62045 = n62033 & n62044;
  assign n62046 = ~n61828 & ~n62045;
  assign n62047 = n62030 & ~n62046;
  assign n62048 = ~pi1766 & ~n62047;
  assign n62049 = pi1766 & n62030;
  assign n62050 = ~n62046 & n62049;
  assign po1862 = n62048 | n62050;
  assign n62052 = n61608 & n61636;
  assign n62053 = ~n61655 & ~n61664;
  assign n62054 = n61614 & ~n62053;
  assign n62055 = ~n62052 & ~n62054;
  assign n62056 = ~n61650 & n62055;
  assign n62057 = ~n61614 & n61653;
  assign n62058 = ~n61642 & ~n62057;
  assign n62059 = ~n61672 & n62058;
  assign n62060 = n62056 & n62059;
  assign n62061 = n61589 & ~n62060;
  assign n62062 = n61622 & n61629;
  assign n62063 = n61608 & n62062;
  assign n62064 = ~n61627 & ~n62063;
  assign n62065 = ~n61608 & n61671;
  assign n62066 = ~n61637 & ~n62065;
  assign n62067 = n61602 & n61622;
  assign n62068 = n61614 & n62067;
  assign n62069 = n61608 & n61641;
  assign n62070 = ~n62068 & ~n62069;
  assign n62071 = n61601 & ~n61622;
  assign n62072 = ~n61595 & n61608;
  assign n62073 = ~n62071 & ~n62072;
  assign n62074 = ~n61677 & n62073;
  assign n62075 = ~n61614 & ~n62074;
  assign n62076 = n62070 & ~n62075;
  assign n62077 = n62066 & n62076;
  assign n62078 = n62064 & n62077;
  assign n62079 = ~n61589 & ~n62078;
  assign n62080 = ~n62061 & ~n62079;
  assign n62081 = pi1774 & ~n62080;
  assign n62082 = ~pi1774 & ~n62061;
  assign n62083 = ~n62079 & n62082;
  assign po1863 = n62081 | n62083;
  assign n62085 = ~n61301 & n61559;
  assign n62086 = ~n61329 & ~n62085;
  assign n62087 = ~n61279 & n61550;
  assign n62088 = ~n61294 & ~n62087;
  assign n62089 = ~n61271 & ~n62088;
  assign n62090 = n61301 & n61318;
  assign n62091 = ~n61309 & ~n62090;
  assign n62092 = n61271 & ~n62091;
  assign n62093 = ~n62089 & ~n62092;
  assign n62094 = ~n61544 & n62093;
  assign n62095 = n62086 & n62094;
  assign n62096 = ~n61304 & ~n61317;
  assign n62097 = n62095 & n62096;
  assign n62098 = n61260 & ~n62097;
  assign n62099 = n61285 & n61550;
  assign n62100 = n61293 & n61301;
  assign n62101 = ~n62099 & ~n62100;
  assign n62102 = n61271 & ~n62101;
  assign n62103 = n61271 & n61318;
  assign n62104 = ~n61301 & n62103;
  assign n62105 = ~n62102 & ~n62104;
  assign n62106 = n61302 & n61323;
  assign n62107 = n61545 & ~n62106;
  assign n62108 = n61271 & ~n62107;
  assign n62109 = ~n61301 & n61540;
  assign n62110 = ~n62108 & ~n62109;
  assign n62111 = n62105 & n62110;
  assign n62112 = ~n61260 & ~n62111;
  assign n62113 = ~n61559 & ~n61564;
  assign n62114 = ~n61310 & n62113;
  assign n62115 = n61572 & ~n62114;
  assign n62116 = ~n62112 & ~n62115;
  assign n62117 = ~n61304 & ~n61544;
  assign n62118 = ~n61271 & ~n62117;
  assign n62119 = n62116 & ~n62118;
  assign n62120 = ~n62098 & n62119;
  assign n62121 = ~pi1778 & n62120;
  assign n62122 = pi1778 & ~n62120;
  assign po1864 = n62121 | n62122;
  assign n62124 = ~n62027 & ~n62032;
  assign n62125 = ~n61892 & ~n61903;
  assign n62126 = ~n62037 & n62125;
  assign n62127 = ~n61868 & ~n62126;
  assign n62128 = ~n61834 & n61871;
  assign n62129 = ~n62016 & ~n62128;
  assign n62130 = ~n61918 & n62129;
  assign n62131 = n61857 & n61868;
  assign n62132 = n62130 & ~n62131;
  assign n62133 = ~n62127 & n62132;
  assign n62134 = n61828 & ~n62133;
  assign n62135 = n61834 & n61878;
  assign n62136 = ~n61846 & n61886;
  assign n62137 = ~n61903 & ~n62136;
  assign n62138 = n61868 & ~n62137;
  assign n62139 = ~n62135 & ~n62138;
  assign n62140 = ~n61868 & n61869;
  assign n62141 = n61834 & n62140;
  assign n62142 = ~n61868 & n61876;
  assign n62143 = ~n62141 & ~n62142;
  assign n62144 = n62139 & n62143;
  assign n62145 = ~n61846 & n61890;
  assign n62146 = ~n62003 & ~n62145;
  assign n62147 = ~n62041 & n62146;
  assign n62148 = n62144 & n62147;
  assign n62149 = ~n61828 & ~n62148;
  assign n62150 = ~n62003 & n62129;
  assign n62151 = ~n61868 & ~n62150;
  assign n62152 = ~n62149 & ~n62151;
  assign n62153 = ~n62134 & n62152;
  assign n62154 = n62124 & n62153;
  assign n62155 = pi1773 & ~n62154;
  assign n62156 = ~pi1773 & n62154;
  assign po1865 = n62155 | n62156;
  assign n62158 = ~n61750 & ~n61755;
  assign n62159 = ~n61691 & ~n62158;
  assign n62160 = n61704 & n61739;
  assign n62161 = ~n62159 & ~n62160;
  assign n62162 = n61704 & n61710;
  assign n62163 = ~n61970 & ~n62162;
  assign n62164 = ~n61735 & n62163;
  assign n62165 = n61691 & ~n62164;
  assign n62166 = n62161 & ~n62165;
  assign n62167 = ~n61697 & ~n62166;
  assign n62168 = ~n61691 & n61983;
  assign n62169 = ~n61958 & ~n62168;
  assign n62170 = ~n61960 & n62169;
  assign n62171 = ~n61704 & n61716;
  assign n62172 = ~n61724 & n62171;
  assign n62173 = ~n61768 & ~n62172;
  assign n62174 = n61691 & n61965;
  assign n62175 = n61704 & n61755;
  assign n62176 = ~n61691 & n61970;
  assign n62177 = ~n62175 & ~n62176;
  assign n62178 = ~n61762 & n62177;
  assign n62179 = ~n62174 & n62178;
  assign n62180 = n62173 & n62179;
  assign n62181 = ~n61973 & n62180;
  assign n62182 = n61697 & ~n62181;
  assign n62183 = n62170 & ~n62182;
  assign n62184 = ~n62167 & n62183;
  assign n62185 = ~pi1762 & ~n62184;
  assign n62186 = ~n62167 & n62170;
  assign n62187 = pi1762 & n62186;
  assign n62188 = ~n62182 & n62187;
  assign po1866 = n62185 | n62188;
  assign n62190 = n61691 & n61728;
  assign n62191 = ~n61704 & n62190;
  assign n62192 = ~n61993 & ~n62191;
  assign n62193 = n61716 & n61763;
  assign n62194 = ~n61704 & ~n61710;
  assign n62195 = ~n62172 & ~n62194;
  assign n62196 = ~n61691 & ~n62195;
  assign n62197 = ~n62193 & ~n62196;
  assign n62198 = n62192 & n62197;
  assign n62199 = n61697 & ~n62198;
  assign n62200 = ~n61726 & ~n61765;
  assign n62201 = ~n61704 & n61743;
  assign n62202 = n62200 & ~n62201;
  assign n62203 = n61691 & ~n62202;
  assign n62204 = n61728 & n61760;
  assign n62205 = ~n61776 & ~n62204;
  assign n62206 = ~n62203 & n62205;
  assign n62207 = ~n61735 & ~n61745;
  assign n62208 = ~n61691 & ~n62207;
  assign n62209 = n62206 & ~n62208;
  assign n62210 = ~n61697 & ~n62209;
  assign n62211 = ~n62199 & ~n62210;
  assign n62212 = ~n61704 & n61749;
  assign n62213 = n61704 & ~n61740;
  assign n62214 = ~n62212 & ~n62213;
  assign n62215 = ~n61691 & ~n62214;
  assign n62216 = ~n61726 & n62158;
  assign n62217 = n61971 & ~n62216;
  assign n62218 = ~n62215 & ~n62217;
  assign n62219 = n62211 & n62218;
  assign n62220 = ~pi1767 & ~n62219;
  assign n62221 = ~n62210 & n62218;
  assign n62222 = pi1767 & n62221;
  assign n62223 = ~n62199 & n62222;
  assign po1869 = n62220 | n62223;
  assign n62225 = ~n61855 & ~n61887;
  assign n62226 = n61828 & ~n62225;
  assign n62227 = ~n61891 & ~n62008;
  assign n62228 = ~n61861 & n62227;
  assign n62229 = ~n61868 & ~n62228;
  assign n62230 = n61828 & n62229;
  assign n62231 = ~n62226 & ~n62230;
  assign n62232 = n61854 & n62011;
  assign n62233 = ~n62013 & ~n62232;
  assign n62234 = ~n61894 & ~n62038;
  assign n62235 = n61868 & ~n62234;
  assign n62236 = n61828 & n62235;
  assign n62237 = n62233 & ~n62236;
  assign n62238 = n61834 & n61854;
  assign n62239 = n61834 & n61856;
  assign n62240 = ~n62004 & ~n62239;
  assign n62241 = n61868 & ~n62240;
  assign n62242 = ~n61892 & ~n62016;
  assign n62243 = n61834 & n61853;
  assign n62244 = ~n61916 & ~n62243;
  assign n62245 = ~n61868 & ~n62244;
  assign n62246 = n62242 & ~n62245;
  assign n62247 = ~n62241 & n62246;
  assign n62248 = ~n62238 & n62247;
  assign n62249 = ~n61828 & ~n62248;
  assign n62250 = ~n62041 & n62129;
  assign n62251 = n61868 & ~n62250;
  assign n62252 = ~n62249 & ~n62251;
  assign n62253 = n62237 & n62252;
  assign n62254 = n62231 & n62253;
  assign n62255 = ~pi1784 & ~n62254;
  assign n62256 = pi1784 & n62237;
  assign n62257 = n62231 & n62256;
  assign n62258 = n62252 & n62257;
  assign po1870 = n62255 | n62258;
  assign n62260 = ~n61039 & n61069;
  assign n62261 = n61039 & n61080;
  assign n62262 = ~n61066 & ~n62261;
  assign n62263 = ~n61013 & ~n62262;
  assign n62264 = ~n62260 & ~n62263;
  assign n62265 = n61013 & ~n61039;
  assign n62266 = ~n61031 & n62265;
  assign n62267 = n61025 & n62266;
  assign n62268 = n61048 & n61081;
  assign n62269 = ~n62267 & ~n62268;
  assign n62270 = n61013 & n61088;
  assign n62271 = n62269 & ~n62270;
  assign n62272 = ~n61043 & ~n61056;
  assign n62273 = n61031 & n61046;
  assign n62274 = n62272 & ~n62273;
  assign n62275 = n62271 & n62274;
  assign n62276 = n62264 & n62275;
  assign n62277 = ~n61078 & ~n62276;
  assign n62278 = ~n61019 & n61045;
  assign n62279 = ~n61066 & ~n62278;
  assign n62280 = n61039 & ~n62279;
  assign n62281 = n61025 & n61041;
  assign n62282 = ~n61093 & ~n62281;
  assign n62283 = n61019 & ~n61031;
  assign n62284 = n61039 & n62283;
  assign n62285 = n62282 & ~n62284;
  assign n62286 = ~n61013 & ~n62285;
  assign n62287 = ~n61039 & n61054;
  assign n62288 = ~n61019 & n61039;
  assign n62289 = ~n61031 & n62288;
  assign n62290 = n61025 & n62289;
  assign n62291 = ~n62287 & ~n62290;
  assign n62292 = n61013 & ~n62291;
  assign n62293 = ~n61039 & n61049;
  assign n62294 = ~n62292 & ~n62293;
  assign n62295 = ~n62286 & n62294;
  assign n62296 = ~n62280 & n62295;
  assign n62297 = n61078 & ~n62296;
  assign n62298 = ~n61013 & n61042;
  assign n62299 = ~n62297 & ~n62298;
  assign n62300 = n61061 & n62265;
  assign n62301 = ~n61031 & n62300;
  assign n62302 = n62299 & ~n62301;
  assign n62303 = ~n62277 & n62302;
  assign n62304 = ~pi1793 & ~n62303;
  assign n62305 = pi1793 & n62299;
  assign n62306 = ~n62277 & n62305;
  assign n62307 = ~n62301 & n62306;
  assign po1871 = n62304 | n62307;
  assign n62309 = ~n61040 & ~n61047;
  assign n62310 = n61013 & ~n62309;
  assign n62311 = ~n61100 & ~n62310;
  assign n62312 = ~n61019 & ~n61025;
  assign n62313 = ~n61013 & n62312;
  assign n62314 = n61039 & n62313;
  assign n62315 = n61039 & n61054;
  assign n62316 = ~n62312 & ~n62315;
  assign n62317 = n61019 & ~n61039;
  assign n62318 = n61025 & n62317;
  assign n62319 = n62316 & ~n62318;
  assign n62320 = ~n61013 & ~n62319;
  assign n62321 = ~n61050 & ~n62320;
  assign n62322 = ~n61078 & ~n62321;
  assign n62323 = n61013 & n61032;
  assign n62324 = n61039 & n62323;
  assign n62325 = ~n62270 & ~n62324;
  assign n62326 = ~n61078 & ~n62325;
  assign n62327 = ~n62322 & ~n62326;
  assign n62328 = ~n62314 & n62327;
  assign n62329 = ~n61042 & ~n61066;
  assign n62330 = ~n61093 & n62329;
  assign n62331 = n61013 & ~n62330;
  assign n62332 = ~n61039 & n61088;
  assign n62333 = ~n61069 & ~n62332;
  assign n62334 = ~n61013 & ~n62333;
  assign n62335 = ~n62281 & ~n62334;
  assign n62336 = ~n62331 & n62335;
  assign n62337 = ~n61056 & ~n61094;
  assign n62338 = n62336 & n62337;
  assign n62339 = n61078 & ~n62338;
  assign n62340 = n62328 & ~n62339;
  assign n62341 = n62311 & n62340;
  assign n62342 = ~pi1810 & ~n62341;
  assign n62343 = pi1810 & n62328;
  assign n62344 = n62311 & n62343;
  assign n62345 = ~n62339 & n62344;
  assign po1872 = n62342 | n62345;
  assign n62347 = ~n61393 & ~n61482;
  assign n62348 = ~n61462 & n62347;
  assign n62349 = n61400 & ~n62348;
  assign n62350 = ~n61412 & ~n61439;
  assign n62351 = ~n61409 & ~n61470;
  assign n62352 = ~n61383 & ~n61475;
  assign n62353 = ~n61400 & ~n62352;
  assign n62354 = ~n61449 & ~n62353;
  assign n62355 = n62351 & n62354;
  assign n62356 = n61357 & ~n62355;
  assign n62357 = ~n61369 & n61381;
  assign n62358 = ~n61500 & ~n62357;
  assign n62359 = ~n61363 & ~n62358;
  assign n62360 = ~n61418 & ~n61422;
  assign n62361 = ~n61400 & ~n62360;
  assign n62362 = ~n61363 & n61381;
  assign n62363 = ~n61390 & ~n62362;
  assign n62364 = ~n61382 & n62363;
  assign n62365 = n61400 & ~n62364;
  assign n62366 = ~n62361 & ~n62365;
  assign n62367 = ~n62359 & n62366;
  assign n62368 = ~n61357 & ~n62367;
  assign n62369 = ~n62356 & ~n62368;
  assign n62370 = n62350 & n62369;
  assign n62371 = ~n62349 & n62370;
  assign n62372 = ~pi1795 & ~n62371;
  assign n62373 = pi1795 & n62350;
  assign n62374 = ~n62349 & n62373;
  assign n62375 = n62369 & n62374;
  assign po1873 = n62372 | n62375;
  assign n62377 = ~n61608 & n61629;
  assign n62378 = ~n62065 & ~n62377;
  assign n62379 = n61614 & n62378;
  assign n62380 = n61608 & n61666;
  assign n62381 = ~n61602 & ~n61623;
  assign n62382 = ~n61622 & ~n62381;
  assign n62383 = n61595 & n61648;
  assign n62384 = n61608 & n61623;
  assign n62385 = ~n62383 & ~n62384;
  assign n62386 = ~n62382 & n62385;
  assign n62387 = ~n62380 & n62386;
  assign n62388 = ~n61614 & n62387;
  assign n62389 = ~n62379 & ~n62388;
  assign n62390 = n61608 & n62382;
  assign n62391 = ~n62063 & ~n62390;
  assign n62392 = ~n62389 & n62391;
  assign n62393 = n61589 & ~n62392;
  assign n62394 = n61614 & ~n62381;
  assign n62395 = ~n61608 & n62394;
  assign n62396 = ~n61643 & ~n61670;
  assign n62397 = n61608 & ~n62396;
  assign n62398 = n61614 & n62397;
  assign n62399 = n61622 & n62394;
  assign n62400 = ~n62398 & ~n62399;
  assign n62401 = ~n62395 & n62400;
  assign n62402 = ~n61589 & ~n62401;
  assign n62403 = ~n62393 & ~n62402;
  assign n62404 = ~n61614 & ~n62378;
  assign n62405 = ~n61627 & ~n62404;
  assign n62406 = ~n61589 & ~n62405;
  assign n62407 = n61614 & n61627;
  assign n62408 = ~n61614 & ~n62391;
  assign n62409 = ~n62407 & ~n62408;
  assign n62410 = ~n62406 & n62409;
  assign n62411 = n62403 & n62410;
  assign n62412 = pi1789 & ~n62411;
  assign n62413 = ~n62393 & n62410;
  assign n62414 = ~n62402 & n62413;
  assign n62415 = ~pi1789 & n62414;
  assign po1874 = n62412 | n62415;
  assign n62417 = n61608 & n62067;
  assign n62418 = n61614 & n62417;
  assign n62419 = n61648 & ~n62381;
  assign n62420 = ~n61671 & ~n62419;
  assign n62421 = ~n62063 & n62420;
  assign n62422 = ~n61614 & ~n62421;
  assign n62423 = n61608 & n61624;
  assign n62424 = ~n62422 & ~n62423;
  assign n62425 = n61622 & n61670;
  assign n62426 = ~n61608 & n62071;
  assign n62427 = ~n62425 & ~n62426;
  assign n62428 = ~n62384 & n62427;
  assign n62429 = n61614 & ~n62428;
  assign n62430 = n62424 & ~n62429;
  assign n62431 = n61589 & ~n62430;
  assign n62432 = ~n62418 & ~n62431;
  assign n62433 = ~n61608 & n61623;
  assign n62434 = ~n62062 & ~n62433;
  assign n62435 = n61614 & ~n62434;
  assign n62436 = ~n61672 & ~n62435;
  assign n62437 = ~n61644 & ~n62417;
  assign n62438 = ~n61608 & n61624;
  assign n62439 = n61608 & n61677;
  assign n62440 = ~n62071 & ~n62439;
  assign n62441 = ~n62425 & n62440;
  assign n62442 = ~n61614 & ~n62441;
  assign n62443 = ~n62438 & ~n62442;
  assign n62444 = n62437 & n62443;
  assign n62445 = n62436 & n62444;
  assign n62446 = ~n61589 & ~n62445;
  assign n62447 = ~n61658 & ~n62380;
  assign n62448 = ~n61614 & ~n62447;
  assign n62449 = ~n62446 & ~n62448;
  assign n62450 = n62432 & n62449;
  assign n62451 = pi1788 & n62450;
  assign n62452 = ~pi1788 & ~n62450;
  assign po1875 = n62451 | n62452;
  assign n62454 = pi5827 & ~pi9040;
  assign n62455 = pi6076 & pi9040;
  assign n62456 = ~n62454 & ~n62455;
  assign n62457 = ~pi1750 & n62456;
  assign n62458 = pi1750 & ~n62456;
  assign n62459 = ~n62457 & ~n62458;
  assign n62460 = pi5838 & pi9040;
  assign n62461 = pi5922 & ~pi9040;
  assign n62462 = ~n62460 & ~n62461;
  assign n62463 = ~pi1739 & n62462;
  assign n62464 = pi1739 & ~n62462;
  assign n62465 = ~n62463 & ~n62464;
  assign n62466 = pi5828 & pi9040;
  assign n62467 = pi5911 & ~pi9040;
  assign n62468 = ~n62466 & ~n62467;
  assign n62469 = ~pi1743 & n62468;
  assign n62470 = pi1743 & ~n62468;
  assign n62471 = ~n62469 & ~n62470;
  assign n62472 = pi5833 & ~pi9040;
  assign n62473 = pi5918 & pi9040;
  assign n62474 = ~n62472 & ~n62473;
  assign n62475 = ~pi1755 & n62474;
  assign n62476 = pi1755 & ~n62474;
  assign n62477 = ~n62475 & ~n62476;
  assign n62478 = ~n62471 & n62477;
  assign n62479 = n62465 & n62478;
  assign n62480 = ~n62459 & n62479;
  assign n62481 = pi5917 & pi9040;
  assign n62482 = pi5836 & ~pi9040;
  assign n62483 = ~n62481 & ~n62482;
  assign n62484 = ~pi1723 & ~n62483;
  assign n62485 = pi1723 & n62483;
  assign n62486 = ~n62484 & ~n62485;
  assign n62487 = pi5822 & ~pi9040;
  assign n62488 = pi5946 & pi9040;
  assign n62489 = ~n62487 & ~n62488;
  assign n62490 = ~pi1751 & ~n62489;
  assign n62491 = pi1751 & n62489;
  assign n62492 = ~n62490 & ~n62491;
  assign n62493 = ~n62471 & n62492;
  assign n62494 = ~n62477 & n62493;
  assign n62495 = n62471 & n62492;
  assign n62496 = n62477 & n62495;
  assign n62497 = n62471 & ~n62492;
  assign n62498 = n62459 & n62497;
  assign n62499 = ~n62496 & ~n62498;
  assign n62500 = ~n62494 & n62499;
  assign n62501 = n62465 & ~n62500;
  assign n62502 = ~n62477 & n62495;
  assign n62503 = n62477 & n62493;
  assign n62504 = ~n62502 & ~n62503;
  assign n62505 = ~n62465 & ~n62504;
  assign n62506 = ~n62501 & ~n62505;
  assign n62507 = ~n62471 & ~n62492;
  assign n62508 = ~n62477 & n62507;
  assign n62509 = ~n62465 & n62508;
  assign n62510 = n62477 & n62498;
  assign n62511 = ~n62509 & ~n62510;
  assign n62512 = n62506 & n62511;
  assign n62513 = ~n62486 & ~n62512;
  assign n62514 = ~n62459 & n62502;
  assign n62515 = n62459 & n62507;
  assign n62516 = ~n62459 & n62497;
  assign n62517 = ~n62515 & ~n62516;
  assign n62518 = n62465 & ~n62517;
  assign n62519 = ~n62514 & ~n62518;
  assign n62520 = ~n62477 & n62497;
  assign n62521 = ~n62465 & n62520;
  assign n62522 = n62477 & n62507;
  assign n62523 = ~n62494 & ~n62522;
  assign n62524 = ~n62521 & n62523;
  assign n62525 = ~n62496 & n62524;
  assign n62526 = n62459 & ~n62525;
  assign n62527 = n62519 & ~n62526;
  assign n62528 = n62486 & ~n62527;
  assign n62529 = ~n62513 & ~n62528;
  assign n62530 = ~n62480 & n62529;
  assign n62531 = ~n62459 & n62508;
  assign n62532 = n62477 & n62516;
  assign n62533 = ~n62531 & ~n62532;
  assign n62534 = ~n62465 & ~n62533;
  assign n62535 = n62530 & ~n62534;
  assign n62536 = ~pi1777 & ~n62535;
  assign n62537 = n62529 & ~n62534;
  assign n62538 = pi1777 & n62537;
  assign n62539 = ~n62480 & n62538;
  assign po1876 = n62536 | n62539;
  assign n62541 = n61293 & ~n61301;
  assign n62542 = ~n61556 & ~n62541;
  assign n62543 = ~n61271 & ~n62542;
  assign n62544 = n61271 & ~n61331;
  assign n62545 = ~n61342 & ~n62544;
  assign n62546 = ~n62543 & n62545;
  assign n62547 = n61260 & ~n62546;
  assign n62548 = ~n61271 & n61540;
  assign n62549 = ~n62547 & ~n62548;
  assign n62550 = ~n62085 & ~n62100;
  assign n62551 = n61271 & ~n62550;
  assign n62552 = n61271 & n61557;
  assign n62553 = n61294 & n61301;
  assign n62554 = n61273 & ~n61292;
  assign n62555 = ~n61308 & ~n62554;
  assign n62556 = ~n61285 & ~n62555;
  assign n62557 = ~n61309 & ~n62556;
  assign n62558 = ~n61544 & n62557;
  assign n62559 = ~n62553 & n62558;
  assign n62560 = ~n62552 & n62559;
  assign n62561 = ~n61260 & ~n62560;
  assign n62562 = ~n62551 & ~n62561;
  assign n62563 = n62549 & n62562;
  assign n62564 = pi1796 & ~n62563;
  assign n62565 = ~pi1796 & n62563;
  assign po1877 = n62564 | n62565;
  assign n62567 = ~n61094 & ~n62293;
  assign n62568 = ~n61013 & ~n62567;
  assign n62569 = ~n61078 & n61080;
  assign n62570 = n61013 & n62569;
  assign n62571 = ~n61025 & n62317;
  assign n62572 = ~n62283 & ~n62571;
  assign n62573 = ~n61049 & n62572;
  assign n62574 = ~n61013 & ~n62573;
  assign n62575 = ~n61039 & n61055;
  assign n62576 = ~n62574 & ~n62575;
  assign n62577 = ~n61078 & ~n62576;
  assign n62578 = ~n62570 & ~n62577;
  assign n62579 = ~n61043 & ~n61047;
  assign n62580 = ~n61039 & n61093;
  assign n62581 = ~n62261 & ~n62580;
  assign n62582 = n62579 & n62581;
  assign n62583 = n61013 & ~n62582;
  assign n62584 = ~n61019 & n61025;
  assign n62585 = n61013 & n62584;
  assign n62586 = n61039 & n62585;
  assign n62587 = ~n61039 & n62283;
  assign n62588 = ~n61047 & ~n62587;
  assign n62589 = ~n62290 & n62588;
  assign n62590 = ~n62586 & n62589;
  assign n62591 = ~n61013 & n62278;
  assign n62592 = n62590 & ~n62591;
  assign n62593 = n61078 & ~n62592;
  assign n62594 = ~n62583 & ~n62593;
  assign n62595 = n62578 & n62594;
  assign n62596 = ~n62568 & n62595;
  assign n62597 = pi1814 & n62596;
  assign n62598 = ~pi1814 & ~n62596;
  assign po1878 = n62597 | n62598;
  assign n62600 = ~n62465 & n62502;
  assign n62601 = n62459 & n62600;
  assign n62602 = n62459 & ~n62465;
  assign n62603 = n62507 & n62602;
  assign n62604 = n62477 & n62603;
  assign n62605 = ~n62601 & ~n62604;
  assign n62606 = n62465 & n62496;
  assign n62607 = n62459 & n62606;
  assign n62608 = n62459 & n62477;
  assign n62609 = ~n62492 & n62608;
  assign n62610 = ~n62471 & n62609;
  assign n62611 = ~n62607 & ~n62610;
  assign n62612 = ~n62493 & ~n62497;
  assign n62613 = n62465 & ~n62608;
  assign n62614 = ~n62612 & n62613;
  assign n62615 = ~n62471 & ~n62477;
  assign n62616 = ~n62459 & n62615;
  assign n62617 = ~n62459 & n62495;
  assign n62618 = ~n62616 & ~n62617;
  assign n62619 = ~n62465 & ~n62618;
  assign n62620 = n62459 & ~n62495;
  assign n62621 = ~n62465 & n62620;
  assign n62622 = n62477 & n62621;
  assign n62623 = ~n62619 & ~n62622;
  assign n62624 = ~n62614 & n62623;
  assign n62625 = n62611 & n62624;
  assign n62626 = n62486 & ~n62625;
  assign n62627 = n62605 & ~n62626;
  assign n62628 = n62465 & n62494;
  assign n62629 = ~n62459 & n62628;
  assign n62630 = n62465 & ~n62486;
  assign n62631 = ~n62508 & ~n62617;
  assign n62632 = n62608 & ~n62612;
  assign n62633 = n62631 & ~n62632;
  assign n62634 = n62630 & ~n62633;
  assign n62635 = ~n62459 & n62522;
  assign n62636 = n62459 & n62495;
  assign n62637 = ~n62520 & ~n62636;
  assign n62638 = ~n62459 & ~n62471;
  assign n62639 = n62477 & n62638;
  assign n62640 = ~n62516 & ~n62639;
  assign n62641 = n62637 & n62640;
  assign n62642 = ~n62465 & ~n62641;
  assign n62643 = ~n62635 & ~n62642;
  assign n62644 = ~n62486 & ~n62643;
  assign n62645 = ~n62634 & ~n62644;
  assign n62646 = ~n62629 & n62645;
  assign n62647 = n62627 & n62646;
  assign n62648 = pi1782 & ~n62647;
  assign n62649 = ~pi1782 & n62627;
  assign n62650 = n62646 & n62649;
  assign po1879 = n62648 | n62650;
  assign n62652 = ~n62516 & ~n62636;
  assign n62653 = ~n62465 & ~n62652;
  assign n62654 = ~n62604 & ~n62653;
  assign n62655 = n62486 & ~n62654;
  assign n62656 = ~n62478 & ~n62493;
  assign n62657 = n62459 & ~n62656;
  assign n62658 = ~n62502 & ~n62657;
  assign n62659 = n62465 & ~n62658;
  assign n62660 = ~n62632 & ~n62659;
  assign n62661 = ~n62459 & n62496;
  assign n62662 = n62459 & ~n62477;
  assign n62663 = ~n62492 & n62662;
  assign n62664 = ~n62459 & ~n62656;
  assign n62665 = ~n62663 & ~n62664;
  assign n62666 = ~n62465 & ~n62665;
  assign n62667 = ~n62661 & ~n62666;
  assign n62668 = n62660 & n62667;
  assign n62669 = ~n62486 & ~n62668;
  assign n62670 = ~n62459 & ~n62477;
  assign n62671 = ~n62493 & n62670;
  assign n62672 = n62486 & n62671;
  assign n62673 = ~n62459 & n62477;
  assign n62674 = n62493 & n62673;
  assign n62675 = ~n62465 & n62674;
  assign n62676 = ~n62459 & n62465;
  assign n62677 = ~n62477 & n62676;
  assign n62678 = ~n62492 & n62677;
  assign n62679 = ~n62675 & ~n62678;
  assign n62680 = ~n62672 & n62679;
  assign n62681 = ~n62520 & ~n62638;
  assign n62682 = n62465 & n62486;
  assign n62683 = ~n62681 & n62682;
  assign n62684 = n62680 & ~n62683;
  assign n62685 = ~n62669 & n62684;
  assign n62686 = ~n62655 & n62685;
  assign n62687 = pi1790 & ~n62686;
  assign n62688 = ~pi1790 & n62686;
  assign po1880 = n62687 | n62688;
  assign n62690 = n62492 & n62662;
  assign n62691 = n62523 & ~n62690;
  assign n62692 = n62682 & ~n62691;
  assign n62693 = n62486 & n62520;
  assign n62694 = ~n62459 & n62693;
  assign n62695 = n62477 & n62492;
  assign n62696 = ~n62617 & ~n62695;
  assign n62697 = ~n62465 & ~n62696;
  assign n62698 = ~n62509 & ~n62697;
  assign n62699 = n62486 & ~n62698;
  assign n62700 = ~n62694 & ~n62699;
  assign n62701 = n62492 & n62673;
  assign n62702 = ~n62510 & ~n62701;
  assign n62703 = ~n62465 & ~n62702;
  assign n62704 = n62700 & ~n62703;
  assign n62705 = n62495 & n62676;
  assign n62706 = ~n62477 & n62705;
  assign n62707 = ~n62612 & n62673;
  assign n62708 = ~n62706 & ~n62707;
  assign n62709 = ~n62531 & n62708;
  assign n62710 = ~n62612 & n62662;
  assign n62711 = ~n62610 & ~n62710;
  assign n62712 = ~n62477 & n62602;
  assign n62713 = n62471 & n62712;
  assign n62714 = ~n62607 & ~n62713;
  assign n62715 = n62711 & n62714;
  assign n62716 = n62709 & n62715;
  assign n62717 = ~n62486 & ~n62716;
  assign n62718 = n62704 & ~n62717;
  assign n62719 = ~n62692 & n62718;
  assign n62720 = ~pi1781 & ~n62719;
  assign n62721 = pi1781 & n62704;
  assign n62722 = ~n62692 & n62721;
  assign n62723 = ~n62717 & n62722;
  assign po1881 = n62720 | n62723;
  assign n62725 = pi6063 & pi9040;
  assign n62726 = pi6150 & ~pi9040;
  assign n62727 = ~n62725 & ~n62726;
  assign n62728 = ~pi1791 & ~n62727;
  assign n62729 = pi1791 & n62727;
  assign n62730 = ~n62728 & ~n62729;
  assign n62731 = pi6031 & pi9040;
  assign n62732 = pi6050 & ~pi9040;
  assign n62733 = ~n62731 & ~n62732;
  assign n62734 = ~pi1775 & ~n62733;
  assign n62735 = pi1775 & n62733;
  assign n62736 = ~n62734 & ~n62735;
  assign n62737 = pi6168 & ~pi9040;
  assign n62738 = pi6058 & pi9040;
  assign n62739 = ~n62737 & ~n62738;
  assign n62740 = ~pi1815 & n62739;
  assign n62741 = pi1815 & ~n62739;
  assign n62742 = ~n62740 & ~n62741;
  assign n62743 = pi6257 & pi9040;
  assign n62744 = pi6233 & ~pi9040;
  assign n62745 = ~n62743 & ~n62744;
  assign n62746 = ~pi1803 & ~n62745;
  assign n62747 = pi1803 & n62745;
  assign n62748 = ~n62746 & ~n62747;
  assign n62749 = ~n62742 & n62748;
  assign n62750 = ~n62736 & n62749;
  assign n62751 = pi6027 & ~pi9040;
  assign n62752 = pi6152 & pi9040;
  assign n62753 = ~n62751 & ~n62752;
  assign n62754 = pi1817 & n62753;
  assign n62755 = ~pi1817 & ~n62753;
  assign n62756 = ~n62754 & ~n62755;
  assign n62757 = n62750 & ~n62756;
  assign n62758 = n62742 & ~n62748;
  assign n62759 = ~n62736 & n62758;
  assign n62760 = ~n62756 & n62759;
  assign n62761 = ~n62757 & ~n62760;
  assign n62762 = n62736 & n62758;
  assign n62763 = n62756 & n62762;
  assign n62764 = ~n62742 & ~n62748;
  assign n62765 = ~n62736 & n62764;
  assign n62766 = n62756 & n62765;
  assign n62767 = ~n62763 & ~n62766;
  assign n62768 = n62761 & n62767;
  assign n62769 = n62730 & ~n62768;
  assign n62770 = ~n62736 & n62756;
  assign n62771 = n62748 & n62770;
  assign n62772 = n62742 & n62771;
  assign n62773 = ~n62765 & ~n62772;
  assign n62774 = n62730 & ~n62773;
  assign n62775 = ~n62730 & n62748;
  assign n62776 = ~n62756 & n62775;
  assign n62777 = n62736 & ~n62742;
  assign n62778 = n62756 & n62758;
  assign n62779 = ~n62777 & ~n62778;
  assign n62780 = ~n62730 & ~n62779;
  assign n62781 = ~n62776 & ~n62780;
  assign n62782 = n62742 & n62748;
  assign n62783 = n62736 & n62782;
  assign n62784 = ~n62756 & n62783;
  assign n62785 = n62781 & ~n62784;
  assign n62786 = n62748 & n62777;
  assign n62787 = n62756 & n62786;
  assign n62788 = n62785 & ~n62787;
  assign n62789 = ~n62774 & n62788;
  assign n62790 = pi6148 & pi9040;
  assign n62791 = pi6083 & ~pi9040;
  assign n62792 = ~n62790 & ~n62791;
  assign n62793 = ~pi1820 & ~n62792;
  assign n62794 = pi1820 & n62792;
  assign n62795 = ~n62793 & ~n62794;
  assign n62796 = ~n62789 & ~n62795;
  assign n62797 = ~n62736 & n62748;
  assign n62798 = ~n62730 & n62756;
  assign n62799 = n62795 & n62798;
  assign n62800 = n62797 & n62799;
  assign n62801 = ~n62736 & ~n62756;
  assign n62802 = ~n62748 & n62801;
  assign n62803 = ~n62730 & ~n62802;
  assign n62804 = n62736 & n62756;
  assign n62805 = n62742 & n62804;
  assign n62806 = ~n62749 & ~n62797;
  assign n62807 = ~n62756 & ~n62806;
  assign n62808 = n62730 & ~n62762;
  assign n62809 = ~n62807 & n62808;
  assign n62810 = ~n62805 & n62809;
  assign n62811 = ~n62803 & ~n62810;
  assign n62812 = n62736 & n62764;
  assign n62813 = n62756 & n62812;
  assign n62814 = ~n62811 & ~n62813;
  assign n62815 = n62795 & ~n62814;
  assign n62816 = ~n62800 & ~n62815;
  assign n62817 = ~n62796 & n62816;
  assign n62818 = ~n62769 & n62817;
  assign n62819 = ~n62730 & n62784;
  assign n62820 = n62818 & ~n62819;
  assign n62821 = pi1824 & ~n62820;
  assign n62822 = ~pi1824 & ~n62819;
  assign n62823 = n62817 & n62822;
  assign n62824 = ~n62769 & n62823;
  assign po1888 = n62821 | n62824;
  assign n62826 = pi6049 & ~pi9040;
  assign n62827 = pi6061 & pi9040;
  assign n62828 = ~n62826 & ~n62827;
  assign n62829 = ~pi1803 & ~n62828;
  assign n62830 = pi1803 & n62828;
  assign n62831 = ~n62829 & ~n62830;
  assign n62832 = pi6225 & ~pi9040;
  assign n62833 = pi6026 & pi9040;
  assign n62834 = ~n62832 & ~n62833;
  assign n62835 = ~pi1813 & n62834;
  assign n62836 = pi1813 & ~n62834;
  assign n62837 = ~n62835 & ~n62836;
  assign n62838 = pi6061 & ~pi9040;
  assign n62839 = pi6225 & pi9040;
  assign n62840 = ~n62838 & ~n62839;
  assign n62841 = pi1775 & n62840;
  assign n62842 = ~pi1775 & ~n62840;
  assign n62843 = ~n62841 & ~n62842;
  assign n62844 = n62837 & n62843;
  assign n62845 = pi6174 & ~pi9040;
  assign n62846 = pi6175 & pi9040;
  assign n62847 = ~n62845 & ~n62846;
  assign n62848 = pi1802 & n62847;
  assign n62849 = ~pi1802 & ~n62847;
  assign n62850 = ~n62848 & ~n62849;
  assign n62851 = pi6133 & pi9040;
  assign n62852 = pi6066 & ~pi9040;
  assign n62853 = ~n62851 & ~n62852;
  assign n62854 = pi1819 & n62853;
  assign n62855 = ~pi1819 & ~n62853;
  assign n62856 = ~n62854 & ~n62855;
  assign n62857 = ~n62850 & ~n62856;
  assign n62858 = n62844 & n62857;
  assign n62859 = pi6056 & ~pi9040;
  assign n62860 = pi6153 & pi9040;
  assign n62861 = ~n62859 & ~n62860;
  assign n62862 = ~pi1787 & n62861;
  assign n62863 = pi1787 & ~n62861;
  assign n62864 = ~n62862 & ~n62863;
  assign n62865 = ~n62837 & n62864;
  assign n62866 = ~n62850 & n62856;
  assign n62867 = n62865 & n62866;
  assign n62868 = ~n62837 & ~n62843;
  assign n62869 = ~n62864 & n62868;
  assign n62870 = n62850 & n62864;
  assign n62871 = ~n62843 & n62870;
  assign n62872 = n62837 & n62871;
  assign n62873 = ~n62869 & ~n62872;
  assign n62874 = ~n62837 & n62843;
  assign n62875 = n62850 & n62874;
  assign n62876 = n62873 & ~n62875;
  assign n62877 = ~n62856 & ~n62876;
  assign n62878 = n62864 & n62868;
  assign n62879 = ~n62850 & n62878;
  assign n62880 = ~n62877 & ~n62879;
  assign n62881 = ~n62867 & n62880;
  assign n62882 = ~n62858 & n62881;
  assign n62883 = n62844 & ~n62864;
  assign n62884 = ~n62850 & n62883;
  assign n62885 = ~n62864 & n62874;
  assign n62886 = n62850 & n62885;
  assign n62887 = ~n62884 & ~n62886;
  assign n62888 = n62882 & n62887;
  assign n62889 = ~n62831 & ~n62888;
  assign n62890 = ~n62850 & n62864;
  assign n62891 = n62843 & n62890;
  assign n62892 = ~n62837 & n62891;
  assign n62893 = ~n62883 & ~n62892;
  assign n62894 = ~n62856 & ~n62893;
  assign n62895 = ~n62837 & n62870;
  assign n62896 = ~n62850 & n62885;
  assign n62897 = ~n62895 & ~n62896;
  assign n62898 = n62856 & ~n62897;
  assign n62899 = n62844 & n62870;
  assign n62900 = ~n62843 & n62890;
  assign n62901 = n62837 & n62900;
  assign n62902 = ~n62899 & ~n62901;
  assign n62903 = ~n62898 & n62902;
  assign n62904 = ~n62894 & n62903;
  assign n62905 = n62831 & ~n62904;
  assign n62906 = ~n62837 & ~n62864;
  assign n62907 = n62850 & n62906;
  assign n62908 = n62837 & ~n62864;
  assign n62909 = ~n62850 & n62908;
  assign n62910 = ~n62907 & ~n62909;
  assign n62911 = ~n62856 & ~n62910;
  assign n62912 = n62837 & ~n62843;
  assign n62913 = ~n62864 & n62912;
  assign n62914 = n62850 & n62913;
  assign n62915 = ~n62899 & ~n62914;
  assign n62916 = ~n62878 & n62915;
  assign n62917 = n62856 & ~n62916;
  assign n62918 = ~n62911 & ~n62917;
  assign n62919 = ~n62843 & n62864;
  assign n62920 = n62856 & n62919;
  assign n62921 = ~n62850 & n62920;
  assign n62922 = n62918 & ~n62921;
  assign n62923 = ~n62905 & n62922;
  assign n62924 = ~n62889 & n62923;
  assign n62925 = ~pi1826 & ~n62924;
  assign n62926 = pi1826 & n62924;
  assign po1895 = n62925 | n62926;
  assign n62928 = n62850 & n62878;
  assign n62929 = ~n62901 & ~n62906;
  assign n62930 = n62856 & ~n62929;
  assign n62931 = ~n62928 & ~n62930;
  assign n62932 = ~n62892 & n62931;
  assign n62933 = ~n62856 & n62899;
  assign n62934 = ~n62884 & ~n62933;
  assign n62935 = ~n62914 & n62934;
  assign n62936 = n62932 & n62935;
  assign n62937 = n62831 & ~n62936;
  assign n62938 = n62864 & n62874;
  assign n62939 = n62850 & n62938;
  assign n62940 = ~n62872 & ~n62939;
  assign n62941 = n62844 & n62864;
  assign n62942 = n62856 & n62941;
  assign n62943 = n62850 & n62883;
  assign n62944 = ~n62942 & ~n62943;
  assign n62945 = n62843 & ~n62864;
  assign n62946 = ~n62837 & n62850;
  assign n62947 = ~n62945 & ~n62946;
  assign n62948 = ~n62919 & n62947;
  assign n62949 = ~n62856 & ~n62948;
  assign n62950 = ~n62850 & n62913;
  assign n62951 = ~n62879 & ~n62950;
  assign n62952 = ~n62949 & n62951;
  assign n62953 = n62944 & n62952;
  assign n62954 = n62940 & n62953;
  assign n62955 = ~n62831 & ~n62954;
  assign n62956 = ~n62937 & ~n62955;
  assign n62957 = pi1828 & ~n62956;
  assign n62958 = ~pi1828 & ~n62937;
  assign n62959 = ~n62955 & n62958;
  assign po1909 = n62957 | n62959;
  assign n62961 = ~n62756 & n62786;
  assign n62962 = n62756 & n62797;
  assign n62963 = ~n62783 & ~n62962;
  assign n62964 = n62730 & ~n62963;
  assign n62965 = ~n62961 & ~n62964;
  assign n62966 = ~n62730 & ~n62756;
  assign n62967 = n62748 & n62966;
  assign n62968 = ~n62742 & n62967;
  assign n62969 = n62764 & n62798;
  assign n62970 = ~n62968 & ~n62969;
  assign n62971 = ~n62730 & n62736;
  assign n62972 = n62758 & n62971;
  assign n62973 = n62970 & ~n62972;
  assign n62974 = ~n62760 & ~n62772;
  assign n62975 = ~n62748 & n62804;
  assign n62976 = n62974 & ~n62975;
  assign n62977 = n62973 & n62976;
  assign n62978 = n62965 & n62977;
  assign n62979 = ~n62795 & ~n62978;
  assign n62980 = ~n62759 & ~n62783;
  assign n62981 = n62756 & ~n62980;
  assign n62982 = ~n62742 & n62801;
  assign n62983 = ~n62812 & ~n62982;
  assign n62984 = n62736 & n62748;
  assign n62985 = n62756 & n62984;
  assign n62986 = n62983 & ~n62985;
  assign n62987 = n62730 & ~n62986;
  assign n62988 = ~n62756 & n62782;
  assign n62989 = ~n62742 & n62771;
  assign n62990 = ~n62988 & ~n62989;
  assign n62991 = ~n62730 & ~n62990;
  assign n62992 = ~n62756 & n62765;
  assign n62993 = ~n62991 & ~n62992;
  assign n62994 = ~n62987 & n62993;
  assign n62995 = ~n62981 & n62994;
  assign n62996 = n62795 & ~n62995;
  assign n62997 = n62730 & n62802;
  assign n62998 = ~n62996 & ~n62997;
  assign n62999 = n62777 & n62966;
  assign n63000 = n62748 & n62999;
  assign n63001 = n62998 & ~n63000;
  assign n63002 = ~n62979 & n63001;
  assign n63003 = ~pi1850 & ~n63002;
  assign n63004 = pi1850 & n62998;
  assign n63005 = ~n62979 & n63004;
  assign n63006 = ~n63000 & n63005;
  assign po1910 = n63003 | n63006;
  assign n63008 = pi6067 & ~pi9040;
  assign n63009 = pi6150 & pi9040;
  assign n63010 = ~n63008 & ~n63009;
  assign n63011 = ~pi1809 & ~n63010;
  assign n63012 = pi1809 & n63010;
  assign n63013 = ~n63011 & ~n63012;
  assign n63014 = pi6081 & pi9040;
  assign n63015 = pi6031 & ~pi9040;
  assign n63016 = ~n63014 & ~n63015;
  assign n63017 = ~pi1813 & ~n63016;
  assign n63018 = pi1813 & n63016;
  assign n63019 = ~n63017 & ~n63018;
  assign n63020 = ~n63013 & ~n63019;
  assign n63021 = pi6058 & ~pi9040;
  assign n63022 = pi6050 & pi9040;
  assign n63023 = ~n63021 & ~n63022;
  assign n63024 = pi1792 & n63023;
  assign n63025 = ~pi1792 & ~n63023;
  assign n63026 = ~n63024 & ~n63025;
  assign n63027 = pi6057 & pi9040;
  assign n63028 = pi6153 & ~pi9040;
  assign n63029 = ~n63027 & ~n63028;
  assign n63030 = ~pi1818 & ~n63029;
  assign n63031 = pi1818 & n63029;
  assign n63032 = ~n63030 & ~n63031;
  assign n63033 = pi6175 & ~pi9040;
  assign n63034 = pi6056 & pi9040;
  assign n63035 = ~n63033 & ~n63034;
  assign n63036 = pi1799 & n63035;
  assign n63037 = ~pi1799 & ~n63035;
  assign n63038 = ~n63036 & ~n63037;
  assign n63039 = n63032 & ~n63038;
  assign n63040 = ~n63026 & n63039;
  assign n63041 = pi6174 & pi9040;
  assign n63042 = pi6148 & ~pi9040;
  assign n63043 = ~n63041 & ~n63042;
  assign n63044 = ~pi1787 & n63043;
  assign n63045 = pi1787 & ~n63043;
  assign n63046 = ~n63044 & ~n63045;
  assign n63047 = n63038 & n63046;
  assign n63048 = n63032 & n63047;
  assign n63049 = n63026 & n63048;
  assign n63050 = n63038 & ~n63046;
  assign n63051 = ~n63026 & n63050;
  assign n63052 = ~n63049 & ~n63051;
  assign n63053 = ~n63040 & n63052;
  assign n63054 = n63020 & ~n63053;
  assign n63055 = ~n63026 & ~n63032;
  assign n63056 = n63046 & n63055;
  assign n63057 = ~n63038 & n63046;
  assign n63058 = n63032 & n63057;
  assign n63059 = n63026 & n63058;
  assign n63060 = ~n63056 & ~n63059;
  assign n63061 = ~n63032 & n63047;
  assign n63062 = n63032 & n63050;
  assign n63063 = ~n63061 & ~n63062;
  assign n63064 = n63060 & n63063;
  assign n63065 = n63013 & ~n63064;
  assign n63066 = n63026 & ~n63032;
  assign n63067 = ~n63046 & n63066;
  assign n63068 = ~n63038 & n63067;
  assign n63069 = ~n63065 & ~n63068;
  assign n63070 = ~n63019 & ~n63069;
  assign n63071 = ~n63054 & ~n63070;
  assign n63072 = n63013 & ~n63026;
  assign n63073 = n63032 & n63072;
  assign n63074 = ~n63046 & n63073;
  assign n63075 = n63038 & n63056;
  assign n63076 = ~n63074 & ~n63075;
  assign n63077 = ~n63032 & n63057;
  assign n63078 = ~n63050 & ~n63057;
  assign n63079 = n63026 & ~n63078;
  assign n63080 = ~n63077 & ~n63079;
  assign n63081 = ~n63013 & ~n63080;
  assign n63082 = ~n63038 & ~n63046;
  assign n63083 = n63032 & n63082;
  assign n63084 = ~n63040 & ~n63083;
  assign n63085 = ~n63049 & n63084;
  assign n63086 = n63013 & ~n63085;
  assign n63087 = ~n63081 & ~n63086;
  assign n63088 = ~n63013 & ~n63026;
  assign n63089 = n63047 & n63088;
  assign n63090 = n63026 & n63077;
  assign n63091 = ~n63032 & n63038;
  assign n63092 = ~n63046 & n63091;
  assign n63093 = n63026 & n63092;
  assign n63094 = ~n63090 & ~n63093;
  assign n63095 = ~n63046 & n63055;
  assign n63096 = ~n63038 & n63095;
  assign n63097 = n63094 & ~n63096;
  assign n63098 = ~n63089 & n63097;
  assign n63099 = n63087 & n63098;
  assign n63100 = n63019 & ~n63099;
  assign n63101 = n63076 & ~n63100;
  assign n63102 = n63071 & n63101;
  assign n63103 = pi1836 & ~n63102;
  assign n63104 = ~pi1836 & n63076;
  assign n63105 = n63071 & n63104;
  assign n63106 = ~n63100 & n63105;
  assign po1911 = n63103 | n63106;
  assign n63108 = ~n62757 & ~n62763;
  assign n63109 = ~n62730 & ~n63108;
  assign n63110 = ~n62819 & ~n63109;
  assign n63111 = ~n62736 & n62742;
  assign n63112 = n62730 & n63111;
  assign n63113 = n62756 & n63112;
  assign n63114 = n62756 & n62782;
  assign n63115 = ~n63111 & ~n63114;
  assign n63116 = n62736 & ~n62756;
  assign n63117 = ~n62742 & n63116;
  assign n63118 = n63115 & ~n63117;
  assign n63119 = n62730 & ~n63118;
  assign n63120 = ~n62766 & ~n63119;
  assign n63121 = ~n62795 & ~n63120;
  assign n63122 = ~n62730 & n62749;
  assign n63123 = n62756 & n63122;
  assign n63124 = ~n62972 & ~n63123;
  assign n63125 = ~n62795 & ~n63124;
  assign n63126 = ~n63121 & ~n63125;
  assign n63127 = ~n63113 & n63126;
  assign n63128 = ~n62783 & ~n62802;
  assign n63129 = ~n62812 & n63128;
  assign n63130 = ~n62730 & ~n63129;
  assign n63131 = ~n62756 & n62762;
  assign n63132 = ~n62786 & ~n63131;
  assign n63133 = n62730 & ~n63132;
  assign n63134 = ~n63130 & ~n63133;
  assign n63135 = ~n62982 & n63134;
  assign n63136 = ~n62772 & ~n62813;
  assign n63137 = n63135 & n63136;
  assign n63138 = n62795 & ~n63137;
  assign n63139 = n63127 & ~n63138;
  assign n63140 = n63110 & n63139;
  assign n63141 = ~pi1863 & ~n63140;
  assign n63142 = pi1863 & n63127;
  assign n63143 = n63110 & n63142;
  assign n63144 = ~n63138 & n63143;
  assign po1914 = n63141 | n63144;
  assign n63146 = pi6065 & pi9040;
  assign n63147 = pi6133 & ~pi9040;
  assign n63148 = ~n63146 & ~n63147;
  assign n63149 = pi1799 & n63148;
  assign n63150 = ~pi1799 & ~n63148;
  assign n63151 = ~n63149 & ~n63150;
  assign n63152 = pi6057 & ~pi9040;
  assign n63153 = pi6027 & pi9040;
  assign n63154 = ~n63152 & ~n63153;
  assign n63155 = pi1822 & n63154;
  assign n63156 = ~pi1822 & ~n63154;
  assign n63157 = ~n63155 & ~n63156;
  assign n63158 = pi6168 & pi9040;
  assign n63159 = pi6152 & ~pi9040;
  assign n63160 = ~n63158 & ~n63159;
  assign n63161 = ~pi1805 & n63160;
  assign n63162 = pi1805 & ~n63160;
  assign n63163 = ~n63161 & ~n63162;
  assign n63164 = pi6081 & ~pi9040;
  assign n63165 = pi6169 & pi9040;
  assign n63166 = ~n63164 & ~n63165;
  assign n63167 = ~pi1798 & ~n63166;
  assign n63168 = pi1798 & n63166;
  assign n63169 = ~n63167 & ~n63168;
  assign n63170 = pi6063 & ~pi9040;
  assign n63171 = pi6233 & pi9040;
  assign n63172 = ~n63170 & ~n63171;
  assign n63173 = ~pi1818 & ~n63172;
  assign n63174 = pi1818 & n63172;
  assign n63175 = ~n63173 & ~n63174;
  assign n63176 = n63169 & ~n63175;
  assign n63177 = ~n63163 & n63176;
  assign n63178 = n63157 & n63177;
  assign n63179 = pi6257 & ~pi9040;
  assign n63180 = pi6066 & pi9040;
  assign n63181 = ~n63179 & ~n63180;
  assign n63182 = pi1786 & n63181;
  assign n63183 = ~pi1786 & ~n63181;
  assign n63184 = ~n63182 & ~n63183;
  assign n63185 = ~n63163 & n63175;
  assign n63186 = n63169 & n63185;
  assign n63187 = n63163 & ~n63169;
  assign n63188 = ~n63169 & ~n63175;
  assign n63189 = ~n63157 & n63188;
  assign n63190 = n63163 & ~n63175;
  assign n63191 = n63157 & n63190;
  assign n63192 = ~n63189 & ~n63191;
  assign n63193 = ~n63187 & n63192;
  assign n63194 = ~n63186 & n63193;
  assign n63195 = n63184 & ~n63194;
  assign n63196 = ~n63157 & n63169;
  assign n63197 = n63175 & n63196;
  assign n63198 = n63163 & n63196;
  assign n63199 = ~n63169 & n63185;
  assign n63200 = ~n63198 & ~n63199;
  assign n63201 = ~n63184 & ~n63200;
  assign n63202 = ~n63197 & ~n63201;
  assign n63203 = ~n63195 & n63202;
  assign n63204 = ~n63178 & n63203;
  assign n63205 = n63151 & ~n63204;
  assign n63206 = n63163 & n63175;
  assign n63207 = ~n63169 & n63206;
  assign n63208 = ~n63157 & n63207;
  assign n63209 = ~n63169 & n63190;
  assign n63210 = n63157 & n63209;
  assign n63211 = ~n63178 & ~n63210;
  assign n63212 = ~n63208 & n63211;
  assign n63213 = n63184 & ~n63212;
  assign n63214 = ~n63205 & ~n63213;
  assign n63215 = ~n63163 & n63197;
  assign n63216 = ~n63163 & ~n63169;
  assign n63217 = ~n63184 & n63216;
  assign n63218 = n63157 & n63217;
  assign n63219 = ~n63157 & n63184;
  assign n63220 = n63169 & n63219;
  assign n63221 = ~n63175 & n63220;
  assign n63222 = n63169 & n63206;
  assign n63223 = n63157 & n63222;
  assign n63224 = ~n63221 & ~n63223;
  assign n63225 = n63163 & n63169;
  assign n63226 = n63157 & n63225;
  assign n63227 = ~n63163 & ~n63175;
  assign n63228 = ~n63169 & n63227;
  assign n63229 = ~n63226 & ~n63228;
  assign n63230 = ~n63184 & ~n63229;
  assign n63231 = ~n63184 & n63187;
  assign n63232 = ~n63157 & n63231;
  assign n63233 = ~n63230 & ~n63232;
  assign n63234 = n63224 & n63233;
  assign n63235 = ~n63151 & ~n63234;
  assign n63236 = ~n63218 & ~n63235;
  assign n63237 = ~n63215 & n63236;
  assign n63238 = n63214 & n63237;
  assign n63239 = ~pi1830 & ~n63238;
  assign n63240 = ~n63205 & ~n63215;
  assign n63241 = ~n63213 & n63240;
  assign n63242 = n63236 & n63241;
  assign n63243 = pi1830 & n63242;
  assign po1917 = n63239 | n63243;
  assign n63245 = pi6052 & pi9040;
  assign n63246 = pi6082 & ~pi9040;
  assign n63247 = ~n63245 & ~n63246;
  assign n63248 = pi1816 & n63247;
  assign n63249 = ~pi1816 & ~n63247;
  assign n63250 = ~n63248 & ~n63249;
  assign n63251 = pi6294 & ~pi9040;
  assign n63252 = pi6143 & pi9040;
  assign n63253 = ~n63251 & ~n63252;
  assign n63254 = ~pi1794 & ~n63253;
  assign n63255 = pi1794 & n63253;
  assign n63256 = ~n63254 & ~n63255;
  assign n63257 = pi6078 & ~pi9040;
  assign n63258 = pi6176 & pi9040;
  assign n63259 = ~n63257 & ~n63258;
  assign n63260 = ~pi1812 & n63259;
  assign n63261 = pi1812 & ~n63259;
  assign n63262 = ~n63260 & ~n63261;
  assign n63263 = n63256 & n63262;
  assign n63264 = pi6064 & ~pi9040;
  assign n63265 = pi6082 & pi9040;
  assign n63266 = ~n63264 & ~n63265;
  assign n63267 = ~pi1811 & ~n63266;
  assign n63268 = pi1811 & n63266;
  assign n63269 = ~n63267 & ~n63268;
  assign n63270 = pi6038 & ~pi9040;
  assign n63271 = pi6154 & pi9040;
  assign n63272 = ~n63270 & ~n63271;
  assign n63273 = ~pi1785 & n63272;
  assign n63274 = pi1785 & ~n63272;
  assign n63275 = ~n63273 & ~n63274;
  assign n63276 = n63269 & ~n63275;
  assign n63277 = n63263 & n63276;
  assign n63278 = n63269 & n63275;
  assign n63279 = ~n63256 & n63278;
  assign n63280 = ~n63277 & ~n63279;
  assign n63281 = ~n63250 & ~n63280;
  assign n63282 = pi6147 & pi9040;
  assign n63283 = pi6159 & ~pi9040;
  assign n63284 = ~n63282 & ~n63283;
  assign n63285 = ~pi1804 & ~n63284;
  assign n63286 = pi1804 & n63284;
  assign n63287 = ~n63285 & ~n63286;
  assign n63288 = n63250 & ~n63269;
  assign n63289 = n63256 & n63288;
  assign n63290 = n63263 & n63275;
  assign n63291 = n63256 & ~n63262;
  assign n63292 = ~n63275 & n63291;
  assign n63293 = ~n63290 & ~n63292;
  assign n63294 = ~n63256 & n63262;
  assign n63295 = ~n63275 & n63294;
  assign n63296 = n63269 & n63295;
  assign n63297 = n63293 & ~n63296;
  assign n63298 = n63250 & ~n63297;
  assign n63299 = ~n63289 & ~n63298;
  assign n63300 = ~n63256 & ~n63262;
  assign n63301 = n63275 & n63300;
  assign n63302 = n63269 & n63301;
  assign n63303 = n63299 & ~n63302;
  assign n63304 = ~n63269 & n63294;
  assign n63305 = ~n63275 & n63300;
  assign n63306 = ~n63304 & ~n63305;
  assign n63307 = ~n63250 & ~n63306;
  assign n63308 = n63275 & n63291;
  assign n63309 = ~n63269 & n63308;
  assign n63310 = ~n63307 & ~n63309;
  assign n63311 = n63303 & n63310;
  assign n63312 = n63287 & ~n63311;
  assign n63313 = ~n63281 & ~n63312;
  assign n63314 = n63250 & ~n63287;
  assign n63315 = ~n63306 & n63314;
  assign n63316 = n63275 & n63294;
  assign n63317 = ~n63308 & ~n63316;
  assign n63318 = n63269 & ~n63317;
  assign n63319 = ~n63277 & ~n63318;
  assign n63320 = ~n63287 & ~n63319;
  assign n63321 = ~n63315 & ~n63320;
  assign n63322 = ~n63250 & ~n63287;
  assign n63323 = n63263 & ~n63269;
  assign n63324 = ~n63301 & ~n63323;
  assign n63325 = n63256 & ~n63275;
  assign n63326 = n63324 & ~n63325;
  assign n63327 = n63322 & ~n63326;
  assign n63328 = n63321 & ~n63327;
  assign n63329 = n63313 & n63328;
  assign n63330 = ~pi1829 & ~n63329;
  assign n63331 = pi1829 & n63321;
  assign n63332 = n63313 & n63331;
  assign n63333 = ~n63327 & n63332;
  assign po1918 = n63330 | n63333;
  assign n63335 = ~n63077 & ~n63083;
  assign n63336 = ~n63013 & ~n63335;
  assign n63337 = n63026 & n63062;
  assign n63338 = ~n63336 & ~n63337;
  assign n63339 = n63026 & n63038;
  assign n63340 = ~n63091 & ~n63339;
  assign n63341 = ~n63058 & n63340;
  assign n63342 = n63013 & ~n63341;
  assign n63343 = n63338 & ~n63342;
  assign n63344 = ~n63019 & ~n63343;
  assign n63345 = ~n63026 & n63092;
  assign n63346 = ~n63013 & n63345;
  assign n63347 = ~n63026 & n63048;
  assign n63348 = ~n63013 & n63347;
  assign n63349 = ~n63346 & ~n63348;
  assign n63350 = n63013 & n63096;
  assign n63351 = n63349 & ~n63350;
  assign n63352 = ~n63032 & n63082;
  assign n63353 = n63013 & n63352;
  assign n63354 = ~n63026 & n63032;
  assign n63355 = n63046 & n63354;
  assign n63356 = ~n63096 & ~n63355;
  assign n63357 = ~n63026 & n63038;
  assign n63358 = n63032 & n63357;
  assign n63359 = n63013 & n63358;
  assign n63360 = n63026 & n63083;
  assign n63361 = ~n63013 & n63091;
  assign n63362 = ~n63360 & ~n63361;
  assign n63363 = ~n63090 & n63362;
  assign n63364 = ~n63359 & n63363;
  assign n63365 = n63356 & n63364;
  assign n63366 = ~n63353 & n63365;
  assign n63367 = n63019 & ~n63366;
  assign n63368 = n63351 & ~n63367;
  assign n63369 = ~n63344 & n63368;
  assign n63370 = ~pi1845 & ~n63369;
  assign n63371 = pi1845 & n63351;
  assign n63372 = ~n63344 & n63371;
  assign n63373 = ~n63367 & n63372;
  assign po1920 = n63370 | n63373;
  assign n63375 = ~n62850 & n62874;
  assign n63376 = ~n62950 & ~n63375;
  assign n63377 = n62856 & n63376;
  assign n63378 = n62850 & n62908;
  assign n63379 = ~n62844 & ~n62868;
  assign n63380 = ~n62864 & ~n63379;
  assign n63381 = n62837 & n62890;
  assign n63382 = n62850 & n62868;
  assign n63383 = ~n63381 & ~n63382;
  assign n63384 = ~n63380 & n63383;
  assign n63385 = ~n62856 & n63384;
  assign n63386 = ~n63378 & n63385;
  assign n63387 = ~n63377 & ~n63386;
  assign n63388 = n62850 & n63380;
  assign n63389 = ~n62939 & ~n63388;
  assign n63390 = ~n63387 & n63389;
  assign n63391 = n62831 & ~n63390;
  assign n63392 = n62856 & ~n63379;
  assign n63393 = ~n62850 & n63392;
  assign n63394 = ~n62885 & ~n62912;
  assign n63395 = n62850 & ~n63394;
  assign n63396 = n62856 & n63395;
  assign n63397 = n62864 & n63392;
  assign n63398 = ~n63396 & ~n63397;
  assign n63399 = ~n63393 & n63398;
  assign n63400 = ~n62831 & ~n63399;
  assign n63401 = ~n63391 & ~n63400;
  assign n63402 = ~n62856 & ~n63376;
  assign n63403 = ~n62872 & ~n63402;
  assign n63404 = ~n62831 & ~n63403;
  assign n63405 = n62856 & n62872;
  assign n63406 = ~n62856 & ~n63389;
  assign n63407 = ~n63405 & ~n63406;
  assign n63408 = ~n63404 & n63407;
  assign n63409 = n63401 & n63408;
  assign n63410 = pi1846 & ~n63409;
  assign n63411 = ~pi1846 & n63408;
  assign n63412 = ~n63400 & n63411;
  assign n63413 = ~n63391 & n63412;
  assign po1922 = n63410 | n63413;
  assign n63415 = pi6062 & pi9040;
  assign n63416 = pi6176 & ~pi9040;
  assign n63417 = ~n63415 & ~n63416;
  assign n63418 = ~pi1794 & ~n63417;
  assign n63419 = pi1794 & n63417;
  assign n63420 = ~n63418 & ~n63419;
  assign n63421 = pi6051 & ~pi9040;
  assign n63422 = pi6084 & pi9040;
  assign n63423 = ~n63421 & ~n63422;
  assign n63424 = ~pi1815 & ~n63423;
  assign n63425 = pi1815 & n63423;
  assign n63426 = ~n63424 & ~n63425;
  assign n63427 = pi6298 & pi9040;
  assign n63428 = pi6041 & ~pi9040;
  assign n63429 = ~n63427 & ~n63428;
  assign n63430 = ~pi1820 & n63429;
  assign n63431 = pi1820 & ~n63429;
  assign n63432 = ~n63430 & ~n63431;
  assign n63433 = pi6298 & ~pi9040;
  assign n63434 = pi6070 & pi9040;
  assign n63435 = ~n63433 & ~n63434;
  assign n63436 = ~pi1785 & n63435;
  assign n63437 = pi1785 & ~n63435;
  assign n63438 = ~n63436 & ~n63437;
  assign n63439 = n63432 & ~n63438;
  assign n63440 = pi6149 & pi9040;
  assign n63441 = pi6259 & ~pi9040;
  assign n63442 = ~n63440 & ~n63441;
  assign n63443 = ~pi1800 & ~n63442;
  assign n63444 = pi1800 & n63442;
  assign n63445 = ~n63443 & ~n63444;
  assign n63446 = pi6070 & ~pi9040;
  assign n63447 = pi6064 & pi9040;
  assign n63448 = ~n63446 & ~n63447;
  assign n63449 = pi1821 & n63448;
  assign n63450 = ~pi1821 & ~n63448;
  assign n63451 = ~n63449 & ~n63450;
  assign n63452 = n63445 & n63451;
  assign n63453 = n63439 & n63452;
  assign n63454 = n63426 & n63453;
  assign n63455 = ~n63445 & n63451;
  assign n63456 = ~n63432 & ~n63438;
  assign n63457 = n63455 & n63456;
  assign n63458 = n63426 & ~n63445;
  assign n63459 = n63438 & n63458;
  assign n63460 = n63432 & n63459;
  assign n63461 = ~n63432 & n63438;
  assign n63462 = n63426 & n63461;
  assign n63463 = n63451 & n63462;
  assign n63464 = n63445 & n63463;
  assign n63465 = ~n63460 & ~n63464;
  assign n63466 = ~n63457 & n63465;
  assign n63467 = ~n63454 & n63466;
  assign n63468 = ~n63426 & ~n63445;
  assign n63469 = ~n63438 & n63468;
  assign n63470 = ~n63432 & n63469;
  assign n63471 = n63467 & ~n63470;
  assign n63472 = ~n63420 & ~n63471;
  assign n63473 = n63426 & ~n63432;
  assign n63474 = ~n63438 & n63473;
  assign n63475 = n63445 & n63474;
  assign n63476 = ~n63459 & ~n63475;
  assign n63477 = ~n63426 & n63439;
  assign n63478 = n63445 & n63477;
  assign n63479 = n63476 & ~n63478;
  assign n63480 = ~n63451 & ~n63479;
  assign n63481 = ~n63426 & n63438;
  assign n63482 = ~n63432 & n63481;
  assign n63483 = ~n63451 & n63482;
  assign n63484 = n63445 & n63483;
  assign n63485 = n63432 & n63458;
  assign n63486 = n63432 & n63438;
  assign n63487 = ~n63445 & n63486;
  assign n63488 = ~n63485 & ~n63487;
  assign n63489 = ~n63451 & ~n63488;
  assign n63490 = ~n63484 & ~n63489;
  assign n63491 = ~n63420 & ~n63490;
  assign n63492 = ~n63480 & ~n63491;
  assign n63493 = ~n63472 & n63492;
  assign n63494 = ~n63426 & n63445;
  assign n63495 = n63451 & n63494;
  assign n63496 = n63486 & n63495;
  assign n63497 = ~n63426 & ~n63432;
  assign n63498 = n63455 & n63497;
  assign n63499 = ~n63445 & n63482;
  assign n63500 = n63426 & ~n63451;
  assign n63501 = ~n63432 & n63500;
  assign n63502 = n63432 & n63445;
  assign n63503 = ~n63426 & n63502;
  assign n63504 = ~n63501 & ~n63503;
  assign n63505 = ~n63499 & n63504;
  assign n63506 = ~n63477 & n63505;
  assign n63507 = n63439 & n63451;
  assign n63508 = ~n63445 & n63507;
  assign n63509 = n63445 & n63486;
  assign n63510 = ~n63426 & ~n63438;
  assign n63511 = ~n63509 & ~n63510;
  assign n63512 = n63451 & ~n63511;
  assign n63513 = ~n63508 & ~n63512;
  assign n63514 = n63506 & n63513;
  assign n63515 = n63420 & ~n63514;
  assign n63516 = ~n63498 & ~n63515;
  assign n63517 = ~n63496 & n63516;
  assign n63518 = n63493 & n63517;
  assign n63519 = pi1825 & n63518;
  assign n63520 = ~pi1825 & ~n63518;
  assign po1924 = n63519 | n63520;
  assign n63522 = ~n63032 & ~n63038;
  assign n63523 = ~n63047 & ~n63522;
  assign n63524 = n63026 & ~n63523;
  assign n63525 = ~n63026 & n63083;
  assign n63526 = ~n63524 & ~n63525;
  assign n63527 = ~n63345 & n63526;
  assign n63528 = ~n63013 & ~n63527;
  assign n63529 = n63026 & n63039;
  assign n63530 = ~n63062 & ~n63529;
  assign n63531 = ~n63075 & n63530;
  assign n63532 = n63013 & ~n63531;
  assign n63533 = ~n63528 & ~n63532;
  assign n63534 = n63019 & ~n63533;
  assign n63535 = ~n63038 & n63072;
  assign n63536 = ~n63358 & ~n63529;
  assign n63537 = ~n63013 & ~n63536;
  assign n63538 = ~n63089 & ~n63537;
  assign n63539 = ~n63093 & ~n63347;
  assign n63540 = n63013 & n63026;
  assign n63541 = n63091 & n63540;
  assign n63542 = ~n63353 & ~n63541;
  assign n63543 = n63539 & n63542;
  assign n63544 = n63538 & n63543;
  assign n63545 = ~n63535 & n63544;
  assign n63546 = ~n63019 & ~n63545;
  assign n63547 = ~n63013 & n63077;
  assign n63548 = ~n63026 & n63547;
  assign n63549 = ~n63348 & ~n63548;
  assign n63550 = ~n63350 & n63549;
  assign n63551 = ~n63026 & n63058;
  assign n63552 = n63026 & n63050;
  assign n63553 = ~n63551 & ~n63552;
  assign n63554 = n63013 & ~n63553;
  assign n63555 = n63550 & ~n63554;
  assign n63556 = ~n63546 & n63555;
  assign n63557 = ~n63534 & n63556;
  assign n63558 = ~pi1839 & ~n63557;
  assign n63559 = pi1839 & n63557;
  assign po1925 = n63558 | n63559;
  assign n63561 = ~n62813 & ~n62992;
  assign n63562 = n62730 & ~n63561;
  assign n63563 = ~n62760 & ~n62763;
  assign n63564 = ~n62756 & n62812;
  assign n63565 = ~n62962 & ~n63564;
  assign n63566 = n63563 & n63565;
  assign n63567 = ~n62730 & ~n63566;
  assign n63568 = ~n62795 & n62797;
  assign n63569 = ~n62730 & n63568;
  assign n63570 = n62742 & n63116;
  assign n63571 = ~n62984 & ~n63570;
  assign n63572 = ~n62765 & n63571;
  assign n63573 = n62730 & ~n63572;
  assign n63574 = ~n62736 & n62782;
  assign n63575 = ~n62756 & n63574;
  assign n63576 = ~n63573 & ~n63575;
  assign n63577 = ~n62795 & ~n63576;
  assign n63578 = ~n63569 & ~n63577;
  assign n63579 = ~n62736 & ~n62742;
  assign n63580 = ~n62730 & n63579;
  assign n63581 = n62756 & n63580;
  assign n63582 = ~n62756 & n62984;
  assign n63583 = ~n62763 & ~n63582;
  assign n63584 = ~n62989 & n63583;
  assign n63585 = ~n63581 & n63584;
  assign n63586 = n62730 & n62759;
  assign n63587 = n63585 & ~n63586;
  assign n63588 = n62795 & ~n63587;
  assign n63589 = n63578 & ~n63588;
  assign n63590 = ~n63567 & n63589;
  assign n63591 = ~n63562 & n63590;
  assign n63592 = pi1870 & n63591;
  assign n63593 = ~pi1870 & ~n63591;
  assign po1926 = n63592 | n63593;
  assign n63595 = pi6054 & ~pi9040;
  assign n63596 = pi6071 & pi9040;
  assign n63597 = ~n63595 & ~n63596;
  assign n63598 = ~pi1805 & ~n63597;
  assign n63599 = pi1805 & n63597;
  assign n63600 = ~n63598 & ~n63599;
  assign n63601 = pi6060 & pi9040;
  assign n63602 = pi6059 & ~pi9040;
  assign n63603 = ~n63601 & ~n63602;
  assign n63604 = ~pi1808 & n63603;
  assign n63605 = pi1808 & ~n63603;
  assign n63606 = ~n63604 & ~n63605;
  assign n63607 = pi6151 & pi9040;
  assign n63608 = pi6297 & ~pi9040;
  assign n63609 = ~n63607 & ~n63608;
  assign n63610 = pi1807 & n63609;
  assign n63611 = ~pi1807 & ~n63609;
  assign n63612 = ~n63610 & ~n63611;
  assign n63613 = pi6053 & ~pi9040;
  assign n63614 = pi6297 & pi9040;
  assign n63615 = ~n63613 & ~n63614;
  assign n63616 = pi1806 & n63615;
  assign n63617 = ~pi1806 & ~n63615;
  assign n63618 = ~n63616 & ~n63617;
  assign n63619 = pi6149 & ~pi9040;
  assign n63620 = pi6159 & pi9040;
  assign n63621 = ~n63619 & ~n63620;
  assign n63622 = ~pi1798 & n63621;
  assign n63623 = pi1798 & ~n63621;
  assign n63624 = ~n63622 & ~n63623;
  assign n63625 = ~n63618 & ~n63624;
  assign n63626 = n63612 & n63625;
  assign n63627 = ~n63606 & n63626;
  assign n63628 = pi6062 & ~pi9040;
  assign n63629 = pi6259 & pi9040;
  assign n63630 = ~n63628 & ~n63629;
  assign n63631 = ~pi1823 & ~n63630;
  assign n63632 = pi1823 & n63630;
  assign n63633 = ~n63631 & ~n63632;
  assign n63634 = ~pi1806 & n63615;
  assign n63635 = pi1806 & ~n63615;
  assign n63636 = ~n63634 & ~n63635;
  assign n63637 = ~n63624 & ~n63636;
  assign n63638 = ~n63606 & n63637;
  assign n63639 = ~n63612 & n63625;
  assign n63640 = n63606 & n63639;
  assign n63641 = ~n63638 & ~n63640;
  assign n63642 = ~n63633 & ~n63641;
  assign n63643 = ~n63627 & ~n63642;
  assign n63644 = ~n63618 & n63624;
  assign n63645 = ~n63612 & n63644;
  assign n63646 = n63633 & n63645;
  assign n63647 = n63625 & n63633;
  assign n63648 = ~n63606 & n63647;
  assign n63649 = ~n63646 & ~n63648;
  assign n63650 = n63643 & n63649;
  assign n63651 = n63624 & ~n63636;
  assign n63652 = n63612 & n63651;
  assign n63653 = ~n63606 & n63652;
  assign n63654 = n63612 & n63644;
  assign n63655 = n63606 & n63654;
  assign n63656 = ~n63653 & ~n63655;
  assign n63657 = n63650 & n63656;
  assign n63658 = n63600 & ~n63657;
  assign n63659 = ~n63600 & ~n63633;
  assign n63660 = ~n63606 & ~n63612;
  assign n63661 = n63636 & n63660;
  assign n63662 = ~n63612 & n63624;
  assign n63663 = ~n63661 & ~n63662;
  assign n63664 = n63659 & ~n63663;
  assign n63665 = n63606 & n63612;
  assign n63666 = ~n63624 & n63665;
  assign n63667 = ~n63618 & n63666;
  assign n63668 = n63606 & ~n63636;
  assign n63669 = ~n63612 & n63668;
  assign n63670 = ~n63667 & ~n63669;
  assign n63671 = ~n63606 & n63633;
  assign n63672 = ~n63625 & n63671;
  assign n63673 = n63612 & n63672;
  assign n63674 = n63633 & n63652;
  assign n63675 = ~n63673 & ~n63674;
  assign n63676 = n63670 & n63675;
  assign n63677 = ~n63600 & ~n63676;
  assign n63678 = ~n63612 & n63651;
  assign n63679 = ~n63633 & n63678;
  assign n63680 = n63606 & n63679;
  assign n63681 = n63612 & n63637;
  assign n63682 = n63606 & n63681;
  assign n63683 = ~n63655 & ~n63682;
  assign n63684 = ~n63633 & ~n63683;
  assign n63685 = ~n63680 & ~n63684;
  assign n63686 = n63633 & n63667;
  assign n63687 = n63685 & ~n63686;
  assign n63688 = ~n63677 & n63687;
  assign n63689 = ~n63664 & n63688;
  assign n63690 = ~n63658 & n63689;
  assign n63691 = ~n63612 & n63637;
  assign n63692 = n63606 & n63633;
  assign n63693 = n63691 & n63692;
  assign n63694 = n63690 & ~n63693;
  assign n63695 = ~pi1835 & ~n63694;
  assign n63696 = ~n63658 & ~n63693;
  assign n63697 = n63689 & n63696;
  assign n63698 = pi1835 & n63697;
  assign po1927 = n63695 | n63698;
  assign n63700 = n62850 & n62941;
  assign n63701 = n62856 & n63700;
  assign n63702 = n62890 & ~n63379;
  assign n63703 = ~n62913 & ~n63702;
  assign n63704 = ~n62939 & n63703;
  assign n63705 = ~n62856 & ~n63704;
  assign n63706 = n62850 & n62869;
  assign n63707 = ~n63705 & ~n63706;
  assign n63708 = n62864 & n62912;
  assign n63709 = ~n62850 & n62945;
  assign n63710 = ~n63708 & ~n63709;
  assign n63711 = ~n63382 & n63710;
  assign n63712 = n62856 & ~n63711;
  assign n63713 = n63707 & ~n63712;
  assign n63714 = n62831 & ~n63713;
  assign n63715 = ~n63701 & ~n63714;
  assign n63716 = ~n62914 & ~n63700;
  assign n63717 = n62850 & n62919;
  assign n63718 = ~n62945 & ~n63717;
  assign n63719 = ~n63708 & n63718;
  assign n63720 = ~n62856 & ~n63719;
  assign n63721 = ~n62850 & n62869;
  assign n63722 = ~n62850 & n62868;
  assign n63723 = ~n62938 & ~n63722;
  assign n63724 = n62856 & ~n63723;
  assign n63725 = ~n63721 & ~n63724;
  assign n63726 = ~n63720 & n63725;
  assign n63727 = n63716 & n63726;
  assign n63728 = ~n62886 & n63727;
  assign n63729 = ~n62831 & ~n63728;
  assign n63730 = ~n62896 & ~n63378;
  assign n63731 = ~n62856 & ~n63730;
  assign n63732 = ~n63729 & ~n63731;
  assign n63733 = n63715 & n63732;
  assign n63734 = pi1851 & n63733;
  assign n63735 = ~pi1851 & ~n63733;
  assign po1928 = n63734 | n63735;
  assign n63737 = ~n63157 & ~n63184;
  assign n63738 = ~n63163 & n63737;
  assign n63739 = n63169 & n63190;
  assign n63740 = n63157 & n63739;
  assign n63741 = n63157 & n63207;
  assign n63742 = ~n63740 & ~n63741;
  assign n63743 = ~n63157 & n63209;
  assign n63744 = ~n63199 & ~n63743;
  assign n63745 = n63184 & ~n63744;
  assign n63746 = n63742 & ~n63745;
  assign n63747 = ~n63738 & n63746;
  assign n63748 = n63151 & ~n63747;
  assign n63749 = n63157 & n63228;
  assign n63750 = ~n63184 & n63749;
  assign n63751 = n63219 & n63228;
  assign n63752 = ~n63198 & ~n63751;
  assign n63753 = ~n63199 & ~n63222;
  assign n63754 = ~n63157 & n63206;
  assign n63755 = n63753 & ~n63754;
  assign n63756 = ~n63184 & ~n63755;
  assign n63757 = n63184 & n63186;
  assign n63758 = n63211 & ~n63757;
  assign n63759 = ~n63756 & n63758;
  assign n63760 = n63752 & n63759;
  assign n63761 = ~n63151 & ~n63760;
  assign n63762 = ~n63750 & ~n63761;
  assign n63763 = ~n63748 & n63762;
  assign n63764 = n63219 & n63222;
  assign n63765 = n63176 & n63184;
  assign n63766 = n63157 & n63765;
  assign n63767 = ~n63764 & ~n63766;
  assign n63768 = n63184 & n63741;
  assign n63769 = n63767 & ~n63768;
  assign n63770 = n63763 & n63769;
  assign n63771 = ~pi1834 & ~n63770;
  assign n63772 = pi1834 & n63769;
  assign n63773 = n63762 & n63772;
  assign n63774 = ~n63748 & n63773;
  assign po1929 = n63771 | n63774;
  assign n63776 = n63606 & n63645;
  assign n63777 = n63624 & n63660;
  assign n63778 = ~n63636 & n63777;
  assign n63779 = ~n63776 & ~n63778;
  assign n63780 = n63633 & ~n63779;
  assign n63781 = ~n63667 & ~n63674;
  assign n63782 = ~n63606 & n63612;
  assign n63783 = ~n63624 & n63782;
  assign n63784 = ~n63636 & n63783;
  assign n63785 = ~n63606 & ~n63633;
  assign n63786 = n63644 & n63785;
  assign n63787 = ~n63612 & n63786;
  assign n63788 = ~n63618 & n63665;
  assign n63789 = ~n63669 & ~n63788;
  assign n63790 = ~n63633 & ~n63789;
  assign n63791 = ~n63612 & n63633;
  assign n63792 = ~n63624 & n63791;
  assign n63793 = ~n63618 & n63792;
  assign n63794 = ~n63790 & ~n63793;
  assign n63795 = ~n63787 & n63794;
  assign n63796 = ~n63784 & n63795;
  assign n63797 = n63781 & n63796;
  assign n63798 = n63600 & ~n63797;
  assign n63799 = ~n63633 & n63667;
  assign n63800 = n63606 & n63674;
  assign n63801 = ~n63799 & ~n63800;
  assign n63802 = ~n63798 & n63801;
  assign n63803 = ~n63780 & n63802;
  assign n63804 = n63612 & ~n63618;
  assign n63805 = n63671 & n63804;
  assign n63806 = ~n63646 & ~n63805;
  assign n63807 = n63633 & n63681;
  assign n63808 = n63606 & n63691;
  assign n63809 = ~n63807 & ~n63808;
  assign n63810 = ~n63606 & n63654;
  assign n63811 = ~n63776 & ~n63810;
  assign n63812 = ~n63606 & n63651;
  assign n63813 = ~n63612 & ~n63624;
  assign n63814 = ~n63812 & ~n63813;
  assign n63815 = ~n63633 & ~n63814;
  assign n63816 = n63811 & ~n63815;
  assign n63817 = n63809 & n63816;
  assign n63818 = n63806 & n63817;
  assign n63819 = ~n63600 & ~n63818;
  assign n63820 = n63803 & ~n63819;
  assign n63821 = ~pi1827 & ~n63820;
  assign n63822 = pi1827 & n63803;
  assign n63823 = ~n63819 & n63822;
  assign po1930 = n63821 | n63823;
  assign n63825 = ~n63157 & n63739;
  assign n63826 = ~n63207 & ~n63215;
  assign n63827 = n63157 & n63176;
  assign n63828 = ~n63157 & n63228;
  assign n63829 = ~n63827 & ~n63828;
  assign n63830 = n63826 & n63829;
  assign n63831 = ~n63184 & ~n63830;
  assign n63832 = n63157 & n63185;
  assign n63833 = ~n63198 & ~n63832;
  assign n63834 = ~n63209 & n63833;
  assign n63835 = n63184 & ~n63834;
  assign n63836 = n63157 & ~n63169;
  assign n63837 = n63175 & n63836;
  assign n63838 = ~n63163 & n63837;
  assign n63839 = ~n63835 & ~n63838;
  assign n63840 = ~n63831 & n63839;
  assign n63841 = ~n63825 & n63840;
  assign n63842 = ~n63151 & ~n63841;
  assign n63843 = n63157 & ~n63184;
  assign n63844 = n63186 & n63843;
  assign n63845 = ~n63184 & n63209;
  assign n63846 = ~n63184 & n63222;
  assign n63847 = ~n63845 & ~n63846;
  assign n63848 = ~n63157 & ~n63847;
  assign n63849 = ~n63844 & ~n63848;
  assign n63850 = ~n63157 & n63177;
  assign n63851 = ~n63749 & ~n63850;
  assign n63852 = n63157 & n63206;
  assign n63853 = ~n63157 & n63185;
  assign n63854 = ~n63852 & ~n63853;
  assign n63855 = ~n63177 & n63854;
  assign n63856 = ~n63207 & n63855;
  assign n63857 = n63184 & ~n63856;
  assign n63858 = ~n63157 & n63199;
  assign n63859 = ~n63857 & ~n63858;
  assign n63860 = n63851 & n63859;
  assign n63861 = n63849 & n63860;
  assign n63862 = n63151 & ~n63861;
  assign n63863 = ~n63184 & ~n63742;
  assign n63864 = ~n63862 & ~n63863;
  assign n63865 = ~n63210 & ~n63850;
  assign n63866 = n63184 & ~n63865;
  assign n63867 = n63864 & ~n63866;
  assign n63868 = ~n63842 & n63867;
  assign n63869 = pi1840 & ~n63868;
  assign n63870 = ~pi1840 & n63868;
  assign po1931 = n63869 | n63870;
  assign n63872 = n63426 & n63432;
  assign n63873 = ~n63470 & ~n63872;
  assign n63874 = ~n63502 & n63873;
  assign n63875 = n63451 & ~n63874;
  assign n63876 = n63445 & ~n63451;
  assign n63877 = ~n63432 & n63876;
  assign n63878 = ~n63426 & n63432;
  assign n63879 = ~n63445 & ~n63451;
  assign n63880 = n63878 & n63879;
  assign n63881 = n63426 & n63445;
  assign n63882 = ~n63438 & n63881;
  assign n63883 = ~n63445 & n63462;
  assign n63884 = ~n63882 & ~n63883;
  assign n63885 = ~n63880 & n63884;
  assign n63886 = ~n63877 & n63885;
  assign n63887 = ~n63875 & n63886;
  assign n63888 = n63420 & ~n63887;
  assign n63889 = n63426 & n63439;
  assign n63890 = ~n63445 & n63889;
  assign n63891 = n63426 & n63486;
  assign n63892 = n63445 & n63891;
  assign n63893 = ~n63890 & ~n63892;
  assign n63894 = n63451 & ~n63893;
  assign n63895 = ~n63888 & ~n63894;
  assign n63896 = n63445 & n63462;
  assign n63897 = ~n63474 & ~n63482;
  assign n63898 = n63451 & ~n63897;
  assign n63899 = ~n63896 & ~n63898;
  assign n63900 = ~n63478 & n63899;
  assign n63901 = ~n63420 & ~n63900;
  assign n63902 = ~n63456 & ~n63486;
  assign n63903 = ~n63426 & ~n63902;
  assign n63904 = ~n63487 & ~n63903;
  assign n63905 = ~n63451 & ~n63904;
  assign n63906 = ~n63420 & n63905;
  assign n63907 = ~n63901 & ~n63906;
  assign n63908 = n63895 & n63907;
  assign n63909 = pi1831 & ~n63908;
  assign n63910 = ~pi1831 & n63895;
  assign n63911 = n63907 & n63910;
  assign po1932 = n63909 | n63911;
  assign n63913 = ~n63250 & n63269;
  assign n63914 = ~n63294 & ~n63308;
  assign n63915 = n63913 & ~n63914;
  assign n63916 = ~n63250 & n63275;
  assign n63917 = n63294 & n63916;
  assign n63918 = ~n63915 & ~n63917;
  assign n63919 = n63287 & ~n63918;
  assign n63920 = ~n63269 & ~n63275;
  assign n63921 = ~n63262 & n63920;
  assign n63922 = n63256 & n63921;
  assign n63923 = ~n63325 & ~n63920;
  assign n63924 = n63250 & ~n63923;
  assign n63925 = ~n63269 & n63275;
  assign n63926 = n63262 & n63925;
  assign n63927 = n63256 & n63926;
  assign n63928 = ~n63924 & ~n63927;
  assign n63929 = ~n63922 & n63928;
  assign n63930 = n63287 & ~n63929;
  assign n63931 = ~n63919 & ~n63930;
  assign n63932 = ~n63262 & n63276;
  assign n63933 = ~n63256 & n63932;
  assign n63934 = ~n63269 & n63301;
  assign n63935 = ~n63933 & ~n63934;
  assign n63936 = ~n63250 & ~n63935;
  assign n63937 = n63269 & n63316;
  assign n63938 = ~n63269 & n63325;
  assign n63939 = ~n63937 & ~n63938;
  assign n63940 = n63250 & ~n63939;
  assign n63941 = ~n63263 & ~n63325;
  assign n63942 = n63269 & ~n63941;
  assign n63943 = ~n63301 & ~n63942;
  assign n63944 = ~n63250 & ~n63943;
  assign n63945 = ~n63262 & ~n63269;
  assign n63946 = n63916 & n63945;
  assign n63947 = n63262 & ~n63275;
  assign n63948 = ~n63301 & ~n63947;
  assign n63949 = ~n63269 & ~n63948;
  assign n63950 = n63250 & n63269;
  assign n63951 = n63291 & n63950;
  assign n63952 = n63275 & n63951;
  assign n63953 = ~n63949 & ~n63952;
  assign n63954 = ~n63946 & n63953;
  assign n63955 = ~n63944 & n63954;
  assign n63956 = ~n63933 & n63955;
  assign n63957 = ~n63287 & ~n63956;
  assign n63958 = ~n63940 & ~n63957;
  assign n63959 = ~n63936 & n63958;
  assign n63960 = n63931 & n63959;
  assign n63961 = pi1832 & n63960;
  assign n63962 = ~pi1832 & ~n63960;
  assign po1933 = n63961 | n63962;
  assign n63964 = n63013 & n63050;
  assign n63965 = ~n63026 & n63964;
  assign n63966 = ~n63551 & ~n63965;
  assign n63967 = n63026 & ~n63046;
  assign n63968 = n63032 & n63967;
  assign n63969 = ~n63026 & ~n63038;
  assign n63970 = ~n63355 & ~n63969;
  assign n63971 = ~n63013 & ~n63970;
  assign n63972 = ~n63968 & ~n63971;
  assign n63973 = n63966 & n63972;
  assign n63974 = n63019 & ~n63973;
  assign n63975 = ~n63048 & ~n63093;
  assign n63976 = ~n63026 & n63082;
  assign n63977 = n63975 & ~n63976;
  assign n63978 = n63013 & ~n63977;
  assign n63979 = n63050 & n63088;
  assign n63980 = ~n63075 & ~n63979;
  assign n63981 = ~n63978 & n63980;
  assign n63982 = ~n63058 & ~n63068;
  assign n63983 = ~n63013 & ~n63982;
  assign n63984 = n63981 & ~n63983;
  assign n63985 = ~n63019 & ~n63984;
  assign n63986 = ~n63974 & ~n63985;
  assign n63987 = ~n63026 & n63057;
  assign n63988 = n63026 & ~n63063;
  assign n63989 = ~n63987 & ~n63988;
  assign n63990 = ~n63013 & ~n63989;
  assign n63991 = ~n63048 & n63335;
  assign n63992 = n63540 & ~n63991;
  assign n63993 = ~n63990 & ~n63992;
  assign n63994 = n63986 & n63993;
  assign n63995 = ~pi1833 & ~n63994;
  assign n63996 = ~n63985 & n63993;
  assign n63997 = pi1833 & n63996;
  assign n63998 = ~n63974 & n63997;
  assign po1934 = n63995 | n63998;
  assign n64000 = ~n63445 & n63477;
  assign n64001 = ~n63883 & ~n64000;
  assign n64002 = ~n63451 & ~n64001;
  assign n64003 = n63474 & n63876;
  assign n64004 = ~n64002 & ~n64003;
  assign n64005 = ~n63498 & n64004;
  assign n64006 = n63426 & n63451;
  assign n64007 = n63438 & n64006;
  assign n64008 = n63432 & n64007;
  assign n64009 = ~n63445 & n64008;
  assign n64010 = n63451 & n63889;
  assign n64011 = ~n63470 & ~n63496;
  assign n64012 = ~n63464 & n64011;
  assign n64013 = ~n64010 & n64012;
  assign n64014 = n63420 & ~n64013;
  assign n64015 = n63445 & n63482;
  assign n64016 = ~n63477 & ~n64015;
  assign n64017 = ~n63891 & n64016;
  assign n64018 = ~n63451 & ~n64017;
  assign n64019 = n63420 & n64018;
  assign n64020 = n63445 & n63507;
  assign n64021 = ~n64008 & ~n64020;
  assign n64022 = ~n63882 & n64021;
  assign n64023 = n63438 & n63468;
  assign n64024 = n63445 & n63456;
  assign n64025 = ~n63473 & ~n64024;
  assign n64026 = ~n63451 & ~n64025;
  assign n64027 = ~n64023 & ~n64026;
  assign n64028 = n64022 & n64027;
  assign n64029 = ~n63420 & ~n64028;
  assign n64030 = ~n64019 & ~n64029;
  assign n64031 = ~n64014 & n64030;
  assign n64032 = ~n64009 & n64031;
  assign n64033 = n64005 & n64032;
  assign n64034 = pi1837 & ~n64033;
  assign n64035 = ~pi1837 & n64005;
  assign n64036 = n64032 & n64035;
  assign po1935 = n64034 | n64036;
  assign n64038 = ~n63800 & ~n63805;
  assign n64039 = ~n63606 & n63639;
  assign n64040 = ~n63784 & ~n64039;
  assign n64041 = ~n63776 & n64040;
  assign n64042 = ~n63633 & ~n64041;
  assign n64043 = ~n63667 & ~n63678;
  assign n64044 = ~n63812 & n64043;
  assign n64045 = ~n63633 & ~n64044;
  assign n64046 = ~n63693 & n64040;
  assign n64047 = n63633 & n63654;
  assign n64048 = n64046 & ~n64047;
  assign n64049 = ~n64045 & n64048;
  assign n64050 = n63600 & ~n64049;
  assign n64051 = n63618 & n63665;
  assign n64052 = ~n63810 & ~n64051;
  assign n64053 = ~n63633 & n63637;
  assign n64054 = n63606 & n64053;
  assign n64055 = ~n63633 & n63645;
  assign n64056 = ~n64054 & ~n64055;
  assign n64057 = n63606 & n63647;
  assign n64058 = n63618 & n63660;
  assign n64059 = ~n63678 & ~n64058;
  assign n64060 = n63633 & ~n64059;
  assign n64061 = ~n64057 & ~n64060;
  assign n64062 = n64056 & n64061;
  assign n64063 = n64052 & n64062;
  assign n64064 = ~n63776 & n64063;
  assign n64065 = ~n63600 & ~n64064;
  assign n64066 = ~n64050 & ~n64065;
  assign n64067 = ~n64042 & n64066;
  assign n64068 = n64038 & n64067;
  assign n64069 = pi1841 & ~n64068;
  assign n64070 = ~pi1841 & n64068;
  assign po1936 = n64069 | n64070;
  assign n64072 = n63262 & n63278;
  assign n64073 = ~n63308 & ~n64072;
  assign n64074 = ~n63250 & ~n64073;
  assign n64075 = n63269 & n63300;
  assign n64076 = ~n63926 & ~n64075;
  assign n64077 = n63250 & ~n64076;
  assign n64078 = ~n63269 & n63295;
  assign n64079 = ~n63946 & ~n64078;
  assign n64080 = ~n63277 & n64079;
  assign n64081 = ~n64077 & n64080;
  assign n64082 = ~n64074 & n64081;
  assign n64083 = ~n63922 & ~n63933;
  assign n64084 = n64082 & n64083;
  assign n64085 = n63287 & ~n64084;
  assign n64086 = n63263 & n63920;
  assign n64087 = n63317 & ~n64086;
  assign n64088 = n63250 & ~n64087;
  assign n64089 = ~n63269 & n63305;
  assign n64090 = ~n64088 & ~n64089;
  assign n64091 = n63256 & n63278;
  assign n64092 = n63269 & n63291;
  assign n64093 = ~n64091 & ~n64092;
  assign n64094 = n63250 & ~n64093;
  assign n64095 = n63250 & n63300;
  assign n64096 = ~n63269 & n64095;
  assign n64097 = ~n64094 & ~n64096;
  assign n64098 = n64090 & n64097;
  assign n64099 = ~n63287 & ~n64098;
  assign n64100 = ~n63295 & ~n63302;
  assign n64101 = ~n63927 & n64100;
  assign n64102 = n63322 & ~n64101;
  assign n64103 = ~n64099 & ~n64102;
  assign n64104 = ~n63277 & ~n63922;
  assign n64105 = ~n63250 & ~n64104;
  assign n64106 = n64103 & ~n64105;
  assign n64107 = ~n64085 & n64106;
  assign n64108 = ~pi1844 & n64107;
  assign n64109 = pi1844 & ~n64107;
  assign po1937 = n64108 | n64109;
  assign n64111 = pi6078 & pi9040;
  assign n64112 = pi6154 & ~pi9040;
  assign n64113 = ~n64111 & ~n64112;
  assign n64114 = ~pi1812 & ~n64113;
  assign n64115 = pi1812 & n64113;
  assign n64116 = ~n64114 & ~n64115;
  assign n64117 = pi6084 & ~pi9040;
  assign n64118 = pi6059 & pi9040;
  assign n64119 = ~n64117 & ~n64118;
  assign n64120 = ~pi1807 & ~n64119;
  assign n64121 = pi1807 & n64119;
  assign n64122 = ~n64120 & ~n64121;
  assign n64123 = pi6035 & ~pi9040;
  assign n64124 = pi6041 & pi9040;
  assign n64125 = ~n64123 & ~n64124;
  assign n64126 = ~pi1804 & n64125;
  assign n64127 = pi1804 & ~n64125;
  assign n64128 = ~n64126 & ~n64127;
  assign n64129 = ~n64122 & ~n64128;
  assign n64130 = ~n64116 & n64129;
  assign n64131 = n64122 & ~n64128;
  assign n64132 = n64116 & n64131;
  assign n64133 = ~n64130 & ~n64132;
  assign n64134 = pi6294 & pi9040;
  assign n64135 = pi6147 & ~pi9040;
  assign n64136 = ~n64134 & ~n64135;
  assign n64137 = pi1801 & n64136;
  assign n64138 = ~pi1801 & ~n64136;
  assign n64139 = ~n64137 & ~n64138;
  assign n64140 = n64116 & ~n64139;
  assign n64141 = n64122 & n64140;
  assign n64142 = n64133 & ~n64141;
  assign n64143 = pi6071 & ~pi9040;
  assign n64144 = pi6035 & pi9040;
  assign n64145 = ~n64143 & ~n64144;
  assign n64146 = ~pi1797 & ~n64145;
  assign n64147 = pi1797 & n64145;
  assign n64148 = ~n64146 & ~n64147;
  assign n64149 = pi6051 & pi9040;
  assign n64150 = pi6151 & ~pi9040;
  assign n64151 = ~n64149 & ~n64150;
  assign n64152 = ~pi1806 & ~n64151;
  assign n64153 = pi1806 & n64151;
  assign n64154 = ~n64152 & ~n64153;
  assign n64155 = ~n64148 & n64154;
  assign n64156 = ~n64142 & n64155;
  assign n64157 = ~n64122 & n64128;
  assign n64158 = n64116 & n64157;
  assign n64159 = n64139 & n64154;
  assign n64160 = n64158 & n64159;
  assign n64161 = n64116 & n64129;
  assign n64162 = n64148 & n64161;
  assign n64163 = n64122 & n64128;
  assign n64164 = n64139 & n64163;
  assign n64165 = ~n64116 & n64122;
  assign n64166 = ~n64164 & ~n64165;
  assign n64167 = n64148 & ~n64166;
  assign n64168 = ~n64162 & ~n64167;
  assign n64169 = n64154 & ~n64168;
  assign n64170 = ~n64160 & ~n64169;
  assign n64171 = ~n64139 & n64157;
  assign n64172 = ~n64116 & n64171;
  assign n64173 = ~n64116 & n64139;
  assign n64174 = n64122 & n64173;
  assign n64175 = ~n64172 & ~n64174;
  assign n64176 = n64148 & ~n64175;
  assign n64177 = n64170 & ~n64176;
  assign n64178 = n64139 & ~n64148;
  assign n64179 = n64163 & n64178;
  assign n64180 = n64116 & n64179;
  assign n64181 = ~n64116 & n64163;
  assign n64182 = ~n64139 & ~n64148;
  assign n64183 = n64181 & n64182;
  assign n64184 = ~n64131 & ~n64157;
  assign n64185 = n64173 & ~n64184;
  assign n64186 = n64139 & n64161;
  assign n64187 = ~n64185 & ~n64186;
  assign n64188 = n64140 & ~n64184;
  assign n64189 = n64130 & ~n64139;
  assign n64190 = ~n64188 & ~n64189;
  assign n64191 = n64187 & n64190;
  assign n64192 = ~n64183 & n64191;
  assign n64193 = ~n64180 & n64192;
  assign n64194 = ~n64139 & n64148;
  assign n64195 = n64116 & n64194;
  assign n64196 = n64128 & n64195;
  assign n64197 = n64193 & ~n64196;
  assign n64198 = ~n64154 & ~n64197;
  assign n64199 = n64177 & ~n64198;
  assign n64200 = ~n64156 & n64199;
  assign n64201 = ~pi1865 & ~n64200;
  assign n64202 = pi1865 & n64177;
  assign n64203 = ~n64156 & n64202;
  assign n64204 = ~n64198 & n64203;
  assign po1938 = n64201 | n64204;
  assign n64206 = n64116 & n64163;
  assign n64207 = n64148 & n64206;
  assign n64208 = ~n64139 & n64207;
  assign n64209 = n64129 & n64194;
  assign n64210 = ~n64116 & n64209;
  assign n64211 = ~n64208 & ~n64210;
  assign n64212 = ~n64183 & ~n64189;
  assign n64213 = n64116 & ~n64128;
  assign n64214 = n64139 & n64213;
  assign n64215 = ~n64164 & ~n64214;
  assign n64216 = n64148 & ~n64215;
  assign n64217 = ~n64116 & ~n64139;
  assign n64218 = ~n64148 & ~n64217;
  assign n64219 = ~n64184 & n64218;
  assign n64220 = ~n64139 & ~n64163;
  assign n64221 = n64148 & n64220;
  assign n64222 = ~n64116 & n64221;
  assign n64223 = ~n64219 & ~n64222;
  assign n64224 = ~n64216 & n64223;
  assign n64225 = n64212 & n64224;
  assign n64226 = n64154 & ~n64225;
  assign n64227 = n64211 & ~n64226;
  assign n64228 = n64132 & ~n64148;
  assign n64229 = n64139 & n64228;
  assign n64230 = ~n64148 & ~n64154;
  assign n64231 = ~n64161 & ~n64164;
  assign n64232 = ~n64184 & n64217;
  assign n64233 = n64231 & ~n64232;
  assign n64234 = n64230 & ~n64233;
  assign n64235 = n64130 & n64139;
  assign n64236 = ~n64128 & n64139;
  assign n64237 = ~n64116 & n64236;
  assign n64238 = n64139 & n64157;
  assign n64239 = ~n64237 & ~n64238;
  assign n64240 = ~n64139 & n64163;
  assign n64241 = ~n64158 & ~n64240;
  assign n64242 = n64239 & n64241;
  assign n64243 = n64148 & ~n64242;
  assign n64244 = ~n64235 & ~n64243;
  assign n64245 = ~n64154 & ~n64244;
  assign n64246 = ~n64234 & ~n64245;
  assign n64247 = ~n64229 & n64246;
  assign n64248 = n64227 & n64247;
  assign n64249 = pi1859 & ~n64248;
  assign n64250 = ~pi1859 & n64227;
  assign n64251 = n64247 & n64250;
  assign po1939 = n64249 | n64251;
  assign n64253 = ~n64238 & ~n64240;
  assign n64254 = n64148 & ~n64253;
  assign n64255 = ~n64210 & ~n64254;
  assign n64256 = n64154 & ~n64255;
  assign n64257 = ~n64116 & ~n64128;
  assign n64258 = ~n64131 & ~n64257;
  assign n64259 = ~n64139 & ~n64258;
  assign n64260 = ~n64206 & ~n64259;
  assign n64261 = ~n64148 & ~n64260;
  assign n64262 = ~n64232 & ~n64261;
  assign n64263 = n64139 & n64181;
  assign n64264 = ~n64122 & n64140;
  assign n64265 = n64139 & ~n64258;
  assign n64266 = ~n64264 & ~n64265;
  assign n64267 = n64148 & ~n64266;
  assign n64268 = ~n64263 & ~n64267;
  assign n64269 = n64262 & n64268;
  assign n64270 = ~n64154 & ~n64269;
  assign n64271 = n64116 & n64139;
  assign n64272 = ~n64131 & n64271;
  assign n64273 = n64154 & n64272;
  assign n64274 = n64131 & n64173;
  assign n64275 = n64148 & n64274;
  assign n64276 = n64116 & ~n64122;
  assign n64277 = n64178 & n64276;
  assign n64278 = ~n64275 & ~n64277;
  assign n64279 = ~n64273 & n64278;
  assign n64280 = ~n64158 & ~n64236;
  assign n64281 = n64155 & ~n64280;
  assign n64282 = n64279 & ~n64281;
  assign n64283 = ~n64270 & n64282;
  assign n64284 = ~n64256 & n64283;
  assign n64285 = pi1867 & ~n64284;
  assign n64286 = ~pi1867 & n64284;
  assign po1940 = n64285 | n64286;
  assign n64288 = ~n63481 & ~n63889;
  assign n64289 = n63455 & ~n64288;
  assign n64290 = ~n63477 & ~n63482;
  assign n64291 = ~n63474 & ~n63891;
  assign n64292 = n64290 & n64291;
  assign n64293 = n63445 & ~n64292;
  assign n64294 = ~n64289 & ~n64293;
  assign n64295 = ~n63883 & n64294;
  assign n64296 = n63420 & ~n64295;
  assign n64297 = n63445 & ~n63902;
  assign n64298 = ~n63426 & n64297;
  assign n64299 = n63438 & n63881;
  assign n64300 = ~n63510 & ~n64299;
  assign n64301 = ~n63891 & n64300;
  assign n64302 = n63451 & ~n64301;
  assign n64303 = ~n63451 & ~n64288;
  assign n64304 = ~n64302 & ~n64303;
  assign n64305 = ~n64298 & n64304;
  assign n64306 = ~n63445 & n63474;
  assign n64307 = n64305 & ~n64306;
  assign n64308 = ~n63420 & ~n64307;
  assign n64309 = n63445 & n63889;
  assign n64310 = ~n64306 & ~n64309;
  assign n64311 = ~n63451 & ~n64310;
  assign n64312 = ~n64308 & ~n64311;
  assign n64313 = ~n64296 & n64312;
  assign n64314 = ~pi1838 & ~n64313;
  assign n64315 = pi1838 & ~n64311;
  assign n64316 = ~n64296 & n64315;
  assign n64317 = ~n64308 & n64316;
  assign po1941 = n64314 | n64317;
  assign n64319 = ~n63653 & ~n63661;
  assign n64320 = n63600 & ~n64319;
  assign n64321 = ~n63666 & ~n63788;
  assign n64322 = ~n63626 & n64321;
  assign n64323 = ~n63633 & ~n64322;
  assign n64324 = n63600 & n64323;
  assign n64325 = ~n64320 & ~n64324;
  assign n64326 = n63652 & n63785;
  assign n64327 = ~n63787 & ~n64326;
  assign n64328 = ~n63669 & ~n63813;
  assign n64329 = n63633 & ~n64328;
  assign n64330 = n63600 & n64329;
  assign n64331 = n64327 & ~n64330;
  assign n64332 = n63606 & n63652;
  assign n64333 = n63606 & n63644;
  assign n64334 = ~n63778 & ~n64333;
  assign n64335 = n63633 & ~n64334;
  assign n64336 = ~n63667 & ~n63784;
  assign n64337 = n63606 & n63651;
  assign n64338 = ~n63691 & ~n64337;
  assign n64339 = ~n63633 & ~n64338;
  assign n64340 = n64336 & ~n64339;
  assign n64341 = ~n64335 & n64340;
  assign n64342 = ~n64332 & n64341;
  assign n64343 = ~n63600 & ~n64342;
  assign n64344 = ~n63810 & n64040;
  assign n64345 = n63633 & ~n64344;
  assign n64346 = ~n64343 & ~n64345;
  assign n64347 = n64331 & n64346;
  assign n64348 = n64325 & n64347;
  assign n64349 = ~pi1842 & ~n64348;
  assign n64350 = pi1842 & n64331;
  assign n64351 = n64325 & n64350;
  assign n64352 = n64346 & n64351;
  assign po1942 = n64349 | n64352;
  assign n64354 = ~n64116 & n64131;
  assign n64355 = ~n64206 & ~n64354;
  assign n64356 = n64148 & ~n64355;
  assign n64357 = ~n64132 & ~n64171;
  assign n64358 = ~n64181 & n64357;
  assign n64359 = ~n64148 & ~n64358;
  assign n64360 = ~n64356 & ~n64359;
  assign n64361 = ~n64162 & ~n64172;
  assign n64362 = n64360 & n64361;
  assign n64363 = ~n64154 & ~n64362;
  assign n64364 = n64139 & n64206;
  assign n64365 = n64129 & ~n64139;
  assign n64366 = ~n64238 & ~n64365;
  assign n64367 = ~n64148 & ~n64366;
  assign n64368 = ~n64364 & ~n64367;
  assign n64369 = n64116 & n64148;
  assign n64370 = ~n64122 & n64369;
  assign n64371 = n64128 & n64370;
  assign n64372 = n64133 & ~n64371;
  assign n64373 = ~n64181 & n64372;
  assign n64374 = ~n64139 & ~n64373;
  assign n64375 = n64368 & ~n64374;
  assign n64376 = n64154 & ~n64375;
  assign n64377 = ~n64363 & ~n64376;
  assign n64378 = ~n64116 & n64238;
  assign n64379 = ~n64186 & ~n64378;
  assign n64380 = n64148 & ~n64379;
  assign n64381 = ~n64148 & n64257;
  assign n64382 = n64139 & n64381;
  assign n64383 = ~n64380 & ~n64382;
  assign n64384 = n64377 & n64383;
  assign n64385 = ~pi1852 & ~n64384;
  assign n64386 = pi1852 & ~n64380;
  assign n64387 = n64377 & n64386;
  assign n64388 = ~n64382 & n64387;
  assign po1943 = n64385 | n64388;
  assign n64390 = ~n63743 & ~n63850;
  assign n64391 = ~n63838 & n64390;
  assign n64392 = ~n63184 & ~n64391;
  assign n64393 = ~n63751 & ~n63768;
  assign n64394 = ~n63749 & ~n63846;
  assign n64395 = ~n63739 & ~n63853;
  assign n64396 = n63184 & ~n64395;
  assign n64397 = ~n63215 & ~n64396;
  assign n64398 = n64394 & n64397;
  assign n64399 = n63151 & ~n64398;
  assign n64400 = ~n63169 & n63175;
  assign n64401 = ~n63187 & ~n64400;
  assign n64402 = n63157 & ~n64401;
  assign n64403 = ~n63177 & ~n63754;
  assign n64404 = n63184 & ~n64403;
  assign n64405 = n63157 & n63175;
  assign n64406 = ~n63199 & ~n64405;
  assign n64407 = ~n63190 & n64406;
  assign n64408 = ~n63184 & ~n64407;
  assign n64409 = ~n64404 & ~n64408;
  assign n64410 = ~n64402 & n64409;
  assign n64411 = ~n63151 & ~n64410;
  assign n64412 = ~n64399 & ~n64411;
  assign n64413 = n64393 & n64412;
  assign n64414 = ~n64392 & n64413;
  assign n64415 = ~pi1847 & ~n64414;
  assign n64416 = pi1847 & n64393;
  assign n64417 = ~n64392 & n64416;
  assign n64418 = n64412 & n64417;
  assign po1944 = n64415 | n64418;
  assign n64420 = ~n63269 & n63291;
  assign n64421 = ~n63290 & ~n64420;
  assign n64422 = ~n63250 & ~n64421;
  assign n64423 = n63250 & ~n63948;
  assign n64424 = ~n63937 & ~n64423;
  assign n64425 = ~n64422 & n64424;
  assign n64426 = n63287 & ~n64425;
  assign n64427 = ~n63250 & n63305;
  assign n64428 = ~n64426 & ~n64427;
  assign n64429 = ~n64078 & ~n64092;
  assign n64430 = n63250 & ~n64429;
  assign n64431 = n63250 & n63292;
  assign n64432 = n63269 & n63308;
  assign n64433 = ~n63250 & n63276;
  assign n64434 = ~n63925 & ~n64433;
  assign n64435 = ~n63256 & ~n64434;
  assign n64436 = ~n63926 & ~n64435;
  assign n64437 = ~n63277 & n64436;
  assign n64438 = ~n64432 & n64437;
  assign n64439 = ~n64431 & n64438;
  assign n64440 = ~n63287 & ~n64439;
  assign n64441 = ~n64430 & ~n64440;
  assign n64442 = n64428 & n64441;
  assign n64443 = pi1853 & ~n64442;
  assign n64444 = ~pi1853 & n64442;
  assign po1945 = n64443 | n64444;
  assign n64446 = pi6403 & pi9040;
  assign n64447 = pi6311 & ~pi9040;
  assign n64448 = ~n64446 & ~n64447;
  assign n64449 = pi1861 & n64448;
  assign n64450 = ~pi1861 & ~n64448;
  assign n64451 = ~n64449 & ~n64450;
  assign n64452 = pi6261 & ~pi9040;
  assign n64453 = pi6293 & pi9040;
  assign n64454 = ~n64452 & ~n64453;
  assign n64455 = ~pi1879 & n64454;
  assign n64456 = pi1879 & ~n64454;
  assign n64457 = ~n64455 & ~n64456;
  assign n64458 = pi6304 & ~pi9040;
  assign n64459 = pi6369 & pi9040;
  assign n64460 = ~n64458 & ~n64459;
  assign n64461 = pi1848 & n64460;
  assign n64462 = ~pi1848 & ~n64460;
  assign n64463 = ~n64461 & ~n64462;
  assign n64464 = pi6372 & ~pi9040;
  assign n64465 = pi6286 & pi9040;
  assign n64466 = ~n64464 & ~n64465;
  assign n64467 = pi1866 & n64466;
  assign n64468 = ~pi1866 & ~n64466;
  assign n64469 = ~n64467 & ~n64468;
  assign n64470 = ~n64463 & n64469;
  assign n64471 = ~n64457 & n64470;
  assign n64472 = n64451 & n64471;
  assign n64473 = pi6372 & pi9040;
  assign n64474 = pi6397 & ~pi9040;
  assign n64475 = ~n64473 & ~n64474;
  assign n64476 = ~pi1855 & ~n64475;
  assign n64477 = pi1855 & n64475;
  assign n64478 = ~n64476 & ~n64477;
  assign n64479 = n64457 & ~n64463;
  assign n64480 = ~n64451 & n64479;
  assign n64481 = n64478 & n64480;
  assign n64482 = ~n64472 & ~n64481;
  assign n64483 = pi6311 & pi9040;
  assign n64484 = pi6296 & ~pi9040;
  assign n64485 = ~n64483 & ~n64484;
  assign n64486 = ~pi1885 & n64485;
  assign n64487 = pi1885 & ~n64485;
  assign n64488 = ~n64486 & ~n64487;
  assign n64489 = ~n64469 & n64488;
  assign n64490 = n64451 & n64478;
  assign n64491 = ~n64463 & n64490;
  assign n64492 = ~n64451 & n64478;
  assign n64493 = ~n64457 & n64492;
  assign n64494 = n64463 & n64493;
  assign n64495 = ~n64491 & ~n64494;
  assign n64496 = ~n64457 & ~n64478;
  assign n64497 = ~n64463 & n64496;
  assign n64498 = n64495 & ~n64497;
  assign n64499 = n64489 & ~n64498;
  assign n64500 = ~n64451 & ~n64478;
  assign n64501 = ~n64457 & n64500;
  assign n64502 = n64463 & n64501;
  assign n64503 = ~n64480 & ~n64502;
  assign n64504 = n64457 & n64492;
  assign n64505 = ~n64457 & n64490;
  assign n64506 = ~n64504 & ~n64505;
  assign n64507 = n64503 & n64506;
  assign n64508 = n64469 & ~n64507;
  assign n64509 = n64451 & ~n64478;
  assign n64510 = n64457 & n64509;
  assign n64511 = n64463 & n64510;
  assign n64512 = ~n64508 & ~n64511;
  assign n64513 = n64488 & ~n64512;
  assign n64514 = ~n64499 & ~n64513;
  assign n64515 = n64457 & n64500;
  assign n64516 = ~n64490 & ~n64500;
  assign n64517 = n64463 & ~n64516;
  assign n64518 = ~n64515 & ~n64517;
  assign n64519 = ~n64469 & ~n64518;
  assign n64520 = ~n64457 & n64509;
  assign n64521 = ~n64497 & ~n64520;
  assign n64522 = ~n64494 & n64521;
  assign n64523 = n64469 & ~n64522;
  assign n64524 = ~n64519 & ~n64523;
  assign n64525 = ~n64463 & ~n64469;
  assign n64526 = n64492 & n64525;
  assign n64527 = n64463 & n64515;
  assign n64528 = n64457 & n64478;
  assign n64529 = n64451 & n64528;
  assign n64530 = n64463 & n64529;
  assign n64531 = ~n64527 & ~n64530;
  assign n64532 = n64451 & n64479;
  assign n64533 = ~n64478 & n64532;
  assign n64534 = n64531 & ~n64533;
  assign n64535 = ~n64526 & n64534;
  assign n64536 = n64524 & n64535;
  assign n64537 = ~n64488 & ~n64536;
  assign n64538 = n64514 & ~n64537;
  assign n64539 = n64482 & n64538;
  assign n64540 = pi1891 & ~n64539;
  assign n64541 = ~pi1891 & n64482;
  assign n64542 = n64514 & n64541;
  assign n64543 = ~n64537 & n64542;
  assign po1961 = n64540 | n64543;
  assign n64545 = pi6304 & pi9040;
  assign n64546 = pi6278 & ~pi9040;
  assign n64547 = ~n64545 & ~n64546;
  assign n64548 = ~pi1849 & n64547;
  assign n64549 = pi1849 & ~n64547;
  assign n64550 = ~n64548 & ~n64549;
  assign n64551 = pi6467 & ~pi9040;
  assign n64552 = pi6300 & pi9040;
  assign n64553 = ~n64551 & ~n64552;
  assign n64554 = ~pi1864 & n64553;
  assign n64555 = pi1864 & ~n64553;
  assign n64556 = ~n64554 & ~n64555;
  assign n64557 = pi6286 & ~pi9040;
  assign n64558 = pi6314 & pi9040;
  assign n64559 = ~n64557 & ~n64558;
  assign n64560 = ~pi1873 & n64559;
  assign n64561 = pi1873 & ~n64559;
  assign n64562 = ~n64560 & ~n64561;
  assign n64563 = pi6296 & pi9040;
  assign n64564 = pi6322 & ~pi9040;
  assign n64565 = ~n64563 & ~n64564;
  assign n64566 = ~pi1857 & n64565;
  assign n64567 = pi1857 & ~n64565;
  assign n64568 = ~n64566 & ~n64567;
  assign n64569 = ~n64562 & ~n64568;
  assign n64570 = n64556 & n64569;
  assign n64571 = pi6396 & pi9040;
  assign n64572 = pi6291 & ~pi9040;
  assign n64573 = ~n64571 & ~n64572;
  assign n64574 = pi1887 & n64573;
  assign n64575 = ~pi1887 & ~n64573;
  assign n64576 = ~n64574 & ~n64575;
  assign n64577 = n64570 & ~n64576;
  assign n64578 = n64562 & n64568;
  assign n64579 = n64556 & ~n64576;
  assign n64580 = n64578 & n64579;
  assign n64581 = ~n64577 & ~n64580;
  assign n64582 = ~n64556 & n64578;
  assign n64583 = n64576 & n64582;
  assign n64584 = ~n64562 & n64568;
  assign n64585 = n64556 & n64584;
  assign n64586 = n64576 & n64585;
  assign n64587 = ~n64583 & ~n64586;
  assign n64588 = n64581 & n64587;
  assign n64589 = ~n64550 & ~n64588;
  assign n64590 = n64562 & ~n64568;
  assign n64591 = n64556 & n64590;
  assign n64592 = n64576 & n64591;
  assign n64593 = ~n64585 & ~n64592;
  assign n64594 = ~n64550 & ~n64593;
  assign n64595 = n64550 & ~n64568;
  assign n64596 = ~n64576 & n64595;
  assign n64597 = ~n64556 & ~n64562;
  assign n64598 = n64576 & n64578;
  assign n64599 = ~n64597 & ~n64598;
  assign n64600 = n64550 & ~n64599;
  assign n64601 = ~n64596 & ~n64600;
  assign n64602 = ~n64556 & n64590;
  assign n64603 = ~n64576 & n64602;
  assign n64604 = n64601 & ~n64603;
  assign n64605 = ~n64568 & n64597;
  assign n64606 = n64576 & n64605;
  assign n64607 = n64604 & ~n64606;
  assign n64608 = ~n64594 & n64607;
  assign n64609 = ~pi6466 & pi9040;
  assign n64610 = ~pi6300 & ~pi9040;
  assign n64611 = ~n64609 & ~n64610;
  assign n64612 = ~pi1881 & n64611;
  assign n64613 = pi1881 & ~n64611;
  assign n64614 = ~n64612 & ~n64613;
  assign n64615 = ~n64608 & ~n64614;
  assign n64616 = n64556 & ~n64568;
  assign n64617 = n64550 & n64576;
  assign n64618 = n64614 & n64617;
  assign n64619 = n64616 & n64618;
  assign n64620 = n64568 & n64579;
  assign n64621 = n64550 & ~n64620;
  assign n64622 = ~n64556 & n64576;
  assign n64623 = n64562 & n64622;
  assign n64624 = ~n64569 & ~n64616;
  assign n64625 = ~n64576 & ~n64624;
  assign n64626 = ~n64550 & ~n64582;
  assign n64627 = ~n64625 & n64626;
  assign n64628 = ~n64623 & n64627;
  assign n64629 = ~n64621 & ~n64628;
  assign n64630 = n64568 & n64622;
  assign n64631 = ~n64562 & n64630;
  assign n64632 = ~n64629 & ~n64631;
  assign n64633 = n64614 & ~n64632;
  assign n64634 = ~n64619 & ~n64633;
  assign n64635 = ~n64615 & n64634;
  assign n64636 = ~n64589 & n64635;
  assign n64637 = n64550 & n64603;
  assign n64638 = n64636 & ~n64637;
  assign n64639 = pi1888 & ~n64638;
  assign n64640 = ~pi1888 & ~n64637;
  assign n64641 = n64635 & n64640;
  assign n64642 = ~n64589 & n64641;
  assign po1971 = n64639 | n64642;
  assign n64644 = ~n64515 & ~n64520;
  assign n64645 = ~n64469 & ~n64644;
  assign n64646 = n64463 & n64505;
  assign n64647 = ~n64645 & ~n64646;
  assign n64648 = n64463 & n64478;
  assign n64649 = ~n64528 & ~n64648;
  assign n64650 = ~n64501 & n64649;
  assign n64651 = n64469 & ~n64650;
  assign n64652 = n64647 & ~n64651;
  assign n64653 = n64488 & ~n64652;
  assign n64654 = ~n64463 & n64529;
  assign n64655 = ~n64469 & n64654;
  assign n64656 = ~n64457 & ~n64463;
  assign n64657 = ~n64451 & n64656;
  assign n64658 = n64478 & n64657;
  assign n64659 = ~n64469 & n64658;
  assign n64660 = ~n64655 & ~n64659;
  assign n64661 = n64469 & n64533;
  assign n64662 = n64660 & ~n64661;
  assign n64663 = n64457 & n64469;
  assign n64664 = n64451 & n64663;
  assign n64665 = ~n64478 & n64664;
  assign n64666 = ~n64533 & ~n64657;
  assign n64667 = n64478 & n64656;
  assign n64668 = n64469 & n64667;
  assign n64669 = n64463 & n64520;
  assign n64670 = ~n64469 & n64528;
  assign n64671 = ~n64669 & ~n64670;
  assign n64672 = ~n64527 & n64671;
  assign n64673 = ~n64668 & n64672;
  assign n64674 = n64666 & n64673;
  assign n64675 = ~n64665 & n64674;
  assign n64676 = ~n64488 & ~n64675;
  assign n64677 = n64662 & ~n64676;
  assign n64678 = ~n64653 & n64677;
  assign n64679 = ~pi1907 & ~n64678;
  assign n64680 = pi1907 & n64662;
  assign n64681 = ~n64653 & n64680;
  assign n64682 = ~n64676 & n64681;
  assign po1972 = n64679 | n64682;
  assign n64684 = ~pi6315 & pi9040;
  assign n64685 = pi6314 & ~pi9040;
  assign n64686 = ~n64684 & ~n64685;
  assign n64687 = ~pi1855 & ~n64686;
  assign n64688 = pi1855 & n64686;
  assign n64689 = ~n64687 & ~n64688;
  assign n64690 = pi6260 & ~pi9040;
  assign n64691 = pi6322 & pi9040;
  assign n64692 = ~n64690 & ~n64691;
  assign n64693 = pi1883 & n64692;
  assign n64694 = ~pi1883 & ~n64692;
  assign n64695 = ~n64693 & ~n64694;
  assign n64696 = pi6402 & ~pi9040;
  assign n64697 = pi6395 & pi9040;
  assign n64698 = ~n64696 & ~n64697;
  assign n64699 = ~pi1882 & ~n64698;
  assign n64700 = pi1882 & n64698;
  assign n64701 = ~n64699 & ~n64700;
  assign n64702 = pi6277 & ~pi9040;
  assign n64703 = pi6375 & pi9040;
  assign n64704 = ~n64702 & ~n64703;
  assign n64705 = pi1856 & n64704;
  assign n64706 = ~pi1856 & ~n64704;
  assign n64707 = ~n64705 & ~n64706;
  assign n64708 = pi6467 & pi9040;
  assign n64709 = pi6293 & ~pi9040;
  assign n64710 = ~n64708 & ~n64709;
  assign n64711 = ~pi1879 & ~n64710;
  assign n64712 = pi1879 & n64710;
  assign n64713 = ~n64711 & ~n64712;
  assign n64714 = n64707 & ~n64713;
  assign n64715 = n64701 & n64714;
  assign n64716 = n64695 & n64715;
  assign n64717 = pi6396 & ~pi9040;
  assign n64718 = pi6277 & pi9040;
  assign n64719 = ~n64717 & ~n64718;
  assign n64720 = ~pi1876 & n64719;
  assign n64721 = pi1876 & ~n64719;
  assign n64722 = ~n64720 & ~n64721;
  assign n64723 = n64701 & n64713;
  assign n64724 = n64707 & n64723;
  assign n64725 = ~n64701 & ~n64707;
  assign n64726 = ~n64707 & ~n64713;
  assign n64727 = ~n64695 & n64726;
  assign n64728 = ~n64701 & ~n64713;
  assign n64729 = n64695 & n64728;
  assign n64730 = ~n64727 & ~n64729;
  assign n64731 = ~n64725 & n64730;
  assign n64732 = ~n64724 & n64731;
  assign n64733 = ~n64722 & ~n64732;
  assign n64734 = ~n64695 & n64707;
  assign n64735 = n64713 & n64734;
  assign n64736 = ~n64701 & n64734;
  assign n64737 = ~n64707 & n64723;
  assign n64738 = ~n64736 & ~n64737;
  assign n64739 = n64722 & ~n64738;
  assign n64740 = ~n64735 & ~n64739;
  assign n64741 = ~n64733 & n64740;
  assign n64742 = ~n64716 & n64741;
  assign n64743 = n64689 & ~n64742;
  assign n64744 = ~n64701 & n64713;
  assign n64745 = ~n64707 & n64744;
  assign n64746 = ~n64695 & n64745;
  assign n64747 = n64695 & ~n64707;
  assign n64748 = ~n64713 & n64747;
  assign n64749 = ~n64701 & n64748;
  assign n64750 = ~n64716 & ~n64749;
  assign n64751 = ~n64746 & n64750;
  assign n64752 = ~n64722 & ~n64751;
  assign n64753 = ~n64743 & ~n64752;
  assign n64754 = ~n64695 & n64724;
  assign n64755 = n64701 & ~n64707;
  assign n64756 = n64722 & n64755;
  assign n64757 = n64695 & n64756;
  assign n64758 = n64707 & n64744;
  assign n64759 = n64695 & n64758;
  assign n64760 = n64714 & ~n64722;
  assign n64761 = ~n64695 & n64760;
  assign n64762 = ~n64759 & ~n64761;
  assign n64763 = ~n64701 & n64707;
  assign n64764 = n64695 & n64763;
  assign n64765 = n64701 & ~n64713;
  assign n64766 = ~n64707 & n64765;
  assign n64767 = ~n64764 & ~n64766;
  assign n64768 = n64722 & ~n64767;
  assign n64769 = n64722 & n64725;
  assign n64770 = ~n64695 & n64769;
  assign n64771 = ~n64768 & ~n64770;
  assign n64772 = n64762 & n64771;
  assign n64773 = ~n64689 & ~n64772;
  assign n64774 = ~n64757 & ~n64773;
  assign n64775 = ~n64754 & n64774;
  assign n64776 = n64753 & n64775;
  assign n64777 = ~pi1895 & ~n64776;
  assign n64778 = ~n64743 & ~n64754;
  assign n64779 = ~n64752 & n64778;
  assign n64780 = n64774 & n64779;
  assign n64781 = pi1895 & n64780;
  assign po1973 = n64777 | n64781;
  assign n64783 = pi6263 & pi9040;
  assign n64784 = pi6533 & ~pi9040;
  assign n64785 = ~n64783 & ~n64784;
  assign n64786 = ~pi1874 & ~n64785;
  assign n64787 = pi1874 & n64785;
  assign n64788 = ~n64786 & ~n64787;
  assign n64789 = pi6295 & pi9040;
  assign n64790 = pi6382 & ~pi9040;
  assign n64791 = ~n64789 & ~n64790;
  assign n64792 = pi1873 & n64791;
  assign n64793 = ~pi1873 & ~n64791;
  assign n64794 = ~n64792 & ~n64793;
  assign n64795 = pi6282 & ~pi9040;
  assign n64796 = pi6533 & pi9040;
  assign n64797 = ~n64795 & ~n64796;
  assign n64798 = ~pi1881 & ~n64797;
  assign n64799 = pi1881 & n64797;
  assign n64800 = ~n64798 & ~n64799;
  assign n64801 = pi6367 & pi9040;
  assign n64802 = pi6531 & ~pi9040;
  assign n64803 = ~n64801 & ~n64802;
  assign n64804 = ~pi1843 & n64803;
  assign n64805 = pi1843 & ~n64803;
  assign n64806 = ~n64804 & ~n64805;
  assign n64807 = ~n64800 & ~n64806;
  assign n64808 = pi6306 & ~pi9040;
  assign n64809 = pi6287 & pi9040;
  assign n64810 = ~n64808 & ~n64809;
  assign n64811 = ~pi1858 & n64810;
  assign n64812 = pi1858 & ~n64810;
  assign n64813 = ~n64811 & ~n64812;
  assign n64814 = pi6319 & ~pi9040;
  assign n64815 = pi6306 & pi9040;
  assign n64816 = ~n64814 & ~n64815;
  assign n64817 = pi1878 & n64816;
  assign n64818 = ~pi1878 & ~n64816;
  assign n64819 = ~n64817 & ~n64818;
  assign n64820 = ~n64813 & n64819;
  assign n64821 = n64807 & n64820;
  assign n64822 = n64794 & n64821;
  assign n64823 = n64813 & n64819;
  assign n64824 = n64800 & ~n64806;
  assign n64825 = n64823 & n64824;
  assign n64826 = n64800 & n64806;
  assign n64827 = n64794 & n64826;
  assign n64828 = n64819 & n64827;
  assign n64829 = ~n64813 & n64828;
  assign n64830 = n64794 & n64813;
  assign n64831 = n64806 & n64830;
  assign n64832 = ~n64800 & n64831;
  assign n64833 = ~n64829 & ~n64832;
  assign n64834 = ~n64825 & n64833;
  assign n64835 = ~n64822 & n64834;
  assign n64836 = ~n64794 & n64813;
  assign n64837 = ~n64806 & n64836;
  assign n64838 = n64800 & n64837;
  assign n64839 = n64835 & ~n64838;
  assign n64840 = ~n64788 & ~n64839;
  assign n64841 = n64794 & n64800;
  assign n64842 = ~n64806 & n64841;
  assign n64843 = ~n64813 & n64842;
  assign n64844 = ~n64831 & ~n64843;
  assign n64845 = ~n64794 & n64807;
  assign n64846 = ~n64813 & n64845;
  assign n64847 = n64844 & ~n64846;
  assign n64848 = ~n64819 & ~n64847;
  assign n64849 = ~n64794 & n64806;
  assign n64850 = n64800 & n64849;
  assign n64851 = ~n64819 & n64850;
  assign n64852 = ~n64813 & n64851;
  assign n64853 = ~n64800 & n64830;
  assign n64854 = ~n64800 & n64806;
  assign n64855 = n64813 & n64854;
  assign n64856 = ~n64853 & ~n64855;
  assign n64857 = ~n64819 & ~n64856;
  assign n64858 = ~n64852 & ~n64857;
  assign n64859 = ~n64788 & ~n64858;
  assign n64860 = ~n64848 & ~n64859;
  assign n64861 = ~n64840 & n64860;
  assign n64862 = ~n64794 & ~n64813;
  assign n64863 = n64819 & n64862;
  assign n64864 = n64854 & n64863;
  assign n64865 = ~n64794 & n64800;
  assign n64866 = n64823 & n64865;
  assign n64867 = n64813 & n64850;
  assign n64868 = n64794 & ~n64819;
  assign n64869 = n64800 & n64868;
  assign n64870 = ~n64800 & ~n64813;
  assign n64871 = ~n64794 & n64870;
  assign n64872 = ~n64869 & ~n64871;
  assign n64873 = ~n64867 & n64872;
  assign n64874 = ~n64845 & n64873;
  assign n64875 = n64807 & n64819;
  assign n64876 = n64813 & n64875;
  assign n64877 = ~n64813 & n64854;
  assign n64878 = ~n64794 & ~n64806;
  assign n64879 = ~n64877 & ~n64878;
  assign n64880 = n64819 & ~n64879;
  assign n64881 = ~n64876 & ~n64880;
  assign n64882 = n64874 & n64881;
  assign n64883 = n64788 & ~n64882;
  assign n64884 = ~n64866 & ~n64883;
  assign n64885 = ~n64864 & n64884;
  assign n64886 = n64861 & n64885;
  assign n64887 = pi1897 & n64886;
  assign n64888 = ~pi1897 & ~n64886;
  assign po1977 = n64887 | n64888;
  assign n64890 = pi6270 & pi9040;
  assign n64891 = ~pi6315 & ~pi9040;
  assign n64892 = ~n64890 & ~n64891;
  assign n64893 = pi1857 & n64892;
  assign n64894 = ~pi1857 & ~n64892;
  assign n64895 = ~n64893 & ~n64894;
  assign n64896 = pi6260 & pi9040;
  assign n64897 = pi6466 & ~pi9040;
  assign n64898 = ~n64896 & ~n64897;
  assign n64899 = ~pi1885 & n64898;
  assign n64900 = pi1885 & ~n64898;
  assign n64901 = ~n64899 & ~n64900;
  assign n64902 = pi6288 & ~pi9040;
  assign n64903 = pi6261 & pi9040;
  assign n64904 = ~n64902 & ~n64903;
  assign n64905 = pi1864 & n64904;
  assign n64906 = ~pi1864 & ~n64904;
  assign n64907 = ~n64905 & ~n64906;
  assign n64908 = n64901 & n64907;
  assign n64909 = pi6375 & ~pi9040;
  assign n64910 = pi6271 & pi9040;
  assign n64911 = ~n64909 & ~n64910;
  assign n64912 = pi1862 & n64911;
  assign n64913 = ~pi1862 & ~n64911;
  assign n64914 = ~n64912 & ~n64913;
  assign n64915 = pi6290 & pi9040;
  assign n64916 = pi6395 & ~pi9040;
  assign n64917 = ~n64915 & ~n64916;
  assign n64918 = pi1880 & n64917;
  assign n64919 = ~pi1880 & ~n64917;
  assign n64920 = ~n64918 & ~n64919;
  assign n64921 = ~n64914 & ~n64920;
  assign n64922 = n64908 & n64921;
  assign n64923 = pi6270 & ~pi9040;
  assign n64924 = pi6278 & pi9040;
  assign n64925 = ~n64923 & ~n64924;
  assign n64926 = ~pi1861 & n64925;
  assign n64927 = pi1861 & ~n64925;
  assign n64928 = ~n64926 & ~n64927;
  assign n64929 = ~n64901 & n64928;
  assign n64930 = ~n64914 & n64920;
  assign n64931 = n64929 & n64930;
  assign n64932 = ~n64901 & ~n64907;
  assign n64933 = ~n64928 & n64932;
  assign n64934 = n64914 & n64928;
  assign n64935 = ~n64907 & n64934;
  assign n64936 = n64901 & n64935;
  assign n64937 = ~n64933 & ~n64936;
  assign n64938 = ~n64901 & n64907;
  assign n64939 = n64914 & n64938;
  assign n64940 = n64937 & ~n64939;
  assign n64941 = ~n64920 & ~n64940;
  assign n64942 = n64928 & n64932;
  assign n64943 = ~n64914 & n64942;
  assign n64944 = ~n64941 & ~n64943;
  assign n64945 = ~n64931 & n64944;
  assign n64946 = ~n64922 & n64945;
  assign n64947 = n64908 & ~n64928;
  assign n64948 = ~n64914 & n64947;
  assign n64949 = ~n64928 & n64938;
  assign n64950 = n64914 & n64949;
  assign n64951 = ~n64948 & ~n64950;
  assign n64952 = n64946 & n64951;
  assign n64953 = ~n64895 & ~n64952;
  assign n64954 = ~n64914 & n64928;
  assign n64955 = n64907 & n64954;
  assign n64956 = ~n64901 & n64955;
  assign n64957 = ~n64947 & ~n64956;
  assign n64958 = ~n64920 & ~n64957;
  assign n64959 = n64908 & n64934;
  assign n64960 = ~n64907 & n64954;
  assign n64961 = n64901 & n64960;
  assign n64962 = ~n64959 & ~n64961;
  assign n64963 = ~n64901 & n64934;
  assign n64964 = ~n64914 & n64949;
  assign n64965 = ~n64963 & ~n64964;
  assign n64966 = n64920 & ~n64965;
  assign n64967 = n64962 & ~n64966;
  assign n64968 = ~n64958 & n64967;
  assign n64969 = n64895 & ~n64968;
  assign n64970 = ~n64901 & ~n64928;
  assign n64971 = n64914 & n64970;
  assign n64972 = n64901 & ~n64928;
  assign n64973 = ~n64914 & n64972;
  assign n64974 = ~n64971 & ~n64973;
  assign n64975 = ~n64920 & ~n64974;
  assign n64976 = n64901 & ~n64907;
  assign n64977 = ~n64928 & n64976;
  assign n64978 = n64914 & n64977;
  assign n64979 = ~n64959 & ~n64978;
  assign n64980 = ~n64942 & n64979;
  assign n64981 = n64920 & ~n64980;
  assign n64982 = ~n64975 & ~n64981;
  assign n64983 = ~n64907 & n64928;
  assign n64984 = n64920 & n64983;
  assign n64985 = ~n64914 & n64984;
  assign n64986 = n64982 & ~n64985;
  assign n64987 = ~n64969 & n64986;
  assign n64988 = ~n64953 & n64987;
  assign n64989 = ~pi1889 & ~n64988;
  assign n64990 = pi1889 & n64988;
  assign po1978 = n64989 | n64990;
  assign n64992 = n64451 & n64463;
  assign n64993 = ~n64457 & n64992;
  assign n64994 = ~n64463 & ~n64478;
  assign n64995 = ~n64657 & ~n64994;
  assign n64996 = ~n64469 & ~n64995;
  assign n64997 = ~n64993 & ~n64996;
  assign n64998 = n64469 & n64490;
  assign n64999 = ~n64463 & n64998;
  assign n65000 = ~n64463 & n64501;
  assign n65001 = ~n64999 & ~n65000;
  assign n65002 = n64997 & n65001;
  assign n65003 = ~n64488 & ~n65002;
  assign n65004 = ~n64493 & ~n64530;
  assign n65005 = ~n64463 & n64509;
  assign n65006 = n65004 & ~n65005;
  assign n65007 = n64469 & ~n65006;
  assign n65008 = n64490 & n64525;
  assign n65009 = ~n64481 & ~n65008;
  assign n65010 = ~n65007 & n65009;
  assign n65011 = ~n64501 & ~n64511;
  assign n65012 = ~n64469 & ~n65011;
  assign n65013 = n65010 & ~n65012;
  assign n65014 = n64488 & ~n65013;
  assign n65015 = ~n65003 & ~n65014;
  assign n65016 = n64463 & n64506;
  assign n65017 = ~n64463 & ~n64500;
  assign n65018 = ~n65016 & ~n65017;
  assign n65019 = ~n64469 & n65018;
  assign n65020 = n64463 & n64469;
  assign n65021 = ~n64493 & n64644;
  assign n65022 = n65020 & ~n65021;
  assign n65023 = ~n65019 & ~n65022;
  assign n65024 = n65015 & n65023;
  assign n65025 = ~pi1898 & ~n65024;
  assign n65026 = pi1898 & n65023;
  assign n65027 = ~n65014 & n65026;
  assign n65028 = ~n65003 & n65027;
  assign po1980 = n65025 | n65028;
  assign n65030 = ~n64463 & ~n64520;
  assign n65031 = n64457 & ~n64478;
  assign n65032 = ~n64492 & ~n65031;
  assign n65033 = n64463 & n65032;
  assign n65034 = ~n65030 & ~n65033;
  assign n65035 = ~n64654 & ~n65034;
  assign n65036 = ~n64469 & ~n65035;
  assign n65037 = n64463 & n64496;
  assign n65038 = ~n64505 & ~n65037;
  assign n65039 = ~n64481 & n65038;
  assign n65040 = n64469 & ~n65039;
  assign n65041 = ~n65036 & ~n65040;
  assign n65042 = ~n64488 & ~n65041;
  assign n65043 = n64470 & ~n64478;
  assign n65044 = ~n64667 & ~n65037;
  assign n65045 = ~n64469 & ~n65044;
  assign n65046 = ~n64526 & ~n65045;
  assign n65047 = ~n64530 & ~n64658;
  assign n65048 = n64528 & n65020;
  assign n65049 = ~n64665 & ~n65048;
  assign n65050 = n65047 & n65049;
  assign n65051 = n65046 & n65050;
  assign n65052 = ~n65043 & n65051;
  assign n65053 = n64488 & ~n65052;
  assign n65054 = ~n64469 & n64515;
  assign n65055 = ~n64463 & n65054;
  assign n65056 = ~n64659 & ~n65055;
  assign n65057 = ~n64661 & n65056;
  assign n65058 = n64463 & n64490;
  assign n65059 = ~n65000 & ~n65058;
  assign n65060 = n64469 & ~n65059;
  assign n65061 = n65057 & ~n65060;
  assign n65062 = ~n65053 & n65061;
  assign n65063 = ~n65042 & n65062;
  assign n65064 = ~pi1890 & n65063;
  assign n65065 = pi1890 & ~n65063;
  assign po1983 = n65064 | n65065;
  assign n65067 = n64794 & ~n64800;
  assign n65068 = ~n64838 & ~n65067;
  assign n65069 = ~n64870 & n65068;
  assign n65070 = n64819 & ~n65069;
  assign n65071 = ~n64813 & ~n64819;
  assign n65072 = n64800 & n65071;
  assign n65073 = n64794 & ~n64813;
  assign n65074 = ~n64806 & n65073;
  assign n65075 = n64813 & n64827;
  assign n65076 = ~n65074 & ~n65075;
  assign n65077 = ~n64794 & ~n64800;
  assign n65078 = n64813 & ~n64819;
  assign n65079 = n65077 & n65078;
  assign n65080 = n65076 & ~n65079;
  assign n65081 = ~n65072 & n65080;
  assign n65082 = ~n65070 & n65081;
  assign n65083 = n64788 & ~n65082;
  assign n65084 = n64794 & n64807;
  assign n65085 = n64813 & n65084;
  assign n65086 = n64794 & n64854;
  assign n65087 = ~n64813 & n65086;
  assign n65088 = ~n65085 & ~n65087;
  assign n65089 = n64819 & ~n65088;
  assign n65090 = ~n65083 & ~n65089;
  assign n65091 = ~n64813 & n64827;
  assign n65092 = ~n64842 & ~n64850;
  assign n65093 = n64819 & ~n65092;
  assign n65094 = ~n65091 & ~n65093;
  assign n65095 = ~n64846 & n65094;
  assign n65096 = ~n64788 & ~n65095;
  assign n65097 = ~n64824 & ~n64854;
  assign n65098 = ~n64794 & ~n65097;
  assign n65099 = ~n64855 & ~n65098;
  assign n65100 = ~n64819 & ~n65099;
  assign n65101 = ~n64788 & n65100;
  assign n65102 = ~n65096 & ~n65101;
  assign n65103 = n65090 & n65102;
  assign n65104 = pi1905 & ~n65103;
  assign n65105 = ~pi1905 & n65102;
  assign n65106 = n65090 & n65105;
  assign po1984 = n65104 | n65106;
  assign n65108 = pi6367 & ~pi9040;
  assign n65109 = pi6309 & pi9040;
  assign n65110 = ~n65108 & ~n65109;
  assign n65111 = ~pi1884 & ~n65110;
  assign n65112 = pi1884 & n65110;
  assign n65113 = ~n65111 & ~n65112;
  assign n65114 = pi6282 & pi9040;
  assign n65115 = pi6401 & ~pi9040;
  assign n65116 = ~n65114 & ~n65115;
  assign n65117 = ~pi1872 & n65116;
  assign n65118 = pi1872 & ~n65116;
  assign n65119 = ~n65117 & ~n65118;
  assign n65120 = pi6308 & pi9040;
  assign n65121 = pi6309 & ~pi9040;
  assign n65122 = ~n65120 & ~n65121;
  assign n65123 = ~pi1875 & n65122;
  assign n65124 = pi1875 & ~n65122;
  assign n65125 = ~n65123 & ~n65124;
  assign n65126 = pi6292 & ~pi9040;
  assign n65127 = pi6382 & pi9040;
  assign n65128 = ~n65126 & ~n65127;
  assign n65129 = ~pi1856 & n65128;
  assign n65130 = pi1856 & ~n65128;
  assign n65131 = ~n65129 & ~n65130;
  assign n65132 = pi6263 & ~pi9040;
  assign n65133 = pi6535 & pi9040;
  assign n65134 = ~n65132 & ~n65133;
  assign n65135 = ~pi1860 & ~n65134;
  assign n65136 = pi1860 & n65134;
  assign n65137 = ~n65135 & ~n65136;
  assign n65138 = n65131 & ~n65137;
  assign n65139 = n65125 & n65138;
  assign n65140 = n65119 & n65139;
  assign n65141 = ~n65119 & n65125;
  assign n65142 = n65131 & n65141;
  assign n65143 = n65137 & n65142;
  assign n65144 = ~n65140 & ~n65143;
  assign n65145 = n65113 & ~n65144;
  assign n65146 = pi6312 & pi9040;
  assign n65147 = pi6284 & ~pi9040;
  assign n65148 = ~n65146 & ~n65147;
  assign n65149 = ~pi1882 & ~n65148;
  assign n65150 = pi1882 & n65148;
  assign n65151 = ~n65149 & ~n65150;
  assign n65152 = n65119 & ~n65125;
  assign n65153 = ~n65131 & n65152;
  assign n65154 = ~n65137 & n65153;
  assign n65155 = n65131 & n65137;
  assign n65156 = ~n65125 & n65155;
  assign n65157 = n65113 & n65156;
  assign n65158 = ~n65154 & ~n65157;
  assign n65159 = ~n65125 & n65137;
  assign n65160 = ~n65131 & n65159;
  assign n65161 = ~n65119 & n65160;
  assign n65162 = ~n65113 & ~n65119;
  assign n65163 = n65138 & n65162;
  assign n65164 = n65125 & n65163;
  assign n65165 = n65119 & n65137;
  assign n65166 = n65125 & n65165;
  assign n65167 = ~n65137 & n65152;
  assign n65168 = ~n65166 & ~n65167;
  assign n65169 = ~n65113 & ~n65168;
  assign n65170 = n65113 & n65125;
  assign n65171 = ~n65131 & n65170;
  assign n65172 = ~n65137 & n65171;
  assign n65173 = ~n65169 & ~n65172;
  assign n65174 = ~n65164 & n65173;
  assign n65175 = ~n65161 & n65174;
  assign n65176 = n65158 & n65175;
  assign n65177 = n65151 & ~n65176;
  assign n65178 = ~n65113 & n65154;
  assign n65179 = n65119 & n65157;
  assign n65180 = ~n65178 & ~n65179;
  assign n65181 = ~n65177 & n65180;
  assign n65182 = ~n65145 & n65181;
  assign n65183 = n65113 & ~n65119;
  assign n65184 = ~n65125 & ~n65137;
  assign n65185 = n65183 & n65184;
  assign n65186 = n65113 & n65139;
  assign n65187 = ~n65185 & ~n65186;
  assign n65188 = ~n65131 & n65137;
  assign n65189 = ~n65125 & n65188;
  assign n65190 = n65113 & n65189;
  assign n65191 = n65125 & n65188;
  assign n65192 = n65119 & n65191;
  assign n65193 = ~n65190 & ~n65192;
  assign n65194 = ~n65125 & n65138;
  assign n65195 = ~n65119 & n65194;
  assign n65196 = ~n65140 & ~n65195;
  assign n65197 = ~n65119 & n65155;
  assign n65198 = n65125 & ~n65131;
  assign n65199 = ~n65197 & ~n65198;
  assign n65200 = ~n65113 & ~n65199;
  assign n65201 = n65196 & ~n65200;
  assign n65202 = n65193 & n65201;
  assign n65203 = n65187 & n65202;
  assign n65204 = ~n65151 & ~n65203;
  assign n65205 = n65182 & ~n65204;
  assign n65206 = ~pi1892 & ~n65205;
  assign n65207 = pi1892 & n65182;
  assign n65208 = ~n65204 & n65207;
  assign po1985 = n65206 | n65208;
  assign n65210 = pi6272 & pi9040;
  assign n65211 = pi6281 & ~pi9040;
  assign n65212 = ~n65210 & ~n65211;
  assign n65213 = ~pi1868 & ~n65212;
  assign n65214 = pi1868 & n65212;
  assign n65215 = ~n65213 & ~n65214;
  assign n65216 = pi6289 & ~pi9040;
  assign n65217 = pi6292 & pi9040;
  assign n65218 = ~n65216 & ~n65217;
  assign n65219 = pi1886 & n65218;
  assign n65220 = ~pi1886 & ~n65218;
  assign n65221 = ~n65219 & ~n65220;
  assign n65222 = pi6281 & pi9040;
  assign n65223 = pi6307 & ~pi9040;
  assign n65224 = ~n65222 & ~n65223;
  assign n65225 = pi1877 & n65224;
  assign n65226 = ~pi1877 & ~n65224;
  assign n65227 = ~n65225 & ~n65226;
  assign n65228 = n65221 & ~n65227;
  assign n65229 = pi6535 & ~pi9040;
  assign n65230 = pi6268 & pi9040;
  assign n65231 = ~n65229 & ~n65230;
  assign n65232 = pi1874 & n65231;
  assign n65233 = ~pi1874 & ~n65231;
  assign n65234 = ~n65232 & ~n65233;
  assign n65235 = pi6374 & ~pi9040;
  assign n65236 = pi6285 & pi9040;
  assign n65237 = ~n65235 & ~n65236;
  assign n65238 = ~pi1869 & n65237;
  assign n65239 = pi1869 & ~n65237;
  assign n65240 = ~n65238 & ~n65239;
  assign n65241 = ~n65234 & n65240;
  assign n65242 = pi6289 & pi9040;
  assign n65243 = pi6312 & ~pi9040;
  assign n65244 = ~n65242 & ~n65243;
  assign n65245 = pi1843 & n65244;
  assign n65246 = ~pi1843 & ~n65244;
  assign n65247 = ~n65245 & ~n65246;
  assign n65248 = n65234 & ~n65240;
  assign n65249 = ~n65247 & n65248;
  assign n65250 = ~n65241 & ~n65249;
  assign n65251 = n65228 & ~n65250;
  assign n65252 = ~n65227 & ~n65247;
  assign n65253 = n65241 & n65252;
  assign n65254 = ~n65251 & ~n65253;
  assign n65255 = n65215 & ~n65254;
  assign n65256 = ~n65221 & n65247;
  assign n65257 = ~n65240 & n65256;
  assign n65258 = n65234 & n65257;
  assign n65259 = n65234 & n65247;
  assign n65260 = ~n65256 & ~n65259;
  assign n65261 = n65227 & ~n65260;
  assign n65262 = ~n65221 & ~n65247;
  assign n65263 = n65240 & n65262;
  assign n65264 = n65234 & n65263;
  assign n65265 = ~n65261 & ~n65264;
  assign n65266 = ~n65258 & n65265;
  assign n65267 = n65215 & ~n65266;
  assign n65268 = ~n65255 & ~n65267;
  assign n65269 = n65221 & n65247;
  assign n65270 = ~n65240 & n65269;
  assign n65271 = ~n65234 & n65270;
  assign n65272 = ~n65234 & ~n65240;
  assign n65273 = ~n65247 & n65272;
  assign n65274 = ~n65221 & n65273;
  assign n65275 = ~n65271 & ~n65274;
  assign n65276 = ~n65227 & ~n65275;
  assign n65277 = n65241 & ~n65247;
  assign n65278 = n65221 & n65277;
  assign n65279 = ~n65221 & n65259;
  assign n65280 = ~n65278 & ~n65279;
  assign n65281 = n65227 & ~n65280;
  assign n65282 = n65234 & n65240;
  assign n65283 = ~n65259 & ~n65282;
  assign n65284 = n65221 & ~n65283;
  assign n65285 = ~n65273 & ~n65284;
  assign n65286 = ~n65227 & ~n65285;
  assign n65287 = ~n65221 & ~n65240;
  assign n65288 = n65252 & n65287;
  assign n65289 = n65240 & n65247;
  assign n65290 = ~n65273 & ~n65289;
  assign n65291 = ~n65221 & ~n65290;
  assign n65292 = n65221 & n65227;
  assign n65293 = n65248 & n65292;
  assign n65294 = ~n65247 & n65293;
  assign n65295 = ~n65291 & ~n65294;
  assign n65296 = ~n65288 & n65295;
  assign n65297 = ~n65286 & n65296;
  assign n65298 = ~n65271 & n65297;
  assign n65299 = ~n65215 & ~n65298;
  assign n65300 = ~n65281 & ~n65299;
  assign n65301 = ~n65276 & n65300;
  assign n65302 = n65268 & n65301;
  assign n65303 = pi1910 & n65302;
  assign n65304 = ~pi1910 & ~n65302;
  assign po1986 = n65303 | n65304;
  assign n65306 = ~n65179 & ~n65185;
  assign n65307 = ~n65131 & ~n65137;
  assign n65308 = n65113 & n65307;
  assign n65309 = n65119 & n65308;
  assign n65310 = n65125 & n65155;
  assign n65311 = n65137 & n65141;
  assign n65312 = ~n65310 & ~n65311;
  assign n65313 = n65113 & ~n65312;
  assign n65314 = ~n65309 & ~n65313;
  assign n65315 = ~n65113 & n65188;
  assign n65316 = n65119 & n65315;
  assign n65317 = ~n65113 & n65139;
  assign n65318 = ~n65316 & ~n65317;
  assign n65319 = n65314 & n65318;
  assign n65320 = n65137 & n65152;
  assign n65321 = ~n65140 & ~n65320;
  assign n65322 = ~n65195 & n65321;
  assign n65323 = n65319 & n65322;
  assign n65324 = ~n65151 & ~n65323;
  assign n65325 = ~n65154 & ~n65310;
  assign n65326 = ~n65197 & n65325;
  assign n65327 = ~n65113 & ~n65326;
  assign n65328 = ~n65131 & n65141;
  assign n65329 = ~n65137 & n65328;
  assign n65330 = ~n65161 & ~n65329;
  assign n65331 = n65113 & n65119;
  assign n65332 = n65191 & n65331;
  assign n65333 = n65330 & ~n65332;
  assign n65334 = n65113 & n65194;
  assign n65335 = n65333 & ~n65334;
  assign n65336 = ~n65327 & n65335;
  assign n65337 = n65151 & ~n65336;
  assign n65338 = ~n65140 & n65330;
  assign n65339 = ~n65113 & ~n65338;
  assign n65340 = ~n65337 & ~n65339;
  assign n65341 = ~n65324 & n65340;
  assign n65342 = n65306 & n65341;
  assign n65343 = pi1899 & ~n65342;
  assign n65344 = ~pi1899 & n65342;
  assign po1987 = n65343 | n65344;
  assign n65346 = ~n65125 & n65307;
  assign n65347 = ~n65119 & n65346;
  assign n65348 = ~n65119 & n65188;
  assign n65349 = n65125 & n65307;
  assign n65350 = n65119 & n65349;
  assign n65351 = ~n65348 & ~n65350;
  assign n65352 = ~n65113 & ~n65351;
  assign n65353 = ~n65347 & ~n65352;
  assign n65354 = ~n65119 & n65308;
  assign n65355 = ~n65186 & ~n65354;
  assign n65356 = n65353 & n65355;
  assign n65357 = ~n65119 & n65156;
  assign n65358 = n65119 & n65194;
  assign n65359 = ~n65357 & ~n65358;
  assign n65360 = n65356 & n65359;
  assign n65361 = n65151 & ~n65360;
  assign n65362 = ~n65113 & ~n65151;
  assign n65363 = ~n65137 & n65141;
  assign n65364 = n65125 & n65131;
  assign n65365 = ~n65363 & ~n65364;
  assign n65366 = n65362 & ~n65365;
  assign n65367 = ~n65154 & ~n65166;
  assign n65368 = ~n65125 & n65183;
  assign n65369 = ~n65307 & n65368;
  assign n65370 = ~n65157 & ~n65369;
  assign n65371 = n65367 & n65370;
  assign n65372 = ~n65151 & ~n65371;
  assign n65373 = ~n65113 & n65310;
  assign n65374 = n65119 & n65373;
  assign n65375 = n65119 & n65189;
  assign n65376 = ~n65358 & ~n65375;
  assign n65377 = ~n65113 & ~n65376;
  assign n65378 = ~n65374 & ~n65377;
  assign n65379 = n65113 & n65154;
  assign n65380 = n65378 & ~n65379;
  assign n65381 = ~n65372 & n65380;
  assign n65382 = ~n65366 & n65381;
  assign n65383 = ~n65361 & n65382;
  assign n65384 = ~n65332 & n65383;
  assign n65385 = ~pi1894 & ~n65384;
  assign n65386 = pi1894 & ~n65332;
  assign n65387 = n65383 & n65386;
  assign po1988 = n65385 | n65387;
  assign n65389 = n65269 & n65282;
  assign n65390 = n65221 & ~n65247;
  assign n65391 = ~n65234 & n65390;
  assign n65392 = ~n65389 & ~n65391;
  assign n65393 = ~n65227 & ~n65392;
  assign n65394 = ~n65221 & n65227;
  assign n65395 = n65234 & n65394;
  assign n65396 = ~n65247 & n65282;
  assign n65397 = n65247 & n65248;
  assign n65398 = ~n65396 & ~n65397;
  assign n65399 = n65241 & n65247;
  assign n65400 = n65221 & n65399;
  assign n65401 = n65398 & ~n65400;
  assign n65402 = n65227 & ~n65401;
  assign n65403 = ~n65395 & ~n65402;
  assign n65404 = n65221 & n65273;
  assign n65405 = n65403 & ~n65404;
  assign n65406 = ~n65221 & n65241;
  assign n65407 = n65247 & n65272;
  assign n65408 = ~n65406 & ~n65407;
  assign n65409 = ~n65227 & ~n65408;
  assign n65410 = ~n65221 & n65249;
  assign n65411 = ~n65409 & ~n65410;
  assign n65412 = n65405 & n65411;
  assign n65413 = n65215 & ~n65412;
  assign n65414 = ~n65393 & ~n65413;
  assign n65415 = ~n65215 & n65227;
  assign n65416 = ~n65408 & n65415;
  assign n65417 = ~n65249 & ~n65277;
  assign n65418 = n65221 & ~n65417;
  assign n65419 = ~n65389 & ~n65418;
  assign n65420 = ~n65215 & ~n65419;
  assign n65421 = ~n65416 & ~n65420;
  assign n65422 = ~n65215 & ~n65227;
  assign n65423 = ~n65221 & n65282;
  assign n65424 = ~n65273 & ~n65423;
  assign n65425 = ~n65259 & n65424;
  assign n65426 = n65422 & ~n65425;
  assign n65427 = n65421 & ~n65426;
  assign n65428 = n65414 & n65427;
  assign n65429 = ~pi1896 & ~n65428;
  assign n65430 = pi1896 & n65421;
  assign n65431 = n65414 & n65430;
  assign n65432 = ~n65426 & n65431;
  assign po1989 = n65429 | n65432;
  assign n65434 = ~n64695 & n64722;
  assign n65435 = n64701 & n65434;
  assign n65436 = n64707 & n64728;
  assign n65437 = n64695 & n65436;
  assign n65438 = n64744 & n64747;
  assign n65439 = ~n65437 & ~n65438;
  assign n65440 = ~n64695 & ~n64707;
  assign n65441 = ~n64713 & n65440;
  assign n65442 = ~n64701 & n65441;
  assign n65443 = ~n64737 & ~n65442;
  assign n65444 = ~n64722 & ~n65443;
  assign n65445 = n65439 & ~n65444;
  assign n65446 = ~n65435 & n65445;
  assign n65447 = n64689 & ~n65446;
  assign n65448 = n64695 & n64766;
  assign n65449 = n64722 & n65448;
  assign n65450 = ~n64695 & ~n64722;
  assign n65451 = n64766 & n65450;
  assign n65452 = ~n64736 & ~n65451;
  assign n65453 = ~n64737 & ~n64758;
  assign n65454 = ~n64695 & n64744;
  assign n65455 = n65453 & ~n65454;
  assign n65456 = n64722 & ~n65455;
  assign n65457 = ~n64722 & n64724;
  assign n65458 = n64750 & ~n65457;
  assign n65459 = ~n65456 & n65458;
  assign n65460 = n65452 & n65459;
  assign n65461 = ~n64689 & ~n65460;
  assign n65462 = ~n65449 & ~n65461;
  assign n65463 = ~n65447 & n65462;
  assign n65464 = n64758 & n65450;
  assign n65465 = n64695 & n64760;
  assign n65466 = ~n65464 & ~n65465;
  assign n65467 = ~n64722 & n65438;
  assign n65468 = n65466 & ~n65467;
  assign n65469 = n65463 & n65468;
  assign n65470 = ~pi1901 & ~n65469;
  assign n65471 = pi1901 & n65468;
  assign n65472 = n65462 & n65471;
  assign n65473 = ~n65447 & n65472;
  assign po1990 = n65470 | n65473;
  assign n65475 = pi6280 & ~pi9040;
  assign n65476 = pi6401 & pi9040;
  assign n65477 = ~n65475 & ~n65476;
  assign n65478 = ~pi1871 & n65477;
  assign n65479 = pi1871 & ~n65477;
  assign n65480 = ~n65478 & ~n65479;
  assign n65481 = pi6295 & ~pi9040;
  assign n65482 = pi6368 & pi9040;
  assign n65483 = ~n65481 & ~n65482;
  assign n65484 = pi1854 & n65483;
  assign n65485 = ~pi1854 & ~n65483;
  assign n65486 = ~n65484 & ~n65485;
  assign n65487 = pi6313 & ~pi9040;
  assign n65488 = pi6374 & pi9040;
  assign n65489 = ~n65487 & ~n65488;
  assign n65490 = pi1868 & n65489;
  assign n65491 = ~pi1868 & ~n65489;
  assign n65492 = ~n65490 & ~n65491;
  assign n65493 = pi6368 & ~pi9040;
  assign n65494 = pi6307 & pi9040;
  assign n65495 = ~n65493 & ~n65494;
  assign n65496 = pi1869 & n65495;
  assign n65497 = ~pi1869 & ~n65495;
  assign n65498 = ~n65496 & ~n65497;
  assign n65499 = n65492 & ~n65498;
  assign n65500 = ~n65486 & n65499;
  assign n65501 = ~n65480 & n65500;
  assign n65502 = pi6284 & pi9040;
  assign n65503 = pi6287 & ~pi9040;
  assign n65504 = ~n65502 & ~n65503;
  assign n65505 = ~pi1860 & n65504;
  assign n65506 = pi1860 & ~n65504;
  assign n65507 = ~n65505 & ~n65506;
  assign n65508 = pi6272 & ~pi9040;
  assign n65509 = pi6313 & pi9040;
  assign n65510 = ~n65508 & ~n65509;
  assign n65511 = ~pi1875 & n65510;
  assign n65512 = pi1875 & ~n65510;
  assign n65513 = ~n65511 & ~n65512;
  assign n65514 = n65492 & ~n65513;
  assign n65515 = n65498 & n65514;
  assign n65516 = ~n65492 & ~n65513;
  assign n65517 = ~n65498 & n65516;
  assign n65518 = ~n65492 & n65513;
  assign n65519 = n65480 & n65518;
  assign n65520 = ~n65517 & ~n65519;
  assign n65521 = ~n65515 & n65520;
  assign n65522 = ~n65486 & ~n65521;
  assign n65523 = n65498 & n65516;
  assign n65524 = ~n65498 & n65514;
  assign n65525 = ~n65523 & ~n65524;
  assign n65526 = n65486 & ~n65525;
  assign n65527 = ~n65522 & ~n65526;
  assign n65528 = n65492 & n65513;
  assign n65529 = n65498 & n65528;
  assign n65530 = n65486 & n65529;
  assign n65531 = ~n65498 & n65519;
  assign n65532 = ~n65530 & ~n65531;
  assign n65533 = n65527 & n65532;
  assign n65534 = n65507 & ~n65533;
  assign n65535 = ~n65480 & n65523;
  assign n65536 = n65480 & n65528;
  assign n65537 = ~n65480 & n65518;
  assign n65538 = ~n65536 & ~n65537;
  assign n65539 = ~n65486 & ~n65538;
  assign n65540 = ~n65535 & ~n65539;
  assign n65541 = n65498 & n65518;
  assign n65542 = n65486 & n65541;
  assign n65543 = ~n65498 & n65528;
  assign n65544 = ~n65515 & ~n65543;
  assign n65545 = ~n65542 & n65544;
  assign n65546 = ~n65517 & n65545;
  assign n65547 = n65480 & ~n65546;
  assign n65548 = n65540 & ~n65547;
  assign n65549 = ~n65507 & ~n65548;
  assign n65550 = ~n65534 & ~n65549;
  assign n65551 = ~n65501 & n65550;
  assign n65552 = ~n65480 & n65498;
  assign n65553 = n65513 & n65552;
  assign n65554 = n65492 & n65553;
  assign n65555 = ~n65498 & n65537;
  assign n65556 = ~n65554 & ~n65555;
  assign n65557 = n65486 & ~n65556;
  assign n65558 = n65551 & ~n65557;
  assign n65559 = ~pi1918 & ~n65558;
  assign n65560 = pi1918 & ~n65557;
  assign n65561 = n65550 & n65560;
  assign n65562 = ~n65501 & n65561;
  assign po1991 = n65559 | n65562;
  assign n65564 = n64914 & n64942;
  assign n65565 = ~n64961 & ~n64970;
  assign n65566 = n64920 & ~n65565;
  assign n65567 = ~n65564 & ~n65566;
  assign n65568 = ~n64956 & n65567;
  assign n65569 = ~n64920 & n64959;
  assign n65570 = ~n64948 & ~n65569;
  assign n65571 = ~n64978 & n65570;
  assign n65572 = n65568 & n65571;
  assign n65573 = n64895 & ~n65572;
  assign n65574 = n64928 & n64938;
  assign n65575 = n64914 & n65574;
  assign n65576 = ~n64936 & ~n65575;
  assign n65577 = ~n64914 & n64977;
  assign n65578 = n64907 & ~n64928;
  assign n65579 = ~n64901 & n64914;
  assign n65580 = ~n65578 & ~n65579;
  assign n65581 = ~n64983 & n65580;
  assign n65582 = ~n64920 & ~n65581;
  assign n65583 = n64908 & n64928;
  assign n65584 = n64920 & n65583;
  assign n65585 = ~n64943 & ~n65584;
  assign n65586 = n64914 & n64947;
  assign n65587 = n65585 & ~n65586;
  assign n65588 = ~n65582 & n65587;
  assign n65589 = ~n65577 & n65588;
  assign n65590 = n65576 & n65589;
  assign n65591 = ~n64895 & ~n65590;
  assign n65592 = ~n65573 & ~n65591;
  assign n65593 = pi1893 & ~n65592;
  assign n65594 = ~pi1893 & ~n65573;
  assign n65595 = ~n65591 & n65594;
  assign po1992 = n65593 | n65595;
  assign n65597 = n65240 & n65390;
  assign n65598 = ~n65249 & ~n65597;
  assign n65599 = ~n65227 & ~n65598;
  assign n65600 = n65221 & n65272;
  assign n65601 = ~n65263 & ~n65600;
  assign n65602 = n65227 & ~n65601;
  assign n65603 = ~n65221 & n65399;
  assign n65604 = ~n65288 & ~n65603;
  assign n65605 = ~n65389 & n65604;
  assign n65606 = ~n65602 & n65605;
  assign n65607 = ~n65599 & n65606;
  assign n65608 = ~n65258 & ~n65271;
  assign n65609 = n65607 & n65608;
  assign n65610 = n65215 & ~n65609;
  assign n65611 = n65256 & n65282;
  assign n65612 = n65417 & ~n65611;
  assign n65613 = n65227 & ~n65612;
  assign n65614 = ~n65221 & n65407;
  assign n65615 = ~n65613 & ~n65614;
  assign n65616 = n65234 & n65390;
  assign n65617 = n65221 & n65248;
  assign n65618 = ~n65616 & ~n65617;
  assign n65619 = n65227 & ~n65618;
  assign n65620 = n65227 & n65272;
  assign n65621 = ~n65221 & n65620;
  assign n65622 = ~n65619 & ~n65621;
  assign n65623 = n65615 & n65622;
  assign n65624 = ~n65215 & ~n65623;
  assign n65625 = ~n65399 & ~n65404;
  assign n65626 = ~n65264 & n65625;
  assign n65627 = n65422 & ~n65626;
  assign n65628 = ~n65624 & ~n65627;
  assign n65629 = ~n65258 & ~n65389;
  assign n65630 = ~n65227 & ~n65629;
  assign n65631 = n65628 & ~n65630;
  assign n65632 = ~n65610 & n65631;
  assign n65633 = ~pi1921 & n65632;
  assign n65634 = pi1921 & ~n65632;
  assign po1993 = n65633 | n65634;
  assign n65636 = ~n64695 & n65436;
  assign n65637 = ~n64745 & ~n64754;
  assign n65638 = n64695 & n64714;
  assign n65639 = ~n64695 & n64766;
  assign n65640 = ~n65638 & ~n65639;
  assign n65641 = n65637 & n65640;
  assign n65642 = n64722 & ~n65641;
  assign n65643 = ~n64707 & n64728;
  assign n65644 = n64695 & n64723;
  assign n65645 = ~n64736 & ~n65644;
  assign n65646 = ~n65643 & n65645;
  assign n65647 = ~n64722 & ~n65646;
  assign n65648 = n64713 & n64747;
  assign n65649 = n64701 & n65648;
  assign n65650 = ~n65647 & ~n65649;
  assign n65651 = ~n65642 & n65650;
  assign n65652 = ~n65636 & n65651;
  assign n65653 = ~n64689 & ~n65652;
  assign n65654 = n64695 & n64722;
  assign n65655 = n64724 & n65654;
  assign n65656 = n64722 & n65643;
  assign n65657 = n64722 & n64758;
  assign n65658 = ~n65656 & ~n65657;
  assign n65659 = ~n64695 & ~n65658;
  assign n65660 = ~n65655 & ~n65659;
  assign n65661 = ~n64695 & n64715;
  assign n65662 = ~n65448 & ~n65661;
  assign n65663 = n64695 & n64744;
  assign n65664 = ~n64695 & n64723;
  assign n65665 = ~n65663 & ~n65664;
  assign n65666 = ~n64715 & n65665;
  assign n65667 = ~n64745 & n65666;
  assign n65668 = ~n64722 & ~n65667;
  assign n65669 = ~n64695 & n64737;
  assign n65670 = ~n65668 & ~n65669;
  assign n65671 = n65662 & n65670;
  assign n65672 = n65660 & n65671;
  assign n65673 = n64689 & ~n65672;
  assign n65674 = n64722 & ~n65439;
  assign n65675 = ~n65673 & ~n65674;
  assign n65676 = ~n64749 & ~n65661;
  assign n65677 = ~n64722 & ~n65676;
  assign n65678 = n65675 & ~n65677;
  assign n65679 = ~n65653 & n65678;
  assign n65680 = pi1911 & ~n65679;
  assign n65681 = ~pi1911 & n65679;
  assign po1994 = n65680 | n65681;
  assign n65683 = n64813 & n64845;
  assign n65684 = ~n65075 & ~n65683;
  assign n65685 = ~n64819 & ~n65684;
  assign n65686 = n64842 & n65071;
  assign n65687 = ~n65685 & ~n65686;
  assign n65688 = ~n64866 & n65687;
  assign n65689 = n64794 & n64819;
  assign n65690 = n64806 & n65689;
  assign n65691 = ~n64800 & n65690;
  assign n65692 = n64813 & n65691;
  assign n65693 = n64819 & n65084;
  assign n65694 = ~n64838 & ~n64864;
  assign n65695 = ~n64829 & n65694;
  assign n65696 = ~n65693 & n65695;
  assign n65697 = n64788 & ~n65696;
  assign n65698 = ~n64813 & n64875;
  assign n65699 = ~n65691 & ~n65698;
  assign n65700 = ~n65074 & n65699;
  assign n65701 = n64806 & n64836;
  assign n65702 = ~n64813 & n64824;
  assign n65703 = ~n64841 & ~n65702;
  assign n65704 = ~n64819 & ~n65703;
  assign n65705 = ~n65701 & ~n65704;
  assign n65706 = n65700 & n65705;
  assign n65707 = ~n64788 & ~n65706;
  assign n65708 = ~n64813 & n64850;
  assign n65709 = ~n64845 & ~n65708;
  assign n65710 = ~n65086 & n65709;
  assign n65711 = ~n64819 & ~n65710;
  assign n65712 = n64788 & n65711;
  assign n65713 = ~n65707 & ~n65712;
  assign n65714 = ~n65697 & n65713;
  assign n65715 = ~n65692 & n65714;
  assign n65716 = n65688 & n65715;
  assign n65717 = pi1913 & ~n65716;
  assign n65718 = ~pi1913 & n65688;
  assign n65719 = n65715 & n65718;
  assign po1995 = n65717 | n65719;
  assign n65721 = n65480 & n65498;
  assign n65722 = ~n65513 & n65721;
  assign n65723 = n65544 & ~n65722;
  assign n65724 = ~n65486 & ~n65507;
  assign n65725 = ~n65723 & n65724;
  assign n65726 = ~n65507 & n65541;
  assign n65727 = ~n65480 & n65726;
  assign n65728 = ~n65498 & ~n65513;
  assign n65729 = ~n65480 & n65516;
  assign n65730 = ~n65728 & ~n65729;
  assign n65731 = n65486 & ~n65730;
  assign n65732 = ~n65530 & ~n65731;
  assign n65733 = ~n65507 & ~n65732;
  assign n65734 = ~n65727 & ~n65733;
  assign n65735 = ~n65480 & ~n65498;
  assign n65736 = ~n65513 & n65735;
  assign n65737 = ~n65531 & ~n65736;
  assign n65738 = n65486 & ~n65737;
  assign n65739 = n65734 & ~n65738;
  assign n65740 = ~n65480 & ~n65486;
  assign n65741 = n65516 & n65740;
  assign n65742 = n65498 & n65741;
  assign n65743 = ~n65514 & ~n65518;
  assign n65744 = n65735 & ~n65743;
  assign n65745 = ~n65742 & ~n65744;
  assign n65746 = ~n65554 & n65745;
  assign n65747 = n65721 & ~n65743;
  assign n65748 = n65480 & n65543;
  assign n65749 = ~n65747 & ~n65748;
  assign n65750 = n65486 & n65721;
  assign n65751 = ~n65492 & n65750;
  assign n65752 = ~n65486 & n65517;
  assign n65753 = n65480 & n65752;
  assign n65754 = ~n65751 & ~n65753;
  assign n65755 = n65749 & n65754;
  assign n65756 = n65746 & n65755;
  assign n65757 = n65507 & ~n65756;
  assign n65758 = n65739 & ~n65757;
  assign n65759 = ~n65725 & n65758;
  assign n65760 = ~pi1916 & ~n65759;
  assign n65761 = pi1916 & n65739;
  assign n65762 = ~n65725 & n65761;
  assign n65763 = ~n65757 & n65762;
  assign po1997 = n65760 | n65763;
  assign n65765 = ~n64813 & n65098;
  assign n65766 = ~n64849 & ~n65084;
  assign n65767 = ~n64819 & ~n65766;
  assign n65768 = ~n65765 & ~n65767;
  assign n65769 = n64806 & n65073;
  assign n65770 = ~n64878 & ~n65769;
  assign n65771 = ~n65086 & n65770;
  assign n65772 = n64819 & ~n65771;
  assign n65773 = n65768 & ~n65772;
  assign n65774 = n64813 & n64842;
  assign n65775 = n65773 & ~n65774;
  assign n65776 = ~n64788 & ~n65775;
  assign n65777 = n64823 & ~n65766;
  assign n65778 = ~n64845 & ~n64850;
  assign n65779 = ~n64842 & ~n65086;
  assign n65780 = n65778 & n65779;
  assign n65781 = ~n64813 & ~n65780;
  assign n65782 = ~n65777 & ~n65781;
  assign n65783 = ~n65075 & n65782;
  assign n65784 = n64788 & ~n65783;
  assign n65785 = ~n65776 & ~n65784;
  assign n65786 = ~n64813 & n65084;
  assign n65787 = ~n65774 & ~n65786;
  assign n65788 = ~n64819 & ~n65787;
  assign n65789 = n65785 & ~n65788;
  assign n65790 = pi1917 & ~n65789;
  assign n65791 = ~pi1917 & ~n65788;
  assign n65792 = ~n65784 & n65791;
  assign n65793 = ~n65776 & n65792;
  assign po1998 = n65790 | n65793;
  assign n65795 = n65486 & n65523;
  assign n65796 = n65480 & n65795;
  assign n65797 = n65480 & n65486;
  assign n65798 = n65528 & n65797;
  assign n65799 = ~n65498 & n65798;
  assign n65800 = ~n65796 & ~n65799;
  assign n65801 = ~n65748 & ~n65753;
  assign n65802 = n65492 & n65498;
  assign n65803 = ~n65480 & n65802;
  assign n65804 = ~n65729 & ~n65803;
  assign n65805 = n65486 & ~n65804;
  assign n65806 = n65480 & ~n65498;
  assign n65807 = ~n65486 & ~n65806;
  assign n65808 = ~n65743 & n65807;
  assign n65809 = ~n65516 & n65797;
  assign n65810 = ~n65498 & n65809;
  assign n65811 = ~n65808 & ~n65810;
  assign n65812 = ~n65805 & n65811;
  assign n65813 = n65801 & n65812;
  assign n65814 = ~n65507 & ~n65813;
  assign n65815 = n65800 & ~n65814;
  assign n65816 = ~n65486 & n65515;
  assign n65817 = ~n65480 & n65816;
  assign n65818 = ~n65486 & n65507;
  assign n65819 = ~n65529 & ~n65729;
  assign n65820 = ~n65743 & n65806;
  assign n65821 = n65819 & ~n65820;
  assign n65822 = n65818 & ~n65821;
  assign n65823 = ~n65480 & n65543;
  assign n65824 = ~n65480 & n65492;
  assign n65825 = ~n65498 & n65824;
  assign n65826 = ~n65537 & ~n65825;
  assign n65827 = n65480 & n65516;
  assign n65828 = ~n65541 & ~n65827;
  assign n65829 = n65826 & n65828;
  assign n65830 = n65486 & ~n65829;
  assign n65831 = ~n65823 & ~n65830;
  assign n65832 = n65507 & ~n65831;
  assign n65833 = ~n65822 & ~n65832;
  assign n65834 = ~n65817 & n65833;
  assign n65835 = n65815 & n65834;
  assign n65836 = pi1908 & ~n65835;
  assign n65837 = ~pi1908 & n65815;
  assign n65838 = n65834 & n65837;
  assign po1999 = n65836 | n65838;
  assign n65840 = ~n65357 & ~n65363;
  assign n65841 = n65151 & ~n65840;
  assign n65842 = ~n65153 & ~n65167;
  assign n65843 = ~n65346 & n65842;
  assign n65844 = ~n65113 & ~n65843;
  assign n65845 = n65151 & n65844;
  assign n65846 = ~n65841 & ~n65845;
  assign n65847 = n65156 & n65162;
  assign n65848 = ~n65164 & ~n65847;
  assign n65849 = ~n65166 & ~n65198;
  assign n65850 = n65113 & ~n65849;
  assign n65851 = n65151 & n65850;
  assign n65852 = n65848 & ~n65851;
  assign n65853 = n65119 & n65156;
  assign n65854 = ~n65154 & ~n65161;
  assign n65855 = n65119 & n65138;
  assign n65856 = ~n65143 & ~n65855;
  assign n65857 = n65113 & ~n65856;
  assign n65858 = n65119 & n65155;
  assign n65859 = ~n65191 & ~n65858;
  assign n65860 = ~n65113 & ~n65859;
  assign n65861 = ~n65857 & ~n65860;
  assign n65862 = n65854 & n65861;
  assign n65863 = ~n65853 & n65862;
  assign n65864 = ~n65151 & ~n65863;
  assign n65865 = ~n65195 & n65330;
  assign n65866 = n65113 & ~n65865;
  assign n65867 = ~n65864 & ~n65866;
  assign n65868 = n65852 & n65867;
  assign n65869 = n65846 & n65868;
  assign n65870 = ~pi1912 & ~n65869;
  assign n65871 = pi1912 & n65852;
  assign n65872 = n65846 & n65871;
  assign n65873 = n65867 & n65872;
  assign po2001 = n65870 | n65873;
  assign n65875 = ~n64914 & n64938;
  assign n65876 = ~n65577 & ~n65875;
  assign n65877 = n64920 & n65876;
  assign n65878 = ~n64908 & ~n64932;
  assign n65879 = ~n64928 & ~n65878;
  assign n65880 = n64914 & n64972;
  assign n65881 = n64901 & n64954;
  assign n65882 = n64914 & n64932;
  assign n65883 = ~n65881 & ~n65882;
  assign n65884 = ~n65880 & n65883;
  assign n65885 = ~n65879 & n65884;
  assign n65886 = ~n64920 & n65885;
  assign n65887 = ~n65877 & ~n65886;
  assign n65888 = n64914 & n65879;
  assign n65889 = ~n65575 & ~n65888;
  assign n65890 = ~n65887 & n65889;
  assign n65891 = n64895 & ~n65890;
  assign n65892 = n64920 & ~n65878;
  assign n65893 = ~n64914 & n65892;
  assign n65894 = ~n64949 & ~n64976;
  assign n65895 = n64914 & ~n65894;
  assign n65896 = n64920 & n65895;
  assign n65897 = n64928 & n65892;
  assign n65898 = ~n65896 & ~n65897;
  assign n65899 = ~n65893 & n65898;
  assign n65900 = ~n64895 & ~n65899;
  assign n65901 = ~n65891 & ~n65900;
  assign n65902 = ~n64920 & ~n65876;
  assign n65903 = ~n64936 & ~n65902;
  assign n65904 = ~n64895 & ~n65903;
  assign n65905 = n64920 & n64936;
  assign n65906 = ~n64920 & ~n65889;
  assign n65907 = ~n65905 & ~n65906;
  assign n65908 = ~n65904 & n65907;
  assign n65909 = n65901 & n65908;
  assign n65910 = pi1904 & ~n65909;
  assign n65911 = ~n65891 & n65908;
  assign n65912 = ~n65900 & n65911;
  assign n65913 = ~pi1904 & n65912;
  assign po2002 = n65910 | n65913;
  assign n65915 = ~n65537 & ~n65827;
  assign n65916 = n65486 & ~n65915;
  assign n65917 = ~n65799 & ~n65916;
  assign n65918 = ~n65507 & ~n65917;
  assign n65919 = ~n65499 & ~n65514;
  assign n65920 = n65480 & ~n65919;
  assign n65921 = ~n65523 & ~n65920;
  assign n65922 = ~n65486 & ~n65921;
  assign n65923 = ~n65820 & ~n65922;
  assign n65924 = ~n65480 & n65517;
  assign n65925 = n65513 & n65721;
  assign n65926 = ~n65480 & ~n65919;
  assign n65927 = ~n65925 & ~n65926;
  assign n65928 = n65486 & ~n65927;
  assign n65929 = ~n65924 & ~n65928;
  assign n65930 = n65923 & n65929;
  assign n65931 = n65507 & ~n65930;
  assign n65932 = ~n65514 & n65552;
  assign n65933 = ~n65507 & n65932;
  assign n65934 = n65514 & n65735;
  assign n65935 = n65486 & n65934;
  assign n65936 = n65498 & n65740;
  assign n65937 = n65513 & n65936;
  assign n65938 = ~n65935 & ~n65937;
  assign n65939 = ~n65933 & n65938;
  assign n65940 = ~n65541 & ~n65824;
  assign n65941 = n65724 & ~n65940;
  assign n65942 = n65939 & ~n65941;
  assign n65943 = ~n65931 & n65942;
  assign n65944 = ~n65918 & n65943;
  assign n65945 = pi1909 & ~n65944;
  assign n65946 = ~pi1909 & n65944;
  assign po2003 = n65945 | n65946;
  assign n65948 = n64550 & ~n64576;
  assign n65949 = n64597 & n65948;
  assign n65950 = ~n64568 & n65949;
  assign n65951 = n64556 & n64578;
  assign n65952 = ~n64602 & ~n65951;
  assign n65953 = n64576 & ~n65952;
  assign n65954 = ~n64562 & n64579;
  assign n65955 = ~n64556 & n64584;
  assign n65956 = ~n65954 & ~n65955;
  assign n65957 = ~n64556 & ~n64568;
  assign n65958 = n64576 & n65957;
  assign n65959 = n65956 & ~n65958;
  assign n65960 = ~n64550 & ~n65959;
  assign n65961 = ~n64576 & n64590;
  assign n65962 = n64556 & n64576;
  assign n65963 = ~n64568 & n65962;
  assign n65964 = ~n64562 & n65963;
  assign n65965 = ~n65961 & ~n65964;
  assign n65966 = n64550 & ~n65965;
  assign n65967 = ~n64576 & n64585;
  assign n65968 = ~n65966 & ~n65967;
  assign n65969 = ~n65960 & n65968;
  assign n65970 = ~n65953 & n65969;
  assign n65971 = n64614 & ~n65970;
  assign n65972 = ~n64550 & n64620;
  assign n65973 = ~n65971 & ~n65972;
  assign n65974 = ~n64576 & n64605;
  assign n65975 = n64576 & n64616;
  assign n65976 = ~n64602 & ~n65975;
  assign n65977 = ~n64550 & ~n65976;
  assign n65978 = ~n65974 & ~n65977;
  assign n65979 = ~n64568 & n65948;
  assign n65980 = ~n64562 & n65979;
  assign n65981 = n64584 & n64617;
  assign n65982 = ~n65980 & ~n65981;
  assign n65983 = n64550 & n64582;
  assign n65984 = n65982 & ~n65983;
  assign n65985 = ~n64580 & ~n64592;
  assign n65986 = ~n64630 & n65985;
  assign n65987 = n65984 & n65986;
  assign n65988 = n65978 & n65987;
  assign n65989 = ~n64614 & ~n65988;
  assign n65990 = n65973 & ~n65989;
  assign n65991 = ~n65950 & n65990;
  assign n65992 = ~pi1902 & ~n65991;
  assign n65993 = pi1902 & n65991;
  assign po2004 = n65992 | n65993;
  assign n65995 = ~n64577 & ~n64583;
  assign n65996 = n64550 & ~n65995;
  assign n65997 = ~n64637 & ~n65996;
  assign n65998 = n64556 & n64562;
  assign n65999 = ~n64550 & n65998;
  assign n66000 = n64576 & n65999;
  assign n66001 = n64576 & n64590;
  assign n66002 = ~n65998 & ~n66001;
  assign n66003 = ~n64556 & ~n64576;
  assign n66004 = ~n64562 & n66003;
  assign n66005 = n66002 & ~n66004;
  assign n66006 = ~n64550 & ~n66005;
  assign n66007 = ~n64586 & ~n66006;
  assign n66008 = ~n64614 & ~n66007;
  assign n66009 = n64550 & n64569;
  assign n66010 = n64576 & n66009;
  assign n66011 = ~n65983 & ~n66010;
  assign n66012 = ~n64614 & ~n66011;
  assign n66013 = ~n66008 & ~n66012;
  assign n66014 = ~n66000 & n66013;
  assign n66015 = ~n64602 & ~n64620;
  assign n66016 = ~n65955 & n66015;
  assign n66017 = n64550 & ~n66016;
  assign n66018 = n64578 & n66003;
  assign n66019 = ~n64605 & ~n66018;
  assign n66020 = ~n64550 & ~n66019;
  assign n66021 = ~n65954 & ~n66020;
  assign n66022 = ~n66017 & n66021;
  assign n66023 = ~n64592 & ~n64631;
  assign n66024 = n66022 & n66023;
  assign n66025 = n64614 & ~n66024;
  assign n66026 = n66014 & ~n66025;
  assign n66027 = n65997 & n66026;
  assign n66028 = ~pi1915 & ~n66027;
  assign n66029 = pi1915 & n66014;
  assign n66030 = n65997 & n66029;
  assign n66031 = ~n66025 & n66030;
  assign po2005 = n66028 | n66031;
  assign n66033 = n64914 & n65583;
  assign n66034 = n64920 & n66033;
  assign n66035 = n64954 & ~n65878;
  assign n66036 = ~n64977 & ~n66035;
  assign n66037 = ~n65575 & n66036;
  assign n66038 = ~n64920 & ~n66037;
  assign n66039 = n64914 & n64933;
  assign n66040 = ~n66038 & ~n66039;
  assign n66041 = n64928 & n64976;
  assign n66042 = ~n64914 & n65578;
  assign n66043 = ~n66041 & ~n66042;
  assign n66044 = ~n65882 & n66043;
  assign n66045 = n64920 & ~n66044;
  assign n66046 = n66040 & ~n66045;
  assign n66047 = n64895 & ~n66046;
  assign n66048 = ~n66034 & ~n66047;
  assign n66049 = ~n64964 & ~n65880;
  assign n66050 = ~n64920 & ~n66049;
  assign n66051 = ~n64950 & ~n64978;
  assign n66052 = n64914 & n64983;
  assign n66053 = ~n65578 & ~n66052;
  assign n66054 = ~n66041 & n66053;
  assign n66055 = ~n64920 & ~n66054;
  assign n66056 = ~n64914 & n64933;
  assign n66057 = ~n64914 & n64932;
  assign n66058 = ~n65574 & ~n66057;
  assign n66059 = n64920 & ~n66058;
  assign n66060 = ~n66033 & ~n66059;
  assign n66061 = ~n66056 & n66060;
  assign n66062 = ~n66055 & n66061;
  assign n66063 = n66051 & n66062;
  assign n66064 = ~n64895 & ~n66063;
  assign n66065 = ~n66050 & ~n66064;
  assign n66066 = n66048 & n66065;
  assign n66067 = pi1903 & n66066;
  assign n66068 = ~pi1903 & ~n66066;
  assign po2006 = n66067 | n66068;
  assign n66070 = ~n65442 & ~n65661;
  assign n66071 = ~n65649 & n66070;
  assign n66072 = n64722 & ~n66071;
  assign n66073 = ~n65451 & ~n65467;
  assign n66074 = ~n65448 & ~n65657;
  assign n66075 = ~n65436 & ~n65664;
  assign n66076 = ~n64722 & ~n66075;
  assign n66077 = ~n64754 & ~n66076;
  assign n66078 = n66074 & n66077;
  assign n66079 = n64689 & ~n66078;
  assign n66080 = ~n64707 & n64713;
  assign n66081 = ~n64725 & ~n66080;
  assign n66082 = n64695 & ~n66081;
  assign n66083 = ~n64715 & ~n65454;
  assign n66084 = ~n64722 & ~n66083;
  assign n66085 = n64695 & n64713;
  assign n66086 = ~n64737 & ~n66085;
  assign n66087 = ~n64728 & n66086;
  assign n66088 = n64722 & ~n66087;
  assign n66089 = ~n66084 & ~n66088;
  assign n66090 = ~n66082 & n66089;
  assign n66091 = ~n64689 & ~n66090;
  assign n66092 = ~n66079 & ~n66091;
  assign n66093 = n66073 & n66092;
  assign n66094 = ~n66072 & n66093;
  assign n66095 = ~pi1930 & ~n66094;
  assign n66096 = pi1930 & n66073;
  assign n66097 = ~n66072 & n66096;
  assign n66098 = n66092 & n66097;
  assign po2007 = n66095 | n66098;
  assign n66100 = ~n65221 & n65248;
  assign n66101 = ~n65396 & ~n66100;
  assign n66102 = ~n65227 & ~n66101;
  assign n66103 = n65227 & ~n65290;
  assign n66104 = ~n65278 & ~n66103;
  assign n66105 = ~n66102 & n66104;
  assign n66106 = n65215 & ~n66105;
  assign n66107 = ~n65227 & n65407;
  assign n66108 = ~n66106 & ~n66107;
  assign n66109 = ~n65603 & ~n65617;
  assign n66110 = n65227 & ~n66109;
  assign n66111 = n65227 & n65397;
  assign n66112 = n65221 & n65249;
  assign n66113 = ~n65227 & n65269;
  assign n66114 = ~n65262 & ~n66113;
  assign n66115 = ~n65234 & ~n66114;
  assign n66116 = ~n65263 & ~n66115;
  assign n66117 = ~n65389 & n66116;
  assign n66118 = ~n66112 & n66117;
  assign n66119 = ~n66111 & n66118;
  assign n66120 = ~n65215 & ~n66119;
  assign n66121 = ~n66110 & ~n66120;
  assign n66122 = n66108 & n66121;
  assign n66123 = pi1931 & ~n66122;
  assign n66124 = ~pi1931 & n66122;
  assign po2008 = n66123 | n66124;
  assign n66126 = ~n64631 & ~n65967;
  assign n66127 = ~n64550 & ~n66126;
  assign n66128 = ~n64614 & n64616;
  assign n66129 = n64550 & n66128;
  assign n66130 = n64562 & n66003;
  assign n66131 = ~n65957 & ~n66130;
  assign n66132 = ~n64585 & n66131;
  assign n66133 = ~n64550 & ~n66132;
  assign n66134 = ~n64576 & n64591;
  assign n66135 = ~n66133 & ~n66134;
  assign n66136 = ~n64614 & ~n66135;
  assign n66137 = ~n66129 & ~n66136;
  assign n66138 = ~n64580 & ~n64583;
  assign n66139 = ~n64576 & n65955;
  assign n66140 = ~n65975 & ~n66139;
  assign n66141 = n66138 & n66140;
  assign n66142 = n64550 & ~n66141;
  assign n66143 = n64556 & ~n64562;
  assign n66144 = n64550 & n66143;
  assign n66145 = n64576 & n66144;
  assign n66146 = ~n64576 & n65957;
  assign n66147 = ~n64583 & ~n66146;
  assign n66148 = ~n65964 & n66147;
  assign n66149 = ~n66145 & n66148;
  assign n66150 = ~n64550 & n65951;
  assign n66151 = n66149 & ~n66150;
  assign n66152 = n64614 & ~n66151;
  assign n66153 = ~n66142 & ~n66152;
  assign n66154 = n66137 & n66153;
  assign n66155 = ~n66127 & n66154;
  assign n66156 = pi1914 & n66155;
  assign n66157 = ~pi1914 & ~n66155;
  assign po2009 = n66156 | n66157;
  assign n66159 = pi6526 & pi9040;
  assign n66160 = pi6609 & ~pi9040;
  assign n66161 = ~n66159 & ~n66160;
  assign n66162 = ~pi1925 & ~n66161;
  assign n66163 = pi1925 & n66161;
  assign n66164 = ~n66162 & ~n66163;
  assign n66165 = pi6527 & pi9040;
  assign n66166 = pi6695 & ~pi9040;
  assign n66167 = ~n66165 & ~n66166;
  assign n66168 = pi1920 & n66167;
  assign n66169 = ~pi1920 & ~n66167;
  assign n66170 = ~n66168 & ~n66169;
  assign n66171 = pi6600 & pi9040;
  assign n66172 = pi6528 & ~pi9040;
  assign n66173 = ~n66171 & ~n66172;
  assign n66174 = ~pi1943 & n66173;
  assign n66175 = pi1943 & ~n66173;
  assign n66176 = ~n66174 & ~n66175;
  assign n66177 = pi6525 & pi9040;
  assign n66178 = pi6540 & ~pi9040;
  assign n66179 = ~n66177 & ~n66178;
  assign n66180 = ~pi1928 & n66179;
  assign n66181 = pi1928 & ~n66179;
  assign n66182 = ~n66180 & ~n66181;
  assign n66183 = ~n66176 & ~n66182;
  assign n66184 = ~n66170 & n66183;
  assign n66185 = pi6629 & pi9040;
  assign n66186 = pi6530 & ~pi9040;
  assign n66187 = ~n66185 & ~n66186;
  assign n66188 = pi1940 & n66187;
  assign n66189 = ~pi1940 & ~n66187;
  assign n66190 = ~n66188 & ~n66189;
  assign n66191 = n66184 & ~n66190;
  assign n66192 = n66176 & n66182;
  assign n66193 = ~n66170 & ~n66190;
  assign n66194 = n66192 & n66193;
  assign n66195 = ~n66191 & ~n66194;
  assign n66196 = n66170 & n66192;
  assign n66197 = n66190 & n66196;
  assign n66198 = ~n66176 & n66182;
  assign n66199 = ~n66170 & n66198;
  assign n66200 = n66190 & n66199;
  assign n66201 = ~n66197 & ~n66200;
  assign n66202 = n66195 & n66201;
  assign n66203 = n66164 & ~n66202;
  assign n66204 = n66176 & ~n66182;
  assign n66205 = ~n66170 & n66204;
  assign n66206 = n66190 & n66205;
  assign n66207 = ~n66199 & ~n66206;
  assign n66208 = n66164 & ~n66207;
  assign n66209 = ~n66164 & ~n66182;
  assign n66210 = ~n66190 & n66209;
  assign n66211 = n66170 & ~n66176;
  assign n66212 = n66190 & n66192;
  assign n66213 = ~n66211 & ~n66212;
  assign n66214 = ~n66164 & ~n66213;
  assign n66215 = ~n66210 & ~n66214;
  assign n66216 = n66170 & n66204;
  assign n66217 = ~n66190 & n66216;
  assign n66218 = n66215 & ~n66217;
  assign n66219 = ~n66182 & n66211;
  assign n66220 = n66190 & n66219;
  assign n66221 = n66218 & ~n66220;
  assign n66222 = ~n66208 & n66221;
  assign n66223 = pi6693 & pi9040;
  assign n66224 = pi6525 & ~pi9040;
  assign n66225 = ~n66223 & ~n66224;
  assign n66226 = ~pi1938 & ~n66225;
  assign n66227 = pi1938 & n66225;
  assign n66228 = ~n66226 & ~n66227;
  assign n66229 = ~n66222 & ~n66228;
  assign n66230 = ~n66170 & ~n66182;
  assign n66231 = ~n66164 & n66190;
  assign n66232 = n66228 & n66231;
  assign n66233 = n66230 & n66232;
  assign n66234 = n66182 & n66193;
  assign n66235 = ~n66164 & ~n66234;
  assign n66236 = n66170 & n66190;
  assign n66237 = n66176 & n66236;
  assign n66238 = ~n66183 & ~n66230;
  assign n66239 = ~n66190 & ~n66238;
  assign n66240 = n66164 & ~n66196;
  assign n66241 = ~n66239 & n66240;
  assign n66242 = ~n66237 & n66241;
  assign n66243 = ~n66235 & ~n66242;
  assign n66244 = n66170 & n66198;
  assign n66245 = n66190 & n66244;
  assign n66246 = ~n66243 & ~n66245;
  assign n66247 = n66228 & ~n66246;
  assign n66248 = ~n66233 & ~n66247;
  assign n66249 = ~n66229 & n66248;
  assign n66250 = ~n66203 & n66249;
  assign n66251 = ~n66164 & n66217;
  assign n66252 = n66250 & ~n66251;
  assign n66253 = pi1954 & ~n66252;
  assign n66254 = ~pi1954 & ~n66251;
  assign n66255 = n66249 & n66254;
  assign n66256 = ~n66203 & n66255;
  assign po2029 = n66253 | n66256;
  assign n66258 = pi6523 & pi9040;
  assign n66259 = pi6497 & ~pi9040;
  assign n66260 = ~n66258 & ~n66259;
  assign n66261 = ~pi1928 & ~n66260;
  assign n66262 = pi1928 & n66260;
  assign n66263 = ~n66261 & ~n66262;
  assign n66264 = pi6543 & pi9040;
  assign n66265 = pi6492 & ~pi9040;
  assign n66266 = ~n66264 & ~n66265;
  assign n66267 = ~pi1939 & n66266;
  assign n66268 = pi1939 & ~n66266;
  assign n66269 = ~n66267 & ~n66268;
  assign n66270 = pi6609 & pi9040;
  assign n66271 = pi6527 & ~pi9040;
  assign n66272 = ~n66270 & ~n66271;
  assign n66273 = ~pi1920 & ~n66272;
  assign n66274 = pi1920 & n66272;
  assign n66275 = ~n66273 & ~n66274;
  assign n66276 = n66269 & n66275;
  assign n66277 = pi6625 & ~pi9040;
  assign n66278 = pi6530 & pi9040;
  assign n66279 = ~n66277 & ~n66278;
  assign n66280 = pi1924 & n66279;
  assign n66281 = ~pi1924 & ~n66279;
  assign n66282 = ~n66280 & ~n66281;
  assign n66283 = pi6626 & ~pi9040;
  assign n66284 = pi6625 & pi9040;
  assign n66285 = ~n66283 & ~n66284;
  assign n66286 = pi1933 & n66285;
  assign n66287 = ~pi1933 & ~n66285;
  assign n66288 = ~n66286 & ~n66287;
  assign n66289 = ~n66282 & ~n66288;
  assign n66290 = n66276 & n66289;
  assign n66291 = pi6532 & ~pi9040;
  assign n66292 = pi6528 & pi9040;
  assign n66293 = ~n66291 & ~n66292;
  assign n66294 = ~pi1923 & n66293;
  assign n66295 = pi1923 & ~n66293;
  assign n66296 = ~n66294 & ~n66295;
  assign n66297 = ~n66269 & n66296;
  assign n66298 = ~n66282 & n66288;
  assign n66299 = n66297 & n66298;
  assign n66300 = ~n66269 & ~n66275;
  assign n66301 = ~n66296 & n66300;
  assign n66302 = n66282 & n66296;
  assign n66303 = ~n66275 & n66302;
  assign n66304 = n66269 & n66303;
  assign n66305 = ~n66301 & ~n66304;
  assign n66306 = ~n66269 & n66275;
  assign n66307 = n66282 & n66306;
  assign n66308 = n66305 & ~n66307;
  assign n66309 = ~n66288 & ~n66308;
  assign n66310 = n66296 & n66300;
  assign n66311 = ~n66282 & n66310;
  assign n66312 = ~n66309 & ~n66311;
  assign n66313 = ~n66299 & n66312;
  assign n66314 = ~n66290 & n66313;
  assign n66315 = n66276 & ~n66296;
  assign n66316 = ~n66282 & n66315;
  assign n66317 = ~n66296 & n66306;
  assign n66318 = n66282 & n66317;
  assign n66319 = ~n66316 & ~n66318;
  assign n66320 = n66314 & n66319;
  assign n66321 = ~n66263 & ~n66320;
  assign n66322 = ~n66282 & n66296;
  assign n66323 = n66275 & n66322;
  assign n66324 = ~n66269 & n66323;
  assign n66325 = ~n66315 & ~n66324;
  assign n66326 = ~n66288 & ~n66325;
  assign n66327 = n66276 & n66302;
  assign n66328 = ~n66275 & n66322;
  assign n66329 = n66269 & n66328;
  assign n66330 = ~n66327 & ~n66329;
  assign n66331 = ~n66269 & n66302;
  assign n66332 = ~n66282 & n66317;
  assign n66333 = ~n66331 & ~n66332;
  assign n66334 = n66288 & ~n66333;
  assign n66335 = n66330 & ~n66334;
  assign n66336 = ~n66326 & n66335;
  assign n66337 = n66263 & ~n66336;
  assign n66338 = ~n66269 & ~n66296;
  assign n66339 = n66282 & n66338;
  assign n66340 = n66269 & ~n66296;
  assign n66341 = ~n66282 & n66340;
  assign n66342 = ~n66339 & ~n66341;
  assign n66343 = ~n66288 & ~n66342;
  assign n66344 = n66269 & ~n66275;
  assign n66345 = ~n66296 & n66344;
  assign n66346 = n66282 & n66345;
  assign n66347 = ~n66327 & ~n66346;
  assign n66348 = ~n66310 & n66347;
  assign n66349 = n66288 & ~n66348;
  assign n66350 = ~n66343 & ~n66349;
  assign n66351 = ~n66275 & n66296;
  assign n66352 = n66288 & n66351;
  assign n66353 = ~n66282 & n66352;
  assign n66354 = n66350 & ~n66353;
  assign n66355 = ~n66337 & n66354;
  assign n66356 = ~n66321 & n66355;
  assign n66357 = ~pi1959 & ~n66356;
  assign n66358 = pi1959 & n66356;
  assign po2034 = n66357 | n66358;
  assign n66360 = pi6512 & pi9040;
  assign n66361 = pi6622 & ~pi9040;
  assign n66362 = ~n66360 & ~n66361;
  assign n66363 = ~pi1927 & ~n66362;
  assign n66364 = pi1927 & n66362;
  assign n66365 = ~n66363 & ~n66364;
  assign n66366 = pi6489 & pi9040;
  assign n66367 = pi6621 & ~pi9040;
  assign n66368 = ~n66366 & ~n66367;
  assign n66369 = pi1943 & n66368;
  assign n66370 = ~pi1943 & ~n66368;
  assign n66371 = ~n66369 & ~n66370;
  assign n66372 = pi6517 & ~pi9040;
  assign n66373 = pi6623 & pi9040;
  assign n66374 = ~n66372 & ~n66373;
  assign n66375 = ~pi1938 & ~n66374;
  assign n66376 = pi1938 & n66374;
  assign n66377 = ~n66375 & ~n66376;
  assign n66378 = pi6539 & pi9040;
  assign n66379 = pi6513 & ~pi9040;
  assign n66380 = ~n66378 & ~n66379;
  assign n66381 = ~pi1900 & n66380;
  assign n66382 = pi1900 & ~n66380;
  assign n66383 = ~n66381 & ~n66382;
  assign n66384 = ~n66377 & ~n66383;
  assign n66385 = pi6546 & pi9040;
  assign n66386 = pi6524 & ~pi9040;
  assign n66387 = ~n66385 & ~n66386;
  assign n66388 = pi1941 & n66387;
  assign n66389 = ~pi1941 & ~n66387;
  assign n66390 = ~n66388 & ~n66389;
  assign n66391 = pi6520 & ~pi9040;
  assign n66392 = pi6608 & pi9040;
  assign n66393 = ~n66391 & ~n66392;
  assign n66394 = ~pi1950 & ~n66393;
  assign n66395 = pi1950 & n66393;
  assign n66396 = ~n66394 & ~n66395;
  assign n66397 = n66390 & n66396;
  assign n66398 = n66384 & n66397;
  assign n66399 = n66371 & n66398;
  assign n66400 = ~n66390 & n66396;
  assign n66401 = n66377 & ~n66383;
  assign n66402 = n66400 & n66401;
  assign n66403 = n66377 & n66383;
  assign n66404 = n66371 & n66403;
  assign n66405 = n66396 & n66404;
  assign n66406 = n66390 & n66405;
  assign n66407 = n66371 & ~n66390;
  assign n66408 = n66383 & n66407;
  assign n66409 = ~n66377 & n66408;
  assign n66410 = ~n66406 & ~n66409;
  assign n66411 = ~n66402 & n66410;
  assign n66412 = ~n66399 & n66411;
  assign n66413 = ~n66371 & ~n66390;
  assign n66414 = ~n66383 & n66413;
  assign n66415 = n66377 & n66414;
  assign n66416 = n66412 & ~n66415;
  assign n66417 = ~n66365 & ~n66416;
  assign n66418 = n66371 & n66377;
  assign n66419 = ~n66383 & n66418;
  assign n66420 = n66390 & n66419;
  assign n66421 = ~n66408 & ~n66420;
  assign n66422 = ~n66371 & n66384;
  assign n66423 = n66390 & n66422;
  assign n66424 = n66421 & ~n66423;
  assign n66425 = ~n66396 & ~n66424;
  assign n66426 = ~n66371 & n66383;
  assign n66427 = n66377 & n66426;
  assign n66428 = ~n66396 & n66427;
  assign n66429 = n66390 & n66428;
  assign n66430 = ~n66377 & n66407;
  assign n66431 = ~n66377 & n66383;
  assign n66432 = ~n66390 & n66431;
  assign n66433 = ~n66430 & ~n66432;
  assign n66434 = ~n66396 & ~n66433;
  assign n66435 = ~n66429 & ~n66434;
  assign n66436 = ~n66365 & ~n66435;
  assign n66437 = ~n66425 & ~n66436;
  assign n66438 = ~n66417 & n66437;
  assign n66439 = ~n66371 & n66390;
  assign n66440 = n66396 & n66439;
  assign n66441 = n66431 & n66440;
  assign n66442 = ~n66371 & n66377;
  assign n66443 = n66400 & n66442;
  assign n66444 = ~n66390 & n66427;
  assign n66445 = n66371 & ~n66396;
  assign n66446 = n66377 & n66445;
  assign n66447 = ~n66377 & n66390;
  assign n66448 = ~n66371 & n66447;
  assign n66449 = ~n66446 & ~n66448;
  assign n66450 = ~n66444 & n66449;
  assign n66451 = ~n66422 & n66450;
  assign n66452 = n66384 & n66396;
  assign n66453 = ~n66390 & n66452;
  assign n66454 = n66390 & n66431;
  assign n66455 = ~n66371 & ~n66383;
  assign n66456 = ~n66454 & ~n66455;
  assign n66457 = n66396 & ~n66456;
  assign n66458 = ~n66453 & ~n66457;
  assign n66459 = n66451 & n66458;
  assign n66460 = n66365 & ~n66459;
  assign n66461 = ~n66443 & ~n66460;
  assign n66462 = ~n66441 & n66461;
  assign n66463 = n66438 & n66462;
  assign n66464 = pi1960 & n66463;
  assign n66465 = ~pi1960 & ~n66463;
  assign po2035 = n66464 | n66465;
  assign n66467 = pi6492 & pi9040;
  assign n66468 = pi6629 & ~pi9040;
  assign n66469 = ~n66467 & ~n66468;
  assign n66470 = ~pi1939 & ~n66469;
  assign n66471 = pi1939 & n66469;
  assign n66472 = ~n66470 & ~n66471;
  assign n66473 = pi6626 & pi9040;
  assign n66474 = pi6523 & ~pi9040;
  assign n66475 = ~n66473 & ~n66474;
  assign n66476 = ~pi1944 & ~n66475;
  assign n66477 = pi1944 & n66475;
  assign n66478 = ~n66476 & ~n66477;
  assign n66479 = pi6488 & ~pi9040;
  assign n66480 = pi6497 & pi9040;
  assign n66481 = ~n66479 & ~n66480;
  assign n66482 = pi1906 & n66481;
  assign n66483 = ~pi1906 & ~n66481;
  assign n66484 = ~n66482 & ~n66483;
  assign n66485 = pi6488 & pi9040;
  assign n66486 = pi6693 & ~pi9040;
  assign n66487 = ~n66485 & ~n66486;
  assign n66488 = ~pi1932 & n66487;
  assign n66489 = pi1932 & ~n66487;
  assign n66490 = ~n66488 & ~n66489;
  assign n66491 = pi6486 & pi9040;
  assign n66492 = pi6518 & ~pi9040;
  assign n66493 = ~n66491 & ~n66492;
  assign n66494 = ~pi1926 & n66493;
  assign n66495 = pi1926 & ~n66493;
  assign n66496 = ~n66494 & ~n66495;
  assign n66497 = ~n66490 & n66496;
  assign n66498 = n66484 & n66497;
  assign n66499 = pi6515 & ~pi9040;
  assign n66500 = pi6493 & pi9040;
  assign n66501 = ~n66499 & ~n66500;
  assign n66502 = ~pi1923 & n66501;
  assign n66503 = pi1923 & ~n66501;
  assign n66504 = ~n66502 & ~n66503;
  assign n66505 = ~n66496 & ~n66504;
  assign n66506 = ~n66490 & n66505;
  assign n66507 = ~n66498 & ~n66506;
  assign n66508 = ~n66484 & n66490;
  assign n66509 = n66504 & n66508;
  assign n66510 = ~n66496 & n66509;
  assign n66511 = n66507 & ~n66510;
  assign n66512 = n66478 & ~n66511;
  assign n66513 = n66490 & ~n66496;
  assign n66514 = ~n66504 & n66513;
  assign n66515 = ~n66484 & n66514;
  assign n66516 = n66496 & ~n66504;
  assign n66517 = ~n66490 & n66516;
  assign n66518 = ~n66484 & n66517;
  assign n66519 = ~n66496 & n66504;
  assign n66520 = n66490 & n66496;
  assign n66521 = ~n66519 & ~n66520;
  assign n66522 = n66484 & ~n66521;
  assign n66523 = ~n66518 & ~n66522;
  assign n66524 = ~n66515 & n66523;
  assign n66525 = ~n66478 & ~n66524;
  assign n66526 = ~n66512 & ~n66525;
  assign n66527 = n66472 & ~n66526;
  assign n66528 = n66478 & ~n66484;
  assign n66529 = n66496 & n66528;
  assign n66530 = ~n66478 & ~n66484;
  assign n66531 = n66519 & n66530;
  assign n66532 = ~n66484 & ~n66496;
  assign n66533 = ~n66490 & n66532;
  assign n66534 = ~n66498 & ~n66533;
  assign n66535 = ~n66478 & ~n66534;
  assign n66536 = ~n66531 & ~n66535;
  assign n66537 = ~n66490 & n66519;
  assign n66538 = ~n66484 & n66537;
  assign n66539 = n66484 & n66514;
  assign n66540 = ~n66538 & ~n66539;
  assign n66541 = n66478 & n66484;
  assign n66542 = n66513 & n66541;
  assign n66543 = n66490 & n66516;
  assign n66544 = n66478 & n66543;
  assign n66545 = ~n66542 & ~n66544;
  assign n66546 = n66540 & n66545;
  assign n66547 = n66536 & n66546;
  assign n66548 = ~n66529 & n66547;
  assign n66549 = ~n66472 & ~n66548;
  assign n66550 = n66496 & n66504;
  assign n66551 = n66490 & n66550;
  assign n66552 = ~n66478 & n66551;
  assign n66553 = ~n66484 & n66552;
  assign n66554 = ~n66478 & n66538;
  assign n66555 = ~n66553 & ~n66554;
  assign n66556 = ~n66504 & n66508;
  assign n66557 = n66496 & n66556;
  assign n66558 = n66478 & n66557;
  assign n66559 = n66555 & ~n66558;
  assign n66560 = ~n66484 & ~n66490;
  assign n66561 = n66504 & n66560;
  assign n66562 = n66496 & n66561;
  assign n66563 = n66484 & n66505;
  assign n66564 = ~n66562 & ~n66563;
  assign n66565 = n66478 & ~n66564;
  assign n66566 = n66559 & ~n66565;
  assign n66567 = ~n66549 & n66566;
  assign n66568 = ~n66527 & n66567;
  assign n66569 = ~pi1953 & ~n66568;
  assign n66570 = pi1953 & n66568;
  assign po2040 = n66569 | n66570;
  assign n66572 = pi6522 & ~pi9040;
  assign n66573 = pi6718 & pi9040;
  assign n66574 = ~n66572 & ~n66573;
  assign n66575 = ~pi1945 & ~n66574;
  assign n66576 = pi1945 & n66574;
  assign n66577 = ~n66575 & ~n66576;
  assign n66578 = pi6729 & pi9040;
  assign n66579 = pi6539 & ~pi9040;
  assign n66580 = ~n66578 & ~n66579;
  assign n66581 = ~pi1922 & n66580;
  assign n66582 = pi1922 & ~n66580;
  assign n66583 = ~n66581 & ~n66582;
  assign n66584 = pi6509 & pi9040;
  assign n66585 = pi6529 & ~pi9040;
  assign n66586 = ~n66584 & ~n66585;
  assign n66587 = ~pi1935 & ~n66586;
  assign n66588 = pi1935 & n66586;
  assign n66589 = ~n66587 & ~n66588;
  assign n66590 = pi6606 & pi9040;
  assign n66591 = pi6608 & ~pi9040;
  assign n66592 = ~n66590 & ~n66591;
  assign n66593 = ~pi1949 & n66592;
  assign n66594 = pi1949 & ~n66592;
  assign n66595 = ~n66593 & ~n66594;
  assign n66596 = pi6729 & ~pi9040;
  assign n66597 = pi6490 & pi9040;
  assign n66598 = ~n66596 & ~n66597;
  assign n66599 = ~pi1942 & n66598;
  assign n66600 = pi1942 & ~n66598;
  assign n66601 = ~n66599 & ~n66600;
  assign n66602 = n66595 & n66601;
  assign n66603 = ~n66589 & n66602;
  assign n66604 = n66583 & n66603;
  assign n66605 = n66595 & ~n66601;
  assign n66606 = ~n66589 & n66605;
  assign n66607 = ~n66583 & n66606;
  assign n66608 = ~n66604 & ~n66607;
  assign n66609 = n66577 & ~n66608;
  assign n66610 = ~n66595 & n66601;
  assign n66611 = n66589 & n66610;
  assign n66612 = n66583 & n66611;
  assign n66613 = ~n66577 & n66612;
  assign n66614 = pi6520 & pi9040;
  assign n66615 = pi6509 & ~pi9040;
  assign n66616 = ~n66614 & ~n66615;
  assign n66617 = ~pi1948 & ~n66616;
  assign n66618 = pi1948 & n66616;
  assign n66619 = ~n66617 & ~n66618;
  assign n66620 = ~n66583 & ~n66589;
  assign n66621 = ~n66595 & n66620;
  assign n66622 = n66577 & n66621;
  assign n66623 = ~n66612 & ~n66622;
  assign n66624 = ~n66583 & n66601;
  assign n66625 = n66595 & n66624;
  assign n66626 = n66583 & n66610;
  assign n66627 = ~n66625 & ~n66626;
  assign n66628 = ~n66577 & ~n66627;
  assign n66629 = n66583 & ~n66589;
  assign n66630 = ~n66577 & ~n66601;
  assign n66631 = n66629 & n66630;
  assign n66632 = n66595 & n66631;
  assign n66633 = ~n66595 & ~n66601;
  assign n66634 = n66589 & n66633;
  assign n66635 = ~n66583 & n66634;
  assign n66636 = n66583 & n66589;
  assign n66637 = n66595 & n66636;
  assign n66638 = n66577 & n66637;
  assign n66639 = ~n66635 & ~n66638;
  assign n66640 = ~n66632 & n66639;
  assign n66641 = ~n66628 & n66640;
  assign n66642 = n66623 & n66641;
  assign n66643 = n66619 & ~n66642;
  assign n66644 = n66601 & n66622;
  assign n66645 = ~n66643 & ~n66644;
  assign n66646 = ~n66613 & n66645;
  assign n66647 = ~n66609 & n66646;
  assign n66648 = n66577 & ~n66601;
  assign n66649 = n66583 & ~n66595;
  assign n66650 = n66648 & n66649;
  assign n66651 = n66595 & n66629;
  assign n66652 = n66577 & n66651;
  assign n66653 = ~n66650 & ~n66652;
  assign n66654 = ~n66583 & n66589;
  assign n66655 = ~n66595 & n66654;
  assign n66656 = n66577 & n66655;
  assign n66657 = n66595 & n66654;
  assign n66658 = n66601 & n66657;
  assign n66659 = ~n66656 & ~n66658;
  assign n66660 = ~n66601 & n66620;
  assign n66661 = n66589 & n66595;
  assign n66662 = ~n66660 & ~n66661;
  assign n66663 = ~n66577 & ~n66662;
  assign n66664 = ~n66595 & n66629;
  assign n66665 = ~n66601 & n66664;
  assign n66666 = ~n66604 & ~n66665;
  assign n66667 = ~n66663 & n66666;
  assign n66668 = n66659 & n66667;
  assign n66669 = n66653 & n66668;
  assign n66670 = ~n66619 & ~n66669;
  assign n66671 = n66647 & ~n66670;
  assign n66672 = ~pi1952 & ~n66671;
  assign n66673 = pi1952 & n66647;
  assign n66674 = ~n66670 & n66673;
  assign po2041 = n66672 | n66674;
  assign n66676 = n66371 & ~n66377;
  assign n66677 = ~n66415 & ~n66676;
  assign n66678 = ~n66447 & n66677;
  assign n66679 = n66396 & ~n66678;
  assign n66680 = n66390 & ~n66396;
  assign n66681 = n66377 & n66680;
  assign n66682 = n66371 & n66390;
  assign n66683 = ~n66383 & n66682;
  assign n66684 = ~n66390 & n66404;
  assign n66685 = ~n66683 & ~n66684;
  assign n66686 = ~n66371 & ~n66377;
  assign n66687 = ~n66390 & ~n66396;
  assign n66688 = n66686 & n66687;
  assign n66689 = n66685 & ~n66688;
  assign n66690 = ~n66681 & n66689;
  assign n66691 = ~n66679 & n66690;
  assign n66692 = n66365 & ~n66691;
  assign n66693 = n66371 & n66384;
  assign n66694 = ~n66390 & n66693;
  assign n66695 = n66371 & n66431;
  assign n66696 = n66390 & n66695;
  assign n66697 = ~n66694 & ~n66696;
  assign n66698 = n66396 & ~n66697;
  assign n66699 = ~n66692 & ~n66698;
  assign n66700 = n66390 & n66404;
  assign n66701 = ~n66419 & ~n66427;
  assign n66702 = n66396 & ~n66701;
  assign n66703 = ~n66700 & ~n66702;
  assign n66704 = ~n66423 & n66703;
  assign n66705 = ~n66365 & ~n66704;
  assign n66706 = ~n66401 & ~n66431;
  assign n66707 = ~n66371 & ~n66706;
  assign n66708 = ~n66432 & ~n66707;
  assign n66709 = ~n66396 & ~n66708;
  assign n66710 = ~n66365 & n66709;
  assign n66711 = ~n66705 & ~n66710;
  assign n66712 = n66699 & n66711;
  assign n66713 = pi1965 & ~n66712;
  assign n66714 = ~pi1965 & n66699;
  assign n66715 = n66711 & n66714;
  assign po2042 = n66713 | n66715;
  assign n66717 = pi6516 & ~pi9040;
  assign n66718 = pi6621 & pi9040;
  assign n66719 = ~n66717 & ~n66718;
  assign n66720 = pi1934 & n66719;
  assign n66721 = ~pi1934 & ~n66719;
  assign n66722 = ~n66720 & ~n66721;
  assign n66723 = pi6517 & pi9040;
  assign n66724 = pi6718 & ~pi9040;
  assign n66725 = ~n66723 & ~n66724;
  assign n66726 = ~pi1927 & ~n66725;
  assign n66727 = pi1927 & n66725;
  assign n66728 = ~n66726 & ~n66727;
  assign n66729 = pi6534 & pi9040;
  assign n66730 = pi6490 & ~pi9040;
  assign n66731 = ~n66729 & ~n66730;
  assign n66732 = ~pi1947 & n66731;
  assign n66733 = pi1947 & ~n66731;
  assign n66734 = ~n66732 & ~n66733;
  assign n66735 = n66728 & n66734;
  assign n66736 = pi6511 & pi9040;
  assign n66737 = pi6620 & ~pi9040;
  assign n66738 = ~n66736 & ~n66737;
  assign n66739 = ~pi1946 & ~n66738;
  assign n66740 = pi1946 & n66738;
  assign n66741 = ~n66739 & ~n66740;
  assign n66742 = pi6489 & ~pi9040;
  assign n66743 = pi6524 & pi9040;
  assign n66744 = ~n66742 & ~n66743;
  assign n66745 = ~pi1900 & n66744;
  assign n66746 = pi1900 & ~n66744;
  assign n66747 = ~n66745 & ~n66746;
  assign n66748 = n66741 & ~n66747;
  assign n66749 = n66735 & n66748;
  assign n66750 = n66741 & n66747;
  assign n66751 = ~n66728 & n66750;
  assign n66752 = ~n66749 & ~n66751;
  assign n66753 = ~n66722 & ~n66752;
  assign n66754 = pi6496 & pi9040;
  assign n66755 = pi6534 & ~pi9040;
  assign n66756 = ~n66754 & ~n66755;
  assign n66757 = ~pi1937 & ~n66756;
  assign n66758 = pi1937 & n66756;
  assign n66759 = ~n66757 & ~n66758;
  assign n66760 = n66722 & ~n66741;
  assign n66761 = n66728 & n66760;
  assign n66762 = n66735 & n66747;
  assign n66763 = n66728 & ~n66734;
  assign n66764 = ~n66747 & n66763;
  assign n66765 = ~n66762 & ~n66764;
  assign n66766 = ~n66728 & n66734;
  assign n66767 = ~n66747 & n66766;
  assign n66768 = n66741 & n66767;
  assign n66769 = n66765 & ~n66768;
  assign n66770 = n66722 & ~n66769;
  assign n66771 = ~n66761 & ~n66770;
  assign n66772 = ~n66728 & ~n66734;
  assign n66773 = n66747 & n66772;
  assign n66774 = n66741 & n66773;
  assign n66775 = n66771 & ~n66774;
  assign n66776 = ~n66741 & n66766;
  assign n66777 = ~n66747 & n66772;
  assign n66778 = ~n66776 & ~n66777;
  assign n66779 = ~n66722 & ~n66778;
  assign n66780 = n66747 & n66763;
  assign n66781 = ~n66741 & n66780;
  assign n66782 = ~n66779 & ~n66781;
  assign n66783 = n66775 & n66782;
  assign n66784 = n66759 & ~n66783;
  assign n66785 = ~n66753 & ~n66784;
  assign n66786 = n66722 & ~n66759;
  assign n66787 = ~n66778 & n66786;
  assign n66788 = n66747 & n66766;
  assign n66789 = ~n66780 & ~n66788;
  assign n66790 = n66741 & ~n66789;
  assign n66791 = ~n66749 & ~n66790;
  assign n66792 = ~n66759 & ~n66791;
  assign n66793 = ~n66787 & ~n66792;
  assign n66794 = ~n66722 & ~n66759;
  assign n66795 = n66735 & ~n66741;
  assign n66796 = ~n66773 & ~n66795;
  assign n66797 = n66728 & ~n66747;
  assign n66798 = n66796 & ~n66797;
  assign n66799 = n66794 & ~n66798;
  assign n66800 = n66793 & ~n66799;
  assign n66801 = n66785 & n66800;
  assign n66802 = ~pi1961 & ~n66801;
  assign n66803 = pi1961 & n66793;
  assign n66804 = n66785 & n66803;
  assign n66805 = ~n66799 & n66804;
  assign po2043 = n66802 | n66805;
  assign n66807 = ~n66722 & n66741;
  assign n66808 = ~n66766 & ~n66780;
  assign n66809 = n66807 & ~n66808;
  assign n66810 = ~n66722 & n66747;
  assign n66811 = n66766 & n66810;
  assign n66812 = ~n66809 & ~n66811;
  assign n66813 = n66759 & ~n66812;
  assign n66814 = ~n66741 & ~n66747;
  assign n66815 = ~n66734 & n66814;
  assign n66816 = n66728 & n66815;
  assign n66817 = ~n66797 & ~n66814;
  assign n66818 = n66722 & ~n66817;
  assign n66819 = ~n66741 & n66747;
  assign n66820 = n66734 & n66819;
  assign n66821 = n66728 & n66820;
  assign n66822 = ~n66818 & ~n66821;
  assign n66823 = ~n66816 & n66822;
  assign n66824 = n66759 & ~n66823;
  assign n66825 = ~n66813 & ~n66824;
  assign n66826 = ~n66734 & n66748;
  assign n66827 = ~n66728 & n66826;
  assign n66828 = ~n66741 & n66773;
  assign n66829 = ~n66827 & ~n66828;
  assign n66830 = ~n66722 & ~n66829;
  assign n66831 = n66741 & n66788;
  assign n66832 = ~n66741 & n66797;
  assign n66833 = ~n66831 & ~n66832;
  assign n66834 = n66722 & ~n66833;
  assign n66835 = ~n66735 & ~n66797;
  assign n66836 = n66741 & ~n66835;
  assign n66837 = ~n66773 & ~n66836;
  assign n66838 = ~n66722 & ~n66837;
  assign n66839 = ~n66734 & ~n66741;
  assign n66840 = n66810 & n66839;
  assign n66841 = n66734 & ~n66747;
  assign n66842 = ~n66773 & ~n66841;
  assign n66843 = ~n66741 & ~n66842;
  assign n66844 = n66722 & n66741;
  assign n66845 = n66763 & n66844;
  assign n66846 = n66747 & n66845;
  assign n66847 = ~n66843 & ~n66846;
  assign n66848 = ~n66840 & n66847;
  assign n66849 = ~n66838 & n66848;
  assign n66850 = ~n66827 & n66849;
  assign n66851 = ~n66759 & ~n66850;
  assign n66852 = ~n66834 & ~n66851;
  assign n66853 = ~n66830 & n66852;
  assign n66854 = n66825 & n66853;
  assign n66855 = pi1969 & n66854;
  assign n66856 = ~pi1969 & ~n66854;
  assign po2044 = n66855 | n66856;
  assign n66858 = n66282 & n66310;
  assign n66859 = ~n66329 & ~n66338;
  assign n66860 = n66288 & ~n66859;
  assign n66861 = ~n66858 & ~n66860;
  assign n66862 = ~n66324 & n66861;
  assign n66863 = ~n66288 & n66327;
  assign n66864 = ~n66316 & ~n66863;
  assign n66865 = ~n66346 & n66864;
  assign n66866 = n66862 & n66865;
  assign n66867 = n66263 & ~n66866;
  assign n66868 = n66296 & n66306;
  assign n66869 = n66282 & n66868;
  assign n66870 = ~n66304 & ~n66869;
  assign n66871 = ~n66282 & n66345;
  assign n66872 = ~n66311 & ~n66871;
  assign n66873 = n66276 & n66296;
  assign n66874 = n66288 & n66873;
  assign n66875 = n66282 & n66315;
  assign n66876 = ~n66874 & ~n66875;
  assign n66877 = n66275 & ~n66296;
  assign n66878 = ~n66269 & n66282;
  assign n66879 = ~n66877 & ~n66878;
  assign n66880 = ~n66351 & n66879;
  assign n66881 = ~n66288 & ~n66880;
  assign n66882 = n66876 & ~n66881;
  assign n66883 = n66872 & n66882;
  assign n66884 = n66870 & n66883;
  assign n66885 = ~n66263 & ~n66884;
  assign n66886 = ~n66867 & ~n66885;
  assign n66887 = pi1955 & ~n66886;
  assign n66888 = ~pi1955 & ~n66867;
  assign n66889 = ~n66885 & n66888;
  assign po2046 = n66887 | n66889;
  assign n66891 = pi6518 & pi9040;
  assign n66892 = pi6526 & ~pi9040;
  assign n66893 = ~n66891 & ~n66892;
  assign n66894 = pi1926 & n66893;
  assign n66895 = ~pi1926 & ~n66893;
  assign n66896 = ~n66894 & ~n66895;
  assign n66897 = pi6493 & ~pi9040;
  assign n66898 = pi6695 & pi9040;
  assign n66899 = ~n66897 & ~n66898;
  assign n66900 = pi1951 & n66899;
  assign n66901 = ~pi1951 & ~n66899;
  assign n66902 = ~n66900 & ~n66901;
  assign n66903 = pi6486 & ~pi9040;
  assign n66904 = pi6536 & pi9040;
  assign n66905 = ~n66903 & ~n66904;
  assign n66906 = ~pi1948 & n66905;
  assign n66907 = pi1948 & ~n66905;
  assign n66908 = ~n66906 & ~n66907;
  assign n66909 = pi6628 & pi9040;
  assign n66910 = pi6536 & ~pi9040;
  assign n66911 = ~n66909 & ~n66910;
  assign n66912 = ~pi1935 & ~n66911;
  assign n66913 = pi1935 & n66911;
  assign n66914 = ~n66912 & ~n66913;
  assign n66915 = pi6543 & ~pi9040;
  assign n66916 = pi6521 & pi9040;
  assign n66917 = ~n66915 & ~n66916;
  assign n66918 = ~pi1932 & ~n66917;
  assign n66919 = pi1932 & n66917;
  assign n66920 = ~n66918 & ~n66919;
  assign n66921 = n66914 & ~n66920;
  assign n66922 = ~n66908 & n66921;
  assign n66923 = n66902 & n66922;
  assign n66924 = ~n66902 & n66914;
  assign n66925 = n66920 & n66924;
  assign n66926 = pi6515 & pi9040;
  assign n66927 = pi6607 & ~pi9040;
  assign n66928 = ~n66926 & ~n66927;
  assign n66929 = pi1936 & n66928;
  assign n66930 = ~pi1936 & ~n66928;
  assign n66931 = ~n66929 & ~n66930;
  assign n66932 = n66908 & n66924;
  assign n66933 = ~n66908 & n66920;
  assign n66934 = ~n66914 & n66933;
  assign n66935 = ~n66932 & ~n66934;
  assign n66936 = ~n66931 & ~n66935;
  assign n66937 = ~n66925 & ~n66936;
  assign n66938 = n66914 & n66933;
  assign n66939 = n66908 & ~n66914;
  assign n66940 = ~n66914 & ~n66920;
  assign n66941 = ~n66902 & n66940;
  assign n66942 = n66908 & ~n66920;
  assign n66943 = n66902 & n66942;
  assign n66944 = ~n66941 & ~n66943;
  assign n66945 = ~n66939 & n66944;
  assign n66946 = ~n66938 & n66945;
  assign n66947 = n66931 & ~n66946;
  assign n66948 = n66937 & ~n66947;
  assign n66949 = ~n66923 & n66948;
  assign n66950 = n66896 & ~n66949;
  assign n66951 = n66908 & n66920;
  assign n66952 = ~n66914 & n66951;
  assign n66953 = ~n66902 & n66952;
  assign n66954 = ~n66914 & n66942;
  assign n66955 = n66902 & n66954;
  assign n66956 = ~n66923 & ~n66955;
  assign n66957 = ~n66953 & n66956;
  assign n66958 = n66931 & ~n66957;
  assign n66959 = ~n66950 & ~n66958;
  assign n66960 = ~n66908 & n66925;
  assign n66961 = ~n66908 & ~n66914;
  assign n66962 = ~n66931 & n66961;
  assign n66963 = n66902 & n66962;
  assign n66964 = ~n66902 & n66931;
  assign n66965 = n66914 & n66964;
  assign n66966 = ~n66920 & n66965;
  assign n66967 = n66914 & n66951;
  assign n66968 = n66902 & n66967;
  assign n66969 = ~n66966 & ~n66968;
  assign n66970 = n66908 & n66914;
  assign n66971 = n66902 & n66970;
  assign n66972 = ~n66908 & ~n66920;
  assign n66973 = ~n66914 & n66972;
  assign n66974 = ~n66971 & ~n66973;
  assign n66975 = ~n66931 & ~n66974;
  assign n66976 = ~n66931 & n66939;
  assign n66977 = ~n66902 & n66976;
  assign n66978 = ~n66975 & ~n66977;
  assign n66979 = n66969 & n66978;
  assign n66980 = ~n66896 & ~n66979;
  assign n66981 = ~n66963 & ~n66980;
  assign n66982 = ~n66960 & n66981;
  assign n66983 = n66959 & n66982;
  assign n66984 = ~pi1967 & ~n66983;
  assign n66985 = ~n66950 & ~n66960;
  assign n66986 = ~n66958 & n66985;
  assign n66987 = n66981 & n66986;
  assign n66988 = pi1967 & n66987;
  assign po2047 = n66984 | n66988;
  assign n66990 = ~n66601 & n66621;
  assign n66991 = n66601 & n66664;
  assign n66992 = ~n66990 & ~n66991;
  assign n66993 = ~n66595 & n66636;
  assign n66994 = ~n66601 & n66993;
  assign n66995 = ~n66601 & n66654;
  assign n66996 = n66601 & n66637;
  assign n66997 = ~n66995 & ~n66996;
  assign n66998 = ~n66577 & ~n66997;
  assign n66999 = ~n66994 & ~n66998;
  assign n67000 = n66577 & n66636;
  assign n67001 = ~n66601 & n67000;
  assign n67002 = ~n66652 & ~n67001;
  assign n67003 = n66999 & n67002;
  assign n67004 = n66992 & n67003;
  assign n67005 = n66619 & ~n67004;
  assign n67006 = ~n66577 & ~n66619;
  assign n67007 = n66583 & n66605;
  assign n67008 = ~n66589 & n66595;
  assign n67009 = ~n67007 & ~n67008;
  assign n67010 = n67006 & ~n67009;
  assign n67011 = ~n66612 & ~n66625;
  assign n67012 = ~n66595 & n66648;
  assign n67013 = ~n66636 & n67012;
  assign n67014 = ~n66622 & ~n67013;
  assign n67015 = n67011 & n67014;
  assign n67016 = ~n66619 & ~n67015;
  assign n67017 = n66595 & n66620;
  assign n67018 = ~n66577 & n67017;
  assign n67019 = n66601 & n67018;
  assign n67020 = n66601 & n66655;
  assign n67021 = ~n66991 & ~n67020;
  assign n67022 = ~n66577 & ~n67021;
  assign n67023 = ~n67019 & ~n67022;
  assign n67024 = n66577 & n66612;
  assign n67025 = n67023 & ~n67024;
  assign n67026 = ~n67016 & n67025;
  assign n67027 = ~n67010 & n67026;
  assign n67028 = ~n67005 & n67027;
  assign n67029 = n66577 & n66601;
  assign n67030 = n66657 & n67029;
  assign n67031 = n67028 & ~n67030;
  assign n67032 = ~pi1956 & ~n67031;
  assign n67033 = pi1956 & ~n67030;
  assign n67034 = n67027 & n67033;
  assign n67035 = ~n67005 & n67034;
  assign po2048 = n67032 | n67035;
  assign n67037 = ~n66490 & n66528;
  assign n67038 = ~n66504 & n67037;
  assign n67039 = ~n66510 & ~n67038;
  assign n67040 = ~n66472 & ~n66478;
  assign n67041 = ~n66484 & n66505;
  assign n67042 = n66484 & n66537;
  assign n67043 = ~n67041 & ~n67042;
  assign n67044 = ~n66484 & n66497;
  assign n67045 = n67043 & ~n67044;
  assign n67046 = n67040 & ~n67045;
  assign n67047 = ~n66490 & n66550;
  assign n67048 = n66484 & n67047;
  assign n67049 = ~n66509 & ~n67048;
  assign n67050 = n66490 & n66519;
  assign n67051 = ~n66506 & ~n67050;
  assign n67052 = n67049 & n67051;
  assign n67053 = n66478 & ~n67052;
  assign n67054 = n66484 & n66543;
  assign n67055 = ~n67053 & ~n67054;
  assign n67056 = ~n66472 & ~n67055;
  assign n67057 = ~n67046 & ~n67056;
  assign n67058 = ~n66505 & ~n66550;
  assign n67059 = n66484 & ~n67058;
  assign n67060 = ~n66551 & ~n67059;
  assign n67061 = ~n66478 & ~n67060;
  assign n67062 = ~n66517 & ~n67044;
  assign n67063 = ~n67042 & n67062;
  assign n67064 = n66478 & ~n67063;
  assign n67065 = ~n67061 & ~n67064;
  assign n67066 = n66484 & n66551;
  assign n67067 = ~n66539 & ~n67066;
  assign n67068 = ~n66557 & n67067;
  assign n67069 = ~n66531 & n67068;
  assign n67070 = n67065 & n67069;
  assign n67071 = n66472 & ~n67070;
  assign n67072 = n67057 & ~n67071;
  assign n67073 = n67039 & n67072;
  assign n67074 = pi1957 & ~n67073;
  assign n67075 = ~pi1957 & n67039;
  assign n67076 = n67057 & n67075;
  assign n67077 = ~n67071 & n67076;
  assign po2050 = n67074 | n67077;
  assign n67079 = ~n66390 & n66422;
  assign n67080 = ~n66684 & ~n67079;
  assign n67081 = ~n66396 & ~n67080;
  assign n67082 = n66419 & n66680;
  assign n67083 = ~n67081 & ~n67082;
  assign n67084 = ~n66443 & n67083;
  assign n67085 = n66371 & n66396;
  assign n67086 = n66383 & n67085;
  assign n67087 = ~n66377 & n67086;
  assign n67088 = ~n66390 & n67087;
  assign n67089 = n66396 & n66693;
  assign n67090 = ~n66415 & ~n66441;
  assign n67091 = ~n66406 & n67090;
  assign n67092 = ~n67089 & n67091;
  assign n67093 = n66365 & ~n67092;
  assign n67094 = n66390 & n66452;
  assign n67095 = ~n67087 & ~n67094;
  assign n67096 = ~n66683 & n67095;
  assign n67097 = n66383 & n66413;
  assign n67098 = n66390 & n66401;
  assign n67099 = ~n66418 & ~n67098;
  assign n67100 = ~n66396 & ~n67099;
  assign n67101 = ~n67097 & ~n67100;
  assign n67102 = n67096 & n67101;
  assign n67103 = ~n66365 & ~n67102;
  assign n67104 = n66390 & n66427;
  assign n67105 = ~n66422 & ~n67104;
  assign n67106 = ~n66695 & n67105;
  assign n67107 = ~n66396 & ~n67106;
  assign n67108 = n66365 & n67107;
  assign n67109 = ~n67103 & ~n67108;
  assign n67110 = ~n67093 & n67109;
  assign n67111 = ~n67088 & n67110;
  assign n67112 = n67084 & n67111;
  assign n67113 = pi1970 & ~n67112;
  assign n67114 = ~pi1970 & n67084;
  assign n67115 = n67111 & n67114;
  assign po2052 = n67113 | n67115;
  assign n67117 = ~n66902 & ~n66931;
  assign n67118 = ~n66908 & n67117;
  assign n67119 = n66914 & n66942;
  assign n67120 = n66902 & n67119;
  assign n67121 = n66902 & n66952;
  assign n67122 = ~n67120 & ~n67121;
  assign n67123 = ~n66902 & n66954;
  assign n67124 = ~n66934 & ~n67123;
  assign n67125 = n66931 & ~n67124;
  assign n67126 = n67122 & ~n67125;
  assign n67127 = ~n67118 & n67126;
  assign n67128 = n66896 & ~n67127;
  assign n67129 = n66902 & n66973;
  assign n67130 = ~n66931 & n67129;
  assign n67131 = n66964 & n66973;
  assign n67132 = ~n66932 & ~n67131;
  assign n67133 = ~n66934 & ~n66967;
  assign n67134 = ~n66902 & n66951;
  assign n67135 = n67133 & ~n67134;
  assign n67136 = ~n66931 & ~n67135;
  assign n67137 = n66931 & n66938;
  assign n67138 = n66956 & ~n67137;
  assign n67139 = ~n67136 & n67138;
  assign n67140 = n67132 & n67139;
  assign n67141 = ~n66896 & ~n67140;
  assign n67142 = ~n67130 & ~n67141;
  assign n67143 = ~n67128 & n67142;
  assign n67144 = n66964 & n66967;
  assign n67145 = n66921 & n66931;
  assign n67146 = n66902 & n67145;
  assign n67147 = ~n67144 & ~n67146;
  assign n67148 = n66931 & n67121;
  assign n67149 = n67147 & ~n67148;
  assign n67150 = n67143 & n67149;
  assign n67151 = ~pi1966 & ~n67150;
  assign n67152 = pi1966 & n67149;
  assign n67153 = n67142 & n67152;
  assign n67154 = ~n67128 & n67153;
  assign po2054 = n67151 | n67154;
  assign n67156 = n66390 & n66707;
  assign n67157 = ~n66426 & ~n66693;
  assign n67158 = ~n66396 & ~n67157;
  assign n67159 = ~n67156 & ~n67158;
  assign n67160 = n66383 & n66682;
  assign n67161 = ~n66455 & ~n67160;
  assign n67162 = ~n66695 & n67161;
  assign n67163 = n66396 & ~n67162;
  assign n67164 = n67159 & ~n67163;
  assign n67165 = ~n66390 & n66419;
  assign n67166 = n67164 & ~n67165;
  assign n67167 = ~n66365 & ~n67166;
  assign n67168 = n66400 & ~n67157;
  assign n67169 = ~n66422 & ~n66427;
  assign n67170 = ~n66419 & ~n66695;
  assign n67171 = n67169 & n67170;
  assign n67172 = n66390 & ~n67171;
  assign n67173 = ~n67168 & ~n67172;
  assign n67174 = ~n66684 & n67173;
  assign n67175 = n66365 & ~n67174;
  assign n67176 = ~n67167 & ~n67175;
  assign n67177 = n66390 & n66693;
  assign n67178 = ~n67165 & ~n67177;
  assign n67179 = ~n66396 & ~n67178;
  assign n67180 = n67176 & ~n67179;
  assign n67181 = pi1963 & ~n67180;
  assign n67182 = ~pi1963 & ~n67179;
  assign n67183 = ~n67175 & n67182;
  assign n67184 = ~n67167 & n67183;
  assign po2055 = n67181 | n67184;
  assign n67186 = n66601 & n67000;
  assign n67187 = ~n66583 & n66605;
  assign n67188 = ~n67017 & ~n67187;
  assign n67189 = n66577 & ~n67188;
  assign n67190 = ~n67186 & ~n67189;
  assign n67191 = ~n66577 & n66654;
  assign n67192 = n66601 & n67191;
  assign n67193 = ~n66577 & n66651;
  assign n67194 = ~n67192 & ~n67193;
  assign n67195 = n67190 & n67194;
  assign n67196 = ~n66583 & n66610;
  assign n67197 = ~n66604 & ~n67196;
  assign n67198 = ~n66665 & n67197;
  assign n67199 = n67195 & n67198;
  assign n67200 = ~n66619 & ~n67199;
  assign n67201 = ~n66612 & ~n67017;
  assign n67202 = ~n66660 & n67201;
  assign n67203 = ~n66577 & ~n67202;
  assign n67204 = ~n66601 & n66637;
  assign n67205 = ~n66635 & ~n67204;
  assign n67206 = ~n67030 & n67205;
  assign n67207 = n66577 & n66664;
  assign n67208 = n67206 & ~n67207;
  assign n67209 = ~n67203 & n67208;
  assign n67210 = n66619 & ~n67209;
  assign n67211 = ~n66644 & ~n66650;
  assign n67212 = ~n66604 & n67205;
  assign n67213 = ~n66577 & ~n67212;
  assign n67214 = n67211 & ~n67213;
  assign n67215 = ~n67210 & n67214;
  assign n67216 = ~n67200 & n67215;
  assign n67217 = pi1964 & ~n67216;
  assign n67218 = ~pi1964 & n67216;
  assign po2057 = n67217 | n67218;
  assign n67220 = ~n66902 & n67119;
  assign n67221 = ~n66952 & ~n66960;
  assign n67222 = n66902 & n66921;
  assign n67223 = ~n66902 & n66973;
  assign n67224 = ~n67222 & ~n67223;
  assign n67225 = n67221 & n67224;
  assign n67226 = ~n66931 & ~n67225;
  assign n67227 = n66902 & n66933;
  assign n67228 = ~n66932 & ~n67227;
  assign n67229 = ~n66954 & n67228;
  assign n67230 = n66931 & ~n67229;
  assign n67231 = n66902 & ~n66914;
  assign n67232 = n66920 & n67231;
  assign n67233 = ~n66908 & n67232;
  assign n67234 = ~n67230 & ~n67233;
  assign n67235 = ~n67226 & n67234;
  assign n67236 = ~n67220 & n67235;
  assign n67237 = ~n66896 & ~n67236;
  assign n67238 = n66902 & ~n66931;
  assign n67239 = n66938 & n67238;
  assign n67240 = ~n66931 & n66954;
  assign n67241 = ~n66931 & n66967;
  assign n67242 = ~n67240 & ~n67241;
  assign n67243 = ~n66902 & ~n67242;
  assign n67244 = ~n67239 & ~n67243;
  assign n67245 = ~n66902 & n66922;
  assign n67246 = ~n67129 & ~n67245;
  assign n67247 = n66902 & n66951;
  assign n67248 = ~n66902 & n66933;
  assign n67249 = ~n67247 & ~n67248;
  assign n67250 = ~n66922 & n67249;
  assign n67251 = ~n66952 & n67250;
  assign n67252 = n66931 & ~n67251;
  assign n67253 = ~n66902 & n66934;
  assign n67254 = ~n67252 & ~n67253;
  assign n67255 = n67246 & n67254;
  assign n67256 = n67244 & n67255;
  assign n67257 = n66896 & ~n67256;
  assign n67258 = ~n66931 & ~n67122;
  assign n67259 = ~n67257 & ~n67258;
  assign n67260 = ~n66955 & ~n67245;
  assign n67261 = n66931 & ~n67260;
  assign n67262 = n67259 & ~n67261;
  assign n67263 = ~n67237 & n67262;
  assign n67264 = pi1968 & ~n67263;
  assign n67265 = ~pi1968 & n67263;
  assign po2058 = n67264 | n67265;
  assign n67267 = ~n66990 & ~n67007;
  assign n67268 = n66619 & ~n67267;
  assign n67269 = ~n66611 & ~n66626;
  assign n67270 = ~n66993 & n67269;
  assign n67271 = ~n66577 & ~n67270;
  assign n67272 = n66619 & n67271;
  assign n67273 = ~n67268 & ~n67272;
  assign n67274 = n66621 & n66630;
  assign n67275 = ~n66632 & ~n67274;
  assign n67276 = ~n66625 & ~n66661;
  assign n67277 = n66577 & ~n67276;
  assign n67278 = n66619 & n67277;
  assign n67279 = n67275 & ~n67278;
  assign n67280 = n66601 & n66621;
  assign n67281 = n66601 & n66629;
  assign n67282 = ~n66607 & ~n67281;
  assign n67283 = n66577 & ~n67282;
  assign n67284 = ~n66612 & ~n66635;
  assign n67285 = n66601 & n66620;
  assign n67286 = ~n66657 & ~n67285;
  assign n67287 = ~n66577 & ~n67286;
  assign n67288 = n67284 & ~n67287;
  assign n67289 = ~n67283 & n67288;
  assign n67290 = ~n67280 & n67289;
  assign n67291 = ~n66619 & ~n67290;
  assign n67292 = ~n66665 & n67205;
  assign n67293 = n66577 & ~n67292;
  assign n67294 = ~n67291 & ~n67293;
  assign n67295 = n67279 & n67294;
  assign n67296 = n67273 & n67295;
  assign n67297 = ~pi1973 & ~n67296;
  assign n67298 = pi1973 & n67279;
  assign n67299 = n67273 & n67298;
  assign n67300 = n67294 & n67299;
  assign po2059 = n67297 | n67300;
  assign n67302 = ~n66484 & n66496;
  assign n67303 = ~n66561 & ~n67302;
  assign n67304 = ~n66478 & ~n67303;
  assign n67305 = n66478 & n66505;
  assign n67306 = ~n66484 & n67305;
  assign n67307 = n66484 & ~n66504;
  assign n67308 = ~n66490 & n67307;
  assign n67309 = ~n67306 & ~n67308;
  assign n67310 = ~n66562 & n67309;
  assign n67311 = ~n67304 & n67310;
  assign n67312 = n66472 & ~n67311;
  assign n67313 = ~n66537 & ~n66539;
  assign n67314 = ~n66484 & n66516;
  assign n67315 = n67313 & ~n67314;
  assign n67316 = n66478 & ~n67315;
  assign n67317 = n66505 & n66530;
  assign n67318 = ~n66510 & ~n67317;
  assign n67319 = ~n67316 & n67318;
  assign n67320 = ~n67047 & ~n67054;
  assign n67321 = ~n66478 & ~n67320;
  assign n67322 = n67319 & ~n67321;
  assign n67323 = ~n66472 & ~n67322;
  assign n67324 = ~n67312 & ~n67323;
  assign n67325 = ~n66484 & n66550;
  assign n67326 = n66484 & ~n67051;
  assign n67327 = ~n67325 & ~n67326;
  assign n67328 = ~n66478 & ~n67327;
  assign n67329 = ~n66517 & ~n66551;
  assign n67330 = ~n66537 & n67329;
  assign n67331 = n66541 & ~n67330;
  assign n67332 = ~n67328 & ~n67331;
  assign n67333 = n67324 & n67332;
  assign n67334 = ~pi1958 & ~n67333;
  assign n67335 = ~n67323 & n67332;
  assign n67336 = pi1958 & n67335;
  assign n67337 = ~n67312 & n67336;
  assign po2060 = n67334 | n67337;
  assign n67339 = n66734 & n66750;
  assign n67340 = ~n66780 & ~n67339;
  assign n67341 = ~n66722 & ~n67340;
  assign n67342 = n66741 & n66772;
  assign n67343 = ~n66820 & ~n67342;
  assign n67344 = n66722 & ~n67343;
  assign n67345 = ~n66741 & n66767;
  assign n67346 = ~n66840 & ~n67345;
  assign n67347 = ~n66749 & n67346;
  assign n67348 = ~n67344 & n67347;
  assign n67349 = ~n67341 & n67348;
  assign n67350 = ~n66816 & ~n66827;
  assign n67351 = n67349 & n67350;
  assign n67352 = n66759 & ~n67351;
  assign n67353 = n66735 & n66814;
  assign n67354 = n66789 & ~n67353;
  assign n67355 = n66722 & ~n67354;
  assign n67356 = ~n66741 & n66777;
  assign n67357 = ~n67355 & ~n67356;
  assign n67358 = n66728 & n66750;
  assign n67359 = n66741 & n66763;
  assign n67360 = ~n67358 & ~n67359;
  assign n67361 = n66722 & ~n67360;
  assign n67362 = n66722 & n66772;
  assign n67363 = ~n66741 & n67362;
  assign n67364 = ~n67361 & ~n67363;
  assign n67365 = n67357 & n67364;
  assign n67366 = ~n66759 & ~n67365;
  assign n67367 = ~n66767 & ~n66774;
  assign n67368 = ~n66821 & n67367;
  assign n67369 = n66794 & ~n67368;
  assign n67370 = ~n67366 & ~n67369;
  assign n67371 = ~n66749 & ~n66816;
  assign n67372 = ~n66722 & ~n67371;
  assign n67373 = n67370 & ~n67372;
  assign n67374 = ~n67352 & n67373;
  assign n67375 = ~pi1986 & n67374;
  assign n67376 = pi1986 & ~n67374;
  assign po2061 = n67375 | n67376;
  assign n67378 = ~n66478 & ~n67329;
  assign n67379 = n66484 & n66506;
  assign n67380 = ~n67378 & ~n67379;
  assign n67381 = n66484 & ~n66496;
  assign n67382 = ~n66513 & ~n67381;
  assign n67383 = ~n67047 & n67382;
  assign n67384 = n66478 & ~n67383;
  assign n67385 = n67380 & ~n67384;
  assign n67386 = ~n66472 & ~n67385;
  assign n67387 = ~n66478 & n66515;
  assign n67388 = ~n66554 & ~n67387;
  assign n67389 = ~n66558 & n67388;
  assign n67390 = ~n66557 & ~n66561;
  assign n67391 = n66478 & n66533;
  assign n67392 = n66484 & n66517;
  assign n67393 = ~n66478 & n66513;
  assign n67394 = ~n67392 & ~n67393;
  assign n67395 = ~n67066 & n67394;
  assign n67396 = ~n67391 & n67395;
  assign n67397 = n67390 & n67396;
  assign n67398 = ~n66544 & n67397;
  assign n67399 = n66472 & ~n67398;
  assign n67400 = n67389 & ~n67399;
  assign n67401 = ~n67386 & n67400;
  assign n67402 = ~pi1962 & ~n67401;
  assign n67403 = pi1962 & n67389;
  assign n67404 = ~n67386 & n67403;
  assign n67405 = ~n67399 & n67404;
  assign po2062 = n67402 | n67405;
  assign n67407 = ~n66282 & n66306;
  assign n67408 = ~n66871 & ~n67407;
  assign n67409 = n66288 & n67408;
  assign n67410 = n66282 & n66340;
  assign n67411 = ~n66276 & ~n66300;
  assign n67412 = ~n66296 & ~n67411;
  assign n67413 = n66269 & n66322;
  assign n67414 = n66282 & n66300;
  assign n67415 = ~n67413 & ~n67414;
  assign n67416 = ~n67412 & n67415;
  assign n67417 = ~n67410 & n67416;
  assign n67418 = ~n66288 & n67417;
  assign n67419 = ~n67409 & ~n67418;
  assign n67420 = n66282 & n67412;
  assign n67421 = ~n66869 & ~n67420;
  assign n67422 = ~n67419 & n67421;
  assign n67423 = n66263 & ~n67422;
  assign n67424 = n66288 & ~n67411;
  assign n67425 = ~n66282 & n67424;
  assign n67426 = ~n66317 & ~n66344;
  assign n67427 = n66282 & ~n67426;
  assign n67428 = n66288 & n67427;
  assign n67429 = n66296 & n67424;
  assign n67430 = ~n67428 & ~n67429;
  assign n67431 = ~n67425 & n67430;
  assign n67432 = ~n66263 & ~n67431;
  assign n67433 = ~n67423 & ~n67432;
  assign n67434 = ~n66288 & ~n67408;
  assign n67435 = ~n66304 & ~n67434;
  assign n67436 = ~n66263 & ~n67435;
  assign n67437 = n66288 & n66304;
  assign n67438 = ~n66288 & ~n67421;
  assign n67439 = ~n67437 & ~n67438;
  assign n67440 = ~n67436 & n67439;
  assign n67441 = n67433 & n67440;
  assign n67442 = pi1971 & ~n67441;
  assign n67443 = ~n67423 & n67440;
  assign n67444 = ~n67432 & n67443;
  assign n67445 = ~pi1971 & n67444;
  assign po2063 = n67442 | n67445;
  assign n67447 = ~n67123 & ~n67245;
  assign n67448 = ~n67233 & n67447;
  assign n67449 = ~n66931 & ~n67448;
  assign n67450 = ~n67129 & ~n67241;
  assign n67451 = ~n67119 & ~n67248;
  assign n67452 = n66931 & ~n67451;
  assign n67453 = ~n66960 & ~n67452;
  assign n67454 = n67450 & n67453;
  assign n67455 = n66896 & ~n67454;
  assign n67456 = ~n66914 & n66920;
  assign n67457 = ~n66939 & ~n67456;
  assign n67458 = n66902 & ~n67457;
  assign n67459 = ~n66922 & ~n67134;
  assign n67460 = n66931 & ~n67459;
  assign n67461 = n66902 & n66920;
  assign n67462 = ~n66934 & ~n67461;
  assign n67463 = ~n66942 & n67462;
  assign n67464 = ~n66931 & ~n67463;
  assign n67465 = ~n67460 & ~n67464;
  assign n67466 = ~n67458 & n67465;
  assign n67467 = ~n66896 & ~n67466;
  assign n67468 = ~n67455 & ~n67467;
  assign n67469 = ~n67131 & ~n67148;
  assign n67470 = n67468 & n67469;
  assign n67471 = ~n67449 & n67470;
  assign n67472 = ~pi1980 & ~n67471;
  assign n67473 = pi1980 & n67469;
  assign n67474 = ~n67449 & n67473;
  assign n67475 = n67468 & n67474;
  assign po2064 = n67472 | n67475;
  assign n67477 = ~n66190 & n66219;
  assign n67478 = ~n66182 & n66190;
  assign n67479 = ~n66170 & n67478;
  assign n67480 = ~n66216 & ~n67479;
  assign n67481 = n66164 & ~n67480;
  assign n67482 = ~n67477 & ~n67481;
  assign n67483 = ~n66164 & ~n66190;
  assign n67484 = ~n66182 & n67483;
  assign n67485 = ~n66176 & n67484;
  assign n67486 = n66198 & n66231;
  assign n67487 = ~n67485 & ~n67486;
  assign n67488 = ~n66164 & n66170;
  assign n67489 = n66192 & n67488;
  assign n67490 = n67487 & ~n67489;
  assign n67491 = ~n66194 & ~n66206;
  assign n67492 = n66182 & n66236;
  assign n67493 = n67491 & ~n67492;
  assign n67494 = n67490 & n67493;
  assign n67495 = n67482 & n67494;
  assign n67496 = ~n66228 & ~n67495;
  assign n67497 = ~n66170 & n66192;
  assign n67498 = ~n66216 & ~n67497;
  assign n67499 = n66190 & ~n67498;
  assign n67500 = ~n66176 & n66193;
  assign n67501 = ~n66244 & ~n67500;
  assign n67502 = n66170 & ~n66182;
  assign n67503 = n66190 & n67502;
  assign n67504 = n67501 & ~n67503;
  assign n67505 = n66164 & ~n67504;
  assign n67506 = ~n66190 & n66204;
  assign n67507 = ~n66170 & n66190;
  assign n67508 = ~n66182 & n67507;
  assign n67509 = ~n66176 & n67508;
  assign n67510 = ~n67506 & ~n67509;
  assign n67511 = ~n66164 & ~n67510;
  assign n67512 = ~n66190 & n66199;
  assign n67513 = ~n67511 & ~n67512;
  assign n67514 = ~n67505 & n67513;
  assign n67515 = ~n67499 & n67514;
  assign n67516 = n66228 & ~n67515;
  assign n67517 = n66164 & n66234;
  assign n67518 = ~n67516 & ~n67517;
  assign n67519 = n66211 & n67483;
  assign n67520 = ~n66182 & n67519;
  assign n67521 = n67518 & ~n67520;
  assign n67522 = ~n67496 & n67521;
  assign n67523 = ~pi1984 & ~n67522;
  assign n67524 = pi1984 & n67518;
  assign n67525 = ~n67496 & n67524;
  assign n67526 = ~n67520 & n67525;
  assign po2065 = n67523 | n67526;
  assign n67528 = ~n66191 & ~n66197;
  assign n67529 = ~n66164 & ~n67528;
  assign n67530 = ~n66251 & ~n67529;
  assign n67531 = ~n66170 & n66176;
  assign n67532 = n66164 & n67531;
  assign n67533 = n66190 & n67532;
  assign n67534 = n66190 & n66204;
  assign n67535 = ~n67531 & ~n67534;
  assign n67536 = n66170 & ~n66190;
  assign n67537 = ~n66176 & n67536;
  assign n67538 = n67535 & ~n67537;
  assign n67539 = n66164 & ~n67538;
  assign n67540 = ~n66200 & ~n67539;
  assign n67541 = ~n66228 & ~n67540;
  assign n67542 = ~n66164 & n66183;
  assign n67543 = n66190 & n67542;
  assign n67544 = ~n67489 & ~n67543;
  assign n67545 = ~n66228 & ~n67544;
  assign n67546 = ~n67541 & ~n67545;
  assign n67547 = ~n67533 & n67546;
  assign n67548 = ~n66216 & ~n66234;
  assign n67549 = ~n66244 & n67548;
  assign n67550 = ~n66164 & ~n67549;
  assign n67551 = ~n66190 & n66196;
  assign n67552 = ~n66219 & ~n67551;
  assign n67553 = n66164 & ~n67552;
  assign n67554 = ~n67550 & ~n67553;
  assign n67555 = ~n67500 & n67554;
  assign n67556 = ~n66206 & ~n66245;
  assign n67557 = n67555 & n67556;
  assign n67558 = n66228 & ~n67557;
  assign n67559 = n67547 & ~n67558;
  assign n67560 = n67530 & n67559;
  assign n67561 = ~pi1996 & ~n67560;
  assign n67562 = pi1996 & n67547;
  assign n67563 = n67530 & n67562;
  assign n67564 = ~n67558 & n67563;
  assign po2066 = n67561 | n67564;
  assign n67566 = n66282 & n66873;
  assign n67567 = n66288 & n67566;
  assign n67568 = n66322 & ~n67411;
  assign n67569 = ~n66345 & ~n67568;
  assign n67570 = ~n66869 & n67569;
  assign n67571 = ~n66288 & ~n67570;
  assign n67572 = n66282 & n66301;
  assign n67573 = ~n67571 & ~n67572;
  assign n67574 = n66296 & n66344;
  assign n67575 = ~n66282 & n66877;
  assign n67576 = ~n67574 & ~n67575;
  assign n67577 = ~n67414 & n67576;
  assign n67578 = n66288 & ~n67577;
  assign n67579 = n67573 & ~n67578;
  assign n67580 = n66263 & ~n67579;
  assign n67581 = ~n67567 & ~n67580;
  assign n67582 = ~n66282 & n66300;
  assign n67583 = ~n66868 & ~n67582;
  assign n67584 = n66288 & ~n67583;
  assign n67585 = ~n66346 & ~n67584;
  assign n67586 = ~n66318 & ~n67566;
  assign n67587 = ~n66282 & n66301;
  assign n67588 = n66282 & n66351;
  assign n67589 = ~n66877 & ~n67588;
  assign n67590 = ~n67574 & n67589;
  assign n67591 = ~n66288 & ~n67590;
  assign n67592 = ~n67587 & ~n67591;
  assign n67593 = n67586 & n67592;
  assign n67594 = n67585 & n67593;
  assign n67595 = ~n66263 & ~n67594;
  assign n67596 = ~n66332 & ~n67410;
  assign n67597 = ~n66288 & ~n67596;
  assign n67598 = ~n67595 & ~n67597;
  assign n67599 = n67581 & n67598;
  assign n67600 = pi1976 & n67599;
  assign n67601 = ~pi1976 & ~n67599;
  assign po2067 = n67600 | n67601;
  assign n67603 = pi6512 & ~pi9040;
  assign n67604 = pi6487 & pi9040;
  assign n67605 = ~n67603 & ~n67604;
  assign n67606 = pi1929 & n67605;
  assign n67607 = ~pi1929 & ~n67605;
  assign n67608 = ~n67606 & ~n67607;
  assign n67609 = pi6496 & ~pi9040;
  assign n67610 = pi6620 & pi9040;
  assign n67611 = ~n67609 & ~n67610;
  assign n67612 = ~pi1919 & n67611;
  assign n67613 = pi1919 & ~n67611;
  assign n67614 = ~n67612 & ~n67613;
  assign n67615 = pi6516 & pi9040;
  assign n67616 = pi6487 & ~pi9040;
  assign n67617 = ~n67615 & ~n67616;
  assign n67618 = ~pi1937 & n67617;
  assign n67619 = pi1937 & ~n67617;
  assign n67620 = ~n67618 & ~n67619;
  assign n67621 = pi6519 & ~pi9040;
  assign n67622 = pi6529 & pi9040;
  assign n67623 = ~n67621 & ~n67622;
  assign n67624 = ~pi1947 & n67623;
  assign n67625 = pi1947 & ~n67623;
  assign n67626 = ~n67624 & ~n67625;
  assign n67627 = ~n67620 & n67626;
  assign n67628 = n67614 & n67627;
  assign n67629 = n67608 & n67628;
  assign n67630 = pi6510 & pi9040;
  assign n67631 = pi6511 & ~pi9040;
  assign n67632 = ~n67630 & ~n67631;
  assign n67633 = ~pi1922 & n67632;
  assign n67634 = pi1922 & ~n67632;
  assign n67635 = ~n67633 & ~n67634;
  assign n67636 = pi6519 & pi9040;
  assign n67637 = pi6605 & ~pi9040;
  assign n67638 = ~n67636 & ~n67637;
  assign n67639 = pi1949 & n67638;
  assign n67640 = ~pi1949 & ~n67638;
  assign n67641 = ~n67639 & ~n67640;
  assign n67642 = ~n67620 & n67641;
  assign n67643 = ~n67626 & n67642;
  assign n67644 = n67620 & n67641;
  assign n67645 = n67626 & n67644;
  assign n67646 = n67620 & ~n67641;
  assign n67647 = ~n67608 & n67646;
  assign n67648 = ~n67645 & ~n67647;
  assign n67649 = ~n67643 & n67648;
  assign n67650 = n67614 & ~n67649;
  assign n67651 = ~n67626 & n67644;
  assign n67652 = n67626 & n67642;
  assign n67653 = ~n67651 & ~n67652;
  assign n67654 = ~n67614 & ~n67653;
  assign n67655 = ~n67650 & ~n67654;
  assign n67656 = ~n67620 & ~n67641;
  assign n67657 = ~n67626 & n67656;
  assign n67658 = ~n67614 & n67657;
  assign n67659 = n67626 & n67647;
  assign n67660 = ~n67658 & ~n67659;
  assign n67661 = n67655 & n67660;
  assign n67662 = n67635 & ~n67661;
  assign n67663 = n67608 & n67651;
  assign n67664 = ~n67608 & n67656;
  assign n67665 = n67608 & n67646;
  assign n67666 = ~n67664 & ~n67665;
  assign n67667 = n67614 & ~n67666;
  assign n67668 = ~n67663 & ~n67667;
  assign n67669 = ~n67626 & n67646;
  assign n67670 = ~n67614 & n67669;
  assign n67671 = n67626 & n67656;
  assign n67672 = ~n67643 & ~n67671;
  assign n67673 = ~n67670 & n67672;
  assign n67674 = ~n67645 & n67673;
  assign n67675 = ~n67608 & ~n67674;
  assign n67676 = n67668 & ~n67675;
  assign n67677 = ~n67635 & ~n67676;
  assign n67678 = ~n67662 & ~n67677;
  assign n67679 = ~n67629 & n67678;
  assign n67680 = n67608 & n67657;
  assign n67681 = n67626 & n67665;
  assign n67682 = ~n67680 & ~n67681;
  assign n67683 = ~n67614 & ~n67682;
  assign n67684 = n67679 & ~n67683;
  assign n67685 = ~pi1987 & ~n67684;
  assign n67686 = n67678 & ~n67683;
  assign n67687 = pi1987 & n67686;
  assign n67688 = ~n67629 & n67687;
  assign po2068 = n67685 | n67688;
  assign n67690 = ~n66741 & n66763;
  assign n67691 = ~n66762 & ~n67690;
  assign n67692 = ~n66722 & ~n67691;
  assign n67693 = n66722 & ~n66842;
  assign n67694 = ~n66831 & ~n67693;
  assign n67695 = ~n67692 & n67694;
  assign n67696 = n66759 & ~n67695;
  assign n67697 = ~n66722 & n66777;
  assign n67698 = ~n67696 & ~n67697;
  assign n67699 = ~n67345 & ~n67359;
  assign n67700 = n66722 & ~n67699;
  assign n67701 = n66722 & n66764;
  assign n67702 = n66741 & n66780;
  assign n67703 = ~n66722 & n66748;
  assign n67704 = ~n66819 & ~n67703;
  assign n67705 = ~n66728 & ~n67704;
  assign n67706 = ~n66820 & ~n67705;
  assign n67707 = ~n66749 & n67706;
  assign n67708 = ~n67702 & n67707;
  assign n67709 = ~n67701 & n67708;
  assign n67710 = ~n66759 & ~n67709;
  assign n67711 = ~n67700 & ~n67710;
  assign n67712 = n67698 & n67711;
  assign n67713 = pi1995 & ~n67712;
  assign n67714 = ~pi1995 & n67712;
  assign po2069 = n67713 | n67714;
  assign n67716 = ~n66245 & ~n67512;
  assign n67717 = n66164 & ~n67716;
  assign n67718 = ~n66228 & n66230;
  assign n67719 = ~n66164 & n67718;
  assign n67720 = n66176 & n67536;
  assign n67721 = ~n67502 & ~n67720;
  assign n67722 = ~n66199 & n67721;
  assign n67723 = n66164 & ~n67722;
  assign n67724 = ~n66190 & n66205;
  assign n67725 = ~n67723 & ~n67724;
  assign n67726 = ~n66228 & ~n67725;
  assign n67727 = ~n67719 & ~n67726;
  assign n67728 = ~n66194 & ~n66197;
  assign n67729 = ~n66190 & n66244;
  assign n67730 = ~n67479 & ~n67729;
  assign n67731 = n67728 & n67730;
  assign n67732 = ~n66164 & ~n67731;
  assign n67733 = ~n66170 & ~n66176;
  assign n67734 = ~n66164 & n67733;
  assign n67735 = n66190 & n67734;
  assign n67736 = ~n66190 & n67502;
  assign n67737 = ~n66197 & ~n67736;
  assign n67738 = ~n67509 & n67737;
  assign n67739 = ~n67735 & n67738;
  assign n67740 = n66164 & n67497;
  assign n67741 = n67739 & ~n67740;
  assign n67742 = n66228 & ~n67741;
  assign n67743 = ~n67732 & ~n67742;
  assign n67744 = n67727 & n67743;
  assign n67745 = ~n67717 & n67744;
  assign n67746 = pi1994 & n67745;
  assign n67747 = ~pi1994 & ~n67745;
  assign po2070 = n67746 | n67747;
  assign n67749 = ~n67614 & n67651;
  assign n67750 = ~n67608 & n67749;
  assign n67751 = ~n67608 & ~n67614;
  assign n67752 = n67656 & n67751;
  assign n67753 = n67626 & n67752;
  assign n67754 = ~n67750 & ~n67753;
  assign n67755 = ~n67608 & n67614;
  assign n67756 = n67644 & n67755;
  assign n67757 = n67626 & n67756;
  assign n67758 = ~n67608 & n67626;
  assign n67759 = ~n67620 & n67758;
  assign n67760 = ~n67641 & n67759;
  assign n67761 = ~n67757 & ~n67760;
  assign n67762 = ~n67642 & ~n67646;
  assign n67763 = n67614 & ~n67758;
  assign n67764 = ~n67762 & n67763;
  assign n67765 = ~n67620 & ~n67626;
  assign n67766 = n67608 & n67765;
  assign n67767 = n67608 & n67644;
  assign n67768 = ~n67766 & ~n67767;
  assign n67769 = ~n67614 & ~n67768;
  assign n67770 = ~n67608 & ~n67644;
  assign n67771 = ~n67614 & n67770;
  assign n67772 = n67626 & n67771;
  assign n67773 = ~n67769 & ~n67772;
  assign n67774 = ~n67764 & n67773;
  assign n67775 = n67761 & n67774;
  assign n67776 = ~n67635 & ~n67775;
  assign n67777 = n67754 & ~n67776;
  assign n67778 = n67614 & n67643;
  assign n67779 = n67608 & n67778;
  assign n67780 = n67614 & n67635;
  assign n67781 = ~n67657 & ~n67767;
  assign n67782 = n67758 & ~n67762;
  assign n67783 = n67781 & ~n67782;
  assign n67784 = n67780 & ~n67783;
  assign n67785 = n67608 & n67671;
  assign n67786 = n67608 & ~n67620;
  assign n67787 = n67626 & n67786;
  assign n67788 = ~n67665 & ~n67787;
  assign n67789 = ~n67608 & n67644;
  assign n67790 = ~n67669 & ~n67789;
  assign n67791 = n67788 & n67790;
  assign n67792 = ~n67614 & ~n67791;
  assign n67793 = ~n67785 & ~n67792;
  assign n67794 = n67635 & ~n67793;
  assign n67795 = ~n67784 & ~n67794;
  assign n67796 = ~n67779 & n67795;
  assign n67797 = n67777 & n67796;
  assign n67798 = pi1979 & ~n67797;
  assign n67799 = ~pi1979 & n67777;
  assign n67800 = n67796 & n67799;
  assign po2071 = n67798 | n67800;
  assign n67802 = ~n67608 & ~n67626;
  assign n67803 = n67641 & n67802;
  assign n67804 = n67672 & ~n67803;
  assign n67805 = n67614 & ~n67635;
  assign n67806 = ~n67804 & n67805;
  assign n67807 = ~n67635 & n67669;
  assign n67808 = n67608 & n67807;
  assign n67809 = n67626 & n67641;
  assign n67810 = ~n67767 & ~n67809;
  assign n67811 = ~n67614 & ~n67810;
  assign n67812 = ~n67658 & ~n67811;
  assign n67813 = ~n67635 & ~n67812;
  assign n67814 = ~n67808 & ~n67813;
  assign n67815 = n67608 & n67626;
  assign n67816 = n67641 & n67815;
  assign n67817 = ~n67659 & ~n67816;
  assign n67818 = ~n67614 & ~n67817;
  assign n67819 = n67814 & ~n67818;
  assign n67820 = n67608 & n67614;
  assign n67821 = n67644 & n67820;
  assign n67822 = ~n67626 & n67821;
  assign n67823 = ~n67762 & n67815;
  assign n67824 = ~n67822 & ~n67823;
  assign n67825 = ~n67680 & n67824;
  assign n67826 = ~n67762 & n67802;
  assign n67827 = ~n67760 & ~n67826;
  assign n67828 = ~n67614 & n67802;
  assign n67829 = n67620 & n67828;
  assign n67830 = ~n67757 & ~n67829;
  assign n67831 = n67827 & n67830;
  assign n67832 = n67825 & n67831;
  assign n67833 = n67635 & ~n67832;
  assign n67834 = n67819 & ~n67833;
  assign n67835 = ~n67806 & n67834;
  assign n67836 = ~pi1977 & ~n67835;
  assign n67837 = pi1977 & n67819;
  assign n67838 = ~n67806 & n67837;
  assign n67839 = ~n67833 & n67838;
  assign po2072 = n67836 | n67839;
  assign n67841 = ~n67665 & ~n67789;
  assign n67842 = ~n67614 & ~n67841;
  assign n67843 = ~n67753 & ~n67842;
  assign n67844 = ~n67635 & ~n67843;
  assign n67845 = ~n67627 & ~n67642;
  assign n67846 = ~n67608 & ~n67845;
  assign n67847 = ~n67651 & ~n67846;
  assign n67848 = n67614 & ~n67847;
  assign n67849 = ~n67782 & ~n67848;
  assign n67850 = n67608 & n67645;
  assign n67851 = ~n67641 & n67802;
  assign n67852 = n67608 & ~n67845;
  assign n67853 = ~n67851 & ~n67852;
  assign n67854 = ~n67614 & ~n67853;
  assign n67855 = ~n67850 & ~n67854;
  assign n67856 = n67849 & n67855;
  assign n67857 = n67635 & ~n67856;
  assign n67858 = n67608 & ~n67626;
  assign n67859 = ~n67642 & n67858;
  assign n67860 = ~n67635 & n67859;
  assign n67861 = ~n67614 & n67815;
  assign n67862 = n67642 & n67861;
  assign n67863 = ~n67626 & ~n67641;
  assign n67864 = n67820 & n67863;
  assign n67865 = ~n67862 & ~n67864;
  assign n67866 = ~n67860 & n67865;
  assign n67867 = ~n67669 & ~n67786;
  assign n67868 = n67805 & ~n67867;
  assign n67869 = n67866 & ~n67868;
  assign n67870 = ~n67857 & n67869;
  assign n67871 = ~n67844 & n67870;
  assign n67872 = pi1988 & ~n67871;
  assign n67873 = ~pi1988 & n67871;
  assign po2073 = n67872 | n67873;
  assign n67875 = pi6759 & ~pi9040;
  assign n67876 = pi6720 & pi9040;
  assign n67877 = ~n67875 & ~n67876;
  assign n67878 = pi1985 & n67877;
  assign n67879 = ~pi1985 & ~n67877;
  assign n67880 = ~n67878 & ~n67879;
  assign n67881 = pi6724 & pi9040;
  assign n67882 = pi6779 & ~pi9040;
  assign n67883 = ~n67881 & ~n67882;
  assign n67884 = pi1972 & n67883;
  assign n67885 = ~pi1972 & ~n67883;
  assign n67886 = ~n67884 & ~n67885;
  assign n67887 = pi6758 & pi9040;
  assign n67888 = pi6725 & ~pi9040;
  assign n67889 = ~n67887 & ~n67888;
  assign n67890 = ~pi2003 & n67889;
  assign n67891 = pi2003 & ~n67889;
  assign n67892 = ~n67890 & ~n67891;
  assign n67893 = pi6761 & ~pi9040;
  assign n67894 = pi6767 & pi9040;
  assign n67895 = ~n67893 & ~n67894;
  assign n67896 = ~pi1991 & ~n67895;
  assign n67897 = pi1991 & n67895;
  assign n67898 = ~n67896 & ~n67897;
  assign n67899 = ~n67892 & n67898;
  assign n67900 = ~n67886 & n67899;
  assign n67901 = pi6742 & pi9040;
  assign n67902 = pi6775 & ~pi9040;
  assign n67903 = ~n67901 & ~n67902;
  assign n67904 = pi2008 & n67903;
  assign n67905 = ~pi2008 & ~n67903;
  assign n67906 = ~n67904 & ~n67905;
  assign n67907 = n67900 & ~n67906;
  assign n67908 = ~n67886 & ~n67906;
  assign n67909 = ~n67898 & n67908;
  assign n67910 = n67892 & n67909;
  assign n67911 = ~n67907 & ~n67910;
  assign n67912 = n67892 & ~n67898;
  assign n67913 = n67886 & n67906;
  assign n67914 = n67912 & n67913;
  assign n67915 = ~n67892 & ~n67898;
  assign n67916 = ~n67886 & n67915;
  assign n67917 = n67906 & n67916;
  assign n67918 = ~n67914 & ~n67917;
  assign n67919 = n67911 & n67918;
  assign n67920 = n67880 & ~n67919;
  assign n67921 = n67892 & n67898;
  assign n67922 = ~n67886 & n67921;
  assign n67923 = n67906 & n67922;
  assign n67924 = ~n67916 & ~n67923;
  assign n67925 = n67880 & ~n67924;
  assign n67926 = n67886 & n67921;
  assign n67927 = ~n67906 & n67926;
  assign n67928 = ~n67880 & n67898;
  assign n67929 = ~n67906 & n67928;
  assign n67930 = n67886 & ~n67892;
  assign n67931 = n67906 & n67912;
  assign n67932 = ~n67930 & ~n67931;
  assign n67933 = ~n67880 & ~n67932;
  assign n67934 = ~n67929 & ~n67933;
  assign n67935 = ~n67927 & n67934;
  assign n67936 = n67898 & n67930;
  assign n67937 = n67906 & n67936;
  assign n67938 = n67935 & ~n67937;
  assign n67939 = ~n67925 & n67938;
  assign n67940 = pi6759 & pi9040;
  assign n67941 = pi6742 & ~pi9040;
  assign n67942 = ~n67940 & ~n67941;
  assign n67943 = ~pi2013 & ~n67942;
  assign n67944 = pi2013 & n67942;
  assign n67945 = ~n67943 & ~n67944;
  assign n67946 = ~n67939 & ~n67945;
  assign n67947 = ~n67886 & n67898;
  assign n67948 = ~n67880 & n67906;
  assign n67949 = n67945 & n67948;
  assign n67950 = n67947 & n67949;
  assign n67951 = ~n67880 & ~n67909;
  assign n67952 = n67892 & n67913;
  assign n67953 = ~n67899 & ~n67947;
  assign n67954 = ~n67906 & ~n67953;
  assign n67955 = n67886 & n67912;
  assign n67956 = n67880 & ~n67955;
  assign n67957 = ~n67954 & n67956;
  assign n67958 = ~n67952 & n67957;
  assign n67959 = ~n67951 & ~n67958;
  assign n67960 = n67886 & ~n67898;
  assign n67961 = n67906 & n67960;
  assign n67962 = ~n67892 & n67961;
  assign n67963 = ~n67959 & ~n67962;
  assign n67964 = n67945 & ~n67963;
  assign n67965 = ~n67950 & ~n67964;
  assign n67966 = ~n67946 & n67965;
  assign n67967 = ~n67920 & n67966;
  assign n67968 = ~n67880 & n67927;
  assign n67969 = n67967 & ~n67968;
  assign n67970 = pi2019 & ~n67969;
  assign n67971 = ~pi2019 & ~n67968;
  assign n67972 = n67966 & n67971;
  assign n67973 = ~n67920 & n67972;
  assign po2086 = n67970 | n67973;
  assign n67975 = pi6821 & ~pi9040;
  assign n67976 = pi6778 & pi9040;
  assign n67977 = ~n67975 & ~n67976;
  assign n67978 = ~pi1991 & ~n67977;
  assign n67979 = pi1991 & n67977;
  assign n67980 = ~n67978 & ~n67979;
  assign n67981 = pi6762 & ~pi9040;
  assign n67982 = pi6773 & pi9040;
  assign n67983 = ~n67981 & ~n67982;
  assign n67984 = ~pi2006 & n67983;
  assign n67985 = pi2006 & ~n67983;
  assign n67986 = ~n67984 & ~n67985;
  assign n67987 = pi6767 & ~pi9040;
  assign n67988 = pi6725 & pi9040;
  assign n67989 = ~n67987 & ~n67988;
  assign n67990 = pi1972 & n67989;
  assign n67991 = ~pi1972 & ~n67989;
  assign n67992 = ~n67990 & ~n67991;
  assign n67993 = n67986 & n67992;
  assign n67994 = pi6758 & ~pi9040;
  assign n67995 = pi6761 & pi9040;
  assign n67996 = ~n67994 & ~n67995;
  assign n67997 = pi1975 & n67996;
  assign n67998 = ~pi1975 & ~n67996;
  assign n67999 = ~n67997 & ~n67998;
  assign n68000 = pi6757 & ~pi9040;
  assign n68001 = pi6827 & pi9040;
  assign n68002 = ~n68000 & ~n68001;
  assign n68003 = pi2009 & n68002;
  assign n68004 = ~pi2009 & ~n68002;
  assign n68005 = ~n68003 & ~n68004;
  assign n68006 = ~n67999 & ~n68005;
  assign n68007 = n67993 & n68006;
  assign n68008 = pi6724 & ~pi9040;
  assign n68009 = pi6757 & pi9040;
  assign n68010 = ~n68008 & ~n68009;
  assign n68011 = ~pi1999 & n68010;
  assign n68012 = pi1999 & ~n68010;
  assign n68013 = ~n68011 & ~n68012;
  assign n68014 = ~n67986 & ~n67992;
  assign n68015 = ~n68013 & n68014;
  assign n68016 = n67999 & n68013;
  assign n68017 = ~n67992 & n68016;
  assign n68018 = n67986 & n68017;
  assign n68019 = ~n68015 & ~n68018;
  assign n68020 = ~n67986 & n67992;
  assign n68021 = n67999 & n68020;
  assign n68022 = n68019 & ~n68021;
  assign n68023 = ~n68005 & ~n68022;
  assign n68024 = ~n67986 & n68013;
  assign n68025 = ~n67999 & n68005;
  assign n68026 = n68024 & n68025;
  assign n68027 = n68013 & n68014;
  assign n68028 = ~n67999 & n68027;
  assign n68029 = ~n68026 & ~n68028;
  assign n68030 = ~n68023 & n68029;
  assign n68031 = ~n68007 & n68030;
  assign n68032 = n67993 & ~n68013;
  assign n68033 = ~n67999 & n68032;
  assign n68034 = ~n68013 & n68020;
  assign n68035 = n67999 & n68034;
  assign n68036 = ~n68033 & ~n68035;
  assign n68037 = n68031 & n68036;
  assign n68038 = ~n67980 & ~n68037;
  assign n68039 = ~n67999 & n68013;
  assign n68040 = n67992 & n68039;
  assign n68041 = ~n67986 & n68040;
  assign n68042 = ~n68032 & ~n68041;
  assign n68043 = ~n68005 & ~n68042;
  assign n68044 = n67993 & n68016;
  assign n68045 = ~n67992 & n68039;
  assign n68046 = n67986 & n68045;
  assign n68047 = ~n68044 & ~n68046;
  assign n68048 = ~n67986 & n68016;
  assign n68049 = ~n67999 & n68034;
  assign n68050 = ~n68048 & ~n68049;
  assign n68051 = n68005 & ~n68050;
  assign n68052 = n68047 & ~n68051;
  assign n68053 = ~n68043 & n68052;
  assign n68054 = n67980 & ~n68053;
  assign n68055 = ~n67986 & ~n68013;
  assign n68056 = n67999 & n68055;
  assign n68057 = n67986 & ~n68013;
  assign n68058 = ~n67999 & n68057;
  assign n68059 = ~n68056 & ~n68058;
  assign n68060 = ~n68005 & ~n68059;
  assign n68061 = n67986 & ~n67992;
  assign n68062 = ~n68013 & n68061;
  assign n68063 = n67999 & n68062;
  assign n68064 = ~n68044 & ~n68063;
  assign n68065 = ~n68027 & n68064;
  assign n68066 = n68005 & ~n68065;
  assign n68067 = ~n68060 & ~n68066;
  assign n68068 = ~n67992 & n68013;
  assign n68069 = n68005 & n68068;
  assign n68070 = ~n67999 & n68069;
  assign n68071 = n68067 & ~n68070;
  assign n68072 = ~n68054 & n68071;
  assign n68073 = ~n68038 & n68072;
  assign n68074 = ~pi2028 & ~n68073;
  assign n68075 = pi2028 & n68073;
  assign po2092 = n68074 | n68075;
  assign n68077 = pi6854 & pi9040;
  assign n68078 = pi6776 & ~pi9040;
  assign n68079 = ~n68077 & ~n68078;
  assign n68080 = ~pi2006 & ~n68079;
  assign n68081 = pi2006 & n68079;
  assign n68082 = ~n68080 & ~n68081;
  assign n68083 = pi6753 & ~pi9040;
  assign n68084 = pi6719 & pi9040;
  assign n68085 = ~n68083 & ~n68084;
  assign n68086 = ~pi2002 & ~n68085;
  assign n68087 = pi2002 & n68085;
  assign n68088 = ~n68086 & ~n68087;
  assign n68089 = pi6754 & pi9040;
  assign n68090 = pi6773 & ~pi9040;
  assign n68091 = ~n68089 & ~n68090;
  assign n68092 = pi1982 & n68091;
  assign n68093 = ~pi1982 & ~n68091;
  assign n68094 = ~n68092 & ~n68093;
  assign n68095 = pi6754 & ~pi9040;
  assign n68096 = pi6855 & pi9040;
  assign n68097 = ~n68095 & ~n68096;
  assign n68098 = ~pi1983 & n68097;
  assign n68099 = pi1983 & ~n68097;
  assign n68100 = ~n68098 & ~n68099;
  assign n68101 = pi6733 & pi9040;
  assign n68102 = pi6854 & ~pi9040;
  assign n68103 = ~n68101 & ~n68102;
  assign n68104 = ~pi2010 & n68103;
  assign n68105 = pi2010 & ~n68103;
  assign n68106 = ~n68104 & ~n68105;
  assign n68107 = n68100 & ~n68106;
  assign n68108 = n68094 & n68107;
  assign n68109 = pi6764 & pi9040;
  assign n68110 = pi6744 & ~pi9040;
  assign n68111 = ~n68109 & ~n68110;
  assign n68112 = ~pi1999 & n68111;
  assign n68113 = pi1999 & ~n68111;
  assign n68114 = ~n68112 & ~n68113;
  assign n68115 = ~n68100 & ~n68114;
  assign n68116 = ~n68106 & n68115;
  assign n68117 = ~n68108 & ~n68116;
  assign n68118 = ~n68100 & n68114;
  assign n68119 = ~n68094 & n68106;
  assign n68120 = n68118 & n68119;
  assign n68121 = n68117 & ~n68120;
  assign n68122 = n68088 & ~n68121;
  assign n68123 = ~n68100 & n68106;
  assign n68124 = ~n68094 & n68123;
  assign n68125 = ~n68114 & n68124;
  assign n68126 = n68100 & ~n68114;
  assign n68127 = ~n68106 & n68126;
  assign n68128 = ~n68094 & n68127;
  assign n68129 = n68100 & n68106;
  assign n68130 = ~n68118 & ~n68129;
  assign n68131 = n68094 & ~n68130;
  assign n68132 = ~n68128 & ~n68131;
  assign n68133 = ~n68125 & n68132;
  assign n68134 = ~n68088 & ~n68133;
  assign n68135 = ~n68122 & ~n68134;
  assign n68136 = n68082 & ~n68135;
  assign n68137 = n68088 & ~n68094;
  assign n68138 = n68100 & n68137;
  assign n68139 = ~n68088 & ~n68094;
  assign n68140 = n68118 & n68139;
  assign n68141 = ~n68094 & ~n68100;
  assign n68142 = ~n68106 & n68141;
  assign n68143 = ~n68108 & ~n68142;
  assign n68144 = ~n68088 & ~n68143;
  assign n68145 = ~n68140 & ~n68144;
  assign n68146 = ~n68106 & n68118;
  assign n68147 = ~n68094 & n68146;
  assign n68148 = ~n68114 & n68123;
  assign n68149 = n68094 & n68148;
  assign n68150 = ~n68147 & ~n68149;
  assign n68151 = n68088 & n68094;
  assign n68152 = n68123 & n68151;
  assign n68153 = n68106 & n68126;
  assign n68154 = n68088 & n68153;
  assign n68155 = ~n68152 & ~n68154;
  assign n68156 = n68150 & n68155;
  assign n68157 = n68145 & n68156;
  assign n68158 = ~n68138 & n68157;
  assign n68159 = ~n68082 & ~n68158;
  assign n68160 = n68100 & n68114;
  assign n68161 = n68106 & n68160;
  assign n68162 = ~n68088 & n68161;
  assign n68163 = ~n68094 & n68162;
  assign n68164 = ~n68088 & n68147;
  assign n68165 = ~n68163 & ~n68164;
  assign n68166 = ~n68114 & n68119;
  assign n68167 = n68100 & n68166;
  assign n68168 = n68088 & n68167;
  assign n68169 = n68165 & ~n68168;
  assign n68170 = ~n68094 & ~n68106;
  assign n68171 = n68114 & n68170;
  assign n68172 = n68100 & n68171;
  assign n68173 = n68094 & n68115;
  assign n68174 = ~n68172 & ~n68173;
  assign n68175 = n68088 & ~n68174;
  assign n68176 = n68169 & ~n68175;
  assign n68177 = ~n68159 & n68176;
  assign n68178 = ~n68136 & n68177;
  assign n68179 = ~pi2039 & ~n68178;
  assign n68180 = pi2039 & n68178;
  assign po2105 = n68179 | n68180;
  assign n68182 = ~n68082 & ~n68088;
  assign n68183 = ~n68094 & n68107;
  assign n68184 = n68094 & n68146;
  assign n68185 = ~n68094 & n68115;
  assign n68186 = ~n68184 & ~n68185;
  assign n68187 = ~n68183 & n68186;
  assign n68188 = n68182 & ~n68187;
  assign n68189 = n68114 & n68119;
  assign n68190 = ~n68106 & n68160;
  assign n68191 = n68094 & n68190;
  assign n68192 = ~n68189 & ~n68191;
  assign n68193 = n68106 & n68118;
  assign n68194 = ~n68116 & ~n68193;
  assign n68195 = n68192 & n68194;
  assign n68196 = n68088 & ~n68195;
  assign n68197 = n68094 & n68153;
  assign n68198 = ~n68196 & ~n68197;
  assign n68199 = ~n68082 & ~n68198;
  assign n68200 = ~n68188 & ~n68199;
  assign n68201 = ~n68106 & n68137;
  assign n68202 = ~n68114 & n68201;
  assign n68203 = ~n68120 & ~n68202;
  assign n68204 = ~n68115 & ~n68160;
  assign n68205 = n68094 & ~n68204;
  assign n68206 = ~n68161 & ~n68205;
  assign n68207 = ~n68088 & ~n68206;
  assign n68208 = ~n68127 & ~n68183;
  assign n68209 = ~n68184 & n68208;
  assign n68210 = n68088 & ~n68209;
  assign n68211 = ~n68207 & ~n68210;
  assign n68212 = n68094 & n68161;
  assign n68213 = ~n68149 & ~n68212;
  assign n68214 = ~n68167 & n68213;
  assign n68215 = ~n68140 & n68214;
  assign n68216 = n68211 & n68215;
  assign n68217 = n68082 & ~n68216;
  assign n68218 = n68203 & ~n68217;
  assign n68219 = n68200 & n68218;
  assign n68220 = pi2023 & ~n68219;
  assign n68221 = ~pi2023 & n68203;
  assign n68222 = n68200 & n68221;
  assign n68223 = ~n68217 & n68222;
  assign po2106 = n68220 | n68223;
  assign n68225 = n67999 & n68027;
  assign n68226 = ~n68046 & ~n68055;
  assign n68227 = n68005 & ~n68226;
  assign n68228 = ~n68225 & ~n68227;
  assign n68229 = ~n68041 & n68228;
  assign n68230 = ~n68005 & n68044;
  assign n68231 = ~n68033 & ~n68230;
  assign n68232 = ~n68063 & n68231;
  assign n68233 = n68229 & n68232;
  assign n68234 = n67980 & ~n68233;
  assign n68235 = n68013 & n68020;
  assign n68236 = n67999 & n68235;
  assign n68237 = ~n68018 & ~n68236;
  assign n68238 = ~n67999 & n68062;
  assign n68239 = ~n68028 & ~n68238;
  assign n68240 = n67993 & n68013;
  assign n68241 = n68005 & n68240;
  assign n68242 = n67999 & n68032;
  assign n68243 = ~n68241 & ~n68242;
  assign n68244 = n67992 & ~n68013;
  assign n68245 = ~n67986 & n67999;
  assign n68246 = ~n68244 & ~n68245;
  assign n68247 = ~n68068 & n68246;
  assign n68248 = ~n68005 & ~n68247;
  assign n68249 = n68243 & ~n68248;
  assign n68250 = n68239 & n68249;
  assign n68251 = n68237 & n68250;
  assign n68252 = ~n67980 & ~n68251;
  assign n68253 = ~n68234 & ~n68252;
  assign n68254 = pi2040 & ~n68253;
  assign n68255 = ~pi2040 & ~n68234;
  assign n68256 = ~n68252 & n68255;
  assign po2108 = n68254 | n68256;
  assign n68258 = pi6855 & ~pi9040;
  assign n68259 = pi6762 & pi9040;
  assign n68260 = ~n68258 & ~n68259;
  assign n68261 = ~pi1981 & n68260;
  assign n68262 = pi1981 & ~n68260;
  assign n68263 = ~n68261 & ~n68262;
  assign n68264 = pi6858 & ~pi9040;
  assign n68265 = pi6941 & pi9040;
  assign n68266 = ~n68264 & ~n68265;
  assign n68267 = pi2014 & n68266;
  assign n68268 = ~pi2014 & ~n68266;
  assign n68269 = ~n68267 & ~n68268;
  assign n68270 = pi6858 & pi9040;
  assign n68271 = pi6719 & ~pi9040;
  assign n68272 = ~n68270 & ~n68271;
  assign n68273 = pi1992 & n68272;
  assign n68274 = ~pi1992 & ~n68272;
  assign n68275 = ~n68273 & ~n68274;
  assign n68276 = pi6778 & ~pi9040;
  assign n68277 = pi6744 & pi9040;
  assign n68278 = ~n68276 & ~n68277;
  assign n68279 = ~pi2012 & n68278;
  assign n68280 = pi2012 & ~n68278;
  assign n68281 = ~n68279 & ~n68280;
  assign n68282 = pi6764 & ~pi9040;
  assign n68283 = pi6821 & pi9040;
  assign n68284 = ~n68282 & ~n68283;
  assign n68285 = ~pi2010 & ~n68284;
  assign n68286 = pi2010 & n68284;
  assign n68287 = ~n68285 & ~n68286;
  assign n68288 = n68281 & n68287;
  assign n68289 = ~n68275 & n68288;
  assign n68290 = ~n68269 & n68289;
  assign n68291 = n68275 & ~n68287;
  assign n68292 = ~n68281 & n68291;
  assign n68293 = n68269 & n68292;
  assign n68294 = n68269 & ~n68275;
  assign n68295 = ~n68287 & n68294;
  assign n68296 = n68281 & n68295;
  assign n68297 = ~n68293 & ~n68296;
  assign n68298 = ~n68290 & n68297;
  assign n68299 = ~n68263 & ~n68298;
  assign n68300 = ~n68269 & n68275;
  assign n68301 = n68287 & n68300;
  assign n68302 = ~n68281 & n68301;
  assign n68303 = pi6770 & pi9040;
  assign n68304 = pi6733 & ~pi9040;
  assign n68305 = ~n68303 & ~n68304;
  assign n68306 = pi1983 & n68305;
  assign n68307 = ~pi1983 & ~n68305;
  assign n68308 = ~n68306 & ~n68307;
  assign n68309 = n68281 & n68300;
  assign n68310 = ~n68281 & n68287;
  assign n68311 = ~n68275 & n68310;
  assign n68312 = ~n68309 & ~n68311;
  assign n68313 = n68263 & ~n68312;
  assign n68314 = ~n68301 & ~n68313;
  assign n68315 = n68275 & n68310;
  assign n68316 = ~n68275 & n68281;
  assign n68317 = ~n68275 & ~n68287;
  assign n68318 = ~n68269 & n68317;
  assign n68319 = n68281 & ~n68287;
  assign n68320 = n68269 & n68319;
  assign n68321 = ~n68318 & ~n68320;
  assign n68322 = ~n68316 & n68321;
  assign n68323 = ~n68315 & n68322;
  assign n68324 = ~n68263 & ~n68323;
  assign n68325 = n68314 & ~n68324;
  assign n68326 = ~n68293 & n68325;
  assign n68327 = n68308 & ~n68326;
  assign n68328 = ~n68302 & ~n68327;
  assign n68329 = ~n68299 & n68328;
  assign n68330 = ~n68275 & ~n68281;
  assign n68331 = n68263 & n68330;
  assign n68332 = n68269 & n68331;
  assign n68333 = n68275 & n68288;
  assign n68334 = n68269 & n68333;
  assign n68335 = ~n68263 & n68291;
  assign n68336 = ~n68269 & n68335;
  assign n68337 = ~n68334 & ~n68336;
  assign n68338 = n68275 & n68281;
  assign n68339 = n68269 & n68338;
  assign n68340 = ~n68281 & ~n68287;
  assign n68341 = ~n68275 & n68340;
  assign n68342 = ~n68339 & ~n68341;
  assign n68343 = n68263 & ~n68342;
  assign n68344 = n68263 & n68316;
  assign n68345 = ~n68269 & n68344;
  assign n68346 = ~n68343 & ~n68345;
  assign n68347 = n68337 & n68346;
  assign n68348 = ~n68308 & ~n68347;
  assign n68349 = ~n68332 & ~n68348;
  assign n68350 = n68329 & n68349;
  assign n68351 = pi2018 & n68350;
  assign n68352 = ~n68302 & ~n68332;
  assign n68353 = ~n68348 & n68352;
  assign n68354 = ~n68299 & ~n68327;
  assign n68355 = n68353 & n68354;
  assign n68356 = ~pi2018 & ~n68355;
  assign po2109 = n68351 | n68356;
  assign n68358 = pi6716 & ~pi9040;
  assign n68359 = pi6746 & pi9040;
  assign n68360 = ~n68358 & ~n68359;
  assign n68361 = ~pi2012 & ~n68360;
  assign n68362 = pi2012 & n68360;
  assign n68363 = ~n68361 & ~n68362;
  assign n68364 = pi6857 & ~pi9040;
  assign n68365 = pi6782 & pi9040;
  assign n68366 = ~n68364 & ~n68365;
  assign n68367 = ~pi2001 & n68366;
  assign n68368 = pi2001 & ~n68366;
  assign n68369 = ~n68367 & ~n68368;
  assign n68370 = pi6760 & ~pi9040;
  assign n68371 = pi6752 & pi9040;
  assign n68372 = ~n68370 & ~n68371;
  assign n68373 = pi2011 & n68372;
  assign n68374 = ~pi2011 & ~n68372;
  assign n68375 = ~n68373 & ~n68374;
  assign n68376 = pi6780 & ~pi9040;
  assign n68377 = pi6859 & pi9040;
  assign n68378 = ~n68376 & ~n68377;
  assign n68379 = ~pi1990 & ~n68378;
  assign n68380 = pi1990 & n68378;
  assign n68381 = ~n68379 & ~n68380;
  assign n68382 = pi6715 & pi9040;
  assign n68383 = pi6747 & ~pi9040;
  assign n68384 = ~n68382 & ~n68383;
  assign n68385 = ~pi1992 & n68384;
  assign n68386 = pi1992 & ~n68384;
  assign n68387 = ~n68385 & ~n68386;
  assign n68388 = ~n68381 & ~n68387;
  assign n68389 = n68375 & n68388;
  assign n68390 = ~n68369 & n68389;
  assign n68391 = pi6857 & pi9040;
  assign n68392 = pi6746 & ~pi9040;
  assign n68393 = ~n68391 & ~n68392;
  assign n68394 = pi2015 & n68393;
  assign n68395 = ~pi2015 & ~n68393;
  assign n68396 = ~n68394 & ~n68395;
  assign n68397 = n68381 & ~n68387;
  assign n68398 = ~n68369 & n68397;
  assign n68399 = ~n68375 & n68388;
  assign n68400 = n68369 & n68399;
  assign n68401 = ~n68398 & ~n68400;
  assign n68402 = ~n68396 & ~n68401;
  assign n68403 = ~n68390 & ~n68402;
  assign n68404 = ~n68381 & n68387;
  assign n68405 = ~n68375 & n68404;
  assign n68406 = n68396 & n68405;
  assign n68407 = n68388 & n68396;
  assign n68408 = ~n68369 & n68407;
  assign n68409 = ~n68406 & ~n68408;
  assign n68410 = n68403 & n68409;
  assign n68411 = n68381 & n68387;
  assign n68412 = n68375 & n68411;
  assign n68413 = ~n68369 & n68412;
  assign n68414 = n68375 & n68404;
  assign n68415 = n68369 & n68414;
  assign n68416 = ~n68413 & ~n68415;
  assign n68417 = n68410 & n68416;
  assign n68418 = n68363 & ~n68417;
  assign n68419 = ~n68363 & ~n68396;
  assign n68420 = ~n68369 & ~n68375;
  assign n68421 = ~n68381 & n68420;
  assign n68422 = ~n68375 & n68387;
  assign n68423 = ~n68421 & ~n68422;
  assign n68424 = n68419 & ~n68423;
  assign n68425 = n68369 & n68375;
  assign n68426 = ~n68387 & n68425;
  assign n68427 = ~n68381 & n68426;
  assign n68428 = n68369 & n68381;
  assign n68429 = ~n68375 & n68428;
  assign n68430 = ~n68427 & ~n68429;
  assign n68431 = ~n68369 & n68396;
  assign n68432 = n68375 & n68431;
  assign n68433 = ~n68388 & n68432;
  assign n68434 = n68396 & n68412;
  assign n68435 = ~n68433 & ~n68434;
  assign n68436 = n68430 & n68435;
  assign n68437 = ~n68363 & ~n68436;
  assign n68438 = ~n68375 & n68411;
  assign n68439 = ~n68396 & n68438;
  assign n68440 = n68369 & n68439;
  assign n68441 = n68375 & n68397;
  assign n68442 = n68369 & n68441;
  assign n68443 = ~n68415 & ~n68442;
  assign n68444 = ~n68396 & ~n68443;
  assign n68445 = ~n68440 & ~n68444;
  assign n68446 = n68396 & n68427;
  assign n68447 = n68445 & ~n68446;
  assign n68448 = ~n68437 & n68447;
  assign n68449 = ~n68424 & n68448;
  assign n68450 = ~n68418 & n68449;
  assign n68451 = ~n68375 & n68397;
  assign n68452 = n68369 & n68396;
  assign n68453 = n68451 & n68452;
  assign n68454 = n68450 & ~n68453;
  assign n68455 = ~pi2021 & ~n68454;
  assign n68456 = ~n68418 & ~n68453;
  assign n68457 = n68449 & n68456;
  assign n68458 = pi2021 & n68457;
  assign po2110 = n68455 | n68458;
  assign n68460 = pi6771 & pi9040;
  assign n68461 = pi6852 & ~pi9040;
  assign n68462 = ~n68460 & ~n68461;
  assign n68463 = ~pi1989 & ~n68462;
  assign n68464 = pi1989 & n68462;
  assign n68465 = ~n68463 & ~n68464;
  assign n68466 = pi6743 & ~pi9040;
  assign n68467 = pi6741 & pi9040;
  assign n68468 = ~n68466 & ~n68467;
  assign n68469 = ~pi2003 & ~n68468;
  assign n68470 = pi2003 & n68468;
  assign n68471 = ~n68469 & ~n68470;
  assign n68472 = pi6752 & ~pi9040;
  assign n68473 = pi6749 & pi9040;
  assign n68474 = ~n68472 & ~n68473;
  assign n68475 = ~pi2013 & ~n68474;
  assign n68476 = pi2013 & n68474;
  assign n68477 = ~n68475 & ~n68476;
  assign n68478 = pi6751 & pi9040;
  assign n68479 = pi6756 & ~pi9040;
  assign n68480 = ~n68478 & ~n68479;
  assign n68481 = ~pi1974 & n68480;
  assign n68482 = pi1974 & ~n68480;
  assign n68483 = ~n68481 & ~n68482;
  assign n68484 = ~n68477 & ~n68483;
  assign n68485 = pi6772 & ~pi9040;
  assign n68486 = pi6717 & pi9040;
  assign n68487 = ~n68485 & ~n68486;
  assign n68488 = ~pi1998 & n68487;
  assign n68489 = pi1998 & ~n68487;
  assign n68490 = ~n68488 & ~n68489;
  assign n68491 = pi6741 & ~pi9040;
  assign n68492 = pi6750 & pi9040;
  assign n68493 = ~n68491 & ~n68492;
  assign n68494 = pi2007 & n68493;
  assign n68495 = ~pi2007 & ~n68493;
  assign n68496 = ~n68494 & ~n68495;
  assign n68497 = ~n68490 & n68496;
  assign n68498 = n68484 & n68497;
  assign n68499 = n68471 & n68498;
  assign n68500 = n68490 & n68496;
  assign n68501 = n68477 & ~n68483;
  assign n68502 = n68500 & n68501;
  assign n68503 = n68477 & n68483;
  assign n68504 = n68471 & n68503;
  assign n68505 = n68496 & n68504;
  assign n68506 = ~n68490 & n68505;
  assign n68507 = n68471 & n68490;
  assign n68508 = n68483 & n68507;
  assign n68509 = ~n68477 & n68508;
  assign n68510 = ~n68506 & ~n68509;
  assign n68511 = ~n68502 & n68510;
  assign n68512 = ~n68499 & n68511;
  assign n68513 = ~n68471 & n68490;
  assign n68514 = ~n68483 & n68513;
  assign n68515 = n68477 & n68514;
  assign n68516 = n68512 & ~n68515;
  assign n68517 = ~n68465 & ~n68516;
  assign n68518 = n68471 & n68477;
  assign n68519 = ~n68483 & n68518;
  assign n68520 = ~n68490 & n68519;
  assign n68521 = ~n68508 & ~n68520;
  assign n68522 = ~n68471 & n68484;
  assign n68523 = ~n68490 & n68522;
  assign n68524 = n68521 & ~n68523;
  assign n68525 = ~n68496 & ~n68524;
  assign n68526 = ~n68471 & n68483;
  assign n68527 = n68477 & n68526;
  assign n68528 = ~n68496 & n68527;
  assign n68529 = ~n68490 & n68528;
  assign n68530 = ~n68477 & n68507;
  assign n68531 = ~n68477 & n68483;
  assign n68532 = n68490 & n68531;
  assign n68533 = ~n68530 & ~n68532;
  assign n68534 = ~n68496 & ~n68533;
  assign n68535 = ~n68529 & ~n68534;
  assign n68536 = ~n68465 & ~n68535;
  assign n68537 = ~n68525 & ~n68536;
  assign n68538 = ~n68517 & n68537;
  assign n68539 = ~n68471 & ~n68490;
  assign n68540 = n68496 & n68539;
  assign n68541 = n68531 & n68540;
  assign n68542 = ~n68471 & n68477;
  assign n68543 = n68500 & n68542;
  assign n68544 = n68490 & n68527;
  assign n68545 = n68471 & ~n68496;
  assign n68546 = n68477 & n68545;
  assign n68547 = ~n68477 & ~n68490;
  assign n68548 = ~n68471 & n68547;
  assign n68549 = ~n68546 & ~n68548;
  assign n68550 = ~n68544 & n68549;
  assign n68551 = ~n68522 & n68550;
  assign n68552 = n68484 & n68496;
  assign n68553 = n68490 & n68552;
  assign n68554 = ~n68490 & n68531;
  assign n68555 = ~n68471 & ~n68483;
  assign n68556 = ~n68554 & ~n68555;
  assign n68557 = n68496 & ~n68556;
  assign n68558 = ~n68553 & ~n68557;
  assign n68559 = n68551 & n68558;
  assign n68560 = n68465 & ~n68559;
  assign n68561 = ~n68543 & ~n68560;
  assign n68562 = ~n68541 & n68561;
  assign n68563 = n68538 & n68562;
  assign n68564 = pi2038 & n68563;
  assign n68565 = ~pi2038 & ~n68563;
  assign po2111 = n68564 | n68565;
  assign n68567 = n68369 & n68405;
  assign n68568 = n68387 & n68420;
  assign n68569 = n68381 & n68568;
  assign n68570 = ~n68567 & ~n68569;
  assign n68571 = n68396 & ~n68570;
  assign n68572 = ~n68427 & ~n68434;
  assign n68573 = ~n68381 & n68425;
  assign n68574 = ~n68429 & ~n68573;
  assign n68575 = ~n68396 & ~n68574;
  assign n68576 = ~n68369 & ~n68396;
  assign n68577 = n68404 & n68576;
  assign n68578 = ~n68375 & n68577;
  assign n68579 = ~n68369 & n68375;
  assign n68580 = ~n68387 & n68579;
  assign n68581 = n68381 & n68580;
  assign n68582 = n68396 & n68399;
  assign n68583 = ~n68581 & ~n68582;
  assign n68584 = ~n68578 & n68583;
  assign n68585 = ~n68575 & n68584;
  assign n68586 = n68572 & n68585;
  assign n68587 = n68363 & ~n68586;
  assign n68588 = ~n68396 & n68427;
  assign n68589 = n68369 & n68434;
  assign n68590 = ~n68588 & ~n68589;
  assign n68591 = ~n68587 & n68590;
  assign n68592 = ~n68571 & n68591;
  assign n68593 = n68375 & ~n68381;
  assign n68594 = n68431 & n68593;
  assign n68595 = ~n68406 & ~n68594;
  assign n68596 = n68396 & n68441;
  assign n68597 = n68369 & n68451;
  assign n68598 = ~n68596 & ~n68597;
  assign n68599 = ~n68369 & n68414;
  assign n68600 = ~n68567 & ~n68599;
  assign n68601 = ~n68369 & n68411;
  assign n68602 = ~n68375 & ~n68387;
  assign n68603 = ~n68601 & ~n68602;
  assign n68604 = ~n68396 & ~n68603;
  assign n68605 = n68600 & ~n68604;
  assign n68606 = n68598 & n68605;
  assign n68607 = n68595 & n68606;
  assign n68608 = ~n68363 & ~n68607;
  assign n68609 = n68592 & ~n68608;
  assign n68610 = ~pi2017 & ~n68609;
  assign n68611 = pi2017 & n68609;
  assign po2112 = n68610 | n68611;
  assign n68613 = n68088 & n68115;
  assign n68614 = ~n68094 & n68613;
  assign n68615 = ~n68172 & ~n68614;
  assign n68616 = n68094 & ~n68114;
  assign n68617 = ~n68106 & n68616;
  assign n68618 = ~n68094 & n68100;
  assign n68619 = ~n68171 & ~n68618;
  assign n68620 = ~n68088 & ~n68619;
  assign n68621 = ~n68617 & ~n68620;
  assign n68622 = n68615 & n68621;
  assign n68623 = n68082 & ~n68622;
  assign n68624 = ~n68146 & ~n68149;
  assign n68625 = ~n68094 & n68126;
  assign n68626 = n68624 & ~n68625;
  assign n68627 = n68088 & ~n68626;
  assign n68628 = n68115 & n68139;
  assign n68629 = ~n68120 & ~n68628;
  assign n68630 = ~n68627 & n68629;
  assign n68631 = ~n68190 & ~n68197;
  assign n68632 = ~n68088 & ~n68631;
  assign n68633 = n68630 & ~n68632;
  assign n68634 = ~n68082 & ~n68633;
  assign n68635 = ~n68623 & ~n68634;
  assign n68636 = ~n68094 & n68160;
  assign n68637 = n68094 & ~n68194;
  assign n68638 = ~n68636 & ~n68637;
  assign n68639 = ~n68088 & ~n68638;
  assign n68640 = ~n68127 & ~n68161;
  assign n68641 = ~n68146 & n68640;
  assign n68642 = n68151 & ~n68641;
  assign n68643 = ~n68639 & ~n68642;
  assign n68644 = n68635 & n68643;
  assign n68645 = ~pi2027 & ~n68644;
  assign n68646 = ~n68634 & n68643;
  assign n68647 = pi2027 & n68646;
  assign n68648 = ~n68623 & n68647;
  assign po2113 = n68645 | n68648;
  assign n68650 = pi6782 & ~pi9040;
  assign n68651 = pi6716 & pi9040;
  assign n68652 = ~n68650 & ~n68651;
  assign n68653 = pi2005 & n68652;
  assign n68654 = ~pi2005 & ~n68652;
  assign n68655 = ~n68653 & ~n68654;
  assign n68656 = pi6768 & pi9040;
  assign n68657 = pi6750 & ~pi9040;
  assign n68658 = ~n68656 & ~n68657;
  assign n68659 = pi1989 & n68658;
  assign n68660 = ~pi1989 & ~n68658;
  assign n68661 = ~n68659 & ~n68660;
  assign n68662 = pi6768 & ~pi9040;
  assign n68663 = pi6743 & pi9040;
  assign n68664 = ~n68662 & ~n68663;
  assign n68665 = pi1997 & n68664;
  assign n68666 = ~pi1997 & ~n68664;
  assign n68667 = ~n68665 & ~n68666;
  assign n68668 = n68661 & ~n68667;
  assign n68669 = pi6849 & ~pi9040;
  assign n68670 = pi6777 & pi9040;
  assign n68671 = ~n68669 & ~n68670;
  assign n68672 = ~pi2004 & n68671;
  assign n68673 = pi2004 & ~n68671;
  assign n68674 = ~n68672 & ~n68673;
  assign n68675 = pi6728 & ~pi9040;
  assign n68676 = pi6760 & pi9040;
  assign n68677 = ~n68675 & ~n68676;
  assign n68678 = ~pi1974 & n68677;
  assign n68679 = pi1974 & ~n68677;
  assign n68680 = ~n68678 & ~n68679;
  assign n68681 = ~n68674 & ~n68680;
  assign n68682 = n68668 & n68681;
  assign n68683 = ~n68674 & n68680;
  assign n68684 = ~n68661 & n68683;
  assign n68685 = ~n68682 & ~n68684;
  assign n68686 = ~n68655 & ~n68685;
  assign n68687 = pi6728 & pi9040;
  assign n68688 = pi6749 & ~pi9040;
  assign n68689 = ~n68687 & ~n68688;
  assign n68690 = ~pi2000 & ~n68689;
  assign n68691 = pi2000 & n68689;
  assign n68692 = ~n68690 & ~n68691;
  assign n68693 = n68655 & n68674;
  assign n68694 = n68661 & n68693;
  assign n68695 = n68668 & n68680;
  assign n68696 = n68661 & n68667;
  assign n68697 = ~n68680 & n68696;
  assign n68698 = ~n68695 & ~n68697;
  assign n68699 = ~n68661 & ~n68667;
  assign n68700 = ~n68680 & n68699;
  assign n68701 = ~n68674 & n68700;
  assign n68702 = n68698 & ~n68701;
  assign n68703 = n68655 & ~n68702;
  assign n68704 = ~n68694 & ~n68703;
  assign n68705 = ~n68661 & n68667;
  assign n68706 = n68680 & n68705;
  assign n68707 = ~n68674 & n68706;
  assign n68708 = n68704 & ~n68707;
  assign n68709 = n68674 & n68699;
  assign n68710 = ~n68661 & ~n68680;
  assign n68711 = n68667 & n68710;
  assign n68712 = ~n68709 & ~n68711;
  assign n68713 = ~n68655 & ~n68712;
  assign n68714 = n68680 & n68696;
  assign n68715 = n68674 & n68714;
  assign n68716 = ~n68713 & ~n68715;
  assign n68717 = n68708 & n68716;
  assign n68718 = n68692 & ~n68717;
  assign n68719 = ~n68686 & ~n68718;
  assign n68720 = n68655 & ~n68692;
  assign n68721 = ~n68712 & n68720;
  assign n68722 = n68680 & n68699;
  assign n68723 = ~n68714 & ~n68722;
  assign n68724 = ~n68674 & ~n68723;
  assign n68725 = ~n68682 & ~n68724;
  assign n68726 = ~n68692 & ~n68725;
  assign n68727 = ~n68721 & ~n68726;
  assign n68728 = ~n68655 & ~n68692;
  assign n68729 = n68668 & n68674;
  assign n68730 = ~n68706 & ~n68729;
  assign n68731 = n68661 & ~n68680;
  assign n68732 = n68730 & ~n68731;
  assign n68733 = n68728 & ~n68732;
  assign n68734 = n68727 & ~n68733;
  assign n68735 = n68719 & n68734;
  assign n68736 = ~pi2022 & ~n68735;
  assign n68737 = pi2022 & n68727;
  assign n68738 = n68719 & n68737;
  assign n68739 = ~n68733 & n68738;
  assign po2114 = n68736 | n68739;
  assign n68741 = ~n68589 & ~n68594;
  assign n68742 = ~n68387 & n68420;
  assign n68743 = ~n68381 & n68742;
  assign n68744 = ~n68581 & ~n68743;
  assign n68745 = ~n68567 & n68744;
  assign n68746 = ~n68396 & ~n68745;
  assign n68747 = n68369 & n68407;
  assign n68748 = n68381 & n68420;
  assign n68749 = ~n68438 & ~n68748;
  assign n68750 = n68396 & ~n68749;
  assign n68751 = ~n68747 & ~n68750;
  assign n68752 = n68381 & n68425;
  assign n68753 = ~n68567 & ~n68752;
  assign n68754 = ~n68599 & n68753;
  assign n68755 = ~n68396 & n68397;
  assign n68756 = n68369 & n68755;
  assign n68757 = ~n68396 & n68405;
  assign n68758 = ~n68756 & ~n68757;
  assign n68759 = n68754 & n68758;
  assign n68760 = n68751 & n68759;
  assign n68761 = ~n68363 & ~n68760;
  assign n68762 = ~n68427 & ~n68438;
  assign n68763 = ~n68601 & n68762;
  assign n68764 = ~n68396 & ~n68763;
  assign n68765 = ~n68453 & n68744;
  assign n68766 = n68396 & n68414;
  assign n68767 = n68765 & ~n68766;
  assign n68768 = ~n68764 & n68767;
  assign n68769 = n68363 & ~n68768;
  assign n68770 = ~n68761 & ~n68769;
  assign n68771 = ~n68746 & n68770;
  assign n68772 = n68741 & n68771;
  assign n68773 = pi2024 & ~n68772;
  assign n68774 = ~pi2024 & n68772;
  assign po2115 = n68773 | n68774;
  assign n68776 = ~n67906 & n67936;
  assign n68777 = n67906 & n67947;
  assign n68778 = ~n67926 & ~n68777;
  assign n68779 = n67880 & ~n68778;
  assign n68780 = ~n68776 & ~n68779;
  assign n68781 = ~n67880 & n67899;
  assign n68782 = ~n67906 & n68781;
  assign n68783 = n67915 & n67948;
  assign n68784 = ~n68782 & ~n68783;
  assign n68785 = ~n67880 & n67955;
  assign n68786 = n68784 & ~n68785;
  assign n68787 = ~n67910 & ~n67923;
  assign n68788 = ~n67898 & n67913;
  assign n68789 = n68787 & ~n68788;
  assign n68790 = n68786 & n68789;
  assign n68791 = n68780 & n68790;
  assign n68792 = ~n67945 & ~n68791;
  assign n68793 = ~n67886 & n67912;
  assign n68794 = ~n67926 & ~n68793;
  assign n68795 = n67906 & ~n68794;
  assign n68796 = ~n67892 & n67908;
  assign n68797 = n67886 & n67915;
  assign n68798 = ~n68796 & ~n68797;
  assign n68799 = n67886 & n67898;
  assign n68800 = n67906 & n68799;
  assign n68801 = n68798 & ~n68800;
  assign n68802 = n67880 & ~n68801;
  assign n68803 = ~n67906 & n67921;
  assign n68804 = ~n67886 & n67906;
  assign n68805 = n67898 & n68804;
  assign n68806 = ~n67892 & n68805;
  assign n68807 = ~n68803 & ~n68806;
  assign n68808 = ~n67880 & ~n68807;
  assign n68809 = ~n67892 & n67909;
  assign n68810 = ~n68808 & ~n68809;
  assign n68811 = ~n68802 & n68810;
  assign n68812 = ~n68795 & n68811;
  assign n68813 = n67945 & ~n68812;
  assign n68814 = n67880 & n67909;
  assign n68815 = ~n68813 & ~n68814;
  assign n68816 = ~n67880 & n68776;
  assign n68817 = n68815 & ~n68816;
  assign n68818 = ~n68792 & n68817;
  assign n68819 = ~pi2031 & ~n68818;
  assign n68820 = pi2031 & n68815;
  assign n68821 = ~n68792 & n68820;
  assign n68822 = ~n68816 & n68821;
  assign po2118 = n68819 | n68822;
  assign n68824 = ~n67907 & ~n67914;
  assign n68825 = ~n67880 & ~n68824;
  assign n68826 = ~n67968 & ~n68825;
  assign n68827 = ~n67886 & n67892;
  assign n68828 = n67880 & n68827;
  assign n68829 = n67906 & n68828;
  assign n68830 = n67906 & n67921;
  assign n68831 = ~n68827 & ~n68830;
  assign n68832 = n67886 & ~n67906;
  assign n68833 = ~n67892 & n68832;
  assign n68834 = n68831 & ~n68833;
  assign n68835 = n67880 & ~n68834;
  assign n68836 = ~n67917 & ~n68835;
  assign n68837 = ~n67945 & ~n68836;
  assign n68838 = n67906 & n68781;
  assign n68839 = ~n68785 & ~n68838;
  assign n68840 = ~n67945 & ~n68839;
  assign n68841 = ~n68837 & ~n68840;
  assign n68842 = ~n68829 & n68841;
  assign n68843 = ~n67909 & ~n67926;
  assign n68844 = ~n68797 & n68843;
  assign n68845 = ~n67880 & ~n68844;
  assign n68846 = ~n67906 & n67955;
  assign n68847 = ~n67936 & ~n68846;
  assign n68848 = n67880 & ~n68847;
  assign n68849 = ~n68845 & ~n68848;
  assign n68850 = ~n68796 & n68849;
  assign n68851 = ~n67923 & ~n67962;
  assign n68852 = n68850 & n68851;
  assign n68853 = n67945 & ~n68852;
  assign n68854 = n68842 & ~n68853;
  assign n68855 = n68826 & n68854;
  assign n68856 = ~pi2044 & ~n68855;
  assign n68857 = pi2044 & n68842;
  assign n68858 = n68826 & n68857;
  assign n68859 = ~n68853 & n68858;
  assign po2119 = n68856 | n68859;
  assign n68861 = ~n67999 & n68020;
  assign n68862 = ~n68238 & ~n68861;
  assign n68863 = n68005 & n68862;
  assign n68864 = n67999 & n68057;
  assign n68865 = ~n67993 & ~n68014;
  assign n68866 = ~n68013 & ~n68865;
  assign n68867 = n67986 & n68039;
  assign n68868 = n67999 & n68014;
  assign n68869 = ~n68867 & ~n68868;
  assign n68870 = ~n68866 & n68869;
  assign n68871 = ~n68005 & n68870;
  assign n68872 = ~n68864 & n68871;
  assign n68873 = ~n68863 & ~n68872;
  assign n68874 = n67999 & n68866;
  assign n68875 = ~n68236 & ~n68874;
  assign n68876 = ~n68873 & n68875;
  assign n68877 = n67980 & ~n68876;
  assign n68878 = n68005 & ~n68865;
  assign n68879 = ~n67999 & n68878;
  assign n68880 = ~n68034 & ~n68061;
  assign n68881 = n67999 & ~n68880;
  assign n68882 = n68005 & n68881;
  assign n68883 = n68013 & n68878;
  assign n68884 = ~n68882 & ~n68883;
  assign n68885 = ~n68879 & n68884;
  assign n68886 = ~n67980 & ~n68885;
  assign n68887 = ~n68877 & ~n68886;
  assign n68888 = ~n68005 & ~n68862;
  assign n68889 = ~n68018 & ~n68888;
  assign n68890 = ~n67980 & ~n68889;
  assign n68891 = n68005 & n68018;
  assign n68892 = ~n68005 & ~n68875;
  assign n68893 = ~n68891 & ~n68892;
  assign n68894 = ~n68890 & n68893;
  assign n68895 = n68887 & n68894;
  assign n68896 = pi2051 & ~n68895;
  assign n68897 = ~pi2051 & n68894;
  assign n68898 = ~n68886 & n68897;
  assign n68899 = ~n68877 & n68898;
  assign po2120 = n68896 | n68899;
  assign n68901 = n68471 & ~n68477;
  assign n68902 = ~n68515 & ~n68901;
  assign n68903 = ~n68547 & n68902;
  assign n68904 = n68496 & ~n68903;
  assign n68905 = ~n68490 & ~n68496;
  assign n68906 = n68477 & n68905;
  assign n68907 = n68471 & ~n68490;
  assign n68908 = ~n68483 & n68907;
  assign n68909 = n68490 & n68504;
  assign n68910 = ~n68908 & ~n68909;
  assign n68911 = ~n68471 & ~n68477;
  assign n68912 = n68490 & ~n68496;
  assign n68913 = n68911 & n68912;
  assign n68914 = n68910 & ~n68913;
  assign n68915 = ~n68906 & n68914;
  assign n68916 = ~n68904 & n68915;
  assign n68917 = n68465 & ~n68916;
  assign n68918 = n68471 & n68484;
  assign n68919 = n68490 & n68918;
  assign n68920 = n68471 & n68531;
  assign n68921 = ~n68490 & n68920;
  assign n68922 = ~n68919 & ~n68921;
  assign n68923 = n68496 & ~n68922;
  assign n68924 = ~n68917 & ~n68923;
  assign n68925 = ~n68490 & n68504;
  assign n68926 = ~n68519 & ~n68527;
  assign n68927 = n68496 & ~n68926;
  assign n68928 = ~n68925 & ~n68927;
  assign n68929 = ~n68523 & n68928;
  assign n68930 = ~n68465 & ~n68929;
  assign n68931 = ~n68501 & ~n68531;
  assign n68932 = ~n68471 & ~n68931;
  assign n68933 = ~n68532 & ~n68932;
  assign n68934 = ~n68496 & ~n68933;
  assign n68935 = ~n68465 & n68934;
  assign n68936 = ~n68930 & ~n68935;
  assign n68937 = n68924 & n68936;
  assign n68938 = pi2047 & ~n68937;
  assign n68939 = ~pi2047 & n68924;
  assign n68940 = n68936 & n68939;
  assign po2121 = n68938 | n68940;
  assign n68942 = ~n68094 & n68148;
  assign n68943 = ~n68088 & n68942;
  assign n68944 = ~n68164 & ~n68943;
  assign n68945 = ~n68168 & n68944;
  assign n68946 = ~n68167 & ~n68171;
  assign n68947 = n68088 & n68142;
  assign n68948 = n68094 & n68127;
  assign n68949 = ~n68088 & n68123;
  assign n68950 = ~n68948 & ~n68949;
  assign n68951 = ~n68212 & n68950;
  assign n68952 = ~n68947 & n68951;
  assign n68953 = n68946 & n68952;
  assign n68954 = ~n68154 & n68953;
  assign n68955 = n68082 & ~n68954;
  assign n68956 = n68945 & ~n68955;
  assign n68957 = ~n68088 & ~n68640;
  assign n68958 = n68094 & n68116;
  assign n68959 = ~n68957 & ~n68958;
  assign n68960 = n68094 & ~n68100;
  assign n68961 = ~n68123 & ~n68960;
  assign n68962 = ~n68190 & n68961;
  assign n68963 = n68088 & ~n68962;
  assign n68964 = n68959 & ~n68963;
  assign n68965 = ~n68082 & ~n68964;
  assign n68966 = n68956 & ~n68965;
  assign n68967 = ~pi2046 & ~n68966;
  assign n68968 = n68945 & ~n68965;
  assign n68969 = ~n68955 & n68968;
  assign n68970 = pi2046 & n68969;
  assign po2122 = n68967 | n68970;
  assign n68972 = n68263 & ~n68269;
  assign n68973 = ~n68281 & n68972;
  assign n68974 = n68275 & n68319;
  assign n68975 = n68269 & n68974;
  assign n68976 = n68288 & n68294;
  assign n68977 = ~n68975 & ~n68976;
  assign n68978 = ~n68275 & n68319;
  assign n68979 = ~n68269 & n68978;
  assign n68980 = ~n68311 & ~n68979;
  assign n68981 = ~n68263 & ~n68980;
  assign n68982 = n68977 & ~n68981;
  assign n68983 = ~n68973 & n68982;
  assign n68984 = n68308 & ~n68983;
  assign n68985 = n68269 & n68341;
  assign n68986 = n68263 & n68985;
  assign n68987 = ~n68263 & ~n68269;
  assign n68988 = n68341 & n68987;
  assign n68989 = ~n68309 & ~n68988;
  assign n68990 = ~n68311 & ~n68333;
  assign n68991 = ~n68269 & n68288;
  assign n68992 = n68990 & ~n68991;
  assign n68993 = n68263 & ~n68992;
  assign n68994 = ~n68263 & n68315;
  assign n68995 = n68297 & ~n68994;
  assign n68996 = ~n68993 & n68995;
  assign n68997 = n68989 & n68996;
  assign n68998 = ~n68308 & ~n68997;
  assign n68999 = ~n68986 & ~n68998;
  assign n69000 = ~n68984 & n68999;
  assign n69001 = n68333 & n68987;
  assign n69002 = n68269 & n68335;
  assign n69003 = ~n69001 & ~n69002;
  assign n69004 = ~n68263 & n68976;
  assign n69005 = n69003 & ~n69004;
  assign n69006 = n69000 & n69005;
  assign n69007 = ~pi2020 & ~n69006;
  assign n69008 = pi2020 & n69005;
  assign n69009 = n68999 & n69008;
  assign n69010 = ~n68984 & n69009;
  assign po2123 = n69007 | n69010;
  assign n69012 = n67999 & n68240;
  assign n69013 = n68005 & n69012;
  assign n69014 = n68039 & ~n68865;
  assign n69015 = ~n68062 & ~n69014;
  assign n69016 = ~n68236 & n69015;
  assign n69017 = ~n68005 & ~n69016;
  assign n69018 = n67999 & n68015;
  assign n69019 = ~n69017 & ~n69018;
  assign n69020 = n68013 & n68061;
  assign n69021 = ~n67999 & n68244;
  assign n69022 = ~n69020 & ~n69021;
  assign n69023 = ~n68868 & n69022;
  assign n69024 = n68005 & ~n69023;
  assign n69025 = n69019 & ~n69024;
  assign n69026 = n67980 & ~n69025;
  assign n69027 = ~n69013 & ~n69026;
  assign n69028 = ~n67999 & n68014;
  assign n69029 = ~n68235 & ~n69028;
  assign n69030 = n68005 & ~n69029;
  assign n69031 = ~n68063 & ~n69030;
  assign n69032 = ~n68035 & ~n69012;
  assign n69033 = n67999 & n68068;
  assign n69034 = ~n68244 & ~n69033;
  assign n69035 = ~n69020 & n69034;
  assign n69036 = ~n68005 & ~n69035;
  assign n69037 = ~n67999 & n68015;
  assign n69038 = ~n69036 & ~n69037;
  assign n69039 = n69032 & n69038;
  assign n69040 = n69031 & n69039;
  assign n69041 = ~n67980 & ~n69040;
  assign n69042 = ~n68049 & ~n68864;
  assign n69043 = ~n68005 & ~n69042;
  assign n69044 = ~n69041 & ~n69043;
  assign n69045 = n69027 & n69044;
  assign n69046 = pi2041 & n69045;
  assign n69047 = ~pi2041 & ~n69045;
  assign po2124 = n69046 | n69047;
  assign n69049 = pi6751 & ~pi9040;
  assign n69050 = pi6748 & pi9040;
  assign n69051 = ~n69049 & ~n69050;
  assign n69052 = pi1993 & n69051;
  assign n69053 = ~pi1993 & ~n69051;
  assign n69054 = ~n69052 & ~n69053;
  assign n69055 = pi6723 & ~pi9040;
  assign n69056 = pi6772 & pi9040;
  assign n69057 = ~n69055 & ~n69056;
  assign n69058 = ~pi1978 & n69057;
  assign n69059 = pi1978 & ~n69057;
  assign n69060 = ~n69058 & ~n69059;
  assign n69061 = pi6748 & ~pi9040;
  assign n69062 = pi6755 & pi9040;
  assign n69063 = ~n69061 & ~n69062;
  assign n69064 = pi1997 & n69063;
  assign n69065 = ~pi1997 & ~n69063;
  assign n69066 = ~n69064 & ~n69065;
  assign n69067 = pi6859 & ~pi9040;
  assign n69068 = pi6747 & pi9040;
  assign n69069 = ~n69067 & ~n69068;
  assign n69070 = ~pi2000 & n69069;
  assign n69071 = pi2000 & ~n69069;
  assign n69072 = ~n69070 & ~n69071;
  assign n69073 = pi6771 & ~pi9040;
  assign n69074 = pi6849 & pi9040;
  assign n69075 = ~n69073 & ~n69074;
  assign n69076 = ~pi2011 & ~n69075;
  assign n69077 = pi2011 & n69075;
  assign n69078 = ~n69076 & ~n69077;
  assign n69079 = n69072 & n69078;
  assign n69080 = n69066 & n69079;
  assign n69081 = ~n69060 & n69080;
  assign n69082 = ~n69054 & n69081;
  assign n69083 = ~n69072 & ~n69078;
  assign n69084 = ~n69054 & ~n69060;
  assign n69085 = n69083 & n69084;
  assign n69086 = ~n69066 & n69085;
  assign n69087 = ~n69082 & ~n69086;
  assign n69088 = ~n69066 & n69079;
  assign n69089 = ~n69054 & n69060;
  assign n69090 = n69088 & n69089;
  assign n69091 = ~n69066 & n69083;
  assign n69092 = ~n69054 & n69091;
  assign n69093 = ~n69090 & ~n69092;
  assign n69094 = n69066 & ~n69072;
  assign n69095 = n69054 & n69094;
  assign n69096 = n69054 & n69079;
  assign n69097 = ~n69095 & ~n69096;
  assign n69098 = ~n69060 & ~n69097;
  assign n69099 = ~n69072 & n69078;
  assign n69100 = n69072 & ~n69078;
  assign n69101 = ~n69099 & ~n69100;
  assign n69102 = ~n69054 & ~n69066;
  assign n69103 = n69060 & ~n69102;
  assign n69104 = ~n69101 & n69103;
  assign n69105 = ~n69054 & ~n69079;
  assign n69106 = ~n69060 & n69105;
  assign n69107 = ~n69066 & n69106;
  assign n69108 = ~n69104 & ~n69107;
  assign n69109 = ~n69098 & n69108;
  assign n69110 = n69093 & n69109;
  assign n69111 = pi6756 & pi9040;
  assign n69112 = pi6755 & ~pi9040;
  assign n69113 = ~n69111 & ~n69112;
  assign n69114 = ~pi1990 & ~n69113;
  assign n69115 = pi1990 & n69113;
  assign n69116 = ~n69114 & ~n69115;
  assign n69117 = ~n69110 & n69116;
  assign n69118 = n69087 & ~n69117;
  assign n69119 = n69066 & n69099;
  assign n69120 = n69060 & n69119;
  assign n69121 = n69054 & n69120;
  assign n69122 = n69060 & ~n69116;
  assign n69123 = n69066 & n69083;
  assign n69124 = ~n69096 & ~n69123;
  assign n69125 = ~n69101 & n69102;
  assign n69126 = n69124 & ~n69125;
  assign n69127 = n69122 & ~n69126;
  assign n69128 = n69054 & n69091;
  assign n69129 = n69054 & ~n69072;
  assign n69130 = ~n69066 & n69129;
  assign n69131 = n69054 & n69100;
  assign n69132 = ~n69130 & ~n69131;
  assign n69133 = ~n69054 & n69079;
  assign n69134 = n69066 & n69100;
  assign n69135 = ~n69133 & ~n69134;
  assign n69136 = n69132 & n69135;
  assign n69137 = ~n69060 & ~n69136;
  assign n69138 = ~n69128 & ~n69137;
  assign n69139 = ~n69116 & ~n69138;
  assign n69140 = ~n69127 & ~n69139;
  assign n69141 = ~n69121 & n69140;
  assign n69142 = n69118 & n69141;
  assign n69143 = pi2034 & ~n69142;
  assign n69144 = ~pi2034 & n69118;
  assign n69145 = n69141 & n69144;
  assign po2125 = n69143 | n69145;
  assign n69147 = ~n69131 & ~n69133;
  assign n69148 = ~n69060 & ~n69147;
  assign n69149 = ~n69086 & ~n69148;
  assign n69150 = n69116 & ~n69149;
  assign n69151 = ~n69066 & ~n69072;
  assign n69152 = ~n69099 & ~n69151;
  assign n69153 = ~n69054 & ~n69152;
  assign n69154 = ~n69080 & ~n69153;
  assign n69155 = n69060 & ~n69154;
  assign n69156 = ~n69125 & ~n69155;
  assign n69157 = n69054 & n69088;
  assign n69158 = ~n69054 & n69066;
  assign n69159 = ~n69078 & n69158;
  assign n69160 = n69054 & ~n69152;
  assign n69161 = ~n69159 & ~n69160;
  assign n69162 = ~n69060 & ~n69161;
  assign n69163 = ~n69157 & ~n69162;
  assign n69164 = n69156 & n69163;
  assign n69165 = ~n69116 & ~n69164;
  assign n69166 = n69054 & n69066;
  assign n69167 = ~n69099 & n69166;
  assign n69168 = n69116 & n69167;
  assign n69169 = n69054 & ~n69066;
  assign n69170 = n69099 & n69169;
  assign n69171 = ~n69060 & n69170;
  assign n69172 = n69054 & n69060;
  assign n69173 = n69066 & n69172;
  assign n69174 = ~n69078 & n69173;
  assign n69175 = ~n69171 & ~n69174;
  assign n69176 = ~n69168 & n69175;
  assign n69177 = ~n69129 & ~n69134;
  assign n69178 = n69060 & n69116;
  assign n69179 = ~n69177 & n69178;
  assign n69180 = n69176 & ~n69179;
  assign n69181 = ~n69165 & n69180;
  assign n69182 = ~n69150 & n69181;
  assign n69183 = pi2048 & ~n69182;
  assign n69184 = ~pi2048 & n69182;
  assign po2126 = n69183 | n69184;
  assign n69186 = ~n68655 & ~n68674;
  assign n69187 = ~n68699 & ~n68714;
  assign n69188 = n69186 & ~n69187;
  assign n69189 = ~n68655 & n68680;
  assign n69190 = n68699 & n69189;
  assign n69191 = ~n69188 & ~n69190;
  assign n69192 = n68692 & ~n69191;
  assign n69193 = n68674 & n68697;
  assign n69194 = n68674 & ~n68680;
  assign n69195 = ~n68731 & ~n69194;
  assign n69196 = n68655 & ~n69195;
  assign n69197 = n68674 & n68680;
  assign n69198 = ~n68667 & n69197;
  assign n69199 = n68661 & n69198;
  assign n69200 = ~n69196 & ~n69199;
  assign n69201 = ~n69193 & n69200;
  assign n69202 = n68692 & ~n69201;
  assign n69203 = ~n69192 & ~n69202;
  assign n69204 = n68667 & n68681;
  assign n69205 = ~n68661 & n69204;
  assign n69206 = n68674 & n68706;
  assign n69207 = ~n69205 & ~n69206;
  assign n69208 = ~n68655 & ~n69207;
  assign n69209 = ~n68674 & n68722;
  assign n69210 = n68674 & n68731;
  assign n69211 = ~n69209 & ~n69210;
  assign n69212 = n68655 & ~n69211;
  assign n69213 = ~n68668 & ~n68731;
  assign n69214 = ~n68674 & ~n69213;
  assign n69215 = ~n68706 & ~n69214;
  assign n69216 = ~n68655 & ~n69215;
  assign n69217 = n68667 & n68674;
  assign n69218 = n69189 & n69217;
  assign n69219 = ~n68667 & ~n68680;
  assign n69220 = ~n68706 & ~n69219;
  assign n69221 = n68674 & ~n69220;
  assign n69222 = n68655 & ~n68674;
  assign n69223 = n68696 & n69222;
  assign n69224 = n68680 & n69223;
  assign n69225 = ~n69221 & ~n69224;
  assign n69226 = ~n69218 & n69225;
  assign n69227 = ~n69216 & n69226;
  assign n69228 = ~n69205 & n69227;
  assign n69229 = ~n68692 & ~n69228;
  assign n69230 = ~n69212 & ~n69229;
  assign n69231 = ~n69208 & n69230;
  assign n69232 = n69203 & n69231;
  assign n69233 = pi2029 & n69232;
  assign n69234 = ~pi2029 & ~n69232;
  assign po2127 = n69233 | n69234;
  assign n69236 = ~n68269 & n68974;
  assign n69237 = ~n68289 & ~n68302;
  assign n69238 = n68269 & n68291;
  assign n69239 = ~n68269 & n68341;
  assign n69240 = ~n69238 & ~n69239;
  assign n69241 = n69237 & n69240;
  assign n69242 = n68263 & ~n69241;
  assign n69243 = n68269 & n68310;
  assign n69244 = ~n68309 & ~n69243;
  assign n69245 = ~n68978 & n69244;
  assign n69246 = ~n68263 & ~n69245;
  assign n69247 = n68287 & n68294;
  assign n69248 = ~n68281 & n69247;
  assign n69249 = ~n69246 & ~n69248;
  assign n69250 = ~n69242 & n69249;
  assign n69251 = ~n69236 & n69250;
  assign n69252 = ~n68308 & ~n69251;
  assign n69253 = n68263 & n68269;
  assign n69254 = n68315 & n69253;
  assign n69255 = n68263 & n68978;
  assign n69256 = n68263 & n68333;
  assign n69257 = ~n69255 & ~n69256;
  assign n69258 = ~n68269 & ~n69257;
  assign n69259 = ~n69254 & ~n69258;
  assign n69260 = ~n68269 & n68292;
  assign n69261 = ~n68985 & ~n69260;
  assign n69262 = n68269 & n68288;
  assign n69263 = ~n68269 & n68310;
  assign n69264 = ~n69262 & ~n69263;
  assign n69265 = ~n68292 & n69264;
  assign n69266 = ~n68289 & n69265;
  assign n69267 = ~n68263 & ~n69266;
  assign n69268 = ~n68269 & n68311;
  assign n69269 = ~n69267 & ~n69268;
  assign n69270 = n69261 & n69269;
  assign n69271 = n69259 & n69270;
  assign n69272 = n68308 & ~n69271;
  assign n69273 = n68263 & ~n68977;
  assign n69274 = ~n69272 & ~n69273;
  assign n69275 = ~n68296 & ~n69260;
  assign n69276 = ~n68263 & ~n69275;
  assign n69277 = n69274 & ~n69276;
  assign n69278 = ~n69252 & n69277;
  assign n69279 = pi2016 & ~n69278;
  assign n69280 = ~pi2016 & n69278;
  assign po2128 = n69279 | n69280;
  assign n69282 = ~n68413 & ~n68421;
  assign n69283 = n68363 & ~n69282;
  assign n69284 = ~n68426 & ~n68573;
  assign n69285 = ~n68389 & n69284;
  assign n69286 = ~n68396 & ~n69285;
  assign n69287 = n68363 & n69286;
  assign n69288 = ~n69283 & ~n69287;
  assign n69289 = n68412 & n68576;
  assign n69290 = ~n68578 & ~n69289;
  assign n69291 = ~n68429 & ~n68602;
  assign n69292 = n68396 & ~n69291;
  assign n69293 = n68363 & n69292;
  assign n69294 = n69290 & ~n69293;
  assign n69295 = n68369 & n68412;
  assign n69296 = n68369 & n68404;
  assign n69297 = ~n68569 & ~n69296;
  assign n69298 = n68396 & ~n69297;
  assign n69299 = ~n68427 & ~n68581;
  assign n69300 = n68369 & n68411;
  assign n69301 = ~n68451 & ~n69300;
  assign n69302 = ~n68396 & ~n69301;
  assign n69303 = n69299 & ~n69302;
  assign n69304 = ~n69298 & n69303;
  assign n69305 = ~n69295 & n69304;
  assign n69306 = ~n68363 & ~n69305;
  assign n69307 = ~n68599 & n68744;
  assign n69308 = n68396 & ~n69307;
  assign n69309 = ~n69306 & ~n69308;
  assign n69310 = n69294 & n69309;
  assign n69311 = n69288 & n69310;
  assign n69312 = ~pi2030 & ~n69311;
  assign n69313 = pi2030 & n69294;
  assign n69314 = n69288 & n69313;
  assign n69315 = n69309 & n69314;
  assign po2129 = n69312 | n69315;
  assign n69317 = n68490 & n68522;
  assign n69318 = ~n68909 & ~n69317;
  assign n69319 = ~n68496 & ~n69318;
  assign n69320 = n68519 & n68905;
  assign n69321 = ~n69319 & ~n69320;
  assign n69322 = ~n68543 & n69321;
  assign n69323 = n68471 & n68496;
  assign n69324 = n68483 & n69323;
  assign n69325 = ~n68477 & n69324;
  assign n69326 = n68490 & n69325;
  assign n69327 = n68496 & n68918;
  assign n69328 = ~n68515 & ~n68541;
  assign n69329 = ~n68506 & n69328;
  assign n69330 = ~n69327 & n69329;
  assign n69331 = n68465 & ~n69330;
  assign n69332 = ~n68490 & n68552;
  assign n69333 = ~n69325 & ~n69332;
  assign n69334 = ~n68908 & n69333;
  assign n69335 = n68483 & n68513;
  assign n69336 = ~n68490 & n68501;
  assign n69337 = ~n68518 & ~n69336;
  assign n69338 = ~n68496 & ~n69337;
  assign n69339 = ~n69335 & ~n69338;
  assign n69340 = n69334 & n69339;
  assign n69341 = ~n68465 & ~n69340;
  assign n69342 = ~n68490 & n68527;
  assign n69343 = ~n68522 & ~n69342;
  assign n69344 = ~n68920 & n69343;
  assign n69345 = ~n68496 & ~n69344;
  assign n69346 = n68465 & n69345;
  assign n69347 = ~n69341 & ~n69346;
  assign n69348 = ~n69331 & n69347;
  assign n69349 = ~n69326 & n69348;
  assign n69350 = n69322 & n69349;
  assign n69351 = pi2050 & ~n69350;
  assign n69352 = ~pi2050 & n69322;
  assign n69353 = n69349 & n69352;
  assign po2130 = n69351 | n69353;
  assign n69355 = ~n67962 & ~n68809;
  assign n69356 = n67880 & ~n69355;
  assign n69357 = ~n67945 & n67947;
  assign n69358 = ~n67880 & n69357;
  assign n69359 = n67892 & n68832;
  assign n69360 = ~n68799 & ~n69359;
  assign n69361 = ~n67916 & n69360;
  assign n69362 = n67880 & ~n69361;
  assign n69363 = ~n67906 & n67922;
  assign n69364 = ~n69362 & ~n69363;
  assign n69365 = ~n67945 & ~n69364;
  assign n69366 = ~n69358 & ~n69365;
  assign n69367 = ~n67910 & ~n67914;
  assign n69368 = ~n67906 & n68797;
  assign n69369 = ~n68777 & ~n69368;
  assign n69370 = n69367 & n69369;
  assign n69371 = ~n67880 & ~n69370;
  assign n69372 = ~n67886 & ~n67892;
  assign n69373 = ~n67880 & n69372;
  assign n69374 = n67906 & n69373;
  assign n69375 = ~n67906 & n68799;
  assign n69376 = ~n67914 & ~n69375;
  assign n69377 = ~n68806 & n69376;
  assign n69378 = ~n69374 & n69377;
  assign n69379 = n67880 & n68793;
  assign n69380 = n69378 & ~n69379;
  assign n69381 = n67945 & ~n69380;
  assign n69382 = ~n69371 & ~n69381;
  assign n69383 = n69366 & n69382;
  assign n69384 = ~n69356 & n69383;
  assign n69385 = pi2063 & n69384;
  assign n69386 = ~pi2063 & ~n69384;
  assign po2131 = n69385 | n69386;
  assign n69388 = n69078 & n69158;
  assign n69389 = ~n69091 & ~n69119;
  assign n69390 = ~n69388 & n69389;
  assign n69391 = n69178 & ~n69390;
  assign n69392 = n69054 & n69116;
  assign n69393 = n69134 & n69392;
  assign n69394 = ~n69060 & n69123;
  assign n69395 = ~n69066 & n69078;
  assign n69396 = ~n69096 & ~n69395;
  assign n69397 = ~n69060 & ~n69396;
  assign n69398 = ~n69394 & ~n69397;
  assign n69399 = n69116 & ~n69398;
  assign n69400 = ~n69393 & ~n69399;
  assign n69401 = n69078 & n69169;
  assign n69402 = ~n69054 & n69100;
  assign n69403 = ~n69066 & n69402;
  assign n69404 = ~n69401 & ~n69403;
  assign n69405 = ~n69060 & ~n69404;
  assign n69406 = n69400 & ~n69405;
  assign n69407 = n69079 & n69172;
  assign n69408 = n69066 & n69407;
  assign n69409 = ~n69101 & n69169;
  assign n69410 = n69054 & n69123;
  assign n69411 = ~n69409 & ~n69410;
  assign n69412 = ~n69101 & n69158;
  assign n69413 = ~n69092 & ~n69412;
  assign n69414 = n69411 & n69413;
  assign n69415 = ~n69090 & n69414;
  assign n69416 = ~n69408 & n69415;
  assign n69417 = n69066 & n69084;
  assign n69418 = n69072 & n69417;
  assign n69419 = n69416 & ~n69418;
  assign n69420 = ~n69116 & ~n69419;
  assign n69421 = n69406 & ~n69420;
  assign n69422 = ~n69391 & n69421;
  assign n69423 = ~pi2042 & ~n69422;
  assign n69424 = pi2042 & n69406;
  assign n69425 = ~n69391 & n69424;
  assign n69426 = ~n69420 & n69425;
  assign po2132 = n69423 | n69426;
  assign n69428 = ~n68490 & n68932;
  assign n69429 = ~n68526 & ~n68918;
  assign n69430 = ~n68496 & ~n69429;
  assign n69431 = ~n69428 & ~n69430;
  assign n69432 = n68483 & n68907;
  assign n69433 = ~n68555 & ~n69432;
  assign n69434 = ~n68920 & n69433;
  assign n69435 = n68496 & ~n69434;
  assign n69436 = n69431 & ~n69435;
  assign n69437 = n68490 & n68519;
  assign n69438 = n69436 & ~n69437;
  assign n69439 = ~n68465 & ~n69438;
  assign n69440 = n68500 & ~n69429;
  assign n69441 = ~n68522 & ~n68527;
  assign n69442 = ~n68519 & ~n68920;
  assign n69443 = n69441 & n69442;
  assign n69444 = ~n68490 & ~n69443;
  assign n69445 = ~n69440 & ~n69444;
  assign n69446 = ~n68909 & n69445;
  assign n69447 = n68465 & ~n69446;
  assign n69448 = ~n69439 & ~n69447;
  assign n69449 = ~n68490 & n68918;
  assign n69450 = ~n69437 & ~n69449;
  assign n69451 = ~n68496 & ~n69450;
  assign n69452 = n69448 & ~n69451;
  assign n69453 = pi2033 & ~n69452;
  assign n69454 = ~pi2033 & ~n69451;
  assign n69455 = ~n69447 & n69454;
  assign n69456 = ~n69439 & n69455;
  assign po2133 = n69453 | n69456;
  assign n69458 = ~n69066 & n69099;
  assign n69459 = ~n69080 & ~n69458;
  assign n69460 = ~n69060 & ~n69459;
  assign n69461 = ~n69119 & ~n69402;
  assign n69462 = ~n69088 & n69461;
  assign n69463 = n69060 & ~n69462;
  assign n69464 = ~n69460 & ~n69463;
  assign n69465 = ~n69394 & ~n69403;
  assign n69466 = n69464 & n69465;
  assign n69467 = ~n69116 & ~n69466;
  assign n69468 = n69054 & n69080;
  assign n69469 = ~n69054 & n69083;
  assign n69470 = ~n69131 & ~n69469;
  assign n69471 = n69060 & ~n69470;
  assign n69472 = ~n69468 & ~n69471;
  assign n69473 = ~n69060 & n69066;
  assign n69474 = ~n69078 & n69473;
  assign n69475 = n69072 & n69474;
  assign n69476 = n69389 & ~n69475;
  assign n69477 = ~n69088 & n69476;
  assign n69478 = ~n69054 & ~n69477;
  assign n69479 = n69472 & ~n69478;
  assign n69480 = n69116 & ~n69479;
  assign n69481 = ~n69467 & ~n69480;
  assign n69482 = ~n69066 & n69131;
  assign n69483 = ~n69410 & ~n69482;
  assign n69484 = ~n69060 & ~n69483;
  assign n69485 = n69060 & n69151;
  assign n69486 = n69054 & n69485;
  assign n69487 = ~n69484 & ~n69486;
  assign n69488 = n69481 & n69487;
  assign n69489 = ~pi2026 & ~n69488;
  assign n69490 = pi2026 & ~n69484;
  assign n69491 = n69481 & n69490;
  assign n69492 = ~n69486 & n69491;
  assign po2134 = n69489 | n69492;
  assign n69494 = ~n68667 & n68683;
  assign n69495 = ~n68714 & ~n69494;
  assign n69496 = ~n68655 & ~n69495;
  assign n69497 = ~n68674 & n68705;
  assign n69498 = ~n68667 & n68674;
  assign n69499 = n68680 & n69498;
  assign n69500 = ~n69497 & ~n69499;
  assign n69501 = n68655 & ~n69500;
  assign n69502 = n68674 & n68700;
  assign n69503 = ~n69218 & ~n69502;
  assign n69504 = ~n68682 & n69503;
  assign n69505 = ~n69501 & n69504;
  assign n69506 = ~n69496 & n69505;
  assign n69507 = ~n69193 & ~n69205;
  assign n69508 = n69506 & n69507;
  assign n69509 = n68692 & ~n69508;
  assign n69510 = n68668 & n69194;
  assign n69511 = n68723 & ~n69510;
  assign n69512 = n68655 & ~n69511;
  assign n69513 = n68674 & n68711;
  assign n69514 = ~n69512 & ~n69513;
  assign n69515 = n68661 & n68683;
  assign n69516 = ~n68674 & n68696;
  assign n69517 = ~n69515 & ~n69516;
  assign n69518 = n68655 & ~n69517;
  assign n69519 = n68655 & n68705;
  assign n69520 = n68674 & n69519;
  assign n69521 = ~n69518 & ~n69520;
  assign n69522 = n69514 & n69521;
  assign n69523 = ~n68692 & ~n69522;
  assign n69524 = ~n68700 & ~n68707;
  assign n69525 = ~n69199 & n69524;
  assign n69526 = n68728 & ~n69525;
  assign n69527 = ~n69523 & ~n69526;
  assign n69528 = ~n68682 & ~n69193;
  assign n69529 = ~n68655 & ~n69528;
  assign n69530 = n69527 & ~n69529;
  assign n69531 = ~n69509 & n69530;
  assign n69532 = ~pi2035 & n69531;
  assign n69533 = pi2035 & ~n69531;
  assign po2135 = n69532 | n69533;
  assign n69535 = ~n68979 & ~n69260;
  assign n69536 = ~n69248 & n69535;
  assign n69537 = n68263 & ~n69536;
  assign n69538 = ~n68988 & ~n69004;
  assign n69539 = ~n68985 & ~n69256;
  assign n69540 = ~n68974 & ~n69263;
  assign n69541 = ~n68263 & ~n69540;
  assign n69542 = ~n68302 & ~n69541;
  assign n69543 = n69539 & n69542;
  assign n69544 = n68308 & ~n69543;
  assign n69545 = ~n68275 & n68287;
  assign n69546 = ~n68316 & ~n69545;
  assign n69547 = n68269 & ~n69546;
  assign n69548 = ~n68292 & ~n68991;
  assign n69549 = ~n68263 & ~n69548;
  assign n69550 = n68269 & n68287;
  assign n69551 = ~n68311 & ~n69550;
  assign n69552 = ~n68319 & n69551;
  assign n69553 = n68263 & ~n69552;
  assign n69554 = ~n69549 & ~n69553;
  assign n69555 = ~n69547 & n69554;
  assign n69556 = ~n68308 & ~n69555;
  assign n69557 = ~n69544 & ~n69556;
  assign n69558 = n69538 & n69557;
  assign n69559 = ~n69537 & n69558;
  assign n69560 = ~pi2025 & ~n69559;
  assign n69561 = pi2025 & n69538;
  assign n69562 = ~n69537 & n69561;
  assign n69563 = n69557 & n69562;
  assign po2136 = n69560 | n69563;
  assign n69565 = n68674 & n68696;
  assign n69566 = ~n68695 & ~n69565;
  assign n69567 = ~n68655 & ~n69566;
  assign n69568 = n68655 & ~n69220;
  assign n69569 = ~n69209 & ~n69568;
  assign n69570 = ~n69567 & n69569;
  assign n69571 = n68692 & ~n69570;
  assign n69572 = ~n68655 & n68711;
  assign n69573 = ~n69571 & ~n69572;
  assign n69574 = ~n69502 & ~n69516;
  assign n69575 = n68655 & ~n69574;
  assign n69576 = n68655 & n68697;
  assign n69577 = ~n68674 & n68714;
  assign n69578 = ~n68655 & n68681;
  assign n69579 = ~n69197 & ~n69578;
  assign n69580 = ~n68661 & ~n69579;
  assign n69581 = ~n69499 & ~n69580;
  assign n69582 = ~n68682 & n69581;
  assign n69583 = ~n69577 & n69582;
  assign n69584 = ~n69576 & n69583;
  assign n69585 = ~n68692 & ~n69584;
  assign n69586 = ~n69575 & ~n69585;
  assign n69587 = n69573 & n69586;
  assign n69588 = pi2057 & ~n69587;
  assign n69589 = ~pi2057 & n69587;
  assign po2137 = n69588 | n69589;
  assign n69591 = pi6980 & ~pi9040;
  assign n69592 = pi7002 & pi9040;
  assign n69593 = ~n69591 & ~n69592;
  assign n69594 = ~pi2076 & ~n69593;
  assign n69595 = pi2076 & n69593;
  assign n69596 = ~n69594 & ~n69595;
  assign n69597 = pi6960 & ~pi9040;
  assign n69598 = pi7084 & pi9040;
  assign n69599 = ~n69597 & ~n69598;
  assign n69600 = ~pi2074 & ~n69599;
  assign n69601 = pi2074 & n69599;
  assign n69602 = ~n69600 & ~n69601;
  assign n69603 = ~n69596 & ~n69602;
  assign n69604 = pi6958 & ~pi9040;
  assign n69605 = pi6979 & pi9040;
  assign n69606 = ~n69604 & ~n69605;
  assign n69607 = pi2061 & n69606;
  assign n69608 = ~pi2061 & ~n69606;
  assign n69609 = ~n69607 & ~n69608;
  assign n69610 = pi6956 & pi9040;
  assign n69611 = pi6946 & ~pi9040;
  assign n69612 = ~n69610 & ~n69611;
  assign n69613 = ~pi2065 & ~n69612;
  assign n69614 = pi2065 & n69612;
  assign n69615 = ~n69613 & ~n69614;
  assign n69616 = pi6960 & pi9040;
  assign n69617 = pi6975 & ~pi9040;
  assign n69618 = ~n69616 & ~n69617;
  assign n69619 = ~pi2043 & n69618;
  assign n69620 = pi2043 & ~n69618;
  assign n69621 = ~n69619 & ~n69620;
  assign n69622 = n69615 & n69621;
  assign n69623 = ~n69609 & n69622;
  assign n69624 = pi6958 & pi9040;
  assign n69625 = pi7002 & ~pi9040;
  assign n69626 = ~n69624 & ~n69625;
  assign n69627 = ~pi2037 & ~n69626;
  assign n69628 = pi2037 & n69626;
  assign n69629 = ~n69627 & ~n69628;
  assign n69630 = ~n69621 & ~n69629;
  assign n69631 = n69615 & n69630;
  assign n69632 = n69609 & n69631;
  assign n69633 = ~n69621 & n69629;
  assign n69634 = ~n69609 & n69633;
  assign n69635 = ~n69632 & ~n69634;
  assign n69636 = ~n69623 & n69635;
  assign n69637 = n69603 & ~n69636;
  assign n69638 = ~n69609 & ~n69615;
  assign n69639 = ~n69629 & n69638;
  assign n69640 = n69622 & ~n69629;
  assign n69641 = n69609 & n69640;
  assign n69642 = ~n69639 & ~n69641;
  assign n69643 = ~n69615 & n69630;
  assign n69644 = n69615 & n69633;
  assign n69645 = ~n69643 & ~n69644;
  assign n69646 = n69642 & n69645;
  assign n69647 = n69596 & ~n69646;
  assign n69648 = n69621 & n69629;
  assign n69649 = ~n69615 & n69648;
  assign n69650 = n69609 & n69649;
  assign n69651 = ~n69647 & ~n69650;
  assign n69652 = ~n69602 & ~n69651;
  assign n69653 = ~n69637 & ~n69652;
  assign n69654 = n69596 & ~n69609;
  assign n69655 = n69615 & n69654;
  assign n69656 = n69629 & n69655;
  assign n69657 = ~n69609 & n69643;
  assign n69658 = ~n69656 & ~n69657;
  assign n69659 = n69621 & ~n69629;
  assign n69660 = ~n69633 & ~n69659;
  assign n69661 = n69609 & ~n69660;
  assign n69662 = ~n69615 & n69659;
  assign n69663 = ~n69661 & ~n69662;
  assign n69664 = ~n69596 & ~n69663;
  assign n69665 = n69615 & n69648;
  assign n69666 = ~n69623 & ~n69665;
  assign n69667 = ~n69632 & n69666;
  assign n69668 = n69596 & ~n69667;
  assign n69669 = ~n69664 & ~n69668;
  assign n69670 = ~n69596 & ~n69609;
  assign n69671 = n69630 & n69670;
  assign n69672 = n69609 & ~n69615;
  assign n69673 = ~n69629 & n69672;
  assign n69674 = n69621 & n69673;
  assign n69675 = ~n69615 & ~n69621;
  assign n69676 = n69629 & n69675;
  assign n69677 = n69609 & n69676;
  assign n69678 = ~n69674 & ~n69677;
  assign n69679 = n69629 & n69638;
  assign n69680 = n69621 & n69679;
  assign n69681 = n69678 & ~n69680;
  assign n69682 = ~n69671 & n69681;
  assign n69683 = n69669 & n69682;
  assign n69684 = n69602 & ~n69683;
  assign n69685 = n69658 & ~n69684;
  assign n69686 = n69653 & n69685;
  assign n69687 = pi2153 & ~n69686;
  assign n69688 = ~pi2153 & n69658;
  assign n69689 = n69653 & n69688;
  assign n69690 = ~n69684 & n69689;
  assign po2158 = n69687 | n69690;
  assign n69692 = pi6984 & pi9040;
  assign n69693 = pi7084 & ~pi9040;
  assign n69694 = ~n69692 & ~n69693;
  assign n69695 = ~pi2066 & ~n69694;
  assign n69696 = pi2066 & n69694;
  assign n69697 = ~n69695 & ~n69696;
  assign n69698 = pi6980 & pi9040;
  assign n69699 = pi7009 & ~pi9040;
  assign n69700 = ~n69698 & ~n69699;
  assign n69701 = pi2049 & n69700;
  assign n69702 = ~pi2049 & ~n69700;
  assign n69703 = ~n69701 & ~n69702;
  assign n69704 = pi7083 & pi9040;
  assign n69705 = pi6982 & ~pi9040;
  assign n69706 = ~n69704 & ~n69705;
  assign n69707 = ~pi2060 & n69706;
  assign n69708 = pi2060 & ~n69706;
  assign n69709 = ~n69707 & ~n69708;
  assign n69710 = pi6973 & ~pi9040;
  assign n69711 = pi7005 & pi9040;
  assign n69712 = ~n69710 & ~n69711;
  assign n69713 = ~pi2055 & n69712;
  assign n69714 = pi2055 & ~n69712;
  assign n69715 = ~n69713 & ~n69714;
  assign n69716 = ~n69709 & ~n69715;
  assign n69717 = ~n69703 & n69716;
  assign n69718 = pi7004 & pi9040;
  assign n69719 = pi6993 & ~pi9040;
  assign n69720 = ~n69718 & ~n69719;
  assign n69721 = pi2075 & n69720;
  assign n69722 = ~pi2075 & ~n69720;
  assign n69723 = ~n69721 & ~n69722;
  assign n69724 = n69717 & ~n69723;
  assign n69725 = n69709 & n69715;
  assign n69726 = ~n69703 & ~n69723;
  assign n69727 = n69725 & n69726;
  assign n69728 = ~n69724 & ~n69727;
  assign n69729 = n69703 & n69725;
  assign n69730 = n69723 & n69729;
  assign n69731 = ~n69709 & n69715;
  assign n69732 = ~n69703 & n69731;
  assign n69733 = n69723 & n69732;
  assign n69734 = ~n69730 & ~n69733;
  assign n69735 = n69728 & n69734;
  assign n69736 = n69697 & ~n69735;
  assign n69737 = n69709 & ~n69715;
  assign n69738 = ~n69703 & n69737;
  assign n69739 = n69723 & n69738;
  assign n69740 = ~n69732 & ~n69739;
  assign n69741 = n69697 & ~n69740;
  assign n69742 = ~n69697 & ~n69715;
  assign n69743 = ~n69723 & n69742;
  assign n69744 = n69703 & ~n69709;
  assign n69745 = n69723 & n69725;
  assign n69746 = ~n69744 & ~n69745;
  assign n69747 = ~n69697 & ~n69746;
  assign n69748 = ~n69743 & ~n69747;
  assign n69749 = n69703 & n69737;
  assign n69750 = ~n69723 & n69749;
  assign n69751 = n69748 & ~n69750;
  assign n69752 = ~n69715 & n69744;
  assign n69753 = n69723 & n69752;
  assign n69754 = n69751 & ~n69753;
  assign n69755 = ~n69741 & n69754;
  assign n69756 = pi6982 & pi9040;
  assign n69757 = pi6978 & ~pi9040;
  assign n69758 = ~n69756 & ~n69757;
  assign n69759 = ~pi2077 & ~n69758;
  assign n69760 = pi2077 & n69758;
  assign n69761 = ~n69759 & ~n69760;
  assign n69762 = ~n69755 & ~n69761;
  assign n69763 = ~n69703 & ~n69715;
  assign n69764 = ~n69697 & n69723;
  assign n69765 = n69761 & n69764;
  assign n69766 = n69763 & n69765;
  assign n69767 = n69715 & n69726;
  assign n69768 = ~n69697 & ~n69767;
  assign n69769 = n69703 & n69723;
  assign n69770 = n69709 & n69769;
  assign n69771 = ~n69716 & ~n69763;
  assign n69772 = ~n69723 & ~n69771;
  assign n69773 = n69697 & ~n69729;
  assign n69774 = ~n69772 & n69773;
  assign n69775 = ~n69770 & n69774;
  assign n69776 = ~n69768 & ~n69775;
  assign n69777 = n69703 & n69731;
  assign n69778 = n69723 & n69777;
  assign n69779 = ~n69776 & ~n69778;
  assign n69780 = n69761 & ~n69779;
  assign n69781 = ~n69766 & ~n69780;
  assign n69782 = ~n69762 & n69781;
  assign n69783 = ~n69736 & n69782;
  assign n69784 = ~n69697 & n69750;
  assign n69785 = n69783 & ~n69784;
  assign n69786 = pi2152 & ~n69785;
  assign n69787 = ~pi2152 & ~n69784;
  assign n69788 = n69782 & n69787;
  assign n69789 = ~n69736 & n69788;
  assign po2160 = n69786 | n69789;
  assign n69791 = pi6990 & ~pi9040;
  assign n69792 = pi6962 & pi9040;
  assign n69793 = ~n69791 & ~n69792;
  assign n69794 = ~pi2069 & ~n69793;
  assign n69795 = pi2069 & n69793;
  assign n69796 = ~n69794 & ~n69795;
  assign n69797 = pi6945 & pi9040;
  assign n69798 = pi7081 & ~pi9040;
  assign n69799 = ~n69797 & ~n69798;
  assign n69800 = ~pi2032 & n69799;
  assign n69801 = pi2032 & ~n69799;
  assign n69802 = ~n69800 & ~n69801;
  assign n69803 = pi7012 & pi9040;
  assign n69804 = pi6947 & ~pi9040;
  assign n69805 = ~n69803 & ~n69804;
  assign n69806 = pi2067 & n69805;
  assign n69807 = ~pi2067 & ~n69805;
  assign n69808 = ~n69806 & ~n69807;
  assign n69809 = pi6962 & ~pi9040;
  assign n69810 = pi6968 & pi9040;
  assign n69811 = ~n69809 & ~n69810;
  assign n69812 = pi2073 & n69811;
  assign n69813 = ~pi2073 & ~n69811;
  assign n69814 = ~n69812 & ~n69813;
  assign n69815 = pi6945 & ~pi9040;
  assign n69816 = pi7008 & pi9040;
  assign n69817 = ~n69815 & ~n69816;
  assign n69818 = ~pi2070 & n69817;
  assign n69819 = pi2070 & ~n69817;
  assign n69820 = ~n69818 & ~n69819;
  assign n69821 = ~n69814 & ~n69820;
  assign n69822 = n69808 & n69821;
  assign n69823 = ~n69802 & n69822;
  assign n69824 = pi7082 & pi9040;
  assign n69825 = pi7006 & ~pi9040;
  assign n69826 = ~n69824 & ~n69825;
  assign n69827 = ~pi2071 & ~n69826;
  assign n69828 = pi2071 & n69826;
  assign n69829 = ~n69827 & ~n69828;
  assign n69830 = ~pi2073 & n69811;
  assign n69831 = pi2073 & ~n69811;
  assign n69832 = ~n69830 & ~n69831;
  assign n69833 = ~n69820 & ~n69832;
  assign n69834 = ~n69802 & n69833;
  assign n69835 = ~n69808 & n69821;
  assign n69836 = n69802 & n69835;
  assign n69837 = ~n69834 & ~n69836;
  assign n69838 = ~n69829 & ~n69837;
  assign n69839 = ~n69823 & ~n69838;
  assign n69840 = ~n69814 & n69820;
  assign n69841 = ~n69808 & n69840;
  assign n69842 = n69829 & n69841;
  assign n69843 = n69821 & n69829;
  assign n69844 = ~n69802 & n69843;
  assign n69845 = ~n69842 & ~n69844;
  assign n69846 = n69839 & n69845;
  assign n69847 = n69820 & ~n69832;
  assign n69848 = n69808 & n69847;
  assign n69849 = ~n69802 & n69848;
  assign n69850 = n69808 & n69840;
  assign n69851 = n69802 & n69850;
  assign n69852 = ~n69849 & ~n69851;
  assign n69853 = n69846 & n69852;
  assign n69854 = n69796 & ~n69853;
  assign n69855 = ~n69796 & ~n69829;
  assign n69856 = ~n69802 & ~n69808;
  assign n69857 = n69832 & n69856;
  assign n69858 = ~n69808 & n69820;
  assign n69859 = ~n69857 & ~n69858;
  assign n69860 = n69855 & ~n69859;
  assign n69861 = n69802 & n69808;
  assign n69862 = ~n69820 & n69861;
  assign n69863 = ~n69814 & n69862;
  assign n69864 = n69802 & ~n69832;
  assign n69865 = ~n69808 & n69864;
  assign n69866 = ~n69863 & ~n69865;
  assign n69867 = ~n69802 & n69829;
  assign n69868 = ~n69821 & n69867;
  assign n69869 = n69808 & n69868;
  assign n69870 = n69829 & n69848;
  assign n69871 = ~n69869 & ~n69870;
  assign n69872 = n69866 & n69871;
  assign n69873 = ~n69796 & ~n69872;
  assign n69874 = ~n69808 & n69847;
  assign n69875 = ~n69829 & n69874;
  assign n69876 = n69802 & n69875;
  assign n69877 = n69808 & n69833;
  assign n69878 = n69802 & n69877;
  assign n69879 = ~n69851 & ~n69878;
  assign n69880 = ~n69829 & ~n69879;
  assign n69881 = ~n69876 & ~n69880;
  assign n69882 = n69829 & n69863;
  assign n69883 = n69881 & ~n69882;
  assign n69884 = ~n69873 & n69883;
  assign n69885 = ~n69860 & n69884;
  assign n69886 = ~n69854 & n69885;
  assign n69887 = ~n69808 & n69833;
  assign n69888 = n69802 & n69829;
  assign n69889 = n69887 & n69888;
  assign n69890 = n69886 & ~n69889;
  assign n69891 = ~pi2173 & ~n69890;
  assign n69892 = ~n69854 & ~n69889;
  assign n69893 = n69885 & n69892;
  assign n69894 = pi2173 & n69893;
  assign po2161 = n69891 | n69894;
  assign n69896 = n69609 & n69622;
  assign n69897 = ~n69644 & ~n69896;
  assign n69898 = ~n69657 & n69897;
  assign n69899 = n69596 & ~n69898;
  assign n69900 = ~n69609 & n69676;
  assign n69901 = ~n69609 & n69665;
  assign n69902 = ~n69615 & n69621;
  assign n69903 = ~n69630 & ~n69902;
  assign n69904 = n69609 & ~n69903;
  assign n69905 = ~n69901 & ~n69904;
  assign n69906 = ~n69900 & n69905;
  assign n69907 = ~n69596 & ~n69906;
  assign n69908 = ~n69899 & ~n69907;
  assign n69909 = n69602 & ~n69908;
  assign n69910 = n69621 & n69654;
  assign n69911 = ~n69609 & ~n69621;
  assign n69912 = n69615 & n69911;
  assign n69913 = ~n69896 & ~n69912;
  assign n69914 = ~n69596 & ~n69913;
  assign n69915 = ~n69671 & ~n69914;
  assign n69916 = ~n69609 & n69631;
  assign n69917 = ~n69677 & ~n69916;
  assign n69918 = n69596 & n69609;
  assign n69919 = n69675 & n69918;
  assign n69920 = n69596 & n69649;
  assign n69921 = ~n69919 & ~n69920;
  assign n69922 = n69917 & n69921;
  assign n69923 = n69915 & n69922;
  assign n69924 = ~n69910 & n69923;
  assign n69925 = ~n69602 & ~n69924;
  assign n69926 = ~n69596 & n69662;
  assign n69927 = ~n69609 & n69926;
  assign n69928 = ~n69596 & n69916;
  assign n69929 = ~n69927 & ~n69928;
  assign n69930 = n69596 & n69680;
  assign n69931 = n69929 & ~n69930;
  assign n69932 = ~n69609 & n69640;
  assign n69933 = n69609 & n69633;
  assign n69934 = ~n69932 & ~n69933;
  assign n69935 = n69596 & ~n69934;
  assign n69936 = n69931 & ~n69935;
  assign n69937 = ~n69925 & n69936;
  assign n69938 = ~n69909 & n69937;
  assign n69939 = ~pi2169 & ~n69938;
  assign n69940 = pi2169 & n69938;
  assign po2164 = n69939 | n69940;
  assign n69942 = ~n69596 & n69900;
  assign n69943 = ~n69928 & ~n69942;
  assign n69944 = ~n69930 & n69943;
  assign n69945 = ~n69662 & ~n69665;
  assign n69946 = ~n69596 & ~n69945;
  assign n69947 = n69609 & n69644;
  assign n69948 = ~n69946 & ~n69947;
  assign n69949 = n69609 & ~n69621;
  assign n69950 = ~n69675 & ~n69949;
  assign n69951 = ~n69640 & n69950;
  assign n69952 = n69596 & ~n69951;
  assign n69953 = n69948 & ~n69952;
  assign n69954 = ~n69602 & ~n69953;
  assign n69955 = ~n69609 & n69615;
  assign n69956 = ~n69629 & n69955;
  assign n69957 = ~n69680 & ~n69956;
  assign n69958 = n69596 & n69912;
  assign n69959 = n69609 & n69665;
  assign n69960 = ~n69596 & n69675;
  assign n69961 = ~n69959 & ~n69960;
  assign n69962 = ~n69674 & n69961;
  assign n69963 = ~n69958 & n69962;
  assign n69964 = n69957 & n69963;
  assign n69965 = ~n69920 & n69964;
  assign n69966 = n69602 & ~n69965;
  assign n69967 = ~n69954 & ~n69966;
  assign n69968 = n69944 & n69967;
  assign n69969 = ~pi2163 & ~n69968;
  assign n69970 = pi2163 & n69944;
  assign n69971 = ~n69954 & n69970;
  assign n69972 = ~n69966 & n69971;
  assign po2167 = n69969 | n69972;
  assign n69974 = pi6953 & pi9040;
  assign n69975 = pi6983 & ~pi9040;
  assign n69976 = ~n69974 & ~n69975;
  assign n69977 = pi2062 & n69976;
  assign n69978 = ~pi2062 & ~n69976;
  assign n69979 = ~n69977 & ~n69978;
  assign n69980 = pi7004 & ~pi9040;
  assign n69981 = pi6983 & pi9040;
  assign n69982 = ~n69980 & ~n69981;
  assign n69983 = pi2049 & n69982;
  assign n69984 = ~pi2049 & ~n69982;
  assign n69985 = ~n69983 & ~n69984;
  assign n69986 = pi6992 & pi9040;
  assign n69987 = pi6988 & ~pi9040;
  assign n69988 = ~n69986 & ~n69987;
  assign n69989 = pi2074 & n69988;
  assign n69990 = ~pi2074 & ~n69988;
  assign n69991 = ~n69989 & ~n69990;
  assign n69992 = n69985 & ~n69991;
  assign n69993 = pi6984 & ~pi9040;
  assign n69994 = pi7009 & pi9040;
  assign n69995 = ~n69993 & ~n69994;
  assign n69996 = pi2045 & n69995;
  assign n69997 = ~pi2045 & ~n69995;
  assign n69998 = ~n69996 & ~n69997;
  assign n69999 = pi6966 & pi9040;
  assign n70000 = pi7005 & ~pi9040;
  assign n70001 = ~n69999 & ~n70000;
  assign n70002 = ~pi2037 & n70001;
  assign n70003 = pi2037 & ~n70001;
  assign n70004 = ~n70002 & ~n70003;
  assign n70005 = n69998 & n70004;
  assign n70006 = n69992 & n70005;
  assign n70007 = ~n69985 & ~n69991;
  assign n70008 = ~n70004 & n70007;
  assign n70009 = n69998 & n70008;
  assign n70010 = ~n70006 & ~n70009;
  assign n70011 = ~n69985 & n69991;
  assign n70012 = n70004 & n70011;
  assign n70013 = n70010 & ~n70012;
  assign n70014 = n69979 & ~n70013;
  assign n70015 = pi6959 & pi9040;
  assign n70016 = pi7003 & ~pi9040;
  assign n70017 = ~n70015 & ~n70016;
  assign n70018 = pi2055 & n70017;
  assign n70019 = ~pi2055 & ~n70017;
  assign n70020 = ~n70018 & ~n70019;
  assign n70021 = ~n69979 & ~n69998;
  assign n70022 = n69992 & n70021;
  assign n70023 = ~n69998 & n70004;
  assign n70024 = ~n69985 & n70023;
  assign n70025 = n69991 & n70024;
  assign n70026 = ~n70004 & n70011;
  assign n70027 = ~n69991 & n70004;
  assign n70028 = ~n69985 & n70027;
  assign n70029 = n69998 & n70028;
  assign n70030 = ~n70026 & ~n70029;
  assign n70031 = n69985 & n69991;
  assign n70032 = n69998 & n70031;
  assign n70033 = n70030 & ~n70032;
  assign n70034 = ~n69979 & ~n70033;
  assign n70035 = n69991 & n70004;
  assign n70036 = n69979 & ~n69998;
  assign n70037 = n70035 & n70036;
  assign n70038 = ~n70034 & ~n70037;
  assign n70039 = ~n70025 & n70038;
  assign n70040 = ~n70022 & n70039;
  assign n70041 = ~n70004 & n70031;
  assign n70042 = n69998 & n70041;
  assign n70043 = n69992 & ~n70004;
  assign n70044 = ~n69998 & n70043;
  assign n70045 = ~n70042 & ~n70044;
  assign n70046 = n70040 & n70045;
  assign n70047 = ~n70020 & ~n70046;
  assign n70048 = ~n69985 & n70004;
  assign n70049 = n69979 & n70048;
  assign n70050 = ~n69998 & n70049;
  assign n70051 = n69991 & ~n70004;
  assign n70052 = n69998 & n70051;
  assign n70053 = ~n69991 & ~n70004;
  assign n70054 = ~n69998 & n70053;
  assign n70055 = ~n70052 & ~n70054;
  assign n70056 = ~n69979 & ~n70055;
  assign n70057 = ~n70050 & ~n70056;
  assign n70058 = n69985 & n70023;
  assign n70059 = n69991 & n70058;
  assign n70060 = ~n70043 & ~n70059;
  assign n70061 = ~n69979 & ~n70060;
  assign n70062 = ~n69991 & n70024;
  assign n70063 = ~n70006 & ~n70062;
  assign n70064 = n69991 & n70005;
  assign n70065 = ~n69998 & n70041;
  assign n70066 = ~n70064 & ~n70065;
  assign n70067 = n69979 & ~n70066;
  assign n70068 = n70063 & ~n70067;
  assign n70069 = ~n70061 & n70068;
  assign n70070 = n70020 & ~n70069;
  assign n70071 = n70057 & ~n70070;
  assign n70072 = ~n70047 & n70071;
  assign n70073 = ~n70014 & n70072;
  assign n70074 = ~pi2197 & ~n70073;
  assign n70075 = pi2197 & n70073;
  assign po2168 = n70074 | n70075;
  assign n70077 = n69802 & n69841;
  assign n70078 = n69820 & n69856;
  assign n70079 = ~n69832 & n70078;
  assign n70080 = ~n70077 & ~n70079;
  assign n70081 = n69829 & ~n70080;
  assign n70082 = ~n69863 & ~n69870;
  assign n70083 = ~n69814 & n69861;
  assign n70084 = ~n69865 & ~n70083;
  assign n70085 = ~n69829 & ~n70084;
  assign n70086 = ~n69802 & ~n69829;
  assign n70087 = n69840 & n70086;
  assign n70088 = ~n69808 & n70087;
  assign n70089 = ~n69808 & n69829;
  assign n70090 = ~n69820 & n70089;
  assign n70091 = ~n69814 & n70090;
  assign n70092 = ~n69802 & n69808;
  assign n70093 = ~n69820 & n70092;
  assign n70094 = ~n69832 & n70093;
  assign n70095 = ~n70091 & ~n70094;
  assign n70096 = ~n70088 & n70095;
  assign n70097 = ~n70085 & n70096;
  assign n70098 = n70082 & n70097;
  assign n70099 = n69796 & ~n70098;
  assign n70100 = ~n69829 & n69863;
  assign n70101 = n69802 & n69870;
  assign n70102 = ~n70100 & ~n70101;
  assign n70103 = ~n70099 & n70102;
  assign n70104 = ~n70081 & n70103;
  assign n70105 = n69808 & ~n69814;
  assign n70106 = n69867 & n70105;
  assign n70107 = ~n69842 & ~n70106;
  assign n70108 = n69829 & n69877;
  assign n70109 = n69802 & n69887;
  assign n70110 = ~n70108 & ~n70109;
  assign n70111 = ~n69802 & n69850;
  assign n70112 = ~n70077 & ~n70111;
  assign n70113 = ~n69802 & n69847;
  assign n70114 = ~n69808 & ~n69820;
  assign n70115 = ~n70113 & ~n70114;
  assign n70116 = ~n69829 & ~n70115;
  assign n70117 = n70112 & ~n70116;
  assign n70118 = n70110 & n70117;
  assign n70119 = n70107 & n70118;
  assign n70120 = ~n69796 & ~n70119;
  assign n70121 = n70104 & ~n70120;
  assign n70122 = ~pi2145 & ~n70121;
  assign n70123 = pi2145 & n70104;
  assign n70124 = ~n70120 & n70123;
  assign po2169 = n70122 | n70124;
  assign n70126 = pi6954 & pi9040;
  assign n70127 = pi6986 & ~pi9040;
  assign n70128 = ~n70126 & ~n70127;
  assign n70129 = ~pi2058 & ~n70128;
  assign n70130 = pi2058 & n70128;
  assign n70131 = ~n70129 & ~n70130;
  assign n70132 = pi6948 & ~pi9040;
  assign n70133 = pi7006 & pi9040;
  assign n70134 = ~n70132 & ~n70133;
  assign n70135 = ~pi2060 & n70134;
  assign n70136 = pi2060 & ~n70134;
  assign n70137 = ~n70135 & ~n70136;
  assign n70138 = pi6948 & pi9040;
  assign n70139 = pi7068 & ~pi9040;
  assign n70140 = ~n70138 & ~n70139;
  assign n70141 = pi2077 & n70140;
  assign n70142 = ~pi2077 & ~n70140;
  assign n70143 = ~n70141 & ~n70142;
  assign n70144 = pi6974 & pi9040;
  assign n70145 = pi7008 & ~pi9040;
  assign n70146 = ~n70144 & ~n70145;
  assign n70147 = ~pi2036 & ~n70146;
  assign n70148 = pi2036 & n70146;
  assign n70149 = ~n70147 & ~n70148;
  assign n70150 = ~n70143 & n70149;
  assign n70151 = pi7068 & pi9040;
  assign n70152 = pi6972 & ~pi9040;
  assign n70153 = ~n70151 & ~n70152;
  assign n70154 = pi2059 & n70153;
  assign n70155 = ~pi2059 & ~n70153;
  assign n70156 = ~n70154 & ~n70155;
  assign n70157 = pi6952 & ~pi9040;
  assign n70158 = pi7081 & pi9040;
  assign n70159 = ~n70157 & ~n70158;
  assign n70160 = pi2052 & n70159;
  assign n70161 = ~pi2052 & ~n70159;
  assign n70162 = ~n70160 & ~n70161;
  assign n70163 = n70156 & n70162;
  assign n70164 = n70150 & n70163;
  assign n70165 = ~n70137 & n70164;
  assign n70166 = ~n70156 & n70162;
  assign n70167 = n70143 & n70149;
  assign n70168 = n70166 & n70167;
  assign n70169 = ~n70137 & ~n70156;
  assign n70170 = ~n70149 & n70169;
  assign n70171 = ~n70143 & n70170;
  assign n70172 = n70143 & ~n70149;
  assign n70173 = ~n70137 & n70172;
  assign n70174 = n70162 & n70173;
  assign n70175 = n70156 & n70174;
  assign n70176 = ~n70171 & ~n70175;
  assign n70177 = ~n70168 & n70176;
  assign n70178 = ~n70165 & n70177;
  assign n70179 = n70137 & ~n70156;
  assign n70180 = n70149 & n70179;
  assign n70181 = n70143 & n70180;
  assign n70182 = n70178 & ~n70181;
  assign n70183 = ~n70131 & ~n70182;
  assign n70184 = ~n70137 & n70143;
  assign n70185 = n70149 & n70184;
  assign n70186 = n70156 & n70185;
  assign n70187 = ~n70170 & ~n70186;
  assign n70188 = n70137 & n70150;
  assign n70189 = n70156 & n70188;
  assign n70190 = n70187 & ~n70189;
  assign n70191 = ~n70162 & ~n70190;
  assign n70192 = n70137 & ~n70149;
  assign n70193 = n70143 & n70192;
  assign n70194 = ~n70162 & n70193;
  assign n70195 = n70156 & n70194;
  assign n70196 = ~n70143 & n70169;
  assign n70197 = ~n70143 & ~n70149;
  assign n70198 = ~n70156 & n70197;
  assign n70199 = ~n70196 & ~n70198;
  assign n70200 = ~n70162 & ~n70199;
  assign n70201 = ~n70195 & ~n70200;
  assign n70202 = ~n70131 & ~n70201;
  assign n70203 = ~n70191 & ~n70202;
  assign n70204 = ~n70183 & n70203;
  assign n70205 = n70137 & n70156;
  assign n70206 = n70162 & n70205;
  assign n70207 = n70197 & n70206;
  assign n70208 = n70137 & n70143;
  assign n70209 = n70166 & n70208;
  assign n70210 = ~n70156 & n70193;
  assign n70211 = ~n70137 & ~n70162;
  assign n70212 = n70143 & n70211;
  assign n70213 = ~n70143 & n70156;
  assign n70214 = n70137 & n70213;
  assign n70215 = ~n70212 & ~n70214;
  assign n70216 = ~n70210 & n70215;
  assign n70217 = ~n70188 & n70216;
  assign n70218 = n70150 & n70162;
  assign n70219 = ~n70156 & n70218;
  assign n70220 = n70156 & n70197;
  assign n70221 = n70137 & n70149;
  assign n70222 = ~n70220 & ~n70221;
  assign n70223 = n70162 & ~n70222;
  assign n70224 = ~n70219 & ~n70223;
  assign n70225 = n70217 & n70224;
  assign n70226 = n70131 & ~n70225;
  assign n70227 = ~n70209 & ~n70226;
  assign n70228 = ~n70207 & n70227;
  assign n70229 = n70204 & n70228;
  assign n70230 = pi2147 & n70229;
  assign n70231 = ~pi2147 & ~n70229;
  assign po2171 = n70230 | n70231;
  assign n70233 = n69596 & n69633;
  assign n70234 = ~n69609 & n70233;
  assign n70235 = ~n69932 & ~n70234;
  assign n70236 = n69609 & n69629;
  assign n70237 = n69615 & n70236;
  assign n70238 = ~n69609 & n69621;
  assign n70239 = ~n69956 & ~n70238;
  assign n70240 = ~n69596 & ~n70239;
  assign n70241 = ~n70237 & ~n70240;
  assign n70242 = n70235 & n70241;
  assign n70243 = n69602 & ~n70242;
  assign n70244 = ~n69631 & ~n69677;
  assign n70245 = ~n69609 & n69648;
  assign n70246 = n70244 & ~n70245;
  assign n70247 = n69596 & ~n70246;
  assign n70248 = n69633 & n69670;
  assign n70249 = ~n69657 & ~n70248;
  assign n70250 = ~n70247 & n70249;
  assign n70251 = ~n69640 & ~n69650;
  assign n70252 = ~n69596 & ~n70251;
  assign n70253 = n70250 & ~n70252;
  assign n70254 = ~n69602 & ~n70253;
  assign n70255 = ~n70243 & ~n70254;
  assign n70256 = ~n69609 & n69659;
  assign n70257 = n69609 & ~n69645;
  assign n70258 = ~n70256 & ~n70257;
  assign n70259 = ~n69596 & ~n70258;
  assign n70260 = ~n69631 & n69945;
  assign n70261 = n69918 & ~n70260;
  assign n70262 = ~n70259 & ~n70261;
  assign n70263 = n70255 & n70262;
  assign n70264 = ~pi2150 & ~n70263;
  assign n70265 = ~n70254 & n70262;
  assign n70266 = pi2150 & n70265;
  assign n70267 = ~n70243 & n70266;
  assign po2175 = n70264 | n70267;
  assign n70269 = n69998 & n70012;
  assign n70270 = ~n70051 & ~n70062;
  assign n70271 = n69979 & ~n70270;
  assign n70272 = ~n70269 & ~n70271;
  assign n70273 = ~n70059 & n70272;
  assign n70274 = ~n69979 & n70006;
  assign n70275 = ~n70044 & ~n70274;
  assign n70276 = ~n70009 & n70275;
  assign n70277 = n70273 & n70276;
  assign n70278 = n70020 & ~n70277;
  assign n70279 = n70004 & n70031;
  assign n70280 = n69998 & n70279;
  assign n70281 = ~n70029 & ~n70280;
  assign n70282 = n69992 & n70004;
  assign n70283 = n69979 & n70282;
  assign n70284 = n69998 & n70043;
  assign n70285 = ~n70283 & ~n70284;
  assign n70286 = n69985 & ~n70004;
  assign n70287 = n69991 & n69998;
  assign n70288 = ~n70286 & ~n70287;
  assign n70289 = ~n70048 & n70288;
  assign n70290 = ~n69979 & ~n70289;
  assign n70291 = ~n69998 & n70008;
  assign n70292 = ~n70025 & ~n70291;
  assign n70293 = ~n70290 & n70292;
  assign n70294 = n70285 & n70293;
  assign n70295 = n70281 & n70294;
  assign n70296 = ~n70020 & ~n70295;
  assign n70297 = ~n70278 & ~n70296;
  assign n70298 = pi2154 & ~n70297;
  assign n70299 = ~pi2154 & ~n70278;
  assign n70300 = ~n70296 & n70299;
  assign po2176 = n70298 | n70300;
  assign n70302 = pi6952 & pi9040;
  assign n70303 = pi6996 & ~pi9040;
  assign n70304 = ~n70302 & ~n70303;
  assign n70305 = pi2056 & n70304;
  assign n70306 = ~pi2056 & ~n70304;
  assign n70307 = ~n70305 & ~n70306;
  assign n70308 = pi6985 & pi9040;
  assign n70309 = pi6967 & ~pi9040;
  assign n70310 = ~n70308 & ~n70309;
  assign n70311 = ~pi2058 & ~n70310;
  assign n70312 = pi2058 & n70310;
  assign n70313 = ~n70311 & ~n70312;
  assign n70314 = pi7012 & ~pi9040;
  assign n70315 = pi6990 & pi9040;
  assign n70316 = ~n70314 & ~n70315;
  assign n70317 = pi2072 & n70316;
  assign n70318 = ~pi2072 & ~n70316;
  assign n70319 = ~n70317 & ~n70318;
  assign n70320 = n70313 & ~n70319;
  assign n70321 = pi6994 & pi9040;
  assign n70322 = pi6969 & ~pi9040;
  assign n70323 = ~n70321 & ~n70322;
  assign n70324 = ~pi2068 & ~n70323;
  assign n70325 = pi2068 & n70323;
  assign n70326 = ~n70324 & ~n70325;
  assign n70327 = pi6950 & ~pi9040;
  assign n70328 = pi6967 & pi9040;
  assign n70329 = ~n70327 & ~n70328;
  assign n70330 = ~pi2036 & n70329;
  assign n70331 = pi2036 & ~n70329;
  assign n70332 = ~n70330 & ~n70331;
  assign n70333 = n70326 & ~n70332;
  assign n70334 = n70320 & n70333;
  assign n70335 = n70313 & n70319;
  assign n70336 = n70332 & n70335;
  assign n70337 = ~n70313 & ~n70319;
  assign n70338 = n70332 & n70337;
  assign n70339 = ~n70336 & ~n70338;
  assign n70340 = n70326 & ~n70339;
  assign n70341 = ~n70334 & ~n70340;
  assign n70342 = ~n70307 & ~n70341;
  assign n70343 = ~n70326 & n70337;
  assign n70344 = ~n70313 & ~n70332;
  assign n70345 = n70319 & n70344;
  assign n70346 = ~n70343 & ~n70345;
  assign n70347 = pi6951 & pi9040;
  assign n70348 = pi6985 & ~pi9040;
  assign n70349 = ~n70347 & ~n70348;
  assign n70350 = pi2078 & n70349;
  assign n70351 = ~pi2078 & ~n70349;
  assign n70352 = ~n70350 & ~n70351;
  assign n70353 = ~n70307 & n70352;
  assign n70354 = ~n70346 & n70353;
  assign n70355 = ~n70342 & ~n70354;
  assign n70356 = n70326 & n70332;
  assign n70357 = ~n70313 & n70356;
  assign n70358 = ~n70334 & ~n70357;
  assign n70359 = ~n70352 & ~n70358;
  assign n70360 = ~n70326 & n70352;
  assign n70361 = n70313 & n70360;
  assign n70362 = n70320 & n70332;
  assign n70363 = ~n70332 & n70335;
  assign n70364 = ~n70362 & ~n70363;
  assign n70365 = ~n70332 & n70337;
  assign n70366 = n70326 & n70365;
  assign n70367 = n70364 & ~n70366;
  assign n70368 = n70352 & ~n70367;
  assign n70369 = ~n70361 & ~n70368;
  assign n70370 = ~n70313 & n70319;
  assign n70371 = n70332 & n70370;
  assign n70372 = n70326 & n70371;
  assign n70373 = n70369 & ~n70372;
  assign n70374 = ~n70346 & ~n70352;
  assign n70375 = ~n70326 & n70336;
  assign n70376 = ~n70374 & ~n70375;
  assign n70377 = n70373 & n70376;
  assign n70378 = n70307 & ~n70377;
  assign n70379 = ~n70359 & ~n70378;
  assign n70380 = ~n70307 & ~n70352;
  assign n70381 = n70320 & ~n70326;
  assign n70382 = ~n70371 & ~n70381;
  assign n70383 = n70313 & ~n70332;
  assign n70384 = n70382 & ~n70383;
  assign n70385 = n70380 & ~n70384;
  assign n70386 = n70379 & ~n70385;
  assign n70387 = n70355 & n70386;
  assign n70388 = ~pi2144 & ~n70387;
  assign n70389 = pi2144 & n70355;
  assign n70390 = n70379 & n70389;
  assign n70391 = ~n70385 & n70390;
  assign po2177 = n70388 | n70391;
  assign n70393 = ~n70137 & ~n70143;
  assign n70394 = ~n70181 & ~n70393;
  assign n70395 = ~n70213 & n70394;
  assign n70396 = n70162 & ~n70395;
  assign n70397 = n70156 & ~n70162;
  assign n70398 = n70143 & n70397;
  assign n70399 = n70137 & ~n70143;
  assign n70400 = ~n70156 & ~n70162;
  assign n70401 = n70399 & n70400;
  assign n70402 = ~n70137 & n70149;
  assign n70403 = n70156 & n70402;
  assign n70404 = ~n70156 & n70173;
  assign n70405 = ~n70403 & ~n70404;
  assign n70406 = ~n70401 & n70405;
  assign n70407 = ~n70398 & n70406;
  assign n70408 = ~n70396 & n70407;
  assign n70409 = n70131 & ~n70408;
  assign n70410 = ~n70137 & n70150;
  assign n70411 = ~n70156 & n70410;
  assign n70412 = ~n70137 & n70197;
  assign n70413 = n70156 & n70412;
  assign n70414 = ~n70411 & ~n70413;
  assign n70415 = n70162 & ~n70414;
  assign n70416 = ~n70409 & ~n70415;
  assign n70417 = n70156 & n70173;
  assign n70418 = ~n70185 & ~n70193;
  assign n70419 = n70162 & ~n70418;
  assign n70420 = ~n70417 & ~n70419;
  assign n70421 = ~n70189 & n70420;
  assign n70422 = ~n70131 & ~n70421;
  assign n70423 = ~n70167 & ~n70197;
  assign n70424 = n70137 & ~n70423;
  assign n70425 = ~n70198 & ~n70424;
  assign n70426 = ~n70162 & ~n70425;
  assign n70427 = ~n70131 & n70426;
  assign n70428 = ~n70422 & ~n70427;
  assign n70429 = n70416 & n70428;
  assign n70430 = pi2146 & ~n70429;
  assign n70431 = ~pi2146 & n70416;
  assign n70432 = n70428 & n70431;
  assign po2178 = n70430 | n70432;
  assign n70434 = ~n70101 & ~n70106;
  assign n70435 = ~n69802 & n69835;
  assign n70436 = ~n70094 & ~n70435;
  assign n70437 = ~n70077 & n70436;
  assign n70438 = ~n69829 & ~n70437;
  assign n70439 = ~n69863 & ~n69874;
  assign n70440 = ~n70113 & n70439;
  assign n70441 = ~n69829 & ~n70440;
  assign n70442 = ~n69889 & n70436;
  assign n70443 = n69829 & n69850;
  assign n70444 = n70442 & ~n70443;
  assign n70445 = ~n70441 & n70444;
  assign n70446 = n69796 & ~n70445;
  assign n70447 = n69814 & n69861;
  assign n70448 = ~n70111 & ~n70447;
  assign n70449 = ~n69829 & n69833;
  assign n70450 = n69802 & n70449;
  assign n70451 = ~n69829 & n69841;
  assign n70452 = ~n70450 & ~n70451;
  assign n70453 = n69802 & n69843;
  assign n70454 = n69814 & n69856;
  assign n70455 = ~n69874 & ~n70454;
  assign n70456 = n69829 & ~n70455;
  assign n70457 = ~n70453 & ~n70456;
  assign n70458 = n70452 & n70457;
  assign n70459 = n70448 & n70458;
  assign n70460 = ~n70077 & n70459;
  assign n70461 = ~n69796 & ~n70460;
  assign n70462 = ~n70446 & ~n70461;
  assign n70463 = ~n70438 & n70462;
  assign n70464 = n70434 & n70463;
  assign n70465 = pi2171 & ~n70464;
  assign n70466 = ~pi2171 & n70464;
  assign po2179 = n70465 | n70466;
  assign n70468 = n70156 & n70424;
  assign n70469 = ~n70192 & ~n70410;
  assign n70470 = ~n70162 & ~n70469;
  assign n70471 = ~n70468 & ~n70470;
  assign n70472 = ~n70137 & n70156;
  assign n70473 = ~n70149 & n70472;
  assign n70474 = ~n70221 & ~n70473;
  assign n70475 = ~n70412 & n70474;
  assign n70476 = n70162 & ~n70475;
  assign n70477 = n70471 & ~n70476;
  assign n70478 = ~n70156 & n70185;
  assign n70479 = n70477 & ~n70478;
  assign n70480 = ~n70131 & ~n70479;
  assign n70481 = n70166 & ~n70469;
  assign n70482 = ~n70188 & ~n70193;
  assign n70483 = ~n70185 & ~n70412;
  assign n70484 = n70482 & n70483;
  assign n70485 = n70156 & ~n70484;
  assign n70486 = ~n70481 & ~n70485;
  assign n70487 = ~n70404 & n70486;
  assign n70488 = n70131 & ~n70487;
  assign n70489 = ~n70480 & ~n70488;
  assign n70490 = n70156 & n70410;
  assign n70491 = ~n70478 & ~n70490;
  assign n70492 = ~n70162 & ~n70491;
  assign n70493 = n70489 & ~n70492;
  assign n70494 = pi2149 & ~n70493;
  assign n70495 = ~pi2149 & ~n70492;
  assign n70496 = ~n70488 & n70495;
  assign n70497 = ~n70480 & n70496;
  assign po2183 = n70494 | n70497;
  assign n70499 = n70326 & ~n70352;
  assign n70500 = ~n70336 & ~n70337;
  assign n70501 = n70499 & ~n70500;
  assign n70502 = n70332 & ~n70352;
  assign n70503 = n70337 & n70502;
  assign n70504 = ~n70501 & ~n70503;
  assign n70505 = n70307 & ~n70504;
  assign n70506 = ~n70326 & n70363;
  assign n70507 = ~n70326 & ~n70332;
  assign n70508 = ~n70383 & ~n70507;
  assign n70509 = n70352 & ~n70508;
  assign n70510 = ~n70326 & n70332;
  assign n70511 = ~n70319 & n70510;
  assign n70512 = n70313 & n70511;
  assign n70513 = ~n70509 & ~n70512;
  assign n70514 = ~n70506 & n70513;
  assign n70515 = n70307 & ~n70514;
  assign n70516 = ~n70505 & ~n70515;
  assign n70517 = n70319 & n70333;
  assign n70518 = ~n70313 & n70517;
  assign n70519 = ~n70326 & n70371;
  assign n70520 = ~n70518 & ~n70519;
  assign n70521 = ~n70352 & ~n70520;
  assign n70522 = n70326 & n70338;
  assign n70523 = ~n70326 & n70383;
  assign n70524 = ~n70522 & ~n70523;
  assign n70525 = n70352 & ~n70524;
  assign n70526 = ~n70320 & ~n70383;
  assign n70527 = n70326 & ~n70526;
  assign n70528 = ~n70371 & ~n70527;
  assign n70529 = ~n70352 & ~n70528;
  assign n70530 = n70319 & ~n70326;
  assign n70531 = n70502 & n70530;
  assign n70532 = ~n70319 & ~n70332;
  assign n70533 = ~n70371 & ~n70532;
  assign n70534 = ~n70326 & ~n70533;
  assign n70535 = n70326 & n70352;
  assign n70536 = n70335 & n70535;
  assign n70537 = n70332 & n70536;
  assign n70538 = ~n70534 & ~n70537;
  assign n70539 = ~n70531 & n70538;
  assign n70540 = ~n70529 & n70539;
  assign n70541 = ~n70518 & n70540;
  assign n70542 = ~n70307 & ~n70541;
  assign n70543 = ~n70525 & ~n70542;
  assign n70544 = ~n70521 & n70543;
  assign n70545 = n70516 & n70544;
  assign n70546 = pi2155 & n70545;
  assign n70547 = ~pi2155 & ~n70545;
  assign po2184 = n70546 | n70547;
  assign n70549 = pi6993 & pi9040;
  assign n70550 = pi6992 & ~pi9040;
  assign n70551 = ~n70549 & ~n70550;
  assign n70552 = pi2043 & n70551;
  assign n70553 = ~pi2043 & ~n70551;
  assign n70554 = ~n70552 & ~n70553;
  assign n70555 = pi6955 & ~pi9040;
  assign n70556 = pi6975 & pi9040;
  assign n70557 = ~n70555 & ~n70556;
  assign n70558 = pi2065 & n70557;
  assign n70559 = ~pi2065 & ~n70557;
  assign n70560 = ~n70558 & ~n70559;
  assign n70561 = pi6966 & ~pi9040;
  assign n70562 = pi6955 & pi9040;
  assign n70563 = ~n70561 & ~n70562;
  assign n70564 = pi2070 & n70563;
  assign n70565 = ~pi2070 & ~n70563;
  assign n70566 = ~n70564 & ~n70565;
  assign n70567 = pi6953 & ~pi9040;
  assign n70568 = pi7003 & pi9040;
  assign n70569 = ~n70567 & ~n70568;
  assign n70570 = pi2079 & n70569;
  assign n70571 = ~pi2079 & ~n70569;
  assign n70572 = ~n70570 & ~n70571;
  assign n70573 = n70566 & ~n70572;
  assign n70574 = n70560 & n70573;
  assign n70575 = pi6988 & pi9040;
  assign n70576 = pi6961 & ~pi9040;
  assign n70577 = ~n70575 & ~n70576;
  assign n70578 = pi2069 & n70577;
  assign n70579 = ~pi2069 & ~n70577;
  assign n70580 = ~n70578 & ~n70579;
  assign n70581 = ~n70560 & n70566;
  assign n70582 = n70580 & n70581;
  assign n70583 = n70572 & n70582;
  assign n70584 = ~n70574 & ~n70583;
  assign n70585 = pi6959 & ~pi9040;
  assign n70586 = pi6946 & pi9040;
  assign n70587 = ~n70585 & ~n70586;
  assign n70588 = ~pi2064 & n70587;
  assign n70589 = pi2064 & ~n70587;
  assign n70590 = ~n70588 & ~n70589;
  assign n70591 = n70573 & ~n70580;
  assign n70592 = n70560 & n70580;
  assign n70593 = ~n70566 & n70592;
  assign n70594 = ~n70591 & ~n70593;
  assign n70595 = n70590 & ~n70594;
  assign n70596 = n70584 & ~n70595;
  assign n70597 = n70566 & n70592;
  assign n70598 = ~n70566 & ~n70580;
  assign n70599 = ~n70560 & ~n70566;
  assign n70600 = ~n70572 & n70599;
  assign n70601 = ~n70560 & ~n70580;
  assign n70602 = n70572 & n70601;
  assign n70603 = ~n70600 & ~n70602;
  assign n70604 = ~n70598 & n70603;
  assign n70605 = ~n70597 & n70604;
  assign n70606 = ~n70590 & ~n70605;
  assign n70607 = n70596 & ~n70606;
  assign n70608 = n70554 & ~n70607;
  assign n70609 = n70560 & ~n70580;
  assign n70610 = ~n70566 & n70609;
  assign n70611 = ~n70572 & n70610;
  assign n70612 = ~n70566 & n70601;
  assign n70613 = n70572 & n70612;
  assign n70614 = ~n70583 & ~n70613;
  assign n70615 = ~n70611 & n70614;
  assign n70616 = ~n70590 & ~n70615;
  assign n70617 = ~n70608 & ~n70616;
  assign n70618 = n70574 & n70580;
  assign n70619 = ~n70566 & n70580;
  assign n70620 = n70590 & n70619;
  assign n70621 = n70572 & n70620;
  assign n70622 = ~n70572 & ~n70590;
  assign n70623 = n70566 & n70622;
  assign n70624 = ~n70560 & n70623;
  assign n70625 = n70566 & n70609;
  assign n70626 = n70572 & n70625;
  assign n70627 = ~n70624 & ~n70626;
  assign n70628 = n70566 & ~n70580;
  assign n70629 = n70572 & n70628;
  assign n70630 = ~n70560 & n70580;
  assign n70631 = ~n70566 & n70630;
  assign n70632 = ~n70629 & ~n70631;
  assign n70633 = n70590 & ~n70632;
  assign n70634 = n70590 & n70598;
  assign n70635 = ~n70572 & n70634;
  assign n70636 = ~n70633 & ~n70635;
  assign n70637 = n70627 & n70636;
  assign n70638 = ~n70554 & ~n70637;
  assign n70639 = ~n70621 & ~n70638;
  assign n70640 = ~n70618 & n70639;
  assign n70641 = n70617 & n70640;
  assign n70642 = ~pi2156 & ~n70641;
  assign n70643 = ~n70608 & ~n70618;
  assign n70644 = ~n70616 & n70643;
  assign n70645 = n70639 & n70644;
  assign n70646 = pi2156 & n70645;
  assign po2185 = n70642 | n70646;
  assign n70648 = ~n70572 & n70590;
  assign n70649 = n70580 & n70648;
  assign n70650 = n70566 & n70601;
  assign n70651 = n70572 & n70650;
  assign n70652 = n70572 & n70610;
  assign n70653 = ~n70651 & ~n70652;
  assign n70654 = ~n70566 & ~n70572;
  assign n70655 = ~n70560 & n70654;
  assign n70656 = ~n70580 & n70655;
  assign n70657 = ~n70593 & ~n70656;
  assign n70658 = ~n70590 & ~n70657;
  assign n70659 = n70653 & ~n70658;
  assign n70660 = ~n70649 & n70659;
  assign n70661 = n70554 & ~n70660;
  assign n70662 = n70572 & n70631;
  assign n70663 = n70590 & n70662;
  assign n70664 = n70622 & n70631;
  assign n70665 = ~n70591 & ~n70664;
  assign n70666 = ~n70593 & ~n70625;
  assign n70667 = ~n70572 & n70609;
  assign n70668 = n70666 & ~n70667;
  assign n70669 = n70590 & ~n70668;
  assign n70670 = ~n70590 & n70597;
  assign n70671 = n70614 & ~n70670;
  assign n70672 = ~n70669 & n70671;
  assign n70673 = n70665 & n70672;
  assign n70674 = ~n70554 & ~n70673;
  assign n70675 = ~n70663 & ~n70674;
  assign n70676 = ~n70661 & n70675;
  assign n70677 = n70622 & n70625;
  assign n70678 = n70581 & ~n70590;
  assign n70679 = n70572 & n70678;
  assign n70680 = ~n70677 & ~n70679;
  assign n70681 = ~n70590 & n70652;
  assign n70682 = n70680 & ~n70681;
  assign n70683 = n70676 & n70682;
  assign n70684 = ~pi2148 & ~n70683;
  assign n70685 = n70675 & n70682;
  assign n70686 = pi2148 & n70685;
  assign n70687 = ~n70661 & n70686;
  assign po2186 = n70684 | n70687;
  assign n70689 = ~n70572 & n70650;
  assign n70690 = n70572 & n70581;
  assign n70691 = ~n70572 & n70631;
  assign n70692 = ~n70690 & ~n70691;
  assign n70693 = ~n70610 & ~n70618;
  assign n70694 = n70692 & n70693;
  assign n70695 = n70590 & ~n70694;
  assign n70696 = n70572 & n70592;
  assign n70697 = ~n70591 & ~n70696;
  assign n70698 = ~n70612 & n70697;
  assign n70699 = ~n70590 & ~n70698;
  assign n70700 = n70572 & n70593;
  assign n70701 = ~n70699 & ~n70700;
  assign n70702 = ~n70695 & n70701;
  assign n70703 = ~n70689 & n70702;
  assign n70704 = ~n70554 & ~n70703;
  assign n70705 = n70572 & n70590;
  assign n70706 = n70597 & n70705;
  assign n70707 = n70590 & n70612;
  assign n70708 = n70590 & n70625;
  assign n70709 = ~n70707 & ~n70708;
  assign n70710 = ~n70572 & ~n70709;
  assign n70711 = ~n70706 & ~n70710;
  assign n70712 = ~n70572 & n70582;
  assign n70713 = ~n70662 & ~n70712;
  assign n70714 = n70572 & n70609;
  assign n70715 = ~n70572 & n70592;
  assign n70716 = ~n70714 & ~n70715;
  assign n70717 = ~n70582 & n70716;
  assign n70718 = ~n70610 & n70717;
  assign n70719 = ~n70590 & ~n70718;
  assign n70720 = ~n70572 & n70593;
  assign n70721 = ~n70719 & ~n70720;
  assign n70722 = n70713 & n70721;
  assign n70723 = n70711 & n70722;
  assign n70724 = n70554 & ~n70723;
  assign n70725 = n70590 & ~n70653;
  assign n70726 = ~n70724 & ~n70725;
  assign n70727 = ~n70613 & ~n70712;
  assign n70728 = ~n70590 & ~n70727;
  assign n70729 = n70726 & ~n70728;
  assign n70730 = ~n70704 & n70729;
  assign n70731 = pi2165 & ~n70730;
  assign n70732 = ~pi2165 & n70730;
  assign po2187 = n70731 | n70732;
  assign n70734 = ~n70156 & n70188;
  assign n70735 = ~n70404 & ~n70734;
  assign n70736 = ~n70162 & ~n70735;
  assign n70737 = n70185 & n70397;
  assign n70738 = ~n70736 & ~n70737;
  assign n70739 = ~n70209 & n70738;
  assign n70740 = ~n70137 & n70162;
  assign n70741 = ~n70149 & n70740;
  assign n70742 = ~n70143 & n70741;
  assign n70743 = ~n70156 & n70742;
  assign n70744 = n70162 & n70410;
  assign n70745 = ~n70181 & ~n70207;
  assign n70746 = ~n70175 & n70745;
  assign n70747 = ~n70744 & n70746;
  assign n70748 = n70131 & ~n70747;
  assign n70749 = n70156 & n70193;
  assign n70750 = ~n70188 & ~n70749;
  assign n70751 = ~n70412 & n70750;
  assign n70752 = ~n70162 & ~n70751;
  assign n70753 = n70131 & n70752;
  assign n70754 = n70156 & n70218;
  assign n70755 = ~n70742 & ~n70754;
  assign n70756 = ~n70403 & n70755;
  assign n70757 = ~n70149 & n70179;
  assign n70758 = n70156 & n70167;
  assign n70759 = ~n70184 & ~n70758;
  assign n70760 = ~n70162 & ~n70759;
  assign n70761 = ~n70757 & ~n70760;
  assign n70762 = n70756 & n70761;
  assign n70763 = ~n70131 & ~n70762;
  assign n70764 = ~n70753 & ~n70763;
  assign n70765 = ~n70748 & n70764;
  assign n70766 = ~n70743 & n70765;
  assign n70767 = n70739 & n70766;
  assign n70768 = pi2151 & ~n70767;
  assign n70769 = ~pi2151 & n70739;
  assign n70770 = n70766 & n70769;
  assign po2188 = n70768 | n70770;
  assign n70772 = ~n69849 & ~n69857;
  assign n70773 = n69796 & ~n70772;
  assign n70774 = ~n69862 & ~n70083;
  assign n70775 = ~n69822 & n70774;
  assign n70776 = ~n69829 & ~n70775;
  assign n70777 = n69796 & n70776;
  assign n70778 = ~n70773 & ~n70777;
  assign n70779 = n69848 & n70086;
  assign n70780 = ~n70088 & ~n70779;
  assign n70781 = ~n69865 & ~n70114;
  assign n70782 = n69829 & ~n70781;
  assign n70783 = n69796 & n70782;
  assign n70784 = n70780 & ~n70783;
  assign n70785 = n69802 & n69848;
  assign n70786 = n69802 & n69840;
  assign n70787 = ~n70079 & ~n70786;
  assign n70788 = n69829 & ~n70787;
  assign n70789 = ~n69863 & ~n70094;
  assign n70790 = n69802 & n69847;
  assign n70791 = ~n69887 & ~n70790;
  assign n70792 = ~n69829 & ~n70791;
  assign n70793 = n70789 & ~n70792;
  assign n70794 = ~n70788 & n70793;
  assign n70795 = ~n70785 & n70794;
  assign n70796 = ~n69796 & ~n70795;
  assign n70797 = ~n70111 & n70436;
  assign n70798 = n69829 & ~n70797;
  assign n70799 = ~n70796 & ~n70798;
  assign n70800 = n70784 & n70799;
  assign n70801 = n70778 & n70800;
  assign n70802 = ~pi2161 & ~n70801;
  assign n70803 = pi2161 & n70784;
  assign n70804 = n70778 & n70803;
  assign n70805 = n70799 & n70804;
  assign po2189 = n70802 | n70805;
  assign n70807 = pi6957 & pi9040;
  assign n70808 = pi6968 & ~pi9040;
  assign n70809 = ~n70807 & ~n70808;
  assign n70810 = ~pi2072 & n70809;
  assign n70811 = pi2072 & ~n70809;
  assign n70812 = ~n70810 & ~n70811;
  assign n70813 = pi6974 & ~pi9040;
  assign n70814 = pi6972 & pi9040;
  assign n70815 = ~n70813 & ~n70814;
  assign n70816 = ~pi2067 & ~n70815;
  assign n70817 = pi2067 & n70815;
  assign n70818 = ~n70816 & ~n70817;
  assign n70819 = pi6965 & pi9040;
  assign n70820 = pi7082 & ~pi9040;
  assign n70821 = ~n70819 & ~n70820;
  assign n70822 = ~pi2056 & n70821;
  assign n70823 = pi2056 & ~n70821;
  assign n70824 = ~n70822 & ~n70823;
  assign n70825 = ~n70818 & ~n70824;
  assign n70826 = n70812 & n70825;
  assign n70827 = n70818 & ~n70824;
  assign n70828 = ~n70812 & n70827;
  assign n70829 = ~n70826 & ~n70828;
  assign n70830 = pi6969 & pi9040;
  assign n70831 = pi6981 & ~pi9040;
  assign n70832 = ~n70830 & ~n70831;
  assign n70833 = pi2054 & n70832;
  assign n70834 = ~pi2054 & ~n70832;
  assign n70835 = ~n70833 & ~n70834;
  assign n70836 = ~n70812 & ~n70835;
  assign n70837 = n70818 & n70836;
  assign n70838 = n70829 & ~n70837;
  assign n70839 = pi6947 & pi9040;
  assign n70840 = pi6954 & ~pi9040;
  assign n70841 = ~n70839 & ~n70840;
  assign n70842 = ~pi2053 & n70841;
  assign n70843 = pi2053 & ~n70841;
  assign n70844 = ~n70842 & ~n70843;
  assign n70845 = pi6986 & pi9040;
  assign n70846 = pi6965 & ~pi9040;
  assign n70847 = ~n70845 & ~n70846;
  assign n70848 = ~pi2073 & ~n70847;
  assign n70849 = pi2073 & n70847;
  assign n70850 = ~n70848 & ~n70849;
  assign n70851 = n70844 & n70850;
  assign n70852 = ~n70838 & n70851;
  assign n70853 = ~n70818 & n70824;
  assign n70854 = ~n70812 & n70853;
  assign n70855 = n70835 & n70850;
  assign n70856 = n70854 & n70855;
  assign n70857 = ~n70812 & n70825;
  assign n70858 = ~n70844 & n70857;
  assign n70859 = n70818 & n70824;
  assign n70860 = n70835 & n70859;
  assign n70861 = n70812 & n70818;
  assign n70862 = ~n70860 & ~n70861;
  assign n70863 = ~n70844 & ~n70862;
  assign n70864 = ~n70858 & ~n70863;
  assign n70865 = n70850 & ~n70864;
  assign n70866 = ~n70856 & ~n70865;
  assign n70867 = n70812 & ~n70835;
  assign n70868 = ~n70818 & n70867;
  assign n70869 = n70824 & n70868;
  assign n70870 = n70812 & n70835;
  assign n70871 = n70818 & n70870;
  assign n70872 = ~n70869 & ~n70871;
  assign n70873 = ~n70844 & ~n70872;
  assign n70874 = n70866 & ~n70873;
  assign n70875 = n70835 & n70844;
  assign n70876 = n70859 & n70875;
  assign n70877 = ~n70812 & n70876;
  assign n70878 = n70812 & n70859;
  assign n70879 = ~n70835 & n70844;
  assign n70880 = n70878 & n70879;
  assign n70881 = ~n70827 & ~n70853;
  assign n70882 = n70836 & ~n70881;
  assign n70883 = n70826 & ~n70835;
  assign n70884 = ~n70882 & ~n70883;
  assign n70885 = n70870 & ~n70881;
  assign n70886 = n70835 & n70857;
  assign n70887 = ~n70885 & ~n70886;
  assign n70888 = n70884 & n70887;
  assign n70889 = ~n70880 & n70888;
  assign n70890 = ~n70877 & n70889;
  assign n70891 = ~n70835 & ~n70844;
  assign n70892 = ~n70812 & n70891;
  assign n70893 = n70824 & n70892;
  assign n70894 = n70890 & ~n70893;
  assign n70895 = ~n70850 & ~n70894;
  assign n70896 = n70874 & ~n70895;
  assign n70897 = ~n70852 & n70896;
  assign n70898 = ~pi2195 & ~n70897;
  assign n70899 = pi2195 & n70874;
  assign n70900 = ~n70852 & n70899;
  assign n70901 = ~n70895 & n70900;
  assign po2190 = n70898 | n70901;
  assign n70903 = ~n69998 & n70031;
  assign n70904 = ~n70291 & ~n70903;
  assign n70905 = n69979 & n70904;
  assign n70906 = ~n69992 & ~n70011;
  assign n70907 = ~n70004 & ~n70906;
  assign n70908 = n69998 & n70053;
  assign n70909 = ~n69991 & n70023;
  assign n70910 = n69998 & n70011;
  assign n70911 = ~n70909 & ~n70910;
  assign n70912 = ~n70908 & n70911;
  assign n70913 = ~n70907 & n70912;
  assign n70914 = ~n69979 & n70913;
  assign n70915 = ~n70905 & ~n70914;
  assign n70916 = n69998 & n70907;
  assign n70917 = ~n70280 & ~n70916;
  assign n70918 = ~n70915 & n70917;
  assign n70919 = n70020 & ~n70918;
  assign n70920 = n69979 & ~n70906;
  assign n70921 = ~n69998 & n70920;
  assign n70922 = ~n70007 & ~n70041;
  assign n70923 = n69998 & ~n70922;
  assign n70924 = n69979 & n70923;
  assign n70925 = n70004 & n70920;
  assign n70926 = ~n70924 & ~n70925;
  assign n70927 = ~n70921 & n70926;
  assign n70928 = ~n70020 & ~n70927;
  assign n70929 = ~n70919 & ~n70928;
  assign n70930 = n69979 & n70029;
  assign n70931 = ~n69979 & ~n70917;
  assign n70932 = ~n70930 & ~n70931;
  assign n70933 = ~n69979 & ~n70904;
  assign n70934 = ~n70029 & ~n70933;
  assign n70935 = ~n70020 & ~n70934;
  assign n70936 = n70932 & ~n70935;
  assign n70937 = n70929 & n70936;
  assign n70938 = pi2201 & ~n70937;
  assign n70939 = ~pi2201 & n70936;
  assign n70940 = ~n70928 & n70939;
  assign n70941 = ~n70919 & n70940;
  assign po2191 = n70938 | n70941;
  assign n70943 = ~n70812 & n70859;
  assign n70944 = ~n70844 & n70943;
  assign n70945 = ~n70835 & n70944;
  assign n70946 = n70825 & n70891;
  assign n70947 = n70812 & n70946;
  assign n70948 = ~n70945 & ~n70947;
  assign n70949 = ~n70880 & ~n70883;
  assign n70950 = ~n70812 & ~n70824;
  assign n70951 = n70835 & n70950;
  assign n70952 = ~n70860 & ~n70951;
  assign n70953 = ~n70844 & ~n70952;
  assign n70954 = n70844 & ~n70867;
  assign n70955 = ~n70881 & n70954;
  assign n70956 = ~n70859 & n70891;
  assign n70957 = n70812 & n70956;
  assign n70958 = ~n70955 & ~n70957;
  assign n70959 = ~n70953 & n70958;
  assign n70960 = n70949 & n70959;
  assign n70961 = n70850 & ~n70960;
  assign n70962 = n70948 & ~n70961;
  assign n70963 = n70828 & n70844;
  assign n70964 = n70835 & n70963;
  assign n70965 = n70844 & ~n70850;
  assign n70966 = ~n70857 & ~n70860;
  assign n70967 = n70867 & ~n70881;
  assign n70968 = n70966 & ~n70967;
  assign n70969 = n70965 & ~n70968;
  assign n70970 = n70826 & n70835;
  assign n70971 = ~n70824 & n70835;
  assign n70972 = n70812 & n70971;
  assign n70973 = n70835 & n70853;
  assign n70974 = ~n70972 & ~n70973;
  assign n70975 = ~n70835 & n70859;
  assign n70976 = ~n70854 & ~n70975;
  assign n70977 = n70974 & n70976;
  assign n70978 = ~n70844 & ~n70977;
  assign n70979 = ~n70970 & ~n70978;
  assign n70980 = ~n70850 & ~n70979;
  assign n70981 = ~n70969 & ~n70980;
  assign n70982 = ~n70964 & n70981;
  assign n70983 = n70962 & n70982;
  assign n70984 = pi2186 & ~n70983;
  assign n70985 = ~pi2186 & n70962;
  assign n70986 = n70982 & n70985;
  assign po2192 = n70984 | n70986;
  assign n70988 = ~n70656 & ~n70712;
  assign n70989 = ~n70700 & n70988;
  assign n70990 = n70590 & ~n70989;
  assign n70991 = ~n70662 & ~n70708;
  assign n70992 = ~n70650 & ~n70715;
  assign n70993 = ~n70590 & ~n70992;
  assign n70994 = ~n70618 & ~n70993;
  assign n70995 = n70991 & n70994;
  assign n70996 = n70554 & ~n70995;
  assign n70997 = n70560 & ~n70566;
  assign n70998 = ~n70598 & ~n70997;
  assign n70999 = n70572 & ~n70998;
  assign n71000 = ~n70582 & ~n70667;
  assign n71001 = ~n70590 & ~n71000;
  assign n71002 = n70560 & n70572;
  assign n71003 = ~n70593 & ~n71002;
  assign n71004 = ~n70601 & n71003;
  assign n71005 = n70590 & ~n71004;
  assign n71006 = ~n71001 & ~n71005;
  assign n71007 = ~n70999 & n71006;
  assign n71008 = ~n70554 & ~n71007;
  assign n71009 = ~n70996 & ~n71008;
  assign n71010 = ~n70664 & ~n70681;
  assign n71011 = n71009 & n71010;
  assign n71012 = ~n70990 & n71011;
  assign n71013 = ~pi2179 & ~n71012;
  assign n71014 = pi2179 & n71010;
  assign n71015 = ~n70990 & n71014;
  assign n71016 = n71009 & n71015;
  assign po2193 = n71013 | n71016;
  assign n71018 = ~n70973 & ~n70975;
  assign n71019 = ~n70844 & ~n71018;
  assign n71020 = ~n70947 & ~n71019;
  assign n71021 = n70850 & ~n71020;
  assign n71022 = n70835 & n70878;
  assign n71023 = ~n70818 & n70836;
  assign n71024 = n70812 & ~n70824;
  assign n71025 = ~n70827 & ~n71024;
  assign n71026 = n70835 & ~n71025;
  assign n71027 = ~n71023 & ~n71026;
  assign n71028 = ~n70844 & ~n71027;
  assign n71029 = ~n71022 & ~n71028;
  assign n71030 = ~n70835 & ~n71025;
  assign n71031 = ~n70943 & ~n71030;
  assign n71032 = n70844 & ~n71031;
  assign n71033 = ~n70967 & ~n71032;
  assign n71034 = n71029 & n71033;
  assign n71035 = ~n70850 & ~n71034;
  assign n71036 = ~n70812 & n70835;
  assign n71037 = ~n70827 & n71036;
  assign n71038 = n70850 & n71037;
  assign n71039 = n70827 & n70870;
  assign n71040 = ~n70844 & n71039;
  assign n71041 = ~n70812 & ~n70818;
  assign n71042 = n70875 & n71041;
  assign n71043 = ~n71040 & ~n71042;
  assign n71044 = ~n71038 & n71043;
  assign n71045 = ~n70854 & ~n70971;
  assign n71046 = n70851 & ~n71045;
  assign n71047 = n71044 & ~n71046;
  assign n71048 = ~n71035 & n71047;
  assign n71049 = ~n71021 & n71048;
  assign n71050 = pi2205 & ~n71049;
  assign n71051 = ~pi2205 & n71049;
  assign po2194 = n71050 | n71051;
  assign n71053 = ~n69724 & ~n69730;
  assign n71054 = ~n69697 & ~n71053;
  assign n71055 = ~n69784 & ~n71054;
  assign n71056 = ~n69703 & n69709;
  assign n71057 = n69697 & n71056;
  assign n71058 = n69723 & n71057;
  assign n71059 = n69723 & n69737;
  assign n71060 = ~n71056 & ~n71059;
  assign n71061 = n69703 & ~n69723;
  assign n71062 = ~n69709 & n71061;
  assign n71063 = n71060 & ~n71062;
  assign n71064 = n69697 & ~n71063;
  assign n71065 = ~n69733 & ~n71064;
  assign n71066 = ~n69761 & ~n71065;
  assign n71067 = ~n69697 & n69716;
  assign n71068 = n69723 & n71067;
  assign n71069 = ~n69697 & n69703;
  assign n71070 = n69725 & n71069;
  assign n71071 = ~n71068 & ~n71070;
  assign n71072 = ~n69761 & ~n71071;
  assign n71073 = ~n71066 & ~n71072;
  assign n71074 = ~n71058 & n71073;
  assign n71075 = ~n69709 & n69726;
  assign n71076 = ~n69749 & ~n69767;
  assign n71077 = ~n69777 & n71076;
  assign n71078 = ~n69697 & ~n71077;
  assign n71079 = ~n69723 & n69729;
  assign n71080 = ~n69752 & ~n71079;
  assign n71081 = n69697 & ~n71080;
  assign n71082 = ~n71078 & ~n71081;
  assign n71083 = ~n71075 & n71082;
  assign n71084 = ~n69739 & ~n69778;
  assign n71085 = n71083 & n71084;
  assign n71086 = n69761 & ~n71085;
  assign n71087 = n71074 & ~n71086;
  assign n71088 = n71055 & n71087;
  assign n71089 = ~pi2200 & ~n71088;
  assign n71090 = pi2200 & n71074;
  assign n71091 = n71055 & n71090;
  assign n71092 = ~n71086 & n71091;
  assign po2195 = n71089 | n71092;
  assign n71094 = ~n69723 & n69752;
  assign n71095 = ~n69715 & n69723;
  assign n71096 = ~n69703 & n71095;
  assign n71097 = ~n69749 & ~n71096;
  assign n71098 = n69697 & ~n71097;
  assign n71099 = ~n71094 & ~n71098;
  assign n71100 = ~n69697 & ~n69723;
  assign n71101 = ~n69715 & n71100;
  assign n71102 = ~n69709 & n71101;
  assign n71103 = n69731 & n69764;
  assign n71104 = ~n71102 & ~n71103;
  assign n71105 = ~n71070 & n71104;
  assign n71106 = ~n69727 & ~n69739;
  assign n71107 = n69715 & n69769;
  assign n71108 = n71106 & ~n71107;
  assign n71109 = n71105 & n71108;
  assign n71110 = n71099 & n71109;
  assign n71111 = ~n69761 & ~n71110;
  assign n71112 = ~n69703 & n69725;
  assign n71113 = ~n69749 & ~n71112;
  assign n71114 = n69723 & ~n71113;
  assign n71115 = ~n69777 & ~n71075;
  assign n71116 = n69703 & ~n69715;
  assign n71117 = n69723 & n71116;
  assign n71118 = n71115 & ~n71117;
  assign n71119 = n69697 & ~n71118;
  assign n71120 = ~n69723 & n69737;
  assign n71121 = ~n69703 & n69723;
  assign n71122 = ~n69715 & n71121;
  assign n71123 = ~n69709 & n71122;
  assign n71124 = ~n71120 & ~n71123;
  assign n71125 = ~n69697 & ~n71124;
  assign n71126 = ~n69723 & n69732;
  assign n71127 = ~n71125 & ~n71126;
  assign n71128 = ~n71119 & n71127;
  assign n71129 = ~n71114 & n71128;
  assign n71130 = n69761 & ~n71129;
  assign n71131 = n69697 & n69767;
  assign n71132 = ~n71130 & ~n71131;
  assign n71133 = n69744 & n71100;
  assign n71134 = ~n69715 & n71133;
  assign n71135 = n71132 & ~n71134;
  assign n71136 = ~n71111 & n71135;
  assign n71137 = ~pi2172 & ~n71136;
  assign n71138 = pi2172 & n71132;
  assign n71139 = ~n71111 & n71138;
  assign n71140 = ~n71134 & n71139;
  assign po2196 = n71137 | n71140;
  assign n71142 = ~n70319 & n70356;
  assign n71143 = ~n70336 & ~n71142;
  assign n71144 = ~n70352 & ~n71143;
  assign n71145 = n70326 & n70370;
  assign n71146 = ~n70511 & ~n71145;
  assign n71147 = n70352 & ~n71146;
  assign n71148 = ~n70326 & n70365;
  assign n71149 = ~n70531 & ~n71148;
  assign n71150 = ~n70334 & n71149;
  assign n71151 = ~n71147 & n71150;
  assign n71152 = ~n71144 & n71151;
  assign n71153 = ~n70506 & ~n70518;
  assign n71154 = n71152 & n71153;
  assign n71155 = n70307 & ~n71154;
  assign n71156 = n70320 & n70507;
  assign n71157 = n70339 & ~n71156;
  assign n71158 = n70352 & ~n71157;
  assign n71159 = ~n70326 & n70345;
  assign n71160 = ~n71158 & ~n71159;
  assign n71161 = n70313 & n70356;
  assign n71162 = n70326 & n70335;
  assign n71163 = ~n71161 & ~n71162;
  assign n71164 = n70352 & ~n71163;
  assign n71165 = n70352 & n70370;
  assign n71166 = ~n70326 & n71165;
  assign n71167 = ~n71164 & ~n71166;
  assign n71168 = n71160 & n71167;
  assign n71169 = ~n70307 & ~n71168;
  assign n71170 = ~n70365 & ~n70372;
  assign n71171 = ~n70512 & n71170;
  assign n71172 = n70380 & ~n71171;
  assign n71173 = ~n71169 & ~n71172;
  assign n71174 = ~n70334 & ~n70506;
  assign n71175 = ~n70352 & ~n71174;
  assign n71176 = n71173 & ~n71175;
  assign n71177 = ~n71155 & n71176;
  assign n71178 = ~pi2157 & n71177;
  assign n71179 = pi2157 & ~n71177;
  assign po2197 = n71178 | n71179;
  assign n71181 = n70812 & n70827;
  assign n71182 = ~n70943 & ~n71181;
  assign n71183 = ~n70844 & ~n71182;
  assign n71184 = ~n70835 & n70853;
  assign n71185 = ~n70828 & ~n71184;
  assign n71186 = ~n70878 & n71185;
  assign n71187 = n70844 & ~n71186;
  assign n71188 = ~n71183 & ~n71187;
  assign n71189 = ~n70858 & ~n70869;
  assign n71190 = n71188 & n71189;
  assign n71191 = ~n70850 & ~n71190;
  assign n71192 = n70835 & n70943;
  assign n71193 = n70825 & ~n70835;
  assign n71194 = ~n70973 & ~n71193;
  assign n71195 = n70844 & ~n71194;
  assign n71196 = ~n71192 & ~n71195;
  assign n71197 = ~n70844 & n70854;
  assign n71198 = n70829 & ~n71197;
  assign n71199 = ~n70878 & n71198;
  assign n71200 = ~n70835 & ~n71199;
  assign n71201 = n71196 & ~n71200;
  assign n71202 = n70850 & ~n71201;
  assign n71203 = ~n71191 & ~n71202;
  assign n71204 = n70812 & n70973;
  assign n71205 = ~n70886 & ~n71204;
  assign n71206 = ~n70844 & ~n71205;
  assign n71207 = n70844 & n71024;
  assign n71208 = n70835 & n71207;
  assign n71209 = ~n71206 & ~n71208;
  assign n71210 = n71203 & n71209;
  assign n71211 = ~pi2180 & ~n71210;
  assign n71212 = pi2180 & ~n71206;
  assign n71213 = n71203 & n71212;
  assign n71214 = ~n71208 & n71213;
  assign po2198 = n71211 | n71214;
  assign n71216 = n69998 & n70282;
  assign n71217 = n69979 & n71216;
  assign n71218 = n70023 & ~n70906;
  assign n71219 = ~n70008 & ~n71218;
  assign n71220 = ~n70280 & n71219;
  assign n71221 = ~n69979 & ~n71220;
  assign n71222 = n69998 & n70026;
  assign n71223 = ~n71221 & ~n71222;
  assign n71224 = n70004 & n70007;
  assign n71225 = ~n69998 & n70286;
  assign n71226 = ~n71224 & ~n71225;
  assign n71227 = ~n70910 & n71226;
  assign n71228 = n69979 & ~n71227;
  assign n71229 = n71223 & ~n71228;
  assign n71230 = n70020 & ~n71229;
  assign n71231 = ~n71217 & ~n71230;
  assign n71232 = ~n69998 & n70011;
  assign n71233 = ~n70279 & ~n71232;
  assign n71234 = n69979 & ~n71233;
  assign n71235 = ~n70009 & ~n71234;
  assign n71236 = ~n70042 & ~n71216;
  assign n71237 = n69998 & n70048;
  assign n71238 = ~n70286 & ~n71237;
  assign n71239 = ~n71224 & n71238;
  assign n71240 = ~n69979 & ~n71239;
  assign n71241 = ~n69998 & n70026;
  assign n71242 = ~n71240 & ~n71241;
  assign n71243 = n71236 & n71242;
  assign n71244 = n71235 & n71243;
  assign n71245 = ~n70020 & ~n71244;
  assign n71246 = ~n70065 & ~n70908;
  assign n71247 = ~n69979 & ~n71246;
  assign n71248 = ~n71245 & ~n71247;
  assign n71249 = n71231 & n71248;
  assign n71250 = pi2177 & n71249;
  assign n71251 = ~pi2177 & ~n71249;
  assign po2199 = n71250 | n71251;
  assign n71253 = ~n70326 & n70335;
  assign n71254 = ~n70362 & ~n71253;
  assign n71255 = ~n70352 & ~n71254;
  assign n71256 = n70352 & ~n70533;
  assign n71257 = ~n70522 & ~n71256;
  assign n71258 = ~n71255 & n71257;
  assign n71259 = n70307 & ~n71258;
  assign n71260 = n70345 & ~n70352;
  assign n71261 = ~n71259 & ~n71260;
  assign n71262 = ~n71148 & ~n71162;
  assign n71263 = n70352 & ~n71262;
  assign n71264 = n70352 & n70363;
  assign n71265 = n70326 & n70336;
  assign n71266 = n70333 & ~n70352;
  assign n71267 = ~n70510 & ~n71266;
  assign n71268 = ~n70313 & ~n71267;
  assign n71269 = ~n70511 & ~n71268;
  assign n71270 = ~n70334 & n71269;
  assign n71271 = ~n71265 & n71270;
  assign n71272 = ~n71264 & n71271;
  assign n71273 = ~n70307 & ~n71272;
  assign n71274 = ~n71263 & ~n71273;
  assign n71275 = n71261 & n71274;
  assign n71276 = pi2188 & ~n71275;
  assign n71277 = ~pi2188 & n71275;
  assign po2200 = n71276 | n71277;
  assign n71279 = ~n69778 & ~n71126;
  assign n71280 = n69697 & ~n71279;
  assign n71281 = ~n69761 & n69763;
  assign n71282 = ~n69697 & n71281;
  assign n71283 = n69709 & n71061;
  assign n71284 = ~n71116 & ~n71283;
  assign n71285 = ~n69732 & n71284;
  assign n71286 = n69697 & ~n71285;
  assign n71287 = ~n69723 & n69738;
  assign n71288 = ~n71286 & ~n71287;
  assign n71289 = ~n69761 & ~n71288;
  assign n71290 = ~n71282 & ~n71289;
  assign n71291 = ~n69727 & ~n69730;
  assign n71292 = ~n69723 & n69777;
  assign n71293 = ~n71096 & ~n71292;
  assign n71294 = n71291 & n71293;
  assign n71295 = ~n69697 & ~n71294;
  assign n71296 = ~n69703 & ~n69709;
  assign n71297 = ~n69697 & n71296;
  assign n71298 = n69723 & n71297;
  assign n71299 = ~n69723 & n71116;
  assign n71300 = ~n69730 & ~n71299;
  assign n71301 = ~n71123 & n71300;
  assign n71302 = ~n71298 & n71301;
  assign n71303 = n69697 & n71112;
  assign n71304 = n71302 & ~n71303;
  assign n71305 = n69761 & ~n71304;
  assign n71306 = ~n71295 & ~n71305;
  assign n71307 = n71290 & n71306;
  assign n71308 = ~n71280 & n71307;
  assign n71309 = pi2191 & n71308;
  assign n71310 = ~pi2191 & ~n71308;
  assign po2201 = n71309 | n71310;
  assign n71312 = pi7244 & pi9040;
  assign n71313 = pi7209 & ~pi9040;
  assign n71314 = ~n71312 & ~n71313;
  assign n71315 = ~pi2162 & ~n71314;
  assign n71316 = pi2162 & n71314;
  assign n71317 = ~n71315 & ~n71316;
  assign n71318 = pi7202 & pi9040;
  assign n71319 = pi7185 & ~pi9040;
  assign n71320 = ~n71318 & ~n71319;
  assign n71321 = pi2225 & n71320;
  assign n71322 = ~pi2225 & ~n71320;
  assign n71323 = ~n71321 & ~n71322;
  assign n71324 = pi7196 & pi9040;
  assign n71325 = pi7204 & ~pi9040;
  assign n71326 = ~n71324 & ~n71325;
  assign n71327 = ~pi2158 & ~n71326;
  assign n71328 = pi2158 & n71326;
  assign n71329 = ~n71327 & ~n71328;
  assign n71330 = pi7241 & pi9040;
  assign n71331 = pi7240 & ~pi9040;
  assign n71332 = ~n71330 & ~n71331;
  assign n71333 = ~pi2208 & n71332;
  assign n71334 = pi2208 & ~n71332;
  assign n71335 = ~n71333 & ~n71334;
  assign n71336 = pi7190 & pi9040;
  assign n71337 = pi7200 & ~pi9040;
  assign n71338 = ~n71336 & ~n71337;
  assign n71339 = ~pi2211 & ~n71338;
  assign n71340 = pi2211 & n71338;
  assign n71341 = ~n71339 & ~n71340;
  assign n71342 = n71335 & ~n71341;
  assign n71343 = n71329 & n71342;
  assign n71344 = ~n71323 & n71343;
  assign n71345 = pi7239 & pi9040;
  assign n71346 = pi7237 & ~pi9040;
  assign n71347 = ~n71345 & ~n71346;
  assign n71348 = ~pi2189 & n71347;
  assign n71349 = pi2189 & ~n71347;
  assign n71350 = ~n71348 & ~n71349;
  assign n71351 = n71335 & n71341;
  assign n71352 = ~n71329 & n71351;
  assign n71353 = ~n71323 & n71329;
  assign n71354 = n71341 & n71353;
  assign n71355 = ~n71335 & n71354;
  assign n71356 = ~n71352 & ~n71355;
  assign n71357 = n71329 & ~n71341;
  assign n71358 = n71323 & n71357;
  assign n71359 = ~n71335 & ~n71341;
  assign n71360 = ~n71329 & n71359;
  assign n71361 = ~n71323 & n71360;
  assign n71362 = ~n71358 & ~n71361;
  assign n71363 = n71356 & n71362;
  assign n71364 = n71350 & ~n71363;
  assign n71365 = ~n71329 & n71342;
  assign n71366 = ~n71335 & n71341;
  assign n71367 = n71323 & n71366;
  assign n71368 = n71335 & n71353;
  assign n71369 = ~n71367 & ~n71368;
  assign n71370 = ~n71365 & n71369;
  assign n71371 = ~n71350 & ~n71370;
  assign n71372 = n71323 & ~n71329;
  assign n71373 = n71341 & n71372;
  assign n71374 = ~n71335 & n71373;
  assign n71375 = ~n71371 & ~n71374;
  assign n71376 = ~n71364 & n71375;
  assign n71377 = ~n71344 & n71376;
  assign n71378 = ~n71317 & ~n71377;
  assign n71379 = n71329 & n71366;
  assign n71380 = n71323 & n71350;
  assign n71381 = n71379 & n71380;
  assign n71382 = n71350 & n71365;
  assign n71383 = n71329 & n71351;
  assign n71384 = n71350 & n71383;
  assign n71385 = ~n71382 & ~n71384;
  assign n71386 = ~n71323 & ~n71385;
  assign n71387 = ~n71381 & ~n71386;
  assign n71388 = ~n71335 & n71357;
  assign n71389 = ~n71323 & n71388;
  assign n71390 = n71323 & n71360;
  assign n71391 = ~n71389 & ~n71390;
  assign n71392 = n71323 & n71351;
  assign n71393 = ~n71323 & n71366;
  assign n71394 = ~n71392 & ~n71393;
  assign n71395 = ~n71388 & n71394;
  assign n71396 = ~n71352 & n71395;
  assign n71397 = ~n71350 & ~n71396;
  assign n71398 = ~n71329 & n71366;
  assign n71399 = ~n71323 & n71398;
  assign n71400 = ~n71397 & ~n71399;
  assign n71401 = n71391 & n71400;
  assign n71402 = n71387 & n71401;
  assign n71403 = n71317 & ~n71402;
  assign n71404 = n71323 & n71343;
  assign n71405 = n71351 & n71372;
  assign n71406 = ~n71404 & ~n71405;
  assign n71407 = n71350 & ~n71406;
  assign n71408 = ~n71403 & ~n71407;
  assign n71409 = ~n71341 & n71372;
  assign n71410 = n71335 & n71409;
  assign n71411 = ~n71389 & ~n71410;
  assign n71412 = ~n71350 & ~n71411;
  assign n71413 = n71408 & ~n71412;
  assign n71414 = ~n71378 & n71413;
  assign n71415 = pi2080 & ~n71414;
  assign n71416 = ~pi2080 & n71414;
  assign po2218 = n71415 | n71416;
  assign n71418 = pi7197 & ~pi9040;
  assign n71419 = pi7237 & pi9040;
  assign n71420 = ~n71418 & ~n71419;
  assign n71421 = ~pi2160 & n71420;
  assign n71422 = pi2160 & ~n71420;
  assign n71423 = ~n71421 & ~n71422;
  assign n71424 = pi7186 & pi9040;
  assign n71425 = pi7241 & ~pi9040;
  assign n71426 = ~n71424 & ~n71425;
  assign n71427 = pi2176 & n71426;
  assign n71428 = ~pi2176 & ~n71426;
  assign n71429 = ~n71427 & ~n71428;
  assign n71430 = pi7213 & pi9040;
  assign n71431 = pi7202 & ~pi9040;
  assign n71432 = ~n71430 & ~n71431;
  assign n71433 = ~pi2192 & ~n71432;
  assign n71434 = pi2192 & n71432;
  assign n71435 = ~n71433 & ~n71434;
  assign n71436 = pi7189 & ~pi9040;
  assign n71437 = pi7209 & pi9040;
  assign n71438 = ~n71436 & ~n71437;
  assign n71439 = ~pi2159 & n71438;
  assign n71440 = pi2159 & ~n71438;
  assign n71441 = ~n71439 & ~n71440;
  assign n71442 = n71435 & ~n71441;
  assign n71443 = ~n71429 & n71442;
  assign n71444 = pi7216 & pi9040;
  assign n71445 = pi7223 & ~pi9040;
  assign n71446 = ~n71444 & ~n71445;
  assign n71447 = pi2238 & n71446;
  assign n71448 = ~pi2238 & ~n71446;
  assign n71449 = ~n71447 & ~n71448;
  assign n71450 = n71443 & ~n71449;
  assign n71451 = ~n71429 & ~n71449;
  assign n71452 = n71441 & n71451;
  assign n71453 = ~n71435 & n71452;
  assign n71454 = ~n71450 & ~n71453;
  assign n71455 = ~n71435 & n71441;
  assign n71456 = n71429 & n71449;
  assign n71457 = n71455 & n71456;
  assign n71458 = n71435 & n71441;
  assign n71459 = ~n71429 & n71458;
  assign n71460 = n71449 & n71459;
  assign n71461 = ~n71457 & ~n71460;
  assign n71462 = n71454 & n71461;
  assign n71463 = ~n71423 & ~n71462;
  assign n71464 = ~n71435 & ~n71441;
  assign n71465 = ~n71429 & n71464;
  assign n71466 = n71449 & n71465;
  assign n71467 = ~n71459 & ~n71466;
  assign n71468 = ~n71423 & ~n71467;
  assign n71469 = n71423 & ~n71441;
  assign n71470 = ~n71449 & n71469;
  assign n71471 = n71429 & n71435;
  assign n71472 = n71449 & n71455;
  assign n71473 = ~n71471 & ~n71472;
  assign n71474 = n71423 & ~n71473;
  assign n71475 = ~n71470 & ~n71474;
  assign n71476 = n71429 & n71464;
  assign n71477 = ~n71449 & n71476;
  assign n71478 = n71475 & ~n71477;
  assign n71479 = ~n71441 & n71471;
  assign n71480 = n71449 & n71479;
  assign n71481 = n71478 & ~n71480;
  assign n71482 = ~n71468 & n71481;
  assign n71483 = pi7195 & pi9040;
  assign n71484 = pi7225 & ~pi9040;
  assign n71485 = ~n71483 & ~n71484;
  assign n71486 = ~pi2221 & ~n71485;
  assign n71487 = pi2221 & n71485;
  assign n71488 = ~n71486 & ~n71487;
  assign n71489 = ~n71482 & ~n71488;
  assign n71490 = ~n71429 & ~n71441;
  assign n71491 = n71423 & n71449;
  assign n71492 = n71488 & n71491;
  assign n71493 = n71490 & n71492;
  assign n71494 = n71423 & ~n71452;
  assign n71495 = ~n71435 & n71456;
  assign n71496 = ~n71442 & ~n71490;
  assign n71497 = ~n71449 & ~n71496;
  assign n71498 = n71429 & n71455;
  assign n71499 = ~n71423 & ~n71498;
  assign n71500 = ~n71497 & n71499;
  assign n71501 = ~n71495 & n71500;
  assign n71502 = ~n71494 & ~n71501;
  assign n71503 = n71429 & n71458;
  assign n71504 = n71449 & n71503;
  assign n71505 = ~n71502 & ~n71504;
  assign n71506 = n71488 & ~n71505;
  assign n71507 = ~n71493 & ~n71506;
  assign n71508 = ~n71489 & n71507;
  assign n71509 = ~n71463 & n71508;
  assign n71510 = n71423 & n71477;
  assign n71511 = n71509 & ~n71510;
  assign n71512 = pi2093 & ~n71511;
  assign n71513 = ~pi2093 & ~n71510;
  assign n71514 = n71508 & n71513;
  assign n71515 = ~n71463 & n71514;
  assign po2222 = n71512 | n71515;
  assign n71517 = ~n71368 & ~n71398;
  assign n71518 = n71350 & ~n71517;
  assign n71519 = n71323 & n71388;
  assign n71520 = ~n71354 & ~n71519;
  assign n71521 = ~n71518 & n71520;
  assign n71522 = ~n71329 & n71335;
  assign n71523 = ~n71329 & ~n71341;
  assign n71524 = ~n71323 & n71523;
  assign n71525 = n71323 & n71342;
  assign n71526 = ~n71524 & ~n71525;
  assign n71527 = ~n71522 & n71526;
  assign n71528 = ~n71379 & n71527;
  assign n71529 = ~n71350 & ~n71528;
  assign n71530 = n71521 & ~n71529;
  assign n71531 = n71317 & ~n71530;
  assign n71532 = ~n71323 & n71352;
  assign n71533 = ~n71410 & ~n71519;
  assign n71534 = ~n71532 & n71533;
  assign n71535 = ~n71350 & ~n71534;
  assign n71536 = ~n71531 & ~n71535;
  assign n71537 = ~n71329 & ~n71335;
  assign n71538 = n71350 & n71537;
  assign n71539 = n71323 & n71538;
  assign n71540 = n71323 & n71383;
  assign n71541 = ~n71350 & n71357;
  assign n71542 = ~n71323 & n71541;
  assign n71543 = ~n71540 & ~n71542;
  assign n71544 = n71329 & n71335;
  assign n71545 = n71323 & n71544;
  assign n71546 = ~n71360 & ~n71545;
  assign n71547 = n71350 & ~n71546;
  assign n71548 = n71350 & n71522;
  assign n71549 = ~n71323 & n71548;
  assign n71550 = ~n71547 & ~n71549;
  assign n71551 = n71543 & n71550;
  assign n71552 = ~n71317 & ~n71551;
  assign n71553 = ~n71539 & ~n71552;
  assign n71554 = ~n71355 & n71553;
  assign n71555 = n71536 & n71554;
  assign n71556 = ~pi2081 & ~n71555;
  assign n71557 = ~n71355 & ~n71531;
  assign n71558 = ~n71535 & n71557;
  assign n71559 = n71553 & n71558;
  assign n71560 = pi2081 & n71559;
  assign po2223 = n71556 | n71560;
  assign n71562 = pi7188 & pi9040;
  assign n71563 = pi7203 & ~pi9040;
  assign n71564 = ~n71562 & ~n71563;
  assign n71565 = pi2229 & n71564;
  assign n71566 = ~pi2229 & ~n71564;
  assign n71567 = ~n71565 & ~n71566;
  assign n71568 = pi7242 & pi9040;
  assign n71569 = pi7217 & ~pi9040;
  assign n71570 = ~n71568 & ~n71569;
  assign n71571 = ~pi2196 & n71570;
  assign n71572 = pi2196 & ~n71570;
  assign n71573 = ~n71571 & ~n71572;
  assign n71574 = pi7199 & pi9040;
  assign n71575 = pi7215 & ~pi9040;
  assign n71576 = ~n71574 & ~n71575;
  assign n71577 = ~pi2182 & n71576;
  assign n71578 = pi2182 & ~n71576;
  assign n71579 = ~n71577 & ~n71578;
  assign n71580 = pi7187 & pi9040;
  assign n71581 = pi7208 & ~pi9040;
  assign n71582 = ~n71580 & ~n71581;
  assign n71583 = pi2158 & n71582;
  assign n71584 = ~pi2158 & ~n71582;
  assign n71585 = ~n71583 & ~n71584;
  assign n71586 = pi7219 & ~pi9040;
  assign n71587 = pi7243 & pi9040;
  assign n71588 = ~n71586 & ~n71587;
  assign n71589 = pi2199 & n71588;
  assign n71590 = ~pi2199 & ~n71588;
  assign n71591 = ~n71589 & ~n71590;
  assign n71592 = ~n71585 & ~n71591;
  assign n71593 = n71579 & n71592;
  assign n71594 = n71573 & n71593;
  assign n71595 = ~n71573 & n71579;
  assign n71596 = ~n71585 & n71595;
  assign n71597 = n71591 & n71596;
  assign n71598 = ~n71594 & ~n71597;
  assign n71599 = n71567 & ~n71598;
  assign n71600 = pi7210 & ~pi9040;
  assign n71601 = pi7221 & pi9040;
  assign n71602 = ~n71600 & ~n71601;
  assign n71603 = ~pi2208 & ~n71602;
  assign n71604 = pi2208 & n71602;
  assign n71605 = ~n71603 & ~n71604;
  assign n71606 = n71573 & ~n71579;
  assign n71607 = n71585 & n71606;
  assign n71608 = ~n71591 & n71607;
  assign n71609 = ~n71585 & n71591;
  assign n71610 = ~n71579 & n71609;
  assign n71611 = n71567 & n71610;
  assign n71612 = ~n71608 & ~n71611;
  assign n71613 = n71573 & n71591;
  assign n71614 = n71579 & n71613;
  assign n71615 = ~n71591 & n71606;
  assign n71616 = ~n71614 & ~n71615;
  assign n71617 = ~n71567 & ~n71616;
  assign n71618 = ~n71567 & ~n71573;
  assign n71619 = n71592 & n71618;
  assign n71620 = n71579 & n71619;
  assign n71621 = ~n71573 & ~n71579;
  assign n71622 = n71585 & n71621;
  assign n71623 = n71591 & n71622;
  assign n71624 = ~pi2158 & n71582;
  assign n71625 = pi2158 & ~n71582;
  assign n71626 = ~n71624 & ~n71625;
  assign n71627 = ~n71591 & ~n71626;
  assign n71628 = n71579 & n71627;
  assign n71629 = n71567 & n71628;
  assign n71630 = ~n71623 & ~n71629;
  assign n71631 = ~n71620 & n71630;
  assign n71632 = ~n71617 & n71631;
  assign n71633 = n71612 & n71632;
  assign n71634 = n71605 & ~n71633;
  assign n71635 = ~n71567 & n71608;
  assign n71636 = n71573 & n71611;
  assign n71637 = ~n71635 & ~n71636;
  assign n71638 = ~n71634 & n71637;
  assign n71639 = ~n71599 & n71638;
  assign n71640 = n71567 & ~n71573;
  assign n71641 = ~n71579 & ~n71591;
  assign n71642 = n71640 & n71641;
  assign n71643 = n71567 & n71593;
  assign n71644 = ~n71642 & ~n71643;
  assign n71645 = n71591 & ~n71626;
  assign n71646 = ~n71579 & n71645;
  assign n71647 = n71567 & n71646;
  assign n71648 = n71579 & n71645;
  assign n71649 = n71573 & n71648;
  assign n71650 = ~n71647 & ~n71649;
  assign n71651 = ~n71579 & n71592;
  assign n71652 = ~n71573 & n71651;
  assign n71653 = ~n71594 & ~n71652;
  assign n71654 = ~n71573 & n71609;
  assign n71655 = n71579 & n71585;
  assign n71656 = ~n71654 & ~n71655;
  assign n71657 = ~n71567 & ~n71656;
  assign n71658 = n71653 & ~n71657;
  assign n71659 = n71650 & n71658;
  assign n71660 = n71644 & n71659;
  assign n71661 = ~n71605 & ~n71660;
  assign n71662 = n71639 & ~n71661;
  assign n71663 = ~pi2082 & ~n71662;
  assign n71664 = pi2082 & n71639;
  assign n71665 = ~n71661 & n71664;
  assign po2229 = n71663 | n71665;
  assign n71667 = ~n71579 & n71627;
  assign n71668 = ~n71573 & n71667;
  assign n71669 = ~n71573 & n71645;
  assign n71670 = n71573 & n71628;
  assign n71671 = ~n71669 & ~n71670;
  assign n71672 = ~n71567 & ~n71671;
  assign n71673 = ~n71668 & ~n71672;
  assign n71674 = n71567 & n71627;
  assign n71675 = ~n71573 & n71674;
  assign n71676 = ~n71643 & ~n71675;
  assign n71677 = n71673 & n71676;
  assign n71678 = ~n71573 & n71610;
  assign n71679 = n71573 & n71651;
  assign n71680 = ~n71678 & ~n71679;
  assign n71681 = n71677 & n71680;
  assign n71682 = n71605 & ~n71681;
  assign n71683 = ~n71567 & ~n71605;
  assign n71684 = ~n71591 & n71595;
  assign n71685 = n71579 & ~n71585;
  assign n71686 = ~n71684 & ~n71685;
  assign n71687 = n71683 & ~n71686;
  assign n71688 = ~n71608 & ~n71614;
  assign n71689 = ~n71579 & n71640;
  assign n71690 = ~n71627 & n71689;
  assign n71691 = ~n71611 & ~n71690;
  assign n71692 = n71688 & n71691;
  assign n71693 = ~n71605 & ~n71692;
  assign n71694 = n71579 & n71609;
  assign n71695 = ~n71567 & n71694;
  assign n71696 = n71573 & n71695;
  assign n71697 = n71573 & n71646;
  assign n71698 = ~n71679 & ~n71697;
  assign n71699 = ~n71567 & ~n71698;
  assign n71700 = ~n71696 & ~n71699;
  assign n71701 = n71567 & n71608;
  assign n71702 = n71700 & ~n71701;
  assign n71703 = ~n71693 & n71702;
  assign n71704 = ~n71687 & n71703;
  assign n71705 = ~n71682 & n71704;
  assign n71706 = n71567 & n71573;
  assign n71707 = n71648 & n71706;
  assign n71708 = n71705 & ~n71707;
  assign n71709 = ~pi2099 & ~n71708;
  assign n71710 = ~n71682 & ~n71707;
  assign n71711 = n71704 & n71710;
  assign n71712 = pi2099 & n71711;
  assign po2231 = n71709 | n71712;
  assign n71714 = pi7189 & pi9040;
  assign n71715 = pi7184 & ~pi9040;
  assign n71716 = ~n71714 & ~n71715;
  assign n71717 = ~pi2168 & ~n71716;
  assign n71718 = pi2168 & n71716;
  assign n71719 = ~n71717 & ~n71718;
  assign n71720 = pi7213 & ~pi9040;
  assign n71721 = pi7222 & pi9040;
  assign n71722 = ~n71720 & ~n71721;
  assign n71723 = ~pi2224 & ~n71722;
  assign n71724 = pi2224 & n71722;
  assign n71725 = ~n71723 & ~n71724;
  assign n71726 = ~n71719 & ~n71725;
  assign n71727 = pi7204 & pi9040;
  assign n71728 = pi7216 & ~pi9040;
  assign n71729 = ~n71727 & ~n71728;
  assign n71730 = ~pi2243 & ~n71729;
  assign n71731 = pi2243 & ~n71727;
  assign n71732 = ~n71728 & n71731;
  assign n71733 = ~n71730 & ~n71732;
  assign n71734 = pi7240 & pi9040;
  assign n71735 = pi7192 & ~pi9040;
  assign n71736 = ~n71734 & ~n71735;
  assign n71737 = ~pi2211 & n71736;
  assign n71738 = pi2211 & ~n71736;
  assign n71739 = ~n71737 & ~n71738;
  assign n71740 = pi7195 & ~pi9040;
  assign n71741 = pi7185 & pi9040;
  assign n71742 = ~n71740 & ~n71741;
  assign n71743 = ~pi2162 & n71742;
  assign n71744 = pi2162 & ~n71742;
  assign n71745 = ~n71743 & ~n71744;
  assign n71746 = ~n71739 & n71745;
  assign n71747 = ~n71733 & n71746;
  assign n71748 = pi7206 & pi9040;
  assign n71749 = pi7244 & ~pi9040;
  assign n71750 = ~n71748 & ~n71749;
  assign n71751 = ~pi2184 & n71750;
  assign n71752 = pi2184 & ~n71750;
  assign n71753 = ~n71751 & ~n71752;
  assign n71754 = ~n71745 & n71753;
  assign n71755 = ~n71739 & n71754;
  assign n71756 = n71733 & n71755;
  assign n71757 = ~n71745 & ~n71753;
  assign n71758 = ~n71733 & n71757;
  assign n71759 = ~n71756 & ~n71758;
  assign n71760 = ~n71747 & n71759;
  assign n71761 = n71726 & ~n71760;
  assign n71762 = ~n71733 & n71739;
  assign n71763 = n71753 & n71762;
  assign n71764 = n71745 & n71753;
  assign n71765 = ~n71739 & n71764;
  assign n71766 = n71733 & n71765;
  assign n71767 = ~n71763 & ~n71766;
  assign n71768 = n71739 & n71754;
  assign n71769 = ~n71739 & n71757;
  assign n71770 = ~n71768 & ~n71769;
  assign n71771 = n71767 & n71770;
  assign n71772 = n71719 & ~n71771;
  assign n71773 = n71745 & ~n71753;
  assign n71774 = n71739 & n71773;
  assign n71775 = n71733 & n71774;
  assign n71776 = ~n71772 & ~n71775;
  assign n71777 = ~n71725 & ~n71776;
  assign n71778 = ~n71761 & ~n71777;
  assign n71779 = n71719 & ~n71733;
  assign n71780 = ~n71739 & n71779;
  assign n71781 = ~n71753 & n71780;
  assign n71782 = n71754 & n71762;
  assign n71783 = ~n71781 & ~n71782;
  assign n71784 = n71739 & n71764;
  assign n71785 = ~n71757 & ~n71764;
  assign n71786 = n71733 & ~n71785;
  assign n71787 = ~n71784 & ~n71786;
  assign n71788 = ~n71719 & ~n71787;
  assign n71789 = ~n71739 & n71773;
  assign n71790 = ~n71747 & ~n71789;
  assign n71791 = ~n71756 & n71790;
  assign n71792 = n71719 & ~n71791;
  assign n71793 = ~n71788 & ~n71792;
  assign n71794 = ~n71719 & ~n71733;
  assign n71795 = n71754 & n71794;
  assign n71796 = n71733 & n71784;
  assign n71797 = n71739 & ~n71745;
  assign n71798 = ~n71753 & n71797;
  assign n71799 = n71733 & n71798;
  assign n71800 = ~n71796 & ~n71799;
  assign n71801 = ~n71753 & n71762;
  assign n71802 = n71745 & n71801;
  assign n71803 = n71800 & ~n71802;
  assign n71804 = ~n71795 & n71803;
  assign n71805 = n71793 & n71804;
  assign n71806 = n71725 & ~n71805;
  assign n71807 = n71783 & ~n71806;
  assign n71808 = n71778 & n71807;
  assign n71809 = pi2091 & ~n71808;
  assign n71810 = ~pi2091 & n71783;
  assign n71811 = n71778 & n71810;
  assign n71812 = ~n71806 & n71811;
  assign po2235 = n71809 | n71812;
  assign n71814 = ~n71323 & n71365;
  assign n71815 = ~n71389 & ~n71814;
  assign n71816 = ~n71374 & n71815;
  assign n71817 = n71350 & ~n71816;
  assign n71818 = ~n71323 & ~n71350;
  assign n71819 = n71360 & n71818;
  assign n71820 = ~n71350 & n71405;
  assign n71821 = ~n71819 & ~n71820;
  assign n71822 = ~n71384 & ~n71390;
  assign n71823 = ~n71343 & ~n71393;
  assign n71824 = ~n71350 & ~n71823;
  assign n71825 = ~n71355 & ~n71824;
  assign n71826 = n71822 & n71825;
  assign n71827 = n71317 & ~n71826;
  assign n71828 = ~n71329 & n71341;
  assign n71829 = ~n71522 & ~n71828;
  assign n71830 = n71323 & ~n71829;
  assign n71831 = ~n71323 & n71351;
  assign n71832 = ~n71388 & ~n71831;
  assign n71833 = ~n71350 & ~n71832;
  assign n71834 = n71323 & n71341;
  assign n71835 = ~n71398 & ~n71834;
  assign n71836 = ~n71342 & n71835;
  assign n71837 = n71350 & ~n71836;
  assign n71838 = ~n71833 & ~n71837;
  assign n71839 = ~n71830 & n71838;
  assign n71840 = ~n71317 & ~n71839;
  assign n71841 = ~n71827 & ~n71840;
  assign n71842 = n71821 & n71841;
  assign n71843 = ~n71817 & n71842;
  assign n71844 = ~pi2088 & ~n71843;
  assign n71845 = pi2088 & n71821;
  assign n71846 = ~n71817 & n71845;
  assign n71847 = n71841 & n71846;
  assign po2238 = n71844 | n71847;
  assign n71849 = ~n71733 & ~n71739;
  assign n71850 = n71753 & n71849;
  assign n71851 = n71745 & n71850;
  assign n71852 = n71733 & n71757;
  assign n71853 = ~n71851 & ~n71852;
  assign n71854 = n71719 & ~n71853;
  assign n71855 = n71733 & n71746;
  assign n71856 = ~n71769 & ~n71855;
  assign n71857 = ~n71782 & n71856;
  assign n71858 = n71719 & ~n71857;
  assign n71859 = ~n71733 & ~n71753;
  assign n71860 = n71797 & n71859;
  assign n71861 = ~n71733 & n71789;
  assign n71862 = n71739 & n71745;
  assign n71863 = ~n71754 & ~n71862;
  assign n71864 = n71733 & ~n71863;
  assign n71865 = ~n71861 & ~n71864;
  assign n71866 = ~n71860 & n71865;
  assign n71867 = ~n71719 & ~n71866;
  assign n71868 = ~n71858 & ~n71867;
  assign n71869 = n71725 & ~n71868;
  assign n71870 = n71719 & n71802;
  assign n71871 = ~n71719 & n71784;
  assign n71872 = ~n71733 & n71871;
  assign n71873 = ~n71733 & n71755;
  assign n71874 = ~n71719 & n71873;
  assign n71875 = ~n71872 & ~n71874;
  assign n71876 = ~n71870 & n71875;
  assign n71877 = n71745 & n71779;
  assign n71878 = ~n71733 & ~n71745;
  assign n71879 = ~n71739 & n71878;
  assign n71880 = ~n71855 & ~n71879;
  assign n71881 = ~n71719 & ~n71880;
  assign n71882 = ~n71795 & ~n71881;
  assign n71883 = ~n71799 & ~n71873;
  assign n71884 = n71719 & n71733;
  assign n71885 = n71797 & n71884;
  assign n71886 = n71719 & n71774;
  assign n71887 = ~n71885 & ~n71886;
  assign n71888 = n71883 & n71887;
  assign n71889 = n71882 & n71888;
  assign n71890 = ~n71877 & n71889;
  assign n71891 = ~n71725 & ~n71890;
  assign n71892 = n71876 & ~n71891;
  assign n71893 = ~n71869 & n71892;
  assign n71894 = ~n71854 & n71893;
  assign n71895 = ~pi2104 & ~n71894;
  assign n71896 = pi2104 & n71894;
  assign po2239 = n71895 | n71896;
  assign n71898 = ~n71636 & ~n71642;
  assign n71899 = n71573 & n71674;
  assign n71900 = n71591 & n71595;
  assign n71901 = ~n71694 & ~n71900;
  assign n71902 = n71567 & ~n71901;
  assign n71903 = ~n71899 & ~n71902;
  assign n71904 = ~n71567 & n71645;
  assign n71905 = n71573 & n71904;
  assign n71906 = ~n71567 & n71593;
  assign n71907 = ~n71905 & ~n71906;
  assign n71908 = n71903 & n71907;
  assign n71909 = n71591 & n71606;
  assign n71910 = ~n71594 & ~n71909;
  assign n71911 = ~n71652 & n71910;
  assign n71912 = n71908 & n71911;
  assign n71913 = ~n71605 & ~n71912;
  assign n71914 = ~n71608 & ~n71694;
  assign n71915 = ~n71654 & n71914;
  assign n71916 = ~n71567 & ~n71915;
  assign n71917 = n71585 & n71595;
  assign n71918 = ~n71591 & n71917;
  assign n71919 = ~n71623 & ~n71918;
  assign n71920 = ~n71707 & n71919;
  assign n71921 = n71567 & n71651;
  assign n71922 = n71920 & ~n71921;
  assign n71923 = ~n71916 & n71922;
  assign n71924 = n71605 & ~n71923;
  assign n71925 = ~n71594 & n71919;
  assign n71926 = ~n71567 & ~n71925;
  assign n71927 = ~n71924 & ~n71926;
  assign n71928 = ~n71913 & n71927;
  assign n71929 = n71898 & n71928;
  assign n71930 = pi2085 & ~n71929;
  assign n71931 = ~pi2085 & n71929;
  assign po2240 = n71930 | n71931;
  assign n71933 = pi7215 & pi9040;
  assign n71934 = pi7183 & ~pi9040;
  assign n71935 = ~n71933 & ~n71934;
  assign n71936 = pi2244 & n71935;
  assign n71937 = ~pi2244 & ~n71935;
  assign n71938 = ~n71936 & ~n71937;
  assign n71939 = pi7193 & pi9040;
  assign n71940 = pi7187 & ~pi9040;
  assign n71941 = ~n71939 & ~n71940;
  assign n71942 = pi2185 & n71941;
  assign n71943 = ~pi2185 & ~n71941;
  assign n71944 = ~n71942 & ~n71943;
  assign n71945 = pi7180 & pi9040;
  assign n71946 = pi7198 & ~pi9040;
  assign n71947 = ~n71945 & ~n71946;
  assign n71948 = ~pi2164 & n71947;
  assign n71949 = pi2164 & ~n71947;
  assign n71950 = ~n71948 & ~n71949;
  assign n71951 = n71944 & n71950;
  assign n71952 = pi7219 & pi9040;
  assign n71953 = pi7226 & ~pi9040;
  assign n71954 = ~n71952 & ~n71953;
  assign n71955 = pi2242 & n71954;
  assign n71956 = ~pi2242 & ~n71954;
  assign n71957 = ~n71955 & ~n71956;
  assign n71958 = pi7191 & pi9040;
  assign n71959 = pi7242 & ~pi9040;
  assign n71960 = ~n71958 & ~n71959;
  assign n71961 = ~pi2174 & n71960;
  assign n71962 = pi2174 & ~n71960;
  assign n71963 = ~n71961 & ~n71962;
  assign n71964 = n71957 & ~n71963;
  assign n71965 = n71951 & n71964;
  assign n71966 = n71957 & n71963;
  assign n71967 = ~n71944 & n71966;
  assign n71968 = ~n71965 & ~n71967;
  assign n71969 = ~n71938 & ~n71968;
  assign n71970 = pi7188 & ~pi9040;
  assign n71971 = pi7211 & pi9040;
  assign n71972 = ~n71970 & ~n71971;
  assign n71973 = ~pi2178 & ~n71972;
  assign n71974 = pi2178 & n71972;
  assign n71975 = ~n71973 & ~n71974;
  assign n71976 = n71938 & ~n71957;
  assign n71977 = n71944 & n71976;
  assign n71978 = n71951 & n71963;
  assign n71979 = n71944 & ~n71950;
  assign n71980 = ~n71963 & n71979;
  assign n71981 = ~n71978 & ~n71980;
  assign n71982 = ~n71944 & n71950;
  assign n71983 = ~n71963 & n71982;
  assign n71984 = n71957 & n71983;
  assign n71985 = n71981 & ~n71984;
  assign n71986 = n71938 & ~n71985;
  assign n71987 = ~n71977 & ~n71986;
  assign n71988 = ~n71944 & ~n71950;
  assign n71989 = n71963 & n71988;
  assign n71990 = n71957 & n71989;
  assign n71991 = n71987 & ~n71990;
  assign n71992 = ~n71957 & n71982;
  assign n71993 = ~n71963 & n71988;
  assign n71994 = ~n71992 & ~n71993;
  assign n71995 = ~n71938 & ~n71994;
  assign n71996 = n71963 & n71979;
  assign n71997 = ~n71957 & n71996;
  assign n71998 = ~n71995 & ~n71997;
  assign n71999 = n71991 & n71998;
  assign n72000 = n71975 & ~n71999;
  assign n72001 = ~n71969 & ~n72000;
  assign n72002 = n71938 & ~n71975;
  assign n72003 = ~n71994 & n72002;
  assign n72004 = n71963 & n71982;
  assign n72005 = ~n71996 & ~n72004;
  assign n72006 = n71957 & ~n72005;
  assign n72007 = ~n71965 & ~n72006;
  assign n72008 = ~n71975 & ~n72007;
  assign n72009 = ~n72003 & ~n72008;
  assign n72010 = ~n71938 & ~n71975;
  assign n72011 = n71951 & ~n71957;
  assign n72012 = ~n71989 & ~n72011;
  assign n72013 = n71944 & ~n71963;
  assign n72014 = n72012 & ~n72013;
  assign n72015 = n72010 & ~n72014;
  assign n72016 = n72009 & ~n72015;
  assign n72017 = n72001 & n72016;
  assign n72018 = ~pi2086 & ~n72017;
  assign n72019 = pi2086 & n72009;
  assign n72020 = n72001 & n72019;
  assign n72021 = ~n72015 & n72020;
  assign po2241 = n72018 | n72021;
  assign n72023 = ~n71398 & ~n71814;
  assign n72024 = ~n71350 & ~n72023;
  assign n72025 = n71406 & ~n72024;
  assign n72026 = ~n71323 & n71350;
  assign n72027 = ~n71335 & n72026;
  assign n72028 = n72025 & ~n72027;
  assign n72029 = n71317 & ~n72028;
  assign n72030 = n71350 & n71390;
  assign n72031 = ~n71368 & ~n71819;
  assign n72032 = ~n71383 & ~n71398;
  assign n72033 = ~n71831 & n72032;
  assign n72034 = n71350 & ~n72033;
  assign n72035 = ~n71350 & n71379;
  assign n72036 = n71533 & ~n72035;
  assign n72037 = ~n72034 & n72036;
  assign n72038 = n72031 & n72037;
  assign n72039 = ~n71317 & ~n72038;
  assign n72040 = ~n72030 & ~n72039;
  assign n72041 = ~n72029 & n72040;
  assign n72042 = n71383 & n71818;
  assign n72043 = n71323 & n71541;
  assign n72044 = ~n72042 & ~n72043;
  assign n72045 = ~n71820 & n72044;
  assign n72046 = n72041 & n72045;
  assign n72047 = ~pi2087 & ~n72046;
  assign n72048 = pi2087 & n72045;
  assign n72049 = n72040 & n72048;
  assign n72050 = ~n72029 & n72049;
  assign po2242 = n72047 | n72050;
  assign n72052 = n71719 & n71757;
  assign n72053 = ~n71733 & n72052;
  assign n72054 = ~n71851 & ~n72053;
  assign n72055 = n71733 & ~n71753;
  assign n72056 = ~n71739 & n72055;
  assign n72057 = ~n71733 & n71745;
  assign n72058 = ~n71850 & ~n72057;
  assign n72059 = ~n71719 & ~n72058;
  assign n72060 = ~n72056 & ~n72059;
  assign n72061 = n72054 & n72060;
  assign n72062 = n71725 & ~n72061;
  assign n72063 = ~n71755 & ~n71799;
  assign n72064 = ~n71733 & n71773;
  assign n72065 = n72063 & ~n72064;
  assign n72066 = n71719 & ~n72065;
  assign n72067 = n71757 & n71794;
  assign n72068 = ~n71782 & ~n72067;
  assign n72069 = ~n72066 & n72068;
  assign n72070 = ~n71765 & ~n71775;
  assign n72071 = ~n71719 & ~n72070;
  assign n72072 = n72069 & ~n72071;
  assign n72073 = ~n71725 & ~n72072;
  assign n72074 = ~n72062 & ~n72073;
  assign n72075 = ~n71733 & n71764;
  assign n72076 = n71733 & ~n71770;
  assign n72077 = ~n72075 & ~n72076;
  assign n72078 = ~n71719 & ~n72077;
  assign n72079 = ~n71784 & ~n71789;
  assign n72080 = ~n71755 & n72079;
  assign n72081 = n71884 & ~n72080;
  assign n72082 = ~n72078 & ~n72081;
  assign n72083 = n72074 & n72082;
  assign n72084 = ~pi2095 & ~n72083;
  assign n72085 = ~n72073 & n72082;
  assign n72086 = pi2095 & n72085;
  assign n72087 = ~n72062 & n72086;
  assign po2244 = n72084 | n72087;
  assign n72089 = ~n71938 & n71957;
  assign n72090 = ~n71982 & ~n71996;
  assign n72091 = n72089 & ~n72090;
  assign n72092 = ~n71938 & n71963;
  assign n72093 = n71982 & n72092;
  assign n72094 = ~n72091 & ~n72093;
  assign n72095 = n71975 & ~n72094;
  assign n72096 = ~n71957 & ~n71963;
  assign n72097 = ~n71950 & n72096;
  assign n72098 = n71944 & n72097;
  assign n72099 = ~n72013 & ~n72096;
  assign n72100 = n71938 & ~n72099;
  assign n72101 = ~n71957 & n71963;
  assign n72102 = n71950 & n72101;
  assign n72103 = n71944 & n72102;
  assign n72104 = ~n72100 & ~n72103;
  assign n72105 = ~n72098 & n72104;
  assign n72106 = n71975 & ~n72105;
  assign n72107 = ~n72095 & ~n72106;
  assign n72108 = ~n71950 & n71964;
  assign n72109 = ~n71944 & n72108;
  assign n72110 = ~n71957 & n71989;
  assign n72111 = ~n72109 & ~n72110;
  assign n72112 = ~n71938 & ~n72111;
  assign n72113 = n71957 & n72004;
  assign n72114 = ~n71957 & n72013;
  assign n72115 = ~n72113 & ~n72114;
  assign n72116 = n71938 & ~n72115;
  assign n72117 = ~n71951 & ~n72013;
  assign n72118 = n71957 & ~n72117;
  assign n72119 = ~n71989 & ~n72118;
  assign n72120 = ~n71938 & ~n72119;
  assign n72121 = ~n71950 & ~n71957;
  assign n72122 = n72092 & n72121;
  assign n72123 = n71950 & ~n71963;
  assign n72124 = ~n71989 & ~n72123;
  assign n72125 = ~n71957 & ~n72124;
  assign n72126 = n71938 & n71957;
  assign n72127 = n71979 & n72126;
  assign n72128 = n71963 & n72127;
  assign n72129 = ~n72125 & ~n72128;
  assign n72130 = ~n72122 & n72129;
  assign n72131 = ~n72120 & n72130;
  assign n72132 = ~n72109 & n72131;
  assign n72133 = ~n71975 & ~n72132;
  assign n72134 = ~n72116 & ~n72133;
  assign n72135 = ~n72112 & n72134;
  assign n72136 = n72107 & n72135;
  assign n72137 = pi2084 & n72136;
  assign n72138 = ~pi2084 & ~n72136;
  assign po2245 = n72137 | n72138;
  assign n72140 = ~n71678 & ~n71684;
  assign n72141 = n71605 & ~n72140;
  assign n72142 = ~n71607 & ~n71615;
  assign n72143 = ~n71667 & n72142;
  assign n72144 = ~n71567 & ~n72143;
  assign n72145 = n71605 & n72144;
  assign n72146 = ~n72141 & ~n72145;
  assign n72147 = n71610 & n71618;
  assign n72148 = ~n71620 & ~n72147;
  assign n72149 = ~n71614 & ~n71655;
  assign n72150 = n71567 & ~n72149;
  assign n72151 = n71605 & n72150;
  assign n72152 = n72148 & ~n72151;
  assign n72153 = n71573 & n71610;
  assign n72154 = n71573 & n71592;
  assign n72155 = ~n71597 & ~n72154;
  assign n72156 = n71567 & ~n72155;
  assign n72157 = ~n71608 & ~n71623;
  assign n72158 = n71573 & n71609;
  assign n72159 = ~n71648 & ~n72158;
  assign n72160 = ~n71567 & ~n72159;
  assign n72161 = n72157 & ~n72160;
  assign n72162 = ~n72156 & n72161;
  assign n72163 = ~n72153 & n72162;
  assign n72164 = ~n71605 & ~n72163;
  assign n72165 = ~n71652 & n71919;
  assign n72166 = n71567 & ~n72165;
  assign n72167 = ~n72164 & ~n72166;
  assign n72168 = n72152 & n72167;
  assign n72169 = n72146 & n72168;
  assign n72170 = ~pi2097 & ~n72169;
  assign n72171 = pi2097 & n72152;
  assign n72172 = n72146 & n72171;
  assign n72173 = n72167 & n72172;
  assign po2246 = n72170 | n72173;
  assign n72175 = pi7222 & ~pi9040;
  assign n72176 = pi7179 & pi9040;
  assign n72177 = ~n72175 & ~n72176;
  assign n72178 = pi2159 & n72177;
  assign n72179 = ~pi2159 & ~n72177;
  assign n72180 = ~n72178 & ~n72179;
  assign n72181 = pi7201 & ~pi9040;
  assign n72182 = pi7184 & pi9040;
  assign n72183 = ~n72181 & ~n72182;
  assign n72184 = ~pi2224 & n72183;
  assign n72185 = pi2224 & ~n72183;
  assign n72186 = ~n72184 & ~n72185;
  assign n72187 = pi7182 & pi9040;
  assign n72188 = pi7196 & ~pi9040;
  assign n72189 = ~n72187 & ~n72188;
  assign n72190 = pi2176 & n72189;
  assign n72191 = ~pi2176 & ~n72189;
  assign n72192 = ~n72190 & ~n72191;
  assign n72193 = n72186 & n72192;
  assign n72194 = pi7192 & pi9040;
  assign n72195 = pi7220 & ~pi9040;
  assign n72196 = ~n72194 & ~n72195;
  assign n72197 = pi2212 & n72196;
  assign n72198 = ~pi2212 & ~n72196;
  assign n72199 = ~n72197 & ~n72198;
  assign n72200 = pi7190 & ~pi9040;
  assign n72201 = pi7225 & pi9040;
  assign n72202 = ~n72200 & ~n72201;
  assign n72203 = pi2218 & n72202;
  assign n72204 = ~pi2218 & ~n72202;
  assign n72205 = ~n72203 & ~n72204;
  assign n72206 = ~n72199 & ~n72205;
  assign n72207 = n72193 & n72206;
  assign n72208 = pi7223 & pi9040;
  assign n72209 = pi7206 & ~pi9040;
  assign n72210 = ~n72208 & ~n72209;
  assign n72211 = ~pi2184 & n72210;
  assign n72212 = pi2184 & ~n72210;
  assign n72213 = ~n72211 & ~n72212;
  assign n72214 = ~n72186 & ~n72192;
  assign n72215 = ~n72213 & n72214;
  assign n72216 = n72199 & n72213;
  assign n72217 = ~n72192 & n72216;
  assign n72218 = n72186 & n72217;
  assign n72219 = ~n72215 & ~n72218;
  assign n72220 = ~n72186 & n72192;
  assign n72221 = n72199 & n72220;
  assign n72222 = n72219 & ~n72221;
  assign n72223 = ~n72205 & ~n72222;
  assign n72224 = ~n72186 & n72213;
  assign n72225 = ~n72199 & n72205;
  assign n72226 = n72224 & n72225;
  assign n72227 = n72213 & n72214;
  assign n72228 = ~n72199 & n72227;
  assign n72229 = ~n72226 & ~n72228;
  assign n72230 = ~n72223 & n72229;
  assign n72231 = ~n72207 & n72230;
  assign n72232 = n72193 & ~n72213;
  assign n72233 = ~n72199 & n72232;
  assign n72234 = ~n72213 & n72220;
  assign n72235 = n72199 & n72234;
  assign n72236 = ~n72233 & ~n72235;
  assign n72237 = n72231 & n72236;
  assign n72238 = ~n72180 & ~n72237;
  assign n72239 = ~n72199 & n72213;
  assign n72240 = n72192 & n72239;
  assign n72241 = ~n72186 & n72240;
  assign n72242 = ~n72232 & ~n72241;
  assign n72243 = ~n72205 & ~n72242;
  assign n72244 = n72193 & n72216;
  assign n72245 = ~n72192 & n72239;
  assign n72246 = n72186 & n72245;
  assign n72247 = ~n72244 & ~n72246;
  assign n72248 = ~n72186 & n72216;
  assign n72249 = ~n72199 & n72234;
  assign n72250 = ~n72248 & ~n72249;
  assign n72251 = n72205 & ~n72250;
  assign n72252 = n72247 & ~n72251;
  assign n72253 = ~n72243 & n72252;
  assign n72254 = n72180 & ~n72253;
  assign n72255 = ~n72186 & ~n72213;
  assign n72256 = n72199 & n72255;
  assign n72257 = n72186 & ~n72213;
  assign n72258 = ~n72199 & n72257;
  assign n72259 = ~n72256 & ~n72258;
  assign n72260 = ~n72205 & ~n72259;
  assign n72261 = n72186 & ~n72192;
  assign n72262 = ~n72213 & n72261;
  assign n72263 = n72199 & n72262;
  assign n72264 = ~n72244 & ~n72263;
  assign n72265 = ~n72227 & n72264;
  assign n72266 = n72205 & ~n72265;
  assign n72267 = ~n72260 & ~n72266;
  assign n72268 = ~n72192 & n72213;
  assign n72269 = n72205 & n72268;
  assign n72270 = ~n72199 & n72269;
  assign n72271 = n72267 & ~n72270;
  assign n72272 = ~n72254 & n72271;
  assign n72273 = ~n72238 & n72272;
  assign n72274 = ~pi2094 & ~n72273;
  assign n72275 = pi2094 & n72273;
  assign po2247 = n72274 | n72275;
  assign n72277 = ~n71450 & ~n71457;
  assign n72278 = n71423 & ~n72277;
  assign n72279 = ~n71510 & ~n72278;
  assign n72280 = ~n71429 & ~n71435;
  assign n72281 = ~n71423 & n72280;
  assign n72282 = n71449 & n72281;
  assign n72283 = n71449 & n71464;
  assign n72284 = ~n72280 & ~n72283;
  assign n72285 = n71429 & ~n71449;
  assign n72286 = n71435 & n72285;
  assign n72287 = n72284 & ~n72286;
  assign n72288 = ~n71423 & ~n72287;
  assign n72289 = ~n71460 & ~n72288;
  assign n72290 = ~n71488 & ~n72289;
  assign n72291 = n71423 & n71442;
  assign n72292 = n71449 & n72291;
  assign n72293 = n71423 & n71498;
  assign n72294 = ~n72292 & ~n72293;
  assign n72295 = ~n71488 & ~n72294;
  assign n72296 = ~n72290 & ~n72295;
  assign n72297 = ~n72282 & n72296;
  assign n72298 = ~n71452 & ~n71476;
  assign n72299 = ~n71503 & n72298;
  assign n72300 = n71423 & ~n72299;
  assign n72301 = n71435 & n71451;
  assign n72302 = ~n71449 & n71498;
  assign n72303 = ~n71479 & ~n72302;
  assign n72304 = ~n71423 & ~n72303;
  assign n72305 = ~n72301 & ~n72304;
  assign n72306 = ~n72300 & n72305;
  assign n72307 = ~n71466 & ~n71504;
  assign n72308 = n72306 & n72307;
  assign n72309 = n71488 & ~n72308;
  assign n72310 = n72297 & ~n72309;
  assign n72311 = n72279 & n72310;
  assign n72312 = ~pi2101 & ~n72311;
  assign n72313 = pi2101 & n72297;
  assign n72314 = n72279 & n72313;
  assign n72315 = ~n72309 & n72314;
  assign po2248 = n72312 | n72315;
  assign n72317 = ~n71719 & ~n72079;
  assign n72318 = n71733 & n71769;
  assign n72319 = ~n72317 & ~n72318;
  assign n72320 = n71733 & ~n71745;
  assign n72321 = ~n71797 & ~n72320;
  assign n72322 = ~n71765 & n72321;
  assign n72323 = n71719 & ~n72322;
  assign n72324 = n72319 & ~n72323;
  assign n72325 = ~n71725 & ~n72324;
  assign n72326 = ~n71733 & n71798;
  assign n72327 = ~n71719 & n72326;
  assign n72328 = ~n71874 & ~n72327;
  assign n72329 = ~n71870 & n72328;
  assign n72330 = ~n71802 & ~n71850;
  assign n72331 = n71719 & n71879;
  assign n72332 = n71733 & n71789;
  assign n72333 = ~n71719 & n71797;
  assign n72334 = ~n72332 & ~n72333;
  assign n72335 = ~n71796 & n72334;
  assign n72336 = ~n72331 & n72335;
  assign n72337 = n72330 & n72336;
  assign n72338 = ~n71886 & n72337;
  assign n72339 = n71725 & ~n72338;
  assign n72340 = n72329 & ~n72339;
  assign n72341 = ~n72325 & n72340;
  assign n72342 = ~pi2090 & ~n72341;
  assign n72343 = pi2090 & n72329;
  assign n72344 = ~n72325 & n72343;
  assign n72345 = ~n72339 & n72344;
  assign po2250 = n72342 | n72345;
  assign n72347 = ~n71449 & n71479;
  assign n72348 = n71449 & n71490;
  assign n72349 = ~n71476 & ~n72348;
  assign n72350 = ~n71423 & ~n72349;
  assign n72351 = ~n72347 & ~n72350;
  assign n72352 = n71423 & ~n71449;
  assign n72353 = ~n71441 & n72352;
  assign n72354 = n71435 & n72353;
  assign n72355 = n71458 & n71491;
  assign n72356 = ~n72354 & ~n72355;
  assign n72357 = ~n72293 & n72356;
  assign n72358 = ~n71453 & ~n71466;
  assign n72359 = n71441 & n71456;
  assign n72360 = n72358 & ~n72359;
  assign n72361 = n72357 & n72360;
  assign n72362 = n72351 & n72361;
  assign n72363 = ~n71488 & ~n72362;
  assign n72364 = ~n71429 & n71455;
  assign n72365 = ~n71476 & ~n72364;
  assign n72366 = n71449 & ~n72365;
  assign n72367 = ~n71503 & ~n72301;
  assign n72368 = n71429 & ~n71441;
  assign n72369 = n71449 & n72368;
  assign n72370 = n72367 & ~n72369;
  assign n72371 = ~n71423 & ~n72370;
  assign n72372 = ~n71449 & n71464;
  assign n72373 = ~n71429 & n71449;
  assign n72374 = ~n71441 & n72373;
  assign n72375 = n71435 & n72374;
  assign n72376 = ~n72372 & ~n72375;
  assign n72377 = n71423 & ~n72376;
  assign n72378 = ~n71449 & n71459;
  assign n72379 = ~n72377 & ~n72378;
  assign n72380 = ~n72371 & n72379;
  assign n72381 = ~n72366 & n72380;
  assign n72382 = n71488 & ~n72381;
  assign n72383 = ~n71423 & n71452;
  assign n72384 = ~n72382 & ~n72383;
  assign n72385 = n71471 & n72352;
  assign n72386 = ~n71441 & n72385;
  assign n72387 = n72384 & ~n72386;
  assign n72388 = ~n72363 & n72387;
  assign n72389 = ~pi2098 & ~n72388;
  assign n72390 = pi2098 & n72384;
  assign n72391 = ~n72363 & n72390;
  assign n72392 = ~n72386 & n72391;
  assign po2251 = n72389 | n72392;
  assign n72394 = pi7208 & pi9040;
  assign n72395 = pi7191 & ~pi9040;
  assign n72396 = ~n72394 & ~n72395;
  assign n72397 = ~pi2185 & ~n72396;
  assign n72398 = pi2185 & n72396;
  assign n72399 = ~n72397 & ~n72398;
  assign n72400 = pi7243 & ~pi9040;
  assign n72401 = pi7238 & pi9040;
  assign n72402 = ~n72400 & ~n72401;
  assign n72403 = ~pi2192 & ~n72402;
  assign n72404 = pi2192 & n72402;
  assign n72405 = ~n72403 & ~n72404;
  assign n72406 = pi7226 & pi9040;
  assign n72407 = pi7221 & ~pi9040;
  assign n72408 = ~n72406 & ~n72407;
  assign n72409 = ~pi2221 & ~n72408;
  assign n72410 = pi2221 & n72408;
  assign n72411 = ~n72409 & ~n72410;
  assign n72412 = pi7183 & pi9040;
  assign n72413 = pi7207 & ~pi9040;
  assign n72414 = ~n72412 & ~n72413;
  assign n72415 = ~pi2174 & n72414;
  assign n72416 = pi2174 & ~n72414;
  assign n72417 = ~n72415 & ~n72416;
  assign n72418 = ~n72411 & ~n72417;
  assign n72419 = pi7212 & pi9040;
  assign n72420 = pi7180 & ~pi9040;
  assign n72421 = ~n72419 & ~n72420;
  assign n72422 = ~pi2183 & n72421;
  assign n72423 = pi2183 & ~n72421;
  assign n72424 = ~n72422 & ~n72423;
  assign n72425 = pi7181 & ~pi9040;
  assign n72426 = pi7205 & pi9040;
  assign n72427 = ~n72425 & ~n72426;
  assign n72428 = pi2215 & n72427;
  assign n72429 = ~pi2215 & ~n72427;
  assign n72430 = ~n72428 & ~n72429;
  assign n72431 = ~n72424 & n72430;
  assign n72432 = n72418 & n72431;
  assign n72433 = n72405 & n72432;
  assign n72434 = n72424 & n72430;
  assign n72435 = n72411 & ~n72417;
  assign n72436 = n72434 & n72435;
  assign n72437 = n72411 & n72417;
  assign n72438 = n72405 & n72437;
  assign n72439 = n72430 & n72438;
  assign n72440 = ~n72424 & n72439;
  assign n72441 = n72405 & n72424;
  assign n72442 = n72417 & n72441;
  assign n72443 = ~n72411 & n72442;
  assign n72444 = ~n72440 & ~n72443;
  assign n72445 = ~n72436 & n72444;
  assign n72446 = ~n72433 & n72445;
  assign n72447 = ~n72405 & n72424;
  assign n72448 = ~n72417 & n72447;
  assign n72449 = n72411 & n72448;
  assign n72450 = n72446 & ~n72449;
  assign n72451 = ~n72399 & ~n72450;
  assign n72452 = n72405 & n72411;
  assign n72453 = ~n72417 & n72452;
  assign n72454 = ~n72424 & n72453;
  assign n72455 = ~n72442 & ~n72454;
  assign n72456 = ~n72405 & n72418;
  assign n72457 = ~n72424 & n72456;
  assign n72458 = n72455 & ~n72457;
  assign n72459 = ~n72430 & ~n72458;
  assign n72460 = ~n72405 & n72417;
  assign n72461 = n72411 & n72460;
  assign n72462 = ~n72430 & n72461;
  assign n72463 = ~n72424 & n72462;
  assign n72464 = ~n72411 & n72441;
  assign n72465 = ~n72411 & n72417;
  assign n72466 = n72424 & n72465;
  assign n72467 = ~n72464 & ~n72466;
  assign n72468 = ~n72430 & ~n72467;
  assign n72469 = ~n72463 & ~n72468;
  assign n72470 = ~n72399 & ~n72469;
  assign n72471 = ~n72459 & ~n72470;
  assign n72472 = ~n72451 & n72471;
  assign n72473 = ~n72405 & ~n72424;
  assign n72474 = n72430 & n72473;
  assign n72475 = n72465 & n72474;
  assign n72476 = ~n72405 & n72411;
  assign n72477 = n72434 & n72476;
  assign n72478 = n72424 & n72461;
  assign n72479 = n72405 & ~n72430;
  assign n72480 = n72411 & n72479;
  assign n72481 = ~n72411 & ~n72424;
  assign n72482 = ~n72405 & n72481;
  assign n72483 = ~n72480 & ~n72482;
  assign n72484 = ~n72478 & n72483;
  assign n72485 = ~n72456 & n72484;
  assign n72486 = n72418 & n72430;
  assign n72487 = n72424 & n72486;
  assign n72488 = ~n72424 & n72465;
  assign n72489 = ~n72405 & ~n72417;
  assign n72490 = ~n72488 & ~n72489;
  assign n72491 = n72430 & ~n72490;
  assign n72492 = ~n72487 & ~n72491;
  assign n72493 = n72485 & n72492;
  assign n72494 = n72399 & ~n72493;
  assign n72495 = ~n72477 & ~n72494;
  assign n72496 = ~n72475 & n72495;
  assign n72497 = n72472 & n72496;
  assign n72498 = pi2092 & n72497;
  assign n72499 = ~pi2092 & ~n72497;
  assign po2252 = n72498 | n72499;
  assign n72501 = n71950 & n71966;
  assign n72502 = ~n71996 & ~n72501;
  assign n72503 = ~n71938 & ~n72502;
  assign n72504 = n71957 & n71988;
  assign n72505 = ~n72102 & ~n72504;
  assign n72506 = n71938 & ~n72505;
  assign n72507 = ~n71957 & n71983;
  assign n72508 = ~n72122 & ~n72507;
  assign n72509 = ~n71965 & n72508;
  assign n72510 = ~n72506 & n72509;
  assign n72511 = ~n72503 & n72510;
  assign n72512 = ~n72098 & ~n72109;
  assign n72513 = n72511 & n72512;
  assign n72514 = n71975 & ~n72513;
  assign n72515 = n71951 & n72096;
  assign n72516 = n72005 & ~n72515;
  assign n72517 = n71938 & ~n72516;
  assign n72518 = ~n71957 & n71993;
  assign n72519 = ~n72517 & ~n72518;
  assign n72520 = n71944 & n71966;
  assign n72521 = n71957 & n71979;
  assign n72522 = ~n72520 & ~n72521;
  assign n72523 = n71938 & ~n72522;
  assign n72524 = n71938 & n71988;
  assign n72525 = ~n71957 & n72524;
  assign n72526 = ~n72523 & ~n72525;
  assign n72527 = n72519 & n72526;
  assign n72528 = ~n71975 & ~n72527;
  assign n72529 = ~n71983 & ~n71990;
  assign n72530 = ~n72103 & n72529;
  assign n72531 = n72010 & ~n72530;
  assign n72532 = ~n72528 & ~n72531;
  assign n72533 = ~n71965 & ~n72098;
  assign n72534 = ~n71938 & ~n72533;
  assign n72535 = n72532 & ~n72534;
  assign n72536 = ~n72514 & n72535;
  assign n72537 = ~pi2096 & n72536;
  assign n72538 = pi2096 & ~n72536;
  assign po2253 = n72537 | n72538;
  assign n72540 = pi7227 & pi9040;
  assign n72541 = pi7199 & ~pi9040;
  assign n72542 = ~n72540 & ~n72541;
  assign n72543 = ~pi2182 & n72542;
  assign n72544 = pi2182 & ~n72542;
  assign n72545 = ~n72543 & ~n72544;
  assign n72546 = pi7210 & pi9040;
  assign n72547 = pi7212 & ~pi9040;
  assign n72548 = ~n72546 & ~n72547;
  assign n72549 = pi2210 & n72548;
  assign n72550 = ~pi2210 & ~n72548;
  assign n72551 = ~n72549 & ~n72550;
  assign n72552 = pi7203 & pi9040;
  assign n72553 = pi7214 & ~pi9040;
  assign n72554 = ~n72552 & ~n72553;
  assign n72555 = pi2164 & n72554;
  assign n72556 = ~pi2164 & ~n72554;
  assign n72557 = ~n72555 & ~n72556;
  assign n72558 = ~n72551 & n72557;
  assign n72559 = ~n72545 & n72558;
  assign n72560 = pi7181 & pi9040;
  assign n72561 = pi7245 & ~pi9040;
  assign n72562 = ~n72560 & ~n72561;
  assign n72563 = pi2178 & n72562;
  assign n72564 = ~pi2178 & ~n72562;
  assign n72565 = ~n72563 & ~n72564;
  assign n72566 = n72545 & n72565;
  assign n72567 = ~n72557 & n72566;
  assign n72568 = ~n72545 & n72565;
  assign n72569 = n72557 & n72568;
  assign n72570 = ~n72567 & ~n72569;
  assign n72571 = ~n72559 & n72570;
  assign n72572 = pi7207 & pi9040;
  assign n72573 = pi7193 & ~pi9040;
  assign n72574 = ~n72572 & ~n72573;
  assign n72575 = ~pi2209 & n72574;
  assign n72576 = pi2209 & ~n72574;
  assign n72577 = ~n72575 & ~n72576;
  assign n72578 = pi7217 & pi9040;
  assign n72579 = pi7194 & ~pi9040;
  assign n72580 = ~n72578 & ~n72579;
  assign n72581 = ~pi2199 & n72580;
  assign n72582 = pi2199 & ~n72580;
  assign n72583 = ~n72581 & ~n72582;
  assign n72584 = n72577 & ~n72583;
  assign n72585 = ~n72571 & n72584;
  assign n72586 = n72545 & ~n72565;
  assign n72587 = n72557 & n72586;
  assign n72588 = ~n72583 & n72587;
  assign n72589 = n72551 & n72588;
  assign n72590 = ~n72545 & ~n72557;
  assign n72591 = ~n72545 & ~n72565;
  assign n72592 = n72551 & n72591;
  assign n72593 = ~n72590 & ~n72592;
  assign n72594 = ~n72577 & ~n72593;
  assign n72595 = n72557 & n72566;
  assign n72596 = ~n72577 & n72595;
  assign n72597 = ~n72594 & ~n72596;
  assign n72598 = ~n72583 & ~n72597;
  assign n72599 = ~n72589 & ~n72598;
  assign n72600 = n72551 & ~n72557;
  assign n72601 = ~n72545 & n72600;
  assign n72602 = ~n72551 & n72586;
  assign n72603 = ~n72557 & n72602;
  assign n72604 = ~n72601 & ~n72603;
  assign n72605 = ~n72577 & ~n72604;
  assign n72606 = n72599 & ~n72605;
  assign n72607 = n72551 & n72557;
  assign n72608 = n72545 & n72607;
  assign n72609 = n72565 & n72608;
  assign n72610 = n72551 & n72577;
  assign n72611 = n72591 & n72610;
  assign n72612 = n72557 & n72611;
  assign n72613 = ~n72568 & ~n72586;
  assign n72614 = n72600 & ~n72613;
  assign n72615 = ~n72612 & ~n72614;
  assign n72616 = ~n72609 & n72615;
  assign n72617 = n72558 & ~n72613;
  assign n72618 = ~n72551 & n72567;
  assign n72619 = ~n72617 & ~n72618;
  assign n72620 = ~n72551 & ~n72577;
  assign n72621 = n72557 & n72620;
  assign n72622 = ~n72565 & n72621;
  assign n72623 = ~n72557 & n72591;
  assign n72624 = n72577 & n72623;
  assign n72625 = ~n72551 & n72624;
  assign n72626 = ~n72622 & ~n72625;
  assign n72627 = n72619 & n72626;
  assign n72628 = n72616 & n72627;
  assign n72629 = n72583 & ~n72628;
  assign n72630 = n72606 & ~n72629;
  assign n72631 = ~n72585 & n72630;
  assign n72632 = ~pi2105 & ~n72631;
  assign n72633 = pi2105 & n72606;
  assign n72634 = ~n72585 & n72633;
  assign n72635 = ~n72629 & n72634;
  assign po2254 = n72632 | n72635;
  assign n72637 = ~n72557 & n72565;
  assign n72638 = n72577 & n72637;
  assign n72639 = n72551 & n72638;
  assign n72640 = ~n72602 & ~n72623;
  assign n72641 = ~n72569 & n72640;
  assign n72642 = n72577 & ~n72641;
  assign n72643 = n72557 & n72591;
  assign n72644 = ~n72557 & n72568;
  assign n72645 = ~n72643 & ~n72644;
  assign n72646 = ~n72577 & ~n72645;
  assign n72647 = ~n72642 & ~n72646;
  assign n72648 = ~n72596 & ~n72603;
  assign n72649 = n72647 & n72648;
  assign n72650 = n72583 & ~n72649;
  assign n72651 = n72551 & n72643;
  assign n72652 = ~n72551 & n72566;
  assign n72653 = n72551 & n72586;
  assign n72654 = ~n72652 & ~n72653;
  assign n72655 = n72577 & ~n72654;
  assign n72656 = ~n72651 & ~n72655;
  assign n72657 = ~n72577 & n72587;
  assign n72658 = n72570 & ~n72657;
  assign n72659 = ~n72623 & n72658;
  assign n72660 = ~n72551 & ~n72659;
  assign n72661 = n72656 & ~n72660;
  assign n72662 = ~n72583 & ~n72661;
  assign n72663 = ~n72650 & ~n72662;
  assign n72664 = ~n72639 & n72663;
  assign n72665 = ~n72557 & n72653;
  assign n72666 = ~n72609 & ~n72665;
  assign n72667 = ~n72577 & ~n72666;
  assign n72668 = n72664 & ~n72667;
  assign n72669 = ~pi2125 & ~n72668;
  assign n72670 = pi2125 & ~n72667;
  assign n72671 = n72663 & n72670;
  assign n72672 = ~n72639 & n72671;
  assign po2255 = n72669 | n72672;
  assign n72674 = n72405 & ~n72411;
  assign n72675 = ~n72449 & ~n72674;
  assign n72676 = ~n72481 & n72675;
  assign n72677 = n72430 & ~n72676;
  assign n72678 = ~n72424 & ~n72430;
  assign n72679 = n72411 & n72678;
  assign n72680 = n72405 & ~n72424;
  assign n72681 = ~n72417 & n72680;
  assign n72682 = n72424 & n72438;
  assign n72683 = ~n72681 & ~n72682;
  assign n72684 = ~n72405 & ~n72411;
  assign n72685 = n72424 & ~n72430;
  assign n72686 = n72684 & n72685;
  assign n72687 = n72683 & ~n72686;
  assign n72688 = ~n72679 & n72687;
  assign n72689 = ~n72677 & n72688;
  assign n72690 = n72399 & ~n72689;
  assign n72691 = n72405 & n72418;
  assign n72692 = n72424 & n72691;
  assign n72693 = n72405 & n72465;
  assign n72694 = ~n72424 & n72693;
  assign n72695 = ~n72692 & ~n72694;
  assign n72696 = n72430 & ~n72695;
  assign n72697 = ~n72690 & ~n72696;
  assign n72698 = ~n72424 & n72438;
  assign n72699 = ~n72453 & ~n72461;
  assign n72700 = n72430 & ~n72699;
  assign n72701 = ~n72698 & ~n72700;
  assign n72702 = ~n72457 & n72701;
  assign n72703 = ~n72399 & ~n72702;
  assign n72704 = ~n72435 & ~n72465;
  assign n72705 = ~n72405 & ~n72704;
  assign n72706 = ~n72466 & ~n72705;
  assign n72707 = ~n72430 & ~n72706;
  assign n72708 = ~n72399 & n72707;
  assign n72709 = ~n72703 & ~n72708;
  assign n72710 = n72697 & n72709;
  assign n72711 = pi2112 & ~n72710;
  assign n72712 = ~pi2112 & n72697;
  assign n72713 = n72709 & n72712;
  assign po2256 = n72711 | n72713;
  assign n72715 = ~n71504 & ~n72378;
  assign n72716 = ~n71423 & ~n72715;
  assign n72717 = ~n71488 & n71490;
  assign n72718 = n71423 & n72717;
  assign n72719 = ~n71435 & n72285;
  assign n72720 = ~n72368 & ~n72719;
  assign n72721 = ~n71459 & n72720;
  assign n72722 = ~n71423 & ~n72721;
  assign n72723 = ~n71449 & n71465;
  assign n72724 = ~n72722 & ~n72723;
  assign n72725 = ~n71488 & ~n72724;
  assign n72726 = ~n72718 & ~n72725;
  assign n72727 = ~n71453 & ~n71457;
  assign n72728 = ~n71449 & n71503;
  assign n72729 = ~n72348 & ~n72728;
  assign n72730 = n72727 & n72729;
  assign n72731 = n71423 & ~n72730;
  assign n72732 = ~n71429 & n71435;
  assign n72733 = n71423 & n72732;
  assign n72734 = n71449 & n72733;
  assign n72735 = ~n71449 & n72368;
  assign n72736 = ~n71457 & ~n72735;
  assign n72737 = ~n72375 & n72736;
  assign n72738 = ~n72734 & n72737;
  assign n72739 = ~n71423 & n72364;
  assign n72740 = n72738 & ~n72739;
  assign n72741 = n71488 & ~n72740;
  assign n72742 = ~n72731 & ~n72741;
  assign n72743 = n72726 & n72742;
  assign n72744 = ~n72716 & n72743;
  assign n72745 = pi2103 & n72744;
  assign n72746 = ~pi2103 & ~n72744;
  assign po2257 = n72745 | n72746;
  assign n72748 = ~n72424 & n72705;
  assign n72749 = ~n72460 & ~n72691;
  assign n72750 = ~n72430 & ~n72749;
  assign n72751 = ~n72748 & ~n72750;
  assign n72752 = n72417 & n72680;
  assign n72753 = ~n72489 & ~n72752;
  assign n72754 = ~n72693 & n72753;
  assign n72755 = n72430 & ~n72754;
  assign n72756 = n72751 & ~n72755;
  assign n72757 = n72424 & n72453;
  assign n72758 = n72756 & ~n72757;
  assign n72759 = ~n72399 & ~n72758;
  assign n72760 = n72434 & ~n72749;
  assign n72761 = ~n72456 & ~n72461;
  assign n72762 = ~n72453 & ~n72693;
  assign n72763 = n72761 & n72762;
  assign n72764 = ~n72424 & ~n72763;
  assign n72765 = ~n72760 & ~n72764;
  assign n72766 = ~n72682 & n72765;
  assign n72767 = n72399 & ~n72766;
  assign n72768 = ~n72759 & ~n72767;
  assign n72769 = ~n72424 & n72691;
  assign n72770 = ~n72757 & ~n72769;
  assign n72771 = ~n72430 & ~n72770;
  assign n72772 = n72768 & ~n72771;
  assign n72773 = pi2113 & ~n72772;
  assign n72774 = ~pi2113 & ~n72771;
  assign n72775 = ~n72767 & n72774;
  assign n72776 = ~n72759 & n72775;
  assign po2258 = n72773 | n72776;
  assign n72778 = n72199 & n72227;
  assign n72779 = ~n72246 & ~n72255;
  assign n72780 = n72205 & ~n72779;
  assign n72781 = ~n72778 & ~n72780;
  assign n72782 = ~n72241 & n72781;
  assign n72783 = ~n72205 & n72244;
  assign n72784 = ~n72233 & ~n72783;
  assign n72785 = ~n72263 & n72784;
  assign n72786 = n72782 & n72785;
  assign n72787 = n72180 & ~n72786;
  assign n72788 = n72213 & n72220;
  assign n72789 = n72199 & n72788;
  assign n72790 = ~n72218 & ~n72789;
  assign n72791 = ~n72199 & n72262;
  assign n72792 = ~n72228 & ~n72791;
  assign n72793 = n72193 & n72213;
  assign n72794 = n72205 & n72793;
  assign n72795 = n72199 & n72232;
  assign n72796 = ~n72794 & ~n72795;
  assign n72797 = n72192 & ~n72213;
  assign n72798 = ~n72186 & n72199;
  assign n72799 = ~n72797 & ~n72798;
  assign n72800 = ~n72268 & n72799;
  assign n72801 = ~n72205 & ~n72800;
  assign n72802 = n72796 & ~n72801;
  assign n72803 = n72792 & n72802;
  assign n72804 = n72790 & n72803;
  assign n72805 = ~n72180 & ~n72804;
  assign n72806 = ~n72787 & ~n72805;
  assign n72807 = pi2119 & ~n72806;
  assign n72808 = ~pi2119 & ~n72787;
  assign n72809 = ~n72805 & n72808;
  assign po2259 = n72807 | n72809;
  assign n72811 = ~n72577 & n72643;
  assign n72812 = ~n72551 & n72811;
  assign n72813 = n72566 & n72620;
  assign n72814 = ~n72557 & n72813;
  assign n72815 = ~n72812 & ~n72814;
  assign n72816 = ~n72618 & ~n72625;
  assign n72817 = n72557 & n72565;
  assign n72818 = n72551 & n72817;
  assign n72819 = ~n72592 & ~n72818;
  assign n72820 = ~n72577 & ~n72819;
  assign n72821 = ~n72551 & ~n72557;
  assign n72822 = n72577 & ~n72821;
  assign n72823 = ~n72613 & n72822;
  assign n72824 = ~n72551 & ~n72591;
  assign n72825 = ~n72577 & n72824;
  assign n72826 = ~n72557 & n72825;
  assign n72827 = ~n72823 & ~n72826;
  assign n72828 = ~n72820 & n72827;
  assign n72829 = n72816 & n72828;
  assign n72830 = ~n72583 & ~n72829;
  assign n72831 = n72815 & ~n72830;
  assign n72832 = n72569 & n72577;
  assign n72833 = n72551 & n72832;
  assign n72834 = n72577 & n72583;
  assign n72835 = ~n72592 & ~n72595;
  assign n72836 = ~n72613 & n72821;
  assign n72837 = n72835 & ~n72836;
  assign n72838 = n72834 & ~n72837;
  assign n72839 = n72551 & n72567;
  assign n72840 = n72551 & n72565;
  assign n72841 = ~n72557 & n72840;
  assign n72842 = ~n72653 & ~n72841;
  assign n72843 = ~n72551 & n72591;
  assign n72844 = ~n72587 & ~n72843;
  assign n72845 = n72842 & n72844;
  assign n72846 = ~n72577 & ~n72845;
  assign n72847 = ~n72839 & ~n72846;
  assign n72848 = n72583 & ~n72847;
  assign n72849 = ~n72838 & ~n72848;
  assign n72850 = ~n72833 & n72849;
  assign n72851 = n72831 & n72850;
  assign n72852 = pi2127 & ~n72851;
  assign n72853 = ~pi2127 & n72831;
  assign n72854 = n72850 & n72853;
  assign po2260 = n72852 | n72854;
  assign n72856 = ~n72568 & n72607;
  assign n72857 = ~n72583 & n72856;
  assign n72858 = n72568 & n72600;
  assign n72859 = ~n72577 & n72858;
  assign n72860 = n72557 & n72610;
  assign n72861 = n72545 & n72860;
  assign n72862 = ~n72859 & ~n72861;
  assign n72863 = ~n72857 & n72862;
  assign n72864 = ~n72653 & ~n72843;
  assign n72865 = ~n72577 & ~n72864;
  assign n72866 = ~n72814 & ~n72865;
  assign n72867 = ~n72583 & ~n72866;
  assign n72868 = ~n72568 & ~n72637;
  assign n72869 = ~n72551 & ~n72868;
  assign n72870 = ~n72643 & ~n72869;
  assign n72871 = n72577 & ~n72870;
  assign n72872 = ~n72836 & ~n72871;
  assign n72873 = n72551 & n72623;
  assign n72874 = n72545 & n72558;
  assign n72875 = n72551 & ~n72868;
  assign n72876 = ~n72874 & ~n72875;
  assign n72877 = ~n72577 & ~n72876;
  assign n72878 = ~n72873 & ~n72877;
  assign n72879 = n72872 & n72878;
  assign n72880 = n72583 & ~n72879;
  assign n72881 = ~n72587 & ~n72840;
  assign n72882 = n72584 & ~n72881;
  assign n72883 = ~n72880 & ~n72882;
  assign n72884 = ~n72867 & n72883;
  assign n72885 = n72863 & n72884;
  assign n72886 = ~pi2116 & n72885;
  assign n72887 = pi2116 & ~n72885;
  assign po2261 = n72886 | n72887;
  assign n72889 = n72424 & n72456;
  assign n72890 = ~n72682 & ~n72889;
  assign n72891 = ~n72430 & ~n72890;
  assign n72892 = n72453 & n72678;
  assign n72893 = ~n72891 & ~n72892;
  assign n72894 = ~n72477 & n72893;
  assign n72895 = n72405 & n72430;
  assign n72896 = n72417 & n72895;
  assign n72897 = ~n72411 & n72896;
  assign n72898 = n72424 & n72897;
  assign n72899 = n72430 & n72691;
  assign n72900 = ~n72449 & ~n72475;
  assign n72901 = ~n72440 & n72900;
  assign n72902 = ~n72899 & n72901;
  assign n72903 = n72399 & ~n72902;
  assign n72904 = ~n72424 & n72486;
  assign n72905 = ~n72897 & ~n72904;
  assign n72906 = ~n72681 & n72905;
  assign n72907 = n72417 & n72447;
  assign n72908 = ~n72424 & n72435;
  assign n72909 = ~n72452 & ~n72908;
  assign n72910 = ~n72430 & ~n72909;
  assign n72911 = ~n72907 & ~n72910;
  assign n72912 = n72906 & n72911;
  assign n72913 = ~n72399 & ~n72912;
  assign n72914 = ~n72424 & n72461;
  assign n72915 = ~n72456 & ~n72914;
  assign n72916 = ~n72693 & n72915;
  assign n72917 = ~n72430 & ~n72916;
  assign n72918 = n72399 & n72917;
  assign n72919 = ~n72913 & ~n72918;
  assign n72920 = ~n72903 & n72919;
  assign n72921 = ~n72898 & n72920;
  assign n72922 = n72894 & n72921;
  assign n72923 = pi2131 & ~n72922;
  assign n72924 = ~pi2131 & n72894;
  assign n72925 = n72921 & n72924;
  assign po2262 = n72923 | n72925;
  assign n72927 = ~n72199 & n72214;
  assign n72928 = ~n72788 & ~n72927;
  assign n72929 = n72205 & ~n72928;
  assign n72930 = ~n72263 & ~n72929;
  assign n72931 = n72199 & n72793;
  assign n72932 = ~n72235 & ~n72931;
  assign n72933 = n72199 & n72268;
  assign n72934 = ~n72797 & ~n72933;
  assign n72935 = n72213 & n72261;
  assign n72936 = n72934 & ~n72935;
  assign n72937 = ~n72205 & ~n72936;
  assign n72938 = ~n72199 & n72215;
  assign n72939 = ~n72937 & ~n72938;
  assign n72940 = n72932 & n72939;
  assign n72941 = n72930 & n72940;
  assign n72942 = ~n72180 & ~n72941;
  assign n72943 = n72199 & n72257;
  assign n72944 = ~n72249 & ~n72943;
  assign n72945 = ~n72205 & ~n72944;
  assign n72946 = ~n72942 & ~n72945;
  assign n72947 = n72205 & n72931;
  assign n72948 = ~n72193 & ~n72214;
  assign n72949 = n72239 & ~n72948;
  assign n72950 = ~n72262 & ~n72949;
  assign n72951 = ~n72789 & n72950;
  assign n72952 = ~n72205 & ~n72951;
  assign n72953 = n72199 & n72215;
  assign n72954 = ~n72952 & ~n72953;
  assign n72955 = n72199 & n72214;
  assign n72956 = ~n72199 & n72797;
  assign n72957 = ~n72935 & ~n72956;
  assign n72958 = ~n72955 & n72957;
  assign n72959 = n72205 & ~n72958;
  assign n72960 = n72954 & ~n72959;
  assign n72961 = n72180 & ~n72960;
  assign n72962 = ~n72947 & ~n72961;
  assign n72963 = n72946 & n72962;
  assign n72964 = pi2121 & n72963;
  assign n72965 = ~pi2121 & ~n72963;
  assign po2263 = n72964 | n72965;
  assign n72967 = ~n72199 & n72220;
  assign n72968 = ~n72791 & ~n72967;
  assign n72969 = n72205 & n72968;
  assign n72970 = ~n72213 & ~n72948;
  assign n72971 = n72186 & n72239;
  assign n72972 = ~n72955 & ~n72971;
  assign n72973 = ~n72970 & n72972;
  assign n72974 = ~n72205 & n72973;
  assign n72975 = ~n72943 & n72974;
  assign n72976 = ~n72969 & ~n72975;
  assign n72977 = n72199 & n72970;
  assign n72978 = ~n72789 & ~n72977;
  assign n72979 = ~n72976 & n72978;
  assign n72980 = n72180 & ~n72979;
  assign n72981 = n72205 & ~n72948;
  assign n72982 = ~n72199 & n72981;
  assign n72983 = ~n72234 & ~n72261;
  assign n72984 = n72199 & ~n72983;
  assign n72985 = n72205 & n72984;
  assign n72986 = n72213 & n72981;
  assign n72987 = ~n72985 & ~n72986;
  assign n72988 = ~n72982 & n72987;
  assign n72989 = ~n72180 & ~n72988;
  assign n72990 = ~n72980 & ~n72989;
  assign n72991 = ~n72205 & ~n72968;
  assign n72992 = ~n72218 & ~n72991;
  assign n72993 = ~n72180 & ~n72992;
  assign n72994 = n72205 & n72218;
  assign n72995 = ~n72205 & ~n72978;
  assign n72996 = ~n72994 & ~n72995;
  assign n72997 = ~n72993 & n72996;
  assign n72998 = n72990 & n72997;
  assign n72999 = pi2130 & ~n72998;
  assign n73000 = ~pi2130 & n72997;
  assign n73001 = ~n72989 & n73000;
  assign n73002 = ~n72980 & n73001;
  assign po2264 = n72999 | n73002;
  assign n73004 = ~n71957 & n71979;
  assign n73005 = ~n71978 & ~n73004;
  assign n73006 = ~n71938 & ~n73005;
  assign n73007 = n71938 & ~n72124;
  assign n73008 = ~n72113 & ~n73007;
  assign n73009 = ~n73006 & n73008;
  assign n73010 = n71975 & ~n73009;
  assign n73011 = ~n71938 & n71993;
  assign n73012 = ~n73010 & ~n73011;
  assign n73013 = ~n72507 & ~n72521;
  assign n73014 = n71938 & ~n73013;
  assign n73015 = n71938 & n71980;
  assign n73016 = n71957 & n71996;
  assign n73017 = ~n71938 & n71964;
  assign n73018 = ~n72101 & ~n73017;
  assign n73019 = ~n71944 & ~n73018;
  assign n73020 = ~n72102 & ~n73019;
  assign n73021 = ~n71965 & n73020;
  assign n73022 = ~n73016 & n73021;
  assign n73023 = ~n73015 & n73022;
  assign n73024 = ~n71975 & ~n73023;
  assign n73025 = ~n73014 & ~n73024;
  assign n73026 = n73012 & n73025;
  assign n73027 = pi2126 & ~n73026;
  assign n73028 = ~pi2126 & n73026;
  assign po2265 = n73027 | n73028;
  assign n73030 = pi4757 & pi9040;
  assign n73031 = pi4407 & ~pi9040;
  assign n73032 = ~n73030 & ~n73031;
  assign n73033 = ~pi2227 & n73032;
  assign n73034 = pi2227 & ~n73032;
  assign n73035 = ~n73033 & ~n73034;
  assign n73036 = pi4323 & pi9040;
  assign n73037 = pi4537 & ~pi9040;
  assign n73038 = ~n73036 & ~n73037;
  assign n73039 = pi2247 & ~n73038;
  assign n73040 = ~pi2247 & n73038;
  assign n73041 = ~n73039 & ~n73040;
  assign n73042 = pi4601 & pi9040;
  assign n73043 = pi4474 & ~pi9040;
  assign n73044 = ~n73042 & ~n73043;
  assign n73045 = pi2206 & n73044;
  assign n73046 = ~pi2206 & ~n73044;
  assign n73047 = ~n73045 & ~n73046;
  assign n73048 = pi4395 & pi9040;
  assign n73049 = pi4386 & ~pi9040;
  assign n73050 = ~n73048 & ~n73049;
  assign n73051 = ~pi2264 & n73050;
  assign n73052 = pi2264 & ~n73050;
  assign n73053 = ~n73051 & ~n73052;
  assign n73054 = pi4585 & pi9040;
  assign n73055 = pi4657 & ~pi9040;
  assign n73056 = ~n73054 & ~n73055;
  assign n73057 = ~pi2262 & n73056;
  assign n73058 = pi2262 & ~n73056;
  assign n73059 = ~n73057 & ~n73058;
  assign n73060 = n73053 & ~n73059;
  assign n73061 = ~n73047 & n73060;
  assign n73062 = pi4312 & pi9040;
  assign n73063 = pi4440 & ~pi9040;
  assign n73064 = ~n73062 & ~n73063;
  assign n73065 = pi2261 & n73064;
  assign n73066 = ~pi2261 & ~n73064;
  assign n73067 = ~n73065 & ~n73066;
  assign n73068 = ~n73053 & n73059;
  assign n73069 = ~n73047 & n73068;
  assign n73070 = ~n73067 & n73069;
  assign n73071 = n73047 & n73059;
  assign n73072 = n73067 & n73071;
  assign n73073 = ~n73070 & ~n73072;
  assign n73074 = n73047 & ~n73067;
  assign n73075 = ~n73059 & n73074;
  assign n73076 = ~n73053 & n73075;
  assign n73077 = n73073 & ~n73076;
  assign n73078 = ~n73061 & n73077;
  assign n73079 = ~n73041 & ~n73078;
  assign n73080 = n73053 & n73059;
  assign n73081 = n73047 & n73080;
  assign n73082 = ~n73067 & n73081;
  assign n73083 = ~n73079 & ~n73082;
  assign n73084 = ~n73047 & ~n73059;
  assign n73085 = ~n73053 & n73084;
  assign n73086 = n73067 & n73085;
  assign n73087 = n73083 & ~n73086;
  assign n73088 = ~n73047 & n73080;
  assign n73089 = n73053 & n73074;
  assign n73090 = ~n73053 & ~n73059;
  assign n73091 = n73067 & n73090;
  assign n73092 = ~n73089 & ~n73091;
  assign n73093 = ~n73088 & n73092;
  assign n73094 = n73041 & ~n73093;
  assign n73095 = n73087 & ~n73094;
  assign n73096 = n73035 & ~n73095;
  assign n73097 = n73047 & n73090;
  assign n73098 = ~n73041 & n73067;
  assign n73099 = n73097 & n73098;
  assign n73100 = n73047 & n73060;
  assign n73101 = ~n73041 & n73100;
  assign n73102 = ~n73041 & n73088;
  assign n73103 = ~n73101 & ~n73102;
  assign n73104 = ~n73067 & ~n73103;
  assign n73105 = ~n73067 & n73090;
  assign n73106 = n73060 & n73067;
  assign n73107 = ~n73105 & ~n73106;
  assign n73108 = ~n73053 & n73071;
  assign n73109 = ~n73061 & ~n73108;
  assign n73110 = n73107 & n73109;
  assign n73111 = n73041 & ~n73110;
  assign n73112 = ~n73067 & n73085;
  assign n73113 = ~n73111 & ~n73112;
  assign n73114 = ~n73067 & n73108;
  assign n73115 = n73067 & n73069;
  assign n73116 = ~n73114 & ~n73115;
  assign n73117 = n73113 & n73116;
  assign n73118 = ~n73104 & n73117;
  assign n73119 = ~n73099 & n73118;
  assign n73120 = ~n73035 & ~n73119;
  assign n73121 = n73061 & n73067;
  assign n73122 = n73067 & n73081;
  assign n73123 = ~n73121 & ~n73122;
  assign n73124 = ~n73041 & ~n73123;
  assign n73125 = ~n73120 & ~n73124;
  assign n73126 = n73067 & n73088;
  assign n73127 = ~n73114 & ~n73126;
  assign n73128 = n73041 & ~n73127;
  assign n73129 = n73125 & ~n73128;
  assign po2270 = ~n73096 & n73129;
  assign n73131 = n73061 & ~n73067;
  assign n73132 = n73067 & n73108;
  assign n73133 = ~n73126 & ~n73132;
  assign n73134 = ~n73131 & n73133;
  assign n73135 = n73041 & ~n73134;
  assign n73136 = ~n73085 & ~n73089;
  assign n73137 = ~n73041 & ~n73136;
  assign n73138 = ~n73075 & ~n73137;
  assign n73139 = n73067 & n73080;
  assign n73140 = ~n73047 & n73059;
  assign n73141 = ~n73067 & n73140;
  assign n73142 = ~n73139 & ~n73141;
  assign n73143 = ~n73047 & n73053;
  assign n73144 = ~n73097 & ~n73143;
  assign n73145 = n73142 & n73144;
  assign n73146 = n73041 & ~n73145;
  assign n73147 = ~n73132 & ~n73146;
  assign n73148 = n73138 & n73147;
  assign n73149 = ~n73035 & ~n73148;
  assign n73150 = ~n73135 & ~n73149;
  assign n73151 = ~n73047 & ~n73053;
  assign n73152 = ~n73041 & n73151;
  assign n73153 = n73067 & n73152;
  assign n73154 = n73067 & n73100;
  assign n73155 = n73041 & n73071;
  assign n73156 = ~n73067 & n73155;
  assign n73157 = ~n73154 & ~n73156;
  assign n73158 = n73047 & n73053;
  assign n73159 = n73067 & n73158;
  assign n73160 = ~n73069 & ~n73159;
  assign n73161 = ~n73041 & ~n73160;
  assign n73162 = ~n73041 & n73143;
  assign n73163 = ~n73067 & n73162;
  assign n73164 = ~n73161 & ~n73163;
  assign n73165 = n73157 & n73164;
  assign n73166 = n73035 & ~n73165;
  assign n73167 = ~n73153 & ~n73166;
  assign n73168 = ~n73076 & n73167;
  assign po2278 = ~n73150 | ~n73168;
  assign n73170 = pi4387 & pi9040;
  assign n73171 = pi4534 & ~pi9040;
  assign n73172 = ~n73170 & ~n73171;
  assign n73173 = pi2269 & n73172;
  assign n73174 = ~pi2269 & ~n73172;
  assign n73175 = ~n73173 & ~n73174;
  assign n73176 = pi4803 & pi9040;
  assign n73177 = pi4476 & ~pi9040;
  assign n73178 = ~n73176 & ~n73177;
  assign n73179 = ~pi2245 & ~n73178;
  assign n73180 = pi2245 & ~n73176;
  assign n73181 = ~n73177 & n73180;
  assign n73182 = ~n73179 & ~n73181;
  assign n73183 = pi4656 & pi9040;
  assign n73184 = pi4439 & ~pi9040;
  assign n73185 = ~n73183 & ~n73184;
  assign n73186 = ~pi2240 & n73185;
  assign n73187 = pi2240 & ~n73185;
  assign n73188 = ~n73186 & ~n73187;
  assign n73189 = pi4501 & pi9040;
  assign n73190 = pi4502 & ~pi9040;
  assign n73191 = ~n73189 & ~n73190;
  assign n73192 = ~pi2258 & n73191;
  assign n73193 = pi2258 & ~n73191;
  assign n73194 = ~n73192 & ~n73193;
  assign n73195 = pi4498 & pi9040;
  assign n73196 = pi4822 & ~pi9040;
  assign n73197 = ~n73195 & ~n73196;
  assign n73198 = pi2206 & n73197;
  assign n73199 = ~pi2206 & ~n73197;
  assign n73200 = ~n73198 & ~n73199;
  assign n73201 = n73194 & ~n73200;
  assign n73202 = n73188 & n73201;
  assign n73203 = ~n73182 & n73202;
  assign n73204 = ~n73194 & ~n73200;
  assign n73205 = n73188 & n73204;
  assign n73206 = n73182 & n73205;
  assign n73207 = ~n73203 & ~n73206;
  assign n73208 = ~n73175 & ~n73207;
  assign n73209 = ~n73182 & n73200;
  assign n73210 = ~n73188 & n73209;
  assign n73211 = n73194 & n73210;
  assign n73212 = n73175 & n73211;
  assign n73213 = pi4536 & ~pi9040;
  assign n73214 = pi4496 & pi9040;
  assign n73215 = ~n73213 & ~n73214;
  assign n73216 = ~pi2264 & ~n73215;
  assign n73217 = pi2264 & n73215;
  assign n73218 = ~n73216 & ~n73217;
  assign n73219 = ~n73188 & n73204;
  assign n73220 = ~n73175 & n73219;
  assign n73221 = ~n73211 & ~n73220;
  assign n73222 = ~n73182 & ~n73194;
  assign n73223 = n73188 & n73222;
  assign n73224 = ~n73182 & ~n73188;
  assign n73225 = n73194 & n73224;
  assign n73226 = ~n73223 & ~n73225;
  assign n73227 = n73175 & ~n73226;
  assign n73228 = n73175 & n73182;
  assign n73229 = n73201 & n73228;
  assign n73230 = n73188 & n73229;
  assign n73231 = n73182 & ~n73188;
  assign n73232 = n73200 & n73231;
  assign n73233 = ~n73194 & n73232;
  assign n73234 = n73194 & n73200;
  assign n73235 = n73188 & n73234;
  assign n73236 = ~n73175 & n73235;
  assign n73237 = ~n73233 & ~n73236;
  assign n73238 = ~n73230 & n73237;
  assign n73239 = ~n73227 & n73238;
  assign n73240 = n73221 & n73239;
  assign n73241 = n73218 & ~n73240;
  assign n73242 = ~n73182 & n73220;
  assign n73243 = ~n73241 & ~n73242;
  assign n73244 = ~n73212 & n73243;
  assign n73245 = ~n73208 & n73244;
  assign n73246 = ~n73188 & n73201;
  assign n73247 = n73182 & n73246;
  assign n73248 = ~n73203 & ~n73247;
  assign n73249 = ~n73175 & n73182;
  assign n73250 = ~n73188 & n73194;
  assign n73251 = n73249 & n73250;
  assign n73252 = ~n73175 & n73202;
  assign n73253 = n73182 & n73204;
  assign n73254 = n73188 & n73200;
  assign n73255 = ~n73253 & ~n73254;
  assign n73256 = n73175 & ~n73255;
  assign n73257 = ~n73194 & n73200;
  assign n73258 = ~n73188 & n73257;
  assign n73259 = ~n73175 & n73258;
  assign n73260 = n73188 & n73257;
  assign n73261 = ~n73182 & n73260;
  assign n73262 = ~n73259 & ~n73261;
  assign n73263 = ~n73256 & n73262;
  assign n73264 = ~n73252 & n73263;
  assign n73265 = ~n73251 & n73264;
  assign n73266 = n73248 & n73265;
  assign n73267 = ~n73218 & ~n73266;
  assign po2291 = n73245 & ~n73267;
  assign n73269 = pi4717 & pi9040;
  assign n73270 = pi4387 & ~pi9040;
  assign n73271 = ~n73269 & ~n73270;
  assign n73272 = ~pi2234 & ~n73271;
  assign n73273 = pi2234 & n73271;
  assign n73274 = ~n73272 & ~n73273;
  assign n73275 = pi4502 & pi9040;
  assign n73276 = pi4434 & ~pi9040;
  assign n73277 = ~n73275 & ~n73276;
  assign n73278 = ~pi2267 & n73277;
  assign n73279 = pi2267 & ~n73277;
  assign n73280 = ~n73278 & ~n73279;
  assign n73281 = pi4803 & ~pi9040;
  assign n73282 = pi4324 & pi9040;
  assign n73283 = ~n73281 & ~n73282;
  assign n73284 = ~pi2230 & n73283;
  assign n73285 = pi2230 & ~n73283;
  assign n73286 = ~n73284 & ~n73285;
  assign n73287 = pi4498 & ~pi9040;
  assign n73288 = pi4764 & pi9040;
  assign n73289 = ~n73287 & ~n73288;
  assign n73290 = ~pi2246 & n73289;
  assign n73291 = pi2246 & ~n73289;
  assign n73292 = ~n73290 & ~n73291;
  assign n73293 = pi4321 & pi9040;
  assign n73294 = pi4443 & ~pi9040;
  assign n73295 = ~n73293 & ~n73294;
  assign n73296 = ~pi2217 & ~n73295;
  assign n73297 = pi2217 & n73295;
  assign n73298 = ~n73296 & ~n73297;
  assign n73299 = ~n73292 & n73298;
  assign n73300 = ~n73286 & n73299;
  assign n73301 = n73280 & n73300;
  assign n73302 = ~n73292 & ~n73298;
  assign n73303 = n73286 & n73302;
  assign n73304 = n73280 & n73303;
  assign n73305 = ~n73301 & ~n73304;
  assign n73306 = pi4439 & pi9040;
  assign n73307 = pi4500 & ~pi9040;
  assign n73308 = ~n73306 & ~n73307;
  assign n73309 = pi2270 & n73308;
  assign n73310 = ~pi2270 & ~n73308;
  assign n73311 = ~n73309 & ~n73310;
  assign n73312 = ~n73286 & ~n73292;
  assign n73313 = ~n73311 & n73312;
  assign n73314 = n73280 & ~n73311;
  assign n73315 = ~n73286 & n73314;
  assign n73316 = ~n73313 & ~n73315;
  assign n73317 = n73305 & n73316;
  assign n73318 = ~n73280 & n73311;
  assign n73319 = n73292 & ~n73298;
  assign n73320 = n73286 & ~n73292;
  assign n73321 = n73298 & n73320;
  assign n73322 = ~n73319 & ~n73321;
  assign n73323 = n73318 & ~n73322;
  assign n73324 = n73311 & n73319;
  assign n73325 = n73286 & n73324;
  assign n73326 = ~n73323 & ~n73325;
  assign n73327 = n73317 & n73326;
  assign n73328 = n73274 & ~n73327;
  assign n73329 = n73292 & n73298;
  assign n73330 = ~n73286 & n73329;
  assign n73331 = ~n73280 & n73330;
  assign n73332 = n73286 & n73329;
  assign n73333 = n73280 & n73332;
  assign n73334 = ~n73331 & ~n73333;
  assign n73335 = n73311 & ~n73334;
  assign n73336 = ~n73328 & ~n73335;
  assign n73337 = n73286 & n73319;
  assign n73338 = ~n73280 & n73337;
  assign n73339 = ~n73311 & n73338;
  assign n73340 = n73280 & n73313;
  assign n73341 = ~n73339 & ~n73340;
  assign n73342 = ~n73280 & n73302;
  assign n73343 = ~n73280 & n73312;
  assign n73344 = ~n73342 & ~n73343;
  assign n73345 = ~n73332 & n73344;
  assign n73346 = n73311 & ~n73345;
  assign n73347 = n73280 & n73286;
  assign n73348 = n73311 & n73347;
  assign n73349 = n73298 & n73348;
  assign n73350 = ~n73286 & ~n73298;
  assign n73351 = ~n73332 & ~n73350;
  assign n73352 = n73280 & ~n73351;
  assign n73353 = ~n73311 & n73321;
  assign n73354 = ~n73280 & n73353;
  assign n73355 = ~n73352 & ~n73354;
  assign n73356 = ~n73349 & n73355;
  assign n73357 = ~n73346 & n73356;
  assign n73358 = ~n73331 & n73357;
  assign n73359 = ~n73274 & ~n73358;
  assign n73360 = n73341 & ~n73359;
  assign po2295 = ~n73336 | ~n73360;
  assign n73362 = ~n73194 & n73224;
  assign n73363 = ~n73203 & ~n73362;
  assign n73364 = n73182 & n73188;
  assign n73365 = ~n73194 & n73364;
  assign n73366 = ~n73205 & ~n73365;
  assign n73367 = ~n73175 & ~n73366;
  assign n73368 = ~n73175 & n73234;
  assign n73369 = ~n73182 & n73368;
  assign n73370 = ~n73367 & ~n73369;
  assign n73371 = n73175 & n73202;
  assign n73372 = n73175 & n73257;
  assign n73373 = ~n73182 & n73372;
  assign n73374 = ~n73371 & ~n73373;
  assign n73375 = n73370 & n73374;
  assign n73376 = ~n73247 & n73375;
  assign n73377 = n73363 & n73376;
  assign n73378 = ~n73218 & ~n73377;
  assign n73379 = n73182 & n73235;
  assign n73380 = ~n73233 & ~n73379;
  assign n73381 = ~n73211 & ~n73253;
  assign n73382 = ~n73205 & n73381;
  assign n73383 = n73175 & ~n73382;
  assign n73384 = ~n73175 & n73246;
  assign n73385 = ~n73383 & ~n73384;
  assign n73386 = ~n73175 & ~n73182;
  assign n73387 = n73260 & n73386;
  assign n73388 = n73385 & ~n73387;
  assign n73389 = n73380 & n73388;
  assign n73390 = n73218 & ~n73389;
  assign n73391 = ~n73242 & ~n73251;
  assign n73392 = ~n73203 & n73380;
  assign n73393 = n73175 & ~n73392;
  assign n73394 = n73391 & ~n73393;
  assign n73395 = ~n73390 & n73394;
  assign po2301 = n73378 | ~n73395;
  assign n73397 = n73280 & n73319;
  assign n73398 = ~n73330 & ~n73397;
  assign n73399 = ~n73274 & ~n73311;
  assign n73400 = ~n73398 & n73399;
  assign n73401 = ~n73286 & n73342;
  assign n73402 = ~n73321 & ~n73337;
  assign n73403 = ~n73280 & ~n73402;
  assign n73404 = ~n73401 & ~n73403;
  assign n73405 = ~n73274 & ~n73404;
  assign n73406 = n73311 & ~n73398;
  assign n73407 = n73280 & n73321;
  assign n73408 = ~n73406 & ~n73407;
  assign n73409 = ~n73280 & n73332;
  assign n73410 = n73408 & ~n73409;
  assign n73411 = ~n73286 & n73319;
  assign n73412 = ~n73280 & n73411;
  assign n73413 = ~n73300 & ~n73412;
  assign n73414 = ~n73303 & n73413;
  assign n73415 = ~n73311 & ~n73414;
  assign n73416 = ~n73292 & n73314;
  assign n73417 = ~n73415 & ~n73416;
  assign n73418 = n73410 & n73417;
  assign n73419 = n73274 & ~n73418;
  assign n73420 = ~n73280 & n73286;
  assign n73421 = n73292 & n73420;
  assign n73422 = ~n73401 & ~n73421;
  assign n73423 = n73311 & ~n73422;
  assign n73424 = ~n73419 & ~n73423;
  assign n73425 = ~n73274 & n73311;
  assign n73426 = n73280 & n73302;
  assign n73427 = ~n73312 & ~n73426;
  assign n73428 = ~n73332 & n73427;
  assign n73429 = n73425 & ~n73428;
  assign n73430 = n73424 & ~n73429;
  assign n73431 = ~n73405 & n73430;
  assign po2304 = n73400 | ~n73431;
  assign n73433 = n73067 & n73155;
  assign n73434 = n73041 & n73100;
  assign n73435 = ~n73067 & n73434;
  assign n73436 = ~n73433 & ~n73435;
  assign n73437 = n73041 & n73121;
  assign n73438 = n73041 & n73070;
  assign n73439 = ~n73089 & ~n73438;
  assign n73440 = n73060 & ~n73067;
  assign n73441 = ~n73100 & ~n73440;
  assign n73442 = ~n73085 & n73441;
  assign n73443 = ~n73041 & ~n73442;
  assign n73444 = n73041 & n73097;
  assign n73445 = ~n73443 & ~n73444;
  assign n73446 = n73439 & n73445;
  assign n73447 = n73133 & n73446;
  assign n73448 = n73035 & ~n73447;
  assign n73449 = ~n73041 & n73115;
  assign n73450 = ~n73448 & ~n73449;
  assign n73451 = ~n73053 & ~n73067;
  assign n73452 = ~n73041 & n73451;
  assign n73453 = ~n73067 & n73088;
  assign n73454 = ~n73085 & ~n73453;
  assign n73455 = n73041 & ~n73454;
  assign n73456 = ~n73452 & ~n73455;
  assign n73457 = n73123 & n73456;
  assign n73458 = ~n73035 & ~n73457;
  assign n73459 = n73450 & ~n73458;
  assign n73460 = ~n73437 & n73459;
  assign po2307 = ~n73436 | ~n73460;
  assign n73462 = ~n73086 & ~n73114;
  assign n73463 = ~n73453 & n73462;
  assign n73464 = ~n73041 & ~n73463;
  assign n73465 = ~n73437 & ~n73438;
  assign n73466 = ~n73108 & ~n73440;
  assign n73467 = n73041 & ~n73466;
  assign n73468 = ~n73084 & ~n73143;
  assign n73469 = n73067 & ~n73468;
  assign n73470 = ~n73059 & n73067;
  assign n73471 = ~n73080 & ~n73470;
  assign n73472 = ~n73085 & n73471;
  assign n73473 = ~n73041 & ~n73472;
  assign n73474 = ~n73469 & ~n73473;
  assign n73475 = ~n73467 & n73474;
  assign n73476 = n73035 & ~n73475;
  assign n73477 = ~n73076 & ~n73115;
  assign n73478 = ~n73081 & ~n73105;
  assign n73479 = n73041 & ~n73478;
  assign n73480 = n73477 & ~n73479;
  assign n73481 = ~n73101 & n73480;
  assign n73482 = ~n73035 & ~n73481;
  assign n73483 = ~n73476 & ~n73482;
  assign n73484 = n73465 & n73483;
  assign n73485 = ~n73464 & n73484;
  assign n73486 = pi2331 & n73485;
  assign n73487 = ~pi2331 & ~n73485;
  assign po2309 = n73486 | n73487;
  assign n73489 = pi4537 & pi9040;
  assign n73490 = pi4390 & ~pi9040;
  assign n73491 = ~n73489 & ~n73490;
  assign n73492 = pi2198 & n73491;
  assign n73493 = ~pi2198 & ~n73491;
  assign n73494 = ~n73492 & ~n73493;
  assign n73495 = pi4646 & ~pi9040;
  assign n73496 = pi4546 & pi9040;
  assign n73497 = ~n73495 & ~n73496;
  assign n73498 = pi2265 & n73497;
  assign n73499 = ~pi2265 & ~n73497;
  assign n73500 = ~n73498 & ~n73499;
  assign n73501 = pi4395 & ~pi9040;
  assign n73502 = pi4478 & pi9040;
  assign n73503 = ~n73501 & ~n73502;
  assign n73504 = ~pi2233 & n73503;
  assign n73505 = pi2233 & ~n73503;
  assign n73506 = ~n73504 & ~n73505;
  assign n73507 = pi4312 & ~pi9040;
  assign n73508 = pi4532 & pi9040;
  assign n73509 = ~n73507 & ~n73508;
  assign n73510 = ~pi2254 & ~n73509;
  assign n73511 = pi2254 & n73509;
  assign n73512 = ~n73510 & ~n73511;
  assign n73513 = pi4407 & pi9040;
  assign n73514 = pi4488 & ~pi9040;
  assign n73515 = ~n73513 & ~n73514;
  assign n73516 = pi2222 & n73515;
  assign n73517 = ~pi2222 & ~n73515;
  assign n73518 = ~n73516 & ~n73517;
  assign n73519 = n73512 & ~n73518;
  assign n73520 = n73506 & n73519;
  assign n73521 = n73500 & n73520;
  assign n73522 = ~n73512 & ~n73518;
  assign n73523 = ~n73506 & n73522;
  assign n73524 = n73500 & n73523;
  assign n73525 = n73506 & n73522;
  assign n73526 = ~n73500 & n73525;
  assign n73527 = ~n73524 & ~n73526;
  assign n73528 = ~n73521 & n73527;
  assign n73529 = ~n73500 & n73506;
  assign n73530 = n73518 & n73529;
  assign n73531 = n73512 & n73530;
  assign n73532 = n73528 & ~n73531;
  assign n73533 = ~n73494 & ~n73532;
  assign n73534 = ~n73512 & n73518;
  assign n73535 = ~n73506 & n73534;
  assign n73536 = ~n73500 & n73535;
  assign n73537 = n73506 & n73534;
  assign n73538 = n73500 & n73537;
  assign n73539 = ~n73520 & ~n73538;
  assign n73540 = ~n73494 & ~n73539;
  assign n73541 = ~n73506 & n73512;
  assign n73542 = n73518 & n73541;
  assign n73543 = n73500 & n73542;
  assign n73544 = ~n73540 & ~n73543;
  assign n73545 = n73494 & n73518;
  assign n73546 = ~n73500 & n73545;
  assign n73547 = n73500 & n73522;
  assign n73548 = ~n73541 & ~n73547;
  assign n73549 = n73494 & ~n73548;
  assign n73550 = ~n73546 & ~n73549;
  assign n73551 = n73544 & n73550;
  assign n73552 = ~n73536 & n73551;
  assign n73553 = pi4662 & pi9040;
  assign n73554 = pi4706 & ~pi9040;
  assign n73555 = ~n73553 & ~n73554;
  assign n73556 = ~pi2271 & ~n73555;
  assign n73557 = pi2271 & n73555;
  assign n73558 = ~n73556 & ~n73557;
  assign n73559 = ~n73552 & ~n73558;
  assign n73560 = ~n73533 & ~n73559;
  assign n73561 = ~n73506 & n73519;
  assign n73562 = n73500 & n73561;
  assign n73563 = ~n73518 & n73529;
  assign n73564 = n73494 & ~n73563;
  assign n73565 = n73500 & ~n73506;
  assign n73566 = ~n73512 & n73565;
  assign n73567 = n73512 & n73518;
  assign n73568 = n73506 & n73518;
  assign n73569 = ~n73567 & ~n73568;
  assign n73570 = ~n73500 & ~n73569;
  assign n73571 = ~n73566 & ~n73570;
  assign n73572 = ~n73494 & n73571;
  assign n73573 = ~n73523 & n73572;
  assign n73574 = ~n73564 & ~n73573;
  assign n73575 = ~n73562 & ~n73574;
  assign n73576 = n73494 & n73500;
  assign n73577 = n73568 & n73576;
  assign n73578 = n73575 & ~n73577;
  assign n73579 = n73558 & ~n73578;
  assign n73580 = n73494 & n73536;
  assign n73581 = ~n73579 & ~n73580;
  assign n73582 = n73560 & n73581;
  assign n73583 = ~pi2272 & n73582;
  assign n73584 = pi2272 & ~n73582;
  assign po2310 = n73583 | n73584;
  assign n73586 = n73219 & n73228;
  assign n73587 = ~n73230 & ~n73586;
  assign n73588 = ~n73223 & ~n73254;
  assign n73589 = ~n73175 & ~n73588;
  assign n73590 = n73218 & n73589;
  assign n73591 = ~n73182 & n73204;
  assign n73592 = ~n73260 & ~n73591;
  assign n73593 = n73175 & ~n73592;
  assign n73594 = ~n73182 & n73201;
  assign n73595 = ~n73206 & ~n73594;
  assign n73596 = ~n73175 & ~n73595;
  assign n73597 = ~n73182 & n73219;
  assign n73598 = ~n73596 & ~n73597;
  assign n73599 = ~n73211 & ~n73233;
  assign n73600 = n73598 & n73599;
  assign n73601 = ~n73593 & n73600;
  assign n73602 = ~n73218 & ~n73601;
  assign n73603 = ~n73233 & ~n73247;
  assign n73604 = ~n73379 & n73603;
  assign n73605 = ~n73175 & ~n73604;
  assign n73606 = ~n73602 & ~n73605;
  assign n73607 = n73194 & n73364;
  assign n73608 = n73182 & n73219;
  assign n73609 = ~n73607 & ~n73608;
  assign n73610 = n73218 & ~n73609;
  assign n73611 = n73200 & n73224;
  assign n73612 = ~n73225 & ~n73611;
  assign n73613 = ~n73188 & n73234;
  assign n73614 = n73612 & ~n73613;
  assign n73615 = n73175 & ~n73614;
  assign n73616 = n73218 & n73615;
  assign n73617 = ~n73610 & ~n73616;
  assign n73618 = n73606 & n73617;
  assign n73619 = ~n73590 & n73618;
  assign po2312 = ~n73587 | ~n73619;
  assign n73621 = pi4546 & ~pi9040;
  assign n73622 = pi4474 & pi9040;
  assign n73623 = ~n73621 & ~n73622;
  assign n73624 = pi2268 & n73623;
  assign n73625 = ~pi2268 & ~n73623;
  assign n73626 = ~n73624 & ~n73625;
  assign n73627 = pi4596 & ~pi9040;
  assign n73628 = pi4488 & pi9040;
  assign n73629 = ~n73627 & ~n73628;
  assign n73630 = pi2216 & ~n73629;
  assign n73631 = ~pi2216 & n73629;
  assign n73632 = ~n73630 & ~n73631;
  assign n73633 = ~n73626 & n73632;
  assign n73634 = pi4386 & pi9040;
  assign n73635 = pi4320 & ~pi9040;
  assign n73636 = ~n73634 & ~n73635;
  assign n73637 = pi2262 & n73636;
  assign n73638 = ~pi2262 & ~n73636;
  assign n73639 = ~n73637 & ~n73638;
  assign n73640 = pi4757 & ~pi9040;
  assign n73641 = pi4720 & pi9040;
  assign n73642 = ~n73640 & ~n73641;
  assign n73643 = ~pi2241 & n73642;
  assign n73644 = pi2241 & ~n73642;
  assign n73645 = ~n73643 & ~n73644;
  assign n73646 = n73639 & ~n73645;
  assign n73647 = n73633 & n73646;
  assign n73648 = pi4440 & pi9040;
  assign n73649 = pi4662 & ~pi9040;
  assign n73650 = ~n73648 & ~n73649;
  assign n73651 = pi2227 & n73650;
  assign n73652 = ~pi2227 & ~n73650;
  assign n73653 = ~n73651 & ~n73652;
  assign n73654 = n73645 & n73653;
  assign n73655 = ~n73639 & n73654;
  assign n73656 = ~n73626 & n73655;
  assign n73657 = ~n73639 & n73653;
  assign n73658 = ~n73645 & n73657;
  assign n73659 = n73626 & n73658;
  assign n73660 = n73626 & ~n73639;
  assign n73661 = n73645 & n73660;
  assign n73662 = ~n73653 & n73661;
  assign n73663 = ~n73659 & ~n73662;
  assign n73664 = ~n73626 & ~n73632;
  assign n73665 = n73654 & n73664;
  assign n73666 = ~n73645 & ~n73653;
  assign n73667 = n73639 & n73666;
  assign n73668 = n73639 & ~n73653;
  assign n73669 = ~n73626 & n73668;
  assign n73670 = ~n73667 & ~n73669;
  assign n73671 = n73626 & n73639;
  assign n73672 = n73645 & n73671;
  assign n73673 = n73653 & n73672;
  assign n73674 = n73670 & ~n73673;
  assign n73675 = n73632 & ~n73674;
  assign n73676 = ~n73645 & n73653;
  assign n73677 = n73645 & ~n73653;
  assign n73678 = ~n73676 & ~n73677;
  assign n73679 = n73626 & ~n73678;
  assign n73680 = ~n73639 & n73677;
  assign n73681 = ~n73679 & ~n73680;
  assign n73682 = ~n73632 & ~n73681;
  assign n73683 = ~n73675 & ~n73682;
  assign n73684 = ~n73639 & n73666;
  assign n73685 = ~n73626 & n73684;
  assign n73686 = n73683 & ~n73685;
  assign n73687 = ~n73665 & n73686;
  assign n73688 = n73663 & n73687;
  assign n73689 = pi4532 & ~pi9040;
  assign n73690 = pi4597 & pi9040;
  assign n73691 = ~n73689 & ~n73690;
  assign n73692 = ~pi2266 & ~n73691;
  assign n73693 = pi2266 & n73691;
  assign n73694 = ~n73692 & ~n73693;
  assign n73695 = ~n73688 & n73694;
  assign n73696 = ~n73626 & n73645;
  assign n73697 = ~n73639 & n73696;
  assign n73698 = n73639 & n73677;
  assign n73699 = n73626 & n73698;
  assign n73700 = ~n73697 & ~n73699;
  assign n73701 = n73639 & n73676;
  assign n73702 = ~n73655 & ~n73701;
  assign n73703 = n73700 & n73702;
  assign n73704 = n73632 & ~n73703;
  assign n73705 = n73626 & n73684;
  assign n73706 = ~n73704 & ~n73705;
  assign n73707 = ~n73694 & ~n73706;
  assign n73708 = ~n73632 & ~n73694;
  assign n73709 = ~n73626 & n73676;
  assign n73710 = ~n73673 & ~n73709;
  assign n73711 = ~n73669 & n73710;
  assign n73712 = n73708 & ~n73711;
  assign n73713 = ~n73707 & ~n73712;
  assign n73714 = ~n73695 & n73713;
  assign n73715 = ~n73656 & n73714;
  assign po2317 = n73647 | ~n73715;
  assign n73717 = n73626 & n73701;
  assign n73718 = ~n73632 & n73667;
  assign n73719 = ~n73717 & ~n73718;
  assign n73720 = n73626 & n73653;
  assign n73721 = ~n73657 & ~n73720;
  assign n73722 = ~n73698 & n73721;
  assign n73723 = n73632 & ~n73722;
  assign n73724 = n73719 & ~n73723;
  assign n73725 = ~n73632 & n73680;
  assign n73726 = n73724 & ~n73725;
  assign n73727 = ~n73694 & ~n73726;
  assign n73728 = ~n73626 & n73653;
  assign n73729 = n73639 & n73728;
  assign n73730 = n73632 & n73729;
  assign n73731 = ~n73653 & n73671;
  assign n73732 = ~n73645 & n73731;
  assign n73733 = ~n73632 & n73657;
  assign n73734 = ~n73662 & ~n73733;
  assign n73735 = ~n73732 & n73734;
  assign n73736 = ~n73730 & n73735;
  assign n73737 = n73632 & n73684;
  assign n73738 = ~n73626 & n73639;
  assign n73739 = n73645 & n73738;
  assign n73740 = ~n73685 & ~n73739;
  assign n73741 = ~n73737 & n73740;
  assign n73742 = n73736 & n73741;
  assign n73743 = n73694 & ~n73742;
  assign n73744 = n73632 & n73685;
  assign n73745 = n73639 & n73654;
  assign n73746 = ~n73626 & n73745;
  assign n73747 = ~n73632 & n73746;
  assign n73748 = ~n73744 & ~n73747;
  assign n73749 = ~n73626 & n73658;
  assign n73750 = ~n73632 & n73749;
  assign n73751 = n73748 & ~n73750;
  assign n73752 = ~n73743 & n73751;
  assign po2320 = n73727 | ~n73752;
  assign n73754 = pi4496 & ~pi9040;
  assign n73755 = pi4434 & pi9040;
  assign n73756 = ~n73754 & ~n73755;
  assign n73757 = pi2271 & n73756;
  assign n73758 = ~pi2271 & ~n73756;
  assign n73759 = ~n73757 & ~n73758;
  assign n73760 = pi4504 & ~pi9040;
  assign n73761 = pi4500 & pi9040;
  assign n73762 = ~n73760 & ~n73761;
  assign n73763 = ~pi2230 & ~n73762;
  assign n73764 = pi2230 & n73762;
  assign n73765 = ~n73763 & ~n73764;
  assign n73766 = ~n73759 & ~n73765;
  assign n73767 = pi4804 & ~pi9040;
  assign n73768 = pi4445 & pi9040;
  assign n73769 = ~n73767 & ~n73768;
  assign n73770 = ~pi2255 & n73769;
  assign n73771 = pi2255 & ~n73769;
  assign n73772 = ~n73770 & ~n73771;
  assign n73773 = pi4729 & pi9040;
  assign n73774 = pi4321 & ~pi9040;
  assign n73775 = ~n73773 & ~n73774;
  assign n73776 = ~pi2223 & ~n73775;
  assign n73777 = pi2223 & n73775;
  assign n73778 = ~n73776 & ~n73777;
  assign n73779 = pi4501 & ~pi9040;
  assign n73780 = pi4487 & pi9040;
  assign n73781 = ~n73779 & ~n73780;
  assign n73782 = ~pi2254 & ~n73781;
  assign n73783 = pi2254 & n73781;
  assign n73784 = ~n73782 & ~n73783;
  assign n73785 = n73778 & ~n73784;
  assign n73786 = ~n73772 & n73785;
  assign n73787 = n73766 & n73786;
  assign n73788 = pi4822 & pi9040;
  assign n73789 = pi4324 & ~pi9040;
  assign n73790 = ~n73788 & ~n73789;
  assign n73791 = ~pi2246 & n73790;
  assign n73792 = pi2246 & ~n73790;
  assign n73793 = ~n73791 & ~n73792;
  assign n73794 = ~n73759 & n73765;
  assign n73795 = ~n73772 & n73778;
  assign n73796 = n73794 & n73795;
  assign n73797 = n73784 & n73796;
  assign n73798 = ~n73772 & ~n73778;
  assign n73799 = n73759 & n73765;
  assign n73800 = n73798 & n73799;
  assign n73801 = ~n73778 & n73784;
  assign n73802 = ~n73765 & n73801;
  assign n73803 = ~n73759 & n73802;
  assign n73804 = n73759 & ~n73765;
  assign n73805 = n73784 & n73804;
  assign n73806 = ~n73772 & n73805;
  assign n73807 = n73778 & n73806;
  assign n73808 = ~n73803 & ~n73807;
  assign n73809 = ~n73800 & n73808;
  assign n73810 = ~n73797 & n73809;
  assign n73811 = ~n73778 & ~n73784;
  assign n73812 = n73765 & n73811;
  assign n73813 = n73759 & n73812;
  assign n73814 = n73810 & ~n73813;
  assign n73815 = n73793 & ~n73814;
  assign n73816 = ~n73784 & n73804;
  assign n73817 = n73772 & n73816;
  assign n73818 = n73778 & n73817;
  assign n73819 = ~n73759 & n73801;
  assign n73820 = n73766 & ~n73778;
  assign n73821 = ~n73819 & ~n73820;
  assign n73822 = n73772 & ~n73821;
  assign n73823 = ~n73818 & ~n73822;
  assign n73824 = n73793 & ~n73823;
  assign n73825 = n73759 & n73784;
  assign n73826 = n73765 & n73825;
  assign n73827 = n73778 & n73826;
  assign n73828 = ~n73802 & ~n73827;
  assign n73829 = ~n73784 & n73794;
  assign n73830 = n73778 & n73829;
  assign n73831 = n73828 & ~n73830;
  assign n73832 = n73772 & ~n73831;
  assign n73833 = ~n73824 & ~n73832;
  assign n73834 = ~n73815 & n73833;
  assign n73835 = ~n73787 & n73834;
  assign n73836 = ~n73784 & n73798;
  assign n73837 = n73759 & n73836;
  assign n73838 = ~n73759 & n73778;
  assign n73839 = ~n73784 & n73838;
  assign n73840 = n73772 & n73784;
  assign n73841 = n73759 & n73840;
  assign n73842 = ~n73839 & ~n73841;
  assign n73843 = ~n73772 & n73794;
  assign n73844 = ~n73778 & n73843;
  assign n73845 = n73765 & ~n73784;
  assign n73846 = n73766 & n73778;
  assign n73847 = ~n73845 & ~n73846;
  assign n73848 = ~n73772 & ~n73847;
  assign n73849 = ~n73844 & ~n73848;
  assign n73850 = ~n73778 & n73816;
  assign n73851 = n73849 & ~n73850;
  assign n73852 = ~n73829 & n73851;
  assign n73853 = n73842 & n73852;
  assign n73854 = ~n73793 & ~n73853;
  assign n73855 = ~n73837 & ~n73854;
  assign po2325 = n73835 & n73855;
  assign n73857 = pi4596 & pi9040;
  assign n73858 = pi4389 & ~pi9040;
  assign n73859 = ~n73857 & ~n73858;
  assign n73860 = ~pi2266 & ~n73859;
  assign n73861 = pi2266 & n73859;
  assign n73862 = ~n73860 & ~n73861;
  assign n73863 = pi4601 & ~pi9040;
  assign n73864 = pi4388 & pi9040;
  assign n73865 = ~n73863 & ~n73864;
  assign n73866 = ~pi2233 & n73865;
  assign n73867 = pi2233 & ~n73865;
  assign n73868 = ~n73866 & ~n73867;
  assign n73869 = pi4646 & pi9040;
  assign n73870 = pi4720 & ~pi9040;
  assign n73871 = ~n73869 & ~n73870;
  assign n73872 = ~pi2241 & n73871;
  assign n73873 = pi2241 & ~n73871;
  assign n73874 = ~n73872 & ~n73873;
  assign n73875 = pi4320 & pi9040;
  assign n73876 = pi4499 & ~pi9040;
  assign n73877 = ~n73875 & ~n73876;
  assign n73878 = ~pi2252 & ~n73877;
  assign n73879 = pi2252 & n73877;
  assign n73880 = ~n73878 & ~n73879;
  assign n73881 = n73874 & n73880;
  assign n73882 = ~n73868 & n73881;
  assign n73883 = ~n73862 & n73882;
  assign n73884 = n73862 & n73868;
  assign n73885 = n73874 & n73884;
  assign n73886 = ~n73862 & n73868;
  assign n73887 = ~n73874 & n73886;
  assign n73888 = n73880 & n73887;
  assign n73889 = ~n73885 & ~n73888;
  assign n73890 = ~n73883 & n73889;
  assign n73891 = pi4706 & pi9040;
  assign n73892 = pi4585 & ~pi9040;
  assign n73893 = ~n73891 & ~n73892;
  assign n73894 = pi2263 & n73893;
  assign n73895 = ~pi2263 & ~n73893;
  assign n73896 = ~n73894 & ~n73895;
  assign n73897 = ~n73890 & ~n73896;
  assign n73898 = ~n73862 & ~n73874;
  assign n73899 = ~n73880 & n73898;
  assign n73900 = n73862 & ~n73874;
  assign n73901 = n73880 & n73900;
  assign n73902 = ~n73899 & ~n73901;
  assign n73903 = n73896 & ~n73902;
  assign n73904 = ~n73897 & ~n73903;
  assign n73905 = pi4597 & ~pi9040;
  assign n73906 = ~pi4423 & pi9040;
  assign n73907 = ~n73905 & ~n73906;
  assign n73908 = ~pi2222 & ~n73907;
  assign n73909 = pi2222 & n73907;
  assign n73910 = ~n73908 & ~n73909;
  assign n73911 = n73874 & n73886;
  assign n73912 = ~n73880 & n73911;
  assign n73913 = ~n73883 & ~n73912;
  assign n73914 = n73862 & n73874;
  assign n73915 = n73880 & n73914;
  assign n73916 = n73862 & ~n73868;
  assign n73917 = ~n73874 & n73916;
  assign n73918 = ~n73880 & n73917;
  assign n73919 = ~n73915 & ~n73918;
  assign n73920 = ~n73896 & ~n73919;
  assign n73921 = ~n73862 & ~n73868;
  assign n73922 = ~n73874 & n73921;
  assign n73923 = n73874 & n73916;
  assign n73924 = ~n73880 & n73923;
  assign n73925 = ~n73922 & ~n73924;
  assign n73926 = n73896 & ~n73925;
  assign n73927 = ~n73920 & ~n73926;
  assign n73928 = n73913 & n73927;
  assign n73929 = n73910 & ~n73928;
  assign n73930 = n73868 & n73874;
  assign n73931 = ~n73896 & n73930;
  assign n73932 = ~n73880 & n73931;
  assign n73933 = n73896 & n73921;
  assign n73934 = ~n73880 & n73933;
  assign n73935 = n73880 & n73911;
  assign n73936 = ~n73874 & n73884;
  assign n73937 = ~n73935 & ~n73936;
  assign n73938 = n73880 & n73916;
  assign n73939 = n73937 & ~n73938;
  assign n73940 = n73896 & ~n73939;
  assign n73941 = ~n73880 & ~n73896;
  assign n73942 = n73914 & n73941;
  assign n73943 = ~n73880 & n73885;
  assign n73944 = ~n73942 & ~n73943;
  assign n73945 = ~n73940 & n73944;
  assign n73946 = ~n73934 & n73945;
  assign n73947 = ~n73880 & n73922;
  assign n73948 = n73880 & n73917;
  assign n73949 = ~n73947 & ~n73948;
  assign n73950 = n73946 & n73949;
  assign n73951 = ~n73910 & ~n73950;
  assign n73952 = ~n73932 & ~n73951;
  assign n73953 = ~n73929 & n73952;
  assign po2327 = n73904 & n73953;
  assign n73955 = ~n73626 & n73698;
  assign n73956 = n73632 & n73676;
  assign n73957 = ~n73626 & n73956;
  assign n73958 = ~n73955 & ~n73957;
  assign n73959 = n73626 & n73646;
  assign n73960 = ~n73626 & ~n73653;
  assign n73961 = ~n73739 & ~n73960;
  assign n73962 = ~n73632 & ~n73961;
  assign n73963 = ~n73959 & ~n73962;
  assign n73964 = n73958 & n73963;
  assign n73965 = n73694 & ~n73964;
  assign n73966 = n73664 & n73676;
  assign n73967 = ~n73626 & n73666;
  assign n73968 = ~n73659 & ~n73967;
  assign n73969 = ~n73745 & n73968;
  assign n73970 = n73632 & ~n73969;
  assign n73971 = ~n73698 & ~n73705;
  assign n73972 = ~n73632 & ~n73971;
  assign n73973 = ~n73656 & ~n73972;
  assign n73974 = ~n73970 & n73973;
  assign n73975 = ~n73966 & n73974;
  assign n73976 = ~n73694 & ~n73975;
  assign n73977 = ~n73965 & ~n73976;
  assign n73978 = n73626 & n73702;
  assign n73979 = ~n73626 & ~n73677;
  assign n73980 = ~n73978 & ~n73979;
  assign n73981 = ~n73632 & n73980;
  assign n73982 = n73626 & n73632;
  assign n73983 = ~n73680 & ~n73745;
  assign n73984 = ~n73667 & n73983;
  assign n73985 = n73982 & ~n73984;
  assign n73986 = ~n73981 & ~n73985;
  assign po2331 = n73977 & n73986;
  assign n73988 = ~n73311 & ~n73402;
  assign n73989 = ~n73292 & n73420;
  assign n73990 = ~n73280 & n73299;
  assign n73991 = ~n73989 & ~n73990;
  assign n73992 = ~n73311 & ~n73991;
  assign n73993 = ~n73311 & n73329;
  assign n73994 = n73280 & n73993;
  assign n73995 = ~n73992 & ~n73994;
  assign n73996 = n73280 & n73330;
  assign n73997 = n73302 & ~n73311;
  assign n73998 = n73280 & n73997;
  assign n73999 = ~n73286 & n73998;
  assign n74000 = ~n73996 & ~n73999;
  assign n74001 = n73995 & n74000;
  assign n74002 = ~n73988 & n74001;
  assign n74003 = ~n73274 & ~n74002;
  assign n74004 = ~n73304 & ~n73409;
  assign n74005 = ~n73411 & n74004;
  assign n74006 = n73425 & ~n74005;
  assign n74007 = ~n74003 & ~n74006;
  assign n74008 = ~n73301 & ~n73401;
  assign n74009 = n73280 & n73411;
  assign n74010 = ~n73280 & n73329;
  assign n74011 = n73280 & ~n73298;
  assign n74012 = n73286 & n74011;
  assign n74013 = ~n74010 & ~n74012;
  assign n74014 = ~n73311 & ~n74013;
  assign n74015 = ~n73298 & n73420;
  assign n74016 = ~n73321 & ~n74015;
  assign n74017 = n73311 & ~n74016;
  assign n74018 = ~n74014 & ~n74017;
  assign n74019 = ~n73349 & n74018;
  assign n74020 = ~n74009 & n74019;
  assign n74021 = ~n73331 & n74020;
  assign n74022 = n74008 & n74021;
  assign n74023 = n73274 & ~n74022;
  assign n74024 = n73311 & ~n74008;
  assign n74025 = ~n74023 & ~n74024;
  assign po2335 = ~n74007 | ~n74025;
  assign n74027 = ~n73494 & n73563;
  assign n74028 = ~n73500 & n73520;
  assign n74029 = n73506 & n73567;
  assign n74030 = n73500 & n74029;
  assign n74031 = ~n73500 & n73534;
  assign n74032 = ~n74030 & ~n74031;
  assign n74033 = n73494 & ~n74032;
  assign n74034 = ~n73525 & ~n73535;
  assign n74035 = n73500 & ~n74034;
  assign n74036 = ~n73518 & n73541;
  assign n74037 = ~n73506 & n73518;
  assign n74038 = n73500 & n74037;
  assign n74039 = n73512 & n73529;
  assign n74040 = ~n74038 & ~n74039;
  assign n74041 = ~n74036 & n74040;
  assign n74042 = ~n73494 & ~n74041;
  assign n74043 = ~n74035 & ~n74042;
  assign n74044 = ~n74033 & n74043;
  assign n74045 = ~n74028 & n74044;
  assign n74046 = n73558 & ~n74045;
  assign n74047 = ~n74027 & ~n74046;
  assign n74048 = ~n73526 & ~n73538;
  assign n74049 = n73519 & n73576;
  assign n74050 = n73494 & n73567;
  assign n74051 = ~n73500 & n74050;
  assign n74052 = ~n74049 & ~n74051;
  assign n74053 = n73494 & n73523;
  assign n74054 = n74052 & ~n74053;
  assign n74055 = ~n73500 & n73542;
  assign n74056 = n73500 & n73568;
  assign n74057 = ~n73535 & ~n74056;
  assign n74058 = ~n73494 & ~n74057;
  assign n74059 = ~n74055 & ~n74058;
  assign n74060 = ~n73518 & n73565;
  assign n74061 = n74059 & ~n74060;
  assign n74062 = n74054 & n74061;
  assign n74063 = n74048 & n74062;
  assign n74064 = ~n73558 & ~n74063;
  assign n74065 = n73494 & ~n73500;
  assign n74066 = n73542 & n74065;
  assign n74067 = ~n74064 & ~n74066;
  assign po2337 = n74047 & n74067;
  assign n74069 = ~n73188 & n73249;
  assign n74070 = ~n73234 & n74069;
  assign n74071 = n73221 & ~n73223;
  assign n74072 = ~n74070 & n74071;
  assign n74073 = ~n73218 & ~n74072;
  assign n74074 = n73175 & ~n73218;
  assign n74075 = n73188 & ~n73200;
  assign n74076 = ~n73607 & ~n74075;
  assign n74077 = n74074 & ~n74076;
  assign n74078 = ~n74073 & ~n74077;
  assign n74079 = ~n73175 & n73211;
  assign n74080 = n74078 & ~n74079;
  assign n74081 = ~n73182 & n73246;
  assign n74082 = ~n73182 & n73258;
  assign n74083 = ~n74081 & ~n74082;
  assign n74084 = n73175 & ~n74083;
  assign n74085 = n73175 & n73205;
  assign n74086 = ~n73182 & n74085;
  assign n74087 = ~n74084 & ~n74086;
  assign n74088 = n73182 & n73368;
  assign n74089 = n73182 & n73613;
  assign n74090 = n73182 & n73257;
  assign n74091 = ~n73182 & n73235;
  assign n74092 = ~n74090 & ~n74091;
  assign n74093 = n73175 & ~n74092;
  assign n74094 = ~n74089 & ~n74093;
  assign n74095 = ~n73608 & ~n74081;
  assign n74096 = ~n73252 & n74095;
  assign n74097 = n74094 & n74096;
  assign n74098 = ~n74088 & n74097;
  assign n74099 = n73218 & ~n74098;
  assign n74100 = ~n73387 & ~n74099;
  assign n74101 = n74087 & n74100;
  assign po2341 = ~n74080 | ~n74101;
  assign n74103 = ~n73524 & ~n73531;
  assign n74104 = n73494 & ~n74103;
  assign n74105 = ~n73580 & ~n74104;
  assign n74106 = n73506 & ~n73512;
  assign n74107 = n73500 & n73534;
  assign n74108 = ~n74106 & ~n74107;
  assign n74109 = ~n73500 & ~n73506;
  assign n74110 = n73512 & n74109;
  assign n74111 = n74108 & ~n74110;
  assign n74112 = ~n73494 & ~n74111;
  assign n74113 = ~n73521 & ~n74112;
  assign n74114 = n73500 & n74050;
  assign n74115 = ~n74053 & ~n74114;
  assign n74116 = n74113 & n74115;
  assign n74117 = ~n73558 & ~n74116;
  assign n74118 = ~n73494 & n74106;
  assign n74119 = n73500 & n74118;
  assign n74120 = ~n74117 & ~n74119;
  assign n74121 = ~n73538 & ~n73562;
  assign n74122 = ~n73535 & ~n73563;
  assign n74123 = ~n74036 & n74122;
  assign n74124 = n73494 & ~n74123;
  assign n74125 = ~n73500 & n73523;
  assign n74126 = ~n73542 & ~n74125;
  assign n74127 = ~n73494 & ~n74126;
  assign n74128 = ~n74039 & ~n74127;
  assign n74129 = ~n74124 & n74128;
  assign n74130 = n74121 & n74129;
  assign n74131 = n73558 & ~n74130;
  assign n74132 = n74120 & ~n74131;
  assign n74133 = n74105 & n74132;
  assign n74134 = pi2288 & n74133;
  assign n74135 = ~pi2288 & ~n74133;
  assign po2346 = n74134 | n74135;
  assign n74137 = n73626 & n73668;
  assign n74138 = ~n73701 & ~n74137;
  assign n74139 = ~n73656 & n74138;
  assign n74140 = n73632 & ~n74139;
  assign n74141 = ~n73639 & ~n73653;
  assign n74142 = ~n73654 & ~n74141;
  assign n74143 = n73626 & n74142;
  assign n74144 = ~n73626 & ~n73667;
  assign n74145 = ~n74143 & ~n74144;
  assign n74146 = ~n73749 & ~n74145;
  assign n74147 = ~n73632 & ~n74146;
  assign n74148 = ~n74140 & ~n74147;
  assign n74149 = n73694 & ~n74148;
  assign n74150 = n73657 & n73982;
  assign n74151 = ~n73659 & ~n73746;
  assign n74152 = ~n73729 & ~n74137;
  assign n74153 = ~n73632 & ~n74152;
  assign n74154 = ~n73665 & ~n74153;
  assign n74155 = n73633 & ~n73653;
  assign n74156 = n74154 & ~n74155;
  assign n74157 = n74151 & n74156;
  assign n74158 = ~n73737 & n74157;
  assign n74159 = ~n74150 & n74158;
  assign n74160 = ~n73694 & ~n74159;
  assign n74161 = ~n73626 & n73725;
  assign n74162 = ~n74160 & ~n74161;
  assign n74163 = n73626 & n73676;
  assign n74164 = ~n73955 & ~n74163;
  assign n74165 = n73632 & ~n74164;
  assign n74166 = ~n73744 & ~n74165;
  assign n74167 = n74162 & n74166;
  assign n74168 = ~n73747 & n74167;
  assign po2348 = n74149 | ~n74168;
  assign n74170 = ~n73500 & n74037;
  assign n74171 = n73506 & n73576;
  assign n74172 = n73512 & n74171;
  assign n74173 = ~n73524 & ~n74172;
  assign n74174 = ~n74030 & n74173;
  assign n74175 = ~n74170 & n74174;
  assign n74176 = ~n73494 & n73525;
  assign n74177 = n74175 & ~n74176;
  assign n74178 = n73558 & ~n74177;
  assign n74179 = ~n73500 & n73561;
  assign n74180 = n73527 & ~n74179;
  assign n74181 = ~n74056 & n74180;
  assign n74182 = n73494 & ~n74181;
  assign n74183 = ~n74178 & ~n74182;
  assign n74184 = ~n73562 & ~n74028;
  assign n74185 = ~n73494 & ~n74184;
  assign n74186 = n73494 & ~n73558;
  assign n74187 = n73568 & n74186;
  assign n74188 = ~n73500 & n73537;
  assign n74189 = ~n73512 & n74109;
  assign n74190 = ~n74037 & ~n74189;
  assign n74191 = ~n73520 & n74190;
  assign n74192 = ~n73494 & ~n74191;
  assign n74193 = ~n74188 & ~n74192;
  assign n74194 = ~n73558 & ~n74193;
  assign n74195 = ~n74187 & ~n74194;
  assign n74196 = ~n74185 & n74195;
  assign n74197 = n74183 & n74196;
  assign n74198 = pi2276 & n74197;
  assign n74199 = ~pi2276 & ~n74197;
  assign po2352 = n74198 | n74199;
  assign n74201 = pi4645 & ~pi9040;
  assign n74202 = pi4476 & pi9040;
  assign n74203 = ~n74201 & ~n74202;
  assign n74204 = ~pi2258 & ~n74203;
  assign n74205 = pi2258 & n74203;
  assign n74206 = ~n74204 & ~n74205;
  assign n74207 = pi4504 & pi9040;
  assign n74208 = pi4764 & ~pi9040;
  assign n74209 = ~n74207 & ~n74208;
  assign n74210 = ~pi2251 & ~n74209;
  assign n74211 = pi2251 & n74209;
  assign n74212 = ~n74210 & ~n74211;
  assign n74213 = pi4656 & ~pi9040;
  assign n74214 = pi4313 & pi9040;
  assign n74215 = ~n74213 & ~n74214;
  assign n74216 = ~pi2240 & n74215;
  assign n74217 = pi2240 & ~n74215;
  assign n74218 = ~n74216 & ~n74217;
  assign n74219 = pi4804 & pi9040;
  assign n74220 = pi4584 & ~pi9040;
  assign n74221 = ~n74219 & ~n74220;
  assign n74222 = ~pi2234 & ~n74221;
  assign n74223 = pi2234 & n74221;
  assign n74224 = ~n74222 & ~n74223;
  assign n74225 = pi4534 & pi9040;
  assign n74226 = pi4503 & ~pi9040;
  assign n74227 = ~n74225 & ~n74226;
  assign n74228 = pi2217 & n74227;
  assign n74229 = ~pi2217 & ~n74227;
  assign n74230 = ~n74228 & ~n74229;
  assign n74231 = n74224 & n74230;
  assign n74232 = n74218 & n74231;
  assign n74233 = n74212 & n74232;
  assign n74234 = pi4536 & pi9040;
  assign n74235 = pi4729 & ~pi9040;
  assign n74236 = ~n74234 & ~n74235;
  assign n74237 = pi2253 & n74236;
  assign n74238 = ~pi2253 & ~n74236;
  assign n74239 = ~n74237 & ~n74238;
  assign n74240 = ~n74218 & ~n74224;
  assign n74241 = n74239 & n74240;
  assign n74242 = ~n74218 & ~n74230;
  assign n74243 = ~n74241 & ~n74242;
  assign n74244 = n74212 & ~n74243;
  assign n74245 = ~n74233 & ~n74244;
  assign n74246 = n74206 & ~n74245;
  assign n74247 = n74218 & ~n74224;
  assign n74248 = n74230 & n74247;
  assign n74249 = n74206 & n74248;
  assign n74250 = n74239 & n74249;
  assign n74251 = ~n74246 & ~n74250;
  assign n74252 = ~n74230 & n74239;
  assign n74253 = ~n74218 & n74252;
  assign n74254 = ~n74239 & n74247;
  assign n74255 = ~n74230 & n74254;
  assign n74256 = ~n74253 & ~n74255;
  assign n74257 = n74212 & ~n74256;
  assign n74258 = ~n74218 & n74224;
  assign n74259 = ~n74247 & ~n74258;
  assign n74260 = n74230 & ~n74239;
  assign n74261 = ~n74259 & n74260;
  assign n74262 = ~n74230 & ~n74239;
  assign n74263 = n74218 & n74262;
  assign n74264 = n74224 & n74263;
  assign n74265 = ~n74261 & ~n74264;
  assign n74266 = n74230 & n74240;
  assign n74267 = n74239 & n74266;
  assign n74268 = ~n74212 & n74267;
  assign n74269 = n74265 & ~n74268;
  assign n74270 = n74232 & n74239;
  assign n74271 = ~n74230 & ~n74259;
  assign n74272 = n74239 & n74271;
  assign n74273 = ~n74270 & ~n74272;
  assign n74274 = n74212 & ~n74239;
  assign n74275 = ~n74224 & n74230;
  assign n74276 = n74274 & n74275;
  assign n74277 = ~n74230 & n74240;
  assign n74278 = ~n74212 & ~n74239;
  assign n74279 = n74277 & n74278;
  assign n74280 = ~n74276 & ~n74279;
  assign n74281 = n74273 & n74280;
  assign n74282 = n74269 & n74281;
  assign n74283 = ~n74206 & ~n74282;
  assign n74284 = n74230 & n74258;
  assign n74285 = n74218 & n74224;
  assign n74286 = ~n74230 & n74285;
  assign n74287 = ~n74284 & ~n74286;
  assign n74288 = ~n74218 & n74260;
  assign n74289 = n74287 & ~n74288;
  assign n74290 = n74206 & ~n74212;
  assign n74291 = ~n74289 & n74290;
  assign n74292 = ~n74283 & ~n74291;
  assign n74293 = ~n74257 & n74292;
  assign po2354 = ~n74251 | ~n74293;
  assign n74295 = ~n73900 & ~n73912;
  assign n74296 = ~n73896 & ~n74295;
  assign n74297 = n73880 & n73885;
  assign n74298 = ~n73888 & ~n74297;
  assign n74299 = ~n73924 & n74298;
  assign n74300 = ~n74296 & n74299;
  assign n74301 = n73883 & n73896;
  assign n74302 = n74300 & ~n74301;
  assign n74303 = ~n73947 & n74302;
  assign n74304 = n73910 & ~n74303;
  assign n74305 = ~n73880 & n73887;
  assign n74306 = n73880 & n73923;
  assign n74307 = n73880 & n73922;
  assign n74308 = n73874 & n73921;
  assign n74309 = ~n73896 & n74308;
  assign n74310 = ~n74307 & ~n74309;
  assign n74311 = ~n73935 & n74310;
  assign n74312 = ~n74306 & n74311;
  assign n74313 = ~n73868 & ~n73874;
  assign n74314 = n73862 & n73880;
  assign n74315 = ~n74313 & ~n74314;
  assign n74316 = ~n73930 & n74315;
  assign n74317 = n73896 & ~n74316;
  assign n74318 = n74312 & ~n74317;
  assign n74319 = ~n73943 & n74318;
  assign n74320 = ~n74305 & n74319;
  assign n74321 = ~n73910 & ~n74320;
  assign po2357 = ~n74304 & ~n74321;
  assign n74323 = n73778 & n73784;
  assign n74324 = n73765 & n74323;
  assign n74325 = ~n73759 & ~n73784;
  assign n74326 = n73772 & n74325;
  assign n74327 = ~n73778 & n74326;
  assign n74328 = n73772 & n73778;
  assign n74329 = n73759 & n74328;
  assign n74330 = ~n73759 & n73784;
  assign n74331 = ~n73838 & ~n74330;
  assign n74332 = ~n73813 & n74331;
  assign n74333 = ~n73772 & ~n74332;
  assign n74334 = ~n74329 & ~n74333;
  assign n74335 = ~n73778 & n73805;
  assign n74336 = n74334 & ~n74335;
  assign n74337 = ~n74327 & n74336;
  assign n74338 = ~n74324 & n74337;
  assign n74339 = ~n73793 & ~n74338;
  assign n74340 = n73784 & n73794;
  assign n74341 = ~n73778 & n74340;
  assign n74342 = n73766 & n73784;
  assign n74343 = n73778 & n74342;
  assign n74344 = ~n74341 & ~n74343;
  assign n74345 = ~n73772 & ~n74344;
  assign n74346 = ~n74339 & ~n74345;
  assign n74347 = ~n73816 & ~n73826;
  assign n74348 = ~n73772 & ~n74347;
  assign n74349 = ~n73830 & ~n74348;
  assign n74350 = n73778 & n73805;
  assign n74351 = n74349 & ~n74350;
  assign n74352 = n73793 & ~n74351;
  assign n74353 = ~n73766 & ~n73799;
  assign n74354 = ~n73784 & ~n74353;
  assign n74355 = ~n73820 & ~n74354;
  assign n74356 = n73772 & ~n74355;
  assign n74357 = n73793 & n74356;
  assign n74358 = ~n74352 & ~n74357;
  assign po2360 = ~n74346 | ~n74358;
  assign n74360 = ~n73765 & ~n73784;
  assign n74361 = ~n74340 & ~n74360;
  assign n74362 = n73798 & ~n74361;
  assign n74363 = ~n73816 & ~n73829;
  assign n74364 = ~n73826 & n74363;
  assign n74365 = ~n74342 & n74364;
  assign n74366 = n73778 & ~n74365;
  assign n74367 = ~n74335 & ~n74366;
  assign n74368 = ~n74362 & n74367;
  assign n74369 = ~n73793 & ~n74368;
  assign n74370 = n73778 & n74354;
  assign n74371 = n73772 & ~n74361;
  assign n74372 = ~n74370 & ~n74371;
  assign n74373 = ~n73778 & n73826;
  assign n74374 = ~n73765 & n74323;
  assign n74375 = ~n73845 & ~n74374;
  assign n74376 = ~n74342 & n74375;
  assign n74377 = ~n73772 & ~n74376;
  assign n74378 = ~n74373 & ~n74377;
  assign n74379 = n74372 & n74378;
  assign n74380 = n73793 & ~n74379;
  assign n74381 = ~n74369 & ~n74380;
  assign n74382 = n73778 & n74340;
  assign n74383 = ~n74373 & ~n74382;
  assign n74384 = n73772 & ~n74383;
  assign n74385 = n74381 & ~n74384;
  assign n74386 = pi2306 & n74385;
  assign n74387 = ~pi2306 & ~n74385;
  assign po2362 = n74386 | n74387;
  assign n74389 = ~n73884 & ~n73921;
  assign n74390 = n73874 & ~n73880;
  assign n74391 = ~n74389 & n74390;
  assign n74392 = ~n74306 & ~n74391;
  assign n74393 = ~n73887 & n74392;
  assign n74394 = n73896 & ~n74393;
  assign n74395 = n73880 & n73936;
  assign n74396 = ~n74394 & ~n74395;
  assign n74397 = n73880 & n73884;
  assign n74398 = ~n73880 & n74313;
  assign n74399 = ~n74397 & ~n74398;
  assign n74400 = ~n73911 & n74399;
  assign n74401 = ~n73896 & ~n74400;
  assign n74402 = n74396 & ~n74401;
  assign n74403 = n73910 & ~n74402;
  assign n74404 = n73883 & ~n73896;
  assign n74405 = ~n74403 & ~n74404;
  assign n74406 = n73880 & n73898;
  assign n74407 = ~n73918 & ~n74406;
  assign n74408 = n73896 & ~n74407;
  assign n74409 = ~n73880 & n73884;
  assign n74410 = ~n73923 & ~n74409;
  assign n74411 = ~n73896 & ~n74410;
  assign n74412 = ~n73888 & ~n74411;
  assign n74413 = ~n73883 & ~n73948;
  assign n74414 = n74412 & n74413;
  assign n74415 = ~n73880 & n73936;
  assign n74416 = n74414 & ~n74415;
  assign n74417 = n73880 & n73930;
  assign n74418 = ~n74313 & ~n74417;
  assign n74419 = ~n73911 & n74418;
  assign n74420 = n73896 & ~n74419;
  assign n74421 = n74416 & ~n74420;
  assign n74422 = ~n73910 & ~n74421;
  assign n74423 = ~n74408 & ~n74422;
  assign po2364 = ~n74405 | ~n74423;
  assign n74425 = ~n73311 & n73351;
  assign n74426 = n73280 & n73299;
  assign n74427 = ~n73303 & ~n74426;
  assign n74428 = n73311 & n74427;
  assign n74429 = ~n74425 & ~n74428;
  assign n74430 = ~n73338 & ~n74429;
  assign n74431 = n73274 & ~n74430;
  assign n74432 = n73311 & n73330;
  assign n74433 = ~n74431 & ~n74432;
  assign n74434 = ~n73990 & ~n74009;
  assign n74435 = ~n73311 & ~n74434;
  assign n74436 = ~n73286 & n73318;
  assign n74437 = ~n73347 & ~n74436;
  assign n74438 = n73292 & ~n74437;
  assign n74439 = n73300 & ~n73311;
  assign n74440 = ~n73280 & n73321;
  assign n74441 = ~n74439 & ~n74440;
  assign n74442 = ~n73401 & n74441;
  assign n74443 = ~n74012 & n74442;
  assign n74444 = ~n74438 & n74443;
  assign n74445 = ~n73274 & ~n74444;
  assign n74446 = ~n74435 & ~n74445;
  assign n74447 = n74433 & n74446;
  assign n74448 = pi2321 & n74447;
  assign n74449 = ~pi2321 & ~n74447;
  assign po2366 = n74448 | n74449;
  assign n74451 = ~n74239 & n74240;
  assign n74452 = n74239 & n74247;
  assign n74453 = ~n74451 & ~n74452;
  assign n74454 = n74212 & ~n74453;
  assign n74455 = n74212 & n74264;
  assign n74456 = ~n74454 & ~n74455;
  assign n74457 = n74206 & ~n74456;
  assign n74458 = ~n74259 & n74262;
  assign n74459 = n74224 & ~n74230;
  assign n74460 = ~n74258 & ~n74459;
  assign n74461 = ~n74239 & ~n74460;
  assign n74462 = ~n74266 & ~n74461;
  assign n74463 = ~n74212 & ~n74462;
  assign n74464 = ~n74458 & ~n74463;
  assign n74465 = n74239 & n74277;
  assign n74466 = n74218 & n74260;
  assign n74467 = n74239 & ~n74460;
  assign n74468 = ~n74466 & ~n74467;
  assign n74469 = n74212 & ~n74468;
  assign n74470 = ~n74465 & ~n74469;
  assign n74471 = n74464 & n74470;
  assign n74472 = ~n74206 & ~n74471;
  assign n74473 = n74212 & n74252;
  assign n74474 = n74258 & n74473;
  assign n74475 = ~n74212 & n74239;
  assign n74476 = n74218 & n74230;
  assign n74477 = n74475 & n74476;
  assign n74478 = ~n74474 & ~n74477;
  assign n74479 = n74230 & n74239;
  assign n74480 = n74206 & ~n74258;
  assign n74481 = n74479 & n74480;
  assign n74482 = n74478 & ~n74481;
  assign n74483 = n74224 & n74239;
  assign n74484 = ~n74248 & ~n74483;
  assign n74485 = n74290 & ~n74484;
  assign n74486 = n74482 & ~n74485;
  assign n74487 = ~n74472 & n74486;
  assign n74488 = ~n74457 & n74487;
  assign n74489 = pi2297 & n74488;
  assign n74490 = ~pi2297 & ~n74488;
  assign po2367 = n74489 | n74490;
  assign n74492 = n74212 & n74266;
  assign n74493 = ~n74239 & n74492;
  assign n74494 = ~n74455 & ~n74493;
  assign n74495 = ~n74240 & n74274;
  assign n74496 = ~n74230 & n74495;
  assign n74497 = n74230 & n74483;
  assign n74498 = ~n74241 & ~n74497;
  assign n74499 = n74212 & ~n74498;
  assign n74500 = ~n74496 & ~n74499;
  assign n74501 = ~n74264 & ~n74279;
  assign n74502 = ~n74259 & ~n74262;
  assign n74503 = ~n74212 & n74502;
  assign n74504 = n74501 & ~n74503;
  assign n74505 = n74500 & n74504;
  assign n74506 = n74206 & ~n74505;
  assign n74507 = n74494 & ~n74506;
  assign n74508 = n74239 & n74286;
  assign n74509 = ~n74230 & n74483;
  assign n74510 = ~n74451 & ~n74509;
  assign n74511 = n74247 & ~n74262;
  assign n74512 = n74510 & ~n74511;
  assign n74513 = n74212 & ~n74512;
  assign n74514 = ~n74508 & ~n74513;
  assign n74515 = ~n74206 & ~n74514;
  assign n74516 = ~n74212 & n74284;
  assign n74517 = n74239 & n74516;
  assign n74518 = ~n74206 & ~n74212;
  assign n74519 = ~n74232 & ~n74241;
  assign n74520 = ~n74458 & n74519;
  assign n74521 = n74518 & ~n74520;
  assign n74522 = ~n74517 & ~n74521;
  assign n74523 = ~n74515 & n74522;
  assign n74524 = n74507 & n74523;
  assign n74525 = pi2289 & ~n74524;
  assign n74526 = ~pi2289 & n74524;
  assign po2368 = n74525 | n74526;
  assign n74528 = ~n74254 & ~n74277;
  assign n74529 = ~n74284 & n74528;
  assign n74530 = ~n74212 & ~n74529;
  assign n74531 = ~n74230 & n74258;
  assign n74532 = ~n74266 & ~n74531;
  assign n74533 = n74212 & ~n74532;
  assign n74534 = ~n74530 & ~n74533;
  assign n74535 = ~n74233 & n74534;
  assign n74536 = ~n74255 & n74535;
  assign n74537 = ~n74206 & ~n74536;
  assign n74538 = ~n74239 & n74285;
  assign n74539 = ~n74452 & ~n74538;
  assign n74540 = ~n74212 & ~n74539;
  assign n74541 = ~n74267 & ~n74540;
  assign n74542 = n74212 & n74248;
  assign n74543 = ~n74277 & ~n74542;
  assign n74544 = n74287 & n74543;
  assign n74545 = ~n74239 & ~n74544;
  assign n74546 = n74541 & ~n74545;
  assign n74547 = n74206 & ~n74546;
  assign n74548 = ~n74230 & n74452;
  assign n74549 = ~n74270 & ~n74548;
  assign n74550 = n74212 & ~n74549;
  assign n74551 = n74459 & n74475;
  assign n74552 = ~n74550 & ~n74551;
  assign n74553 = ~n74547 & n74552;
  assign n74554 = ~n74537 & n74553;
  assign n74555 = pi2281 & n74554;
  assign n74556 = ~pi2281 & ~n74554;
  assign po2369 = n74555 | n74556;
  assign n74558 = ~n73778 & n74360;
  assign n74559 = n73778 & n73799;
  assign n74560 = ~n73825 & ~n74559;
  assign n74561 = n73772 & ~n74560;
  assign n74562 = ~n73772 & n74342;
  assign n74563 = n73778 & n73843;
  assign n74564 = ~n74324 & ~n74563;
  assign n74565 = ~n74562 & n74564;
  assign n74566 = ~n74561 & n74565;
  assign n74567 = ~n74558 & n74566;
  assign n74568 = n73793 & ~n74567;
  assign n74569 = n73772 & ~n73793;
  assign n74570 = n73778 & n73816;
  assign n74571 = ~n73829 & ~n74570;
  assign n74572 = ~n74342 & n74571;
  assign n74573 = n74569 & ~n74572;
  assign n74574 = ~n73772 & n74340;
  assign n74575 = ~n73787 & ~n73813;
  assign n74576 = ~n73807 & n74575;
  assign n74577 = ~n74574 & n74576;
  assign n74578 = ~n73793 & ~n74577;
  assign n74579 = ~n74573 & ~n74578;
  assign n74580 = n73826 & n74328;
  assign n74581 = ~n73778 & n73829;
  assign n74582 = ~n74335 & ~n74581;
  assign n74583 = n73772 & ~n74582;
  assign n74584 = ~n74580 & ~n74583;
  assign n74585 = ~n73837 & n74584;
  assign n74586 = ~n73778 & n74562;
  assign n74587 = n74585 & ~n74586;
  assign n74588 = n74579 & n74587;
  assign n74589 = ~n74568 & n74588;
  assign n74590 = pi2311 & n74589;
  assign n74591 = ~pi2311 & ~n74589;
  assign po2370 = n74590 | n74591;
  assign n74593 = ~n73874 & ~n74389;
  assign n74594 = n73880 & n74593;
  assign n74595 = ~n74306 & ~n74594;
  assign n74596 = n73896 & ~n74595;
  assign n74597 = ~n73896 & n73935;
  assign n74598 = ~n74596 & ~n74597;
  assign n74599 = ~n73880 & n73916;
  assign n74600 = ~n74305 & ~n74599;
  assign n74601 = ~n73896 & n74600;
  assign n74602 = ~n73862 & n73874;
  assign n74603 = ~n73880 & n74602;
  assign n74604 = ~n74397 & ~n74406;
  assign n74605 = n73896 & n74604;
  assign n74606 = ~n74593 & n74605;
  assign n74607 = ~n74603 & n74606;
  assign n74608 = ~n74601 & ~n74607;
  assign n74609 = n74595 & ~n74608;
  assign n74610 = n73910 & ~n74609;
  assign n74611 = ~n73896 & ~n74389;
  assign n74612 = n73874 & n74611;
  assign n74613 = n73880 & n73886;
  assign n74614 = ~n73948 & ~n74613;
  assign n74615 = ~n73896 & ~n74614;
  assign n74616 = ~n74612 & ~n74615;
  assign n74617 = ~n73880 & n74611;
  assign n74618 = n74616 & ~n74617;
  assign n74619 = ~n73910 & ~n74618;
  assign n74620 = ~n74610 & ~n74619;
  assign n74621 = n73896 & ~n74600;
  assign n74622 = ~n73935 & ~n74621;
  assign n74623 = ~n73910 & ~n74622;
  assign n74624 = n74620 & ~n74623;
  assign po2372 = ~n74598 | ~n74624;
  assign n74626 = pi4674 & pi9040;
  assign n74627 = pi4969 & ~pi9040;
  assign n74628 = ~n74626 & ~n74627;
  assign n74629 = ~pi2324 & ~n74628;
  assign n74630 = pi2324 & n74628;
  assign n74631 = ~n74629 & ~n74630;
  assign n74632 = pi4756 & pi9040;
  assign n74633 = pi4672 & ~pi9040;
  assign n74634 = ~n74632 & ~n74633;
  assign n74635 = pi2319 & n74634;
  assign n74636 = ~pi2319 & ~n74634;
  assign n74637 = ~n74635 & ~n74636;
  assign n74638 = pi4725 & ~pi9040;
  assign n74639 = pi4873 & pi9040;
  assign n74640 = ~n74638 & ~n74639;
  assign n74641 = pi2335 & n74640;
  assign n74642 = ~pi2335 & ~n74640;
  assign n74643 = ~n74641 & ~n74642;
  assign n74644 = ~n74637 & n74643;
  assign n74645 = pi4732 & pi9040;
  assign n74646 = pi4756 & ~pi9040;
  assign n74647 = ~n74645 & ~n74646;
  assign n74648 = ~pi2312 & ~n74647;
  assign n74649 = pi2312 & n74647;
  assign n74650 = ~n74648 & ~n74649;
  assign n74651 = pi4658 & pi9040;
  assign n74652 = pi4980 & ~pi9040;
  assign n74653 = ~n74651 & ~n74652;
  assign n74654 = ~pi2275 & ~n74653;
  assign n74655 = pi2275 & n74653;
  assign n74656 = ~n74654 & ~n74655;
  assign n74657 = n74650 & n74656;
  assign n74658 = n74644 & n74657;
  assign n74659 = pi4732 & ~pi9040;
  assign n74660 = pi4722 & pi9040;
  assign n74661 = ~n74659 & ~n74660;
  assign n74662 = ~pi2327 & ~n74661;
  assign n74663 = pi2327 & n74661;
  assign n74664 = ~n74662 & ~n74663;
  assign n74665 = ~n74650 & n74656;
  assign n74666 = n74637 & n74643;
  assign n74667 = n74665 & n74666;
  assign n74668 = n74664 & n74667;
  assign n74669 = n74650 & ~n74656;
  assign n74670 = n74664 & n74669;
  assign n74671 = n74643 & n74670;
  assign n74672 = n74637 & n74671;
  assign n74673 = ~n74637 & n74664;
  assign n74674 = ~n74656 & n74673;
  assign n74675 = ~n74650 & n74674;
  assign n74676 = ~n74672 & ~n74675;
  assign n74677 = ~n74668 & n74676;
  assign n74678 = ~n74658 & n74677;
  assign n74679 = ~n74637 & ~n74664;
  assign n74680 = n74657 & n74679;
  assign n74681 = n74678 & ~n74680;
  assign n74682 = ~n74631 & ~n74681;
  assign n74683 = n74650 & n74664;
  assign n74684 = n74656 & n74683;
  assign n74685 = n74637 & n74684;
  assign n74686 = ~n74674 & ~n74685;
  assign n74687 = ~n74664 & n74665;
  assign n74688 = n74637 & n74687;
  assign n74689 = n74686 & ~n74688;
  assign n74690 = ~n74643 & ~n74689;
  assign n74691 = ~n74650 & ~n74656;
  assign n74692 = ~n74637 & n74691;
  assign n74693 = ~n74650 & n74673;
  assign n74694 = ~n74692 & ~n74693;
  assign n74695 = ~n74643 & ~n74694;
  assign n74696 = ~n74656 & ~n74664;
  assign n74697 = n74650 & n74696;
  assign n74698 = ~n74643 & n74697;
  assign n74699 = n74637 & n74698;
  assign n74700 = ~n74695 & ~n74699;
  assign n74701 = ~n74631 & ~n74700;
  assign n74702 = ~n74690 & ~n74701;
  assign n74703 = ~n74682 & n74702;
  assign n74704 = n74637 & ~n74664;
  assign n74705 = n74643 & n74704;
  assign n74706 = n74691 & n74705;
  assign n74707 = n74650 & ~n74664;
  assign n74708 = n74644 & n74707;
  assign n74709 = ~n74643 & n74664;
  assign n74710 = n74650 & n74709;
  assign n74711 = n74637 & ~n74650;
  assign n74712 = ~n74664 & n74711;
  assign n74713 = ~n74710 & ~n74712;
  assign n74714 = ~n74637 & n74697;
  assign n74715 = n74713 & ~n74714;
  assign n74716 = ~n74687 & n74715;
  assign n74717 = n74643 & n74665;
  assign n74718 = ~n74637 & n74717;
  assign n74719 = n74637 & n74691;
  assign n74720 = n74656 & ~n74664;
  assign n74721 = ~n74719 & ~n74720;
  assign n74722 = n74643 & ~n74721;
  assign n74723 = ~n74718 & ~n74722;
  assign n74724 = n74716 & n74723;
  assign n74725 = n74631 & ~n74724;
  assign n74726 = ~n74708 & ~n74725;
  assign n74727 = ~n74706 & n74726;
  assign n74728 = n74703 & n74727;
  assign n74729 = pi2357 & n74728;
  assign n74730 = ~pi2357 & ~n74728;
  assign po2428 = n74729 | n74730;
  assign n74732 = ~n74650 & n74664;
  assign n74733 = ~n74680 & ~n74732;
  assign n74734 = ~n74711 & n74733;
  assign n74735 = n74643 & ~n74734;
  assign n74736 = n74637 & ~n74643;
  assign n74737 = n74650 & n74736;
  assign n74738 = n74637 & n74664;
  assign n74739 = n74656 & n74738;
  assign n74740 = ~n74637 & n74670;
  assign n74741 = ~n74739 & ~n74740;
  assign n74742 = ~n74650 & ~n74664;
  assign n74743 = ~n74637 & ~n74643;
  assign n74744 = n74742 & n74743;
  assign n74745 = n74741 & ~n74744;
  assign n74746 = ~n74737 & n74745;
  assign n74747 = ~n74735 & n74746;
  assign n74748 = n74631 & ~n74747;
  assign n74749 = n74664 & n74665;
  assign n74750 = ~n74637 & n74749;
  assign n74751 = ~n74656 & n74732;
  assign n74752 = n74637 & n74751;
  assign n74753 = ~n74750 & ~n74752;
  assign n74754 = n74643 & ~n74753;
  assign n74755 = ~n74748 & ~n74754;
  assign n74756 = n74637 & n74670;
  assign n74757 = ~n74684 & ~n74697;
  assign n74758 = n74643 & ~n74757;
  assign n74759 = ~n74756 & ~n74758;
  assign n74760 = ~n74688 & n74759;
  assign n74761 = ~n74631 & ~n74760;
  assign n74762 = ~n74657 & ~n74691;
  assign n74763 = ~n74664 & ~n74762;
  assign n74764 = ~n74692 & ~n74763;
  assign n74765 = ~n74643 & ~n74764;
  assign n74766 = ~n74631 & n74765;
  assign n74767 = ~n74761 & ~n74766;
  assign n74768 = n74755 & n74767;
  assign n74769 = pi2363 & ~n74768;
  assign n74770 = ~pi2363 & n74755;
  assign n74771 = n74767 & n74770;
  assign po2436 = n74769 | n74771;
  assign n74773 = ~n74637 & n74687;
  assign n74774 = ~n74740 & ~n74773;
  assign n74775 = ~n74643 & ~n74774;
  assign n74776 = n74684 & n74736;
  assign n74777 = ~n74775 & ~n74776;
  assign n74778 = ~n74708 & n74777;
  assign n74779 = n74643 & n74664;
  assign n74780 = ~n74656 & n74779;
  assign n74781 = ~n74650 & n74780;
  assign n74782 = ~n74637 & n74781;
  assign n74783 = n74643 & n74749;
  assign n74784 = ~n74680 & ~n74706;
  assign n74785 = ~n74672 & n74784;
  assign n74786 = ~n74783 & n74785;
  assign n74787 = n74631 & ~n74786;
  assign n74788 = n74637 & n74697;
  assign n74789 = ~n74687 & ~n74788;
  assign n74790 = ~n74751 & n74789;
  assign n74791 = ~n74643 & ~n74790;
  assign n74792 = n74631 & n74791;
  assign n74793 = n74637 & n74717;
  assign n74794 = ~n74781 & ~n74793;
  assign n74795 = ~n74739 & n74794;
  assign n74796 = ~n74656 & n74679;
  assign n74797 = n74637 & n74657;
  assign n74798 = ~n74683 & ~n74797;
  assign n74799 = ~n74643 & ~n74798;
  assign n74800 = ~n74796 & ~n74799;
  assign n74801 = n74795 & n74800;
  assign n74802 = ~n74631 & ~n74801;
  assign n74803 = ~n74792 & ~n74802;
  assign n74804 = ~n74787 & n74803;
  assign n74805 = ~n74782 & n74804;
  assign n74806 = n74778 & n74805;
  assign n74807 = pi2368 & ~n74806;
  assign n74808 = ~pi2368 & n74778;
  assign n74809 = n74805 & n74808;
  assign po2446 = n74807 | n74809;
  assign n74811 = n74637 & n74763;
  assign n74812 = ~n74696 & ~n74749;
  assign n74813 = ~n74643 & ~n74812;
  assign n74814 = ~n74811 & ~n74813;
  assign n74815 = ~n74656 & n74738;
  assign n74816 = ~n74720 & ~n74815;
  assign n74817 = ~n74751 & n74816;
  assign n74818 = n74643 & ~n74817;
  assign n74819 = n74814 & ~n74818;
  assign n74820 = ~n74637 & n74684;
  assign n74821 = n74819 & ~n74820;
  assign n74822 = ~n74631 & ~n74821;
  assign n74823 = n74644 & ~n74812;
  assign n74824 = ~n74687 & ~n74697;
  assign n74825 = ~n74684 & ~n74751;
  assign n74826 = n74824 & n74825;
  assign n74827 = n74637 & ~n74826;
  assign n74828 = ~n74823 & ~n74827;
  assign n74829 = ~n74740 & n74828;
  assign n74830 = n74631 & ~n74829;
  assign n74831 = ~n74822 & ~n74830;
  assign n74832 = n74637 & n74749;
  assign n74833 = ~n74820 & ~n74832;
  assign n74834 = ~n74643 & ~n74833;
  assign n74835 = n74831 & ~n74834;
  assign n74836 = pi2373 & ~n74835;
  assign n74837 = ~pi2373 & ~n74834;
  assign n74838 = ~n74830 & n74837;
  assign n74839 = ~n74822 & n74838;
  assign po2447 = n74836 | n74839;
  assign n74841 = pi4867 & pi9040;
  assign n74842 = pi4721 & ~pi9040;
  assign n74843 = ~n74841 & ~n74842;
  assign n74844 = pi2308 & n74843;
  assign n74845 = ~pi2308 & ~n74843;
  assign n74846 = ~n74844 & ~n74845;
  assign n74847 = pi4721 & pi9040;
  assign n74848 = pi5054 & ~pi9040;
  assign n74849 = ~n74847 & ~n74848;
  assign n74850 = ~pi2324 & ~n74849;
  assign n74851 = pi2324 & n74849;
  assign n74852 = ~n74850 & ~n74851;
  assign n74853 = pi4542 & ~pi9040;
  assign n74854 = pi4871 & pi9040;
  assign n74855 = ~n74853 & ~n74854;
  assign n74856 = ~pi2329 & n74855;
  assign n74857 = pi2329 & ~n74855;
  assign n74858 = ~n74856 & ~n74857;
  assign n74859 = n74852 & n74858;
  assign n74860 = pi4661 & ~pi9040;
  assign n74861 = pi5054 & pi9040;
  assign n74862 = ~n74860 & ~n74861;
  assign n74863 = ~pi2275 & n74862;
  assign n74864 = pi2275 & ~n74862;
  assign n74865 = ~n74863 & ~n74864;
  assign n74866 = pi4719 & pi9040;
  assign n74867 = pi4724 & ~pi9040;
  assign n74868 = ~n74866 & ~n74867;
  assign n74869 = ~pi2314 & ~n74868;
  assign n74870 = pi2314 & n74868;
  assign n74871 = ~n74869 & ~n74870;
  assign n74872 = ~n74865 & n74871;
  assign n74873 = n74859 & n74872;
  assign n74874 = n74865 & n74871;
  assign n74875 = ~n74852 & n74874;
  assign n74876 = ~n74873 & ~n74875;
  assign n74877 = ~n74846 & ~n74876;
  assign n74878 = pi4666 & ~pi9040;
  assign n74879 = pi4725 & pi9040;
  assign n74880 = ~n74878 & ~n74879;
  assign n74881 = ~pi2334 & ~n74880;
  assign n74882 = pi2334 & n74880;
  assign n74883 = ~n74881 & ~n74882;
  assign n74884 = ~n74852 & ~n74858;
  assign n74885 = n74865 & n74884;
  assign n74886 = n74871 & n74885;
  assign n74887 = n74846 & ~n74871;
  assign n74888 = n74852 & n74887;
  assign n74889 = n74859 & n74865;
  assign n74890 = n74852 & ~n74858;
  assign n74891 = ~n74865 & n74890;
  assign n74892 = ~n74889 & ~n74891;
  assign n74893 = ~n74852 & n74858;
  assign n74894 = ~n74865 & n74893;
  assign n74895 = n74871 & n74894;
  assign n74896 = n74892 & ~n74895;
  assign n74897 = n74846 & ~n74896;
  assign n74898 = ~n74888 & ~n74897;
  assign n74899 = ~n74886 & n74898;
  assign n74900 = ~n74871 & n74893;
  assign n74901 = ~n74865 & n74884;
  assign n74902 = ~n74900 & ~n74901;
  assign n74903 = ~n74846 & ~n74902;
  assign n74904 = n74865 & n74890;
  assign n74905 = ~n74871 & n74904;
  assign n74906 = ~n74903 & ~n74905;
  assign n74907 = n74899 & n74906;
  assign n74908 = n74883 & ~n74907;
  assign n74909 = ~n74877 & ~n74908;
  assign n74910 = n74865 & n74893;
  assign n74911 = ~n74904 & ~n74910;
  assign n74912 = n74871 & ~n74911;
  assign n74913 = ~n74873 & ~n74912;
  assign n74914 = ~n74883 & ~n74913;
  assign n74915 = n74846 & ~n74883;
  assign n74916 = ~n74902 & n74915;
  assign n74917 = ~n74914 & ~n74916;
  assign n74918 = ~n74846 & ~n74883;
  assign n74919 = n74859 & ~n74871;
  assign n74920 = ~n74885 & ~n74919;
  assign n74921 = n74852 & ~n74865;
  assign n74922 = n74920 & ~n74921;
  assign n74923 = n74918 & ~n74922;
  assign n74924 = n74917 & ~n74923;
  assign n74925 = n74909 & n74924;
  assign n74926 = ~pi2349 & ~n74925;
  assign n74927 = pi2349 & n74917;
  assign n74928 = n74909 & n74927;
  assign n74929 = ~n74923 & n74928;
  assign po2452 = n74926 | n74929;
  assign n74931 = ~n74846 & n74871;
  assign n74932 = ~n74893 & ~n74904;
  assign n74933 = n74931 & ~n74932;
  assign n74934 = ~n74846 & n74865;
  assign n74935 = n74893 & n74934;
  assign n74936 = ~n74933 & ~n74935;
  assign n74937 = n74883 & ~n74936;
  assign n74938 = ~n74865 & ~n74871;
  assign n74939 = ~n74858 & n74938;
  assign n74940 = n74852 & n74939;
  assign n74941 = ~n74921 & ~n74938;
  assign n74942 = n74846 & ~n74941;
  assign n74943 = n74865 & ~n74871;
  assign n74944 = n74858 & n74943;
  assign n74945 = n74852 & n74944;
  assign n74946 = ~n74942 & ~n74945;
  assign n74947 = ~n74940 & n74946;
  assign n74948 = n74883 & ~n74947;
  assign n74949 = ~n74937 & ~n74948;
  assign n74950 = ~n74858 & n74872;
  assign n74951 = ~n74852 & n74950;
  assign n74952 = ~n74871 & n74885;
  assign n74953 = ~n74951 & ~n74952;
  assign n74954 = ~n74846 & ~n74953;
  assign n74955 = n74871 & n74910;
  assign n74956 = ~n74871 & n74921;
  assign n74957 = ~n74955 & ~n74956;
  assign n74958 = n74846 & ~n74957;
  assign n74959 = ~n74859 & ~n74921;
  assign n74960 = n74871 & ~n74959;
  assign n74961 = ~n74885 & ~n74960;
  assign n74962 = ~n74846 & ~n74961;
  assign n74963 = ~n74858 & ~n74871;
  assign n74964 = n74934 & n74963;
  assign n74965 = n74858 & ~n74865;
  assign n74966 = ~n74885 & ~n74965;
  assign n74967 = ~n74871 & ~n74966;
  assign n74968 = n74846 & n74871;
  assign n74969 = n74890 & n74968;
  assign n74970 = n74865 & n74969;
  assign n74971 = ~n74967 & ~n74970;
  assign n74972 = ~n74964 & n74971;
  assign n74973 = ~n74962 & n74972;
  assign n74974 = ~n74951 & n74973;
  assign n74975 = ~n74883 & ~n74974;
  assign n74976 = ~n74958 & ~n74975;
  assign n74977 = ~n74954 & n74976;
  assign n74978 = n74949 & n74977;
  assign n74979 = pi2361 & n74978;
  assign n74980 = ~pi2361 & ~n74978;
  assign po2453 = n74979 | n74980;
  assign n74982 = pi4950 & pi9040;
  assign n74983 = pi4722 & ~pi9040;
  assign n74984 = ~n74982 & ~n74983;
  assign n74985 = ~pi2304 & n74984;
  assign n74986 = pi2304 & ~n74984;
  assign n74987 = ~n74985 & ~n74986;
  assign n74988 = pi4540 & pi9040;
  assign n74989 = pi4873 & ~pi9040;
  assign n74990 = ~n74988 & ~n74989;
  assign n74991 = ~pi2333 & n74990;
  assign n74992 = pi2333 & ~n74990;
  assign n74993 = ~n74991 & ~n74992;
  assign n74994 = pi4542 & pi9040;
  assign n74995 = pi4726 & ~pi9040;
  assign n74996 = ~n74994 & ~n74995;
  assign n74997 = ~pi2320 & n74996;
  assign n74998 = pi2320 & ~n74996;
  assign n74999 = ~n74997 & ~n74998;
  assign n75000 = pi4595 & ~pi9040;
  assign n75001 = pi4659 & pi9040;
  assign n75002 = ~n75000 & ~n75001;
  assign n75003 = ~pi2295 & n75002;
  assign n75004 = pi2295 & ~n75002;
  assign n75005 = ~n75003 & ~n75004;
  assign n75006 = pi4540 & ~pi9040;
  assign n75007 = pi4980 & pi9040;
  assign n75008 = ~n75006 & ~n75007;
  assign n75009 = ~pi2326 & ~n75008;
  assign n75010 = pi2326 & n75008;
  assign n75011 = ~n75009 & ~n75010;
  assign n75012 = n75005 & ~n75011;
  assign n75013 = n74999 & n75012;
  assign n75014 = n74993 & n75013;
  assign n75015 = ~n74993 & n74999;
  assign n75016 = ~n75011 & n75015;
  assign n75017 = ~n75005 & n75016;
  assign n75018 = ~n75014 & ~n75017;
  assign n75019 = ~n74987 & ~n75018;
  assign n75020 = pi4871 & ~pi9040;
  assign n75021 = pi4595 & pi9040;
  assign n75022 = ~n75020 & ~n75021;
  assign n75023 = ~pi2313 & ~n75022;
  assign n75024 = pi2313 & n75022;
  assign n75025 = ~n75023 & ~n75024;
  assign n75026 = n75005 & n75011;
  assign n75027 = ~n74999 & n75026;
  assign n75028 = n74993 & n75027;
  assign n75029 = ~n75005 & ~n75011;
  assign n75030 = ~n74999 & n75029;
  assign n75031 = ~n74987 & n75030;
  assign n75032 = ~n75028 & ~n75031;
  assign n75033 = n74993 & ~n75005;
  assign n75034 = n74999 & n75033;
  assign n75035 = n74993 & ~n74999;
  assign n75036 = n75005 & n75035;
  assign n75037 = ~n75034 & ~n75036;
  assign n75038 = n74987 & ~n75037;
  assign n75039 = n74987 & n75012;
  assign n75040 = ~n74993 & n75039;
  assign n75041 = n74999 & n75040;
  assign n75042 = ~n74993 & ~n74999;
  assign n75043 = n75011 & n75042;
  assign n75044 = ~n75005 & n75043;
  assign n75045 = ~n74987 & n74999;
  assign n75046 = n75011 & n75045;
  assign n75047 = n75005 & n75046;
  assign n75048 = ~n75044 & ~n75047;
  assign n75049 = ~n75041 & n75048;
  assign n75050 = ~n75038 & n75049;
  assign n75051 = n75032 & n75050;
  assign n75052 = n75025 & ~n75051;
  assign n75053 = n74987 & n75028;
  assign n75054 = n74993 & n75031;
  assign n75055 = ~n75053 & ~n75054;
  assign n75056 = ~n75052 & n75055;
  assign n75057 = ~n75019 & n75056;
  assign n75058 = ~n74987 & ~n74993;
  assign n75059 = ~n74999 & n75005;
  assign n75060 = n75058 & n75059;
  assign n75061 = ~n74987 & n75013;
  assign n75062 = ~n75060 & ~n75061;
  assign n75063 = ~n75005 & n75011;
  assign n75064 = ~n74999 & n75063;
  assign n75065 = ~n74987 & n75064;
  assign n75066 = n74999 & n75063;
  assign n75067 = n74993 & n75066;
  assign n75068 = ~n75065 & ~n75067;
  assign n75069 = ~n74999 & n75012;
  assign n75070 = ~n74993 & n75069;
  assign n75071 = ~n75014 & ~n75070;
  assign n75072 = ~n74993 & n75029;
  assign n75073 = n74999 & n75011;
  assign n75074 = ~n75072 & ~n75073;
  assign n75075 = n74987 & ~n75074;
  assign n75076 = n75071 & ~n75075;
  assign n75077 = n75068 & n75076;
  assign n75078 = n75062 & n75077;
  assign n75079 = ~n75025 & ~n75078;
  assign n75080 = n75057 & ~n75079;
  assign n75081 = ~pi2343 & ~n75080;
  assign n75082 = pi2343 & n75057;
  assign n75083 = ~n75079 & n75082;
  assign po2457 = n75081 | n75083;
  assign n75085 = pi4541 & pi9040;
  assign n75086 = pi4664 & ~pi9040;
  assign n75087 = ~n75085 & ~n75086;
  assign n75088 = ~pi2298 & n75087;
  assign n75089 = pi2298 & ~n75087;
  assign n75090 = ~n75088 & ~n75089;
  assign n75091 = pi4668 & pi9040;
  assign n75092 = pi4955 & ~pi9040;
  assign n75093 = ~n75091 & ~n75092;
  assign n75094 = ~pi2322 & ~n75093;
  assign n75095 = pi2322 & n75093;
  assign n75096 = ~n75094 & ~n75095;
  assign n75097 = pi4592 & pi9040;
  assign n75098 = pi4599 & ~pi9040;
  assign n75099 = ~n75097 & ~n75098;
  assign n75100 = ~pi2316 & n75099;
  assign n75101 = pi2316 & ~n75099;
  assign n75102 = ~n75100 & ~n75101;
  assign n75103 = pi4723 & pi9040;
  assign n75104 = pi4594 & ~pi9040;
  assign n75105 = ~n75103 & ~n75104;
  assign n75106 = ~pi2327 & n75105;
  assign n75107 = pi2327 & ~n75105;
  assign n75108 = ~n75106 & ~n75107;
  assign n75109 = pi4830 & ~pi9040;
  assign n75110 = pi4975 & pi9040;
  assign n75111 = ~n75109 & ~n75110;
  assign n75112 = ~pi2305 & n75111;
  assign n75113 = pi2305 & ~n75111;
  assign n75114 = ~n75112 & ~n75113;
  assign n75115 = n75108 & n75114;
  assign n75116 = ~n75102 & n75115;
  assign n75117 = n75096 & n75116;
  assign n75118 = ~n75108 & n75114;
  assign n75119 = n75102 & n75118;
  assign n75120 = n75096 & n75119;
  assign n75121 = ~n75117 & ~n75120;
  assign n75122 = ~n75108 & ~n75114;
  assign n75123 = n75102 & n75122;
  assign n75124 = ~n75096 & n75123;
  assign n75125 = n75102 & n75115;
  assign n75126 = ~n75096 & n75125;
  assign n75127 = ~n75124 & ~n75126;
  assign n75128 = n75121 & n75127;
  assign n75129 = ~n75090 & ~n75128;
  assign n75130 = n75108 & ~n75114;
  assign n75131 = n75102 & n75130;
  assign n75132 = n75096 & n75131;
  assign n75133 = ~n75119 & ~n75132;
  assign n75134 = ~n75090 & ~n75133;
  assign n75135 = ~n75102 & n75130;
  assign n75136 = ~n75096 & n75135;
  assign n75137 = n75090 & ~n75114;
  assign n75138 = ~n75096 & n75137;
  assign n75139 = ~n75102 & ~n75108;
  assign n75140 = n75096 & n75115;
  assign n75141 = ~n75139 & ~n75140;
  assign n75142 = n75090 & ~n75141;
  assign n75143 = ~n75138 & ~n75142;
  assign n75144 = ~n75136 & n75143;
  assign n75145 = ~n75114 & n75139;
  assign n75146 = n75096 & n75145;
  assign n75147 = n75144 & ~n75146;
  assign n75148 = ~n75134 & n75147;
  assign n75149 = pi4594 & pi9040;
  assign n75150 = pi4670 & ~pi9040;
  assign n75151 = ~n75149 & ~n75150;
  assign n75152 = ~pi2312 & ~n75151;
  assign n75153 = pi2312 & n75151;
  assign n75154 = ~n75152 & ~n75153;
  assign n75155 = ~n75148 & ~n75154;
  assign n75156 = n75102 & ~n75114;
  assign n75157 = n75090 & n75096;
  assign n75158 = n75154 & n75157;
  assign n75159 = n75156 & n75158;
  assign n75160 = ~n75096 & n75102;
  assign n75161 = n75114 & n75160;
  assign n75162 = n75090 & ~n75161;
  assign n75163 = ~n75122 & ~n75156;
  assign n75164 = ~n75096 & ~n75163;
  assign n75165 = n75096 & ~n75102;
  assign n75166 = n75108 & n75165;
  assign n75167 = ~n75116 & ~n75166;
  assign n75168 = ~n75164 & n75167;
  assign n75169 = ~n75090 & n75168;
  assign n75170 = ~n75162 & ~n75169;
  assign n75171 = ~n75102 & n75118;
  assign n75172 = n75096 & n75171;
  assign n75173 = ~n75170 & ~n75172;
  assign n75174 = n75154 & ~n75173;
  assign n75175 = ~n75159 & ~n75174;
  assign n75176 = ~n75155 & n75175;
  assign n75177 = ~n75129 & n75176;
  assign n75178 = n75090 & ~n75096;
  assign n75179 = n75130 & n75178;
  assign n75180 = ~n75102 & n75179;
  assign n75181 = n75177 & ~n75180;
  assign n75182 = pi2341 & ~n75181;
  assign n75183 = ~pi2341 & ~n75180;
  assign n75184 = n75176 & n75183;
  assign n75185 = ~n75129 & n75184;
  assign po2460 = n75182 | n75185;
  assign n75187 = pi4592 & ~pi9040;
  assign n75188 = pi4663 & pi9040;
  assign n75189 = ~n75187 & ~n75188;
  assign n75190 = pi2323 & n75189;
  assign n75191 = ~pi2323 & ~n75189;
  assign n75192 = ~n75190 & ~n75191;
  assign n75193 = pi4664 & pi9040;
  assign n75194 = pi4543 & ~pi9040;
  assign n75195 = ~n75193 & ~n75194;
  assign n75196 = ~pi2315 & n75195;
  assign n75197 = pi2315 & ~n75195;
  assign n75198 = ~n75196 & ~n75197;
  assign n75199 = ~n75192 & n75198;
  assign n75200 = pi4860 & ~pi9040;
  assign n75201 = pi4823 & pi9040;
  assign n75202 = ~n75200 & ~n75201;
  assign n75203 = ~pi2291 & ~n75202;
  assign n75204 = pi2291 & ~n75200;
  assign n75205 = ~n75201 & n75204;
  assign n75206 = ~n75203 & ~n75205;
  assign n75207 = pi4600 & pi9040;
  assign n75208 = pi4728 & ~pi9040;
  assign n75209 = ~n75207 & ~n75208;
  assign n75210 = ~pi2296 & ~n75209;
  assign n75211 = pi2296 & n75209;
  assign n75212 = ~n75210 & ~n75211;
  assign n75213 = pi4543 & pi9040;
  assign n75214 = pi4872 & ~pi9040;
  assign n75215 = ~n75213 & ~n75214;
  assign n75216 = pi2310 & n75215;
  assign n75217 = ~pi2310 & ~n75215;
  assign n75218 = ~n75216 & ~n75217;
  assign n75219 = n75212 & ~n75218;
  assign n75220 = ~n75206 & n75219;
  assign n75221 = pi4860 & pi9040;
  assign n75222 = pi4663 & ~pi9040;
  assign n75223 = ~n75221 & ~n75222;
  assign n75224 = ~pi2328 & n75223;
  assign n75225 = pi2328 & ~n75223;
  assign n75226 = ~n75224 & ~n75225;
  assign n75227 = n75218 & n75226;
  assign n75228 = n75212 & n75227;
  assign n75229 = n75206 & n75228;
  assign n75230 = n75218 & ~n75226;
  assign n75231 = ~n75206 & n75230;
  assign n75232 = ~n75229 & ~n75231;
  assign n75233 = ~n75220 & n75232;
  assign n75234 = n75199 & ~n75233;
  assign n75235 = ~n75206 & ~n75212;
  assign n75236 = n75226 & n75235;
  assign n75237 = ~n75218 & n75226;
  assign n75238 = n75212 & n75237;
  assign n75239 = n75206 & n75238;
  assign n75240 = ~n75236 & ~n75239;
  assign n75241 = ~n75212 & n75227;
  assign n75242 = n75212 & n75230;
  assign n75243 = ~n75241 & ~n75242;
  assign n75244 = n75240 & n75243;
  assign n75245 = n75192 & ~n75244;
  assign n75246 = ~n75218 & ~n75226;
  assign n75247 = ~n75212 & n75246;
  assign n75248 = n75206 & n75247;
  assign n75249 = ~n75245 & ~n75248;
  assign n75250 = n75198 & ~n75249;
  assign n75251 = ~n75234 & ~n75250;
  assign n75252 = ~n75230 & ~n75237;
  assign n75253 = n75206 & ~n75252;
  assign n75254 = ~n75212 & n75237;
  assign n75255 = ~n75253 & ~n75254;
  assign n75256 = ~n75192 & ~n75255;
  assign n75257 = n75212 & n75246;
  assign n75258 = ~n75220 & ~n75257;
  assign n75259 = ~n75229 & n75258;
  assign n75260 = n75192 & ~n75259;
  assign n75261 = ~n75256 & ~n75260;
  assign n75262 = ~n75192 & ~n75206;
  assign n75263 = n75227 & n75262;
  assign n75264 = n75206 & ~n75212;
  assign n75265 = n75226 & n75264;
  assign n75266 = ~n75218 & n75265;
  assign n75267 = ~n75212 & n75218;
  assign n75268 = ~n75226 & n75267;
  assign n75269 = n75206 & n75268;
  assign n75270 = ~n75266 & ~n75269;
  assign n75271 = ~n75226 & n75235;
  assign n75272 = ~n75218 & n75271;
  assign n75273 = n75270 & ~n75272;
  assign n75274 = ~n75263 & n75273;
  assign n75275 = n75261 & n75274;
  assign n75276 = ~n75198 & ~n75275;
  assign n75277 = n75192 & ~n75206;
  assign n75278 = n75212 & n75277;
  assign n75279 = ~n75226 & n75278;
  assign n75280 = ~n75206 & n75241;
  assign n75281 = ~n75279 & ~n75280;
  assign n75282 = ~n75276 & n75281;
  assign n75283 = n75251 & n75282;
  assign n75284 = pi2336 & ~n75283;
  assign n75285 = ~pi2336 & n75281;
  assign n75286 = n75251 & n75285;
  assign n75287 = ~n75276 & n75286;
  assign po2463 = n75284 | n75287;
  assign n75289 = pi4955 & pi9040;
  assign n75290 = pi4660 & ~pi9040;
  assign n75291 = ~n75289 & ~n75290;
  assign n75292 = ~pi2310 & ~n75291;
  assign n75293 = pi2310 & n75291;
  assign n75294 = ~n75292 & ~n75293;
  assign n75295 = pi4864 & ~pi9040;
  assign n75296 = pi4727 & pi9040;
  assign n75297 = ~n75295 & ~n75296;
  assign n75298 = pi2330 & n75297;
  assign n75299 = ~pi2330 & ~n75297;
  assign n75300 = ~n75298 & ~n75299;
  assign n75301 = pi4514 & ~pi9040;
  assign n75302 = pi4728 & pi9040;
  assign n75303 = ~n75301 & ~n75302;
  assign n75304 = pi2332 & n75303;
  assign n75305 = ~pi2332 & ~n75303;
  assign n75306 = ~n75304 & ~n75305;
  assign n75307 = ~n75300 & ~n75306;
  assign n75308 = pi4667 & pi9040;
  assign n75309 = pi4538 & ~pi9040;
  assign n75310 = ~n75308 & ~n75309;
  assign n75311 = ~pi2313 & ~n75310;
  assign n75312 = pi2313 & n75310;
  assign n75313 = ~n75311 & ~n75312;
  assign n75314 = n75307 & n75313;
  assign n75315 = pi4763 & ~pi9040;
  assign n75316 = pi4598 & pi9040;
  assign n75317 = ~n75315 & ~n75316;
  assign n75318 = pi2326 & n75317;
  assign n75319 = ~pi2326 & ~n75317;
  assign n75320 = ~n75318 & ~n75319;
  assign n75321 = pi4598 & ~pi9040;
  assign n75322 = pi4872 & pi9040;
  assign n75323 = ~n75321 & ~n75322;
  assign n75324 = pi2296 & n75323;
  assign n75325 = ~pi2296 & ~n75323;
  assign n75326 = ~n75324 & ~n75325;
  assign n75327 = ~n75313 & ~n75326;
  assign n75328 = n75320 & n75327;
  assign n75329 = n75300 & n75328;
  assign n75330 = ~n75313 & n75326;
  assign n75331 = ~n75320 & n75330;
  assign n75332 = n75300 & n75331;
  assign n75333 = ~n75329 & ~n75332;
  assign n75334 = n75313 & n75326;
  assign n75335 = ~n75320 & n75334;
  assign n75336 = ~n75300 & ~n75320;
  assign n75337 = ~n75326 & n75336;
  assign n75338 = ~n75313 & n75337;
  assign n75339 = ~n75335 & ~n75338;
  assign n75340 = n75306 & ~n75339;
  assign n75341 = n75333 & ~n75340;
  assign n75342 = ~n75314 & n75341;
  assign n75343 = n75294 & ~n75342;
  assign n75344 = n75313 & ~n75326;
  assign n75345 = ~n75320 & n75344;
  assign n75346 = n75300 & n75345;
  assign n75347 = ~n75306 & n75346;
  assign n75348 = ~n75300 & n75306;
  assign n75349 = n75345 & n75348;
  assign n75350 = ~n75300 & n75320;
  assign n75351 = ~n75313 & n75350;
  assign n75352 = ~n75349 & ~n75351;
  assign n75353 = n75320 & ~n75326;
  assign n75354 = n75313 & n75353;
  assign n75355 = n75300 & n75354;
  assign n75356 = ~n75320 & n75327;
  assign n75357 = n75300 & n75356;
  assign n75358 = ~n75355 & ~n75357;
  assign n75359 = n75320 & n75330;
  assign n75360 = ~n75335 & ~n75359;
  assign n75361 = ~n75300 & n75330;
  assign n75362 = n75360 & ~n75361;
  assign n75363 = ~n75306 & ~n75362;
  assign n75364 = n75320 & n75334;
  assign n75365 = n75306 & n75364;
  assign n75366 = ~n75363 & ~n75365;
  assign n75367 = n75358 & n75366;
  assign n75368 = n75352 & n75367;
  assign n75369 = ~n75294 & ~n75368;
  assign n75370 = ~n75347 & ~n75369;
  assign n75371 = ~n75343 & n75370;
  assign n75372 = n75348 & n75359;
  assign n75373 = n75306 & n75353;
  assign n75374 = n75300 & n75373;
  assign n75375 = ~n75372 & ~n75374;
  assign n75376 = n75306 & n75332;
  assign n75377 = n75375 & ~n75376;
  assign n75378 = n75371 & n75377;
  assign n75379 = ~pi2340 & ~n75378;
  assign n75380 = pi2340 & n75377;
  assign n75381 = n75370 & n75380;
  assign n75382 = ~n75343 & n75381;
  assign po2464 = n75379 | n75382;
  assign n75384 = n74858 & n74874;
  assign n75385 = ~n74904 & ~n75384;
  assign n75386 = ~n74846 & ~n75385;
  assign n75387 = n74871 & n74884;
  assign n75388 = ~n74944 & ~n75387;
  assign n75389 = n74846 & ~n75388;
  assign n75390 = ~n74871 & n74894;
  assign n75391 = ~n74964 & ~n75390;
  assign n75392 = ~n74873 & n75391;
  assign n75393 = ~n75389 & n75392;
  assign n75394 = ~n75386 & n75393;
  assign n75395 = ~n74940 & ~n74951;
  assign n75396 = n75394 & n75395;
  assign n75397 = n74883 & ~n75396;
  assign n75398 = n74852 & n74874;
  assign n75399 = n74871 & n74890;
  assign n75400 = ~n75398 & ~n75399;
  assign n75401 = n74846 & ~n75400;
  assign n75402 = n74846 & n74884;
  assign n75403 = ~n74871 & n75402;
  assign n75404 = ~n75401 & ~n75403;
  assign n75405 = n74859 & n74938;
  assign n75406 = n74911 & ~n75405;
  assign n75407 = n74846 & ~n75406;
  assign n75408 = ~n74871 & n74901;
  assign n75409 = ~n75407 & ~n75408;
  assign n75410 = n75404 & n75409;
  assign n75411 = ~n74883 & ~n75410;
  assign n75412 = ~n74886 & ~n74894;
  assign n75413 = ~n74945 & n75412;
  assign n75414 = n74918 & ~n75413;
  assign n75415 = ~n75411 & ~n75414;
  assign n75416 = ~n74873 & ~n74940;
  assign n75417 = ~n74846 & ~n75416;
  assign n75418 = n75415 & ~n75417;
  assign n75419 = ~n75397 & n75418;
  assign n75420 = ~pi2375 & n75419;
  assign n75421 = pi2375 & ~n75419;
  assign po2470 = n75420 | n75421;
  assign n75423 = n75326 & n75350;
  assign n75424 = ~n75335 & ~n75351;
  assign n75425 = ~n75306 & ~n75424;
  assign n75426 = ~n75423 & ~n75425;
  assign n75427 = ~n75320 & ~n75326;
  assign n75428 = ~n75300 & n75427;
  assign n75429 = n75300 & n75327;
  assign n75430 = ~n75428 & ~n75429;
  assign n75431 = ~n75313 & ~n75320;
  assign n75432 = n75430 & ~n75431;
  assign n75433 = ~n75364 & n75432;
  assign n75434 = n75306 & ~n75433;
  assign n75435 = n75426 & ~n75434;
  assign n75436 = ~n75355 & n75435;
  assign n75437 = n75294 & ~n75436;
  assign n75438 = ~n75300 & n75331;
  assign n75439 = n75358 & ~n75438;
  assign n75440 = n75306 & ~n75439;
  assign n75441 = ~n75437 & ~n75440;
  assign n75442 = ~n75300 & n75364;
  assign n75443 = n75313 & ~n75320;
  assign n75444 = ~n75306 & n75443;
  assign n75445 = n75300 & n75444;
  assign n75446 = n75320 & n75348;
  assign n75447 = ~n75326 & n75446;
  assign n75448 = n75300 & n75359;
  assign n75449 = ~n75447 & ~n75448;
  assign n75450 = ~n75313 & n75320;
  assign n75451 = n75300 & n75450;
  assign n75452 = ~n75345 & ~n75451;
  assign n75453 = ~n75306 & ~n75452;
  assign n75454 = ~n75306 & ~n75313;
  assign n75455 = ~n75320 & n75454;
  assign n75456 = ~n75300 & n75455;
  assign n75457 = ~n75453 & ~n75456;
  assign n75458 = n75449 & n75457;
  assign n75459 = ~n75294 & ~n75458;
  assign n75460 = ~n75445 & ~n75459;
  assign n75461 = ~n75442 & n75460;
  assign n75462 = n75441 & n75461;
  assign n75463 = ~pi2348 & ~n75462;
  assign n75464 = ~n75437 & ~n75442;
  assign n75465 = ~n75440 & n75464;
  assign n75466 = n75460 & n75465;
  assign n75467 = pi2348 & n75466;
  assign po2471 = n75463 | n75467;
  assign n75469 = ~n75300 & n75328;
  assign n75470 = ~n75331 & ~n75442;
  assign n75471 = n75300 & n75353;
  assign n75472 = ~n75300 & n75345;
  assign n75473 = ~n75471 & ~n75472;
  assign n75474 = n75470 & n75473;
  assign n75475 = ~n75306 & ~n75474;
  assign n75476 = n75300 & n75334;
  assign n75477 = ~n75351 & ~n75476;
  assign n75478 = ~n75356 & n75477;
  assign n75479 = n75306 & ~n75478;
  assign n75480 = n75300 & ~n75320;
  assign n75481 = n75326 & n75480;
  assign n75482 = n75313 & n75481;
  assign n75483 = ~n75479 & ~n75482;
  assign n75484 = ~n75475 & n75483;
  assign n75485 = ~n75469 & n75484;
  assign n75486 = ~n75294 & ~n75485;
  assign n75487 = n75300 & ~n75306;
  assign n75488 = n75364 & n75487;
  assign n75489 = ~n75306 & n75356;
  assign n75490 = ~n75306 & n75359;
  assign n75491 = ~n75489 & ~n75490;
  assign n75492 = ~n75300 & ~n75491;
  assign n75493 = ~n75488 & ~n75492;
  assign n75494 = n75300 & n75330;
  assign n75495 = ~n75300 & n75334;
  assign n75496 = ~n75494 & ~n75495;
  assign n75497 = ~n75354 & n75496;
  assign n75498 = ~n75331 & n75497;
  assign n75499 = n75306 & ~n75498;
  assign n75500 = ~n75300 & n75335;
  assign n75501 = ~n75499 & ~n75500;
  assign n75502 = ~n75300 & n75354;
  assign n75503 = ~n75346 & ~n75502;
  assign n75504 = n75501 & n75503;
  assign n75505 = n75493 & n75504;
  assign n75506 = n75294 & ~n75505;
  assign n75507 = ~n75306 & ~n75333;
  assign n75508 = ~n75506 & ~n75507;
  assign n75509 = ~n75357 & ~n75502;
  assign n75510 = n75306 & ~n75509;
  assign n75511 = n75508 & ~n75510;
  assign n75512 = ~n75486 & n75511;
  assign n75513 = pi2353 & ~n75512;
  assign n75514 = ~pi2353 & n75512;
  assign po2475 = n75513 | n75514;
  assign n75516 = n75192 & n75230;
  assign n75517 = ~n75206 & n75516;
  assign n75518 = ~n75206 & n75212;
  assign n75519 = n75226 & n75518;
  assign n75520 = ~n75218 & n75519;
  assign n75521 = ~n75517 & ~n75520;
  assign n75522 = n75206 & ~n75226;
  assign n75523 = n75212 & n75522;
  assign n75524 = ~n75206 & ~n75218;
  assign n75525 = ~n75519 & ~n75524;
  assign n75526 = ~n75192 & ~n75525;
  assign n75527 = ~n75523 & ~n75526;
  assign n75528 = n75521 & n75527;
  assign n75529 = ~n75198 & ~n75528;
  assign n75530 = ~n75228 & ~n75269;
  assign n75531 = ~n75206 & n75246;
  assign n75532 = n75530 & ~n75531;
  assign n75533 = n75192 & ~n75532;
  assign n75534 = n75230 & n75262;
  assign n75535 = ~n75280 & ~n75534;
  assign n75536 = ~n75533 & n75535;
  assign n75537 = ~n75238 & ~n75248;
  assign n75538 = ~n75192 & ~n75537;
  assign n75539 = n75536 & ~n75538;
  assign n75540 = n75198 & ~n75539;
  assign n75541 = ~n75529 & ~n75540;
  assign n75542 = ~n75206 & n75237;
  assign n75543 = n75206 & ~n75243;
  assign n75544 = ~n75542 & ~n75543;
  assign n75545 = ~n75192 & ~n75544;
  assign n75546 = n75192 & n75206;
  assign n75547 = ~n75254 & ~n75257;
  assign n75548 = ~n75228 & n75547;
  assign n75549 = n75546 & ~n75548;
  assign n75550 = ~n75545 & ~n75549;
  assign n75551 = n75541 & n75550;
  assign n75552 = ~pi2337 & ~n75551;
  assign n75553 = ~n75529 & n75550;
  assign n75554 = ~n75540 & n75553;
  assign n75555 = pi2337 & n75554;
  assign po2476 = n75552 | n75555;
  assign n75557 = ~n75192 & ~n75547;
  assign n75558 = n75206 & n75242;
  assign n75559 = ~n75557 & ~n75558;
  assign n75560 = n75206 & n75218;
  assign n75561 = ~n75267 & ~n75560;
  assign n75562 = ~n75238 & n75561;
  assign n75563 = n75192 & ~n75562;
  assign n75564 = n75559 & ~n75563;
  assign n75565 = n75198 & ~n75564;
  assign n75566 = ~n75206 & n75268;
  assign n75567 = ~n75192 & n75566;
  assign n75568 = ~n75206 & n75228;
  assign n75569 = ~n75192 & n75568;
  assign n75570 = ~n75567 & ~n75569;
  assign n75571 = n75192 & n75272;
  assign n75572 = n75570 & ~n75571;
  assign n75573 = n75192 & ~n75212;
  assign n75574 = ~n75226 & n75573;
  assign n75575 = ~n75218 & n75574;
  assign n75576 = ~n75272 & ~n75519;
  assign n75577 = ~n75206 & n75218;
  assign n75578 = n75212 & n75577;
  assign n75579 = n75192 & n75578;
  assign n75580 = n75206 & n75257;
  assign n75581 = ~n75192 & n75267;
  assign n75582 = ~n75580 & ~n75581;
  assign n75583 = ~n75266 & n75582;
  assign n75584 = ~n75579 & n75583;
  assign n75585 = n75576 & n75584;
  assign n75586 = ~n75575 & n75585;
  assign n75587 = ~n75198 & ~n75586;
  assign n75588 = n75572 & ~n75587;
  assign n75589 = ~n75565 & n75588;
  assign n75590 = ~pi2339 & ~n75589;
  assign n75591 = pi2339 & n75572;
  assign n75592 = ~n75565 & n75591;
  assign n75593 = ~n75587 & n75592;
  assign po2477 = n75590 | n75593;
  assign n75595 = n75206 & n75219;
  assign n75596 = ~n75242 & ~n75595;
  assign n75597 = ~n75280 & n75596;
  assign n75598 = n75192 & ~n75597;
  assign n75599 = ~n75212 & ~n75218;
  assign n75600 = ~n75227 & ~n75599;
  assign n75601 = n75206 & ~n75600;
  assign n75602 = ~n75206 & n75257;
  assign n75603 = ~n75601 & ~n75602;
  assign n75604 = ~n75566 & n75603;
  assign n75605 = ~n75192 & ~n75604;
  assign n75606 = ~n75598 & ~n75605;
  assign n75607 = ~n75198 & ~n75606;
  assign n75608 = ~n75218 & n75277;
  assign n75609 = ~n75578 & ~n75595;
  assign n75610 = ~n75192 & ~n75609;
  assign n75611 = ~n75263 & ~n75610;
  assign n75612 = ~n75269 & ~n75568;
  assign n75613 = n75267 & n75546;
  assign n75614 = ~n75575 & ~n75613;
  assign n75615 = n75612 & n75614;
  assign n75616 = n75611 & n75615;
  assign n75617 = ~n75608 & n75616;
  assign n75618 = n75198 & ~n75617;
  assign n75619 = ~n75192 & n75254;
  assign n75620 = ~n75206 & n75619;
  assign n75621 = ~n75569 & ~n75620;
  assign n75622 = ~n75571 & n75621;
  assign n75623 = n75206 & n75230;
  assign n75624 = ~n75520 & ~n75623;
  assign n75625 = n75192 & ~n75624;
  assign n75626 = n75622 & ~n75625;
  assign n75627 = ~n75618 & n75626;
  assign n75628 = ~n75607 & n75627;
  assign n75629 = ~pi2338 & n75628;
  assign n75630 = pi2338 & ~n75628;
  assign po2481 = n75629 | n75630;
  assign n75632 = n74987 & ~n75025;
  assign n75633 = n75005 & n75015;
  assign n75634 = n74999 & ~n75011;
  assign n75635 = ~n75633 & ~n75634;
  assign n75636 = n75632 & ~n75635;
  assign n75637 = ~n75028 & ~n75034;
  assign n75638 = ~n75026 & n75058;
  assign n75639 = ~n74999 & n75638;
  assign n75640 = ~n75031 & ~n75639;
  assign n75641 = n75637 & n75640;
  assign n75642 = ~n75025 & ~n75641;
  assign n75643 = n74993 & n75069;
  assign n75644 = n74993 & n75064;
  assign n75645 = ~n75643 & ~n75644;
  assign n75646 = n74987 & ~n75645;
  assign n75647 = n74999 & n75029;
  assign n75648 = n74987 & n75647;
  assign n75649 = n74993 & n75648;
  assign n75650 = ~n75646 & ~n75649;
  assign n75651 = ~n74987 & n75028;
  assign n75652 = n75650 & ~n75651;
  assign n75653 = ~n75642 & n75652;
  assign n75654 = ~n75636 & n75653;
  assign n75655 = ~n74987 & n75026;
  assign n75656 = ~n74993 & n75655;
  assign n75657 = ~n74993 & n75027;
  assign n75658 = n74999 & n75026;
  assign n75659 = n74993 & n75658;
  assign n75660 = ~n74993 & n75063;
  assign n75661 = ~n75659 & ~n75660;
  assign n75662 = n74987 & ~n75661;
  assign n75663 = ~n75657 & ~n75662;
  assign n75664 = ~n74993 & n75030;
  assign n75665 = ~n75643 & ~n75664;
  assign n75666 = ~n75061 & n75665;
  assign n75667 = n75663 & n75666;
  assign n75668 = ~n75656 & n75667;
  assign n75669 = n75025 & ~n75668;
  assign n75670 = n75654 & ~n75669;
  assign n75671 = ~n74987 & n74993;
  assign n75672 = n75066 & n75671;
  assign n75673 = n75670 & ~n75672;
  assign n75674 = pi2345 & n75673;
  assign n75675 = ~pi2345 & ~n75673;
  assign po2482 = n75674 | n75675;
  assign n75677 = n74993 & n75655;
  assign n75678 = ~n75005 & n75015;
  assign n75679 = ~n75647 & ~n75678;
  assign n75680 = ~n74987 & ~n75679;
  assign n75681 = ~n75677 & ~n75680;
  assign n75682 = n74987 & n75063;
  assign n75683 = n74993 & n75682;
  assign n75684 = n74987 & n75013;
  assign n75685 = ~n75683 & ~n75684;
  assign n75686 = n75681 & n75685;
  assign n75687 = ~n75005 & n75035;
  assign n75688 = ~n75014 & ~n75687;
  assign n75689 = ~n75070 & n75688;
  assign n75690 = n75686 & n75689;
  assign n75691 = ~n75025 & ~n75690;
  assign n75692 = ~n75028 & ~n75647;
  assign n75693 = ~n75072 & n75692;
  assign n75694 = n74987 & ~n75693;
  assign n75695 = ~n74993 & n75658;
  assign n75696 = ~n75044 & ~n75695;
  assign n75697 = ~n75672 & n75696;
  assign n75698 = ~n74987 & n75069;
  assign n75699 = n75697 & ~n75698;
  assign n75700 = ~n75694 & n75699;
  assign n75701 = n75025 & ~n75700;
  assign n75702 = ~n75054 & ~n75060;
  assign n75703 = ~n75014 & n75696;
  assign n75704 = n74987 & ~n75703;
  assign n75705 = n75702 & ~n75704;
  assign n75706 = ~n75701 & n75705;
  assign n75707 = ~n75691 & n75706;
  assign n75708 = pi2350 & ~n75707;
  assign n75709 = ~pi2350 & n75707;
  assign po2483 = n75708 | n75709;
  assign n75711 = ~n75633 & ~n75664;
  assign n75712 = n75025 & ~n75711;
  assign n75713 = n75011 & n75035;
  assign n75714 = ~n75036 & ~n75713;
  assign n75715 = ~n75027 & n75714;
  assign n75716 = n74987 & ~n75715;
  assign n75717 = n75025 & n75716;
  assign n75718 = ~n75712 & ~n75717;
  assign n75719 = n74987 & ~n74993;
  assign n75720 = n75030 & n75719;
  assign n75721 = ~n75041 & ~n75720;
  assign n75722 = ~n75034 & ~n75073;
  assign n75723 = ~n74987 & ~n75722;
  assign n75724 = n75025 & n75723;
  assign n75725 = n75721 & ~n75724;
  assign n75726 = ~n75011 & n75035;
  assign n75727 = ~n75005 & n75726;
  assign n75728 = n74993 & n75012;
  assign n75729 = ~n75017 & ~n75728;
  assign n75730 = ~n74987 & ~n75729;
  assign n75731 = ~n75028 & ~n75044;
  assign n75732 = n74993 & n75029;
  assign n75733 = ~n75066 & ~n75732;
  assign n75734 = n74987 & ~n75733;
  assign n75735 = n75731 & ~n75734;
  assign n75736 = ~n75730 & n75735;
  assign n75737 = ~n75727 & n75736;
  assign n75738 = ~n75025 & ~n75737;
  assign n75739 = ~n75070 & n75696;
  assign n75740 = ~n74987 & ~n75739;
  assign n75741 = ~n75738 & ~n75740;
  assign n75742 = n75725 & n75741;
  assign n75743 = n75718 & n75742;
  assign n75744 = ~pi2362 & ~n75743;
  assign n75745 = pi2362 & n75725;
  assign n75746 = n75718 & n75745;
  assign n75747 = n75741 & n75746;
  assign po2484 = n75744 | n75747;
  assign n75749 = ~n75338 & ~n75502;
  assign n75750 = ~n75482 & n75749;
  assign n75751 = ~n75306 & ~n75750;
  assign n75752 = ~n75346 & ~n75490;
  assign n75753 = ~n75328 & ~n75495;
  assign n75754 = n75306 & ~n75753;
  assign n75755 = ~n75442 & ~n75754;
  assign n75756 = n75752 & n75755;
  assign n75757 = n75294 & ~n75756;
  assign n75758 = ~n75320 & n75326;
  assign n75759 = ~n75431 & ~n75758;
  assign n75760 = n75300 & ~n75759;
  assign n75761 = ~n75354 & ~n75361;
  assign n75762 = n75306 & ~n75761;
  assign n75763 = n75300 & n75326;
  assign n75764 = ~n75335 & ~n75763;
  assign n75765 = ~n75327 & n75764;
  assign n75766 = ~n75306 & ~n75765;
  assign n75767 = ~n75762 & ~n75766;
  assign n75768 = ~n75760 & n75767;
  assign n75769 = ~n75294 & ~n75768;
  assign n75770 = ~n75757 & ~n75769;
  assign n75771 = ~n75349 & ~n75376;
  assign n75772 = n75770 & n75771;
  assign n75773 = ~n75751 & n75772;
  assign n75774 = ~pi2359 & ~n75773;
  assign n75775 = pi2359 & n75771;
  assign n75776 = ~n75751 & n75775;
  assign n75777 = n75770 & n75776;
  assign po2485 = n75774 | n75777;
  assign n75779 = pi4667 & ~pi9040;
  assign n75780 = pi4660 & pi9040;
  assign n75781 = ~n75779 & ~n75780;
  assign n75782 = ~pi2315 & n75781;
  assign n75783 = pi2315 & ~n75781;
  assign n75784 = ~n75782 & ~n75783;
  assign n75785 = pi4668 & ~pi9040;
  assign n75786 = pi4858 & pi9040;
  assign n75787 = ~n75785 & ~n75786;
  assign n75788 = ~pi2316 & n75787;
  assign n75789 = pi2316 & ~n75787;
  assign n75790 = ~n75788 & ~n75789;
  assign n75791 = pi4541 & ~pi9040;
  assign n75792 = pi4599 & pi9040;
  assign n75793 = ~n75791 & ~n75792;
  assign n75794 = ~pi2301 & n75793;
  assign n75795 = pi2301 & ~n75793;
  assign n75796 = ~n75794 & ~n75795;
  assign n75797 = pi4763 & pi9040;
  assign n75798 = pi4975 & ~pi9040;
  assign n75799 = ~n75797 & ~n75798;
  assign n75800 = ~pi2328 & ~n75799;
  assign n75801 = pi2328 & n75799;
  assign n75802 = ~n75800 & ~n75801;
  assign n75803 = n75796 & ~n75802;
  assign n75804 = ~n75790 & n75803;
  assign n75805 = ~n75784 & n75804;
  assign n75806 = ~n75784 & n75790;
  assign n75807 = ~n75802 & n75806;
  assign n75808 = ~n75796 & n75807;
  assign n75809 = pi4864 & pi9040;
  assign n75810 = pi4858 & ~pi9040;
  assign n75811 = ~n75809 & ~n75810;
  assign n75812 = ~pi2307 & ~n75811;
  assign n75813 = pi2307 & n75811;
  assign n75814 = ~n75812 & ~n75813;
  assign n75815 = n75790 & n75803;
  assign n75816 = n75784 & n75815;
  assign n75817 = ~n75784 & n75802;
  assign n75818 = ~n75816 & ~n75817;
  assign n75819 = n75814 & ~n75818;
  assign n75820 = ~n75808 & ~n75819;
  assign n75821 = ~n75805 & n75820;
  assign n75822 = ~n75796 & n75802;
  assign n75823 = n75790 & n75822;
  assign n75824 = n75784 & n75823;
  assign n75825 = n75784 & ~n75790;
  assign n75826 = n75802 & n75825;
  assign n75827 = n75796 & n75826;
  assign n75828 = ~n75802 & n75825;
  assign n75829 = ~n75796 & n75828;
  assign n75830 = ~n75814 & n75829;
  assign n75831 = ~n75827 & ~n75830;
  assign n75832 = ~n75824 & n75831;
  assign n75833 = n75821 & n75832;
  assign n75834 = pi4727 & ~pi9040;
  assign n75835 = pi4514 & pi9040;
  assign n75836 = ~n75834 & ~n75835;
  assign n75837 = ~pi2305 & ~n75836;
  assign n75838 = pi2305 & n75836;
  assign n75839 = ~n75837 & ~n75838;
  assign n75840 = ~n75833 & n75839;
  assign n75841 = ~n75784 & ~n75790;
  assign n75842 = ~n75802 & n75841;
  assign n75843 = ~n75796 & n75842;
  assign n75844 = ~n75796 & ~n75802;
  assign n75845 = n75790 & n75844;
  assign n75846 = n75784 & n75845;
  assign n75847 = ~n75843 & ~n75846;
  assign n75848 = n75814 & n75828;
  assign n75849 = ~n75796 & n75826;
  assign n75850 = ~n75848 & ~n75849;
  assign n75851 = n75796 & n75807;
  assign n75852 = n75784 & n75790;
  assign n75853 = n75802 & n75852;
  assign n75854 = n75796 & n75853;
  assign n75855 = ~n75851 & ~n75854;
  assign n75856 = ~n75790 & n75802;
  assign n75857 = ~n75784 & ~n75796;
  assign n75858 = ~n75856 & ~n75857;
  assign n75859 = n75790 & ~n75802;
  assign n75860 = n75858 & ~n75859;
  assign n75861 = ~n75814 & ~n75860;
  assign n75862 = n75855 & ~n75861;
  assign n75863 = n75850 & n75862;
  assign n75864 = n75847 & n75863;
  assign n75865 = ~n75839 & ~n75864;
  assign n75866 = ~n75840 & ~n75865;
  assign n75867 = pi2344 & ~n75866;
  assign n75868 = ~pi2344 & ~n75840;
  assign n75869 = ~n75865 & n75868;
  assign po2488 = n75867 | n75869;
  assign n75871 = ~n74871 & n74890;
  assign n75872 = ~n74889 & ~n75871;
  assign n75873 = ~n74846 & ~n75872;
  assign n75874 = n74846 & ~n74966;
  assign n75875 = ~n74955 & ~n75874;
  assign n75876 = ~n75873 & n75875;
  assign n75877 = n74883 & ~n75876;
  assign n75878 = ~n74846 & n74901;
  assign n75879 = ~n75877 & ~n75878;
  assign n75880 = ~n75390 & ~n75399;
  assign n75881 = n74846 & ~n75880;
  assign n75882 = n74846 & n74891;
  assign n75883 = n74871 & n74904;
  assign n75884 = ~n74846 & n74872;
  assign n75885 = ~n74943 & ~n75884;
  assign n75886 = ~n74852 & ~n75885;
  assign n75887 = ~n74944 & ~n75886;
  assign n75888 = ~n74873 & n75887;
  assign n75889 = ~n75883 & n75888;
  assign n75890 = ~n75882 & n75889;
  assign n75891 = ~n74883 & ~n75890;
  assign n75892 = ~n75881 & ~n75891;
  assign n75893 = n75879 & n75892;
  assign n75894 = pi2382 & ~n75893;
  assign n75895 = ~pi2382 & n75893;
  assign po2491 = n75894 | n75895;
  assign n75897 = ~n75096 & n75145;
  assign n75898 = n75096 & n75156;
  assign n75899 = ~n75135 & ~n75898;
  assign n75900 = ~n75090 & ~n75899;
  assign n75901 = ~n75897 & ~n75900;
  assign n75902 = ~n75114 & n75178;
  assign n75903 = ~n75108 & n75902;
  assign n75904 = n75118 & n75157;
  assign n75905 = ~n75903 & ~n75904;
  assign n75906 = n75090 & n75115;
  assign n75907 = ~n75102 & n75906;
  assign n75908 = n75905 & ~n75907;
  assign n75909 = ~n75126 & ~n75132;
  assign n75910 = n75114 & n75165;
  assign n75911 = n75909 & ~n75910;
  assign n75912 = n75908 & n75911;
  assign n75913 = n75901 & n75912;
  assign n75914 = ~n75154 & ~n75913;
  assign n75915 = ~n75125 & ~n75135;
  assign n75916 = n75096 & ~n75915;
  assign n75917 = ~n75108 & n75160;
  assign n75918 = ~n75171 & ~n75917;
  assign n75919 = ~n75102 & ~n75114;
  assign n75920 = n75096 & n75919;
  assign n75921 = n75918 & ~n75920;
  assign n75922 = ~n75090 & ~n75921;
  assign n75923 = ~n75096 & n75130;
  assign n75924 = n75096 & n75102;
  assign n75925 = ~n75114 & n75924;
  assign n75926 = ~n75108 & n75925;
  assign n75927 = ~n75923 & ~n75926;
  assign n75928 = n75090 & ~n75927;
  assign n75929 = ~n75096 & n75119;
  assign n75930 = ~n75928 & ~n75929;
  assign n75931 = ~n75922 & n75930;
  assign n75932 = ~n75916 & n75931;
  assign n75933 = n75154 & ~n75932;
  assign n75934 = ~n75090 & n75161;
  assign n75935 = ~n75933 & ~n75934;
  assign n75936 = n75139 & n75178;
  assign n75937 = ~n75114 & n75936;
  assign n75938 = n75935 & ~n75937;
  assign n75939 = ~n75914 & n75938;
  assign n75940 = ~pi2351 & ~n75939;
  assign n75941 = pi2351 & n75935;
  assign n75942 = ~n75914 & n75941;
  assign n75943 = ~n75937 & n75942;
  assign po2492 = n75940 | n75943;
  assign n75945 = ~n75117 & ~n75124;
  assign n75946 = n75090 & ~n75945;
  assign n75947 = ~n75180 & ~n75946;
  assign n75948 = n75090 & n75122;
  assign n75949 = n75096 & n75948;
  assign n75950 = ~n75907 & ~n75949;
  assign n75951 = n75102 & n75108;
  assign n75952 = n75096 & n75130;
  assign n75953 = ~n75951 & ~n75952;
  assign n75954 = ~n75096 & ~n75102;
  assign n75955 = ~n75108 & n75954;
  assign n75956 = n75953 & ~n75955;
  assign n75957 = ~n75090 & ~n75956;
  assign n75958 = ~n75120 & ~n75957;
  assign n75959 = n75950 & n75958;
  assign n75960 = ~n75154 & ~n75959;
  assign n75961 = ~n75090 & n75951;
  assign n75962 = n75096 & n75961;
  assign n75963 = ~n75960 & ~n75962;
  assign n75964 = ~n75135 & ~n75161;
  assign n75965 = ~n75171 & n75964;
  assign n75966 = n75090 & ~n75965;
  assign n75967 = ~n75096 & n75116;
  assign n75968 = ~n75145 & ~n75967;
  assign n75969 = ~n75090 & ~n75968;
  assign n75970 = ~n75917 & ~n75969;
  assign n75971 = ~n75966 & n75970;
  assign n75972 = ~n75132 & ~n75172;
  assign n75973 = n75971 & n75972;
  assign n75974 = n75154 & ~n75973;
  assign n75975 = n75963 & ~n75974;
  assign n75976 = n75947 & n75975;
  assign n75977 = pi2374 & n75976;
  assign n75978 = ~pi2374 & ~n75976;
  assign po2493 = n75977 | n75978;
  assign n75980 = pi4724 & pi9040;
  assign n75981 = pi4544 & ~pi9040;
  assign n75982 = ~n75980 & ~n75981;
  assign n75983 = ~pi2325 & n75982;
  assign n75984 = pi2325 & ~n75982;
  assign n75985 = ~n75983 & ~n75984;
  assign n75986 = pi4726 & pi9040;
  assign n75987 = pi4674 & ~pi9040;
  assign n75988 = ~n75986 & ~n75987;
  assign n75989 = ~pi2318 & n75988;
  assign n75990 = pi2318 & ~n75988;
  assign n75991 = ~n75989 & ~n75990;
  assign n75992 = pi4669 & pi9040;
  assign n75993 = pi4950 & ~pi9040;
  assign n75994 = ~n75992 & ~n75993;
  assign n75995 = pi2334 & n75994;
  assign n75996 = ~pi2334 & ~n75994;
  assign n75997 = ~n75995 & ~n75996;
  assign n75998 = pi4614 & pi9040;
  assign n75999 = pi4659 & ~pi9040;
  assign n76000 = ~n75998 & ~n75999;
  assign n76001 = ~pi2329 & ~n76000;
  assign n76002 = pi2329 & n76000;
  assign n76003 = ~n76001 & ~n76002;
  assign n76004 = n75997 & ~n76003;
  assign n76005 = n75991 & n76004;
  assign n76006 = ~n75985 & n76005;
  assign n76007 = pi4969 & pi9040;
  assign n76008 = pi4669 & ~pi9040;
  assign n76009 = ~n76007 & ~n76008;
  assign n76010 = ~pi2295 & n76009;
  assign n76011 = pi2295 & ~n76009;
  assign n76012 = ~n76010 & ~n76011;
  assign n76013 = pi4658 & ~pi9040;
  assign n76014 = pi4672 & pi9040;
  assign n76015 = ~n76013 & ~n76014;
  assign n76016 = ~pi2320 & n76015;
  assign n76017 = pi2320 & ~n76015;
  assign n76018 = ~n76016 & ~n76017;
  assign n76019 = n75997 & ~n76018;
  assign n76020 = n76003 & n76019;
  assign n76021 = ~n75997 & ~n76018;
  assign n76022 = ~n76003 & n76021;
  assign n76023 = ~n75997 & n76018;
  assign n76024 = n75985 & n76023;
  assign n76025 = ~n76022 & ~n76024;
  assign n76026 = ~n76020 & n76025;
  assign n76027 = n75991 & ~n76026;
  assign n76028 = n76003 & n76021;
  assign n76029 = ~n76003 & n76019;
  assign n76030 = ~n76028 & ~n76029;
  assign n76031 = ~n75991 & ~n76030;
  assign n76032 = ~n76027 & ~n76031;
  assign n76033 = n75997 & n76018;
  assign n76034 = n76003 & n76033;
  assign n76035 = ~n75991 & n76034;
  assign n76036 = ~n76003 & n76024;
  assign n76037 = ~n76035 & ~n76036;
  assign n76038 = n76032 & n76037;
  assign n76039 = n76012 & ~n76038;
  assign n76040 = ~n75985 & n76028;
  assign n76041 = n75985 & n76033;
  assign n76042 = ~n75985 & n76023;
  assign n76043 = ~n76041 & ~n76042;
  assign n76044 = n75991 & ~n76043;
  assign n76045 = ~n76040 & ~n76044;
  assign n76046 = n76003 & n76023;
  assign n76047 = ~n75991 & n76046;
  assign n76048 = ~n76003 & n76033;
  assign n76049 = ~n76020 & ~n76048;
  assign n76050 = ~n76047 & n76049;
  assign n76051 = ~n76022 & n76050;
  assign n76052 = n75985 & ~n76051;
  assign n76053 = n76045 & ~n76052;
  assign n76054 = ~n76012 & ~n76053;
  assign n76055 = ~n76039 & ~n76054;
  assign n76056 = ~n76006 & n76055;
  assign n76057 = ~n75985 & n76003;
  assign n76058 = n76018 & n76057;
  assign n76059 = n75997 & n76058;
  assign n76060 = ~n76003 & n76042;
  assign n76061 = ~n76059 & ~n76060;
  assign n76062 = ~n75991 & ~n76061;
  assign n76063 = n76056 & ~n76062;
  assign n76064 = ~pi2372 & ~n76063;
  assign n76065 = pi2372 & ~n76062;
  assign n76066 = n76055 & n76065;
  assign n76067 = ~n76006 & n76066;
  assign po2494 = n76064 | n76067;
  assign n76069 = n75985 & n76021;
  assign n76070 = ~n76042 & ~n76069;
  assign n76071 = ~n75991 & ~n76070;
  assign n76072 = n75985 & n76048;
  assign n76073 = ~n75991 & n76072;
  assign n76074 = ~n76071 & ~n76073;
  assign n76075 = ~n76012 & ~n76074;
  assign n76076 = n75985 & ~n76003;
  assign n76077 = ~n76019 & ~n76023;
  assign n76078 = n76076 & ~n76077;
  assign n76079 = ~n76004 & ~n76019;
  assign n76080 = n75985 & ~n76079;
  assign n76081 = ~n76028 & ~n76080;
  assign n76082 = n75991 & ~n76081;
  assign n76083 = ~n76078 & ~n76082;
  assign n76084 = ~n75985 & n76022;
  assign n76085 = n75985 & n76003;
  assign n76086 = n76018 & n76085;
  assign n76087 = ~n75985 & ~n76079;
  assign n76088 = ~n76086 & ~n76087;
  assign n76089 = ~n75991 & ~n76088;
  assign n76090 = ~n76084 & ~n76089;
  assign n76091 = n76083 & n76090;
  assign n76092 = n76012 & ~n76091;
  assign n76093 = ~n76019 & n76057;
  assign n76094 = ~n76012 & n76093;
  assign n76095 = ~n75985 & ~n76003;
  assign n76096 = ~n75991 & n76095;
  assign n76097 = n76019 & n76096;
  assign n76098 = ~n75985 & n75991;
  assign n76099 = n76003 & n76018;
  assign n76100 = n76098 & n76099;
  assign n76101 = ~n76097 & ~n76100;
  assign n76102 = ~n76094 & n76101;
  assign n76103 = ~n75985 & n75997;
  assign n76104 = ~n76046 & ~n76103;
  assign n76105 = n75991 & ~n76012;
  assign n76106 = ~n76104 & n76105;
  assign n76107 = n76102 & ~n76106;
  assign n76108 = ~n76092 & n76107;
  assign n76109 = ~n76075 & n76108;
  assign n76110 = pi2358 & ~n76109;
  assign n76111 = ~pi2358 & n76109;
  assign po2495 = n76110 | n76111;
  assign n76113 = ~n75991 & n76028;
  assign n76114 = n75985 & n76113;
  assign n76115 = ~n76073 & ~n76114;
  assign n76116 = n75985 & n75991;
  assign n76117 = n76021 & n76116;
  assign n76118 = ~n76003 & n76117;
  assign n76119 = ~n76072 & ~n76118;
  assign n76120 = n75997 & n76003;
  assign n76121 = ~n75985 & n76120;
  assign n76122 = ~n75985 & n76021;
  assign n76123 = ~n76121 & ~n76122;
  assign n76124 = ~n75991 & ~n76123;
  assign n76125 = n75991 & ~n76076;
  assign n76126 = ~n76077 & n76125;
  assign n76127 = n75985 & ~n75991;
  assign n76128 = ~n76021 & n76127;
  assign n76129 = ~n76003 & n76128;
  assign n76130 = ~n76126 & ~n76129;
  assign n76131 = ~n76124 & n76130;
  assign n76132 = n76119 & n76131;
  assign n76133 = ~n76012 & ~n76132;
  assign n76134 = n76115 & ~n76133;
  assign n76135 = n75991 & n76020;
  assign n76136 = ~n75985 & n76135;
  assign n76137 = n75991 & n76012;
  assign n76138 = ~n76034 & ~n76122;
  assign n76139 = ~n76078 & n76138;
  assign n76140 = n76137 & ~n76139;
  assign n76141 = ~n75985 & n76048;
  assign n76142 = ~n76003 & n76103;
  assign n76143 = ~n76042 & ~n76142;
  assign n76144 = ~n76046 & ~n76069;
  assign n76145 = n76143 & n76144;
  assign n76146 = ~n75991 & ~n76145;
  assign n76147 = ~n76141 & ~n76146;
  assign n76148 = n76012 & ~n76147;
  assign n76149 = ~n76140 & ~n76148;
  assign n76150 = ~n76136 & n76149;
  assign n76151 = n76134 & n76150;
  assign n76152 = pi2356 & ~n76151;
  assign n76153 = ~pi2356 & n76134;
  assign n76154 = n76150 & n76153;
  assign po2496 = n76152 | n76154;
  assign n76156 = ~n76018 & n76085;
  assign n76157 = n76049 & ~n76156;
  assign n76158 = n76105 & ~n76157;
  assign n76159 = ~n76012 & n76046;
  assign n76160 = ~n75985 & n76159;
  assign n76161 = ~n76003 & ~n76018;
  assign n76162 = ~n76122 & ~n76161;
  assign n76163 = ~n75991 & ~n76162;
  assign n76164 = ~n76035 & ~n76163;
  assign n76165 = ~n76012 & ~n76164;
  assign n76166 = ~n76160 & ~n76165;
  assign n76167 = ~n76018 & n76095;
  assign n76168 = ~n76036 & ~n76167;
  assign n76169 = ~n75991 & ~n76168;
  assign n76170 = n76166 & ~n76169;
  assign n76171 = n76021 & n76098;
  assign n76172 = n76003 & n76171;
  assign n76173 = ~n76077 & n76095;
  assign n76174 = ~n76172 & ~n76173;
  assign n76175 = ~n76059 & n76174;
  assign n76176 = ~n76077 & n76085;
  assign n76177 = ~n76072 & ~n76176;
  assign n76178 = ~n75991 & n76085;
  assign n76179 = ~n75997 & n76178;
  assign n76180 = ~n76118 & ~n76179;
  assign n76181 = n76177 & n76180;
  assign n76182 = n76175 & n76181;
  assign n76183 = n76012 & ~n76182;
  assign n76184 = n76170 & ~n76183;
  assign n76185 = ~n76158 & n76184;
  assign n76186 = ~pi2369 & ~n76185;
  assign n76187 = pi2369 & n76170;
  assign n76188 = ~n76158 & n76187;
  assign n76189 = ~n76183 & n76188;
  assign po2497 = n76186 | n76189;
  assign n76191 = n75784 & n75802;
  assign n76192 = n75796 & n76191;
  assign n76193 = ~n75796 & n75817;
  assign n76194 = ~n76192 & ~n76193;
  assign n76195 = ~n75814 & ~n76194;
  assign n76196 = ~n75824 & ~n75829;
  assign n76197 = ~n75807 & n76196;
  assign n76198 = n75814 & ~n76197;
  assign n76199 = ~n76195 & ~n76198;
  assign n76200 = ~n75805 & ~n75826;
  assign n76201 = ~n75814 & ~n76200;
  assign n76202 = ~n75816 & ~n75829;
  assign n76203 = ~n75784 & n75844;
  assign n76204 = n75802 & n75841;
  assign n76205 = n75796 & n76204;
  assign n76206 = ~n76203 & ~n76205;
  assign n76207 = n75814 & ~n76206;
  assign n76208 = n76202 & ~n76207;
  assign n76209 = ~n76201 & n76208;
  assign n76210 = n75839 & ~n76209;
  assign n76211 = ~n75814 & n75825;
  assign n76212 = n75796 & n76211;
  assign n76213 = n75802 & n75806;
  assign n76214 = ~n75846 & ~n76213;
  assign n76215 = ~n75796 & n75841;
  assign n76216 = n76214 & ~n76215;
  assign n76217 = ~n75814 & ~n76216;
  assign n76218 = ~n75784 & ~n75802;
  assign n76219 = n75796 & n75814;
  assign n76220 = n76218 & n76219;
  assign n76221 = ~n75851 & ~n76220;
  assign n76222 = ~n76217 & n76221;
  assign n76223 = ~n76212 & n76222;
  assign n76224 = ~n75796 & n76204;
  assign n76225 = ~n75827 & ~n76224;
  assign n76226 = n76223 & n76225;
  assign n76227 = ~n75839 & ~n76226;
  assign n76228 = n75814 & n75859;
  assign n76229 = n75796 & n76228;
  assign n76230 = ~n76227 & ~n76229;
  assign n76231 = ~n76210 & n76230;
  assign n76232 = n76199 & n76231;
  assign n76233 = pi2342 & n76232;
  assign n76234 = ~pi2342 & ~n76232;
  assign po2498 = n76233 | n76234;
  assign n76236 = ~n75172 & ~n75929;
  assign n76237 = ~n75090 & ~n76236;
  assign n76238 = ~n75154 & n75156;
  assign n76239 = n75090 & n76238;
  assign n76240 = n75108 & n75954;
  assign n76241 = ~n75919 & ~n76240;
  assign n76242 = ~n75119 & n76241;
  assign n76243 = ~n75090 & ~n76242;
  assign n76244 = ~n75096 & n75131;
  assign n76245 = ~n76243 & ~n76244;
  assign n76246 = ~n75154 & ~n76245;
  assign n76247 = ~n76239 & ~n76246;
  assign n76248 = ~n75117 & ~n75126;
  assign n76249 = ~n75096 & n75171;
  assign n76250 = ~n75898 & ~n76249;
  assign n76251 = n76248 & n76250;
  assign n76252 = n75090 & ~n76251;
  assign n76253 = n75102 & ~n75108;
  assign n76254 = n75090 & n76253;
  assign n76255 = n75096 & n76254;
  assign n76256 = ~n75096 & n75919;
  assign n76257 = ~n75117 & ~n76256;
  assign n76258 = ~n75926 & n76257;
  assign n76259 = ~n76255 & n76258;
  assign n76260 = ~n75090 & n75125;
  assign n76261 = n76259 & ~n76260;
  assign n76262 = n75154 & ~n76261;
  assign n76263 = ~n76252 & ~n76262;
  assign n76264 = n76247 & n76263;
  assign n76265 = ~n76237 & n76264;
  assign n76266 = pi2378 & n76265;
  assign n76267 = ~pi2378 & ~n76265;
  assign po2499 = n76266 | n76267;
  assign n76269 = n75796 & n75841;
  assign n76270 = ~n75854 & ~n76269;
  assign n76271 = n75814 & n76270;
  assign n76272 = ~n75796 & n76191;
  assign n76273 = ~n75806 & ~n75825;
  assign n76274 = n75802 & ~n76273;
  assign n76275 = n75784 & n75803;
  assign n76276 = ~n75796 & n75806;
  assign n76277 = ~n76275 & ~n76276;
  assign n76278 = ~n75814 & n76277;
  assign n76279 = ~n76274 & n76278;
  assign n76280 = ~n76272 & n76279;
  assign n76281 = ~n76271 & ~n76280;
  assign n76282 = ~n75796 & n76274;
  assign n76283 = ~n75843 & ~n76282;
  assign n76284 = ~n76281 & n76283;
  assign n76285 = n75839 & ~n76284;
  assign n76286 = n75814 & ~n76273;
  assign n76287 = n75796 & n76286;
  assign n76288 = ~n75852 & ~n76204;
  assign n76289 = ~n75796 & ~n76288;
  assign n76290 = n75814 & n76289;
  assign n76291 = ~n75802 & n76286;
  assign n76292 = ~n76290 & ~n76291;
  assign n76293 = ~n76287 & n76292;
  assign n76294 = ~n75839 & ~n76293;
  assign n76295 = ~n76285 & ~n76294;
  assign n76296 = ~n75814 & ~n76270;
  assign n76297 = ~n75846 & ~n76296;
  assign n76298 = ~n75839 & ~n76297;
  assign n76299 = n75814 & n75846;
  assign n76300 = ~n75814 & ~n76283;
  assign n76301 = ~n76299 & ~n76300;
  assign n76302 = ~n76298 & n76301;
  assign n76303 = n76295 & n76302;
  assign n76304 = pi2347 & ~n76303;
  assign n76305 = ~pi2347 & n76302;
  assign n76306 = ~n76294 & n76305;
  assign n76307 = ~n76285 & n76306;
  assign po2500 = n76304 | n76307;
  assign n76309 = n75814 & n75829;
  assign n76310 = n75803 & ~n76273;
  assign n76311 = ~n75853 & ~n76310;
  assign n76312 = ~n75843 & n76311;
  assign n76313 = ~n75814 & ~n76312;
  assign n76314 = ~n75796 & n76213;
  assign n76315 = ~n76313 & ~n76314;
  assign n76316 = ~n75802 & n75852;
  assign n76317 = n75796 & n75856;
  assign n76318 = ~n76316 & ~n76317;
  assign n76319 = ~n76276 & n76318;
  assign n76320 = n75814 & ~n76319;
  assign n76321 = n76315 & ~n76320;
  assign n76322 = n75839 & ~n76321;
  assign n76323 = ~n76309 & ~n76322;
  assign n76324 = n75796 & n75806;
  assign n76325 = ~n75842 & ~n76324;
  assign n76326 = n75814 & ~n76325;
  assign n76327 = ~n75824 & ~n76326;
  assign n76328 = ~n75829 & ~n76224;
  assign n76329 = ~n75796 & n75859;
  assign n76330 = ~n75856 & ~n76329;
  assign n76331 = ~n76316 & n76330;
  assign n76332 = ~n75814 & ~n76331;
  assign n76333 = n75796 & n76213;
  assign n76334 = ~n76332 & ~n76333;
  assign n76335 = n76328 & n76334;
  assign n76336 = n76327 & n76335;
  assign n76337 = ~n75839 & ~n76336;
  assign n76338 = ~n76205 & ~n76272;
  assign n76339 = ~n75814 & ~n76338;
  assign n76340 = ~n76337 & ~n76339;
  assign n76341 = n76323 & n76340;
  assign n76342 = pi2354 & n76341;
  assign n76343 = ~pi2354 & ~n76341;
  assign po2501 = n76342 | n76343;
  assign n76345 = pi4857 & ~pi9040;
  assign n76346 = pi4752 & pi9040;
  assign n76347 = ~n76345 & ~n76346;
  assign n76348 = ~pi2392 & n76347;
  assign n76349 = pi2392 & ~n76347;
  assign n76350 = ~n76348 & ~n76349;
  assign n76351 = pi4828 & pi9040;
  assign n76352 = pi4863 & ~pi9040;
  assign n76353 = ~n76351 & ~n76352;
  assign n76354 = pi2388 & n76353;
  assign n76355 = ~pi2388 & ~n76353;
  assign n76356 = ~n76354 & ~n76355;
  assign n76357 = pi4941 & pi9040;
  assign n76358 = pi4968 & ~pi9040;
  assign n76359 = ~n76357 & ~n76358;
  assign n76360 = pi2346 & n76359;
  assign n76361 = ~pi2346 & ~n76359;
  assign n76362 = ~n76360 & ~n76361;
  assign n76363 = pi4800 & pi9040;
  assign n76364 = pi5087 & ~pi9040;
  assign n76365 = ~n76363 & ~n76364;
  assign n76366 = ~pi2390 & n76365;
  assign n76367 = pi2390 & ~n76365;
  assign n76368 = ~n76366 & ~n76367;
  assign n76369 = pi4856 & ~pi9040;
  assign n76370 = pi5111 & pi9040;
  assign n76371 = ~n76369 & ~n76370;
  assign n76372 = ~pi2381 & n76371;
  assign n76373 = pi2381 & ~n76371;
  assign n76374 = ~n76372 & ~n76373;
  assign n76375 = n76368 & n76374;
  assign n76376 = n76362 & n76375;
  assign n76377 = n76356 & n76376;
  assign n76378 = ~n76368 & n76374;
  assign n76379 = ~n76362 & n76378;
  assign n76380 = n76356 & n76379;
  assign n76381 = ~n76377 & ~n76380;
  assign n76382 = ~n76368 & ~n76374;
  assign n76383 = ~n76362 & n76382;
  assign n76384 = ~n76356 & n76383;
  assign n76385 = ~n76356 & ~n76362;
  assign n76386 = n76374 & n76385;
  assign n76387 = n76368 & n76386;
  assign n76388 = ~n76384 & ~n76387;
  assign n76389 = n76381 & n76388;
  assign n76390 = ~n76350 & ~n76389;
  assign n76391 = n76368 & ~n76374;
  assign n76392 = ~n76362 & n76391;
  assign n76393 = n76356 & n76392;
  assign n76394 = ~n76379 & ~n76393;
  assign n76395 = ~n76350 & ~n76394;
  assign n76396 = n76350 & ~n76374;
  assign n76397 = ~n76356 & n76396;
  assign n76398 = n76362 & ~n76368;
  assign n76399 = n76356 & n76375;
  assign n76400 = ~n76398 & ~n76399;
  assign n76401 = n76350 & ~n76400;
  assign n76402 = ~n76397 & ~n76401;
  assign n76403 = n76362 & n76391;
  assign n76404 = ~n76356 & n76403;
  assign n76405 = n76402 & ~n76404;
  assign n76406 = ~n76374 & n76398;
  assign n76407 = n76356 & n76406;
  assign n76408 = n76405 & ~n76407;
  assign n76409 = ~n76395 & n76408;
  assign n76410 = pi4857 & pi9040;
  assign n76411 = pi4828 & ~pi9040;
  assign n76412 = ~n76410 & ~n76411;
  assign n76413 = ~pi2384 & ~n76412;
  assign n76414 = pi2384 & n76412;
  assign n76415 = ~n76413 & ~n76414;
  assign n76416 = ~n76409 & ~n76415;
  assign n76417 = n76350 & n76356;
  assign n76418 = ~n76362 & ~n76374;
  assign n76419 = n76415 & n76418;
  assign n76420 = n76417 & n76419;
  assign n76421 = n76350 & ~n76386;
  assign n76422 = n76356 & n76362;
  assign n76423 = n76368 & n76422;
  assign n76424 = ~n76382 & ~n76418;
  assign n76425 = ~n76356 & ~n76424;
  assign n76426 = ~n76350 & ~n76376;
  assign n76427 = ~n76425 & n76426;
  assign n76428 = ~n76423 & n76427;
  assign n76429 = ~n76421 & ~n76428;
  assign n76430 = n76362 & n76378;
  assign n76431 = n76356 & n76430;
  assign n76432 = ~n76429 & ~n76431;
  assign n76433 = n76415 & ~n76432;
  assign n76434 = ~n76420 & ~n76433;
  assign n76435 = ~n76416 & n76434;
  assign n76436 = ~n76390 & n76435;
  assign n76437 = n76350 & ~n76356;
  assign n76438 = n76391 & n76437;
  assign n76439 = n76362 & n76438;
  assign n76440 = n76436 & ~n76439;
  assign n76441 = pi2408 & ~n76440;
  assign n76442 = ~pi2408 & ~n76439;
  assign n76443 = n76435 & n76442;
  assign n76444 = ~n76390 & n76443;
  assign po2505 = n76441 | n76444;
  assign n76446 = pi4759 & pi9040;
  assign n76447 = pi4826 & ~pi9040;
  assign n76448 = ~n76446 & ~n76447;
  assign n76449 = ~pi2381 & ~n76448;
  assign n76450 = pi2381 & n76448;
  assign n76451 = ~n76449 & ~n76450;
  assign n76452 = pi4800 & ~pi9040;
  assign n76453 = pi4856 & pi9040;
  assign n76454 = ~n76452 & ~n76453;
  assign n76455 = ~pi2366 & n76454;
  assign n76456 = pi2366 & ~n76454;
  assign n76457 = ~n76455 & ~n76456;
  assign n76458 = pi5052 & ~pi9040;
  assign n76459 = pi4751 & pi9040;
  assign n76460 = ~n76458 & ~n76459;
  assign n76461 = ~pi2391 & ~n76460;
  assign n76462 = pi2391 & n76460;
  assign n76463 = ~n76461 & ~n76462;
  assign n76464 = pi4819 & ~pi9040;
  assign n76465 = pi5210 & pi9040;
  assign n76466 = ~n76464 & ~n76465;
  assign n76467 = ~pi2383 & n76466;
  assign n76468 = pi2383 & ~n76466;
  assign n76469 = ~n76467 & ~n76468;
  assign n76470 = pi5111 & ~pi9040;
  assign n76471 = pi5087 & pi9040;
  assign n76472 = ~n76470 & ~n76471;
  assign n76473 = ~pi2346 & n76472;
  assign n76474 = pi2346 & ~n76472;
  assign n76475 = ~n76473 & ~n76474;
  assign n76476 = n76469 & ~n76475;
  assign n76477 = ~n76463 & n76476;
  assign n76478 = n76457 & n76477;
  assign n76479 = pi4941 & ~pi9040;
  assign n76480 = pi5052 & pi9040;
  assign n76481 = ~n76479 & ~n76480;
  assign n76482 = ~pi2377 & n76481;
  assign n76483 = pi2377 & ~n76481;
  assign n76484 = ~n76482 & ~n76483;
  assign n76485 = ~n76469 & n76475;
  assign n76486 = ~n76484 & n76485;
  assign n76487 = n76475 & n76484;
  assign n76488 = ~n76457 & n76487;
  assign n76489 = n76469 & n76488;
  assign n76490 = ~n76486 & ~n76489;
  assign n76491 = ~n76469 & ~n76475;
  assign n76492 = ~n76457 & n76491;
  assign n76493 = n76490 & ~n76492;
  assign n76494 = ~n76463 & ~n76493;
  assign n76495 = ~n76469 & n76484;
  assign n76496 = n76457 & n76463;
  assign n76497 = n76495 & n76496;
  assign n76498 = n76457 & n76484;
  assign n76499 = n76475 & n76498;
  assign n76500 = ~n76469 & n76499;
  assign n76501 = ~n76497 & ~n76500;
  assign n76502 = ~n76494 & n76501;
  assign n76503 = ~n76478 & n76502;
  assign n76504 = n76476 & ~n76484;
  assign n76505 = n76457 & n76504;
  assign n76506 = ~n76484 & n76491;
  assign n76507 = ~n76457 & n76506;
  assign n76508 = ~n76505 & ~n76507;
  assign n76509 = n76503 & n76508;
  assign n76510 = ~n76451 & ~n76509;
  assign n76511 = ~n76475 & n76498;
  assign n76512 = ~n76469 & n76511;
  assign n76513 = ~n76504 & ~n76512;
  assign n76514 = ~n76463 & ~n76513;
  assign n76515 = ~n76457 & n76484;
  assign n76516 = n76476 & n76515;
  assign n76517 = n76469 & n76499;
  assign n76518 = ~n76516 & ~n76517;
  assign n76519 = ~n76469 & n76515;
  assign n76520 = n76457 & n76506;
  assign n76521 = ~n76519 & ~n76520;
  assign n76522 = n76463 & ~n76521;
  assign n76523 = n76518 & ~n76522;
  assign n76524 = ~n76514 & n76523;
  assign n76525 = n76451 & ~n76524;
  assign n76526 = n76469 & ~n76484;
  assign n76527 = n76457 & n76526;
  assign n76528 = ~n76469 & ~n76484;
  assign n76529 = ~n76457 & n76528;
  assign n76530 = ~n76527 & ~n76529;
  assign n76531 = ~n76463 & ~n76530;
  assign n76532 = ~n76457 & ~n76484;
  assign n76533 = n76475 & n76532;
  assign n76534 = n76469 & n76533;
  assign n76535 = ~n76516 & ~n76534;
  assign n76536 = n76484 & n76485;
  assign n76537 = n76535 & ~n76536;
  assign n76538 = n76463 & ~n76537;
  assign n76539 = ~n76531 & ~n76538;
  assign n76540 = n76463 & n76487;
  assign n76541 = n76457 & n76540;
  assign n76542 = n76539 & ~n76541;
  assign n76543 = ~n76525 & n76542;
  assign n76544 = ~n76510 & n76543;
  assign n76545 = pi2425 & n76544;
  assign n76546 = ~pi2425 & ~n76544;
  assign po2521 = n76545 | n76546;
  assign n76548 = ~n76517 & ~n76528;
  assign n76549 = n76463 & ~n76548;
  assign n76550 = ~n76457 & n76536;
  assign n76551 = ~n76549 & ~n76550;
  assign n76552 = ~n76512 & n76551;
  assign n76553 = ~n76463 & n76516;
  assign n76554 = ~n76505 & ~n76553;
  assign n76555 = ~n76534 & n76554;
  assign n76556 = n76552 & n76555;
  assign n76557 = n76451 & ~n76556;
  assign n76558 = n76484 & n76491;
  assign n76559 = ~n76457 & n76558;
  assign n76560 = ~n76489 & ~n76559;
  assign n76561 = n76476 & n76484;
  assign n76562 = n76463 & n76561;
  assign n76563 = ~n76457 & n76504;
  assign n76564 = ~n76562 & ~n76563;
  assign n76565 = n76469 & n76475;
  assign n76566 = ~n76484 & n76565;
  assign n76567 = n76457 & n76566;
  assign n76568 = ~n76500 & ~n76567;
  assign n76569 = ~n76475 & ~n76484;
  assign n76570 = ~n76457 & ~n76469;
  assign n76571 = ~n76569 & ~n76570;
  assign n76572 = ~n76487 & n76571;
  assign n76573 = ~n76463 & ~n76572;
  assign n76574 = n76568 & ~n76573;
  assign n76575 = n76564 & n76574;
  assign n76576 = n76560 & n76575;
  assign n76577 = ~n76451 & ~n76576;
  assign n76578 = ~n76557 & ~n76577;
  assign n76579 = pi2420 & ~n76578;
  assign n76580 = ~pi2420 & ~n76557;
  assign n76581 = ~n76577 & n76580;
  assign po2525 = n76579 | n76581;
  assign n76583 = ~n76356 & n76406;
  assign n76584 = n76356 & n76418;
  assign n76585 = ~n76403 & ~n76584;
  assign n76586 = ~n76350 & ~n76585;
  assign n76587 = ~n76583 & ~n76586;
  assign n76588 = ~n76374 & n76437;
  assign n76589 = ~n76368 & n76588;
  assign n76590 = n76378 & n76417;
  assign n76591 = ~n76589 & ~n76590;
  assign n76592 = n76350 & n76376;
  assign n76593 = n76591 & ~n76592;
  assign n76594 = ~n76387 & ~n76393;
  assign n76595 = n76374 & n76422;
  assign n76596 = n76594 & ~n76595;
  assign n76597 = n76593 & n76596;
  assign n76598 = n76587 & n76597;
  assign n76599 = ~n76415 & ~n76598;
  assign n76600 = ~n76362 & n76375;
  assign n76601 = ~n76403 & ~n76600;
  assign n76602 = n76356 & ~n76601;
  assign n76603 = ~n76368 & n76385;
  assign n76604 = ~n76430 & ~n76603;
  assign n76605 = n76362 & ~n76374;
  assign n76606 = n76356 & n76605;
  assign n76607 = n76604 & ~n76606;
  assign n76608 = ~n76350 & ~n76607;
  assign n76609 = ~n76356 & n76391;
  assign n76610 = n76356 & ~n76362;
  assign n76611 = ~n76374 & n76610;
  assign n76612 = ~n76368 & n76611;
  assign n76613 = ~n76609 & ~n76612;
  assign n76614 = n76350 & ~n76613;
  assign n76615 = ~n76356 & n76379;
  assign n76616 = ~n76614 & ~n76615;
  assign n76617 = ~n76608 & n76616;
  assign n76618 = ~n76602 & n76617;
  assign n76619 = n76415 & ~n76618;
  assign n76620 = ~n76350 & n76386;
  assign n76621 = ~n76619 & ~n76620;
  assign n76622 = n76398 & n76437;
  assign n76623 = ~n76374 & n76622;
  assign n76624 = n76621 & ~n76623;
  assign n76625 = ~n76599 & n76624;
  assign n76626 = ~pi2431 & ~n76625;
  assign n76627 = pi2431 & n76621;
  assign n76628 = ~n76599 & n76627;
  assign n76629 = ~n76623 & n76628;
  assign po2526 = n76626 | n76629;
  assign n76631 = pi4750 & ~pi9040;
  assign n76632 = pi4827 & pi9040;
  assign n76633 = ~n76631 & ~n76632;
  assign n76634 = ~pi2384 & ~n76633;
  assign n76635 = pi2384 & n76633;
  assign n76636 = ~n76634 & ~n76635;
  assign n76637 = pi4953 & ~pi9040;
  assign n76638 = pi4829 & pi9040;
  assign n76639 = ~n76637 & ~n76638;
  assign n76640 = ~pi2390 & ~n76639;
  assign n76641 = pi2390 & n76639;
  assign n76642 = ~n76640 & ~n76641;
  assign n76643 = pi4829 & ~pi9040;
  assign n76644 = pi5211 & pi9040;
  assign n76645 = ~n76643 & ~n76644;
  assign n76646 = pi2387 & n76645;
  assign n76647 = ~pi2387 & ~n76645;
  assign n76648 = ~n76646 & ~n76647;
  assign n76649 = n76642 & ~n76648;
  assign n76650 = n76636 & n76649;
  assign n76651 = pi5095 & ~pi9040;
  assign n76652 = pi4825 & pi9040;
  assign n76653 = ~n76651 & ~n76652;
  assign n76654 = ~pi2389 & n76653;
  assign n76655 = pi2389 & ~n76653;
  assign n76656 = ~n76654 & ~n76655;
  assign n76657 = ~n76636 & ~n76656;
  assign n76658 = ~n76642 & n76657;
  assign n76659 = ~n76650 & ~n76658;
  assign n76660 = pi4758 & pi9040;
  assign n76661 = pi5295 & ~pi9040;
  assign n76662 = ~n76660 & ~n76661;
  assign n76663 = ~pi2364 & n76662;
  assign n76664 = pi2364 & ~n76662;
  assign n76665 = ~n76663 & ~n76664;
  assign n76666 = ~n76636 & ~n76665;
  assign n76667 = ~n76642 & n76666;
  assign n76668 = n76659 & ~n76667;
  assign n76669 = ~n76642 & n76665;
  assign n76670 = n76636 & n76669;
  assign n76671 = n76656 & n76670;
  assign n76672 = n76668 & ~n76671;
  assign n76673 = ~n76636 & n76665;
  assign n76674 = ~n76656 & n76673;
  assign n76675 = ~n76642 & ~n76665;
  assign n76676 = ~n76674 & ~n76675;
  assign n76677 = n76648 & ~n76676;
  assign n76678 = n76648 & n76666;
  assign n76679 = n76656 & n76678;
  assign n76680 = ~n76677 & ~n76679;
  assign n76681 = n76672 & n76680;
  assign n76682 = pi4978 & ~pi9040;
  assign n76683 = pi4865 & pi9040;
  assign n76684 = ~n76682 & ~n76683;
  assign n76685 = ~pi2360 & ~n76684;
  assign n76686 = pi2360 & n76684;
  assign n76687 = ~n76685 & ~n76686;
  assign n76688 = ~n76681 & n76687;
  assign n76689 = ~n76642 & ~n76656;
  assign n76690 = n76648 & n76689;
  assign n76691 = n76673 & n76690;
  assign n76692 = n76648 & ~n76656;
  assign n76693 = n76666 & n76692;
  assign n76694 = n76642 & n76693;
  assign n76695 = n76636 & ~n76665;
  assign n76696 = n76648 & n76656;
  assign n76697 = n76695 & n76696;
  assign n76698 = n76642 & n76656;
  assign n76699 = n76665 & n76698;
  assign n76700 = ~n76636 & n76699;
  assign n76701 = n76636 & n76665;
  assign n76702 = n76642 & n76701;
  assign n76703 = n76648 & n76702;
  assign n76704 = ~n76656 & n76703;
  assign n76705 = ~n76700 & ~n76704;
  assign n76706 = ~n76697 & n76705;
  assign n76707 = ~n76694 & n76706;
  assign n76708 = ~n76642 & n76656;
  assign n76709 = ~n76665 & n76708;
  assign n76710 = n76636 & n76709;
  assign n76711 = n76707 & ~n76710;
  assign n76712 = ~n76687 & ~n76711;
  assign n76713 = n76636 & n76642;
  assign n76714 = ~n76665 & n76713;
  assign n76715 = ~n76656 & n76714;
  assign n76716 = ~n76699 & ~n76715;
  assign n76717 = ~n76656 & n76667;
  assign n76718 = n76716 & ~n76717;
  assign n76719 = ~n76648 & ~n76718;
  assign n76720 = ~n76648 & ~n76656;
  assign n76721 = n76670 & n76720;
  assign n76722 = ~n76636 & n76698;
  assign n76723 = n76656 & n76673;
  assign n76724 = ~n76722 & ~n76723;
  assign n76725 = ~n76648 & ~n76724;
  assign n76726 = ~n76721 & ~n76725;
  assign n76727 = ~n76687 & ~n76726;
  assign n76728 = ~n76719 & ~n76727;
  assign n76729 = ~n76712 & n76728;
  assign n76730 = ~n76691 & n76729;
  assign n76731 = ~n76688 & n76730;
  assign n76732 = n76636 & ~n76642;
  assign n76733 = n76696 & n76732;
  assign n76734 = n76731 & ~n76733;
  assign n76735 = ~pi2402 & ~n76734;
  assign n76736 = pi2402 & ~n76733;
  assign n76737 = n76730 & n76736;
  assign n76738 = ~n76688 & n76737;
  assign po2528 = n76735 | n76738;
  assign n76740 = pi4848 & ~pi9040;
  assign n76741 = pi4870 & pi9040;
  assign n76742 = ~n76740 & ~n76741;
  assign n76743 = ~pi2395 & ~n76742;
  assign n76744 = pi2395 & n76742;
  assign n76745 = ~n76743 & ~n76744;
  assign n76746 = pi5114 & ~pi9040;
  assign n76747 = pi4869 & pi9040;
  assign n76748 = ~n76746 & ~n76747;
  assign n76749 = ~pi2379 & n76748;
  assign n76750 = pi2379 & ~n76748;
  assign n76751 = ~n76749 & ~n76750;
  assign n76752 = pi5277 & ~pi9040;
  assign n76753 = pi4750 & pi9040;
  assign n76754 = ~n76752 & ~n76753;
  assign n76755 = ~pi2398 & n76754;
  assign n76756 = pi2398 & ~n76754;
  assign n76757 = ~n76755 & ~n76756;
  assign n76758 = pi4977 & ~pi9040;
  assign n76759 = pi4866 & pi9040;
  assign n76760 = ~n76758 & ~n76759;
  assign n76761 = ~pi2367 & n76760;
  assign n76762 = pi2367 & ~n76760;
  assign n76763 = ~n76761 & ~n76762;
  assign n76764 = pi4951 & pi9040;
  assign n76765 = pi4862 & ~pi9040;
  assign n76766 = ~n76764 & ~n76765;
  assign n76767 = ~pi2386 & n76766;
  assign n76768 = pi2386 & ~n76766;
  assign n76769 = ~n76767 & ~n76768;
  assign n76770 = ~n76763 & n76769;
  assign n76771 = ~n76757 & n76770;
  assign n76772 = ~n76751 & n76771;
  assign n76773 = n76763 & n76769;
  assign n76774 = ~n76757 & n76773;
  assign n76775 = n76751 & n76774;
  assign n76776 = ~n76772 & ~n76775;
  assign n76777 = n76763 & ~n76769;
  assign n76778 = ~n76757 & n76777;
  assign n76779 = ~n76751 & n76778;
  assign n76780 = pi5114 & pi9040;
  assign n76781 = pi4870 & ~pi9040;
  assign n76782 = ~n76780 & ~n76781;
  assign n76783 = ~pi2396 & ~n76782;
  assign n76784 = pi2396 & n76782;
  assign n76785 = ~n76783 & ~n76784;
  assign n76786 = ~n76763 & ~n76769;
  assign n76787 = ~n76751 & n76786;
  assign n76788 = n76757 & n76777;
  assign n76789 = n76751 & n76788;
  assign n76790 = ~n76787 & ~n76789;
  assign n76791 = ~n76785 & ~n76790;
  assign n76792 = ~n76779 & ~n76791;
  assign n76793 = n76757 & n76773;
  assign n76794 = n76785 & n76793;
  assign n76795 = n76777 & n76785;
  assign n76796 = ~n76751 & n76795;
  assign n76797 = ~n76794 & ~n76796;
  assign n76798 = n76792 & n76797;
  assign n76799 = n76776 & n76798;
  assign n76800 = n76745 & ~n76799;
  assign n76801 = ~n76745 & ~n76785;
  assign n76802 = ~n76751 & n76757;
  assign n76803 = n76763 & n76802;
  assign n76804 = n76757 & n76769;
  assign n76805 = ~n76803 & ~n76804;
  assign n76806 = n76801 & ~n76805;
  assign n76807 = n76751 & ~n76757;
  assign n76808 = ~n76769 & n76807;
  assign n76809 = n76763 & n76808;
  assign n76810 = n76751 & ~n76763;
  assign n76811 = n76757 & n76810;
  assign n76812 = ~n76809 & ~n76811;
  assign n76813 = ~n76751 & n76785;
  assign n76814 = ~n76757 & n76813;
  assign n76815 = ~n76777 & n76814;
  assign n76816 = n76771 & n76785;
  assign n76817 = ~n76815 & ~n76816;
  assign n76818 = n76812 & n76817;
  assign n76819 = ~n76745 & ~n76818;
  assign n76820 = n76757 & n76770;
  assign n76821 = ~n76785 & n76820;
  assign n76822 = n76751 & n76821;
  assign n76823 = ~n76757 & n76786;
  assign n76824 = n76751 & n76823;
  assign n76825 = ~n76775 & ~n76824;
  assign n76826 = ~n76785 & ~n76825;
  assign n76827 = ~n76822 & ~n76826;
  assign n76828 = n76785 & n76809;
  assign n76829 = n76827 & ~n76828;
  assign n76830 = ~n76819 & n76829;
  assign n76831 = ~n76806 & n76830;
  assign n76832 = ~n76800 & n76831;
  assign n76833 = n76757 & n76786;
  assign n76834 = n76751 & n76785;
  assign n76835 = n76833 & n76834;
  assign n76836 = n76832 & ~n76835;
  assign n76837 = ~pi2401 & ~n76836;
  assign n76838 = pi2401 & ~n76835;
  assign n76839 = n76831 & n76838;
  assign n76840 = ~n76800 & n76839;
  assign po2531 = n76837 | n76840;
  assign n76842 = ~n76431 & ~n76615;
  assign n76843 = ~n76350 & ~n76842;
  assign n76844 = ~n76415 & n76418;
  assign n76845 = n76350 & n76844;
  assign n76846 = ~n76356 & n76362;
  assign n76847 = n76368 & n76846;
  assign n76848 = ~n76605 & ~n76847;
  assign n76849 = ~n76379 & n76848;
  assign n76850 = ~n76350 & ~n76849;
  assign n76851 = ~n76356 & n76392;
  assign n76852 = ~n76850 & ~n76851;
  assign n76853 = ~n76415 & ~n76852;
  assign n76854 = ~n76845 & ~n76853;
  assign n76855 = ~n76377 & ~n76387;
  assign n76856 = ~n76356 & n76430;
  assign n76857 = ~n76584 & ~n76856;
  assign n76858 = n76855 & n76857;
  assign n76859 = n76350 & ~n76858;
  assign n76860 = ~n76362 & ~n76368;
  assign n76861 = n76350 & n76860;
  assign n76862 = n76356 & n76861;
  assign n76863 = ~n76356 & n76605;
  assign n76864 = ~n76377 & ~n76863;
  assign n76865 = ~n76612 & n76864;
  assign n76866 = ~n76862 & n76865;
  assign n76867 = ~n76350 & n76600;
  assign n76868 = n76866 & ~n76867;
  assign n76869 = n76415 & ~n76868;
  assign n76870 = ~n76859 & ~n76869;
  assign n76871 = n76854 & n76870;
  assign n76872 = ~n76843 & n76871;
  assign n76873 = pi2460 & n76872;
  assign n76874 = ~pi2460 & ~n76872;
  assign po2534 = n76873 | n76874;
  assign n76876 = pi4869 & ~pi9040;
  assign n76877 = pi4848 & pi9040;
  assign n76878 = ~n76876 & ~n76877;
  assign n76879 = pi2371 & n76878;
  assign n76880 = ~pi2371 & ~n76878;
  assign n76881 = ~n76879 & ~n76880;
  assign n76882 = pi4938 & pi9040;
  assign n76883 = pi5211 & ~pi9040;
  assign n76884 = ~n76882 & ~n76883;
  assign n76885 = pi2360 & n76884;
  assign n76886 = ~pi2360 & ~n76884;
  assign n76887 = ~n76885 & ~n76886;
  assign n76888 = pi4938 & ~pi9040;
  assign n76889 = pi4953 & pi9040;
  assign n76890 = ~n76888 & ~n76889;
  assign n76891 = ~pi2393 & n76890;
  assign n76892 = pi2393 & ~n76890;
  assign n76893 = ~n76891 & ~n76892;
  assign n76894 = n76887 & n76893;
  assign n76895 = pi4942 & ~pi9040;
  assign n76896 = pi5277 & pi9040;
  assign n76897 = ~n76895 & ~n76896;
  assign n76898 = pi2364 & n76897;
  assign n76899 = ~pi2364 & ~n76897;
  assign n76900 = ~n76898 & ~n76899;
  assign n76901 = pi4956 & pi9040;
  assign n76902 = pi5092 & ~pi9040;
  assign n76903 = ~n76901 & ~n76902;
  assign n76904 = pi2394 & n76903;
  assign n76905 = ~pi2394 & ~n76903;
  assign n76906 = ~n76904 & ~n76905;
  assign n76907 = n76900 & n76906;
  assign n76908 = n76894 & n76907;
  assign n76909 = ~n76900 & n76906;
  assign n76910 = ~n76887 & n76909;
  assign n76911 = ~n76908 & ~n76910;
  assign n76912 = ~n76881 & ~n76911;
  assign n76913 = pi4827 & ~pi9040;
  assign n76914 = pi4942 & pi9040;
  assign n76915 = ~n76913 & ~n76914;
  assign n76916 = ~pi2370 & ~n76915;
  assign n76917 = pi2370 & n76915;
  assign n76918 = ~n76916 & ~n76917;
  assign n76919 = n76881 & ~n76906;
  assign n76920 = n76887 & n76919;
  assign n76921 = n76894 & ~n76900;
  assign n76922 = n76887 & ~n76893;
  assign n76923 = n76900 & n76922;
  assign n76924 = ~n76921 & ~n76923;
  assign n76925 = ~n76887 & n76893;
  assign n76926 = n76900 & n76925;
  assign n76927 = n76906 & n76926;
  assign n76928 = n76924 & ~n76927;
  assign n76929 = n76881 & ~n76928;
  assign n76930 = ~n76920 & ~n76929;
  assign n76931 = ~n76887 & ~n76893;
  assign n76932 = ~n76900 & n76931;
  assign n76933 = n76906 & n76932;
  assign n76934 = n76930 & ~n76933;
  assign n76935 = ~n76906 & n76925;
  assign n76936 = n76900 & n76931;
  assign n76937 = ~n76935 & ~n76936;
  assign n76938 = ~n76881 & ~n76937;
  assign n76939 = ~n76900 & n76922;
  assign n76940 = ~n76906 & n76939;
  assign n76941 = ~n76938 & ~n76940;
  assign n76942 = n76934 & n76941;
  assign n76943 = n76918 & ~n76942;
  assign n76944 = ~n76912 & ~n76943;
  assign n76945 = ~n76900 & n76925;
  assign n76946 = ~n76939 & ~n76945;
  assign n76947 = n76906 & ~n76946;
  assign n76948 = ~n76908 & ~n76947;
  assign n76949 = ~n76918 & ~n76948;
  assign n76950 = n76881 & ~n76918;
  assign n76951 = ~n76937 & n76950;
  assign n76952 = ~n76949 & ~n76951;
  assign n76953 = ~n76881 & ~n76918;
  assign n76954 = n76894 & ~n76906;
  assign n76955 = ~n76932 & ~n76954;
  assign n76956 = n76887 & n76900;
  assign n76957 = n76955 & ~n76956;
  assign n76958 = n76953 & ~n76957;
  assign n76959 = n76952 & ~n76958;
  assign n76960 = n76944 & n76959;
  assign n76961 = ~pi2407 & ~n76960;
  assign n76962 = pi2407 & n76952;
  assign n76963 = n76944 & n76962;
  assign n76964 = ~n76958 & n76963;
  assign po2535 = n76961 | n76964;
  assign n76966 = ~n76377 & ~n76384;
  assign n76967 = n76350 & ~n76966;
  assign n76968 = ~n76439 & ~n76967;
  assign n76969 = n76350 & n76382;
  assign n76970 = n76356 & n76969;
  assign n76971 = ~n76592 & ~n76970;
  assign n76972 = ~n76362 & n76368;
  assign n76973 = n76356 & n76391;
  assign n76974 = ~n76972 & ~n76973;
  assign n76975 = ~n76368 & n76846;
  assign n76976 = n76974 & ~n76975;
  assign n76977 = ~n76350 & ~n76976;
  assign n76978 = ~n76380 & ~n76977;
  assign n76979 = n76971 & n76978;
  assign n76980 = ~n76415 & ~n76979;
  assign n76981 = ~n76350 & n76972;
  assign n76982 = n76356 & n76981;
  assign n76983 = ~n76980 & ~n76982;
  assign n76984 = ~n76386 & ~n76403;
  assign n76985 = ~n76430 & n76984;
  assign n76986 = n76350 & ~n76985;
  assign n76987 = ~n76356 & n76376;
  assign n76988 = ~n76406 & ~n76987;
  assign n76989 = ~n76350 & ~n76988;
  assign n76990 = ~n76603 & ~n76989;
  assign n76991 = ~n76986 & n76990;
  assign n76992 = ~n76393 & ~n76431;
  assign n76993 = n76991 & n76992;
  assign n76994 = n76415 & ~n76993;
  assign n76995 = n76983 & ~n76994;
  assign n76996 = n76968 & n76995;
  assign n76997 = pi2451 & n76996;
  assign n76998 = ~pi2451 & ~n76996;
  assign po2537 = n76997 | n76998;
  assign n77000 = ~n76476 & ~n76485;
  assign n77001 = n76463 & ~n77000;
  assign n77002 = n76457 & n77001;
  assign n77003 = ~n76506 & ~n76565;
  assign n77004 = ~n76457 & ~n77003;
  assign n77005 = n76463 & n77004;
  assign n77006 = n76484 & n77001;
  assign n77007 = ~n77005 & ~n77006;
  assign n77008 = ~n77002 & n77007;
  assign n77009 = ~n76451 & ~n77008;
  assign n77010 = n76457 & n76491;
  assign n77011 = ~n76567 & ~n77010;
  assign n77012 = n76463 & n77011;
  assign n77013 = ~n76457 & n76526;
  assign n77014 = ~n76484 & ~n77000;
  assign n77015 = n76469 & n76498;
  assign n77016 = ~n76457 & n76485;
  assign n77017 = ~n77015 & ~n77016;
  assign n77018 = ~n76463 & n77017;
  assign n77019 = ~n77014 & n77018;
  assign n77020 = ~n77013 & n77019;
  assign n77021 = ~n77012 & ~n77020;
  assign n77022 = ~n76457 & n77014;
  assign n77023 = ~n76559 & ~n77022;
  assign n77024 = ~n77021 & n77023;
  assign n77025 = n76451 & ~n77024;
  assign n77026 = ~n77009 & ~n77025;
  assign n77027 = n76463 & n76489;
  assign n77028 = ~n76463 & ~n77023;
  assign n77029 = ~n77027 & ~n77028;
  assign n77030 = ~n76463 & ~n77011;
  assign n77031 = ~n76489 & ~n77030;
  assign n77032 = ~n76451 & ~n77031;
  assign n77033 = n77029 & ~n77032;
  assign n77034 = n77026 & n77033;
  assign n77035 = pi2436 & ~n77034;
  assign n77036 = ~pi2436 & n77033;
  assign n77037 = ~n77009 & n77036;
  assign n77038 = ~n77025 & n77037;
  assign po2538 = n77035 | n77038;
  assign n77040 = n76751 & n76757;
  assign n77041 = n76769 & n77040;
  assign n77042 = n76763 & n77041;
  assign n77043 = n76769 & n76802;
  assign n77044 = ~n76763 & n77043;
  assign n77045 = ~n77042 & ~n77044;
  assign n77046 = n76785 & ~n77045;
  assign n77047 = ~n76809 & ~n76816;
  assign n77048 = n76763 & n76807;
  assign n77049 = ~n76811 & ~n77048;
  assign n77050 = ~n76785 & ~n77049;
  assign n77051 = ~n76751 & ~n76785;
  assign n77052 = n76773 & n77051;
  assign n77053 = n76757 & n77052;
  assign n77054 = n76757 & n76785;
  assign n77055 = ~n76769 & n77054;
  assign n77056 = n76763 & n77055;
  assign n77057 = ~n76751 & n76823;
  assign n77058 = ~n77056 & ~n77057;
  assign n77059 = ~n77053 & n77058;
  assign n77060 = ~n77050 & n77059;
  assign n77061 = n77047 & n77060;
  assign n77062 = n76745 & ~n77061;
  assign n77063 = ~n76785 & n76809;
  assign n77064 = n76751 & n76816;
  assign n77065 = ~n77063 & ~n77064;
  assign n77066 = ~n77062 & n77065;
  assign n77067 = ~n77046 & n77066;
  assign n77068 = ~n76757 & n76763;
  assign n77069 = n76813 & n77068;
  assign n77070 = ~n76794 & ~n77069;
  assign n77071 = n76785 & n76823;
  assign n77072 = n76751 & n76833;
  assign n77073 = ~n77071 & ~n77072;
  assign n77074 = ~n76751 & n76770;
  assign n77075 = n76757 & ~n76769;
  assign n77076 = ~n77074 & ~n77075;
  assign n77077 = ~n76785 & ~n77076;
  assign n77078 = ~n76751 & n76774;
  assign n77079 = ~n77042 & ~n77078;
  assign n77080 = ~n77077 & n77079;
  assign n77081 = n77073 & n77080;
  assign n77082 = n77070 & n77081;
  assign n77083 = ~n76745 & ~n77082;
  assign n77084 = n77067 & ~n77083;
  assign n77085 = ~pi2400 & ~n77084;
  assign n77086 = pi2400 & n77067;
  assign n77087 = ~n77083 & n77086;
  assign po2540 = n77085 | n77087;
  assign n77089 = n76457 & n76485;
  assign n77090 = ~n76558 & ~n77089;
  assign n77091 = n76463 & ~n77090;
  assign n77092 = ~n76534 & ~n77091;
  assign n77093 = ~n76507 & ~n76516;
  assign n77094 = ~n76488 & ~n76569;
  assign n77095 = n76484 & n76565;
  assign n77096 = n77094 & ~n77095;
  assign n77097 = ~n76463 & ~n77096;
  assign n77098 = n76457 & n76486;
  assign n77099 = ~n77097 & ~n77098;
  assign n77100 = n77093 & n77099;
  assign n77101 = n77092 & n77100;
  assign n77102 = ~n76451 & ~n77101;
  assign n77103 = ~n76520 & ~n77013;
  assign n77104 = ~n76463 & ~n77103;
  assign n77105 = ~n77102 & ~n77104;
  assign n77106 = n76463 & n76516;
  assign n77107 = n76498 & ~n77000;
  assign n77108 = ~n76559 & ~n76566;
  assign n77109 = ~n77107 & n77108;
  assign n77110 = ~n76463 & ~n77109;
  assign n77111 = ~n76457 & n76486;
  assign n77112 = ~n77110 & ~n77111;
  assign n77113 = n76457 & n76569;
  assign n77114 = ~n77095 & ~n77113;
  assign n77115 = ~n77016 & n77114;
  assign n77116 = n76463 & ~n77115;
  assign n77117 = n77112 & ~n77116;
  assign n77118 = n76451 & ~n77117;
  assign n77119 = ~n77106 & ~n77118;
  assign n77120 = n77105 & n77119;
  assign n77121 = pi2443 & n77120;
  assign n77122 = ~pi2443 & ~n77120;
  assign po2542 = n77121 | n77122;
  assign n77124 = pi4758 & ~pi9040;
  assign n77125 = pi4948 & pi9040;
  assign n77126 = ~n77124 & ~n77125;
  assign n77127 = pi2385 & n77126;
  assign n77128 = ~pi2385 & ~n77126;
  assign n77129 = ~n77127 & ~n77128;
  assign n77130 = pi4761 & ~pi9040;
  assign n77131 = pi5095 & pi9040;
  assign n77132 = ~n77130 & ~n77131;
  assign n77133 = ~pi2352 & n77132;
  assign n77134 = pi2352 & ~n77132;
  assign n77135 = ~n77133 & ~n77134;
  assign n77136 = pi4866 & ~pi9040;
  assign n77137 = pi4862 & pi9040;
  assign n77138 = ~n77136 & ~n77137;
  assign n77139 = pi2370 & n77138;
  assign n77140 = ~pi2370 & ~n77138;
  assign n77141 = ~n77139 & ~n77140;
  assign n77142 = pi4948 & ~pi9040;
  assign n77143 = pi4954 & pi9040;
  assign n77144 = ~n77142 & ~n77143;
  assign n77145 = ~pi2393 & ~n77144;
  assign n77146 = pi2393 & n77144;
  assign n77147 = ~n77145 & ~n77146;
  assign n77148 = n77141 & ~n77147;
  assign n77149 = n77135 & n77148;
  assign n77150 = n77129 & n77149;
  assign n77151 = pi5295 & pi9040;
  assign n77152 = pi4954 & ~pi9040;
  assign n77153 = ~n77151 & ~n77152;
  assign n77154 = ~pi2367 & n77153;
  assign n77155 = pi2367 & ~n77153;
  assign n77156 = ~n77154 & ~n77155;
  assign n77157 = pi4865 & ~pi9040;
  assign n77158 = pi5092 & pi9040;
  assign n77159 = ~n77157 & ~n77158;
  assign n77160 = ~pi2398 & n77159;
  assign n77161 = pi2398 & ~n77159;
  assign n77162 = ~n77160 & ~n77161;
  assign n77163 = n77141 & ~n77162;
  assign n77164 = n77147 & n77163;
  assign n77165 = ~n77141 & ~n77162;
  assign n77166 = ~n77147 & n77165;
  assign n77167 = ~n77141 & n77162;
  assign n77168 = ~n77129 & n77167;
  assign n77169 = ~n77166 & ~n77168;
  assign n77170 = ~n77164 & n77169;
  assign n77171 = n77135 & ~n77170;
  assign n77172 = n77147 & n77165;
  assign n77173 = ~n77147 & n77163;
  assign n77174 = ~n77172 & ~n77173;
  assign n77175 = ~n77135 & ~n77174;
  assign n77176 = ~n77171 & ~n77175;
  assign n77177 = n77141 & n77162;
  assign n77178 = n77147 & n77177;
  assign n77179 = ~n77135 & n77178;
  assign n77180 = ~n77147 & n77168;
  assign n77181 = ~n77179 & ~n77180;
  assign n77182 = n77176 & n77181;
  assign n77183 = n77156 & ~n77182;
  assign n77184 = n77129 & n77172;
  assign n77185 = ~n77129 & n77177;
  assign n77186 = n77129 & n77167;
  assign n77187 = ~n77185 & ~n77186;
  assign n77188 = n77135 & ~n77187;
  assign n77189 = ~n77184 & ~n77188;
  assign n77190 = n77147 & n77167;
  assign n77191 = ~n77135 & n77190;
  assign n77192 = ~n77147 & n77177;
  assign n77193 = ~n77164 & ~n77192;
  assign n77194 = ~n77191 & n77193;
  assign n77195 = ~n77166 & n77194;
  assign n77196 = ~n77129 & ~n77195;
  assign n77197 = n77189 & ~n77196;
  assign n77198 = ~n77156 & ~n77197;
  assign n77199 = ~n77183 & ~n77198;
  assign n77200 = ~n77150 & n77199;
  assign n77201 = ~n77147 & n77186;
  assign n77202 = n77129 & n77147;
  assign n77203 = n77162 & n77202;
  assign n77204 = n77141 & n77203;
  assign n77205 = ~n77201 & ~n77204;
  assign n77206 = ~n77135 & ~n77205;
  assign n77207 = n77200 & ~n77206;
  assign n77208 = ~pi2449 & ~n77207;
  assign n77209 = n77199 & ~n77206;
  assign n77210 = pi2449 & n77209;
  assign n77211 = ~n77150 & n77210;
  assign po2543 = n77208 | n77211;
  assign n77213 = ~n77129 & n77147;
  assign n77214 = ~n77162 & n77213;
  assign n77215 = n77193 & ~n77214;
  assign n77216 = n77135 & ~n77156;
  assign n77217 = ~n77215 & n77216;
  assign n77218 = ~n77156 & n77190;
  assign n77219 = n77129 & n77218;
  assign n77220 = ~n77147 & ~n77162;
  assign n77221 = n77129 & n77165;
  assign n77222 = ~n77220 & ~n77221;
  assign n77223 = ~n77135 & ~n77222;
  assign n77224 = ~n77179 & ~n77223;
  assign n77225 = ~n77156 & ~n77224;
  assign n77226 = ~n77219 & ~n77225;
  assign n77227 = n77129 & ~n77147;
  assign n77228 = ~n77162 & n77227;
  assign n77229 = ~n77180 & ~n77228;
  assign n77230 = ~n77135 & ~n77229;
  assign n77231 = n77226 & ~n77230;
  assign n77232 = n77129 & n77135;
  assign n77233 = n77165 & n77232;
  assign n77234 = n77147 & n77233;
  assign n77235 = ~n77163 & ~n77167;
  assign n77236 = n77227 & ~n77235;
  assign n77237 = ~n77234 & ~n77236;
  assign n77238 = ~n77204 & n77237;
  assign n77239 = n77213 & ~n77235;
  assign n77240 = ~n77129 & n77192;
  assign n77241 = ~n77239 & ~n77240;
  assign n77242 = ~n77135 & n77213;
  assign n77243 = ~n77141 & n77242;
  assign n77244 = n77135 & n77166;
  assign n77245 = ~n77129 & n77244;
  assign n77246 = ~n77243 & ~n77245;
  assign n77247 = n77241 & n77246;
  assign n77248 = n77238 & n77247;
  assign n77249 = n77156 & ~n77248;
  assign n77250 = n77231 & ~n77249;
  assign n77251 = ~n77217 & n77250;
  assign n77252 = ~pi2441 & ~n77251;
  assign n77253 = pi2441 & n77231;
  assign n77254 = ~n77217 & n77253;
  assign n77255 = ~n77249 & n77254;
  assign po2544 = n77252 | n77255;
  assign n77257 = ~n77135 & n77172;
  assign n77258 = ~n77129 & n77257;
  assign n77259 = ~n77129 & ~n77135;
  assign n77260 = n77177 & n77259;
  assign n77261 = ~n77147 & n77260;
  assign n77262 = ~n77258 & ~n77261;
  assign n77263 = ~n77240 & ~n77245;
  assign n77264 = n77141 & n77147;
  assign n77265 = n77129 & n77264;
  assign n77266 = ~n77221 & ~n77265;
  assign n77267 = ~n77135 & ~n77266;
  assign n77268 = ~n77129 & ~n77147;
  assign n77269 = n77135 & ~n77268;
  assign n77270 = ~n77235 & n77269;
  assign n77271 = ~n77129 & ~n77165;
  assign n77272 = ~n77135 & n77271;
  assign n77273 = ~n77147 & n77272;
  assign n77274 = ~n77270 & ~n77273;
  assign n77275 = ~n77267 & n77274;
  assign n77276 = n77263 & n77275;
  assign n77277 = ~n77156 & ~n77276;
  assign n77278 = n77262 & ~n77277;
  assign n77279 = n77135 & n77164;
  assign n77280 = n77129 & n77279;
  assign n77281 = n77135 & n77156;
  assign n77282 = ~n77178 & ~n77221;
  assign n77283 = ~n77235 & n77268;
  assign n77284 = n77282 & ~n77283;
  assign n77285 = n77281 & ~n77284;
  assign n77286 = n77129 & n77192;
  assign n77287 = n77129 & n77141;
  assign n77288 = ~n77147 & n77287;
  assign n77289 = ~n77186 & ~n77288;
  assign n77290 = ~n77129 & n77165;
  assign n77291 = ~n77190 & ~n77290;
  assign n77292 = n77289 & n77291;
  assign n77293 = ~n77135 & ~n77292;
  assign n77294 = ~n77286 & ~n77293;
  assign n77295 = n77156 & ~n77294;
  assign n77296 = ~n77285 & ~n77295;
  assign n77297 = ~n77280 & n77296;
  assign n77298 = n77278 & n77297;
  assign n77299 = pi2445 & ~n77298;
  assign n77300 = ~pi2445 & n77278;
  assign n77301 = n77297 & n77300;
  assign po2545 = n77299 | n77301;
  assign n77303 = pi4820 & ~pi9040;
  assign n77304 = pi5186 & pi9040;
  assign n77305 = ~n77303 & ~n77304;
  assign n77306 = ~pi2397 & ~n77305;
  assign n77307 = pi2397 & n77305;
  assign n77308 = ~n77306 & ~n77307;
  assign n77309 = pi4859 & pi9040;
  assign n77310 = pi4970 & ~pi9040;
  assign n77311 = ~n77309 & ~n77310;
  assign n77312 = ~pi2383 & ~n77311;
  assign n77313 = pi2383 & n77311;
  assign n77314 = ~n77312 & ~n77313;
  assign n77315 = ~n77308 & ~n77314;
  assign n77316 = pi5090 & pi9040;
  assign n77317 = pi5210 & ~pi9040;
  assign n77318 = ~n77316 & ~n77317;
  assign n77319 = pi2365 & n77318;
  assign n77320 = ~pi2365 & ~n77318;
  assign n77321 = ~n77319 & ~n77320;
  assign n77322 = pi4859 & ~pi9040;
  assign n77323 = pi4824 & pi9040;
  assign n77324 = ~n77322 & ~n77323;
  assign n77325 = ~pi2380 & ~n77324;
  assign n77326 = pi2380 & n77324;
  assign n77327 = ~n77325 & ~n77326;
  assign n77328 = pi5090 & ~pi9040;
  assign n77329 = pi4952 & pi9040;
  assign n77330 = ~n77328 & ~n77329;
  assign n77331 = ~pi2376 & n77330;
  assign n77332 = pi2376 & ~n77330;
  assign n77333 = ~n77331 & ~n77332;
  assign n77334 = n77327 & n77333;
  assign n77335 = ~n77321 & n77334;
  assign n77336 = pi4939 & pi9040;
  assign n77337 = pi5081 & ~pi9040;
  assign n77338 = ~n77336 & ~n77337;
  assign n77339 = ~pi2377 & n77338;
  assign n77340 = pi2377 & ~n77338;
  assign n77341 = ~n77339 & ~n77340;
  assign n77342 = ~n77333 & n77341;
  assign n77343 = n77327 & n77342;
  assign n77344 = n77321 & n77343;
  assign n77345 = ~n77333 & ~n77341;
  assign n77346 = ~n77321 & n77345;
  assign n77347 = ~n77344 & ~n77346;
  assign n77348 = ~n77335 & n77347;
  assign n77349 = n77315 & ~n77348;
  assign n77350 = ~n77327 & n77342;
  assign n77351 = n77327 & n77345;
  assign n77352 = ~n77350 & ~n77351;
  assign n77353 = ~n77321 & ~n77327;
  assign n77354 = n77341 & n77353;
  assign n77355 = n77333 & n77341;
  assign n77356 = n77327 & n77355;
  assign n77357 = n77321 & n77356;
  assign n77358 = ~n77354 & ~n77357;
  assign n77359 = n77352 & n77358;
  assign n77360 = n77308 & ~n77359;
  assign n77361 = n77333 & ~n77341;
  assign n77362 = ~n77327 & n77361;
  assign n77363 = n77321 & n77362;
  assign n77364 = ~n77360 & ~n77363;
  assign n77365 = ~n77314 & ~n77364;
  assign n77366 = ~n77349 & ~n77365;
  assign n77367 = n77308 & ~n77321;
  assign n77368 = n77327 & n77367;
  assign n77369 = ~n77341 & n77368;
  assign n77370 = ~n77333 & n77354;
  assign n77371 = ~n77369 & ~n77370;
  assign n77372 = ~n77327 & n77355;
  assign n77373 = ~n77345 & ~n77355;
  assign n77374 = n77321 & ~n77373;
  assign n77375 = ~n77372 & ~n77374;
  assign n77376 = ~n77308 & ~n77375;
  assign n77377 = n77327 & n77361;
  assign n77378 = ~n77335 & ~n77377;
  assign n77379 = ~n77344 & n77378;
  assign n77380 = n77308 & ~n77379;
  assign n77381 = ~n77376 & ~n77380;
  assign n77382 = ~n77308 & ~n77321;
  assign n77383 = n77342 & n77382;
  assign n77384 = n77321 & n77372;
  assign n77385 = ~n77327 & ~n77333;
  assign n77386 = ~n77341 & n77385;
  assign n77387 = n77321 & n77386;
  assign n77388 = ~n77384 & ~n77387;
  assign n77389 = ~n77341 & n77353;
  assign n77390 = n77333 & n77389;
  assign n77391 = n77388 & ~n77390;
  assign n77392 = ~n77383 & n77391;
  assign n77393 = n77381 & n77392;
  assign n77394 = n77314 & ~n77393;
  assign n77395 = n77371 & ~n77394;
  assign n77396 = n77366 & n77395;
  assign n77397 = pi2414 & ~n77396;
  assign n77398 = ~pi2414 & n77371;
  assign n77399 = n77366 & n77398;
  assign n77400 = ~n77394 & n77399;
  assign po2546 = n77397 | n77400;
  assign n77402 = ~n77308 & n77372;
  assign n77403 = ~n77321 & n77402;
  assign n77404 = ~n77321 & n77343;
  assign n77405 = ~n77308 & n77404;
  assign n77406 = ~n77403 & ~n77405;
  assign n77407 = n77308 & n77390;
  assign n77408 = n77406 & ~n77407;
  assign n77409 = n77333 & n77367;
  assign n77410 = n77321 & n77334;
  assign n77411 = ~n77321 & ~n77333;
  assign n77412 = n77327 & n77411;
  assign n77413 = ~n77410 & ~n77412;
  assign n77414 = ~n77308 & ~n77413;
  assign n77415 = ~n77383 & ~n77414;
  assign n77416 = ~n77387 & ~n77404;
  assign n77417 = n77308 & n77321;
  assign n77418 = n77385 & n77417;
  assign n77419 = n77308 & n77362;
  assign n77420 = ~n77418 & ~n77419;
  assign n77421 = n77416 & n77420;
  assign n77422 = n77415 & n77421;
  assign n77423 = ~n77409 & n77422;
  assign n77424 = ~n77314 & ~n77423;
  assign n77425 = ~n77351 & ~n77410;
  assign n77426 = ~n77370 & n77425;
  assign n77427 = n77308 & ~n77426;
  assign n77428 = ~n77321 & n77386;
  assign n77429 = ~n77321 & n77377;
  assign n77430 = ~n77327 & n77333;
  assign n77431 = ~n77342 & ~n77430;
  assign n77432 = n77321 & ~n77431;
  assign n77433 = ~n77429 & ~n77432;
  assign n77434 = ~n77428 & n77433;
  assign n77435 = ~n77308 & ~n77434;
  assign n77436 = ~n77427 & ~n77435;
  assign n77437 = n77314 & ~n77436;
  assign n77438 = ~n77321 & n77327;
  assign n77439 = n77341 & n77438;
  assign n77440 = n77333 & n77439;
  assign n77441 = n77321 & n77345;
  assign n77442 = ~n77440 & ~n77441;
  assign n77443 = n77308 & ~n77442;
  assign n77444 = ~n77437 & ~n77443;
  assign n77445 = ~n77424 & n77444;
  assign n77446 = n77408 & n77445;
  assign n77447 = ~pi2419 & ~n77446;
  assign n77448 = pi2419 & n77446;
  assign po2548 = n77447 | n77448;
  assign n77450 = ~n76881 & n76906;
  assign n77451 = ~n76925 & ~n76939;
  assign n77452 = n77450 & ~n77451;
  assign n77453 = ~n76881 & ~n76900;
  assign n77454 = n76925 & n77453;
  assign n77455 = ~n77452 & ~n77454;
  assign n77456 = n76918 & ~n77455;
  assign n77457 = n76900 & ~n76906;
  assign n77458 = ~n76893 & n77457;
  assign n77459 = n76887 & n77458;
  assign n77460 = ~n76956 & ~n77457;
  assign n77461 = n76881 & ~n77460;
  assign n77462 = ~n76900 & ~n76906;
  assign n77463 = n76893 & n77462;
  assign n77464 = n76887 & n77463;
  assign n77465 = ~n77461 & ~n77464;
  assign n77466 = ~n77459 & n77465;
  assign n77467 = n76918 & ~n77466;
  assign n77468 = ~n77456 & ~n77467;
  assign n77469 = ~n76893 & n76907;
  assign n77470 = ~n76887 & n77469;
  assign n77471 = ~n76906 & n76932;
  assign n77472 = ~n77470 & ~n77471;
  assign n77473 = ~n76881 & ~n77472;
  assign n77474 = n76906 & n76945;
  assign n77475 = ~n76906 & n76956;
  assign n77476 = ~n77474 & ~n77475;
  assign n77477 = n76881 & ~n77476;
  assign n77478 = ~n76894 & ~n76956;
  assign n77479 = n76906 & ~n77478;
  assign n77480 = ~n76932 & ~n77479;
  assign n77481 = ~n76881 & ~n77480;
  assign n77482 = ~n76893 & ~n76906;
  assign n77483 = n77453 & n77482;
  assign n77484 = n76893 & n76900;
  assign n77485 = ~n76932 & ~n77484;
  assign n77486 = ~n76906 & ~n77485;
  assign n77487 = n76881 & n76906;
  assign n77488 = n76922 & n77487;
  assign n77489 = ~n76900 & n77488;
  assign n77490 = ~n77486 & ~n77489;
  assign n77491 = ~n77483 & n77490;
  assign n77492 = ~n77481 & n77491;
  assign n77493 = ~n77470 & n77492;
  assign n77494 = ~n76918 & ~n77493;
  assign n77495 = ~n77477 & ~n77494;
  assign n77496 = ~n77473 & n77495;
  assign n77497 = n77468 & n77496;
  assign n77498 = pi2406 & n77497;
  assign n77499 = ~pi2406 & ~n77497;
  assign po2549 = n77498 | n77499;
  assign n77501 = n76893 & n76909;
  assign n77502 = ~n76939 & ~n77501;
  assign n77503 = ~n76881 & ~n77502;
  assign n77504 = n76906 & n76931;
  assign n77505 = n76893 & ~n76906;
  assign n77506 = ~n76900 & n77505;
  assign n77507 = ~n77504 & ~n77506;
  assign n77508 = n76881 & ~n77507;
  assign n77509 = ~n76906 & n76926;
  assign n77510 = ~n77483 & ~n77509;
  assign n77511 = ~n76908 & n77510;
  assign n77512 = ~n77508 & n77511;
  assign n77513 = ~n77503 & n77512;
  assign n77514 = ~n77459 & ~n77470;
  assign n77515 = n77513 & n77514;
  assign n77516 = n76918 & ~n77515;
  assign n77517 = n76894 & n77457;
  assign n77518 = n76946 & ~n77517;
  assign n77519 = n76881 & ~n77518;
  assign n77520 = ~n76906 & n76936;
  assign n77521 = ~n77519 & ~n77520;
  assign n77522 = n76887 & n76909;
  assign n77523 = n76906 & n76922;
  assign n77524 = ~n77522 & ~n77523;
  assign n77525 = n76881 & ~n77524;
  assign n77526 = n76881 & n76931;
  assign n77527 = ~n76906 & n77526;
  assign n77528 = ~n77525 & ~n77527;
  assign n77529 = n77521 & n77528;
  assign n77530 = ~n76918 & ~n77529;
  assign n77531 = ~n76926 & ~n76933;
  assign n77532 = ~n77464 & n77531;
  assign n77533 = n76953 & ~n77532;
  assign n77534 = ~n77530 & ~n77533;
  assign n77535 = ~n76908 & ~n77459;
  assign n77536 = ~n76881 & ~n77535;
  assign n77537 = n77534 & ~n77536;
  assign n77538 = ~n77516 & n77537;
  assign n77539 = ~pi2416 & n77538;
  assign n77540 = pi2416 & ~n77538;
  assign po2550 = n77539 | n77540;
  assign n77542 = ~n77186 & ~n77290;
  assign n77543 = ~n77135 & ~n77542;
  assign n77544 = ~n77261 & ~n77543;
  assign n77545 = ~n77156 & ~n77544;
  assign n77546 = n77163 & n77227;
  assign n77547 = ~n77135 & n77546;
  assign n77548 = n77147 & n77232;
  assign n77549 = n77162 & n77548;
  assign n77550 = ~n77547 & ~n77549;
  assign n77551 = ~n77190 & ~n77287;
  assign n77552 = n77216 & ~n77551;
  assign n77553 = ~n77163 & n77202;
  assign n77554 = ~n77156 & n77553;
  assign n77555 = ~n77552 & ~n77554;
  assign n77556 = n77550 & n77555;
  assign n77557 = n77129 & n77166;
  assign n77558 = n77162 & n77213;
  assign n77559 = ~n77148 & ~n77163;
  assign n77560 = n77129 & ~n77559;
  assign n77561 = ~n77558 & ~n77560;
  assign n77562 = ~n77135 & ~n77561;
  assign n77563 = ~n77557 & ~n77562;
  assign n77564 = ~n77129 & ~n77559;
  assign n77565 = ~n77172 & ~n77564;
  assign n77566 = n77135 & ~n77565;
  assign n77567 = ~n77283 & ~n77566;
  assign n77568 = n77563 & n77567;
  assign n77569 = n77156 & ~n77568;
  assign n77570 = n77556 & ~n77569;
  assign n77571 = ~n77545 & n77570;
  assign n77572 = pi2446 & ~n77571;
  assign n77573 = ~pi2446 & n77571;
  assign po2552 = n77572 | n77573;
  assign n77575 = n76656 & n76702;
  assign n77576 = n76656 & n76667;
  assign n77577 = ~n77575 & ~n77576;
  assign n77578 = ~n76648 & ~n77577;
  assign n77579 = n76714 & n76720;
  assign n77580 = ~n77578 & ~n77579;
  assign n77581 = ~n76733 & n77580;
  assign n77582 = ~n76656 & n76670;
  assign n77583 = ~n76667 & ~n77582;
  assign n77584 = n76642 & n76673;
  assign n77585 = n77583 & ~n77584;
  assign n77586 = ~n76648 & ~n77585;
  assign n77587 = n76687 & n77586;
  assign n77588 = n76642 & n76666;
  assign n77589 = n76648 & n77588;
  assign n77590 = ~n76691 & ~n76710;
  assign n77591 = ~n76704 & n77590;
  assign n77592 = ~n77589 & n77591;
  assign n77593 = n76687 & ~n77592;
  assign n77594 = n76642 & ~n76656;
  assign n77595 = ~n76665 & n77594;
  assign n77596 = n76642 & n76648;
  assign n77597 = n76665 & n77596;
  assign n77598 = ~n76636 & n77597;
  assign n77599 = ~n76656 & n76678;
  assign n77600 = ~n77598 & ~n77599;
  assign n77601 = ~n77595 & n77600;
  assign n77602 = n76665 & n76708;
  assign n77603 = ~n76656 & n76695;
  assign n77604 = ~n76713 & ~n77603;
  assign n77605 = ~n76648 & ~n77604;
  assign n77606 = ~n77602 & ~n77605;
  assign n77607 = n77601 & n77606;
  assign n77608 = ~n76687 & ~n77607;
  assign n77609 = n76656 & n77598;
  assign n77610 = ~n77608 & ~n77609;
  assign n77611 = ~n77593 & n77610;
  assign n77612 = ~n77587 & n77611;
  assign n77613 = n77581 & n77612;
  assign n77614 = pi2412 & ~n77613;
  assign n77615 = ~pi2412 & n77581;
  assign n77616 = n77612 & n77615;
  assign po2553 = n77614 | n77616;
  assign n77618 = n77308 & n77345;
  assign n77619 = ~n77321 & n77618;
  assign n77620 = ~n77440 & ~n77619;
  assign n77621 = n77321 & ~n77341;
  assign n77622 = n77327 & n77621;
  assign n77623 = ~n77321 & n77333;
  assign n77624 = ~n77439 & ~n77623;
  assign n77625 = ~n77308 & ~n77624;
  assign n77626 = ~n77622 & ~n77625;
  assign n77627 = n77620 & n77626;
  assign n77628 = n77314 & ~n77627;
  assign n77629 = ~n77343 & ~n77387;
  assign n77630 = ~n77321 & n77361;
  assign n77631 = n77629 & ~n77630;
  assign n77632 = n77308 & ~n77631;
  assign n77633 = ~n77308 & n77346;
  assign n77634 = ~n77370 & ~n77633;
  assign n77635 = ~n77632 & n77634;
  assign n77636 = ~n77356 & ~n77363;
  assign n77637 = ~n77308 & ~n77636;
  assign n77638 = n77635 & ~n77637;
  assign n77639 = ~n77314 & ~n77638;
  assign n77640 = ~n77628 & ~n77639;
  assign n77641 = ~n77321 & n77355;
  assign n77642 = n77321 & ~n77352;
  assign n77643 = ~n77641 & ~n77642;
  assign n77644 = ~n77308 & ~n77643;
  assign n77645 = ~n77372 & ~n77377;
  assign n77646 = ~n77343 & n77645;
  assign n77647 = n77417 & ~n77646;
  assign n77648 = ~n77644 & ~n77647;
  assign n77649 = n77640 & n77648;
  assign n77650 = ~pi2415 & ~n77649;
  assign n77651 = ~n77639 & n77648;
  assign n77652 = pi2415 & n77651;
  assign n77653 = ~n77628 & n77652;
  assign po2554 = n77650 | n77653;
  assign n77655 = ~n77064 & ~n77069;
  assign n77656 = ~n76751 & n76788;
  assign n77657 = ~n77057 & ~n77656;
  assign n77658 = ~n77042 & n77657;
  assign n77659 = ~n76785 & ~n77658;
  assign n77660 = n76751 & n76795;
  assign n77661 = ~n76763 & n76802;
  assign n77662 = ~n76820 & ~n77661;
  assign n77663 = n76785 & ~n77662;
  assign n77664 = ~n77660 & ~n77663;
  assign n77665 = ~n76785 & n76786;
  assign n77666 = n76751 & n77665;
  assign n77667 = ~n76785 & n76793;
  assign n77668 = ~n77666 & ~n77667;
  assign n77669 = n77664 & n77668;
  assign n77670 = ~n76763 & n76807;
  assign n77671 = ~n77042 & ~n77670;
  assign n77672 = ~n77078 & n77671;
  assign n77673 = n77669 & n77672;
  assign n77674 = ~n76745 & ~n77673;
  assign n77675 = n76774 & n76785;
  assign n77676 = ~n76835 & n77657;
  assign n77677 = ~n76809 & ~n76820;
  assign n77678 = ~n77074 & n77677;
  assign n77679 = ~n76785 & ~n77678;
  assign n77680 = n77676 & ~n77679;
  assign n77681 = ~n77675 & n77680;
  assign n77682 = n76745 & ~n77681;
  assign n77683 = ~n77674 & ~n77682;
  assign n77684 = ~n77659 & n77683;
  assign n77685 = n77655 & n77684;
  assign n77686 = pi2403 & ~n77685;
  assign n77687 = ~pi2403 & n77685;
  assign po2555 = n77686 | n77687;
  assign n77689 = ~n76636 & n76642;
  assign n77690 = ~n76710 & ~n77689;
  assign n77691 = ~n76657 & n77690;
  assign n77692 = n76648 & ~n77691;
  assign n77693 = n76636 & n76720;
  assign n77694 = ~n77575 & ~n77595;
  assign n77695 = ~n76636 & ~n76642;
  assign n77696 = ~n76648 & n76656;
  assign n77697 = n77695 & n77696;
  assign n77698 = n77694 & ~n77697;
  assign n77699 = ~n77693 & n77698;
  assign n77700 = ~n77692 & n77699;
  assign n77701 = n76687 & ~n77700;
  assign n77702 = ~n76656 & n77584;
  assign n77703 = n76656 & n77588;
  assign n77704 = ~n77702 & ~n77703;
  assign n77705 = n76648 & ~n77704;
  assign n77706 = ~n77701 & ~n77705;
  assign n77707 = ~n76656 & n76702;
  assign n77708 = ~n76670 & ~n76714;
  assign n77709 = n76648 & ~n77708;
  assign n77710 = ~n77707 & ~n77709;
  assign n77711 = ~n76717 & n77710;
  assign n77712 = ~n76687 & ~n77711;
  assign n77713 = ~n76673 & ~n76695;
  assign n77714 = ~n76642 & ~n77713;
  assign n77715 = ~n76723 & ~n77714;
  assign n77716 = ~n76648 & ~n77715;
  assign n77717 = ~n76687 & n77716;
  assign n77718 = ~n77712 & ~n77717;
  assign n77719 = n77706 & n77718;
  assign n77720 = pi2405 & ~n77719;
  assign n77721 = ~pi2405 & n77706;
  assign n77722 = n77718 & n77721;
  assign po2556 = n77720 | n77722;
  assign n77724 = ~n76772 & ~n76803;
  assign n77725 = n76745 & ~n77724;
  assign n77726 = ~n76808 & ~n77048;
  assign n77727 = ~n76778 & n77726;
  assign n77728 = ~n76785 & ~n77727;
  assign n77729 = n76745 & n77728;
  assign n77730 = ~n77725 & ~n77729;
  assign n77731 = n76771 & n77051;
  assign n77732 = ~n77053 & ~n77731;
  assign n77733 = ~n76811 & ~n77075;
  assign n77734 = n76785 & ~n77733;
  assign n77735 = n76745 & n77734;
  assign n77736 = n77732 & ~n77735;
  assign n77737 = n76751 & n76771;
  assign n77738 = n76751 & n76773;
  assign n77739 = ~n77044 & ~n77738;
  assign n77740 = n76785 & ~n77739;
  assign n77741 = ~n76809 & ~n77057;
  assign n77742 = n76751 & n76770;
  assign n77743 = ~n76833 & ~n77742;
  assign n77744 = ~n76785 & ~n77743;
  assign n77745 = n77741 & ~n77744;
  assign n77746 = ~n77740 & n77745;
  assign n77747 = ~n77737 & n77746;
  assign n77748 = ~n76745 & ~n77747;
  assign n77749 = ~n77078 & n77657;
  assign n77750 = n76785 & ~n77749;
  assign n77751 = ~n77748 & ~n77750;
  assign n77752 = n77736 & n77751;
  assign n77753 = n77730 & n77752;
  assign n77754 = ~pi2411 & ~n77753;
  assign n77755 = pi2411 & n77736;
  assign n77756 = n77730 & n77755;
  assign n77757 = n77751 & n77756;
  assign po2557 = n77754 | n77757;
  assign n77759 = pi4893 & pi9040;
  assign n77760 = pi4824 & ~pi9040;
  assign n77761 = ~n77759 & ~n77760;
  assign n77762 = ~pi2376 & ~n77761;
  assign n77763 = pi2376 & n77761;
  assign n77764 = ~n77762 & ~n77763;
  assign n77765 = pi4855 & ~pi9040;
  assign n77766 = pi4868 & pi9040;
  assign n77767 = ~n77765 & ~n77766;
  assign n77768 = pi2399 & n77767;
  assign n77769 = ~pi2399 & ~n77767;
  assign n77770 = ~n77768 & ~n77769;
  assign n77771 = pi4759 & ~pi9040;
  assign n77772 = pi5081 & pi9040;
  assign n77773 = ~n77771 & ~n77772;
  assign n77774 = ~pi2395 & ~n77773;
  assign n77775 = pi2395 & n77773;
  assign n77776 = ~n77774 & ~n77775;
  assign n77777 = pi4855 & pi9040;
  assign n77778 = pi5186 & ~pi9040;
  assign n77779 = ~n77777 & ~n77778;
  assign n77780 = ~pi2386 & ~n77779;
  assign n77781 = pi2386 & n77779;
  assign n77782 = ~n77780 & ~n77781;
  assign n77783 = pi4939 & ~pi9040;
  assign n77784 = pi4826 & pi9040;
  assign n77785 = ~n77783 & ~n77784;
  assign n77786 = pi2380 & n77785;
  assign n77787 = ~pi2380 & ~n77785;
  assign n77788 = ~n77786 & ~n77787;
  assign n77789 = n77782 & ~n77788;
  assign n77790 = n77776 & n77789;
  assign n77791 = n77770 & n77790;
  assign n77792 = ~n77770 & n77782;
  assign n77793 = n77788 & n77792;
  assign n77794 = pi4952 & ~pi9040;
  assign n77795 = pi4819 & pi9040;
  assign n77796 = ~n77794 & ~n77795;
  assign n77797 = ~pi2355 & n77796;
  assign n77798 = pi2355 & ~n77796;
  assign n77799 = ~n77797 & ~n77798;
  assign n77800 = ~n77776 & n77792;
  assign n77801 = n77776 & n77788;
  assign n77802 = ~n77782 & n77801;
  assign n77803 = ~n77800 & ~n77802;
  assign n77804 = n77799 & ~n77803;
  assign n77805 = ~n77793 & ~n77804;
  assign n77806 = n77782 & n77801;
  assign n77807 = ~n77776 & ~n77782;
  assign n77808 = ~n77782 & ~n77788;
  assign n77809 = ~n77770 & n77808;
  assign n77810 = ~n77776 & ~n77788;
  assign n77811 = n77770 & n77810;
  assign n77812 = ~n77809 & ~n77811;
  assign n77813 = ~n77807 & n77812;
  assign n77814 = ~n77806 & n77813;
  assign n77815 = ~n77799 & ~n77814;
  assign n77816 = n77805 & ~n77815;
  assign n77817 = ~n77791 & n77816;
  assign n77818 = n77764 & ~n77817;
  assign n77819 = ~n77776 & n77788;
  assign n77820 = ~n77782 & n77819;
  assign n77821 = ~n77770 & n77820;
  assign n77822 = ~n77788 & n77807;
  assign n77823 = n77770 & n77822;
  assign n77824 = ~n77791 & ~n77823;
  assign n77825 = ~n77821 & n77824;
  assign n77826 = ~n77799 & ~n77825;
  assign n77827 = ~n77818 & ~n77826;
  assign n77828 = n77776 & n77793;
  assign n77829 = n77776 & ~n77782;
  assign n77830 = n77799 & n77829;
  assign n77831 = n77770 & n77830;
  assign n77832 = n77782 & n77819;
  assign n77833 = n77770 & n77832;
  assign n77834 = n77789 & ~n77799;
  assign n77835 = ~n77770 & n77834;
  assign n77836 = ~n77833 & ~n77835;
  assign n77837 = ~n77776 & n77782;
  assign n77838 = n77770 & n77837;
  assign n77839 = n77776 & ~n77788;
  assign n77840 = ~n77782 & n77839;
  assign n77841 = ~n77838 & ~n77840;
  assign n77842 = n77799 & ~n77841;
  assign n77843 = n77799 & n77807;
  assign n77844 = ~n77770 & n77843;
  assign n77845 = ~n77842 & ~n77844;
  assign n77846 = n77836 & n77845;
  assign n77847 = ~n77764 & ~n77846;
  assign n77848 = ~n77831 & ~n77847;
  assign n77849 = ~n77828 & n77848;
  assign n77850 = n77827 & n77849;
  assign n77851 = ~pi2409 & ~n77850;
  assign n77852 = ~n77818 & ~n77828;
  assign n77853 = ~n77826 & n77852;
  assign n77854 = n77848 & n77853;
  assign n77855 = pi2409 & n77854;
  assign po2558 = n77851 | n77855;
  assign n77857 = ~n76656 & n77714;
  assign n77858 = ~n76669 & ~n77588;
  assign n77859 = ~n76648 & ~n77858;
  assign n77860 = ~n77857 & ~n77859;
  assign n77861 = n76665 & n77594;
  assign n77862 = ~n76675 & ~n77861;
  assign n77863 = ~n77584 & n77862;
  assign n77864 = n76648 & ~n77863;
  assign n77865 = n77860 & ~n77864;
  assign n77866 = n76656 & n76714;
  assign n77867 = n77865 & ~n77866;
  assign n77868 = ~n76687 & ~n77867;
  assign n77869 = ~n76667 & ~n76670;
  assign n77870 = ~n76714 & ~n77584;
  assign n77871 = n77869 & n77870;
  assign n77872 = ~n76656 & ~n77871;
  assign n77873 = n76696 & ~n77858;
  assign n77874 = ~n77872 & ~n77873;
  assign n77875 = ~n77575 & n77874;
  assign n77876 = n76687 & ~n77875;
  assign n77877 = ~n77868 & ~n77876;
  assign n77878 = ~n76656 & n77588;
  assign n77879 = ~n77866 & ~n77878;
  assign n77880 = ~n76648 & ~n77879;
  assign n77881 = n77877 & ~n77880;
  assign n77882 = pi2404 & ~n77881;
  assign n77883 = ~pi2404 & ~n77880;
  assign n77884 = ~n77876 & n77883;
  assign n77885 = ~n77868 & n77884;
  assign po2559 = n77882 | n77885;
  assign n77887 = ~n76906 & n76922;
  assign n77888 = ~n76921 & ~n77887;
  assign n77889 = ~n76881 & ~n77888;
  assign n77890 = n76881 & ~n77485;
  assign n77891 = ~n77474 & ~n77890;
  assign n77892 = ~n77889 & n77891;
  assign n77893 = n76918 & ~n77892;
  assign n77894 = ~n76881 & n76936;
  assign n77895 = ~n77893 & ~n77894;
  assign n77896 = ~n77509 & ~n77523;
  assign n77897 = n76881 & ~n77896;
  assign n77898 = n76881 & n76923;
  assign n77899 = n76906 & n76939;
  assign n77900 = ~n76881 & n76907;
  assign n77901 = ~n77462 & ~n77900;
  assign n77902 = ~n76887 & ~n77901;
  assign n77903 = ~n77506 & ~n77902;
  assign n77904 = ~n76908 & n77903;
  assign n77905 = ~n77899 & n77904;
  assign n77906 = ~n77898 & n77905;
  assign n77907 = ~n76918 & ~n77906;
  assign n77908 = ~n77897 & ~n77907;
  assign n77909 = n77895 & n77908;
  assign n77910 = pi2422 & ~n77909;
  assign n77911 = ~pi2422 & n77909;
  assign po2560 = n77910 | n77911;
  assign n77913 = ~n77308 & ~n77645;
  assign n77914 = n77321 & n77351;
  assign n77915 = ~n77913 & ~n77914;
  assign n77916 = n77321 & ~n77333;
  assign n77917 = ~n77385 & ~n77916;
  assign n77918 = ~n77356 & n77917;
  assign n77919 = n77308 & ~n77918;
  assign n77920 = n77915 & ~n77919;
  assign n77921 = ~n77314 & ~n77920;
  assign n77922 = ~n77308 & n77428;
  assign n77923 = ~n77405 & ~n77922;
  assign n77924 = ~n77407 & n77923;
  assign n77925 = ~n77390 & ~n77439;
  assign n77926 = n77308 & n77412;
  assign n77927 = n77321 & n77377;
  assign n77928 = ~n77308 & n77385;
  assign n77929 = ~n77927 & ~n77928;
  assign n77930 = ~n77384 & n77929;
  assign n77931 = ~n77926 & n77930;
  assign n77932 = n77925 & n77931;
  assign n77933 = ~n77419 & n77932;
  assign n77934 = n77314 & ~n77933;
  assign n77935 = n77924 & ~n77934;
  assign n77936 = ~n77921 & n77935;
  assign n77937 = ~pi2427 & ~n77936;
  assign n77938 = pi2427 & n77924;
  assign n77939 = ~n77921 & n77938;
  assign n77940 = ~n77934 & n77939;
  assign po2562 = n77937 | n77940;
  assign n77942 = n77782 & n77810;
  assign n77943 = ~n77770 & n77942;
  assign n77944 = ~n77820 & ~n77828;
  assign n77945 = n77770 & n77789;
  assign n77946 = ~n77770 & n77840;
  assign n77947 = ~n77945 & ~n77946;
  assign n77948 = n77944 & n77947;
  assign n77949 = n77799 & ~n77948;
  assign n77950 = ~n77782 & n77810;
  assign n77951 = n77770 & n77801;
  assign n77952 = ~n77800 & ~n77951;
  assign n77953 = ~n77950 & n77952;
  assign n77954 = ~n77799 & ~n77953;
  assign n77955 = n77770 & n77802;
  assign n77956 = ~n77954 & ~n77955;
  assign n77957 = ~n77949 & n77956;
  assign n77958 = ~n77943 & n77957;
  assign n77959 = ~n77764 & ~n77958;
  assign n77960 = n77770 & n77799;
  assign n77961 = n77806 & n77960;
  assign n77962 = n77799 & n77950;
  assign n77963 = n77799 & n77832;
  assign n77964 = ~n77962 & ~n77963;
  assign n77965 = ~n77770 & ~n77964;
  assign n77966 = ~n77961 & ~n77965;
  assign n77967 = ~n77770 & n77790;
  assign n77968 = n77770 & n77840;
  assign n77969 = ~n77967 & ~n77968;
  assign n77970 = n77770 & n77819;
  assign n77971 = ~n77770 & n77801;
  assign n77972 = ~n77970 & ~n77971;
  assign n77973 = ~n77790 & n77972;
  assign n77974 = ~n77820 & n77973;
  assign n77975 = ~n77799 & ~n77974;
  assign n77976 = ~n77770 & n77802;
  assign n77977 = ~n77975 & ~n77976;
  assign n77978 = n77969 & n77977;
  assign n77979 = n77966 & n77978;
  assign n77980 = n77764 & ~n77979;
  assign n77981 = n77770 & n77942;
  assign n77982 = n77770 & n77820;
  assign n77983 = ~n77981 & ~n77982;
  assign n77984 = n77799 & ~n77983;
  assign n77985 = ~n77980 & ~n77984;
  assign n77986 = ~n77823 & ~n77967;
  assign n77987 = ~n77799 & ~n77986;
  assign n77988 = n77985 & ~n77987;
  assign n77989 = ~n77959 & n77988;
  assign n77990 = pi2410 & ~n77989;
  assign n77991 = ~pi2410 & n77989;
  assign po2563 = n77990 | n77991;
  assign n77993 = ~n77770 & n77799;
  assign n77994 = n77776 & n77993;
  assign n77995 = ~n77770 & ~n77782;
  assign n77996 = ~n77788 & n77995;
  assign n77997 = ~n77776 & n77996;
  assign n77998 = ~n77802 & ~n77997;
  assign n77999 = ~n77799 & ~n77998;
  assign n78000 = n77983 & ~n77999;
  assign n78001 = ~n77994 & n78000;
  assign n78002 = n77764 & ~n78001;
  assign n78003 = n77799 & n77968;
  assign n78004 = ~n77770 & ~n77799;
  assign n78005 = n77840 & n78004;
  assign n78006 = ~n77800 & ~n78005;
  assign n78007 = ~n77802 & ~n77832;
  assign n78008 = ~n77770 & n77819;
  assign n78009 = n78007 & ~n78008;
  assign n78010 = n77799 & ~n78009;
  assign n78011 = ~n77799 & n77806;
  assign n78012 = n77824 & ~n78011;
  assign n78013 = ~n78010 & n78012;
  assign n78014 = n78006 & n78013;
  assign n78015 = ~n77764 & ~n78014;
  assign n78016 = ~n78003 & ~n78015;
  assign n78017 = ~n78002 & n78016;
  assign n78018 = n77832 & n78004;
  assign n78019 = n77770 & n77834;
  assign n78020 = ~n78018 & ~n78019;
  assign n78021 = ~n77799 & n77982;
  assign n78022 = n78020 & ~n78021;
  assign n78023 = n78017 & n78022;
  assign n78024 = ~pi2413 & ~n78023;
  assign n78025 = pi2413 & n78022;
  assign n78026 = n78016 & n78025;
  assign n78027 = ~n78002 & n78026;
  assign po2564 = n78024 | n78027;
  assign n78029 = ~n77967 & ~n77997;
  assign n78030 = ~n77955 & n78029;
  assign n78031 = n77799 & ~n78030;
  assign n78032 = ~n78005 & ~n78021;
  assign n78033 = ~n77963 & ~n77968;
  assign n78034 = ~n77942 & ~n77971;
  assign n78035 = ~n77799 & ~n78034;
  assign n78036 = ~n77828 & ~n78035;
  assign n78037 = n78033 & n78036;
  assign n78038 = n77764 & ~n78037;
  assign n78039 = ~n77782 & n77788;
  assign n78040 = ~n77807 & ~n78039;
  assign n78041 = n77770 & ~n78040;
  assign n78042 = ~n77790 & ~n78008;
  assign n78043 = ~n77799 & ~n78042;
  assign n78044 = n77770 & n77788;
  assign n78045 = ~n77802 & ~n78044;
  assign n78046 = ~n77810 & n78045;
  assign n78047 = n77799 & ~n78046;
  assign n78048 = ~n78043 & ~n78047;
  assign n78049 = ~n78041 & n78048;
  assign n78050 = ~n77764 & ~n78049;
  assign n78051 = ~n78038 & ~n78050;
  assign n78052 = n78032 & n78051;
  assign n78053 = ~n78031 & n78052;
  assign n78054 = ~pi2418 & ~n78053;
  assign n78055 = pi2418 & n78032;
  assign n78056 = ~n78031 & n78055;
  assign n78057 = n78051 & n78056;
  assign po2565 = n78054 | n78057;
  assign n78059 = pi5104 & pi9040;
  assign n78060 = pi4989 & ~pi9040;
  assign n78061 = ~n78059 & ~n78060;
  assign n78062 = pi2440 & n78061;
  assign n78063 = ~pi2440 & ~n78061;
  assign n78064 = ~n78062 & ~n78063;
  assign n78065 = pi5102 & pi9040;
  assign n78066 = pi5053 & ~pi9040;
  assign n78067 = ~n78065 & ~n78066;
  assign n78068 = ~pi2461 & ~n78067;
  assign n78069 = pi2461 & n78067;
  assign n78070 = ~n78068 & ~n78069;
  assign n78071 = ~n78064 & ~n78070;
  assign n78072 = pi5107 & ~pi9040;
  assign n78073 = pi5418 & pi9040;
  assign n78074 = ~n78072 & ~n78073;
  assign n78075 = ~pi2452 & ~n78074;
  assign n78076 = pi2452 & ~n78072;
  assign n78077 = ~n78073 & n78076;
  assign n78078 = ~n78075 & ~n78077;
  assign n78079 = pi5107 & pi9040;
  assign n78080 = pi5101 & ~pi9040;
  assign n78081 = ~n78079 & ~n78080;
  assign n78082 = ~pi2456 & ~n78081;
  assign n78083 = pi2456 & n78081;
  assign n78084 = ~n78082 & ~n78083;
  assign n78085 = pi4979 & pi9040;
  assign n78086 = pi5290 & ~pi9040;
  assign n78087 = ~n78085 & ~n78086;
  assign n78088 = ~pi2424 & ~n78087;
  assign n78089 = pi2424 & n78087;
  assign n78090 = ~n78088 & ~n78089;
  assign n78091 = n78084 & ~n78090;
  assign n78092 = ~n78078 & n78091;
  assign n78093 = pi5094 & ~pi9040;
  assign n78094 = pi5046 & pi9040;
  assign n78095 = ~n78093 & ~n78094;
  assign n78096 = pi2439 & n78095;
  assign n78097 = ~pi2439 & ~n78095;
  assign n78098 = ~n78096 & ~n78097;
  assign n78099 = n78090 & ~n78098;
  assign n78100 = n78084 & n78099;
  assign n78101 = n78078 & n78100;
  assign n78102 = n78090 & n78098;
  assign n78103 = ~n78078 & n78102;
  assign n78104 = ~n78101 & ~n78103;
  assign n78105 = ~n78092 & n78104;
  assign n78106 = n78071 & ~n78105;
  assign n78107 = ~n78078 & ~n78098;
  assign n78108 = ~n78084 & n78107;
  assign n78109 = ~n78090 & ~n78098;
  assign n78110 = n78084 & n78109;
  assign n78111 = n78078 & n78110;
  assign n78112 = ~n78108 & ~n78111;
  assign n78113 = ~n78084 & n78099;
  assign n78114 = n78084 & n78102;
  assign n78115 = ~n78113 & ~n78114;
  assign n78116 = n78112 & n78115;
  assign n78117 = n78064 & ~n78116;
  assign n78118 = ~n78090 & n78098;
  assign n78119 = ~n78084 & n78118;
  assign n78120 = n78078 & n78119;
  assign n78121 = ~n78117 & ~n78120;
  assign n78122 = ~n78070 & ~n78121;
  assign n78123 = ~n78106 & ~n78122;
  assign n78124 = n78064 & ~n78078;
  assign n78125 = n78084 & n78124;
  assign n78126 = n78098 & n78125;
  assign n78127 = ~n78078 & ~n78084;
  assign n78128 = ~n78098 & n78127;
  assign n78129 = n78090 & n78128;
  assign n78130 = ~n78126 & ~n78129;
  assign n78131 = ~n78102 & ~n78109;
  assign n78132 = n78078 & ~n78131;
  assign n78133 = ~n78084 & n78109;
  assign n78134 = ~n78132 & ~n78133;
  assign n78135 = ~n78064 & ~n78134;
  assign n78136 = n78084 & n78118;
  assign n78137 = ~n78092 & ~n78136;
  assign n78138 = ~n78101 & n78137;
  assign n78139 = n78064 & ~n78138;
  assign n78140 = ~n78135 & ~n78139;
  assign n78141 = ~n78064 & ~n78078;
  assign n78142 = n78099 & n78141;
  assign n78143 = n78078 & ~n78084;
  assign n78144 = ~n78098 & n78143;
  assign n78145 = ~n78090 & n78144;
  assign n78146 = ~n78084 & n78090;
  assign n78147 = n78098 & n78146;
  assign n78148 = n78078 & n78147;
  assign n78149 = ~n78145 & ~n78148;
  assign n78150 = n78098 & n78127;
  assign n78151 = ~n78090 & n78150;
  assign n78152 = n78149 & ~n78151;
  assign n78153 = ~n78142 & n78152;
  assign n78154 = n78140 & n78153;
  assign n78155 = n78070 & ~n78154;
  assign n78156 = n78130 & ~n78155;
  assign n78157 = n78123 & n78156;
  assign n78158 = pi2475 & ~n78157;
  assign n78159 = ~pi2475 & n78130;
  assign n78160 = n78123 & n78159;
  assign n78161 = ~n78155 & n78160;
  assign po2576 = n78158 | n78161;
  assign n78163 = ~n78078 & n78147;
  assign n78164 = ~n78084 & ~n78090;
  assign n78165 = ~n78099 & ~n78164;
  assign n78166 = n78078 & ~n78165;
  assign n78167 = ~n78078 & n78136;
  assign n78168 = ~n78166 & ~n78167;
  assign n78169 = ~n78163 & n78168;
  assign n78170 = ~n78064 & ~n78169;
  assign n78171 = n78078 & n78091;
  assign n78172 = ~n78114 & ~n78171;
  assign n78173 = ~n78129 & n78172;
  assign n78174 = n78064 & ~n78173;
  assign n78175 = ~n78170 & ~n78174;
  assign n78176 = n78070 & ~n78175;
  assign n78177 = ~n78090 & n78124;
  assign n78178 = ~n78078 & n78090;
  assign n78179 = n78084 & n78178;
  assign n78180 = ~n78171 & ~n78179;
  assign n78181 = ~n78064 & ~n78180;
  assign n78182 = ~n78142 & ~n78181;
  assign n78183 = ~n78078 & n78100;
  assign n78184 = ~n78148 & ~n78183;
  assign n78185 = n78064 & n78078;
  assign n78186 = n78146 & n78185;
  assign n78187 = n78064 & n78119;
  assign n78188 = ~n78186 & ~n78187;
  assign n78189 = n78184 & n78188;
  assign n78190 = n78182 & n78189;
  assign n78191 = ~n78177 & n78190;
  assign n78192 = ~n78070 & ~n78191;
  assign n78193 = ~n78064 & n78133;
  assign n78194 = ~n78078 & n78193;
  assign n78195 = ~n78064 & n78183;
  assign n78196 = ~n78194 & ~n78195;
  assign n78197 = n78064 & n78151;
  assign n78198 = n78196 & ~n78197;
  assign n78199 = ~n78078 & n78110;
  assign n78200 = n78078 & n78102;
  assign n78201 = ~n78199 & ~n78200;
  assign n78202 = n78064 & ~n78201;
  assign n78203 = n78198 & ~n78202;
  assign n78204 = ~n78192 & n78203;
  assign n78205 = ~n78176 & n78204;
  assign n78206 = ~pi2474 & ~n78205;
  assign n78207 = pi2474 & n78205;
  assign po2582 = n78206 | n78207;
  assign n78209 = ~n78133 & ~n78136;
  assign n78210 = ~n78064 & ~n78209;
  assign n78211 = n78078 & n78114;
  assign n78212 = ~n78210 & ~n78211;
  assign n78213 = n78078 & n78090;
  assign n78214 = ~n78146 & ~n78213;
  assign n78215 = ~n78110 & n78214;
  assign n78216 = n78064 & ~n78215;
  assign n78217 = n78212 & ~n78216;
  assign n78218 = ~n78070 & ~n78217;
  assign n78219 = ~n78064 & n78163;
  assign n78220 = ~n78195 & ~n78219;
  assign n78221 = ~n78197 & n78220;
  assign n78222 = ~n78078 & n78084;
  assign n78223 = ~n78098 & n78222;
  assign n78224 = ~n78151 & ~n78223;
  assign n78225 = n78064 & n78179;
  assign n78226 = n78078 & n78136;
  assign n78227 = ~n78064 & n78146;
  assign n78228 = ~n78226 & ~n78227;
  assign n78229 = ~n78145 & n78228;
  assign n78230 = ~n78225 & n78229;
  assign n78231 = n78224 & n78230;
  assign n78232 = ~n78187 & n78231;
  assign n78233 = n78070 & ~n78232;
  assign n78234 = n78221 & ~n78233;
  assign n78235 = ~n78218 & n78234;
  assign n78236 = ~pi2477 & ~n78235;
  assign n78237 = pi2477 & n78221;
  assign n78238 = ~n78218 & n78237;
  assign n78239 = ~n78233 & n78238;
  assign po2585 = n78236 | n78239;
  assign n78241 = n78064 & n78102;
  assign n78242 = ~n78078 & n78241;
  assign n78243 = ~n78199 & ~n78242;
  assign n78244 = n78078 & n78098;
  assign n78245 = n78084 & n78244;
  assign n78246 = ~n78078 & ~n78090;
  assign n78247 = ~n78223 & ~n78246;
  assign n78248 = ~n78064 & ~n78247;
  assign n78249 = ~n78245 & ~n78248;
  assign n78250 = n78243 & n78249;
  assign n78251 = n78070 & ~n78250;
  assign n78252 = ~n78100 & ~n78148;
  assign n78253 = ~n78078 & n78118;
  assign n78254 = n78252 & ~n78253;
  assign n78255 = n78064 & ~n78254;
  assign n78256 = n78102 & n78141;
  assign n78257 = ~n78129 & ~n78256;
  assign n78258 = ~n78255 & n78257;
  assign n78259 = ~n78110 & ~n78120;
  assign n78260 = ~n78064 & ~n78259;
  assign n78261 = n78258 & ~n78260;
  assign n78262 = ~n78070 & ~n78261;
  assign n78263 = ~n78251 & ~n78262;
  assign n78264 = ~n78078 & n78109;
  assign n78265 = n78078 & ~n78115;
  assign n78266 = ~n78264 & ~n78265;
  assign n78267 = ~n78064 & ~n78266;
  assign n78268 = ~n78100 & n78209;
  assign n78269 = n78185 & ~n78268;
  assign n78270 = ~n78267 & ~n78269;
  assign n78271 = n78263 & n78270;
  assign n78272 = ~pi2495 & ~n78271;
  assign n78273 = pi2495 & n78270;
  assign n78274 = ~n78262 & n78273;
  assign n78275 = ~n78251 & n78274;
  assign po2590 = n78272 | n78275;
  assign n78277 = pi5057 & pi9040;
  assign n78278 = pi5049 & ~pi9040;
  assign n78279 = ~n78277 & ~n78278;
  assign n78280 = pi2423 & n78279;
  assign n78281 = ~pi2423 & ~n78279;
  assign n78282 = ~n78280 & ~n78281;
  assign n78283 = pi5458 & pi9040;
  assign n78284 = pi5106 & ~pi9040;
  assign n78285 = ~n78283 & ~n78284;
  assign n78286 = pi2438 & n78285;
  assign n78287 = ~pi2438 & ~n78285;
  assign n78288 = ~n78286 & ~n78287;
  assign n78289 = pi4974 & pi9040;
  assign n78290 = pi5332 & ~pi9040;
  assign n78291 = ~n78289 & ~n78290;
  assign n78292 = ~pi2433 & n78291;
  assign n78293 = pi2433 & ~n78291;
  assign n78294 = ~n78292 & ~n78293;
  assign n78295 = pi5097 & pi9040;
  assign n78296 = pi5080 & ~pi9040;
  assign n78297 = ~n78295 & ~n78296;
  assign n78298 = ~pi2429 & ~n78297;
  assign n78299 = pi2429 & n78297;
  assign n78300 = ~n78298 & ~n78299;
  assign n78301 = ~n78294 & n78300;
  assign n78302 = ~n78288 & n78301;
  assign n78303 = pi5053 & pi9040;
  assign n78304 = pi5281 & ~pi9040;
  assign n78305 = ~n78303 & ~n78304;
  assign n78306 = ~pi2459 & n78305;
  assign n78307 = pi2459 & ~n78305;
  assign n78308 = ~n78306 & ~n78307;
  assign n78309 = n78302 & n78308;
  assign n78310 = n78294 & ~n78300;
  assign n78311 = ~n78288 & n78310;
  assign n78312 = n78308 & n78311;
  assign n78313 = ~n78309 & ~n78312;
  assign n78314 = n78288 & n78310;
  assign n78315 = ~n78308 & n78314;
  assign n78316 = ~n78288 & ~n78308;
  assign n78317 = ~n78300 & n78316;
  assign n78318 = ~n78294 & n78317;
  assign n78319 = ~n78315 & ~n78318;
  assign n78320 = n78313 & n78319;
  assign n78321 = n78282 & ~n78320;
  assign n78322 = n78294 & n78300;
  assign n78323 = ~n78288 & n78322;
  assign n78324 = ~n78308 & n78323;
  assign n78325 = ~n78294 & ~n78300;
  assign n78326 = ~n78288 & n78325;
  assign n78327 = ~n78324 & ~n78326;
  assign n78328 = n78282 & ~n78327;
  assign n78329 = ~n78282 & n78300;
  assign n78330 = n78308 & n78329;
  assign n78331 = n78288 & ~n78294;
  assign n78332 = ~n78308 & n78310;
  assign n78333 = ~n78331 & ~n78332;
  assign n78334 = ~n78282 & ~n78333;
  assign n78335 = ~n78330 & ~n78334;
  assign n78336 = n78288 & n78322;
  assign n78337 = n78308 & n78336;
  assign n78338 = n78335 & ~n78337;
  assign n78339 = n78300 & ~n78308;
  assign n78340 = n78288 & n78339;
  assign n78341 = ~n78294 & n78340;
  assign n78342 = n78338 & ~n78341;
  assign n78343 = ~n78328 & n78342;
  assign n78344 = pi5101 & pi9040;
  assign n78345 = pi5097 & ~pi9040;
  assign n78346 = ~n78344 & ~n78345;
  assign n78347 = ~pi2458 & ~n78346;
  assign n78348 = pi2458 & n78346;
  assign n78349 = ~n78347 & ~n78348;
  assign n78350 = ~n78343 & ~n78349;
  assign n78351 = ~n78288 & n78300;
  assign n78352 = ~n78282 & ~n78308;
  assign n78353 = n78349 & n78352;
  assign n78354 = n78351 & n78353;
  assign n78355 = ~n78288 & n78308;
  assign n78356 = ~n78300 & n78355;
  assign n78357 = ~n78282 & ~n78356;
  assign n78358 = n78288 & ~n78308;
  assign n78359 = n78294 & n78358;
  assign n78360 = ~n78301 & ~n78351;
  assign n78361 = n78308 & ~n78360;
  assign n78362 = n78282 & ~n78314;
  assign n78363 = ~n78361 & n78362;
  assign n78364 = ~n78359 & n78363;
  assign n78365 = ~n78357 & ~n78364;
  assign n78366 = n78288 & n78325;
  assign n78367 = ~n78308 & n78366;
  assign n78368 = ~n78365 & ~n78367;
  assign n78369 = n78349 & ~n78368;
  assign n78370 = ~n78354 & ~n78369;
  assign n78371 = ~n78350 & n78370;
  assign n78372 = ~n78321 & n78371;
  assign n78373 = ~n78282 & n78337;
  assign n78374 = n78372 & ~n78373;
  assign n78375 = pi2464 & ~n78374;
  assign n78376 = ~pi2464 & ~n78373;
  assign n78377 = n78371 & n78376;
  assign n78378 = ~n78321 & n78377;
  assign po2594 = n78375 | n78378;
  assign n78380 = pi5418 & ~pi9040;
  assign n78381 = pi4989 & pi9040;
  assign n78382 = ~n78380 & ~n78381;
  assign n78383 = ~pi2429 & ~n78382;
  assign n78384 = pi2429 & n78382;
  assign n78385 = ~n78383 & ~n78384;
  assign n78386 = pi5342 & pi9040;
  assign n78387 = pi5102 & ~pi9040;
  assign n78388 = ~n78386 & ~n78387;
  assign n78389 = ~pi2461 & n78388;
  assign n78390 = pi2461 & ~n78388;
  assign n78391 = ~n78389 & ~n78390;
  assign n78392 = pi5458 & ~pi9040;
  assign n78393 = pi5049 & pi9040;
  assign n78394 = ~n78392 & ~n78393;
  assign n78395 = ~pi2438 & ~n78394;
  assign n78396 = pi2438 & n78394;
  assign n78397 = ~n78395 & ~n78396;
  assign n78398 = pi5181 & ~pi9040;
  assign n78399 = pi5281 & pi9040;
  assign n78400 = ~n78398 & ~n78399;
  assign n78401 = ~pi2417 & ~n78400;
  assign n78402 = pi2417 & n78400;
  assign n78403 = ~n78401 & ~n78402;
  assign n78404 = pi5104 & ~pi9040;
  assign n78405 = pi5181 & pi9040;
  assign n78406 = ~n78404 & ~n78405;
  assign n78407 = pi2455 & n78406;
  assign n78408 = ~pi2455 & ~n78406;
  assign n78409 = ~n78407 & ~n78408;
  assign n78410 = ~n78403 & ~n78409;
  assign n78411 = n78397 & n78410;
  assign n78412 = n78391 & n78411;
  assign n78413 = pi5051 & ~pi9040;
  assign n78414 = pi5332 & pi9040;
  assign n78415 = ~n78413 & ~n78414;
  assign n78416 = pi2439 & n78415;
  assign n78417 = ~pi2439 & ~n78415;
  assign n78418 = ~n78416 & ~n78417;
  assign n78419 = ~n78391 & ~n78397;
  assign n78420 = n78418 & n78419;
  assign n78421 = n78403 & ~n78418;
  assign n78422 = ~n78397 & n78421;
  assign n78423 = n78391 & n78422;
  assign n78424 = ~n78420 & ~n78423;
  assign n78425 = ~n78391 & n78397;
  assign n78426 = n78403 & n78425;
  assign n78427 = n78424 & ~n78426;
  assign n78428 = ~n78409 & ~n78427;
  assign n78429 = ~n78391 & ~n78418;
  assign n78430 = ~n78403 & n78409;
  assign n78431 = n78429 & n78430;
  assign n78432 = ~n78418 & n78419;
  assign n78433 = ~n78403 & n78432;
  assign n78434 = ~n78431 & ~n78433;
  assign n78435 = ~n78428 & n78434;
  assign n78436 = ~n78412 & n78435;
  assign n78437 = n78391 & n78397;
  assign n78438 = n78418 & n78437;
  assign n78439 = ~n78403 & n78438;
  assign n78440 = n78418 & n78425;
  assign n78441 = n78403 & n78440;
  assign n78442 = ~n78439 & ~n78441;
  assign n78443 = n78436 & n78442;
  assign n78444 = ~n78385 & ~n78443;
  assign n78445 = ~n78403 & ~n78418;
  assign n78446 = n78397 & n78445;
  assign n78447 = ~n78391 & n78446;
  assign n78448 = ~n78438 & ~n78447;
  assign n78449 = ~n78409 & ~n78448;
  assign n78450 = ~n78391 & n78421;
  assign n78451 = ~n78403 & n78440;
  assign n78452 = ~n78450 & ~n78451;
  assign n78453 = n78409 & ~n78452;
  assign n78454 = n78421 & n78437;
  assign n78455 = ~n78397 & n78445;
  assign n78456 = n78391 & n78455;
  assign n78457 = ~n78454 & ~n78456;
  assign n78458 = ~n78453 & n78457;
  assign n78459 = ~n78449 & n78458;
  assign n78460 = n78385 & ~n78459;
  assign n78461 = ~n78391 & n78418;
  assign n78462 = n78403 & n78461;
  assign n78463 = n78391 & n78418;
  assign n78464 = ~n78403 & n78463;
  assign n78465 = ~n78462 & ~n78464;
  assign n78466 = ~n78409 & ~n78465;
  assign n78467 = n78391 & ~n78397;
  assign n78468 = n78418 & n78467;
  assign n78469 = n78403 & n78468;
  assign n78470 = ~n78454 & ~n78469;
  assign n78471 = ~n78432 & n78470;
  assign n78472 = n78409 & ~n78471;
  assign n78473 = ~n78466 & ~n78472;
  assign n78474 = ~n78397 & ~n78418;
  assign n78475 = n78409 & n78474;
  assign n78476 = ~n78403 & n78475;
  assign n78477 = n78473 & ~n78476;
  assign n78478 = ~n78460 & n78477;
  assign n78479 = ~n78444 & n78478;
  assign n78480 = ~pi2465 & ~n78479;
  assign n78481 = pi2465 & n78479;
  assign po2595 = n78480 | n78481;
  assign n78483 = pi5110 & pi9040;
  assign n78484 = pi5327 & ~pi9040;
  assign n78485 = ~n78483 & ~n78484;
  assign n78486 = ~pi2462 & ~n78485;
  assign n78487 = pi2462 & n78485;
  assign n78488 = ~n78486 & ~n78487;
  assign n78489 = pi5291 & ~pi9040;
  assign n78490 = pi5108 & pi9040;
  assign n78491 = ~n78489 & ~n78490;
  assign n78492 = pi2432 & n78491;
  assign n78493 = ~pi2432 & ~n78491;
  assign n78494 = ~n78492 & ~n78493;
  assign n78495 = pi5208 & pi9040;
  assign n78496 = pi5542 & ~pi9040;
  assign n78497 = ~n78495 & ~n78496;
  assign n78498 = pi2448 & n78497;
  assign n78499 = ~pi2448 & ~n78497;
  assign n78500 = ~n78498 & ~n78499;
  assign n78501 = pi5291 & pi9040;
  assign n78502 = pi4971 & ~pi9040;
  assign n78503 = ~n78501 & ~n78502;
  assign n78504 = pi2453 & n78503;
  assign n78505 = ~pi2453 & ~n78503;
  assign n78506 = ~n78504 & ~n78505;
  assign n78507 = pi5327 & pi9040;
  assign n78508 = pi5103 & ~pi9040;
  assign n78509 = ~n78507 & ~n78508;
  assign n78510 = ~pi2426 & n78509;
  assign n78511 = pi2426 & ~n78509;
  assign n78512 = ~n78510 & ~n78511;
  assign n78513 = ~n78506 & ~n78512;
  assign n78514 = n78500 & n78513;
  assign n78515 = n78494 & n78514;
  assign n78516 = pi5055 & ~pi9040;
  assign n78517 = pi5206 & pi9040;
  assign n78518 = ~n78516 & ~n78517;
  assign n78519 = ~pi2463 & ~n78518;
  assign n78520 = pi2463 & n78518;
  assign n78521 = ~n78519 & ~n78520;
  assign n78522 = n78506 & ~n78512;
  assign n78523 = n78494 & n78522;
  assign n78524 = ~n78500 & n78513;
  assign n78525 = ~n78494 & n78524;
  assign n78526 = ~n78523 & ~n78525;
  assign n78527 = ~n78521 & ~n78526;
  assign n78528 = ~n78515 & ~n78527;
  assign n78529 = ~n78506 & n78512;
  assign n78530 = ~n78500 & n78529;
  assign n78531 = n78521 & n78530;
  assign n78532 = n78513 & n78521;
  assign n78533 = n78494 & n78532;
  assign n78534 = ~n78531 & ~n78533;
  assign n78535 = n78528 & n78534;
  assign n78536 = n78506 & n78512;
  assign n78537 = n78500 & n78536;
  assign n78538 = n78494 & n78537;
  assign n78539 = n78500 & n78529;
  assign n78540 = ~n78494 & n78539;
  assign n78541 = ~n78538 & ~n78540;
  assign n78542 = n78535 & n78541;
  assign n78543 = n78488 & ~n78542;
  assign n78544 = ~n78488 & ~n78521;
  assign n78545 = n78494 & ~n78500;
  assign n78546 = ~n78506 & n78545;
  assign n78547 = ~n78500 & n78512;
  assign n78548 = ~n78546 & ~n78547;
  assign n78549 = n78544 & ~n78548;
  assign n78550 = ~n78494 & n78500;
  assign n78551 = ~n78512 & n78550;
  assign n78552 = ~n78506 & n78551;
  assign n78553 = ~n78494 & n78506;
  assign n78554 = ~n78500 & n78553;
  assign n78555 = ~n78552 & ~n78554;
  assign n78556 = n78494 & n78521;
  assign n78557 = n78500 & n78556;
  assign n78558 = ~n78513 & n78557;
  assign n78559 = n78521 & n78537;
  assign n78560 = ~n78558 & ~n78559;
  assign n78561 = n78555 & n78560;
  assign n78562 = ~n78488 & ~n78561;
  assign n78563 = ~n78500 & n78536;
  assign n78564 = ~n78521 & n78563;
  assign n78565 = ~n78494 & n78564;
  assign n78566 = n78500 & n78522;
  assign n78567 = ~n78494 & n78566;
  assign n78568 = ~n78540 & ~n78567;
  assign n78569 = ~n78521 & ~n78568;
  assign n78570 = ~n78565 & ~n78569;
  assign n78571 = n78521 & n78552;
  assign n78572 = n78570 & ~n78571;
  assign n78573 = ~n78562 & n78572;
  assign n78574 = ~n78549 & n78573;
  assign n78575 = ~n78543 & n78574;
  assign n78576 = ~n78500 & n78522;
  assign n78577 = ~n78494 & n78521;
  assign n78578 = n78576 & n78577;
  assign n78579 = n78575 & ~n78578;
  assign n78580 = ~pi2476 & ~n78579;
  assign n78581 = pi2476 & ~n78578;
  assign n78582 = n78575 & n78581;
  assign po2596 = n78580 | n78582;
  assign n78584 = n78403 & n78432;
  assign n78585 = ~n78456 & ~n78461;
  assign n78586 = n78409 & ~n78585;
  assign n78587 = ~n78584 & ~n78586;
  assign n78588 = ~n78447 & n78587;
  assign n78589 = ~n78409 & n78454;
  assign n78590 = ~n78439 & ~n78589;
  assign n78591 = ~n78469 & n78590;
  assign n78592 = n78588 & n78591;
  assign n78593 = n78385 & ~n78592;
  assign n78594 = ~n78418 & n78425;
  assign n78595 = n78403 & n78594;
  assign n78596 = ~n78423 & ~n78595;
  assign n78597 = ~n78403 & n78468;
  assign n78598 = ~n78433 & ~n78597;
  assign n78599 = ~n78418 & n78437;
  assign n78600 = n78409 & n78599;
  assign n78601 = n78403 & n78438;
  assign n78602 = ~n78600 & ~n78601;
  assign n78603 = n78397 & n78418;
  assign n78604 = ~n78391 & n78403;
  assign n78605 = ~n78603 & ~n78604;
  assign n78606 = ~n78474 & n78605;
  assign n78607 = ~n78409 & ~n78606;
  assign n78608 = n78602 & ~n78607;
  assign n78609 = n78598 & n78608;
  assign n78610 = n78596 & n78609;
  assign n78611 = ~n78385 & ~n78610;
  assign n78612 = ~n78593 & ~n78611;
  assign n78613 = pi2466 & ~n78612;
  assign n78614 = ~pi2466 & ~n78593;
  assign n78615 = ~n78611 & n78614;
  assign po2597 = n78613 | n78615;
  assign n78617 = pi5290 & pi9040;
  assign n78618 = pi5057 & ~pi9040;
  assign n78619 = ~n78617 & ~n78618;
  assign n78620 = ~pi2424 & ~n78619;
  assign n78621 = pi2424 & n78619;
  assign n78622 = ~n78620 & ~n78621;
  assign n78623 = pi5046 & ~pi9040;
  assign n78624 = pi5106 & pi9040;
  assign n78625 = ~n78623 & ~n78624;
  assign n78626 = pi2450 & n78625;
  assign n78627 = ~pi2450 & ~n78625;
  assign n78628 = ~n78626 & ~n78627;
  assign n78629 = pi5094 & pi9040;
  assign n78630 = pi5036 & ~pi9040;
  assign n78631 = ~n78629 & ~n78630;
  assign n78632 = pi2442 & n78631;
  assign n78633 = ~pi2442 & ~n78631;
  assign n78634 = ~n78632 & ~n78633;
  assign n78635 = ~n78628 & ~n78634;
  assign n78636 = pi4979 & ~pi9040;
  assign n78637 = pi5099 & pi9040;
  assign n78638 = ~n78636 & ~n78637;
  assign n78639 = ~pi2462 & n78638;
  assign n78640 = pi2462 & ~n78638;
  assign n78641 = ~n78639 & ~n78640;
  assign n78642 = n78635 & ~n78641;
  assign n78643 = pi5100 & pi9040;
  assign n78644 = pi5099 & ~pi9040;
  assign n78645 = ~n78643 & ~n78644;
  assign n78646 = pi2426 & n78645;
  assign n78647 = ~pi2426 & ~n78645;
  assign n78648 = ~n78646 & ~n78647;
  assign n78649 = pi5342 & ~pi9040;
  assign n78650 = pi5093 & pi9040;
  assign n78651 = ~n78649 & ~n78650;
  assign n78652 = pi2456 & n78651;
  assign n78653 = ~pi2456 & ~n78651;
  assign n78654 = ~n78652 & ~n78653;
  assign n78655 = n78641 & ~n78654;
  assign n78656 = n78648 & n78655;
  assign n78657 = n78628 & n78656;
  assign n78658 = n78641 & n78654;
  assign n78659 = ~n78648 & n78658;
  assign n78660 = n78628 & n78659;
  assign n78661 = ~n78657 & ~n78660;
  assign n78662 = ~n78641 & n78654;
  assign n78663 = ~n78648 & n78662;
  assign n78664 = ~n78628 & ~n78648;
  assign n78665 = ~n78654 & n78664;
  assign n78666 = n78641 & n78665;
  assign n78667 = ~n78663 & ~n78666;
  assign n78668 = n78634 & ~n78667;
  assign n78669 = n78661 & ~n78668;
  assign n78670 = ~n78642 & n78669;
  assign n78671 = n78622 & ~n78670;
  assign n78672 = ~n78641 & ~n78654;
  assign n78673 = ~n78648 & n78672;
  assign n78674 = n78628 & n78673;
  assign n78675 = ~n78634 & n78674;
  assign n78676 = ~n78628 & n78634;
  assign n78677 = n78673 & n78676;
  assign n78678 = ~n78628 & n78648;
  assign n78679 = n78641 & n78678;
  assign n78680 = ~n78677 & ~n78679;
  assign n78681 = n78648 & n78658;
  assign n78682 = ~n78663 & ~n78681;
  assign n78683 = ~n78628 & n78658;
  assign n78684 = n78682 & ~n78683;
  assign n78685 = ~n78634 & ~n78684;
  assign n78686 = n78648 & ~n78654;
  assign n78687 = ~n78641 & n78686;
  assign n78688 = n78628 & n78687;
  assign n78689 = ~n78648 & n78655;
  assign n78690 = n78628 & n78689;
  assign n78691 = ~n78688 & ~n78690;
  assign n78692 = n78648 & n78662;
  assign n78693 = n78634 & n78692;
  assign n78694 = n78691 & ~n78693;
  assign n78695 = ~n78685 & n78694;
  assign n78696 = n78680 & n78695;
  assign n78697 = ~n78622 & ~n78696;
  assign n78698 = ~n78675 & ~n78697;
  assign n78699 = ~n78671 & n78698;
  assign n78700 = n78676 & n78681;
  assign n78701 = n78634 & n78686;
  assign n78702 = n78628 & n78701;
  assign n78703 = ~n78700 & ~n78702;
  assign n78704 = n78634 & n78660;
  assign n78705 = n78703 & ~n78704;
  assign n78706 = n78699 & n78705;
  assign n78707 = ~pi2489 & ~n78706;
  assign n78708 = pi2489 & n78705;
  assign n78709 = n78698 & n78708;
  assign n78710 = ~n78671 & n78709;
  assign po2600 = n78707 | n78710;
  assign n78712 = ~n78403 & n78425;
  assign n78713 = ~n78597 & ~n78712;
  assign n78714 = n78409 & n78713;
  assign n78715 = n78403 & n78463;
  assign n78716 = ~n78419 & ~n78437;
  assign n78717 = n78418 & ~n78716;
  assign n78718 = n78391 & n78445;
  assign n78719 = n78403 & n78419;
  assign n78720 = ~n78718 & ~n78719;
  assign n78721 = ~n78717 & n78720;
  assign n78722 = ~n78409 & n78721;
  assign n78723 = ~n78715 & n78722;
  assign n78724 = ~n78714 & ~n78723;
  assign n78725 = n78403 & n78717;
  assign n78726 = ~n78595 & ~n78725;
  assign n78727 = ~n78724 & n78726;
  assign n78728 = n78385 & ~n78727;
  assign n78729 = n78409 & ~n78716;
  assign n78730 = ~n78403 & n78729;
  assign n78731 = ~n78440 & ~n78467;
  assign n78732 = n78403 & ~n78731;
  assign n78733 = n78409 & n78732;
  assign n78734 = ~n78418 & n78729;
  assign n78735 = ~n78733 & ~n78734;
  assign n78736 = ~n78730 & n78735;
  assign n78737 = ~n78385 & ~n78736;
  assign n78738 = ~n78728 & ~n78737;
  assign n78739 = n78409 & n78423;
  assign n78740 = ~n78409 & ~n78726;
  assign n78741 = ~n78739 & ~n78740;
  assign n78742 = ~n78409 & ~n78713;
  assign n78743 = ~n78423 & ~n78742;
  assign n78744 = ~n78385 & ~n78743;
  assign n78745 = n78741 & ~n78744;
  assign n78746 = n78738 & n78745;
  assign n78747 = pi2468 & ~n78746;
  assign n78748 = ~pi2468 & n78745;
  assign n78749 = ~n78737 & n78748;
  assign n78750 = ~n78728 & n78749;
  assign po2601 = n78747 | n78750;
  assign n78752 = ~n78494 & n78530;
  assign n78753 = n78512 & n78545;
  assign n78754 = n78506 & n78753;
  assign n78755 = ~n78752 & ~n78754;
  assign n78756 = n78521 & ~n78755;
  assign n78757 = ~n78552 & ~n78559;
  assign n78758 = n78494 & n78500;
  assign n78759 = ~n78512 & n78758;
  assign n78760 = n78506 & n78759;
  assign n78761 = ~n78506 & n78550;
  assign n78762 = ~n78554 & ~n78761;
  assign n78763 = ~n78521 & ~n78762;
  assign n78764 = n78494 & ~n78521;
  assign n78765 = n78529 & n78764;
  assign n78766 = ~n78500 & n78765;
  assign n78767 = ~n78500 & n78521;
  assign n78768 = ~n78512 & n78767;
  assign n78769 = ~n78506 & n78768;
  assign n78770 = ~n78766 & ~n78769;
  assign n78771 = ~n78763 & n78770;
  assign n78772 = ~n78760 & n78771;
  assign n78773 = n78757 & n78772;
  assign n78774 = n78488 & ~n78773;
  assign n78775 = ~n78521 & n78552;
  assign n78776 = ~n78494 & n78559;
  assign n78777 = ~n78775 & ~n78776;
  assign n78778 = ~n78774 & n78777;
  assign n78779 = ~n78756 & n78778;
  assign n78780 = n78500 & ~n78506;
  assign n78781 = n78556 & n78780;
  assign n78782 = ~n78531 & ~n78781;
  assign n78783 = n78521 & n78566;
  assign n78784 = ~n78494 & n78576;
  assign n78785 = ~n78783 & ~n78784;
  assign n78786 = n78494 & n78539;
  assign n78787 = ~n78752 & ~n78786;
  assign n78788 = n78494 & n78536;
  assign n78789 = ~n78500 & ~n78512;
  assign n78790 = ~n78788 & ~n78789;
  assign n78791 = ~n78521 & ~n78790;
  assign n78792 = n78787 & ~n78791;
  assign n78793 = n78785 & n78792;
  assign n78794 = n78782 & n78793;
  assign n78795 = ~n78488 & ~n78794;
  assign n78796 = n78779 & ~n78795;
  assign n78797 = ~pi2473 & ~n78796;
  assign n78798 = pi2473 & n78779;
  assign n78799 = ~n78795 & n78798;
  assign po2606 = n78797 | n78799;
  assign n78801 = n78654 & n78678;
  assign n78802 = ~n78663 & ~n78679;
  assign n78803 = ~n78634 & ~n78802;
  assign n78804 = ~n78801 & ~n78803;
  assign n78805 = ~n78648 & ~n78654;
  assign n78806 = ~n78628 & n78805;
  assign n78807 = n78628 & n78655;
  assign n78808 = ~n78806 & ~n78807;
  assign n78809 = n78641 & ~n78648;
  assign n78810 = n78808 & ~n78809;
  assign n78811 = ~n78692 & n78810;
  assign n78812 = n78634 & ~n78811;
  assign n78813 = n78804 & ~n78812;
  assign n78814 = ~n78688 & n78813;
  assign n78815 = n78622 & ~n78814;
  assign n78816 = ~n78628 & n78659;
  assign n78817 = n78691 & ~n78816;
  assign n78818 = n78634 & ~n78817;
  assign n78819 = ~n78815 & ~n78818;
  assign n78820 = ~n78628 & n78692;
  assign n78821 = ~n78641 & ~n78648;
  assign n78822 = ~n78634 & n78821;
  assign n78823 = n78628 & n78822;
  assign n78824 = n78648 & n78676;
  assign n78825 = ~n78654 & n78824;
  assign n78826 = n78628 & n78681;
  assign n78827 = ~n78825 & ~n78826;
  assign n78828 = n78641 & n78648;
  assign n78829 = n78628 & n78828;
  assign n78830 = ~n78673 & ~n78829;
  assign n78831 = ~n78634 & ~n78830;
  assign n78832 = ~n78634 & n78641;
  assign n78833 = ~n78648 & n78832;
  assign n78834 = ~n78628 & n78833;
  assign n78835 = ~n78831 & ~n78834;
  assign n78836 = n78827 & n78835;
  assign n78837 = ~n78622 & ~n78836;
  assign n78838 = ~n78823 & ~n78837;
  assign n78839 = ~n78820 & n78838;
  assign n78840 = n78819 & n78839;
  assign n78841 = ~pi2496 & ~n78840;
  assign n78842 = ~n78815 & ~n78820;
  assign n78843 = ~n78818 & n78842;
  assign n78844 = n78838 & n78843;
  assign n78845 = pi2496 & n78844;
  assign po2607 = n78841 | n78845;
  assign n78847 = ~n78628 & n78656;
  assign n78848 = ~n78659 & ~n78820;
  assign n78849 = n78628 & n78686;
  assign n78850 = ~n78628 & n78673;
  assign n78851 = ~n78849 & ~n78850;
  assign n78852 = n78848 & n78851;
  assign n78853 = ~n78634 & ~n78852;
  assign n78854 = n78628 & n78662;
  assign n78855 = ~n78679 & ~n78854;
  assign n78856 = ~n78689 & n78855;
  assign n78857 = n78634 & ~n78856;
  assign n78858 = n78628 & ~n78648;
  assign n78859 = n78654 & n78858;
  assign n78860 = ~n78641 & n78859;
  assign n78861 = ~n78857 & ~n78860;
  assign n78862 = ~n78853 & n78861;
  assign n78863 = ~n78847 & n78862;
  assign n78864 = ~n78622 & ~n78863;
  assign n78865 = n78628 & ~n78634;
  assign n78866 = n78692 & n78865;
  assign n78867 = ~n78634 & n78689;
  assign n78868 = ~n78634 & n78681;
  assign n78869 = ~n78867 & ~n78868;
  assign n78870 = ~n78628 & ~n78869;
  assign n78871 = ~n78866 & ~n78870;
  assign n78872 = n78628 & n78658;
  assign n78873 = ~n78628 & n78662;
  assign n78874 = ~n78872 & ~n78873;
  assign n78875 = ~n78687 & n78874;
  assign n78876 = ~n78659 & n78875;
  assign n78877 = n78634 & ~n78876;
  assign n78878 = ~n78628 & n78663;
  assign n78879 = ~n78877 & ~n78878;
  assign n78880 = ~n78628 & n78687;
  assign n78881 = ~n78674 & ~n78880;
  assign n78882 = n78879 & n78881;
  assign n78883 = n78871 & n78882;
  assign n78884 = n78622 & ~n78883;
  assign n78885 = ~n78634 & ~n78661;
  assign n78886 = ~n78884 & ~n78885;
  assign n78887 = ~n78690 & ~n78880;
  assign n78888 = n78634 & ~n78887;
  assign n78889 = n78886 & ~n78888;
  assign n78890 = ~n78864 & n78889;
  assign n78891 = pi2502 & ~n78890;
  assign n78892 = ~pi2502 & n78890;
  assign po2609 = n78891 | n78892;
  assign n78894 = n78300 & n78331;
  assign n78895 = n78308 & n78894;
  assign n78896 = ~n78308 & n78351;
  assign n78897 = ~n78336 & ~n78896;
  assign n78898 = n78282 & ~n78897;
  assign n78899 = ~n78895 & ~n78898;
  assign n78900 = ~n78282 & n78308;
  assign n78901 = n78300 & n78900;
  assign n78902 = ~n78294 & n78901;
  assign n78903 = ~n78300 & n78352;
  assign n78904 = ~n78294 & n78903;
  assign n78905 = ~n78902 & ~n78904;
  assign n78906 = ~n78282 & n78288;
  assign n78907 = n78310 & n78906;
  assign n78908 = n78905 & ~n78907;
  assign n78909 = ~n78312 & ~n78324;
  assign n78910 = ~n78300 & n78358;
  assign n78911 = n78909 & ~n78910;
  assign n78912 = n78908 & n78911;
  assign n78913 = n78899 & n78912;
  assign n78914 = ~n78349 & ~n78913;
  assign n78915 = ~n78311 & ~n78336;
  assign n78916 = ~n78308 & ~n78915;
  assign n78917 = ~n78294 & n78308;
  assign n78918 = ~n78288 & n78917;
  assign n78919 = ~n78366 & ~n78918;
  assign n78920 = n78288 & n78300;
  assign n78921 = ~n78308 & n78920;
  assign n78922 = n78919 & ~n78921;
  assign n78923 = n78282 & ~n78922;
  assign n78924 = n78308 & n78322;
  assign n78925 = n78302 & ~n78308;
  assign n78926 = ~n78924 & ~n78925;
  assign n78927 = ~n78282 & ~n78926;
  assign n78928 = n78308 & n78326;
  assign n78929 = ~n78927 & ~n78928;
  assign n78930 = ~n78923 & n78929;
  assign n78931 = ~n78916 & n78930;
  assign n78932 = n78349 & ~n78931;
  assign n78933 = n78282 & n78356;
  assign n78934 = ~n78932 & ~n78933;
  assign n78935 = ~n78282 & n78895;
  assign n78936 = n78934 & ~n78935;
  assign n78937 = ~n78914 & n78936;
  assign n78938 = ~pi2471 & ~n78937;
  assign n78939 = pi2471 & n78934;
  assign n78940 = ~n78914 & n78939;
  assign n78941 = ~n78935 & n78940;
  assign po2610 = n78938 | n78941;
  assign n78943 = pi5096 & pi9040;
  assign n78944 = pi5088 & ~pi9040;
  assign n78945 = ~n78943 & ~n78944;
  assign n78946 = ~pi2434 & ~n78945;
  assign n78947 = pi2434 & n78945;
  assign n78948 = ~n78946 & ~n78947;
  assign n78949 = pi4976 & pi9040;
  assign n78950 = pi5206 & ~pi9040;
  assign n78951 = ~n78949 & ~n78950;
  assign n78952 = pi2447 & n78951;
  assign n78953 = ~pi2447 & ~n78951;
  assign n78954 = ~n78952 & ~n78953;
  assign n78955 = pi5088 & pi9040;
  assign n78956 = pi5108 & ~pi9040;
  assign n78957 = ~n78955 & ~n78956;
  assign n78958 = pi2435 & n78957;
  assign n78959 = ~pi2435 & ~n78957;
  assign n78960 = ~n78958 & ~n78959;
  assign n78961 = n78954 & ~n78960;
  assign n78962 = pi5082 & pi9040;
  assign n78963 = pi5056 & ~pi9040;
  assign n78964 = ~n78962 & ~n78963;
  assign n78965 = ~pi2457 & ~n78964;
  assign n78966 = pi2457 & n78964;
  assign n78967 = ~n78965 & ~n78966;
  assign n78968 = pi5178 & ~pi9040;
  assign n78969 = pi5180 & pi9040;
  assign n78970 = ~n78968 & ~n78969;
  assign n78971 = ~pi2437 & n78970;
  assign n78972 = pi2437 & ~n78970;
  assign n78973 = ~n78971 & ~n78972;
  assign n78974 = n78967 & ~n78973;
  assign n78975 = n78961 & n78974;
  assign n78976 = n78954 & n78960;
  assign n78977 = n78973 & n78976;
  assign n78978 = ~n78954 & ~n78960;
  assign n78979 = n78973 & n78978;
  assign n78980 = ~n78977 & ~n78979;
  assign n78981 = n78967 & ~n78980;
  assign n78982 = ~n78975 & ~n78981;
  assign n78983 = ~n78948 & ~n78982;
  assign n78984 = ~n78967 & n78978;
  assign n78985 = ~n78954 & n78960;
  assign n78986 = ~n78973 & n78985;
  assign n78987 = ~n78984 & ~n78986;
  assign n78988 = pi5042 & ~pi9040;
  assign n78989 = pi5343 & pi9040;
  assign n78990 = ~n78988 & ~n78989;
  assign n78991 = pi2454 & n78990;
  assign n78992 = ~pi2454 & ~n78990;
  assign n78993 = ~n78991 & ~n78992;
  assign n78994 = ~n78948 & n78993;
  assign n78995 = ~n78987 & n78994;
  assign n78996 = ~n78983 & ~n78995;
  assign n78997 = n78967 & n78973;
  assign n78998 = ~n78954 & n78997;
  assign n78999 = ~n78975 & ~n78998;
  assign n79000 = ~n78993 & ~n78999;
  assign n79001 = ~n78967 & n78993;
  assign n79002 = n78954 & n79001;
  assign n79003 = n78961 & n78973;
  assign n79004 = ~n78973 & n78976;
  assign n79005 = ~n79003 & ~n79004;
  assign n79006 = ~n78973 & n78978;
  assign n79007 = n78967 & n79006;
  assign n79008 = n79005 & ~n79007;
  assign n79009 = n78993 & ~n79008;
  assign n79010 = ~n79002 & ~n79009;
  assign n79011 = n78973 & n78985;
  assign n79012 = n78967 & n79011;
  assign n79013 = n79010 & ~n79012;
  assign n79014 = ~n78987 & ~n78993;
  assign n79015 = ~n78967 & n78977;
  assign n79016 = ~n79014 & ~n79015;
  assign n79017 = n79013 & n79016;
  assign n79018 = n78948 & ~n79017;
  assign n79019 = ~n79000 & ~n79018;
  assign n79020 = ~n78948 & ~n78993;
  assign n79021 = n78961 & ~n78967;
  assign n79022 = ~n79011 & ~n79021;
  assign n79023 = n78954 & ~n78973;
  assign n79024 = n79022 & ~n79023;
  assign n79025 = n79020 & ~n79024;
  assign n79026 = n79019 & ~n79025;
  assign n79027 = n78996 & n79026;
  assign n79028 = ~pi2470 & ~n79027;
  assign n79029 = pi2470 & n78996;
  assign n79030 = n79019 & n79029;
  assign n79031 = ~n79025 & n79030;
  assign po2611 = n79028 | n79031;
  assign n79033 = pi5048 & ~pi9040;
  assign n79034 = pi5047 & pi9040;
  assign n79035 = ~n79033 & ~n79034;
  assign n79036 = ~pi2421 & n79035;
  assign n79037 = pi2421 & ~n79035;
  assign n79038 = ~n79036 & ~n79037;
  assign n79039 = pi5096 & ~pi9040;
  assign n79040 = pi5056 & pi9040;
  assign n79041 = ~n79039 & ~n79040;
  assign n79042 = pi2430 & n79041;
  assign n79043 = ~pi2430 & ~n79041;
  assign n79044 = ~n79042 & ~n79043;
  assign n79045 = pi5179 & ~pi9040;
  assign n79046 = pi5103 & pi9040;
  assign n79047 = ~n79045 & ~n79046;
  assign n79048 = pi2435 & n79047;
  assign n79049 = ~pi2435 & ~n79047;
  assign n79050 = ~n79048 & ~n79049;
  assign n79051 = pi5042 & pi9040;
  assign n79052 = pi5047 & ~pi9040;
  assign n79053 = ~n79051 & ~n79052;
  assign n79054 = ~pi2434 & n79053;
  assign n79055 = pi2434 & ~n79053;
  assign n79056 = ~n79054 & ~n79055;
  assign n79057 = pi5179 & pi9040;
  assign n79058 = pi5091 & ~pi9040;
  assign n79059 = ~n79057 & ~n79058;
  assign n79060 = ~pi2448 & n79059;
  assign n79061 = pi2448 & ~n79059;
  assign n79062 = ~n79060 & ~n79061;
  assign n79063 = n79056 & ~n79062;
  assign n79064 = n79050 & n79063;
  assign n79065 = n79044 & n79064;
  assign n79066 = n79038 & n79065;
  assign n79067 = ~n79056 & n79062;
  assign n79068 = n79038 & n79044;
  assign n79069 = n79067 & n79068;
  assign n79070 = ~n79050 & n79069;
  assign n79071 = ~n79066 & ~n79070;
  assign n79072 = ~n79050 & n79063;
  assign n79073 = n79038 & ~n79044;
  assign n79074 = n79072 & n79073;
  assign n79075 = ~n79050 & n79067;
  assign n79076 = n79038 & n79075;
  assign n79077 = ~n79074 & ~n79076;
  assign n79078 = n79050 & ~n79056;
  assign n79079 = ~n79038 & n79078;
  assign n79080 = ~n79038 & n79063;
  assign n79081 = ~n79079 & ~n79080;
  assign n79082 = n79044 & ~n79081;
  assign n79083 = ~n79056 & ~n79062;
  assign n79084 = n79056 & n79062;
  assign n79085 = ~n79083 & ~n79084;
  assign n79086 = n79038 & ~n79050;
  assign n79087 = ~n79044 & ~n79086;
  assign n79088 = ~n79085 & n79087;
  assign n79089 = n79038 & ~n79063;
  assign n79090 = n79044 & n79089;
  assign n79091 = ~n79050 & n79090;
  assign n79092 = ~n79088 & ~n79091;
  assign n79093 = ~n79082 & n79092;
  assign n79094 = n79077 & n79093;
  assign n79095 = pi5339 & pi9040;
  assign n79096 = pi5082 & ~pi9040;
  assign n79097 = ~n79095 & ~n79096;
  assign n79098 = ~pi2453 & ~n79097;
  assign n79099 = pi2453 & n79097;
  assign n79100 = ~n79098 & ~n79099;
  assign n79101 = ~n79094 & n79100;
  assign n79102 = n79071 & ~n79101;
  assign n79103 = n79050 & n79083;
  assign n79104 = ~n79044 & n79103;
  assign n79105 = ~n79038 & n79104;
  assign n79106 = ~n79044 & ~n79100;
  assign n79107 = n79050 & n79067;
  assign n79108 = ~n79080 & ~n79107;
  assign n79109 = ~n79085 & n79086;
  assign n79110 = n79108 & ~n79109;
  assign n79111 = n79106 & ~n79110;
  assign n79112 = ~n79038 & n79075;
  assign n79113 = ~n79038 & ~n79056;
  assign n79114 = ~n79050 & n79113;
  assign n79115 = ~n79038 & n79084;
  assign n79116 = ~n79114 & ~n79115;
  assign n79117 = n79038 & n79063;
  assign n79118 = n79050 & n79084;
  assign n79119 = ~n79117 & ~n79118;
  assign n79120 = n79116 & n79119;
  assign n79121 = n79044 & ~n79120;
  assign n79122 = ~n79112 & ~n79121;
  assign n79123 = ~n79100 & ~n79122;
  assign n79124 = ~n79111 & ~n79123;
  assign n79125 = ~n79105 & n79124;
  assign n79126 = n79102 & n79125;
  assign n79127 = pi2490 & ~n79126;
  assign n79128 = ~pi2490 & n79102;
  assign n79129 = n79125 & n79128;
  assign po2613 = n79127 | n79129;
  assign n79131 = n78403 & n78599;
  assign n79132 = n78409 & n79131;
  assign n79133 = n78445 & ~n78716;
  assign n79134 = ~n78468 & ~n78595;
  assign n79135 = ~n79133 & n79134;
  assign n79136 = ~n78409 & ~n79135;
  assign n79137 = n78403 & n78420;
  assign n79138 = ~n79136 & ~n79137;
  assign n79139 = ~n78418 & n78467;
  assign n79140 = ~n78403 & n78603;
  assign n79141 = ~n79139 & ~n79140;
  assign n79142 = ~n78719 & n79141;
  assign n79143 = n78409 & ~n79142;
  assign n79144 = n79138 & ~n79143;
  assign n79145 = n78385 & ~n79144;
  assign n79146 = ~n79132 & ~n79145;
  assign n79147 = ~n78403 & n78419;
  assign n79148 = ~n78594 & ~n79147;
  assign n79149 = n78409 & ~n79148;
  assign n79150 = ~n78469 & ~n79149;
  assign n79151 = ~n78441 & ~n79131;
  assign n79152 = n78403 & n78474;
  assign n79153 = ~n78603 & ~n79152;
  assign n79154 = ~n79139 & n79153;
  assign n79155 = ~n78409 & ~n79154;
  assign n79156 = ~n78403 & n78420;
  assign n79157 = ~n79155 & ~n79156;
  assign n79158 = n79151 & n79157;
  assign n79159 = n79150 & n79158;
  assign n79160 = ~n78385 & ~n79159;
  assign n79161 = ~n78451 & ~n78715;
  assign n79162 = ~n78409 & ~n79161;
  assign n79163 = ~n79160 & ~n79162;
  assign n79164 = n79146 & n79163;
  assign n79165 = pi2467 & n79164;
  assign n79166 = ~pi2467 & ~n79164;
  assign po2614 = n79165 | n79166;
  assign n79168 = ~n78776 & ~n78781;
  assign n79169 = ~n78494 & n78532;
  assign n79170 = n78506 & n78545;
  assign n79171 = ~n78563 & ~n79170;
  assign n79172 = n78521 & ~n79171;
  assign n79173 = ~n79169 & ~n79172;
  assign n79174 = ~n78521 & n78522;
  assign n79175 = ~n78494 & n79174;
  assign n79176 = ~n78521 & n78530;
  assign n79177 = ~n79175 & ~n79176;
  assign n79178 = n79173 & n79177;
  assign n79179 = n78506 & n78550;
  assign n79180 = ~n78752 & ~n79179;
  assign n79181 = ~n78786 & n79180;
  assign n79182 = n79178 & n79181;
  assign n79183 = ~n78488 & ~n79182;
  assign n79184 = ~n78552 & ~n78563;
  assign n79185 = ~n78788 & n79184;
  assign n79186 = ~n78521 & ~n79185;
  assign n79187 = n78494 & n78524;
  assign n79188 = ~n78760 & ~n79187;
  assign n79189 = ~n78578 & n79188;
  assign n79190 = n78521 & n78539;
  assign n79191 = n79189 & ~n79190;
  assign n79192 = ~n79186 & n79191;
  assign n79193 = n78488 & ~n79192;
  assign n79194 = ~n78752 & n79188;
  assign n79195 = ~n78521 & ~n79194;
  assign n79196 = ~n79193 & ~n79195;
  assign n79197 = ~n79183 & n79196;
  assign n79198 = n79168 & n79197;
  assign n79199 = pi2480 & ~n79198;
  assign n79200 = ~pi2480 & n79198;
  assign po2615 = n79199 | n79200;
  assign n79202 = pi5048 & pi9040;
  assign n79203 = pi5209 & ~pi9040;
  assign n79204 = ~n79202 & ~n79203;
  assign n79205 = ~pi2447 & ~n79204;
  assign n79206 = pi2447 & n79204;
  assign n79207 = ~n79205 & ~n79206;
  assign n79208 = pi5110 & ~pi9040;
  assign n79209 = pi5542 & pi9040;
  assign n79210 = ~n79208 & ~n79209;
  assign n79211 = pi2444 & n79210;
  assign n79212 = ~pi2444 & ~n79210;
  assign n79213 = ~n79211 & ~n79212;
  assign n79214 = pi5178 & pi9040;
  assign n79215 = pi5343 & ~pi9040;
  assign n79216 = ~n79214 & ~n79215;
  assign n79217 = ~pi2433 & ~n79216;
  assign n79218 = pi2433 & n79216;
  assign n79219 = ~n79217 & ~n79218;
  assign n79220 = pi4976 & ~pi9040;
  assign n79221 = pi5109 & pi9040;
  assign n79222 = ~n79220 & ~n79221;
  assign n79223 = ~pi2458 & ~n79222;
  assign n79224 = pi2458 & n79222;
  assign n79225 = ~n79223 & ~n79224;
  assign n79226 = n79219 & ~n79225;
  assign n79227 = pi5447 & ~pi9040;
  assign n79228 = pi4971 & pi9040;
  assign n79229 = ~n79227 & ~n79228;
  assign n79230 = ~pi2437 & n79229;
  assign n79231 = pi2437 & ~n79229;
  assign n79232 = ~n79230 & ~n79231;
  assign n79233 = n79225 & ~n79232;
  assign n79234 = pi5105 & pi9040;
  assign n79235 = pi5180 & ~pi9040;
  assign n79236 = ~n79234 & ~n79235;
  assign n79237 = ~pi2428 & n79236;
  assign n79238 = pi2428 & ~n79236;
  assign n79239 = ~n79237 & ~n79238;
  assign n79240 = ~n79219 & n79239;
  assign n79241 = n79233 & n79240;
  assign n79242 = ~n79226 & ~n79241;
  assign n79243 = ~n79225 & ~n79239;
  assign n79244 = n79242 & ~n79243;
  assign n79245 = n79213 & ~n79244;
  assign n79246 = ~n79213 & ~n79239;
  assign n79247 = n79225 & n79246;
  assign n79248 = n79219 & ~n79239;
  assign n79249 = ~n79232 & n79248;
  assign n79250 = n79225 & n79232;
  assign n79251 = n79219 & n79250;
  assign n79252 = n79239 & n79251;
  assign n79253 = ~n79249 & ~n79252;
  assign n79254 = ~n79219 & ~n79225;
  assign n79255 = ~n79213 & n79239;
  assign n79256 = n79254 & n79255;
  assign n79257 = n79253 & ~n79256;
  assign n79258 = ~n79247 & n79257;
  assign n79259 = ~n79245 & n79258;
  assign n79260 = n79207 & ~n79259;
  assign n79261 = ~n79225 & ~n79232;
  assign n79262 = n79219 & n79261;
  assign n79263 = n79239 & n79262;
  assign n79264 = ~n79225 & n79232;
  assign n79265 = n79219 & n79264;
  assign n79266 = ~n79239 & n79265;
  assign n79267 = ~n79263 & ~n79266;
  assign n79268 = n79213 & ~n79267;
  assign n79269 = ~n79260 & ~n79268;
  assign n79270 = ~n79239 & n79251;
  assign n79271 = n79219 & n79225;
  assign n79272 = ~n79232 & n79271;
  assign n79273 = ~n79219 & n79232;
  assign n79274 = n79225 & n79273;
  assign n79275 = ~n79272 & ~n79274;
  assign n79276 = n79213 & ~n79275;
  assign n79277 = ~n79270 & ~n79276;
  assign n79278 = ~n79219 & n79261;
  assign n79279 = ~n79239 & n79278;
  assign n79280 = n79277 & ~n79279;
  assign n79281 = ~n79207 & ~n79280;
  assign n79282 = ~n79233 & ~n79264;
  assign n79283 = ~n79219 & ~n79282;
  assign n79284 = n79239 & n79264;
  assign n79285 = ~n79283 & ~n79284;
  assign n79286 = ~n79213 & ~n79285;
  assign n79287 = ~n79207 & n79286;
  assign n79288 = ~n79281 & ~n79287;
  assign n79289 = n79269 & n79288;
  assign n79290 = pi2501 & ~n79289;
  assign n79291 = ~pi2501 & n79269;
  assign n79292 = n79288 & n79291;
  assign po2616 = n79290 | n79292;
  assign n79294 = ~n78666 & ~n78880;
  assign n79295 = ~n78860 & n79294;
  assign n79296 = ~n78634 & ~n79295;
  assign n79297 = ~n78674 & ~n78868;
  assign n79298 = ~n78656 & ~n78873;
  assign n79299 = n78634 & ~n79298;
  assign n79300 = ~n78820 & ~n79299;
  assign n79301 = n79297 & n79300;
  assign n79302 = n78622 & ~n79301;
  assign n79303 = ~n78648 & n78654;
  assign n79304 = ~n78809 & ~n79303;
  assign n79305 = n78628 & ~n79304;
  assign n79306 = ~n78683 & ~n78687;
  assign n79307 = n78634 & ~n79306;
  assign n79308 = n78628 & n78654;
  assign n79309 = ~n78663 & ~n79308;
  assign n79310 = ~n78655 & n79309;
  assign n79311 = ~n78634 & ~n79310;
  assign n79312 = ~n79307 & ~n79311;
  assign n79313 = ~n79305 & n79312;
  assign n79314 = ~n78622 & ~n79313;
  assign n79315 = ~n79302 & ~n79314;
  assign n79316 = ~n78677 & ~n78704;
  assign n79317 = n79315 & n79316;
  assign n79318 = ~n79296 & n79317;
  assign n79319 = ~pi2509 & ~n79318;
  assign n79320 = pi2509 & n79316;
  assign n79321 = ~n79296 & n79320;
  assign n79322 = n79315 & n79321;
  assign po2617 = n79319 | n79322;
  assign n79324 = ~n79115 & ~n79117;
  assign n79325 = n79044 & ~n79324;
  assign n79326 = ~n79070 & ~n79325;
  assign n79327 = n79100 & ~n79326;
  assign n79328 = ~n79050 & ~n79056;
  assign n79329 = ~n79083 & ~n79328;
  assign n79330 = n79038 & ~n79329;
  assign n79331 = ~n79064 & ~n79330;
  assign n79332 = ~n79044 & ~n79331;
  assign n79333 = ~n79109 & ~n79332;
  assign n79334 = ~n79038 & n79072;
  assign n79335 = n79038 & n79050;
  assign n79336 = n79062 & n79335;
  assign n79337 = ~n79038 & ~n79329;
  assign n79338 = ~n79336 & ~n79337;
  assign n79339 = n79044 & ~n79338;
  assign n79340 = ~n79334 & ~n79339;
  assign n79341 = n79333 & n79340;
  assign n79342 = ~n79100 & ~n79341;
  assign n79343 = ~n79038 & n79050;
  assign n79344 = ~n79083 & n79343;
  assign n79345 = n79100 & n79344;
  assign n79346 = ~n79038 & ~n79050;
  assign n79347 = n79083 & n79346;
  assign n79348 = n79044 & n79347;
  assign n79349 = ~n79038 & ~n79044;
  assign n79350 = n79050 & n79062;
  assign n79351 = n79349 & n79350;
  assign n79352 = ~n79348 & ~n79351;
  assign n79353 = ~n79345 & n79352;
  assign n79354 = ~n79113 & ~n79118;
  assign n79355 = ~n79044 & n79100;
  assign n79356 = ~n79354 & n79355;
  assign n79357 = n79353 & ~n79356;
  assign n79358 = ~n79342 & n79357;
  assign n79359 = ~n79327 & n79358;
  assign n79360 = pi2492 & ~n79359;
  assign n79361 = ~pi2492 & n79359;
  assign po2618 = n79360 | n79361;
  assign n79363 = n78967 & ~n78993;
  assign n79364 = ~n78977 & ~n78978;
  assign n79365 = n79363 & ~n79364;
  assign n79366 = n78973 & ~n78993;
  assign n79367 = n78978 & n79366;
  assign n79368 = ~n79365 & ~n79367;
  assign n79369 = n78948 & ~n79368;
  assign n79370 = ~n78967 & ~n78973;
  assign n79371 = n78960 & n79370;
  assign n79372 = n78954 & n79371;
  assign n79373 = ~n79023 & ~n79370;
  assign n79374 = n78993 & ~n79373;
  assign n79375 = ~n78967 & n78973;
  assign n79376 = ~n78960 & n79375;
  assign n79377 = n78954 & n79376;
  assign n79378 = ~n79374 & ~n79377;
  assign n79379 = ~n79372 & n79378;
  assign n79380 = n78948 & ~n79379;
  assign n79381 = ~n79369 & ~n79380;
  assign n79382 = ~n78954 & ~n78973;
  assign n79383 = n78967 & n79382;
  assign n79384 = n78960 & n79383;
  assign n79385 = ~n78967 & n79011;
  assign n79386 = ~n79384 & ~n79385;
  assign n79387 = ~n78993 & ~n79386;
  assign n79388 = ~n78961 & ~n79023;
  assign n79389 = n78967 & ~n79388;
  assign n79390 = ~n79011 & ~n79389;
  assign n79391 = ~n78993 & ~n79390;
  assign n79392 = n78960 & ~n78967;
  assign n79393 = n79366 & n79392;
  assign n79394 = ~n78960 & ~n78973;
  assign n79395 = ~n79011 & ~n79394;
  assign n79396 = ~n78967 & ~n79395;
  assign n79397 = n78967 & n78993;
  assign n79398 = n78976 & n79397;
  assign n79399 = n78973 & n79398;
  assign n79400 = ~n79396 & ~n79399;
  assign n79401 = ~n79393 & n79400;
  assign n79402 = ~n79391 & n79401;
  assign n79403 = ~n79384 & n79402;
  assign n79404 = ~n78948 & ~n79403;
  assign n79405 = n78967 & n78979;
  assign n79406 = ~n78967 & n79023;
  assign n79407 = ~n79405 & ~n79406;
  assign n79408 = n78993 & ~n79407;
  assign n79409 = ~n79404 & ~n79408;
  assign n79410 = ~n79387 & n79409;
  assign n79411 = n79381 & n79410;
  assign n79412 = pi2479 & n79411;
  assign n79413 = ~pi2479 & ~n79411;
  assign po2619 = n79412 | n79413;
  assign n79415 = ~n78538 & ~n78546;
  assign n79416 = n78488 & ~n79415;
  assign n79417 = ~n78551 & ~n78761;
  assign n79418 = ~n78514 & n79417;
  assign n79419 = ~n78521 & ~n79418;
  assign n79420 = n78488 & n79419;
  assign n79421 = ~n79416 & ~n79420;
  assign n79422 = n78537 & n78764;
  assign n79423 = ~n78766 & ~n79422;
  assign n79424 = ~n78554 & ~n78789;
  assign n79425 = n78521 & ~n79424;
  assign n79426 = n78488 & n79425;
  assign n79427 = n79423 & ~n79426;
  assign n79428 = n78512 & n78550;
  assign n79429 = n78506 & n79428;
  assign n79430 = ~n78494 & n78529;
  assign n79431 = ~n78754 & ~n79430;
  assign n79432 = n78521 & ~n79431;
  assign n79433 = ~n78552 & ~n78760;
  assign n79434 = ~n78494 & n78536;
  assign n79435 = ~n78576 & ~n79434;
  assign n79436 = ~n78521 & ~n79435;
  assign n79437 = n79433 & ~n79436;
  assign n79438 = ~n79432 & n79437;
  assign n79439 = ~n79429 & n79438;
  assign n79440 = ~n78488 & ~n79439;
  assign n79441 = ~n78786 & n79188;
  assign n79442 = n78521 & ~n79441;
  assign n79443 = ~n79440 & ~n79442;
  assign n79444 = n79427 & n79443;
  assign n79445 = n79421 & n79444;
  assign n79446 = ~pi2497 & ~n79445;
  assign n79447 = pi2497 & n79427;
  assign n79448 = n79421 & n79447;
  assign n79449 = n79443 & n79448;
  assign po2620 = n79446 | n79449;
  assign n79451 = ~n78309 & ~n78315;
  assign n79452 = ~n78282 & ~n79451;
  assign n79453 = ~n78373 & ~n79452;
  assign n79454 = ~n78288 & n78294;
  assign n79455 = n78282 & n79454;
  assign n79456 = ~n78308 & n79455;
  assign n79457 = ~n78308 & n78322;
  assign n79458 = ~n79454 & ~n79457;
  assign n79459 = n78288 & n78308;
  assign n79460 = ~n78294 & n79459;
  assign n79461 = n79458 & ~n79460;
  assign n79462 = n78282 & ~n79461;
  assign n79463 = ~n78318 & ~n79462;
  assign n79464 = ~n78349 & ~n79463;
  assign n79465 = ~n78282 & n78301;
  assign n79466 = ~n78308 & n79465;
  assign n79467 = ~n78907 & ~n79466;
  assign n79468 = ~n78349 & ~n79467;
  assign n79469 = ~n79464 & ~n79468;
  assign n79470 = ~n79456 & n79469;
  assign n79471 = ~n78336 & ~n78356;
  assign n79472 = ~n78366 & n79471;
  assign n79473 = ~n78282 & ~n79472;
  assign n79474 = n78308 & n78314;
  assign n79475 = ~n78894 & ~n79474;
  assign n79476 = n78282 & ~n79475;
  assign n79477 = ~n79473 & ~n79476;
  assign n79478 = ~n78918 & n79477;
  assign n79479 = ~n78324 & ~n78367;
  assign n79480 = n79478 & n79479;
  assign n79481 = n78349 & ~n79480;
  assign n79482 = n79470 & ~n79481;
  assign n79483 = n79453 & n79482;
  assign n79484 = ~pi2478 & ~n79483;
  assign n79485 = pi2478 & n79470;
  assign n79486 = n79453 & n79485;
  assign n79487 = ~n79481 & n79486;
  assign po2621 = n79484 | n79487;
  assign n79489 = n79213 & ~n79239;
  assign n79490 = n79261 & n79489;
  assign n79491 = n79219 & n79490;
  assign n79492 = n79213 & n79239;
  assign n79493 = ~n79232 & n79492;
  assign n79494 = n79225 & n79493;
  assign n79495 = n79219 & n79239;
  assign n79496 = n79232 & n79495;
  assign n79497 = ~n79225 & n79496;
  assign n79498 = n79213 & n79251;
  assign n79499 = ~n79239 & n79498;
  assign n79500 = ~n79497 & ~n79499;
  assign n79501 = ~n79494 & n79500;
  assign n79502 = ~n79491 & n79501;
  assign n79503 = ~n79241 & n79502;
  assign n79504 = ~n79207 & ~n79503;
  assign n79505 = ~n79213 & n79274;
  assign n79506 = ~n79239 & n79505;
  assign n79507 = ~n79225 & n79495;
  assign n79508 = ~n79284 & ~n79507;
  assign n79509 = ~n79213 & ~n79508;
  assign n79510 = ~n79506 & ~n79509;
  assign n79511 = ~n79207 & ~n79510;
  assign n79512 = ~n79239 & n79272;
  assign n79513 = ~n79496 & ~n79512;
  assign n79514 = ~n79279 & n79513;
  assign n79515 = ~n79213 & ~n79514;
  assign n79516 = ~n79511 & ~n79515;
  assign n79517 = ~n79504 & n79516;
  assign n79518 = ~n79219 & ~n79239;
  assign n79519 = n79213 & n79518;
  assign n79520 = n79264 & n79519;
  assign n79521 = ~n79219 & n79492;
  assign n79522 = n79225 & n79521;
  assign n79523 = n79239 & n79274;
  assign n79524 = ~n79213 & n79219;
  assign n79525 = n79225 & n79524;
  assign n79526 = ~n79219 & n79243;
  assign n79527 = ~n79525 & ~n79526;
  assign n79528 = ~n79523 & n79527;
  assign n79529 = ~n79278 & n79528;
  assign n79530 = n79213 & n79261;
  assign n79531 = n79239 & n79530;
  assign n79532 = ~n79239 & n79264;
  assign n79533 = ~n79219 & ~n79232;
  assign n79534 = ~n79532 & ~n79533;
  assign n79535 = n79213 & ~n79534;
  assign n79536 = ~n79531 & ~n79535;
  assign n79537 = n79529 & n79536;
  assign n79538 = n79207 & ~n79537;
  assign n79539 = ~n79522 & ~n79538;
  assign n79540 = ~n79520 & n79539;
  assign n79541 = n79517 & n79540;
  assign n79542 = pi2483 & n79541;
  assign n79543 = ~pi2483 & ~n79541;
  assign po2622 = n79542 | n79543;
  assign n79545 = ~n79239 & n79283;
  assign n79546 = ~n79262 & ~n79273;
  assign n79547 = ~n79213 & ~n79546;
  assign n79548 = ~n79545 & ~n79547;
  assign n79549 = n79232 & n79248;
  assign n79550 = ~n79533 & ~n79549;
  assign n79551 = ~n79265 & n79550;
  assign n79552 = n79213 & ~n79551;
  assign n79553 = n79548 & ~n79552;
  assign n79554 = n79239 & n79272;
  assign n79555 = n79553 & ~n79554;
  assign n79556 = ~n79207 & ~n79555;
  assign n79557 = n79492 & ~n79546;
  assign n79558 = ~n79274 & ~n79278;
  assign n79559 = ~n79265 & ~n79272;
  assign n79560 = n79558 & n79559;
  assign n79561 = ~n79239 & ~n79560;
  assign n79562 = ~n79557 & ~n79561;
  assign n79563 = ~n79252 & n79562;
  assign n79564 = n79207 & ~n79563;
  assign n79565 = ~n79556 & ~n79564;
  assign n79566 = ~n79239 & n79262;
  assign n79567 = ~n79554 & ~n79566;
  assign n79568 = ~n79213 & ~n79567;
  assign n79569 = n79565 & ~n79568;
  assign n79570 = pi2494 & ~n79569;
  assign n79571 = ~pi2494 & ~n79568;
  assign n79572 = ~n79564 & n79571;
  assign n79573 = ~n79556 & n79572;
  assign po2623 = n79570 | n79573;
  assign n79575 = ~n79075 & ~n79103;
  assign n79576 = ~n79062 & n79335;
  assign n79577 = n79575 & ~n79576;
  assign n79578 = n79355 & ~n79577;
  assign n79579 = ~n79038 & n79100;
  assign n79580 = n79118 & n79579;
  assign n79581 = n79044 & n79107;
  assign n79582 = ~n79050 & ~n79062;
  assign n79583 = ~n79080 & ~n79582;
  assign n79584 = n79044 & ~n79583;
  assign n79585 = ~n79581 & ~n79584;
  assign n79586 = n79100 & ~n79585;
  assign n79587 = ~n79580 & ~n79586;
  assign n79588 = n79062 & n79086;
  assign n79589 = n79056 & n79588;
  assign n79590 = ~n79062 & n79346;
  assign n79591 = ~n79589 & ~n79590;
  assign n79592 = n79044 & ~n79591;
  assign n79593 = n79587 & ~n79592;
  assign n79594 = n79063 & n79349;
  assign n79595 = n79050 & n79594;
  assign n79596 = ~n79085 & n79335;
  assign n79597 = ~n79076 & ~n79596;
  assign n79598 = ~n79085 & n79346;
  assign n79599 = ~n79038 & n79107;
  assign n79600 = ~n79598 & ~n79599;
  assign n79601 = ~n79074 & n79600;
  assign n79602 = n79597 & n79601;
  assign n79603 = ~n79595 & n79602;
  assign n79604 = n79050 & n79068;
  assign n79605 = n79056 & n79604;
  assign n79606 = n79603 & ~n79605;
  assign n79607 = ~n79100 & ~n79606;
  assign n79608 = n79593 & ~n79607;
  assign n79609 = ~n79578 & n79608;
  assign n79610 = ~pi2485 & ~n79609;
  assign n79611 = pi2485 & n79593;
  assign n79612 = ~n79578 & n79611;
  assign n79613 = ~n79607 & n79612;
  assign po2624 = n79610 | n79613;
  assign n79615 = ~n79050 & n79083;
  assign n79616 = ~n79064 & ~n79615;
  assign n79617 = n79044 & ~n79616;
  assign n79618 = n79038 & n79084;
  assign n79619 = ~n79103 & ~n79618;
  assign n79620 = ~n79072 & n79619;
  assign n79621 = ~n79044 & ~n79620;
  assign n79622 = ~n79617 & ~n79621;
  assign n79623 = ~n79581 & ~n79589;
  assign n79624 = n79622 & n79623;
  assign n79625 = ~n79100 & ~n79624;
  assign n79626 = ~n79038 & n79064;
  assign n79627 = n79038 & n79067;
  assign n79628 = ~n79115 & ~n79627;
  assign n79629 = ~n79044 & ~n79628;
  assign n79630 = ~n79626 & ~n79629;
  assign n79631 = n79044 & n79050;
  assign n79632 = n79062 & n79631;
  assign n79633 = n79056 & n79632;
  assign n79634 = n79575 & ~n79633;
  assign n79635 = ~n79072 & n79634;
  assign n79636 = n79038 & ~n79635;
  assign n79637 = n79630 & ~n79636;
  assign n79638 = n79100 & ~n79637;
  assign n79639 = ~n79625 & ~n79638;
  assign n79640 = ~n79050 & n79115;
  assign n79641 = ~n79599 & ~n79640;
  assign n79642 = n79044 & ~n79641;
  assign n79643 = n79328 & n79349;
  assign n79644 = ~n79642 & ~n79643;
  assign n79645 = n79639 & n79644;
  assign n79646 = ~pi2503 & ~n79645;
  assign n79647 = n79639 & ~n79642;
  assign n79648 = pi2503 & n79647;
  assign n79649 = ~n79643 & n79648;
  assign po2625 = n79646 | n79649;
  assign n79651 = ~n78367 & ~n78928;
  assign n79652 = n78282 & ~n79651;
  assign n79653 = ~n78349 & n78351;
  assign n79654 = ~n78282 & n79653;
  assign n79655 = n78294 & n79459;
  assign n79656 = ~n78920 & ~n79655;
  assign n79657 = ~n78326 & n79656;
  assign n79658 = n78282 & ~n79657;
  assign n79659 = n78308 & n78323;
  assign n79660 = ~n79658 & ~n79659;
  assign n79661 = ~n78349 & ~n79660;
  assign n79662 = ~n79654 & ~n79661;
  assign n79663 = ~n78312 & ~n78315;
  assign n79664 = n78308 & n78366;
  assign n79665 = ~n78896 & ~n79664;
  assign n79666 = n79663 & n79665;
  assign n79667 = ~n78282 & ~n79666;
  assign n79668 = ~n78288 & ~n78294;
  assign n79669 = ~n78282 & n79668;
  assign n79670 = ~n78308 & n79669;
  assign n79671 = n78308 & n78920;
  assign n79672 = ~n78315 & ~n79671;
  assign n79673 = ~n78925 & n79672;
  assign n79674 = ~n79670 & n79673;
  assign n79675 = n78282 & n78311;
  assign n79676 = n79674 & ~n79675;
  assign n79677 = n78349 & ~n79676;
  assign n79678 = ~n79667 & ~n79677;
  assign n79679 = n79662 & n79678;
  assign n79680 = ~n79652 & n79679;
  assign n79681 = pi2484 & n79680;
  assign n79682 = ~pi2484 & ~n79680;
  assign po2626 = n79681 | n79682;
  assign n79684 = n79239 & n79278;
  assign n79685 = ~n79252 & ~n79684;
  assign n79686 = ~n79213 & ~n79685;
  assign n79687 = n79246 & n79272;
  assign n79688 = ~n79686 & ~n79687;
  assign n79689 = ~n79522 & n79688;
  assign n79690 = n79213 & n79219;
  assign n79691 = n79232 & n79690;
  assign n79692 = ~n79225 & n79691;
  assign n79693 = n79239 & n79692;
  assign n79694 = ~n79239 & n79274;
  assign n79695 = ~n79278 & ~n79694;
  assign n79696 = ~n79265 & n79695;
  assign n79697 = n79207 & ~n79696;
  assign n79698 = ~n79213 & n79697;
  assign n79699 = ~n79239 & n79530;
  assign n79700 = ~n79692 & ~n79699;
  assign n79701 = ~n79249 & n79700;
  assign n79702 = n79232 & n79240;
  assign n79703 = n79233 & ~n79239;
  assign n79704 = ~n79271 & ~n79703;
  assign n79705 = ~n79213 & ~n79704;
  assign n79706 = ~n79702 & ~n79705;
  assign n79707 = n79701 & n79706;
  assign n79708 = ~n79207 & ~n79707;
  assign n79709 = ~n79241 & ~n79520;
  assign n79710 = n79213 & n79262;
  assign n79711 = n79709 & ~n79710;
  assign n79712 = ~n79499 & n79711;
  assign n79713 = n79207 & ~n79712;
  assign n79714 = ~n79708 & ~n79713;
  assign n79715 = ~n79698 & n79714;
  assign n79716 = ~n79693 & n79715;
  assign n79717 = n79689 & n79716;
  assign n79718 = pi2488 & ~n79717;
  assign n79719 = ~pi2488 & n79689;
  assign n79720 = n79716 & n79719;
  assign po2627 = n79718 | n79720;
  assign n79722 = ~n78960 & n78997;
  assign n79723 = ~n78977 & ~n79722;
  assign n79724 = ~n78993 & ~n79723;
  assign n79725 = n78967 & n78985;
  assign n79726 = ~n79376 & ~n79725;
  assign n79727 = n78993 & ~n79726;
  assign n79728 = ~n78967 & n79006;
  assign n79729 = ~n79393 & ~n79728;
  assign n79730 = ~n78975 & n79729;
  assign n79731 = ~n79727 & n79730;
  assign n79732 = ~n79724 & n79731;
  assign n79733 = ~n79372 & ~n79384;
  assign n79734 = n79732 & n79733;
  assign n79735 = n78948 & ~n79734;
  assign n79736 = n78961 & n79370;
  assign n79737 = n78980 & ~n79736;
  assign n79738 = n78993 & ~n79737;
  assign n79739 = ~n78967 & n78986;
  assign n79740 = ~n79738 & ~n79739;
  assign n79741 = n78954 & n78997;
  assign n79742 = n78967 & n78976;
  assign n79743 = ~n79741 & ~n79742;
  assign n79744 = n78993 & ~n79743;
  assign n79745 = n78985 & n78993;
  assign n79746 = ~n78967 & n79745;
  assign n79747 = ~n79744 & ~n79746;
  assign n79748 = n79740 & n79747;
  assign n79749 = ~n78948 & ~n79748;
  assign n79750 = ~n79006 & ~n79012;
  assign n79751 = ~n79377 & n79750;
  assign n79752 = n79020 & ~n79751;
  assign n79753 = ~n79749 & ~n79752;
  assign n79754 = ~n78975 & ~n79372;
  assign n79755 = ~n78993 & ~n79754;
  assign n79756 = n79753 & ~n79755;
  assign n79757 = ~n79735 & n79756;
  assign n79758 = ~pi2486 & n79757;
  assign n79759 = pi2486 & ~n79757;
  assign po2628 = n79758 | n79759;
  assign n79761 = ~n78967 & n78976;
  assign n79762 = ~n79003 & ~n79761;
  assign n79763 = ~n78993 & ~n79762;
  assign n79764 = n78993 & ~n79395;
  assign n79765 = ~n79405 & ~n79764;
  assign n79766 = ~n79763 & n79765;
  assign n79767 = n78948 & ~n79766;
  assign n79768 = n78986 & ~n78993;
  assign n79769 = ~n79767 & ~n79768;
  assign n79770 = ~n79728 & ~n79742;
  assign n79771 = n78993 & ~n79770;
  assign n79772 = n78993 & n79004;
  assign n79773 = n78967 & n78977;
  assign n79774 = n78974 & ~n78993;
  assign n79775 = ~n79375 & ~n79774;
  assign n79776 = ~n78954 & ~n79775;
  assign n79777 = ~n79376 & ~n79776;
  assign n79778 = ~n78975 & n79777;
  assign n79779 = ~n79773 & n79778;
  assign n79780 = ~n79772 & n79779;
  assign n79781 = ~n78948 & ~n79780;
  assign n79782 = ~n79771 & ~n79781;
  assign n79783 = n79769 & n79782;
  assign n79784 = pi2500 & ~n79783;
  assign n79785 = ~pi2500 & n79783;
  assign po2629 = n79784 | n79785;
  assign n79787 = pi5205 & pi9040;
  assign n79788 = pi5294 & ~pi9040;
  assign n79789 = ~n79787 & ~n79788;
  assign n79790 = ~pi2525 & ~n79789;
  assign n79791 = pi2525 & n79789;
  assign n79792 = ~n79790 & ~n79791;
  assign n79793 = pi5289 & pi9040;
  assign n79794 = pi5340 & ~pi9040;
  assign n79795 = ~n79793 & ~n79794;
  assign n79796 = ~pi2521 & n79795;
  assign n79797 = pi2521 & ~n79795;
  assign n79798 = ~n79796 & ~n79797;
  assign n79799 = pi5286 & pi9040;
  assign n79800 = pi5738 & ~pi9040;
  assign n79801 = ~n79799 & ~n79800;
  assign n79802 = ~pi2514 & ~n79801;
  assign n79803 = pi2514 & n79801;
  assign n79804 = ~n79802 & ~n79803;
  assign n79805 = pi5215 & ~pi9040;
  assign n79806 = pi5506 & pi9040;
  assign n79807 = ~n79805 & ~n79806;
  assign n79808 = ~pi2482 & ~n79807;
  assign n79809 = pi2482 & n79807;
  assign n79810 = ~n79808 & ~n79809;
  assign n79811 = pi5430 & ~pi9040;
  assign n79812 = pi5284 & pi9040;
  assign n79813 = ~n79811 & ~n79812;
  assign n79814 = ~pi2524 & n79813;
  assign n79815 = pi2524 & ~n79813;
  assign n79816 = ~n79814 & ~n79815;
  assign n79817 = n79810 & n79816;
  assign n79818 = n79804 & n79817;
  assign n79819 = ~n79798 & n79818;
  assign n79820 = ~n79810 & n79816;
  assign n79821 = n79804 & n79820;
  assign n79822 = n79798 & n79821;
  assign n79823 = ~n79819 & ~n79822;
  assign n79824 = ~n79810 & ~n79816;
  assign n79825 = n79804 & n79824;
  assign n79826 = ~n79798 & n79825;
  assign n79827 = pi5456 & ~pi9040;
  assign n79828 = pi5738 & pi9040;
  assign n79829 = ~n79827 & ~n79828;
  assign n79830 = ~pi2507 & ~n79829;
  assign n79831 = pi2507 & n79829;
  assign n79832 = ~n79830 & ~n79831;
  assign n79833 = n79810 & ~n79816;
  assign n79834 = ~n79798 & n79833;
  assign n79835 = ~n79804 & n79824;
  assign n79836 = n79798 & n79835;
  assign n79837 = ~n79834 & ~n79836;
  assign n79838 = ~n79832 & ~n79837;
  assign n79839 = ~n79826 & ~n79838;
  assign n79840 = ~n79804 & n79820;
  assign n79841 = n79832 & n79840;
  assign n79842 = n79824 & n79832;
  assign n79843 = ~n79798 & n79842;
  assign n79844 = ~n79841 & ~n79843;
  assign n79845 = n79839 & n79844;
  assign n79846 = n79823 & n79845;
  assign n79847 = n79792 & ~n79846;
  assign n79848 = ~n79792 & ~n79832;
  assign n79849 = ~n79798 & ~n79804;
  assign n79850 = ~n79810 & n79849;
  assign n79851 = ~n79804 & n79816;
  assign n79852 = ~n79850 & ~n79851;
  assign n79853 = n79848 & ~n79852;
  assign n79854 = n79798 & n79804;
  assign n79855 = ~n79816 & n79854;
  assign n79856 = ~n79810 & n79855;
  assign n79857 = n79798 & n79810;
  assign n79858 = ~n79804 & n79857;
  assign n79859 = ~n79856 & ~n79858;
  assign n79860 = ~n79798 & n79832;
  assign n79861 = n79804 & n79860;
  assign n79862 = ~n79824 & n79861;
  assign n79863 = n79818 & n79832;
  assign n79864 = ~n79862 & ~n79863;
  assign n79865 = n79859 & n79864;
  assign n79866 = ~n79792 & ~n79865;
  assign n79867 = ~n79804 & n79817;
  assign n79868 = ~n79832 & n79867;
  assign n79869 = n79798 & n79868;
  assign n79870 = n79804 & n79833;
  assign n79871 = n79798 & n79870;
  assign n79872 = ~n79822 & ~n79871;
  assign n79873 = ~n79832 & ~n79872;
  assign n79874 = ~n79869 & ~n79873;
  assign n79875 = n79832 & n79856;
  assign n79876 = n79874 & ~n79875;
  assign n79877 = ~n79866 & n79876;
  assign n79878 = ~n79853 & n79877;
  assign n79879 = ~n79847 & n79878;
  assign n79880 = ~n79804 & n79833;
  assign n79881 = n79798 & n79832;
  assign n79882 = n79880 & n79881;
  assign n79883 = n79879 & ~n79882;
  assign n79884 = ~pi2536 & ~n79883;
  assign n79885 = pi2536 & ~n79882;
  assign n79886 = n79879 & n79885;
  assign po2647 = n79884 | n79886;
  assign n79888 = n79804 & ~n79810;
  assign n79889 = n79860 & n79888;
  assign n79890 = n79798 & n79863;
  assign n79891 = ~n79889 & ~n79890;
  assign n79892 = ~n79856 & ~n79867;
  assign n79893 = ~n79798 & n79817;
  assign n79894 = n79892 & ~n79893;
  assign n79895 = ~n79832 & ~n79894;
  assign n79896 = ~n79798 & n79835;
  assign n79897 = ~n79798 & n79870;
  assign n79898 = ~n79896 & ~n79897;
  assign n79899 = ~n79882 & n79898;
  assign n79900 = n79821 & n79832;
  assign n79901 = n79899 & ~n79900;
  assign n79902 = ~n79895 & n79901;
  assign n79903 = n79792 & ~n79902;
  assign n79904 = n79798 & n79842;
  assign n79905 = n79810 & n79849;
  assign n79906 = ~n79867 & ~n79905;
  assign n79907 = n79832 & ~n79906;
  assign n79908 = ~n79904 & ~n79907;
  assign n79909 = ~n79832 & n79833;
  assign n79910 = n79798 & n79909;
  assign n79911 = ~n79832 & n79840;
  assign n79912 = ~n79910 & ~n79911;
  assign n79913 = n79908 & n79912;
  assign n79914 = ~n79798 & n79821;
  assign n79915 = n79798 & n79840;
  assign n79916 = n79810 & n79854;
  assign n79917 = ~n79915 & ~n79916;
  assign n79918 = ~n79914 & n79917;
  assign n79919 = n79913 & n79918;
  assign n79920 = ~n79792 & ~n79919;
  assign n79921 = n79898 & ~n79915;
  assign n79922 = ~n79832 & ~n79921;
  assign n79923 = ~n79920 & ~n79922;
  assign n79924 = ~n79903 & n79923;
  assign n79925 = n79891 & n79924;
  assign n79926 = pi2538 & ~n79925;
  assign n79927 = ~pi2538 & n79925;
  assign po2651 = n79926 | n79927;
  assign n79929 = pi5545 & ~pi9040;
  assign n79930 = pi5215 & pi9040;
  assign n79931 = ~n79929 & ~n79930;
  assign n79932 = ~pi2517 & ~n79931;
  assign n79933 = pi2517 & n79931;
  assign n79934 = ~n79932 & ~n79933;
  assign n79935 = pi5341 & pi9040;
  assign n79936 = pi5284 & ~pi9040;
  assign n79937 = ~n79935 & ~n79936;
  assign n79938 = ~pi2522 & ~n79937;
  assign n79939 = pi2522 & n79937;
  assign n79940 = ~n79938 & ~n79939;
  assign n79941 = pi5289 & ~pi9040;
  assign n79942 = pi5545 & pi9040;
  assign n79943 = ~n79941 & ~n79942;
  assign n79944 = ~pi2493 & ~n79943;
  assign n79945 = pi2493 & n79943;
  assign n79946 = ~n79944 & ~n79945;
  assign n79947 = pi5456 & pi9040;
  assign n79948 = pi5461 & ~pi9040;
  assign n79949 = ~n79947 & ~n79948;
  assign n79950 = ~pi2469 & n79949;
  assign n79951 = pi2469 & ~n79949;
  assign n79952 = ~n79950 & ~n79951;
  assign n79953 = ~n79946 & ~n79952;
  assign n79954 = pi5630 & ~pi9040;
  assign n79955 = pi5292 & pi9040;
  assign n79956 = ~n79954 & ~n79955;
  assign n79957 = ~pi2506 & n79956;
  assign n79958 = pi2506 & ~n79956;
  assign n79959 = ~n79957 & ~n79958;
  assign n79960 = pi5422 & ~pi9040;
  assign n79961 = pi5630 & pi9040;
  assign n79962 = ~n79960 & ~n79961;
  assign n79963 = pi2527 & n79962;
  assign n79964 = ~pi2527 & ~n79962;
  assign n79965 = ~n79963 & ~n79964;
  assign n79966 = ~n79959 & n79965;
  assign n79967 = n79953 & n79966;
  assign n79968 = n79940 & n79967;
  assign n79969 = n79959 & n79965;
  assign n79970 = n79946 & ~n79952;
  assign n79971 = n79969 & n79970;
  assign n79972 = n79946 & n79952;
  assign n79973 = n79940 & n79972;
  assign n79974 = n79965 & n79973;
  assign n79975 = ~n79959 & n79974;
  assign n79976 = n79940 & n79959;
  assign n79977 = n79952 & n79976;
  assign n79978 = ~n79946 & n79977;
  assign n79979 = ~n79975 & ~n79978;
  assign n79980 = ~n79971 & n79979;
  assign n79981 = ~n79968 & n79980;
  assign n79982 = ~n79940 & n79959;
  assign n79983 = ~n79952 & n79982;
  assign n79984 = n79946 & n79983;
  assign n79985 = n79981 & ~n79984;
  assign n79986 = ~n79934 & ~n79985;
  assign n79987 = n79940 & n79946;
  assign n79988 = ~n79952 & n79987;
  assign n79989 = ~n79959 & n79988;
  assign n79990 = ~n79977 & ~n79989;
  assign n79991 = ~n79940 & n79953;
  assign n79992 = ~n79959 & n79991;
  assign n79993 = n79990 & ~n79992;
  assign n79994 = ~n79965 & ~n79993;
  assign n79995 = ~n79940 & n79952;
  assign n79996 = n79946 & n79995;
  assign n79997 = ~n79965 & n79996;
  assign n79998 = ~n79959 & n79997;
  assign n79999 = ~n79946 & n79976;
  assign n80000 = ~n79946 & n79952;
  assign n80001 = n79959 & n80000;
  assign n80002 = ~n79999 & ~n80001;
  assign n80003 = ~n79965 & ~n80002;
  assign n80004 = ~n79998 & ~n80003;
  assign n80005 = ~n79934 & ~n80004;
  assign n80006 = ~n79994 & ~n80005;
  assign n80007 = ~n79986 & n80006;
  assign n80008 = ~n79940 & ~n79959;
  assign n80009 = n79965 & n80008;
  assign n80010 = n80000 & n80009;
  assign n80011 = ~n79940 & n79946;
  assign n80012 = n79969 & n80011;
  assign n80013 = n79959 & n79996;
  assign n80014 = n79940 & ~n79965;
  assign n80015 = n79946 & n80014;
  assign n80016 = ~n79946 & ~n79959;
  assign n80017 = ~n79940 & n80016;
  assign n80018 = ~n80015 & ~n80017;
  assign n80019 = ~n80013 & n80018;
  assign n80020 = ~n79991 & n80019;
  assign n80021 = n79953 & n79965;
  assign n80022 = n79959 & n80021;
  assign n80023 = ~n79959 & n80000;
  assign n80024 = ~n79940 & ~n79952;
  assign n80025 = ~n80023 & ~n80024;
  assign n80026 = n79965 & ~n80025;
  assign n80027 = ~n80022 & ~n80026;
  assign n80028 = n80020 & n80027;
  assign n80029 = n79934 & ~n80028;
  assign n80030 = ~n80012 & ~n80029;
  assign n80031 = ~n80010 & n80030;
  assign n80032 = n80007 & n80031;
  assign n80033 = pi2540 & n80032;
  assign n80034 = ~pi2540 & ~n80032;
  assign po2653 = n80033 | n80034;
  assign n80036 = n79816 & n79849;
  assign n80037 = n79810 & n80036;
  assign n80038 = ~n79915 & ~n80037;
  assign n80039 = n79832 & ~n80038;
  assign n80040 = ~n79856 & ~n79863;
  assign n80041 = ~n79810 & n79854;
  assign n80042 = ~n79858 & ~n80041;
  assign n80043 = ~n79832 & ~n80042;
  assign n80044 = ~n79798 & ~n79832;
  assign n80045 = n79820 & n80044;
  assign n80046 = ~n79804 & n80045;
  assign n80047 = ~n79804 & n79832;
  assign n80048 = ~n79816 & n80047;
  assign n80049 = ~n79810 & n80048;
  assign n80050 = ~n79897 & ~n80049;
  assign n80051 = ~n80046 & n80050;
  assign n80052 = ~n80043 & n80051;
  assign n80053 = n80040 & n80052;
  assign n80054 = n79792 & ~n80053;
  assign n80055 = ~n79832 & n79856;
  assign n80056 = ~n79890 & ~n80055;
  assign n80057 = ~n80054 & n80056;
  assign n80058 = ~n80039 & n80057;
  assign n80059 = ~n79841 & ~n79889;
  assign n80060 = n79832 & n79870;
  assign n80061 = n79798 & n79880;
  assign n80062 = ~n80060 & ~n80061;
  assign n80063 = ~n79914 & ~n79915;
  assign n80064 = ~n79804 & ~n79816;
  assign n80065 = ~n79893 & ~n80064;
  assign n80066 = ~n79832 & ~n80065;
  assign n80067 = n80063 & ~n80066;
  assign n80068 = n80062 & n80067;
  assign n80069 = n80059 & n80068;
  assign n80070 = ~n79792 & ~n80069;
  assign n80071 = n80058 & ~n80070;
  assign n80072 = ~pi2532 & ~n80071;
  assign n80073 = pi2532 & n80058;
  assign n80074 = ~n80070 & n80073;
  assign po2654 = n80072 | n80074;
  assign n80076 = n79940 & ~n79946;
  assign n80077 = ~n79984 & ~n80076;
  assign n80078 = ~n80016 & n80077;
  assign n80079 = n79965 & ~n80078;
  assign n80080 = ~n79959 & ~n79965;
  assign n80081 = n79946 & n80080;
  assign n80082 = n79940 & ~n79959;
  assign n80083 = ~n79952 & n80082;
  assign n80084 = n79959 & n79973;
  assign n80085 = ~n80083 & ~n80084;
  assign n80086 = ~n79940 & ~n79946;
  assign n80087 = n79959 & ~n79965;
  assign n80088 = n80086 & n80087;
  assign n80089 = n80085 & ~n80088;
  assign n80090 = ~n80081 & n80089;
  assign n80091 = ~n80079 & n80090;
  assign n80092 = n79934 & ~n80091;
  assign n80093 = n79940 & n79953;
  assign n80094 = n79959 & n80093;
  assign n80095 = n79940 & n80000;
  assign n80096 = ~n79959 & n80095;
  assign n80097 = ~n80094 & ~n80096;
  assign n80098 = n79965 & ~n80097;
  assign n80099 = ~n80092 & ~n80098;
  assign n80100 = ~n79959 & n79973;
  assign n80101 = ~n79988 & ~n79996;
  assign n80102 = n79965 & ~n80101;
  assign n80103 = ~n80100 & ~n80102;
  assign n80104 = ~n79992 & n80103;
  assign n80105 = ~n79934 & ~n80104;
  assign n80106 = ~n79970 & ~n80000;
  assign n80107 = ~n79940 & ~n80106;
  assign n80108 = ~n80001 & ~n80107;
  assign n80109 = ~n79965 & ~n80108;
  assign n80110 = ~n79934 & n80109;
  assign n80111 = ~n80105 & ~n80110;
  assign n80112 = n80099 & n80111;
  assign n80113 = pi2553 & ~n80112;
  assign n80114 = ~pi2553 & n80099;
  assign n80115 = n80111 & n80114;
  assign po2656 = n80113 | n80115;
  assign n80117 = pi5347 & ~pi9040;
  assign n80118 = pi5212 & pi9040;
  assign n80119 = ~n80117 & ~n80118;
  assign n80120 = ~pi2513 & ~n80119;
  assign n80121 = pi2513 & n80119;
  assign n80122 = ~n80120 & ~n80121;
  assign n80123 = pi5544 & ~pi9040;
  assign n80124 = pi5430 & pi9040;
  assign n80125 = ~n80123 & ~n80124;
  assign n80126 = pi2515 & n80125;
  assign n80127 = ~pi2515 & ~n80125;
  assign n80128 = ~n80126 & ~n80127;
  assign n80129 = pi5347 & pi9040;
  assign n80130 = pi5338 & ~pi9040;
  assign n80131 = ~n80129 & ~n80130;
  assign n80132 = pi2481 & n80131;
  assign n80133 = ~pi2481 & ~n80131;
  assign n80134 = ~n80132 & ~n80133;
  assign n80135 = n80128 & ~n80134;
  assign n80136 = pi5506 & ~pi9040;
  assign n80137 = pi5214 & pi9040;
  assign n80138 = ~n80136 & ~n80137;
  assign n80139 = ~pi2517 & ~n80138;
  assign n80140 = pi2517 & n80138;
  assign n80141 = ~n80139 & ~n80140;
  assign n80142 = pi5346 & ~pi9040;
  assign n80143 = pi5287 & pi9040;
  assign n80144 = ~n80142 & ~n80143;
  assign n80145 = pi2526 & n80144;
  assign n80146 = ~pi2526 & ~n80144;
  assign n80147 = ~n80145 & ~n80146;
  assign n80148 = ~n80141 & ~n80147;
  assign n80149 = pi5205 & ~pi9040;
  assign n80150 = pi5544 & pi9040;
  assign n80151 = ~n80149 & ~n80150;
  assign n80152 = ~pi2469 & n80151;
  assign n80153 = pi2469 & ~n80151;
  assign n80154 = ~n80152 & ~n80153;
  assign n80155 = n80141 & n80147;
  assign n80156 = n80154 & n80155;
  assign n80157 = ~n80148 & ~n80156;
  assign n80158 = n80135 & ~n80157;
  assign n80159 = ~n80134 & n80154;
  assign n80160 = n80148 & n80159;
  assign n80161 = ~n80158 & ~n80160;
  assign n80162 = n80122 & ~n80161;
  assign n80163 = ~n80154 & n80155;
  assign n80164 = ~n80128 & n80163;
  assign n80165 = n80141 & ~n80154;
  assign n80166 = ~n80128 & ~n80154;
  assign n80167 = ~n80165 & ~n80166;
  assign n80168 = n80134 & ~n80167;
  assign n80169 = ~n80128 & n80154;
  assign n80170 = ~n80147 & n80169;
  assign n80171 = n80141 & n80170;
  assign n80172 = ~n80168 & ~n80171;
  assign n80173 = ~n80164 & n80172;
  assign n80174 = n80122 & ~n80173;
  assign n80175 = ~n80162 & ~n80174;
  assign n80176 = n80128 & ~n80154;
  assign n80177 = n80147 & n80176;
  assign n80178 = ~n80141 & n80177;
  assign n80179 = ~n80141 & n80147;
  assign n80180 = n80154 & n80179;
  assign n80181 = ~n80128 & n80180;
  assign n80182 = ~n80178 & ~n80181;
  assign n80183 = ~n80134 & ~n80182;
  assign n80184 = n80148 & n80154;
  assign n80185 = n80128 & n80184;
  assign n80186 = ~n80128 & n80165;
  assign n80187 = ~n80185 & ~n80186;
  assign n80188 = n80134 & ~n80187;
  assign n80189 = n80141 & ~n80147;
  assign n80190 = ~n80165 & ~n80189;
  assign n80191 = n80128 & ~n80190;
  assign n80192 = ~n80180 & ~n80191;
  assign n80193 = ~n80134 & ~n80192;
  assign n80194 = ~n80128 & n80147;
  assign n80195 = n80159 & n80194;
  assign n80196 = ~n80147 & ~n80154;
  assign n80197 = ~n80180 & ~n80196;
  assign n80198 = ~n80128 & ~n80197;
  assign n80199 = n80128 & n80134;
  assign n80200 = n80155 & n80199;
  assign n80201 = n80154 & n80200;
  assign n80202 = ~n80198 & ~n80201;
  assign n80203 = ~n80195 & n80202;
  assign n80204 = ~n80193 & n80203;
  assign n80205 = ~n80178 & n80204;
  assign n80206 = ~n80122 & ~n80205;
  assign n80207 = ~n80188 & ~n80206;
  assign n80208 = ~n80183 & n80207;
  assign n80209 = n80175 & n80208;
  assign n80210 = pi2552 & n80209;
  assign n80211 = ~pi2552 & ~n80209;
  assign po2658 = n80210 | n80211;
  assign n80213 = n80176 & n80189;
  assign n80214 = n80128 & n80154;
  assign n80215 = ~n80141 & n80214;
  assign n80216 = ~n80213 & ~n80215;
  assign n80217 = ~n80134 & ~n80216;
  assign n80218 = ~n80128 & n80134;
  assign n80219 = n80141 & n80218;
  assign n80220 = n80154 & n80189;
  assign n80221 = ~n80163 & ~n80220;
  assign n80222 = n80148 & ~n80154;
  assign n80223 = n80128 & n80222;
  assign n80224 = n80221 & ~n80223;
  assign n80225 = n80134 & ~n80224;
  assign n80226 = ~n80219 & ~n80225;
  assign n80227 = n80128 & n80180;
  assign n80228 = n80226 & ~n80227;
  assign n80229 = ~n80128 & n80148;
  assign n80230 = ~n80154 & n80179;
  assign n80231 = ~n80229 & ~n80230;
  assign n80232 = ~n80134 & ~n80231;
  assign n80233 = ~n80128 & n80156;
  assign n80234 = ~n80232 & ~n80233;
  assign n80235 = n80228 & n80234;
  assign n80236 = n80122 & ~n80235;
  assign n80237 = ~n80217 & ~n80236;
  assign n80238 = ~n80156 & ~n80184;
  assign n80239 = n80128 & ~n80238;
  assign n80240 = ~n80213 & ~n80239;
  assign n80241 = ~n80122 & ~n80240;
  assign n80242 = ~n80122 & n80134;
  assign n80243 = ~n80231 & n80242;
  assign n80244 = ~n80241 & ~n80243;
  assign n80245 = ~n80122 & ~n80134;
  assign n80246 = ~n80128 & n80189;
  assign n80247 = ~n80180 & ~n80246;
  assign n80248 = ~n80165 & n80247;
  assign n80249 = n80245 & ~n80248;
  assign n80250 = n80244 & ~n80249;
  assign n80251 = n80237 & n80250;
  assign n80252 = ~pi2546 & ~n80251;
  assign n80253 = pi2546 & n80244;
  assign n80254 = n80237 & n80253;
  assign n80255 = ~n80249 & n80254;
  assign po2659 = n80252 | n80255;
  assign n80257 = pi5298 & pi9040;
  assign n80258 = pi5288 & ~pi9040;
  assign n80259 = ~n80257 & ~n80258;
  assign n80260 = ~pi2516 & n80259;
  assign n80261 = pi2516 & ~n80259;
  assign n80262 = ~n80260 & ~n80261;
  assign n80263 = pi5213 & pi9040;
  assign n80264 = pi5330 & ~pi9040;
  assign n80265 = ~n80263 & ~n80264;
  assign n80266 = ~pi2504 & ~n80265;
  assign n80267 = pi2504 & n80265;
  assign n80268 = ~n80266 & ~n80267;
  assign n80269 = pi5213 & ~pi9040;
  assign n80270 = pi5583 & pi9040;
  assign n80271 = ~n80269 & ~n80270;
  assign n80272 = pi2518 & n80271;
  assign n80273 = ~pi2518 & ~n80271;
  assign n80274 = ~n80272 & ~n80273;
  assign n80275 = pi5296 & ~pi9040;
  assign n80276 = pi5297 & pi9040;
  assign n80277 = ~n80275 & ~n80276;
  assign n80278 = ~pi2472 & ~n80277;
  assign n80279 = pi2472 & n80277;
  assign n80280 = ~n80278 & ~n80279;
  assign n80281 = n80274 & ~n80280;
  assign n80282 = ~n80268 & n80281;
  assign n80283 = pi5283 & pi9040;
  assign n80284 = pi5298 & ~pi9040;
  assign n80285 = ~n80283 & ~n80284;
  assign n80286 = ~pi2520 & ~n80285;
  assign n80287 = pi2520 & n80285;
  assign n80288 = ~n80286 & ~n80287;
  assign n80289 = n80268 & ~n80288;
  assign n80290 = ~n80274 & ~n80280;
  assign n80291 = n80289 & n80290;
  assign n80292 = pi5378 & ~pi9040;
  assign n80293 = pi5736 & pi9040;
  assign n80294 = ~n80292 & ~n80293;
  assign n80295 = ~pi2487 & ~n80294;
  assign n80296 = pi2487 & n80294;
  assign n80297 = ~n80295 & ~n80296;
  assign n80298 = ~n80268 & n80297;
  assign n80299 = n80280 & n80298;
  assign n80300 = n80268 & ~n80280;
  assign n80301 = n80297 & n80300;
  assign n80302 = ~n80299 & ~n80301;
  assign n80303 = ~n80274 & ~n80302;
  assign n80304 = ~n80291 & ~n80303;
  assign n80305 = n80289 & n80297;
  assign n80306 = ~n80280 & n80305;
  assign n80307 = n80268 & ~n80297;
  assign n80308 = n80288 & n80307;
  assign n80309 = n80280 & n80308;
  assign n80310 = ~n80306 & ~n80309;
  assign n80311 = n80274 & n80280;
  assign n80312 = n80307 & n80311;
  assign n80313 = n80274 & ~n80297;
  assign n80314 = n80288 & n80313;
  assign n80315 = ~n80268 & n80314;
  assign n80316 = ~n80312 & ~n80315;
  assign n80317 = n80310 & n80316;
  assign n80318 = n80304 & n80317;
  assign n80319 = ~n80282 & n80318;
  assign n80320 = n80262 & ~n80319;
  assign n80321 = n80268 & n80288;
  assign n80322 = n80297 & n80321;
  assign n80323 = ~n80299 & ~n80322;
  assign n80324 = n80289 & ~n80297;
  assign n80325 = ~n80280 & n80324;
  assign n80326 = n80323 & ~n80325;
  assign n80327 = n80274 & ~n80326;
  assign n80328 = ~n80280 & n80308;
  assign n80329 = ~n80268 & n80288;
  assign n80330 = n80297 & n80329;
  assign n80331 = ~n80280 & n80330;
  assign n80332 = ~n80268 & ~n80297;
  assign n80333 = ~n80289 & ~n80332;
  assign n80334 = n80280 & ~n80333;
  assign n80335 = ~n80331 & ~n80334;
  assign n80336 = ~n80328 & n80335;
  assign n80337 = ~n80274 & ~n80336;
  assign n80338 = ~n80327 & ~n80337;
  assign n80339 = ~n80262 & ~n80338;
  assign n80340 = ~n80268 & ~n80288;
  assign n80341 = ~n80297 & n80340;
  assign n80342 = ~n80274 & n80341;
  assign n80343 = ~n80280 & n80342;
  assign n80344 = ~n80274 & n80306;
  assign n80345 = ~n80343 & ~n80344;
  assign n80346 = ~n80280 & ~n80297;
  assign n80347 = n80288 & n80346;
  assign n80348 = ~n80268 & n80347;
  assign n80349 = n80274 & n80348;
  assign n80350 = n80345 & ~n80349;
  assign n80351 = ~n80280 & n80297;
  assign n80352 = ~n80288 & n80351;
  assign n80353 = ~n80268 & n80352;
  assign n80354 = n80280 & n80321;
  assign n80355 = ~n80353 & ~n80354;
  assign n80356 = n80274 & ~n80355;
  assign n80357 = n80350 & ~n80356;
  assign n80358 = ~n80339 & n80357;
  assign n80359 = ~n80320 & n80358;
  assign n80360 = ~pi2544 & n80359;
  assign n80361 = pi2544 & ~n80359;
  assign po2660 = n80360 | n80361;
  assign n80363 = ~pi5204 & ~pi9040;
  assign n80364 = pi5546 & pi9040;
  assign n80365 = ~n80363 & ~n80364;
  assign n80366 = ~pi2504 & n80365;
  assign n80367 = pi2504 & ~n80365;
  assign n80368 = ~n80366 & ~n80367;
  assign n80369 = pi5337 & ~pi9040;
  assign n80370 = pi5335 & pi9040;
  assign n80371 = ~n80369 & ~n80370;
  assign n80372 = ~pi2523 & ~n80371;
  assign n80373 = pi2523 & n80371;
  assign n80374 = ~n80372 & ~n80373;
  assign n80375 = pi5584 & ~pi9040;
  assign n80376 = pi5203 & pi9040;
  assign n80377 = ~n80375 & ~n80376;
  assign n80378 = ~pi2524 & ~n80377;
  assign n80379 = pi2524 & n80377;
  assign n80380 = ~n80378 & ~n80379;
  assign n80381 = pi5429 & ~pi9040;
  assign n80382 = pi5543 & pi9040;
  assign n80383 = ~n80381 & ~n80382;
  assign n80384 = pi2525 & n80383;
  assign n80385 = ~pi2525 & ~n80383;
  assign n80386 = ~n80384 & ~n80385;
  assign n80387 = pi5344 & pi9040;
  assign n80388 = pi5736 & ~pi9040;
  assign n80389 = ~n80387 & ~n80388;
  assign n80390 = ~pi2487 & ~n80389;
  assign n80391 = pi2487 & n80389;
  assign n80392 = ~n80390 & ~n80391;
  assign n80393 = ~n80386 & ~n80392;
  assign n80394 = n80380 & n80393;
  assign n80395 = ~n80374 & n80394;
  assign n80396 = pi5345 & ~pi9040;
  assign n80397 = pi5584 & pi9040;
  assign n80398 = ~n80396 & ~n80397;
  assign n80399 = ~pi2510 & n80398;
  assign n80400 = pi2510 & ~n80398;
  assign n80401 = ~n80399 & ~n80400;
  assign n80402 = ~n80386 & n80392;
  assign n80403 = ~n80380 & n80402;
  assign n80404 = ~n80374 & n80380;
  assign n80405 = n80392 & n80404;
  assign n80406 = n80386 & n80405;
  assign n80407 = ~n80403 & ~n80406;
  assign n80408 = n80380 & ~n80392;
  assign n80409 = n80374 & n80408;
  assign n80410 = n80386 & ~n80392;
  assign n80411 = ~n80380 & n80410;
  assign n80412 = ~n80374 & n80411;
  assign n80413 = ~n80409 & ~n80412;
  assign n80414 = n80407 & n80413;
  assign n80415 = n80401 & ~n80414;
  assign n80416 = ~n80380 & n80393;
  assign n80417 = n80386 & n80392;
  assign n80418 = n80374 & n80417;
  assign n80419 = ~n80386 & n80404;
  assign n80420 = ~n80418 & ~n80419;
  assign n80421 = ~n80416 & n80420;
  assign n80422 = ~n80401 & ~n80421;
  assign n80423 = n80374 & ~n80380;
  assign n80424 = n80392 & n80423;
  assign n80425 = n80386 & n80424;
  assign n80426 = ~n80422 & ~n80425;
  assign n80427 = ~n80415 & n80426;
  assign n80428 = ~n80395 & n80427;
  assign n80429 = ~n80368 & ~n80428;
  assign n80430 = n80380 & n80417;
  assign n80431 = n80374 & n80401;
  assign n80432 = n80430 & n80431;
  assign n80433 = n80401 & n80416;
  assign n80434 = n80380 & n80402;
  assign n80435 = n80401 & n80434;
  assign n80436 = ~n80433 & ~n80435;
  assign n80437 = ~n80374 & ~n80436;
  assign n80438 = ~n80432 & ~n80437;
  assign n80439 = n80374 & n80402;
  assign n80440 = ~n80374 & n80417;
  assign n80441 = ~n80439 & ~n80440;
  assign n80442 = n80386 & n80408;
  assign n80443 = n80441 & ~n80442;
  assign n80444 = ~n80403 & n80443;
  assign n80445 = ~n80401 & ~n80444;
  assign n80446 = ~n80380 & n80417;
  assign n80447 = ~n80374 & n80446;
  assign n80448 = ~n80445 & ~n80447;
  assign n80449 = ~n80374 & n80442;
  assign n80450 = n80374 & n80411;
  assign n80451 = ~n80449 & ~n80450;
  assign n80452 = n80448 & n80451;
  assign n80453 = n80438 & n80452;
  assign n80454 = n80368 & ~n80453;
  assign n80455 = n80374 & n80394;
  assign n80456 = n80402 & n80423;
  assign n80457 = ~n80455 & ~n80456;
  assign n80458 = n80401 & ~n80457;
  assign n80459 = ~n80454 & ~n80458;
  assign n80460 = n80374 & n80416;
  assign n80461 = ~n80449 & ~n80460;
  assign n80462 = ~n80401 & ~n80461;
  assign n80463 = n80459 & ~n80462;
  assign n80464 = ~n80429 & n80463;
  assign n80465 = pi2547 & ~n80464;
  assign n80466 = ~pi2547 & n80464;
  assign po2662 = n80465 | n80466;
  assign n80468 = ~n79819 & ~n79850;
  assign n80469 = n79792 & ~n80468;
  assign n80470 = ~n79855 & ~n80041;
  assign n80471 = ~n79825 & n80470;
  assign n80472 = ~n79832 & ~n80471;
  assign n80473 = n79792 & n80472;
  assign n80474 = ~n80469 & ~n80473;
  assign n80475 = n79818 & n80044;
  assign n80476 = ~n80046 & ~n80475;
  assign n80477 = ~n79858 & ~n80064;
  assign n80478 = n79832 & ~n80477;
  assign n80479 = n79792 & n80478;
  assign n80480 = n80476 & ~n80479;
  assign n80481 = n79816 & n79854;
  assign n80482 = n79810 & n80481;
  assign n80483 = n79798 & n79820;
  assign n80484 = ~n80037 & ~n80483;
  assign n80485 = n79832 & ~n80484;
  assign n80486 = ~n79856 & ~n79897;
  assign n80487 = n79798 & n79817;
  assign n80488 = ~n79880 & ~n80487;
  assign n80489 = ~n79832 & ~n80488;
  assign n80490 = n80486 & ~n80489;
  assign n80491 = ~n80485 & n80490;
  assign n80492 = ~n80482 & n80491;
  assign n80493 = ~n79792 & ~n80492;
  assign n80494 = n79898 & ~n79914;
  assign n80495 = n79832 & ~n80494;
  assign n80496 = ~n80493 & ~n80495;
  assign n80497 = n80480 & n80496;
  assign n80498 = n80474 & n80497;
  assign n80499 = ~pi2542 & ~n80498;
  assign n80500 = pi2542 & n80480;
  assign n80501 = n80474 & n80500;
  assign n80502 = n80496 & n80501;
  assign po2663 = n80499 | n80502;
  assign n80504 = ~n80374 & n80401;
  assign n80505 = n80386 & n80504;
  assign n80506 = ~n80374 & ~n80380;
  assign n80507 = ~n80392 & n80506;
  assign n80508 = ~n80386 & n80507;
  assign n80509 = ~n80446 & ~n80508;
  assign n80510 = ~n80401 & ~n80509;
  assign n80511 = n80457 & ~n80510;
  assign n80512 = ~n80505 & n80511;
  assign n80513 = n80368 & ~n80512;
  assign n80514 = n80401 & n80450;
  assign n80515 = ~n80374 & ~n80401;
  assign n80516 = n80411 & n80515;
  assign n80517 = ~n80419 & ~n80516;
  assign n80518 = ~n80434 & ~n80446;
  assign n80519 = ~n80374 & n80402;
  assign n80520 = n80518 & ~n80519;
  assign n80521 = n80401 & ~n80520;
  assign n80522 = n80374 & n80442;
  assign n80523 = ~n80460 & ~n80522;
  assign n80524 = ~n80401 & n80430;
  assign n80525 = n80523 & ~n80524;
  assign n80526 = ~n80521 & n80525;
  assign n80527 = n80517 & n80526;
  assign n80528 = ~n80368 & ~n80527;
  assign n80529 = ~n80514 & ~n80528;
  assign n80530 = ~n80513 & n80529;
  assign n80531 = n80434 & n80515;
  assign n80532 = ~n80401 & n80408;
  assign n80533 = n80374 & n80532;
  assign n80534 = ~n80531 & ~n80533;
  assign n80535 = ~n80401 & n80456;
  assign n80536 = n80534 & ~n80535;
  assign n80537 = n80530 & n80536;
  assign n80538 = ~pi2541 & ~n80537;
  assign n80539 = pi2541 & n80536;
  assign n80540 = n80529 & n80539;
  assign n80541 = ~n80513 & n80540;
  assign po2664 = n80538 | n80541;
  assign n80543 = ~n79959 & n80107;
  assign n80544 = ~n79995 & ~n80093;
  assign n80545 = ~n79965 & ~n80544;
  assign n80546 = ~n80543 & ~n80545;
  assign n80547 = n79952 & n80082;
  assign n80548 = ~n80024 & ~n80547;
  assign n80549 = ~n80095 & n80548;
  assign n80550 = n79965 & ~n80549;
  assign n80551 = n80546 & ~n80550;
  assign n80552 = n79959 & n79988;
  assign n80553 = n80551 & ~n80552;
  assign n80554 = ~n79934 & ~n80553;
  assign n80555 = n79969 & ~n80544;
  assign n80556 = ~n79991 & ~n79996;
  assign n80557 = ~n79988 & ~n80095;
  assign n80558 = n80556 & n80557;
  assign n80559 = ~n79959 & ~n80558;
  assign n80560 = ~n80555 & ~n80559;
  assign n80561 = ~n80084 & n80560;
  assign n80562 = n79934 & ~n80561;
  assign n80563 = ~n80554 & ~n80562;
  assign n80564 = ~n79959 & n80093;
  assign n80565 = ~n80552 & ~n80564;
  assign n80566 = ~n79965 & ~n80565;
  assign n80567 = n80563 & ~n80566;
  assign n80568 = pi2549 & ~n80567;
  assign n80569 = ~pi2549 & ~n80566;
  assign n80570 = ~n80562 & n80569;
  assign n80571 = ~n80554 & n80570;
  assign po2665 = n80568 | n80571;
  assign n80573 = pi5296 & pi9040;
  assign n80574 = pi5628 & ~pi9040;
  assign n80575 = ~n80573 & ~n80574;
  assign n80576 = ~pi2512 & n80575;
  assign n80577 = pi2512 & ~n80575;
  assign n80578 = ~n80576 & ~n80577;
  assign n80579 = pi5344 & ~pi9040;
  assign n80580 = pi5641 & pi9040;
  assign n80581 = ~n80579 & ~n80580;
  assign n80582 = ~pi2508 & n80581;
  assign n80583 = pi2508 & ~n80581;
  assign n80584 = ~n80582 & ~n80583;
  assign n80585 = pi5583 & ~pi9040;
  assign n80586 = pi5204 & pi9040;
  assign n80587 = ~n80585 & ~n80586;
  assign n80588 = ~pi2522 & n80587;
  assign n80589 = pi2522 & ~n80587;
  assign n80590 = ~n80588 & ~n80589;
  assign n80591 = pi5288 & pi9040;
  assign n80592 = pi5335 & ~pi9040;
  assign n80593 = ~n80591 & ~n80592;
  assign n80594 = ~pi2499 & n80593;
  assign n80595 = pi2499 & ~n80593;
  assign n80596 = ~n80594 & ~n80595;
  assign n80597 = ~n80590 & ~n80596;
  assign n80598 = n80584 & n80597;
  assign n80599 = pi5345 & pi9040;
  assign n80600 = pi5336 & ~pi9040;
  assign n80601 = ~n80599 & ~n80600;
  assign n80602 = pi2519 & n80601;
  assign n80603 = ~pi2519 & ~n80601;
  assign n80604 = ~n80602 & ~n80603;
  assign n80605 = n80598 & ~n80604;
  assign n80606 = n80584 & ~n80604;
  assign n80607 = n80596 & n80606;
  assign n80608 = n80590 & n80607;
  assign n80609 = ~n80605 & ~n80608;
  assign n80610 = n80590 & n80596;
  assign n80611 = ~n80584 & n80604;
  assign n80612 = n80610 & n80611;
  assign n80613 = ~n80590 & n80596;
  assign n80614 = n80584 & n80613;
  assign n80615 = n80604 & n80614;
  assign n80616 = ~n80612 & ~n80615;
  assign n80617 = n80609 & n80616;
  assign n80618 = ~n80578 & ~n80617;
  assign n80619 = n80590 & ~n80596;
  assign n80620 = n80584 & n80619;
  assign n80621 = n80604 & n80620;
  assign n80622 = ~n80614 & ~n80621;
  assign n80623 = ~n80578 & ~n80622;
  assign n80624 = ~n80584 & n80619;
  assign n80625 = ~n80604 & n80624;
  assign n80626 = n80578 & ~n80596;
  assign n80627 = ~n80604 & n80626;
  assign n80628 = ~n80584 & ~n80590;
  assign n80629 = n80604 & n80610;
  assign n80630 = ~n80628 & ~n80629;
  assign n80631 = n80578 & ~n80630;
  assign n80632 = ~n80627 & ~n80631;
  assign n80633 = ~n80625 & n80632;
  assign n80634 = ~n80596 & n80628;
  assign n80635 = n80604 & n80634;
  assign n80636 = n80633 & ~n80635;
  assign n80637 = ~n80623 & n80636;
  assign n80638 = pi5334 & pi9040;
  assign n80639 = pi5641 & ~pi9040;
  assign n80640 = ~n80638 & ~n80639;
  assign n80641 = ~pi2493 & ~n80640;
  assign n80642 = pi2493 & n80640;
  assign n80643 = ~n80641 & ~n80642;
  assign n80644 = ~n80637 & ~n80643;
  assign n80645 = n80584 & ~n80596;
  assign n80646 = n80578 & n80604;
  assign n80647 = n80643 & n80646;
  assign n80648 = n80645 & n80647;
  assign n80649 = n80578 & ~n80607;
  assign n80650 = n80590 & n80611;
  assign n80651 = ~n80597 & ~n80645;
  assign n80652 = ~n80604 & ~n80651;
  assign n80653 = ~n80584 & n80610;
  assign n80654 = ~n80578 & ~n80653;
  assign n80655 = ~n80652 & n80654;
  assign n80656 = ~n80650 & n80655;
  assign n80657 = ~n80649 & ~n80656;
  assign n80658 = n80596 & n80611;
  assign n80659 = ~n80590 & n80658;
  assign n80660 = ~n80657 & ~n80659;
  assign n80661 = n80643 & ~n80660;
  assign n80662 = ~n80648 & ~n80661;
  assign n80663 = ~n80644 & n80662;
  assign n80664 = ~n80618 & n80663;
  assign n80665 = n80578 & n80625;
  assign n80666 = n80664 & ~n80665;
  assign n80667 = pi2535 & ~n80666;
  assign n80668 = ~pi2535 & ~n80665;
  assign n80669 = n80663 & n80668;
  assign n80670 = ~n80618 & n80669;
  assign po2667 = n80667 | n80670;
  assign n80672 = n80262 & ~n80274;
  assign n80673 = ~n80280 & n80298;
  assign n80674 = n80280 & n80305;
  assign n80675 = ~n80280 & n80321;
  assign n80676 = ~n80674 & ~n80675;
  assign n80677 = ~n80673 & n80676;
  assign n80678 = n80672 & ~n80677;
  assign n80679 = ~n80288 & n80346;
  assign n80680 = n80297 & n80340;
  assign n80681 = n80280 & n80680;
  assign n80682 = ~n80679 & ~n80681;
  assign n80683 = ~n80322 & ~n80324;
  assign n80684 = n80682 & n80683;
  assign n80685 = n80274 & ~n80684;
  assign n80686 = ~n80297 & n80329;
  assign n80687 = n80280 & n80686;
  assign n80688 = ~n80685 & ~n80687;
  assign n80689 = n80262 & ~n80688;
  assign n80690 = ~n80678 & ~n80689;
  assign n80691 = ~n80321 & ~n80340;
  assign n80692 = n80280 & ~n80691;
  assign n80693 = ~n80341 & ~n80692;
  assign n80694 = ~n80274 & ~n80693;
  assign n80695 = ~n80330 & ~n80673;
  assign n80696 = ~n80674 & n80695;
  assign n80697 = n80274 & ~n80696;
  assign n80698 = ~n80694 & ~n80697;
  assign n80699 = n80280 & ~n80297;
  assign n80700 = ~n80288 & n80699;
  assign n80701 = ~n80268 & n80700;
  assign n80702 = ~n80309 & ~n80701;
  assign n80703 = ~n80348 & n80702;
  assign n80704 = ~n80291 & n80703;
  assign n80705 = n80698 & n80704;
  assign n80706 = ~n80262 & ~n80705;
  assign n80707 = n80281 & n80297;
  assign n80708 = n80288 & n80707;
  assign n80709 = ~n80325 & ~n80708;
  assign n80710 = ~n80706 & n80709;
  assign n80711 = n80690 & n80710;
  assign n80712 = pi2528 & ~n80711;
  assign n80713 = ~pi2528 & n80709;
  assign n80714 = n80690 & n80713;
  assign n80715 = ~n80706 & n80714;
  assign po2668 = n80712 | n80715;
  assign n80717 = ~n80419 & ~n80446;
  assign n80718 = n80401 & ~n80717;
  assign n80719 = ~n80405 & ~n80718;
  assign n80720 = ~n80380 & ~n80386;
  assign n80721 = ~n80380 & ~n80392;
  assign n80722 = ~n80374 & n80721;
  assign n80723 = n80374 & n80393;
  assign n80724 = ~n80722 & ~n80723;
  assign n80725 = ~n80720 & n80724;
  assign n80726 = ~n80430 & n80725;
  assign n80727 = ~n80401 & ~n80726;
  assign n80728 = n80719 & ~n80727;
  assign n80729 = ~n80522 & n80728;
  assign n80730 = n80368 & ~n80729;
  assign n80731 = ~n80374 & n80403;
  assign n80732 = n80523 & ~n80731;
  assign n80733 = ~n80401 & ~n80732;
  assign n80734 = ~n80730 & ~n80733;
  assign n80735 = ~n80380 & n80386;
  assign n80736 = n80401 & n80735;
  assign n80737 = n80374 & n80736;
  assign n80738 = n80374 & n80434;
  assign n80739 = ~n80374 & n80532;
  assign n80740 = ~n80738 & ~n80739;
  assign n80741 = n80380 & ~n80386;
  assign n80742 = n80374 & n80741;
  assign n80743 = ~n80411 & ~n80742;
  assign n80744 = n80401 & ~n80743;
  assign n80745 = n80401 & n80720;
  assign n80746 = ~n80374 & n80745;
  assign n80747 = ~n80744 & ~n80746;
  assign n80748 = n80740 & n80747;
  assign n80749 = ~n80368 & ~n80748;
  assign n80750 = ~n80737 & ~n80749;
  assign n80751 = ~n80406 & n80750;
  assign n80752 = n80734 & n80751;
  assign n80753 = ~pi2533 & ~n80752;
  assign n80754 = ~n80406 & ~n80730;
  assign n80755 = ~n80733 & n80754;
  assign n80756 = n80750 & n80755;
  assign n80757 = pi2533 & n80756;
  assign po2669 = n80753 | n80757;
  assign n80759 = n79988 & n80080;
  assign n80760 = n79959 & n79991;
  assign n80761 = ~n80084 & ~n80760;
  assign n80762 = ~n79965 & ~n80761;
  assign n80763 = ~n80759 & ~n80762;
  assign n80764 = ~n80012 & n80763;
  assign n80765 = ~n79959 & n79996;
  assign n80766 = ~n79991 & ~n80765;
  assign n80767 = ~n80095 & n80766;
  assign n80768 = ~n79965 & ~n80767;
  assign n80769 = n79934 & n80768;
  assign n80770 = n79965 & n80093;
  assign n80771 = ~n79984 & ~n80010;
  assign n80772 = ~n79975 & n80771;
  assign n80773 = ~n80770 & n80772;
  assign n80774 = n79934 & ~n80773;
  assign n80775 = n79940 & n79965;
  assign n80776 = n79952 & n80775;
  assign n80777 = ~n79946 & n80776;
  assign n80778 = ~n79959 & n80021;
  assign n80779 = ~n80777 & ~n80778;
  assign n80780 = ~n80083 & n80779;
  assign n80781 = n79952 & n79982;
  assign n80782 = ~n79959 & n79970;
  assign n80783 = ~n79987 & ~n80782;
  assign n80784 = ~n79965 & ~n80783;
  assign n80785 = ~n80781 & ~n80784;
  assign n80786 = n80780 & n80785;
  assign n80787 = ~n79934 & ~n80786;
  assign n80788 = n79959 & n80777;
  assign n80789 = ~n80787 & ~n80788;
  assign n80790 = ~n80774 & n80789;
  assign n80791 = ~n80769 & n80790;
  assign n80792 = n80764 & n80791;
  assign n80793 = pi2545 & ~n80792;
  assign n80794 = ~pi2545 & n80764;
  assign n80795 = n80791 & n80794;
  assign po2670 = n80793 | n80795;
  assign n80797 = ~n80330 & ~n80341;
  assign n80798 = ~n80274 & ~n80797;
  assign n80799 = n80280 & n80322;
  assign n80800 = ~n80798 & ~n80799;
  assign n80801 = n80268 & n80280;
  assign n80802 = ~n80307 & ~n80801;
  assign n80803 = ~n80680 & n80802;
  assign n80804 = n80274 & ~n80803;
  assign n80805 = n80800 & ~n80804;
  assign n80806 = n80262 & ~n80805;
  assign n80807 = ~n80344 & ~n80349;
  assign n80808 = n80290 & n80308;
  assign n80809 = n80807 & ~n80808;
  assign n80810 = n80274 & n80301;
  assign n80811 = n80280 & n80330;
  assign n80812 = ~n80274 & n80307;
  assign n80813 = ~n80811 & ~n80812;
  assign n80814 = ~n80701 & n80813;
  assign n80815 = ~n80810 & n80814;
  assign n80816 = ~n80348 & ~n80352;
  assign n80817 = n80815 & n80816;
  assign n80818 = ~n80315 & n80817;
  assign n80819 = ~n80262 & ~n80818;
  assign n80820 = n80809 & ~n80819;
  assign n80821 = ~n80806 & n80820;
  assign n80822 = ~pi2530 & ~n80821;
  assign n80823 = pi2530 & n80809;
  assign n80824 = ~n80806 & n80823;
  assign n80825 = ~n80819 & n80824;
  assign po2672 = n80822 | n80825;
  assign n80827 = ~n80449 & ~n80508;
  assign n80828 = ~n80425 & n80827;
  assign n80829 = n80401 & ~n80828;
  assign n80830 = ~n80516 & ~n80535;
  assign n80831 = ~n80435 & ~n80450;
  assign n80832 = ~n80394 & ~n80440;
  assign n80833 = ~n80401 & ~n80832;
  assign n80834 = ~n80406 & ~n80833;
  assign n80835 = n80831 & n80834;
  assign n80836 = n80368 & ~n80835;
  assign n80837 = ~n80380 & n80392;
  assign n80838 = ~n80720 & ~n80837;
  assign n80839 = n80374 & ~n80838;
  assign n80840 = ~n80442 & ~n80519;
  assign n80841 = ~n80401 & ~n80840;
  assign n80842 = n80374 & n80392;
  assign n80843 = ~n80446 & ~n80842;
  assign n80844 = ~n80393 & n80843;
  assign n80845 = n80401 & ~n80844;
  assign n80846 = ~n80841 & ~n80845;
  assign n80847 = ~n80839 & n80846;
  assign n80848 = ~n80368 & ~n80847;
  assign n80849 = ~n80836 & ~n80848;
  assign n80850 = n80830 & n80849;
  assign n80851 = ~n80829 & n80850;
  assign n80852 = ~pi2568 & ~n80851;
  assign n80853 = pi2568 & n80830;
  assign n80854 = ~n80829 & n80853;
  assign n80855 = n80849 & n80854;
  assign po2674 = n80852 | n80855;
  assign n80857 = n80274 & n80321;
  assign n80858 = ~n80280 & n80857;
  assign n80859 = ~n80353 & ~n80858;
  assign n80860 = n80280 & n80297;
  assign n80861 = n80288 & n80860;
  assign n80862 = ~n80268 & ~n80280;
  assign n80863 = ~n80352 & ~n80862;
  assign n80864 = ~n80274 & ~n80863;
  assign n80865 = ~n80861 & ~n80864;
  assign n80866 = n80859 & n80865;
  assign n80867 = ~n80262 & ~n80866;
  assign n80868 = ~n80305 & ~n80309;
  assign n80869 = ~n80280 & n80329;
  assign n80870 = n80868 & ~n80869;
  assign n80871 = n80274 & ~n80870;
  assign n80872 = n80290 & n80321;
  assign n80873 = ~n80325 & ~n80872;
  assign n80874 = ~n80871 & n80873;
  assign n80875 = ~n80680 & ~n80687;
  assign n80876 = ~n80274 & ~n80875;
  assign n80877 = n80874 & ~n80876;
  assign n80878 = n80262 & ~n80877;
  assign n80879 = ~n80867 & ~n80878;
  assign n80880 = ~n80280 & n80340;
  assign n80881 = n80280 & ~n80683;
  assign n80882 = ~n80880 & ~n80881;
  assign n80883 = ~n80274 & ~n80882;
  assign n80884 = ~n80305 & n80797;
  assign n80885 = n80311 & ~n80884;
  assign n80886 = ~n80883 & ~n80885;
  assign n80887 = n80879 & n80886;
  assign n80888 = ~pi2531 & ~n80887;
  assign n80889 = pi2531 & n80886;
  assign n80890 = ~n80878 & n80889;
  assign n80891 = ~n80867 & n80890;
  assign po2677 = n80888 | n80891;
  assign n80893 = ~n80147 & n80214;
  assign n80894 = ~n80156 & ~n80893;
  assign n80895 = ~n80134 & ~n80894;
  assign n80896 = n80128 & n80179;
  assign n80897 = ~n80170 & ~n80896;
  assign n80898 = n80134 & ~n80897;
  assign n80899 = ~n80128 & n80222;
  assign n80900 = ~n80195 & ~n80899;
  assign n80901 = ~n80213 & n80900;
  assign n80902 = ~n80898 & n80901;
  assign n80903 = ~n80895 & n80902;
  assign n80904 = ~n80164 & ~n80178;
  assign n80905 = n80903 & n80904;
  assign n80906 = n80122 & ~n80905;
  assign n80907 = n80166 & n80189;
  assign n80908 = n80238 & ~n80907;
  assign n80909 = n80134 & ~n80908;
  assign n80910 = ~n80128 & n80230;
  assign n80911 = ~n80909 & ~n80910;
  assign n80912 = n80141 & n80214;
  assign n80913 = n80128 & n80155;
  assign n80914 = ~n80912 & ~n80913;
  assign n80915 = n80134 & ~n80914;
  assign n80916 = n80134 & n80179;
  assign n80917 = ~n80128 & n80916;
  assign n80918 = ~n80915 & ~n80917;
  assign n80919 = n80911 & n80918;
  assign n80920 = ~n80122 & ~n80919;
  assign n80921 = ~n80222 & ~n80227;
  assign n80922 = ~n80171 & n80921;
  assign n80923 = n80245 & ~n80922;
  assign n80924 = ~n80920 & ~n80923;
  assign n80925 = ~n80164 & ~n80213;
  assign n80926 = ~n80134 & ~n80925;
  assign n80927 = n80924 & ~n80926;
  assign n80928 = ~n80906 & n80927;
  assign n80929 = ~pi2562 & n80928;
  assign n80930 = pi2562 & ~n80928;
  assign po2678 = n80929 | n80930;
  assign n80932 = ~n80128 & n80155;
  assign n80933 = ~n80220 & ~n80932;
  assign n80934 = ~n80134 & ~n80933;
  assign n80935 = n80134 & ~n80197;
  assign n80936 = ~n80185 & ~n80935;
  assign n80937 = ~n80934 & n80936;
  assign n80938 = n80122 & ~n80937;
  assign n80939 = ~n80134 & n80230;
  assign n80940 = ~n80938 & ~n80939;
  assign n80941 = ~n80899 & ~n80913;
  assign n80942 = n80134 & ~n80941;
  assign n80943 = n80134 & n80163;
  assign n80944 = n80147 & n80214;
  assign n80945 = n80141 & n80944;
  assign n80946 = ~n80134 & n80176;
  assign n80947 = ~n80169 & ~n80946;
  assign n80948 = ~n80141 & ~n80947;
  assign n80949 = ~n80170 & ~n80948;
  assign n80950 = ~n80213 & n80949;
  assign n80951 = ~n80945 & n80950;
  assign n80952 = ~n80943 & n80951;
  assign n80953 = ~n80122 & ~n80952;
  assign n80954 = ~n80942 & ~n80953;
  assign n80955 = n80940 & n80954;
  assign n80956 = pi2574 & ~n80955;
  assign n80957 = ~pi2574 & n80955;
  assign po2680 = n80956 | n80957;
  assign n80959 = pi5285 & pi9040;
  assign n80960 = ~pi5546 & ~pi9040;
  assign n80961 = ~n80959 & ~n80960;
  assign n80962 = ~pi2499 & ~n80961;
  assign n80963 = pi2499 & n80961;
  assign n80964 = ~n80962 & ~n80963;
  assign n80965 = pi5337 & pi9040;
  assign n80966 = pi5334 & ~pi9040;
  assign n80967 = ~n80965 & ~n80966;
  assign n80968 = ~pi2516 & n80967;
  assign n80969 = pi2516 & ~n80967;
  assign n80970 = ~n80968 & ~n80969;
  assign n80971 = pi5358 & ~pi9040;
  assign n80972 = pi5378 & pi9040;
  assign n80973 = ~n80971 & ~n80972;
  assign n80974 = ~pi2508 & n80973;
  assign n80975 = pi2508 & ~n80973;
  assign n80976 = ~n80974 & ~n80975;
  assign n80977 = n80970 & ~n80976;
  assign n80978 = pi5203 & ~pi9040;
  assign n80979 = pi5421 & pi9040;
  assign n80980 = ~n80978 & ~n80979;
  assign n80981 = pi2505 & n80980;
  assign n80982 = ~pi2505 & ~n80980;
  assign n80983 = ~n80981 & ~n80982;
  assign n80984 = pi5207 & pi9040;
  assign n80985 = pi5543 & ~pi9040;
  assign n80986 = ~n80984 & ~n80985;
  assign n80987 = ~pi2491 & ~n80986;
  assign n80988 = pi2491 & n80986;
  assign n80989 = ~n80987 & ~n80988;
  assign n80990 = ~n80983 & ~n80989;
  assign n80991 = n80977 & n80990;
  assign n80992 = pi5285 & ~pi9040;
  assign n80993 = pi5628 & pi9040;
  assign n80994 = ~n80992 & ~n80993;
  assign n80995 = pi2520 & n80994;
  assign n80996 = ~pi2520 & ~n80994;
  assign n80997 = ~n80995 & ~n80996;
  assign n80998 = ~n80970 & n80976;
  assign n80999 = n80997 & n80998;
  assign n81000 = n80983 & ~n80997;
  assign n81001 = n80976 & n81000;
  assign n81002 = n80970 & n81001;
  assign n81003 = ~n80999 & ~n81002;
  assign n81004 = ~n80970 & ~n80976;
  assign n81005 = n80983 & n81004;
  assign n81006 = n81003 & ~n81005;
  assign n81007 = ~n80989 & ~n81006;
  assign n81008 = ~n80970 & ~n80997;
  assign n81009 = ~n80983 & n80989;
  assign n81010 = n81008 & n81009;
  assign n81011 = ~n80997 & n80998;
  assign n81012 = ~n80983 & n81011;
  assign n81013 = ~n81010 & ~n81012;
  assign n81014 = ~n81007 & n81013;
  assign n81015 = ~n80991 & n81014;
  assign n81016 = n80977 & n80997;
  assign n81017 = ~n80983 & n81016;
  assign n81018 = n80997 & n81004;
  assign n81019 = n80983 & n81018;
  assign n81020 = ~n81017 & ~n81019;
  assign n81021 = n81015 & n81020;
  assign n81022 = ~n80964 & ~n81021;
  assign n81023 = ~n80997 & n81004;
  assign n81024 = ~n80983 & n81023;
  assign n81025 = ~n81016 & ~n81024;
  assign n81026 = ~n80989 & ~n81025;
  assign n81027 = n80977 & n81000;
  assign n81028 = ~n80983 & ~n80997;
  assign n81029 = n80976 & n81028;
  assign n81030 = n80970 & n81029;
  assign n81031 = ~n81027 & ~n81030;
  assign n81032 = ~n80970 & n81000;
  assign n81033 = ~n80983 & n81018;
  assign n81034 = ~n81032 & ~n81033;
  assign n81035 = n80989 & ~n81034;
  assign n81036 = n81031 & ~n81035;
  assign n81037 = ~n81026 & n81036;
  assign n81038 = n80964 & ~n81037;
  assign n81039 = ~n80970 & n80997;
  assign n81040 = n80983 & n81039;
  assign n81041 = n80970 & n80997;
  assign n81042 = ~n80983 & n81041;
  assign n81043 = ~n81040 & ~n81042;
  assign n81044 = ~n80989 & ~n81043;
  assign n81045 = n80970 & n80976;
  assign n81046 = n80997 & n81045;
  assign n81047 = n80983 & n81046;
  assign n81048 = ~n81027 & ~n81047;
  assign n81049 = ~n81011 & n81048;
  assign n81050 = n80989 & ~n81049;
  assign n81051 = ~n81044 & ~n81050;
  assign n81052 = n80976 & ~n80997;
  assign n81053 = n80989 & n81052;
  assign n81054 = ~n80983 & n81053;
  assign n81055 = n81051 & ~n81054;
  assign n81056 = ~n81038 & n81055;
  assign n81057 = ~n81022 & n81056;
  assign n81058 = ~pi2534 & ~n81057;
  assign n81059 = pi2534 & n81057;
  assign po2682 = n81058 | n81059;
  assign n81061 = n80983 & n81011;
  assign n81062 = ~n81030 & ~n81039;
  assign n81063 = n80989 & ~n81062;
  assign n81064 = ~n81061 & ~n81063;
  assign n81065 = ~n81024 & n81064;
  assign n81066 = ~n80989 & n81027;
  assign n81067 = ~n81017 & ~n81066;
  assign n81068 = ~n81047 & n81067;
  assign n81069 = n81065 & n81068;
  assign n81070 = n80964 & ~n81069;
  assign n81071 = ~n80976 & n81000;
  assign n81072 = ~n80970 & n81071;
  assign n81073 = ~n81002 & ~n81072;
  assign n81074 = n80977 & ~n80997;
  assign n81075 = n80989 & n81074;
  assign n81076 = n80983 & n81016;
  assign n81077 = ~n81075 & ~n81076;
  assign n81078 = ~n80976 & n80997;
  assign n81079 = ~n80970 & n80983;
  assign n81080 = ~n81078 & ~n81079;
  assign n81081 = ~n81052 & n81080;
  assign n81082 = ~n80989 & ~n81081;
  assign n81083 = ~n80983 & n81046;
  assign n81084 = ~n81012 & ~n81083;
  assign n81085 = ~n81082 & n81084;
  assign n81086 = n81077 & n81085;
  assign n81087 = n81073 & n81086;
  assign n81088 = ~n80964 & ~n81087;
  assign n81089 = ~n81070 & ~n81088;
  assign n81090 = pi2529 & ~n81089;
  assign n81091 = ~pi2529 & ~n81070;
  assign n81092 = ~n81088 & n81091;
  assign po2683 = n81090 | n81092;
  assign n81094 = ~n80983 & n81004;
  assign n81095 = ~n81083 & ~n81094;
  assign n81096 = n80989 & n81095;
  assign n81097 = n80983 & n81041;
  assign n81098 = ~n80977 & ~n80998;
  assign n81099 = n80997 & ~n81098;
  assign n81100 = n80970 & n81028;
  assign n81101 = n80983 & n80998;
  assign n81102 = ~n81100 & ~n81101;
  assign n81103 = ~n80989 & n81102;
  assign n81104 = ~n81099 & n81103;
  assign n81105 = ~n81097 & n81104;
  assign n81106 = ~n81096 & ~n81105;
  assign n81107 = n80983 & n81099;
  assign n81108 = ~n81072 & ~n81107;
  assign n81109 = ~n81106 & n81108;
  assign n81110 = n80964 & ~n81109;
  assign n81111 = n80989 & ~n81098;
  assign n81112 = ~n80983 & n81111;
  assign n81113 = ~n81018 & ~n81045;
  assign n81114 = n80983 & ~n81113;
  assign n81115 = n80989 & n81114;
  assign n81116 = ~n80997 & n81111;
  assign n81117 = ~n81115 & ~n81116;
  assign n81118 = ~n81112 & n81117;
  assign n81119 = ~n80964 & ~n81118;
  assign n81120 = ~n81110 & ~n81119;
  assign n81121 = n80989 & n81002;
  assign n81122 = ~n80989 & ~n81108;
  assign n81123 = ~n81121 & ~n81122;
  assign n81124 = ~n80989 & ~n81095;
  assign n81125 = ~n81002 & ~n81124;
  assign n81126 = ~n80964 & ~n81125;
  assign n81127 = n81123 & ~n81126;
  assign n81128 = n81120 & n81127;
  assign n81129 = pi2539 & ~n81128;
  assign n81130 = ~pi2539 & n81127;
  assign n81131 = ~n81119 & n81130;
  assign n81132 = ~n81110 & n81131;
  assign po2684 = n81129 | n81132;
  assign n81134 = ~n80605 & ~n80612;
  assign n81135 = n80578 & ~n81134;
  assign n81136 = ~n80665 & ~n81135;
  assign n81137 = n80584 & n80590;
  assign n81138 = ~n80578 & n81137;
  assign n81139 = n80604 & n81138;
  assign n81140 = n80604 & n80619;
  assign n81141 = ~n81137 & ~n81140;
  assign n81142 = ~n80584 & ~n80604;
  assign n81143 = ~n80590 & n81142;
  assign n81144 = n81141 & ~n81143;
  assign n81145 = ~n80578 & ~n81144;
  assign n81146 = ~n80615 & ~n81145;
  assign n81147 = ~n80643 & ~n81146;
  assign n81148 = n80578 & n80597;
  assign n81149 = n80604 & n81148;
  assign n81150 = n80578 & n80653;
  assign n81151 = ~n81149 & ~n81150;
  assign n81152 = ~n80643 & ~n81151;
  assign n81153 = ~n81147 & ~n81152;
  assign n81154 = ~n81139 & n81153;
  assign n81155 = ~n80590 & n80606;
  assign n81156 = ~n80607 & ~n80624;
  assign n81157 = ~n80584 & n80613;
  assign n81158 = n81156 & ~n81157;
  assign n81159 = n80578 & ~n81158;
  assign n81160 = ~n80604 & n80653;
  assign n81161 = ~n80634 & ~n81160;
  assign n81162 = ~n80578 & ~n81161;
  assign n81163 = ~n81159 & ~n81162;
  assign n81164 = ~n81155 & n81163;
  assign n81165 = ~n80621 & ~n80659;
  assign n81166 = n81164 & n81165;
  assign n81167 = n80643 & ~n81166;
  assign n81168 = n81154 & ~n81167;
  assign n81169 = n81136 & n81168;
  assign n81170 = ~pi2573 & ~n81169;
  assign n81171 = pi2573 & n81154;
  assign n81172 = n81136 & n81171;
  assign n81173 = ~n81167 & n81172;
  assign po2685 = n81170 | n81173;
  assign n81175 = ~n80604 & n80634;
  assign n81176 = n80604 & n80645;
  assign n81177 = ~n80624 & ~n81176;
  assign n81178 = ~n80578 & ~n81177;
  assign n81179 = ~n81175 & ~n81178;
  assign n81180 = n80578 & ~n80604;
  assign n81181 = ~n80596 & n81180;
  assign n81182 = ~n80590 & n81181;
  assign n81183 = n80613 & n80646;
  assign n81184 = ~n81182 & ~n81183;
  assign n81185 = ~n81150 & n81184;
  assign n81186 = ~n80608 & ~n80621;
  assign n81187 = ~n80658 & n81186;
  assign n81188 = n81185 & n81187;
  assign n81189 = n81179 & n81188;
  assign n81190 = ~n80643 & ~n81189;
  assign n81191 = n80584 & n80610;
  assign n81192 = ~n80624 & ~n81191;
  assign n81193 = n80604 & ~n81192;
  assign n81194 = ~n81155 & ~n81157;
  assign n81195 = ~n80584 & ~n80596;
  assign n81196 = n80604 & n81195;
  assign n81197 = n81194 & ~n81196;
  assign n81198 = ~n80578 & ~n81197;
  assign n81199 = ~n80604 & n80619;
  assign n81200 = n80598 & n80604;
  assign n81201 = ~n81199 & ~n81200;
  assign n81202 = n80578 & ~n81201;
  assign n81203 = ~n80604 & n80614;
  assign n81204 = ~n81202 & ~n81203;
  assign n81205 = ~n81198 & n81204;
  assign n81206 = ~n81193 & n81205;
  assign n81207 = n80643 & ~n81206;
  assign n81208 = ~n80578 & n80607;
  assign n81209 = ~n81207 & ~n81208;
  assign n81210 = n80628 & n81180;
  assign n81211 = ~n80596 & n81210;
  assign n81212 = n81209 & ~n81211;
  assign n81213 = ~n81190 & n81212;
  assign n81214 = ~pi2567 & ~n81213;
  assign n81215 = pi2567 & n81209;
  assign n81216 = ~n81190 & n81215;
  assign n81217 = ~n81211 & n81216;
  assign po2686 = n81214 | n81217;
  assign n81219 = pi5212 & ~pi9040;
  assign n81220 = pi5333 & pi9040;
  assign n81221 = ~n81219 & ~n81220;
  assign n81222 = ~pi2514 & ~n81221;
  assign n81223 = pi2514 & n81221;
  assign n81224 = ~n81222 & ~n81223;
  assign n81225 = pi5348 & ~pi9040;
  assign n81226 = pi5340 & pi9040;
  assign n81227 = ~n81225 & ~n81226;
  assign n81228 = pi2511 & n81227;
  assign n81229 = ~pi2511 & ~n81227;
  assign n81230 = ~n81228 & ~n81229;
  assign n81231 = pi5662 & ~pi9040;
  assign n81232 = pi5338 & pi9040;
  assign n81233 = ~n81231 & ~n81232;
  assign n81234 = pi2526 & n81233;
  assign n81235 = ~pi2526 & ~n81233;
  assign n81236 = ~n81234 & ~n81235;
  assign n81237 = ~n81230 & n81236;
  assign n81238 = n81224 & n81237;
  assign n81239 = pi5333 & ~pi9040;
  assign n81240 = pi5346 & pi9040;
  assign n81241 = ~n81239 & ~n81240;
  assign n81242 = ~pi2513 & n81241;
  assign n81243 = pi2513 & ~n81241;
  assign n81244 = ~n81242 & ~n81243;
  assign n81245 = ~n81224 & ~n81244;
  assign n81246 = ~n81236 & n81245;
  assign n81247 = n81224 & ~n81244;
  assign n81248 = n81236 & n81247;
  assign n81249 = ~n81246 & ~n81248;
  assign n81250 = ~n81238 & n81249;
  assign n81251 = pi5341 & ~pi9040;
  assign n81252 = pi5662 & pi9040;
  assign n81253 = ~n81251 & ~n81252;
  assign n81254 = pi2498 & n81253;
  assign n81255 = ~pi2498 & ~n81253;
  assign n81256 = ~n81254 & ~n81255;
  assign n81257 = pi5292 & ~pi9040;
  assign n81258 = pi5294 & pi9040;
  assign n81259 = ~n81257 & ~n81258;
  assign n81260 = ~pi2482 & ~n81259;
  assign n81261 = pi2482 & n81259;
  assign n81262 = ~n81260 & ~n81261;
  assign n81263 = n81256 & n81262;
  assign n81264 = ~n81250 & n81263;
  assign n81265 = ~n81224 & n81244;
  assign n81266 = n81236 & n81265;
  assign n81267 = n81230 & n81262;
  assign n81268 = n81266 & n81267;
  assign n81269 = n81236 & n81245;
  assign n81270 = ~n81256 & n81269;
  assign n81271 = n81224 & n81244;
  assign n81272 = n81230 & n81271;
  assign n81273 = n81224 & ~n81236;
  assign n81274 = ~n81272 & ~n81273;
  assign n81275 = ~n81256 & ~n81274;
  assign n81276 = ~n81270 & ~n81275;
  assign n81277 = n81262 & ~n81276;
  assign n81278 = ~n81268 & ~n81277;
  assign n81279 = n81230 & ~n81236;
  assign n81280 = n81224 & n81279;
  assign n81281 = ~n81230 & n81265;
  assign n81282 = ~n81236 & n81281;
  assign n81283 = ~n81280 & ~n81282;
  assign n81284 = ~n81256 & ~n81283;
  assign n81285 = n81278 & ~n81284;
  assign n81286 = n81230 & n81256;
  assign n81287 = n81271 & n81286;
  assign n81288 = n81236 & n81287;
  assign n81289 = ~n81236 & n81271;
  assign n81290 = ~n81230 & n81256;
  assign n81291 = n81289 & n81290;
  assign n81292 = ~n81247 & ~n81265;
  assign n81293 = n81279 & ~n81292;
  assign n81294 = n81230 & n81269;
  assign n81295 = ~n81293 & ~n81294;
  assign n81296 = n81237 & ~n81292;
  assign n81297 = ~n81230 & n81246;
  assign n81298 = ~n81296 & ~n81297;
  assign n81299 = n81295 & n81298;
  assign n81300 = ~n81291 & n81299;
  assign n81301 = ~n81288 & n81300;
  assign n81302 = ~n81230 & ~n81256;
  assign n81303 = n81236 & n81302;
  assign n81304 = n81244 & n81303;
  assign n81305 = n81301 & ~n81304;
  assign n81306 = ~n81262 & ~n81305;
  assign n81307 = n81285 & ~n81306;
  assign n81308 = ~n81264 & n81307;
  assign n81309 = ~pi2555 & ~n81308;
  assign n81310 = pi2555 & n81285;
  assign n81311 = ~n81264 & n81310;
  assign n81312 = ~n81306 & n81311;
  assign po2687 = n81309 | n81312;
  assign n81314 = n80983 & n81074;
  assign n81315 = n80989 & n81314;
  assign n81316 = n81028 & ~n81098;
  assign n81317 = ~n81046 & ~n81316;
  assign n81318 = ~n81072 & n81317;
  assign n81319 = ~n80989 & ~n81318;
  assign n81320 = n80983 & n80999;
  assign n81321 = ~n81319 & ~n81320;
  assign n81322 = ~n80997 & n81045;
  assign n81323 = ~n80983 & n81078;
  assign n81324 = ~n81322 & ~n81323;
  assign n81325 = ~n81101 & n81324;
  assign n81326 = n80989 & ~n81325;
  assign n81327 = n81321 & ~n81326;
  assign n81328 = n80964 & ~n81327;
  assign n81329 = ~n81315 & ~n81328;
  assign n81330 = ~n80983 & n80998;
  assign n81331 = ~n81023 & ~n81330;
  assign n81332 = n80989 & ~n81331;
  assign n81333 = ~n81047 & ~n81332;
  assign n81334 = ~n81019 & ~n81314;
  assign n81335 = n80983 & n81052;
  assign n81336 = ~n81078 & ~n81335;
  assign n81337 = ~n81322 & n81336;
  assign n81338 = ~n80989 & ~n81337;
  assign n81339 = ~n80983 & n80999;
  assign n81340 = ~n81338 & ~n81339;
  assign n81341 = n81334 & n81340;
  assign n81342 = n81333 & n81341;
  assign n81343 = ~n80964 & ~n81342;
  assign n81344 = ~n81033 & ~n81097;
  assign n81345 = ~n80989 & ~n81344;
  assign n81346 = ~n81343 & ~n81345;
  assign n81347 = n81329 & n81346;
  assign n81348 = pi2543 & n81347;
  assign n81349 = ~pi2543 & ~n81347;
  assign po2688 = n81348 | n81349;
  assign n81351 = n81230 & n81265;
  assign n81352 = ~n81230 & n81271;
  assign n81353 = ~n81351 & ~n81352;
  assign n81354 = ~n81256 & ~n81353;
  assign n81355 = n81245 & n81302;
  assign n81356 = ~n81236 & n81355;
  assign n81357 = ~n81354 & ~n81356;
  assign n81358 = n81262 & ~n81357;
  assign n81359 = ~n81230 & ~n81236;
  assign n81360 = ~n81292 & n81359;
  assign n81361 = n81236 & n81271;
  assign n81362 = ~n81236 & ~n81244;
  assign n81363 = ~n81247 & ~n81362;
  assign n81364 = ~n81230 & ~n81363;
  assign n81365 = ~n81361 & ~n81364;
  assign n81366 = n81256 & ~n81365;
  assign n81367 = ~n81360 & ~n81366;
  assign n81368 = n81230 & n81289;
  assign n81369 = ~n81224 & n81237;
  assign n81370 = n81230 & ~n81363;
  assign n81371 = ~n81369 & ~n81370;
  assign n81372 = ~n81256 & ~n81371;
  assign n81373 = ~n81368 & ~n81372;
  assign n81374 = n81367 & n81373;
  assign n81375 = ~n81262 & ~n81374;
  assign n81376 = n81236 & n81262;
  assign n81377 = ~n81247 & n81376;
  assign n81378 = n81230 & n81377;
  assign n81379 = n81247 & n81279;
  assign n81380 = ~n81256 & n81379;
  assign n81381 = n81236 & n81286;
  assign n81382 = ~n81224 & n81381;
  assign n81383 = ~n81380 & ~n81382;
  assign n81384 = ~n81378 & n81383;
  assign n81385 = n81230 & ~n81244;
  assign n81386 = ~n81266 & ~n81385;
  assign n81387 = n81263 & ~n81386;
  assign n81388 = n81384 & ~n81387;
  assign n81389 = ~n81375 & n81388;
  assign n81390 = ~n81358 & n81389;
  assign n81391 = pi2550 & ~n81390;
  assign n81392 = ~pi2550 & n81390;
  assign po2689 = n81391 | n81392;
  assign n81394 = ~n81256 & n81361;
  assign n81395 = ~n81230 & n81394;
  assign n81396 = ~n81356 & ~n81395;
  assign n81397 = ~n81291 & ~n81297;
  assign n81398 = n81236 & ~n81244;
  assign n81399 = n81230 & n81398;
  assign n81400 = ~n81272 & ~n81399;
  assign n81401 = ~n81256 & ~n81400;
  assign n81402 = n81256 & ~n81359;
  assign n81403 = ~n81292 & n81402;
  assign n81404 = ~n81230 & ~n81271;
  assign n81405 = ~n81256 & n81404;
  assign n81406 = ~n81236 & n81405;
  assign n81407 = ~n81403 & ~n81406;
  assign n81408 = ~n81401 & n81407;
  assign n81409 = n81397 & n81408;
  assign n81410 = n81262 & ~n81409;
  assign n81411 = n81396 & ~n81410;
  assign n81412 = n81248 & n81256;
  assign n81413 = n81230 & n81412;
  assign n81414 = n81256 & ~n81262;
  assign n81415 = ~n81269 & ~n81272;
  assign n81416 = ~n81360 & n81415;
  assign n81417 = n81414 & ~n81416;
  assign n81418 = n81230 & n81246;
  assign n81419 = ~n81236 & n81385;
  assign n81420 = ~n81351 & ~n81419;
  assign n81421 = ~n81266 & ~n81352;
  assign n81422 = n81420 & n81421;
  assign n81423 = ~n81256 & ~n81422;
  assign n81424 = ~n81418 & ~n81423;
  assign n81425 = ~n81262 & ~n81424;
  assign n81426 = ~n81417 & ~n81425;
  assign n81427 = ~n81413 & n81426;
  assign n81428 = n81411 & n81427;
  assign n81429 = pi2551 & ~n81428;
  assign n81430 = ~pi2551 & n81411;
  assign n81431 = n81427 & n81430;
  assign po2691 = n81429 | n81431;
  assign n81433 = ~n81236 & n81247;
  assign n81434 = ~n81361 & ~n81433;
  assign n81435 = ~n81256 & ~n81434;
  assign n81436 = ~n81248 & ~n81281;
  assign n81437 = ~n81289 & n81436;
  assign n81438 = n81256 & ~n81437;
  assign n81439 = ~n81435 & ~n81438;
  assign n81440 = ~n81270 & ~n81282;
  assign n81441 = n81439 & n81440;
  assign n81442 = ~n81262 & ~n81441;
  assign n81443 = n81230 & n81361;
  assign n81444 = ~n81230 & n81245;
  assign n81445 = ~n81351 & ~n81444;
  assign n81446 = n81256 & ~n81445;
  assign n81447 = ~n81443 & ~n81446;
  assign n81448 = n81236 & ~n81256;
  assign n81449 = ~n81224 & n81448;
  assign n81450 = n81244 & n81449;
  assign n81451 = n81249 & ~n81450;
  assign n81452 = ~n81289 & n81451;
  assign n81453 = ~n81230 & ~n81452;
  assign n81454 = n81447 & ~n81453;
  assign n81455 = n81262 & ~n81454;
  assign n81456 = ~n81442 & ~n81455;
  assign n81457 = ~n81236 & n81351;
  assign n81458 = ~n81294 & ~n81457;
  assign n81459 = ~n81256 & ~n81458;
  assign n81460 = n81256 & n81362;
  assign n81461 = n81230 & n81460;
  assign n81462 = ~n81459 & ~n81461;
  assign n81463 = n81456 & n81462;
  assign n81464 = ~pi2556 & ~n81463;
  assign n81465 = pi2556 & ~n81459;
  assign n81466 = n81456 & n81465;
  assign n81467 = ~n81461 & n81466;
  assign po2692 = n81464 | n81467;
  assign n81469 = ~n80659 & ~n81203;
  assign n81470 = ~n80578 & ~n81469;
  assign n81471 = ~n80643 & n80645;
  assign n81472 = n80578 & n81471;
  assign n81473 = n80590 & n81142;
  assign n81474 = ~n81195 & ~n81473;
  assign n81475 = ~n80614 & n81474;
  assign n81476 = ~n80578 & ~n81475;
  assign n81477 = ~n80604 & n80620;
  assign n81478 = ~n81476 & ~n81477;
  assign n81479 = ~n80643 & ~n81478;
  assign n81480 = ~n81472 & ~n81479;
  assign n81481 = ~n80608 & ~n80612;
  assign n81482 = ~n80604 & n81157;
  assign n81483 = ~n81176 & ~n81482;
  assign n81484 = n81481 & n81483;
  assign n81485 = n80578 & ~n81484;
  assign n81486 = n80584 & ~n80590;
  assign n81487 = n80578 & n81486;
  assign n81488 = n80604 & n81487;
  assign n81489 = ~n80604 & n81195;
  assign n81490 = ~n80612 & ~n81489;
  assign n81491 = ~n81200 & n81490;
  assign n81492 = ~n81488 & n81491;
  assign n81493 = ~n80578 & n81191;
  assign n81494 = n81492 & ~n81493;
  assign n81495 = n80643 & ~n81494;
  assign n81496 = ~n81485 & ~n81495;
  assign n81497 = n81480 & n81496;
  assign n81498 = ~n81470 & n81497;
  assign n81499 = pi2588 & n81498;
  assign n81500 = ~pi2588 & ~n81498;
  assign po2693 = n81499 | n81500;
  assign n81502 = pi5634 & pi9040;
  assign n81503 = pi5793 & ~pi9040;
  assign n81504 = ~n81502 & ~n81503;
  assign n81505 = ~pi2569 & ~n81504;
  assign n81506 = pi2569 & n81504;
  assign n81507 = ~n81505 & ~n81506;
  assign n81508 = pi5532 & pi9040;
  assign n81509 = pi5618 & ~pi9040;
  assign n81510 = ~n81508 & ~n81509;
  assign n81511 = pi2537 & n81510;
  assign n81512 = ~pi2537 & ~n81510;
  assign n81513 = ~n81511 & ~n81512;
  assign n81514 = pi5619 & ~pi9040;
  assign n81515 = pi5537 & pi9040;
  assign n81516 = ~n81514 & ~n81515;
  assign n81517 = ~pi2570 & n81516;
  assign n81518 = pi2570 & ~n81516;
  assign n81519 = ~n81517 & ~n81518;
  assign n81520 = pi5562 & pi9040;
  assign n81521 = pi5626 & ~pi9040;
  assign n81522 = ~n81520 & ~n81521;
  assign n81523 = ~pi2578 & n81522;
  assign n81524 = pi2578 & ~n81522;
  assign n81525 = ~n81523 & ~n81524;
  assign n81526 = ~n81519 & ~n81525;
  assign n81527 = ~n81513 & n81526;
  assign n81528 = pi5530 & ~pi9040;
  assign n81529 = pi5459 & pi9040;
  assign n81530 = ~n81528 & ~n81529;
  assign n81531 = ~pi2577 & ~n81530;
  assign n81532 = pi2577 & n81530;
  assign n81533 = ~n81531 & ~n81532;
  assign n81534 = n81527 & ~n81533;
  assign n81535 = n81519 & n81525;
  assign n81536 = ~n81513 & n81535;
  assign n81537 = ~n81533 & n81536;
  assign n81538 = ~n81534 & ~n81537;
  assign n81539 = n81513 & n81535;
  assign n81540 = n81533 & n81539;
  assign n81541 = ~n81513 & n81533;
  assign n81542 = n81525 & n81541;
  assign n81543 = ~n81519 & n81542;
  assign n81544 = ~n81540 & ~n81543;
  assign n81545 = n81538 & n81544;
  assign n81546 = n81507 & ~n81545;
  assign n81547 = ~n81525 & n81541;
  assign n81548 = n81519 & n81547;
  assign n81549 = ~n81519 & n81525;
  assign n81550 = ~n81513 & n81549;
  assign n81551 = ~n81548 & ~n81550;
  assign n81552 = n81507 & ~n81551;
  assign n81553 = ~n81507 & ~n81525;
  assign n81554 = ~n81533 & n81553;
  assign n81555 = n81513 & ~n81519;
  assign n81556 = n81533 & n81535;
  assign n81557 = ~n81555 & ~n81556;
  assign n81558 = ~n81507 & ~n81557;
  assign n81559 = ~n81554 & ~n81558;
  assign n81560 = n81519 & ~n81525;
  assign n81561 = n81513 & n81560;
  assign n81562 = ~n81533 & n81561;
  assign n81563 = n81559 & ~n81562;
  assign n81564 = ~n81525 & n81555;
  assign n81565 = n81533 & n81564;
  assign n81566 = n81563 & ~n81565;
  assign n81567 = ~n81552 & n81566;
  assign n81568 = pi5608 & pi9040;
  assign n81569 = pi5882 & ~pi9040;
  assign n81570 = ~n81568 & ~n81569;
  assign n81571 = ~pi2575 & ~n81570;
  assign n81572 = pi2575 & n81570;
  assign n81573 = ~n81571 & ~n81572;
  assign n81574 = ~n81567 & ~n81573;
  assign n81575 = ~n81513 & ~n81525;
  assign n81576 = ~n81507 & n81533;
  assign n81577 = n81573 & n81576;
  assign n81578 = n81575 & n81577;
  assign n81579 = ~n81513 & ~n81533;
  assign n81580 = n81525 & n81579;
  assign n81581 = ~n81507 & ~n81580;
  assign n81582 = ~n81526 & ~n81575;
  assign n81583 = ~n81533 & ~n81582;
  assign n81584 = n81513 & n81533;
  assign n81585 = n81519 & n81584;
  assign n81586 = ~n81539 & ~n81585;
  assign n81587 = ~n81583 & n81586;
  assign n81588 = n81507 & n81587;
  assign n81589 = ~n81581 & ~n81588;
  assign n81590 = n81513 & n81549;
  assign n81591 = n81533 & n81590;
  assign n81592 = ~n81589 & ~n81591;
  assign n81593 = n81573 & ~n81592;
  assign n81594 = ~n81578 & ~n81593;
  assign n81595 = ~n81574 & n81594;
  assign n81596 = ~n81546 & n81595;
  assign n81597 = ~n81507 & n81562;
  assign n81598 = n81596 & ~n81597;
  assign n81599 = pi2598 & ~n81598;
  assign n81600 = ~pi2598 & ~n81597;
  assign n81601 = n81595 & n81600;
  assign n81602 = ~n81546 & n81601;
  assign po2699 = n81599 | n81602;
  assign n81604 = pi5464 & pi9040;
  assign n81605 = pi5633 & ~pi9040;
  assign n81606 = ~n81604 & ~n81605;
  assign n81607 = pi2589 & n81606;
  assign n81608 = ~pi2589 & ~n81606;
  assign n81609 = ~n81607 & ~n81608;
  assign n81610 = pi5636 & ~pi9040;
  assign n81611 = pi5802 & pi9040;
  assign n81612 = ~n81610 & ~n81611;
  assign n81613 = ~pi2563 & ~n81612;
  assign n81614 = pi2563 & n81612;
  assign n81615 = ~n81613 & ~n81614;
  assign n81616 = pi5450 & ~pi9040;
  assign n81617 = pi5552 & pi9040;
  assign n81618 = ~n81616 & ~n81617;
  assign n81619 = pi2554 & n81618;
  assign n81620 = ~pi2554 & ~n81618;
  assign n81621 = ~n81619 & ~n81620;
  assign n81622 = pi5625 & ~pi9040;
  assign n81623 = pi5547 & pi9040;
  assign n81624 = ~n81622 & ~n81623;
  assign n81625 = ~pi2576 & n81624;
  assign n81626 = pi2576 & ~n81624;
  assign n81627 = ~n81625 & ~n81626;
  assign n81628 = n81621 & ~n81627;
  assign n81629 = n81615 & n81628;
  assign n81630 = n81621 & n81627;
  assign n81631 = ~n81615 & n81630;
  assign n81632 = ~n81629 & ~n81631;
  assign n81633 = ~n81609 & ~n81632;
  assign n81634 = pi5685 & ~pi9040;
  assign n81635 = pi5449 & pi9040;
  assign n81636 = ~n81634 & ~n81635;
  assign n81637 = ~pi2578 & ~n81636;
  assign n81638 = pi2578 & n81636;
  assign n81639 = ~n81637 & ~n81638;
  assign n81640 = pi5449 & ~pi9040;
  assign n81641 = pi5625 & pi9040;
  assign n81642 = ~n81640 & ~n81641;
  assign n81643 = ~pi2537 & ~n81642;
  assign n81644 = pi2537 & n81642;
  assign n81645 = ~n81643 & ~n81644;
  assign n81646 = n81627 & n81645;
  assign n81647 = n81615 & ~n81621;
  assign n81648 = n81646 & n81647;
  assign n81649 = ~n81615 & ~n81621;
  assign n81650 = ~n81645 & n81649;
  assign n81651 = n81627 & n81650;
  assign n81652 = ~n81648 & ~n81651;
  assign n81653 = ~n81627 & n81647;
  assign n81654 = ~n81627 & n81645;
  assign n81655 = n81621 & n81654;
  assign n81656 = ~n81615 & n81655;
  assign n81657 = ~n81653 & ~n81656;
  assign n81658 = n81609 & ~n81657;
  assign n81659 = n81621 & n81646;
  assign n81660 = n81645 & n81649;
  assign n81661 = ~n81627 & n81660;
  assign n81662 = ~n81659 & ~n81661;
  assign n81663 = ~n81609 & ~n81662;
  assign n81664 = ~n81658 & ~n81663;
  assign n81665 = n81652 & n81664;
  assign n81666 = n81639 & ~n81665;
  assign n81667 = ~n81621 & ~n81645;
  assign n81668 = n81609 & n81667;
  assign n81669 = ~n81615 & n81668;
  assign n81670 = n81627 & ~n81645;
  assign n81671 = n81621 & n81670;
  assign n81672 = n81615 & n81671;
  assign n81673 = ~n81648 & ~n81672;
  assign n81674 = ~n81627 & ~n81645;
  assign n81675 = ~n81621 & n81674;
  assign n81676 = n81673 & ~n81675;
  assign n81677 = n81609 & ~n81676;
  assign n81678 = ~n81669 & ~n81677;
  assign n81679 = ~n81609 & ~n81615;
  assign n81680 = n81646 & n81679;
  assign n81681 = n81621 & n81674;
  assign n81682 = n81615 & n81667;
  assign n81683 = n81627 & n81682;
  assign n81684 = ~n81681 & ~n81683;
  assign n81685 = n81615 & n81654;
  assign n81686 = n81684 & ~n81685;
  assign n81687 = ~n81609 & ~n81686;
  assign n81688 = ~n81621 & ~n81627;
  assign n81689 = n81609 & ~n81615;
  assign n81690 = n81688 & n81689;
  assign n81691 = ~n81615 & n81675;
  assign n81692 = ~n81690 & ~n81691;
  assign n81693 = ~n81687 & n81692;
  assign n81694 = ~n81680 & n81693;
  assign n81695 = ~n81615 & n81659;
  assign n81696 = n81615 & n81655;
  assign n81697 = ~n81695 & ~n81696;
  assign n81698 = n81694 & n81697;
  assign n81699 = ~n81639 & ~n81698;
  assign n81700 = n81678 & ~n81699;
  assign n81701 = ~n81666 & n81700;
  assign n81702 = ~n81633 & n81701;
  assign n81703 = ~pi2605 & ~n81702;
  assign n81704 = pi2605 & n81702;
  assign po2702 = n81703 | n81704;
  assign n81706 = ~n81615 & n81654;
  assign n81707 = ~n81615 & n81671;
  assign n81708 = ~n81706 & ~n81707;
  assign n81709 = n81609 & n81708;
  assign n81710 = n81615 & n81630;
  assign n81711 = ~n81646 & ~n81674;
  assign n81712 = n81621 & ~n81711;
  assign n81713 = n81627 & n81649;
  assign n81714 = n81615 & n81674;
  assign n81715 = ~n81713 & ~n81714;
  assign n81716 = ~n81609 & n81715;
  assign n81717 = ~n81712 & n81716;
  assign n81718 = ~n81710 & n81717;
  assign n81719 = ~n81709 & ~n81718;
  assign n81720 = n81615 & n81712;
  assign n81721 = ~n81621 & n81654;
  assign n81722 = n81615 & n81721;
  assign n81723 = ~n81720 & ~n81722;
  assign n81724 = ~n81719 & n81723;
  assign n81725 = n81639 & ~n81724;
  assign n81726 = n81609 & ~n81711;
  assign n81727 = ~n81615 & n81726;
  assign n81728 = ~n81655 & ~n81670;
  assign n81729 = n81615 & ~n81728;
  assign n81730 = n81609 & n81729;
  assign n81731 = ~n81621 & n81726;
  assign n81732 = ~n81730 & ~n81731;
  assign n81733 = ~n81727 & n81732;
  assign n81734 = ~n81639 & ~n81733;
  assign n81735 = ~n81725 & ~n81734;
  assign n81736 = n81609 & n81683;
  assign n81737 = ~n81609 & ~n81723;
  assign n81738 = ~n81736 & ~n81737;
  assign n81739 = ~n81609 & ~n81708;
  assign n81740 = ~n81683 & ~n81739;
  assign n81741 = ~n81639 & ~n81740;
  assign n81742 = n81738 & ~n81741;
  assign n81743 = n81735 & n81742;
  assign n81744 = pi2614 & ~n81743;
  assign n81745 = ~pi2614 & n81742;
  assign n81746 = ~n81734 & n81745;
  assign n81747 = ~n81725 & n81746;
  assign po2711 = n81744 | n81747;
  assign n81749 = ~n81628 & ~n81651;
  assign n81750 = n81609 & ~n81749;
  assign n81751 = n81615 & n81675;
  assign n81752 = ~n81750 & ~n81751;
  assign n81753 = ~n81661 & n81752;
  assign n81754 = ~n81609 & n81648;
  assign n81755 = ~n81695 & ~n81754;
  assign n81756 = ~n81672 & n81755;
  assign n81757 = n81753 & n81756;
  assign n81758 = n81639 & ~n81757;
  assign n81759 = ~n81683 & ~n81722;
  assign n81760 = ~n81691 & ~n81707;
  assign n81761 = n81621 & n81645;
  assign n81762 = n81615 & ~n81627;
  assign n81763 = ~n81761 & ~n81762;
  assign n81764 = ~n81667 & n81763;
  assign n81765 = ~n81609 & ~n81764;
  assign n81766 = ~n81621 & n81646;
  assign n81767 = n81609 & n81766;
  assign n81768 = n81615 & n81659;
  assign n81769 = ~n81767 & ~n81768;
  assign n81770 = ~n81765 & n81769;
  assign n81771 = n81760 & n81770;
  assign n81772 = n81759 & n81771;
  assign n81773 = ~n81639 & ~n81772;
  assign n81774 = ~n81758 & ~n81773;
  assign n81775 = pi2603 & ~n81774;
  assign n81776 = ~pi2603 & ~n81758;
  assign n81777 = ~n81773 & n81776;
  assign po2712 = n81775 | n81777;
  assign n81779 = ~n81533 & n81564;
  assign n81780 = n81533 & n81575;
  assign n81781 = ~n81561 & ~n81780;
  assign n81782 = n81507 & ~n81781;
  assign n81783 = ~n81779 & ~n81782;
  assign n81784 = ~n81507 & ~n81533;
  assign n81785 = ~n81525 & n81784;
  assign n81786 = ~n81519 & n81785;
  assign n81787 = n81549 & n81576;
  assign n81788 = ~n81786 & ~n81787;
  assign n81789 = ~n81507 & n81513;
  assign n81790 = n81535 & n81789;
  assign n81791 = n81788 & ~n81790;
  assign n81792 = ~n81537 & ~n81548;
  assign n81793 = n81525 & n81584;
  assign n81794 = n81792 & ~n81793;
  assign n81795 = n81791 & n81794;
  assign n81796 = n81783 & n81795;
  assign n81797 = ~n81573 & ~n81796;
  assign n81798 = ~n81536 & ~n81561;
  assign n81799 = n81533 & ~n81798;
  assign n81800 = ~n81519 & n81579;
  assign n81801 = ~n81590 & ~n81800;
  assign n81802 = n81513 & ~n81525;
  assign n81803 = n81533 & n81802;
  assign n81804 = n81801 & ~n81803;
  assign n81805 = n81507 & ~n81804;
  assign n81806 = ~n81533 & n81560;
  assign n81807 = n81527 & n81533;
  assign n81808 = ~n81806 & ~n81807;
  assign n81809 = ~n81507 & ~n81808;
  assign n81810 = ~n81533 & n81550;
  assign n81811 = ~n81809 & ~n81810;
  assign n81812 = ~n81805 & n81811;
  assign n81813 = ~n81799 & n81812;
  assign n81814 = n81573 & ~n81813;
  assign n81815 = n81507 & n81580;
  assign n81816 = ~n81814 & ~n81815;
  assign n81817 = n81555 & n81784;
  assign n81818 = ~n81525 & n81817;
  assign n81819 = n81816 & ~n81818;
  assign n81820 = ~n81797 & n81819;
  assign n81821 = ~pi2623 & ~n81820;
  assign n81822 = pi2623 & n81816;
  assign n81823 = ~n81797 & n81822;
  assign n81824 = ~n81818 & n81823;
  assign po2717 = n81821 | n81824;
  assign n81826 = ~n81534 & ~n81540;
  assign n81827 = ~n81507 & ~n81826;
  assign n81828 = ~n81597 & ~n81827;
  assign n81829 = ~n81513 & n81519;
  assign n81830 = n81507 & n81829;
  assign n81831 = n81533 & n81830;
  assign n81832 = n81533 & n81560;
  assign n81833 = ~n81829 & ~n81832;
  assign n81834 = n81513 & ~n81533;
  assign n81835 = ~n81519 & n81834;
  assign n81836 = n81833 & ~n81835;
  assign n81837 = n81507 & ~n81836;
  assign n81838 = ~n81543 & ~n81837;
  assign n81839 = ~n81573 & ~n81838;
  assign n81840 = ~n81507 & n81526;
  assign n81841 = n81533 & n81840;
  assign n81842 = ~n81790 & ~n81841;
  assign n81843 = ~n81573 & ~n81842;
  assign n81844 = ~n81839 & ~n81843;
  assign n81845 = ~n81831 & n81844;
  assign n81846 = ~n81561 & ~n81580;
  assign n81847 = ~n81590 & n81846;
  assign n81848 = ~n81507 & ~n81847;
  assign n81849 = ~n81533 & n81539;
  assign n81850 = ~n81564 & ~n81849;
  assign n81851 = n81507 & ~n81850;
  assign n81852 = ~n81848 & ~n81851;
  assign n81853 = ~n81800 & n81852;
  assign n81854 = ~n81548 & ~n81591;
  assign n81855 = n81853 & n81854;
  assign n81856 = n81573 & ~n81855;
  assign n81857 = n81845 & ~n81856;
  assign n81858 = n81828 & n81857;
  assign n81859 = ~pi2641 & ~n81858;
  assign n81860 = pi2641 & n81845;
  assign n81861 = n81828 & n81860;
  assign n81862 = ~n81856 & n81861;
  assign po2721 = n81859 | n81862;
  assign n81864 = ~n81615 & n81674;
  assign n81865 = ~n81721 & ~n81864;
  assign n81866 = n81609 & ~n81865;
  assign n81867 = ~n81672 & ~n81866;
  assign n81868 = n81615 & n81766;
  assign n81869 = ~n81696 & ~n81868;
  assign n81870 = ~n81682 & ~n81761;
  assign n81871 = ~n81621 & n81670;
  assign n81872 = n81870 & ~n81871;
  assign n81873 = ~n81609 & ~n81872;
  assign n81874 = ~n81615 & n81681;
  assign n81875 = ~n81873 & ~n81874;
  assign n81876 = n81869 & n81875;
  assign n81877 = n81867 & n81876;
  assign n81878 = ~n81639 & ~n81877;
  assign n81879 = ~n81656 & ~n81710;
  assign n81880 = ~n81609 & ~n81879;
  assign n81881 = ~n81878 & ~n81880;
  assign n81882 = n81609 & n81868;
  assign n81883 = n81649 & ~n81711;
  assign n81884 = ~n81671 & ~n81722;
  assign n81885 = ~n81883 & n81884;
  assign n81886 = ~n81609 & ~n81885;
  assign n81887 = n81615 & n81681;
  assign n81888 = ~n81886 & ~n81887;
  assign n81889 = ~n81615 & n81761;
  assign n81890 = ~n81871 & ~n81889;
  assign n81891 = ~n81714 & n81890;
  assign n81892 = n81609 & ~n81891;
  assign n81893 = n81888 & ~n81892;
  assign n81894 = n81639 & ~n81893;
  assign n81895 = ~n81882 & ~n81894;
  assign n81896 = n81881 & n81895;
  assign n81897 = pi2619 & n81896;
  assign n81898 = ~pi2619 & ~n81896;
  assign po2723 = n81897 | n81898;
  assign n81900 = pi5541 & pi9040;
  assign n81901 = pi5532 & ~pi9040;
  assign n81902 = ~n81900 & ~n81901;
  assign n81903 = ~pi2576 & ~n81902;
  assign n81904 = pi2576 & n81902;
  assign n81905 = ~n81903 & ~n81904;
  assign n81906 = pi5460 & ~pi9040;
  assign n81907 = pi5793 & pi9040;
  assign n81908 = ~n81906 & ~n81907;
  assign n81909 = ~pi2572 & ~n81908;
  assign n81910 = pi2572 & n81908;
  assign n81911 = ~n81909 & ~n81910;
  assign n81912 = pi5537 & ~pi9040;
  assign n81913 = pi5618 & pi9040;
  assign n81914 = ~n81912 & ~n81913;
  assign n81915 = pi2559 & n81914;
  assign n81916 = ~pi2559 & ~n81914;
  assign n81917 = ~n81915 & ~n81916;
  assign n81918 = pi5878 & pi9040;
  assign n81919 = pi5552 & ~pi9040;
  assign n81920 = ~n81918 & ~n81919;
  assign n81921 = ~pi2585 & ~n81920;
  assign n81922 = pi2585 & n81920;
  assign n81923 = ~n81921 & ~n81922;
  assign n81924 = pi5802 & ~pi9040;
  assign n81925 = pi5450 & pi9040;
  assign n81926 = ~n81924 & ~n81925;
  assign n81927 = ~pi2560 & n81926;
  assign n81928 = pi2560 & ~n81926;
  assign n81929 = ~n81927 & ~n81928;
  assign n81930 = n81923 & n81929;
  assign n81931 = n81917 & n81930;
  assign n81932 = pi5636 & pi9040;
  assign n81933 = pi5608 & ~pi9040;
  assign n81934 = ~n81932 & ~n81933;
  assign n81935 = ~pi2554 & n81934;
  assign n81936 = pi2554 & ~n81934;
  assign n81937 = ~n81935 & ~n81936;
  assign n81938 = ~n81929 & ~n81937;
  assign n81939 = n81923 & n81938;
  assign n81940 = ~n81931 & ~n81939;
  assign n81941 = ~n81929 & n81937;
  assign n81942 = ~n81923 & n81941;
  assign n81943 = ~n81917 & n81942;
  assign n81944 = n81940 & ~n81943;
  assign n81945 = n81911 & ~n81944;
  assign n81946 = ~n81923 & ~n81929;
  assign n81947 = ~n81937 & n81946;
  assign n81948 = ~n81917 & n81947;
  assign n81949 = n81929 & ~n81937;
  assign n81950 = n81923 & n81949;
  assign n81951 = ~n81917 & n81950;
  assign n81952 = ~n81923 & n81929;
  assign n81953 = ~n81941 & ~n81952;
  assign n81954 = n81917 & ~n81953;
  assign n81955 = ~n81951 & ~n81954;
  assign n81956 = ~n81948 & n81955;
  assign n81957 = ~n81911 & ~n81956;
  assign n81958 = ~n81945 & ~n81957;
  assign n81959 = n81905 & ~n81958;
  assign n81960 = n81911 & ~n81917;
  assign n81961 = n81929 & n81960;
  assign n81962 = ~n81911 & ~n81917;
  assign n81963 = n81941 & n81962;
  assign n81964 = ~n81917 & ~n81929;
  assign n81965 = n81923 & n81964;
  assign n81966 = ~n81931 & ~n81965;
  assign n81967 = ~n81911 & ~n81966;
  assign n81968 = ~n81963 & ~n81967;
  assign n81969 = n81923 & n81941;
  assign n81970 = ~n81917 & n81969;
  assign n81971 = n81917 & n81947;
  assign n81972 = ~n81970 & ~n81971;
  assign n81973 = n81911 & n81917;
  assign n81974 = n81946 & n81973;
  assign n81975 = ~n81923 & n81949;
  assign n81976 = n81911 & n81975;
  assign n81977 = ~n81974 & ~n81976;
  assign n81978 = n81972 & n81977;
  assign n81979 = n81968 & n81978;
  assign n81980 = ~n81961 & n81979;
  assign n81981 = ~n81905 & ~n81980;
  assign n81982 = n81929 & n81937;
  assign n81983 = ~n81923 & n81982;
  assign n81984 = ~n81911 & n81983;
  assign n81985 = ~n81917 & n81984;
  assign n81986 = ~n81911 & n81970;
  assign n81987 = ~n81985 & ~n81986;
  assign n81988 = ~n81917 & ~n81923;
  assign n81989 = ~n81937 & n81988;
  assign n81990 = n81929 & n81989;
  assign n81991 = n81911 & n81990;
  assign n81992 = n81987 & ~n81991;
  assign n81993 = ~n81917 & n81923;
  assign n81994 = n81937 & n81993;
  assign n81995 = n81929 & n81994;
  assign n81996 = n81917 & n81938;
  assign n81997 = ~n81995 & ~n81996;
  assign n81998 = n81911 & ~n81997;
  assign n81999 = n81992 & ~n81998;
  assign n82000 = ~n81981 & n81999;
  assign n82001 = ~n81959 & n82000;
  assign n82002 = pi2596 & n82001;
  assign n82003 = ~pi2596 & ~n82001;
  assign po2728 = n82002 | n82003;
  assign n82005 = pi5549 & pi9040;
  assign n82006 = pi5809 & ~pi9040;
  assign n82007 = ~n82005 & ~n82006;
  assign n82008 = ~pi2571 & ~n82007;
  assign n82009 = pi2571 & n82007;
  assign n82010 = ~n82008 & ~n82009;
  assign n82011 = pi5794 & ~pi9040;
  assign n82012 = pi5740 & pi9040;
  assign n82013 = ~n82011 & ~n82012;
  assign n82014 = ~pi2557 & ~n82013;
  assign n82015 = pi2557 & n82013;
  assign n82016 = ~n82014 & ~n82015;
  assign n82017 = pi5454 & ~pi9040;
  assign n82018 = pi5631 & pi9040;
  assign n82019 = ~n82017 & ~n82018;
  assign n82020 = pi2587 & n82019;
  assign n82021 = ~pi2587 & ~n82019;
  assign n82022 = ~n82020 & ~n82021;
  assign n82023 = n82016 & ~n82022;
  assign n82024 = pi5536 & ~pi9040;
  assign n82025 = pi5616 & pi9040;
  assign n82026 = ~n82024 & ~n82025;
  assign n82027 = ~pi2583 & ~n82026;
  assign n82028 = pi2583 & n82026;
  assign n82029 = ~n82027 & ~n82028;
  assign n82030 = pi5533 & ~pi9040;
  assign n82031 = pi5538 & pi9040;
  assign n82032 = ~n82030 & ~n82031;
  assign n82033 = ~pi2561 & n82032;
  assign n82034 = pi2561 & ~n82032;
  assign n82035 = ~n82033 & ~n82034;
  assign n82036 = n82029 & ~n82035;
  assign n82037 = n82023 & n82036;
  assign n82038 = n82016 & n82022;
  assign n82039 = n82035 & n82038;
  assign n82040 = ~n82016 & ~n82022;
  assign n82041 = n82035 & n82040;
  assign n82042 = ~n82039 & ~n82041;
  assign n82043 = n82029 & ~n82042;
  assign n82044 = ~n82037 & ~n82043;
  assign n82045 = ~n82010 & ~n82044;
  assign n82046 = ~n82029 & n82040;
  assign n82047 = ~n82016 & ~n82035;
  assign n82048 = n82022 & n82047;
  assign n82049 = ~n82046 & ~n82048;
  assign n82050 = pi5606 & pi9040;
  assign n82051 = pi5616 & ~pi9040;
  assign n82052 = ~n82050 & ~n82051;
  assign n82053 = pi2566 & n82052;
  assign n82054 = ~pi2566 & ~n82052;
  assign n82055 = ~n82053 & ~n82054;
  assign n82056 = ~n82010 & n82055;
  assign n82057 = ~n82049 & n82056;
  assign n82058 = ~n82045 & ~n82057;
  assign n82059 = n82029 & n82035;
  assign n82060 = ~n82016 & n82059;
  assign n82061 = ~n82037 & ~n82060;
  assign n82062 = ~n82055 & ~n82061;
  assign n82063 = ~n82029 & n82055;
  assign n82064 = n82016 & n82063;
  assign n82065 = n82023 & n82035;
  assign n82066 = ~n82035 & n82038;
  assign n82067 = ~n82065 & ~n82066;
  assign n82068 = ~n82035 & n82040;
  assign n82069 = n82029 & n82068;
  assign n82070 = n82067 & ~n82069;
  assign n82071 = n82055 & ~n82070;
  assign n82072 = ~n82064 & ~n82071;
  assign n82073 = ~n82016 & n82022;
  assign n82074 = n82035 & n82073;
  assign n82075 = n82029 & n82074;
  assign n82076 = n82072 & ~n82075;
  assign n82077 = ~n82049 & ~n82055;
  assign n82078 = ~n82029 & n82039;
  assign n82079 = ~n82077 & ~n82078;
  assign n82080 = n82076 & n82079;
  assign n82081 = n82010 & ~n82080;
  assign n82082 = ~n82062 & ~n82081;
  assign n82083 = ~n82010 & ~n82055;
  assign n82084 = n82023 & ~n82029;
  assign n82085 = ~n82074 & ~n82084;
  assign n82086 = n82016 & ~n82035;
  assign n82087 = n82085 & ~n82086;
  assign n82088 = n82083 & ~n82087;
  assign n82089 = n82082 & ~n82088;
  assign n82090 = n82058 & n82089;
  assign n82091 = ~pi2601 & ~n82090;
  assign n82092 = pi2601 & n82058;
  assign n82093 = n82082 & n82092;
  assign n82094 = ~n82088 & n82093;
  assign po2729 = n82091 | n82094;
  assign n82096 = pi5453 & ~pi9040;
  assign n82097 = pi5936 & pi9040;
  assign n82098 = ~n82096 & ~n82097;
  assign n82099 = ~pi2590 & ~n82098;
  assign n82100 = pi2590 & n82098;
  assign n82101 = ~n82099 & ~n82100;
  assign n82102 = pi5452 & pi9040;
  assign n82103 = pi5535 & ~pi9040;
  assign n82104 = ~n82102 & ~n82103;
  assign n82105 = ~pi2579 & n82104;
  assign n82106 = pi2579 & ~n82104;
  assign n82107 = ~n82105 & ~n82106;
  assign n82108 = pi5540 & pi9040;
  assign n82109 = pi5734 & ~pi9040;
  assign n82110 = ~n82108 & ~n82109;
  assign n82111 = ~pi2584 & n82110;
  assign n82112 = pi2584 & ~n82110;
  assign n82113 = ~n82111 & ~n82112;
  assign n82114 = pi5455 & ~pi9040;
  assign n82115 = pi5809 & pi9040;
  assign n82116 = ~n82114 & ~n82115;
  assign n82117 = ~pi2580 & n82116;
  assign n82118 = pi2580 & ~n82116;
  assign n82119 = ~n82117 & ~n82118;
  assign n82120 = pi5548 & ~pi9040;
  assign n82121 = pi5734 & pi9040;
  assign n82122 = ~n82120 & ~n82121;
  assign n82123 = ~pi2564 & ~n82122;
  assign n82124 = pi2564 & n82122;
  assign n82125 = ~n82123 & ~n82124;
  assign n82126 = n82119 & ~n82125;
  assign n82127 = n82113 & n82126;
  assign n82128 = n82107 & n82127;
  assign n82129 = ~pi2564 & n82122;
  assign n82130 = pi2564 & ~n82122;
  assign n82131 = ~n82129 & ~n82130;
  assign n82132 = n82119 & ~n82131;
  assign n82133 = n82113 & n82132;
  assign n82134 = ~n82107 & n82133;
  assign n82135 = ~n82128 & ~n82134;
  assign n82136 = n82101 & ~n82135;
  assign n82137 = n82107 & ~n82113;
  assign n82138 = ~n82119 & n82137;
  assign n82139 = ~n82125 & n82138;
  assign n82140 = ~n82101 & n82139;
  assign n82141 = pi5733 & ~pi9040;
  assign n82142 = pi5670 & pi9040;
  assign n82143 = ~n82141 & ~n82142;
  assign n82144 = ~pi2581 & ~n82143;
  assign n82145 = pi2581 & n82143;
  assign n82146 = ~n82144 & ~n82145;
  assign n82147 = ~n82113 & n82132;
  assign n82148 = n82101 & n82147;
  assign n82149 = ~n82139 & ~n82148;
  assign n82150 = n82107 & ~n82131;
  assign n82151 = n82113 & n82150;
  assign n82152 = ~n82125 & n82137;
  assign n82153 = ~n82151 & ~n82152;
  assign n82154 = ~n82101 & ~n82153;
  assign n82155 = ~n82101 & ~n82107;
  assign n82156 = n82126 & n82155;
  assign n82157 = n82113 & n82156;
  assign n82158 = ~n82107 & ~n82113;
  assign n82159 = ~n82119 & n82158;
  assign n82160 = ~n82131 & n82159;
  assign n82161 = n82101 & n82113;
  assign n82162 = ~n82119 & n82161;
  assign n82163 = ~n82125 & n82162;
  assign n82164 = ~n82160 & ~n82163;
  assign n82165 = ~n82157 & n82164;
  assign n82166 = ~n82154 & n82165;
  assign n82167 = n82149 & n82166;
  assign n82168 = n82146 & ~n82167;
  assign n82169 = n82107 & n82148;
  assign n82170 = ~n82168 & ~n82169;
  assign n82171 = ~n82140 & n82170;
  assign n82172 = ~n82136 & n82171;
  assign n82173 = n82101 & ~n82107;
  assign n82174 = ~n82113 & ~n82125;
  assign n82175 = n82173 & n82174;
  assign n82176 = n82101 & n82127;
  assign n82177 = ~n82175 & ~n82176;
  assign n82178 = ~n82119 & ~n82131;
  assign n82179 = ~n82113 & n82178;
  assign n82180 = n82101 & n82179;
  assign n82181 = n82113 & n82178;
  assign n82182 = n82107 & n82181;
  assign n82183 = ~n82180 & ~n82182;
  assign n82184 = ~n82113 & n82126;
  assign n82185 = ~n82107 & n82184;
  assign n82186 = ~n82128 & ~n82185;
  assign n82187 = ~n82107 & n82132;
  assign n82188 = n82113 & ~n82119;
  assign n82189 = ~n82187 & ~n82188;
  assign n82190 = ~n82101 & ~n82189;
  assign n82191 = n82186 & ~n82190;
  assign n82192 = n82183 & n82191;
  assign n82193 = n82177 & n82192;
  assign n82194 = ~n82146 & ~n82193;
  assign n82195 = n82172 & ~n82194;
  assign n82196 = ~pi2592 & ~n82195;
  assign n82197 = pi2592 & n82172;
  assign n82198 = ~n82194 & n82197;
  assign po2734 = n82196 | n82198;
  assign n82200 = ~n82107 & n82147;
  assign n82201 = n82107 & n82184;
  assign n82202 = ~n82200 & ~n82201;
  assign n82203 = ~n82119 & ~n82125;
  assign n82204 = ~n82113 & n82203;
  assign n82205 = ~n82107 & n82204;
  assign n82206 = ~n82107 & n82178;
  assign n82207 = n82113 & n82203;
  assign n82208 = n82107 & n82207;
  assign n82209 = ~n82206 & ~n82208;
  assign n82210 = ~n82101 & ~n82209;
  assign n82211 = ~n82205 & ~n82210;
  assign n82212 = n82101 & n82203;
  assign n82213 = ~n82107 & n82212;
  assign n82214 = ~n82176 & ~n82213;
  assign n82215 = n82211 & n82214;
  assign n82216 = n82202 & n82215;
  assign n82217 = n82146 & ~n82216;
  assign n82218 = ~n82101 & ~n82146;
  assign n82219 = ~n82107 & n82113;
  assign n82220 = n82131 & n82219;
  assign n82221 = n82113 & n82119;
  assign n82222 = ~n82220 & ~n82221;
  assign n82223 = n82218 & ~n82222;
  assign n82224 = ~n82139 & ~n82151;
  assign n82225 = ~n82113 & n82173;
  assign n82226 = ~n82203 & n82225;
  assign n82227 = ~n82148 & ~n82226;
  assign n82228 = n82224 & n82227;
  assign n82229 = ~n82146 & ~n82228;
  assign n82230 = ~n82101 & n82133;
  assign n82231 = n82107 & n82230;
  assign n82232 = n82107 & n82179;
  assign n82233 = ~n82201 & ~n82232;
  assign n82234 = ~n82101 & ~n82233;
  assign n82235 = ~n82231 & ~n82234;
  assign n82236 = n82101 & n82139;
  assign n82237 = n82235 & ~n82236;
  assign n82238 = ~n82229 & n82237;
  assign n82239 = ~n82223 & n82238;
  assign n82240 = ~n82217 & n82239;
  assign n82241 = n82101 & n82107;
  assign n82242 = n82181 & n82241;
  assign n82243 = n82240 & ~n82242;
  assign n82244 = ~pi2593 & ~n82243;
  assign n82245 = pi2593 & ~n82242;
  assign n82246 = n82239 & n82245;
  assign n82247 = ~n82217 & n82246;
  assign po2735 = n82244 | n82247;
  assign n82249 = n82029 & ~n82055;
  assign n82250 = ~n82039 & ~n82040;
  assign n82251 = n82249 & ~n82250;
  assign n82252 = n82035 & ~n82055;
  assign n82253 = n82040 & n82252;
  assign n82254 = ~n82251 & ~n82253;
  assign n82255 = n82010 & ~n82254;
  assign n82256 = ~n82029 & n82066;
  assign n82257 = ~n82029 & ~n82035;
  assign n82258 = ~n82086 & ~n82257;
  assign n82259 = n82055 & ~n82258;
  assign n82260 = ~n82029 & n82035;
  assign n82261 = ~n82022 & n82260;
  assign n82262 = n82016 & n82261;
  assign n82263 = ~n82259 & ~n82262;
  assign n82264 = ~n82256 & n82263;
  assign n82265 = n82010 & ~n82264;
  assign n82266 = ~n82255 & ~n82265;
  assign n82267 = n82029 & n82048;
  assign n82268 = ~n82029 & n82074;
  assign n82269 = ~n82267 & ~n82268;
  assign n82270 = ~n82055 & ~n82269;
  assign n82271 = n82029 & n82041;
  assign n82272 = ~n82029 & n82086;
  assign n82273 = ~n82271 & ~n82272;
  assign n82274 = n82055 & ~n82273;
  assign n82275 = ~n82023 & ~n82086;
  assign n82276 = n82029 & ~n82275;
  assign n82277 = ~n82074 & ~n82276;
  assign n82278 = ~n82055 & ~n82277;
  assign n82279 = n82022 & ~n82029;
  assign n82280 = n82252 & n82279;
  assign n82281 = ~n82022 & ~n82035;
  assign n82282 = ~n82074 & ~n82281;
  assign n82283 = ~n82029 & ~n82282;
  assign n82284 = n82029 & n82055;
  assign n82285 = n82038 & n82284;
  assign n82286 = n82035 & n82285;
  assign n82287 = ~n82283 & ~n82286;
  assign n82288 = ~n82280 & n82287;
  assign n82289 = ~n82278 & n82288;
  assign n82290 = ~n82267 & n82289;
  assign n82291 = ~n82010 & ~n82290;
  assign n82292 = ~n82274 & ~n82291;
  assign n82293 = ~n82270 & n82292;
  assign n82294 = n82266 & n82293;
  assign n82295 = pi2607 & n82294;
  assign n82296 = ~pi2607 & ~n82294;
  assign po2736 = n82295 | n82296;
  assign n82298 = ~n81591 & ~n81810;
  assign n82299 = n81507 & ~n82298;
  assign n82300 = ~n81573 & n81575;
  assign n82301 = ~n81507 & n82300;
  assign n82302 = n81519 & n81834;
  assign n82303 = ~n81802 & ~n82302;
  assign n82304 = ~n81550 & n82303;
  assign n82305 = n81507 & ~n82304;
  assign n82306 = ~n81513 & n81560;
  assign n82307 = ~n81533 & n82306;
  assign n82308 = ~n82305 & ~n82307;
  assign n82309 = ~n81573 & ~n82308;
  assign n82310 = ~n82301 & ~n82309;
  assign n82311 = ~n81537 & ~n81540;
  assign n82312 = ~n81533 & n81590;
  assign n82313 = ~n81780 & ~n82312;
  assign n82314 = n82311 & n82313;
  assign n82315 = ~n81507 & ~n82314;
  assign n82316 = ~n81513 & ~n81519;
  assign n82317 = ~n81507 & n82316;
  assign n82318 = n81533 & n82317;
  assign n82319 = ~n81533 & n81802;
  assign n82320 = ~n81540 & ~n82319;
  assign n82321 = ~n81807 & n82320;
  assign n82322 = ~n82318 & n82321;
  assign n82323 = n81507 & n81536;
  assign n82324 = n82322 & ~n82323;
  assign n82325 = n81573 & ~n82324;
  assign n82326 = ~n82315 & ~n82325;
  assign n82327 = n82310 & n82326;
  assign n82328 = ~n82299 & n82327;
  assign n82329 = pi2652 & n82328;
  assign n82330 = ~pi2652 & ~n82328;
  assign po2737 = n82329 | n82330;
  assign n82332 = ~n81905 & ~n81911;
  assign n82333 = ~n81917 & n81930;
  assign n82334 = n81917 & n81969;
  assign n82335 = ~n81917 & n81938;
  assign n82336 = ~n82334 & ~n82335;
  assign n82337 = ~n82333 & n82336;
  assign n82338 = n82332 & ~n82337;
  assign n82339 = n81937 & n81988;
  assign n82340 = n81923 & n81982;
  assign n82341 = n81917 & n82340;
  assign n82342 = ~n82339 & ~n82341;
  assign n82343 = ~n81939 & ~n81942;
  assign n82344 = n82342 & n82343;
  assign n82345 = n81911 & ~n82344;
  assign n82346 = n81917 & n81975;
  assign n82347 = ~n82345 & ~n82346;
  assign n82348 = ~n81905 & ~n82347;
  assign n82349 = ~n82338 & ~n82348;
  assign n82350 = n81923 & n81960;
  assign n82351 = ~n81937 & n82350;
  assign n82352 = ~n81943 & ~n82351;
  assign n82353 = ~n81938 & ~n81982;
  assign n82354 = n81917 & ~n82353;
  assign n82355 = ~n81983 & ~n82354;
  assign n82356 = ~n81911 & ~n82355;
  assign n82357 = ~n81950 & ~n82333;
  assign n82358 = ~n82334 & n82357;
  assign n82359 = n81911 & ~n82358;
  assign n82360 = ~n82356 & ~n82359;
  assign n82361 = n81917 & ~n81923;
  assign n82362 = n81937 & n82361;
  assign n82363 = n81929 & n82362;
  assign n82364 = ~n81971 & ~n82363;
  assign n82365 = ~n81990 & n82364;
  assign n82366 = ~n81963 & n82365;
  assign n82367 = n82360 & n82366;
  assign n82368 = n81905 & ~n82367;
  assign n82369 = n82352 & ~n82368;
  assign n82370 = n82349 & n82369;
  assign n82371 = pi2600 & ~n82370;
  assign n82372 = ~pi2600 & n82352;
  assign n82373 = n82349 & n82372;
  assign n82374 = ~n82368 & n82373;
  assign po2738 = n82371 | n82374;
  assign n82376 = ~n81950 & ~n81983;
  assign n82377 = ~n81911 & ~n82376;
  assign n82378 = n81917 & n81939;
  assign n82379 = ~n82377 & ~n82378;
  assign n82380 = n81917 & ~n81929;
  assign n82381 = ~n81946 & ~n82380;
  assign n82382 = ~n82340 & n82381;
  assign n82383 = n81911 & ~n82382;
  assign n82384 = n82379 & ~n82383;
  assign n82385 = ~n81905 & ~n82384;
  assign n82386 = ~n81911 & n81948;
  assign n82387 = ~n81986 & ~n82386;
  assign n82388 = ~n81991 & n82387;
  assign n82389 = ~n81976 & ~n81994;
  assign n82390 = n81911 & n81965;
  assign n82391 = n82389 & ~n82390;
  assign n82392 = n81917 & n81950;
  assign n82393 = ~n81911 & n81946;
  assign n82394 = ~n82392 & ~n82393;
  assign n82395 = ~n82363 & n82394;
  assign n82396 = n82391 & n82395;
  assign n82397 = ~n81990 & n82396;
  assign n82398 = n81905 & ~n82397;
  assign n82399 = n82388 & ~n82398;
  assign n82400 = ~n82385 & n82399;
  assign n82401 = ~pi2609 & ~n82400;
  assign n82402 = pi2609 & n82388;
  assign n82403 = ~n82385 & n82402;
  assign n82404 = ~n82398 & n82403;
  assign po2740 = n82401 | n82404;
  assign n82406 = ~n82169 & ~n82175;
  assign n82407 = ~n82133 & ~n82139;
  assign n82408 = ~n82187 & n82407;
  assign n82409 = ~n82101 & ~n82408;
  assign n82410 = ~n82107 & n82207;
  assign n82411 = ~n82160 & ~n82410;
  assign n82412 = ~n82242 & n82411;
  assign n82413 = n82101 & n82184;
  assign n82414 = n82412 & ~n82413;
  assign n82415 = ~n82409 & n82414;
  assign n82416 = n82146 & ~n82415;
  assign n82417 = n82107 & n82212;
  assign n82418 = n82125 & n82219;
  assign n82419 = ~n82133 & ~n82418;
  assign n82420 = n82101 & ~n82419;
  assign n82421 = ~n82417 & ~n82420;
  assign n82422 = ~n82101 & n82178;
  assign n82423 = n82107 & n82422;
  assign n82424 = ~n82101 & n82127;
  assign n82425 = ~n82423 & ~n82424;
  assign n82426 = n82421 & n82425;
  assign n82427 = n82125 & n82137;
  assign n82428 = ~n82128 & ~n82427;
  assign n82429 = ~n82185 & n82428;
  assign n82430 = n82426 & n82429;
  assign n82431 = ~n82146 & ~n82430;
  assign n82432 = ~n82128 & n82411;
  assign n82433 = ~n82101 & ~n82432;
  assign n82434 = ~n82431 & ~n82433;
  assign n82435 = ~n82416 & n82434;
  assign n82436 = n82406 & n82435;
  assign n82437 = pi2594 & ~n82436;
  assign n82438 = ~pi2594 & n82436;
  assign po2741 = n82437 | n82438;
  assign n82440 = pi5453 & pi9040;
  assign n82441 = pi5631 & ~pi9040;
  assign n82442 = ~n82440 & ~n82441;
  assign n82443 = ~pi2557 & ~n82442;
  assign n82444 = pi2557 & n82442;
  assign n82445 = ~n82443 & ~n82444;
  assign n82446 = pi5808 & ~pi9040;
  assign n82447 = pi5624 & pi9040;
  assign n82448 = ~n82446 & ~n82447;
  assign n82449 = ~pi2570 & ~n82448;
  assign n82450 = pi2570 & n82448;
  assign n82451 = ~n82449 & ~n82450;
  assign n82452 = pi5722 & pi9040;
  assign n82453 = pi5609 & ~pi9040;
  assign n82454 = ~n82452 & ~n82453;
  assign n82455 = ~pi2575 & ~n82454;
  assign n82456 = pi2575 & n82454;
  assign n82457 = ~n82455 & ~n82456;
  assign n82458 = pi5722 & ~pi9040;
  assign n82459 = pi5539 & pi9040;
  assign n82460 = ~n82458 & ~n82459;
  assign n82461 = ~pi2561 & n82460;
  assign n82462 = pi2561 & ~n82460;
  assign n82463 = ~n82461 & ~n82462;
  assign n82464 = ~n82457 & ~n82463;
  assign n82465 = pi5455 & pi9040;
  assign n82466 = pi5936 & ~pi9040;
  assign n82467 = ~n82465 & ~n82466;
  assign n82468 = ~pi2582 & ~n82467;
  assign n82469 = pi2582 & n82467;
  assign n82470 = ~n82468 & ~n82469;
  assign n82471 = pi5539 & ~pi9040;
  assign n82472 = pi5536 & pi9040;
  assign n82473 = ~n82471 & ~n82472;
  assign n82474 = pi2586 & n82473;
  assign n82475 = ~pi2586 & ~n82473;
  assign n82476 = ~n82474 & ~n82475;
  assign n82477 = n82470 & n82476;
  assign n82478 = n82464 & n82477;
  assign n82479 = n82451 & n82478;
  assign n82480 = ~n82470 & n82476;
  assign n82481 = n82457 & ~n82463;
  assign n82482 = n82480 & n82481;
  assign n82483 = n82451 & ~n82470;
  assign n82484 = n82463 & n82483;
  assign n82485 = ~n82457 & n82484;
  assign n82486 = n82457 & n82463;
  assign n82487 = n82451 & n82486;
  assign n82488 = n82476 & n82487;
  assign n82489 = n82470 & n82488;
  assign n82490 = ~n82485 & ~n82489;
  assign n82491 = ~n82482 & n82490;
  assign n82492 = ~n82479 & n82491;
  assign n82493 = ~n82451 & ~n82470;
  assign n82494 = ~n82463 & n82493;
  assign n82495 = n82457 & n82494;
  assign n82496 = n82492 & ~n82495;
  assign n82497 = ~n82445 & ~n82496;
  assign n82498 = n82451 & n82457;
  assign n82499 = ~n82463 & n82498;
  assign n82500 = n82470 & n82499;
  assign n82501 = ~n82484 & ~n82500;
  assign n82502 = ~n82451 & n82464;
  assign n82503 = n82470 & n82502;
  assign n82504 = n82501 & ~n82503;
  assign n82505 = ~n82476 & ~n82504;
  assign n82506 = ~n82451 & n82463;
  assign n82507 = n82457 & n82506;
  assign n82508 = ~n82476 & n82507;
  assign n82509 = n82470 & n82508;
  assign n82510 = ~n82457 & n82483;
  assign n82511 = ~n82457 & n82463;
  assign n82512 = ~n82470 & n82511;
  assign n82513 = ~n82510 & ~n82512;
  assign n82514 = ~n82476 & ~n82513;
  assign n82515 = ~n82509 & ~n82514;
  assign n82516 = ~n82445 & ~n82515;
  assign n82517 = ~n82505 & ~n82516;
  assign n82518 = ~n82497 & n82517;
  assign n82519 = ~n82451 & n82470;
  assign n82520 = n82476 & n82519;
  assign n82521 = n82511 & n82520;
  assign n82522 = ~n82451 & n82480;
  assign n82523 = n82457 & n82522;
  assign n82524 = ~n82470 & n82507;
  assign n82525 = n82451 & ~n82476;
  assign n82526 = n82457 & n82525;
  assign n82527 = ~n82457 & n82470;
  assign n82528 = ~n82451 & n82527;
  assign n82529 = ~n82526 & ~n82528;
  assign n82530 = ~n82524 & n82529;
  assign n82531 = ~n82502 & n82530;
  assign n82532 = n82464 & n82476;
  assign n82533 = ~n82470 & n82532;
  assign n82534 = n82470 & n82511;
  assign n82535 = ~n82451 & ~n82463;
  assign n82536 = ~n82534 & ~n82535;
  assign n82537 = n82476 & ~n82536;
  assign n82538 = ~n82533 & ~n82537;
  assign n82539 = n82531 & n82538;
  assign n82540 = n82445 & ~n82539;
  assign n82541 = ~n82523 & ~n82540;
  assign n82542 = ~n82521 & n82541;
  assign n82543 = n82518 & n82542;
  assign n82544 = pi2597 & n82543;
  assign n82545 = ~pi2597 & ~n82543;
  assign po2742 = n82544 | n82545;
  assign n82547 = pi5742 & pi9040;
  assign n82548 = pi5464 & ~pi9040;
  assign n82549 = ~n82547 & ~n82548;
  assign n82550 = pi2560 & n82549;
  assign n82551 = ~pi2560 & ~n82549;
  assign n82552 = ~n82550 & ~n82551;
  assign n82553 = pi5878 & ~pi9040;
  assign n82554 = pi5530 & pi9040;
  assign n82555 = ~n82553 & ~n82554;
  assign n82556 = pi2591 & n82555;
  assign n82557 = ~pi2591 & ~n82555;
  assign n82558 = ~n82556 & ~n82557;
  assign n82559 = pi5562 & ~pi9040;
  assign n82560 = pi5633 & pi9040;
  assign n82561 = ~n82559 & ~n82560;
  assign n82562 = pi2548 & n82561;
  assign n82563 = ~pi2548 & ~n82561;
  assign n82564 = ~n82562 & ~n82563;
  assign n82565 = ~n82558 & ~n82564;
  assign n82566 = pi5619 & pi9040;
  assign n82567 = pi5459 & ~pi9040;
  assign n82568 = ~n82566 & ~n82567;
  assign n82569 = ~pi2581 & ~n82568;
  assign n82570 = pi2581 & n82568;
  assign n82571 = ~n82569 & ~n82570;
  assign n82572 = n82565 & n82571;
  assign n82573 = pi5541 & ~pi9040;
  assign n82574 = pi5687 & pi9040;
  assign n82575 = ~n82573 & ~n82574;
  assign n82576 = pi2580 & n82575;
  assign n82577 = ~pi2580 & ~n82575;
  assign n82578 = ~n82576 & ~n82577;
  assign n82579 = pi5634 & ~pi9040;
  assign n82580 = pi5626 & pi9040;
  assign n82581 = ~n82579 & ~n82580;
  assign n82582 = pi2585 & n82581;
  assign n82583 = ~pi2585 & ~n82581;
  assign n82584 = ~n82582 & ~n82583;
  assign n82585 = ~n82571 & ~n82584;
  assign n82586 = n82578 & n82585;
  assign n82587 = n82558 & n82586;
  assign n82588 = ~n82571 & n82584;
  assign n82589 = ~n82578 & n82588;
  assign n82590 = n82558 & n82589;
  assign n82591 = ~n82587 & ~n82590;
  assign n82592 = n82571 & n82584;
  assign n82593 = ~n82578 & n82592;
  assign n82594 = ~n82558 & ~n82578;
  assign n82595 = ~n82584 & n82594;
  assign n82596 = ~n82571 & n82595;
  assign n82597 = ~n82593 & ~n82596;
  assign n82598 = n82564 & ~n82597;
  assign n82599 = n82591 & ~n82598;
  assign n82600 = ~n82572 & n82599;
  assign n82601 = n82552 & ~n82600;
  assign n82602 = n82571 & ~n82584;
  assign n82603 = ~n82578 & n82602;
  assign n82604 = n82558 & n82603;
  assign n82605 = ~n82564 & n82604;
  assign n82606 = ~n82558 & n82564;
  assign n82607 = n82603 & n82606;
  assign n82608 = ~n82558 & n82578;
  assign n82609 = ~n82571 & n82608;
  assign n82610 = ~n82607 & ~n82609;
  assign n82611 = n82578 & ~n82584;
  assign n82612 = n82571 & n82611;
  assign n82613 = n82558 & n82612;
  assign n82614 = ~n82578 & n82585;
  assign n82615 = n82558 & n82614;
  assign n82616 = ~n82613 & ~n82615;
  assign n82617 = n82578 & n82588;
  assign n82618 = ~n82593 & ~n82617;
  assign n82619 = ~n82558 & n82588;
  assign n82620 = n82618 & ~n82619;
  assign n82621 = ~n82564 & ~n82620;
  assign n82622 = n82578 & n82592;
  assign n82623 = n82564 & n82622;
  assign n82624 = ~n82621 & ~n82623;
  assign n82625 = n82616 & n82624;
  assign n82626 = n82610 & n82625;
  assign n82627 = ~n82552 & ~n82626;
  assign n82628 = ~n82605 & ~n82627;
  assign n82629 = ~n82601 & n82628;
  assign n82630 = n82606 & n82617;
  assign n82631 = n82564 & n82611;
  assign n82632 = n82558 & n82631;
  assign n82633 = ~n82630 & ~n82632;
  assign n82634 = n82564 & n82590;
  assign n82635 = n82633 & ~n82634;
  assign n82636 = n82629 & n82635;
  assign n82637 = ~pi2604 & ~n82636;
  assign n82638 = pi2604 & n82635;
  assign n82639 = n82628 & n82638;
  assign n82640 = ~n82601 & n82639;
  assign po2743 = n82637 | n82640;
  assign n82642 = ~n82022 & n82059;
  assign n82643 = ~n82039 & ~n82642;
  assign n82644 = ~n82055 & ~n82643;
  assign n82645 = n82029 & n82073;
  assign n82646 = ~n82261 & ~n82645;
  assign n82647 = n82055 & ~n82646;
  assign n82648 = ~n82029 & n82068;
  assign n82649 = ~n82280 & ~n82648;
  assign n82650 = ~n82037 & n82649;
  assign n82651 = ~n82647 & n82650;
  assign n82652 = ~n82644 & n82651;
  assign n82653 = ~n82256 & ~n82267;
  assign n82654 = n82652 & n82653;
  assign n82655 = n82010 & ~n82654;
  assign n82656 = n82016 & n82059;
  assign n82657 = n82029 & n82038;
  assign n82658 = ~n82656 & ~n82657;
  assign n82659 = n82055 & ~n82658;
  assign n82660 = n82055 & n82073;
  assign n82661 = ~n82029 & n82660;
  assign n82662 = ~n82659 & ~n82661;
  assign n82663 = n82023 & n82257;
  assign n82664 = n82042 & ~n82663;
  assign n82665 = n82055 & ~n82664;
  assign n82666 = ~n82029 & n82048;
  assign n82667 = ~n82665 & ~n82666;
  assign n82668 = n82662 & n82667;
  assign n82669 = ~n82010 & ~n82668;
  assign n82670 = ~n82068 & ~n82075;
  assign n82671 = ~n82262 & n82670;
  assign n82672 = n82083 & ~n82671;
  assign n82673 = ~n82669 & ~n82672;
  assign n82674 = ~n82037 & ~n82256;
  assign n82675 = ~n82055 & ~n82674;
  assign n82676 = n82673 & ~n82675;
  assign n82677 = ~n82655 & n82676;
  assign n82678 = ~pi2615 & n82677;
  assign n82679 = pi2615 & ~n82677;
  assign po2744 = n82678 | n82679;
  assign n82681 = pi5454 & pi9040;
  assign n82682 = pi5538 & ~pi9040;
  assign n82683 = ~n82681 & ~n82682;
  assign n82684 = ~pi2587 & ~n82683;
  assign n82685 = pi2587 & n82683;
  assign n82686 = ~n82684 & ~n82685;
  assign n82687 = pi5624 & ~pi9040;
  assign n82688 = pi5535 & pi9040;
  assign n82689 = ~n82687 & ~n82688;
  assign n82690 = ~pi2584 & ~n82689;
  assign n82691 = pi2584 & n82689;
  assign n82692 = ~n82690 & ~n82691;
  assign n82693 = pi5668 & ~pi9040;
  assign n82694 = pi5609 & pi9040;
  assign n82695 = ~n82693 & ~n82694;
  assign n82696 = ~pi2571 & ~n82695;
  assign n82697 = pi2571 & n82695;
  assign n82698 = ~n82696 & ~n82697;
  assign n82699 = ~n82692 & n82698;
  assign n82700 = ~n82686 & n82699;
  assign n82701 = n82692 & n82698;
  assign n82702 = n82686 & n82701;
  assign n82703 = ~n82700 & ~n82702;
  assign n82704 = pi5794 & pi9040;
  assign n82705 = pi5549 & ~pi9040;
  assign n82706 = ~n82704 & ~n82705;
  assign n82707 = ~pi2565 & n82706;
  assign n82708 = pi2565 & ~n82706;
  assign n82709 = ~n82707 & ~n82708;
  assign n82710 = n82686 & n82709;
  assign n82711 = n82692 & n82710;
  assign n82712 = n82703 & ~n82711;
  assign n82713 = pi5670 & ~pi9040;
  assign n82714 = pi5668 & pi9040;
  assign n82715 = ~n82713 & ~n82714;
  assign n82716 = ~pi2558 & ~n82715;
  assign n82717 = pi2558 & n82715;
  assign n82718 = ~n82716 & ~n82717;
  assign n82719 = pi5540 & ~pi9040;
  assign n82720 = pi5808 & pi9040;
  assign n82721 = ~n82719 & ~n82720;
  assign n82722 = ~pi2564 & ~n82721;
  assign n82723 = pi2564 & n82721;
  assign n82724 = ~n82722 & ~n82723;
  assign n82725 = ~n82718 & n82724;
  assign n82726 = ~n82712 & n82725;
  assign n82727 = ~n82692 & ~n82698;
  assign n82728 = n82686 & n82727;
  assign n82729 = ~n82709 & n82724;
  assign n82730 = n82728 & n82729;
  assign n82731 = n82686 & n82699;
  assign n82732 = n82718 & n82731;
  assign n82733 = n82692 & ~n82698;
  assign n82734 = ~n82709 & n82733;
  assign n82735 = ~n82686 & n82692;
  assign n82736 = ~n82734 & ~n82735;
  assign n82737 = n82718 & ~n82736;
  assign n82738 = ~n82732 & ~n82737;
  assign n82739 = n82724 & ~n82738;
  assign n82740 = ~n82730 & ~n82739;
  assign n82741 = ~n82686 & n82709;
  assign n82742 = ~n82698 & n82741;
  assign n82743 = ~n82692 & n82742;
  assign n82744 = ~n82686 & ~n82709;
  assign n82745 = n82692 & n82744;
  assign n82746 = ~n82743 & ~n82745;
  assign n82747 = n82718 & ~n82746;
  assign n82748 = n82740 & ~n82747;
  assign n82749 = ~n82709 & ~n82718;
  assign n82750 = n82733 & n82749;
  assign n82751 = n82686 & n82750;
  assign n82752 = ~n82701 & ~n82727;
  assign n82753 = n82710 & ~n82752;
  assign n82754 = n82698 & n82741;
  assign n82755 = ~n82692 & n82754;
  assign n82756 = ~n82753 & ~n82755;
  assign n82757 = n82744 & ~n82752;
  assign n82758 = ~n82709 & n82731;
  assign n82759 = ~n82757 & ~n82758;
  assign n82760 = ~n82686 & n82733;
  assign n82761 = n82709 & ~n82718;
  assign n82762 = n82760 & n82761;
  assign n82763 = n82759 & ~n82762;
  assign n82764 = n82756 & n82763;
  assign n82765 = ~n82751 & n82764;
  assign n82766 = n82709 & n82718;
  assign n82767 = n82686 & n82766;
  assign n82768 = ~n82698 & n82767;
  assign n82769 = n82765 & ~n82768;
  assign n82770 = ~n82724 & ~n82769;
  assign n82771 = n82748 & ~n82770;
  assign n82772 = ~n82726 & n82771;
  assign n82773 = ~pi2618 & ~n82772;
  assign n82774 = pi2618 & n82748;
  assign n82775 = ~n82726 & n82774;
  assign n82776 = ~n82770 & n82775;
  assign po2745 = n82773 | n82776;
  assign n82778 = n82686 & n82733;
  assign n82779 = n82718 & n82778;
  assign n82780 = n82709 & n82779;
  assign n82781 = n82699 & n82766;
  assign n82782 = ~n82686 & n82781;
  assign n82783 = ~n82780 & ~n82782;
  assign n82784 = ~n82755 & ~n82762;
  assign n82785 = n82686 & n82698;
  assign n82786 = ~n82709 & n82785;
  assign n82787 = ~n82734 & ~n82786;
  assign n82788 = n82718 & ~n82787;
  assign n82789 = ~n82718 & ~n82741;
  assign n82790 = ~n82752 & n82789;
  assign n82791 = n82709 & ~n82733;
  assign n82792 = n82718 & n82791;
  assign n82793 = ~n82686 & n82792;
  assign n82794 = ~n82790 & ~n82793;
  assign n82795 = ~n82788 & n82794;
  assign n82796 = n82784 & n82795;
  assign n82797 = n82724 & ~n82796;
  assign n82798 = n82783 & ~n82797;
  assign n82799 = n82702 & ~n82718;
  assign n82800 = ~n82709 & n82799;
  assign n82801 = ~n82718 & ~n82724;
  assign n82802 = ~n82731 & ~n82734;
  assign n82803 = n82741 & ~n82752;
  assign n82804 = n82802 & ~n82803;
  assign n82805 = n82801 & ~n82804;
  assign n82806 = n82700 & ~n82709;
  assign n82807 = n82698 & ~n82709;
  assign n82808 = ~n82686 & n82807;
  assign n82809 = ~n82709 & n82727;
  assign n82810 = ~n82808 & ~n82809;
  assign n82811 = n82709 & n82733;
  assign n82812 = ~n82728 & ~n82811;
  assign n82813 = n82810 & n82812;
  assign n82814 = n82718 & ~n82813;
  assign n82815 = ~n82806 & ~n82814;
  assign n82816 = ~n82724 & ~n82815;
  assign n82817 = ~n82805 & ~n82816;
  assign n82818 = ~n82800 & n82817;
  assign n82819 = n82798 & n82818;
  assign n82820 = pi2620 & ~n82819;
  assign n82821 = ~pi2620 & n82798;
  assign n82822 = n82818 & n82821;
  assign po2746 = n82820 | n82822;
  assign n82824 = n81911 & n81938;
  assign n82825 = ~n81917 & n82824;
  assign n82826 = ~n81995 & ~n82825;
  assign n82827 = n81917 & ~n81937;
  assign n82828 = n81923 & n82827;
  assign n82829 = ~n81917 & n81929;
  assign n82830 = ~n81994 & ~n82829;
  assign n82831 = ~n81911 & ~n82830;
  assign n82832 = ~n82828 & ~n82831;
  assign n82833 = n82826 & n82832;
  assign n82834 = n81905 & ~n82833;
  assign n82835 = ~n81917 & n81949;
  assign n82836 = ~n81969 & ~n81971;
  assign n82837 = ~n82835 & n82836;
  assign n82838 = n81911 & ~n82837;
  assign n82839 = n81938 & n81962;
  assign n82840 = ~n81943 & ~n82839;
  assign n82841 = ~n82838 & n82840;
  assign n82842 = ~n82340 & ~n82346;
  assign n82843 = ~n81911 & ~n82842;
  assign n82844 = n82841 & ~n82843;
  assign n82845 = ~n81905 & ~n82844;
  assign n82846 = ~n82834 & ~n82845;
  assign n82847 = ~n81917 & n81982;
  assign n82848 = n81917 & ~n82343;
  assign n82849 = ~n82847 & ~n82848;
  assign n82850 = ~n81911 & ~n82849;
  assign n82851 = ~n81969 & n82376;
  assign n82852 = n81973 & ~n82851;
  assign n82853 = ~n82850 & ~n82852;
  assign n82854 = n82846 & n82853;
  assign n82855 = ~pi2608 & ~n82854;
  assign n82856 = ~n82834 & n82853;
  assign n82857 = ~n82845 & n82856;
  assign n82858 = pi2608 & n82857;
  assign po2747 = n82855 | n82858;
  assign n82860 = ~n82470 & n82487;
  assign n82861 = ~n82470 & n82502;
  assign n82862 = ~n82860 & ~n82861;
  assign n82863 = ~n82476 & ~n82862;
  assign n82864 = n82470 & ~n82476;
  assign n82865 = n82499 & n82864;
  assign n82866 = ~n82863 & ~n82865;
  assign n82867 = ~n82523 & n82866;
  assign n82868 = n82451 & n82476;
  assign n82869 = n82463 & n82868;
  assign n82870 = ~n82457 & n82869;
  assign n82871 = ~n82470 & n82870;
  assign n82872 = n82451 & n82464;
  assign n82873 = n82476 & n82872;
  assign n82874 = ~n82495 & ~n82521;
  assign n82875 = ~n82489 & n82874;
  assign n82876 = ~n82873 & n82875;
  assign n82877 = n82445 & ~n82876;
  assign n82878 = n82451 & n82470;
  assign n82879 = ~n82463 & n82878;
  assign n82880 = n82470 & n82532;
  assign n82881 = ~n82870 & ~n82880;
  assign n82882 = ~n82879 & n82881;
  assign n82883 = n82463 & n82493;
  assign n82884 = n82470 & n82481;
  assign n82885 = ~n82498 & ~n82884;
  assign n82886 = ~n82476 & ~n82885;
  assign n82887 = ~n82883 & ~n82886;
  assign n82888 = n82882 & n82887;
  assign n82889 = ~n82445 & ~n82888;
  assign n82890 = n82470 & n82507;
  assign n82891 = ~n82502 & ~n82890;
  assign n82892 = n82451 & n82511;
  assign n82893 = n82891 & ~n82892;
  assign n82894 = ~n82476 & ~n82893;
  assign n82895 = n82445 & n82894;
  assign n82896 = ~n82889 & ~n82895;
  assign n82897 = ~n82877 & n82896;
  assign n82898 = ~n82871 & n82897;
  assign n82899 = n82867 & n82898;
  assign n82900 = pi2611 & ~n82899;
  assign n82901 = ~pi2611 & n82867;
  assign n82902 = n82898 & n82901;
  assign po2748 = n82900 | n82902;
  assign n82904 = ~n82809 & ~n82811;
  assign n82905 = n82718 & ~n82904;
  assign n82906 = ~n82782 & ~n82905;
  assign n82907 = n82724 & ~n82906;
  assign n82908 = n82686 & n82724;
  assign n82909 = ~n82701 & n82908;
  assign n82910 = ~n82709 & n82909;
  assign n82911 = n82701 & n82744;
  assign n82912 = n82718 & n82911;
  assign n82913 = n82686 & ~n82692;
  assign n82914 = n82749 & n82913;
  assign n82915 = ~n82912 & ~n82914;
  assign n82916 = ~n82910 & n82915;
  assign n82917 = ~n82686 & n82698;
  assign n82918 = ~n82701 & ~n82917;
  assign n82919 = n82709 & ~n82918;
  assign n82920 = ~n82778 & ~n82919;
  assign n82921 = ~n82718 & ~n82920;
  assign n82922 = ~n82803 & ~n82921;
  assign n82923 = ~n82709 & n82760;
  assign n82924 = ~n82692 & n82710;
  assign n82925 = ~n82709 & ~n82918;
  assign n82926 = ~n82924 & ~n82925;
  assign n82927 = n82718 & ~n82926;
  assign n82928 = ~n82923 & ~n82927;
  assign n82929 = n82922 & n82928;
  assign n82930 = ~n82724 & ~n82929;
  assign n82931 = ~n82728 & ~n82807;
  assign n82932 = n82725 & ~n82931;
  assign n82933 = ~n82930 & ~n82932;
  assign n82934 = n82916 & n82933;
  assign n82935 = ~n82907 & n82934;
  assign n82936 = pi2621 & ~n82935;
  assign n82937 = ~pi2621 & n82935;
  assign po2749 = n82936 | n82937;
  assign n82939 = n82584 & n82608;
  assign n82940 = ~n82593 & ~n82609;
  assign n82941 = ~n82564 & ~n82940;
  assign n82942 = ~n82939 & ~n82941;
  assign n82943 = ~n82578 & ~n82584;
  assign n82944 = ~n82558 & n82943;
  assign n82945 = n82558 & n82585;
  assign n82946 = ~n82944 & ~n82945;
  assign n82947 = ~n82571 & ~n82578;
  assign n82948 = n82946 & ~n82947;
  assign n82949 = ~n82622 & n82948;
  assign n82950 = n82564 & ~n82949;
  assign n82951 = n82942 & ~n82950;
  assign n82952 = ~n82613 & n82951;
  assign n82953 = n82552 & ~n82952;
  assign n82954 = ~n82558 & n82589;
  assign n82955 = n82616 & ~n82954;
  assign n82956 = n82564 & ~n82955;
  assign n82957 = ~n82953 & ~n82956;
  assign n82958 = ~n82558 & n82622;
  assign n82959 = n82571 & ~n82578;
  assign n82960 = ~n82564 & n82959;
  assign n82961 = n82558 & n82960;
  assign n82962 = n82578 & n82606;
  assign n82963 = ~n82584 & n82962;
  assign n82964 = n82558 & n82617;
  assign n82965 = ~n82963 & ~n82964;
  assign n82966 = ~n82571 & n82578;
  assign n82967 = n82558 & n82966;
  assign n82968 = ~n82603 & ~n82967;
  assign n82969 = ~n82564 & ~n82968;
  assign n82970 = ~n82564 & ~n82571;
  assign n82971 = ~n82578 & n82970;
  assign n82972 = ~n82558 & n82971;
  assign n82973 = ~n82969 & ~n82972;
  assign n82974 = n82965 & n82973;
  assign n82975 = ~n82552 & ~n82974;
  assign n82976 = ~n82961 & ~n82975;
  assign n82977 = ~n82958 & n82976;
  assign n82978 = n82957 & n82977;
  assign n82979 = ~pi2606 & ~n82978;
  assign n82980 = ~n82953 & ~n82958;
  assign n82981 = ~n82956 & n82980;
  assign n82982 = n82976 & n82981;
  assign n82983 = pi2606 & n82982;
  assign po2750 = n82979 | n82983;
  assign n82985 = ~n82558 & n82586;
  assign n82986 = ~n82589 & ~n82958;
  assign n82987 = n82558 & n82611;
  assign n82988 = ~n82558 & n82603;
  assign n82989 = ~n82987 & ~n82988;
  assign n82990 = n82986 & n82989;
  assign n82991 = ~n82564 & ~n82990;
  assign n82992 = n82558 & n82592;
  assign n82993 = ~n82609 & ~n82992;
  assign n82994 = ~n82614 & n82993;
  assign n82995 = n82564 & ~n82994;
  assign n82996 = n82558 & ~n82578;
  assign n82997 = n82584 & n82996;
  assign n82998 = n82571 & n82997;
  assign n82999 = ~n82995 & ~n82998;
  assign n83000 = ~n82991 & n82999;
  assign n83001 = ~n82985 & n83000;
  assign n83002 = ~n82552 & ~n83001;
  assign n83003 = n82558 & ~n82564;
  assign n83004 = n82622 & n83003;
  assign n83005 = ~n82564 & n82614;
  assign n83006 = ~n82564 & n82617;
  assign n83007 = ~n83005 & ~n83006;
  assign n83008 = ~n82558 & ~n83007;
  assign n83009 = ~n83004 & ~n83008;
  assign n83010 = n82558 & n82588;
  assign n83011 = ~n82558 & n82592;
  assign n83012 = ~n83010 & ~n83011;
  assign n83013 = ~n82612 & n83012;
  assign n83014 = ~n82589 & n83013;
  assign n83015 = n82564 & ~n83014;
  assign n83016 = ~n82558 & n82593;
  assign n83017 = ~n83015 & ~n83016;
  assign n83018 = ~n82558 & n82612;
  assign n83019 = ~n82604 & ~n83018;
  assign n83020 = n83017 & n83019;
  assign n83021 = n83009 & n83020;
  assign n83022 = n82552 & ~n83021;
  assign n83023 = ~n82564 & ~n82591;
  assign n83024 = ~n83022 & ~n83023;
  assign n83025 = ~n82615 & ~n83018;
  assign n83026 = n82564 & ~n83025;
  assign n83027 = n83024 & ~n83026;
  assign n83028 = ~n83002 & n83027;
  assign n83029 = pi2612 & ~n83028;
  assign n83030 = ~pi2612 & n83028;
  assign po2751 = n83029 | n83030;
  assign n83032 = ~n82200 & ~n82220;
  assign n83033 = n82146 & ~n83032;
  assign n83034 = ~n82138 & ~n82152;
  assign n83035 = ~n82204 & n83034;
  assign n83036 = ~n82101 & ~n83035;
  assign n83037 = n82146 & n83036;
  assign n83038 = ~n83033 & ~n83037;
  assign n83039 = n82147 & n82155;
  assign n83040 = ~n82157 & ~n83039;
  assign n83041 = ~n82151 & ~n82188;
  assign n83042 = n82101 & ~n83041;
  assign n83043 = n82146 & n83042;
  assign n83044 = n83040 & ~n83043;
  assign n83045 = n82119 & n82137;
  assign n83046 = ~n82131 & n83045;
  assign n83047 = n82107 & n82126;
  assign n83048 = ~n82134 & ~n83047;
  assign n83049 = n82101 & ~n83048;
  assign n83050 = ~n82139 & ~n82160;
  assign n83051 = n82107 & n82132;
  assign n83052 = ~n82181 & ~n83051;
  assign n83053 = ~n82101 & ~n83052;
  assign n83054 = n83050 & ~n83053;
  assign n83055 = ~n83049 & n83054;
  assign n83056 = ~n83046 & n83055;
  assign n83057 = ~n82146 & ~n83056;
  assign n83058 = ~n82185 & n82411;
  assign n83059 = n82101 & ~n83058;
  assign n83060 = ~n83057 & ~n83059;
  assign n83061 = n83044 & n83060;
  assign n83062 = n83038 & n83061;
  assign n83063 = ~pi2599 & ~n83062;
  assign n83064 = pi2599 & n83044;
  assign n83065 = n83038 & n83064;
  assign n83066 = n83060 & n83065;
  assign po2752 = n83063 | n83066;
  assign n83068 = ~n82029 & n82038;
  assign n83069 = ~n82065 & ~n83068;
  assign n83070 = ~n82055 & ~n83069;
  assign n83071 = n82055 & ~n82282;
  assign n83072 = ~n82271 & ~n83071;
  assign n83073 = ~n83070 & n83072;
  assign n83074 = n82010 & ~n83073;
  assign n83075 = n82048 & ~n82055;
  assign n83076 = ~n83074 & ~n83075;
  assign n83077 = ~n82648 & ~n82657;
  assign n83078 = n82055 & ~n83077;
  assign n83079 = n82055 & n82066;
  assign n83080 = n82029 & n82039;
  assign n83081 = n82036 & ~n82055;
  assign n83082 = ~n82260 & ~n83081;
  assign n83083 = ~n82016 & ~n83082;
  assign n83084 = ~n82261 & ~n83083;
  assign n83085 = ~n82037 & n83084;
  assign n83086 = ~n83080 & n83085;
  assign n83087 = ~n83079 & n83086;
  assign n83088 = ~n82010 & ~n83087;
  assign n83089 = ~n83078 & ~n83088;
  assign n83090 = n83076 & n83089;
  assign n83091 = pi2635 & ~n83090;
  assign n83092 = ~pi2635 & n83090;
  assign po2753 = n83091 | n83092;
  assign n83094 = n82451 & ~n82457;
  assign n83095 = ~n82495 & ~n83094;
  assign n83096 = ~n82527 & n83095;
  assign n83097 = n82476 & ~n83096;
  assign n83098 = n82457 & n82864;
  assign n83099 = ~n82860 & ~n82879;
  assign n83100 = ~n82451 & ~n82457;
  assign n83101 = ~n82470 & ~n82476;
  assign n83102 = n83100 & n83101;
  assign n83103 = n83099 & ~n83102;
  assign n83104 = ~n83098 & n83103;
  assign n83105 = ~n83097 & n83104;
  assign n83106 = n82445 & ~n83105;
  assign n83107 = ~n82470 & n82872;
  assign n83108 = n82470 & n82892;
  assign n83109 = ~n83107 & ~n83108;
  assign n83110 = n82476 & ~n83109;
  assign n83111 = ~n83106 & ~n83110;
  assign n83112 = n82470 & n82487;
  assign n83113 = ~n82499 & ~n82507;
  assign n83114 = n82476 & ~n83113;
  assign n83115 = ~n83112 & ~n83114;
  assign n83116 = ~n82503 & n83115;
  assign n83117 = ~n82445 & ~n83116;
  assign n83118 = ~n82481 & ~n82511;
  assign n83119 = ~n82451 & ~n83118;
  assign n83120 = ~n82512 & ~n83119;
  assign n83121 = ~n82476 & ~n83120;
  assign n83122 = ~n82445 & n83121;
  assign n83123 = ~n83117 & ~n83122;
  assign n83124 = n83111 & n83123;
  assign n83125 = pi2602 & ~n83124;
  assign n83126 = ~pi2602 & n83111;
  assign n83127 = n83123 & n83126;
  assign po2754 = n83125 | n83127;
  assign n83129 = ~n82686 & n82809;
  assign n83130 = ~n82758 & ~n83129;
  assign n83131 = n82718 & ~n83130;
  assign n83132 = ~n82686 & n82701;
  assign n83133 = ~n82778 & ~n83132;
  assign n83134 = n82718 & ~n83133;
  assign n83135 = n82709 & n82727;
  assign n83136 = ~n82702 & ~n83135;
  assign n83137 = ~n82760 & n83136;
  assign n83138 = ~n82718 & ~n83137;
  assign n83139 = ~n83134 & ~n83138;
  assign n83140 = ~n82732 & ~n82743;
  assign n83141 = n83139 & n83140;
  assign n83142 = ~n82724 & ~n83141;
  assign n83143 = n82718 & n82728;
  assign n83144 = n82703 & ~n83143;
  assign n83145 = ~n82760 & n83144;
  assign n83146 = n82709 & ~n83145;
  assign n83147 = ~n82709 & n82778;
  assign n83148 = n82699 & n82709;
  assign n83149 = ~n82809 & ~n83148;
  assign n83150 = ~n82718 & ~n83149;
  assign n83151 = ~n83147 & ~n83150;
  assign n83152 = ~n83146 & n83151;
  assign n83153 = n82724 & ~n83152;
  assign n83154 = ~n83142 & ~n83153;
  assign n83155 = n82749 & n82917;
  assign n83156 = n83154 & ~n83155;
  assign n83157 = ~n83131 & n83156;
  assign n83158 = ~pi2627 & ~n83157;
  assign n83159 = pi2627 & ~n83131;
  assign n83160 = n83154 & n83159;
  assign n83161 = ~n83155 & n83160;
  assign po2755 = n83158 | n83161;
  assign n83163 = ~n82470 & n82499;
  assign n83164 = n82470 & n82872;
  assign n83165 = ~n83163 & ~n83164;
  assign n83166 = ~n82476 & ~n83165;
  assign n83167 = n82470 & n83119;
  assign n83168 = ~n82506 & ~n82872;
  assign n83169 = ~n82476 & ~n83168;
  assign n83170 = ~n83167 & ~n83169;
  assign n83171 = n82463 & n82878;
  assign n83172 = ~n82535 & ~n83171;
  assign n83173 = ~n82892 & n83172;
  assign n83174 = n82476 & ~n83173;
  assign n83175 = n83170 & ~n83174;
  assign n83176 = ~n83163 & n83175;
  assign n83177 = ~n82445 & ~n83176;
  assign n83178 = n82480 & ~n83168;
  assign n83179 = ~n82502 & ~n82507;
  assign n83180 = ~n82499 & ~n82892;
  assign n83181 = n83179 & n83180;
  assign n83182 = n82470 & ~n83181;
  assign n83183 = ~n83178 & ~n83182;
  assign n83184 = ~n82860 & n83183;
  assign n83185 = n82445 & ~n83184;
  assign n83186 = ~n83177 & ~n83185;
  assign n83187 = ~n83166 & n83186;
  assign n83188 = pi2595 & ~n83187;
  assign n83189 = ~pi2595 & ~n83185;
  assign n83190 = ~n83166 & n83189;
  assign n83191 = ~n83177 & n83190;
  assign po2756 = n83188 | n83191;
  assign n83193 = ~n82596 & ~n83018;
  assign n83194 = ~n82998 & n83193;
  assign n83195 = ~n82564 & ~n83194;
  assign n83196 = ~n82604 & ~n83006;
  assign n83197 = ~n82586 & ~n83011;
  assign n83198 = n82564 & ~n83197;
  assign n83199 = ~n82958 & ~n83198;
  assign n83200 = n83196 & n83199;
  assign n83201 = n82552 & ~n83200;
  assign n83202 = ~n82578 & n82584;
  assign n83203 = ~n82947 & ~n83202;
  assign n83204 = n82558 & ~n83203;
  assign n83205 = ~n82612 & ~n82619;
  assign n83206 = n82564 & ~n83205;
  assign n83207 = n82558 & n82584;
  assign n83208 = ~n82593 & ~n83207;
  assign n83209 = ~n82585 & n83208;
  assign n83210 = ~n82564 & ~n83209;
  assign n83211 = ~n83206 & ~n83210;
  assign n83212 = ~n83204 & n83211;
  assign n83213 = ~n82552 & ~n83212;
  assign n83214 = ~n83201 & ~n83213;
  assign n83215 = ~n82607 & ~n82634;
  assign n83216 = n83214 & n83215;
  assign n83217 = ~n83195 & n83216;
  assign n83218 = ~pi2622 & ~n83217;
  assign n83219 = pi2622 & n83215;
  assign n83220 = ~n83195 & n83219;
  assign n83221 = n83214 & n83220;
  assign po2757 = n83218 | n83221;
  assign n83223 = pi5934 & pi9040;
  assign n83224 = pi6018 & ~pi9040;
  assign n83225 = ~n83223 & ~n83224;
  assign n83226 = ~pi2649 & ~n83225;
  assign n83227 = pi2649 & n83225;
  assign n83228 = ~n83226 & ~n83227;
  assign n83229 = pi5932 & ~pi9040;
  assign n83230 = pi6011 & pi9040;
  assign n83231 = ~n83229 & ~n83230;
  assign n83232 = pi2640 & n83231;
  assign n83233 = ~pi2640 & ~n83231;
  assign n83234 = ~n83232 & ~n83233;
  assign n83235 = pi5737 & pi9040;
  assign n83236 = pi5873 & ~pi9040;
  assign n83237 = ~n83235 & ~n83236;
  assign n83238 = ~pi2639 & ~n83237;
  assign n83239 = pi2639 & n83237;
  assign n83240 = ~n83238 & ~n83239;
  assign n83241 = pi5849 & pi9040;
  assign n83242 = pi5781 & ~pi9040;
  assign n83243 = ~n83241 & ~n83242;
  assign n83244 = ~pi2631 & ~n83243;
  assign n83245 = pi2631 & n83243;
  assign n83246 = ~n83244 & ~n83245;
  assign n83247 = pi5810 & pi9040;
  assign n83248 = pi6011 & ~pi9040;
  assign n83249 = ~n83247 & ~n83248;
  assign n83250 = pi2645 & n83249;
  assign n83251 = ~pi2645 & ~n83249;
  assign n83252 = ~n83250 & ~n83251;
  assign n83253 = ~n83246 & ~n83252;
  assign n83254 = ~n83240 & n83253;
  assign n83255 = pi5910 & ~pi9040;
  assign n83256 = pi5811 & pi9040;
  assign n83257 = ~n83255 & ~n83256;
  assign n83258 = ~pi2613 & ~n83257;
  assign n83259 = pi2613 & n83257;
  assign n83260 = ~n83258 & ~n83259;
  assign n83261 = ~n83240 & ~n83260;
  assign n83262 = n83252 & n83261;
  assign n83263 = n83246 & n83262;
  assign n83264 = ~n83254 & ~n83263;
  assign n83265 = ~n83240 & n83260;
  assign n83266 = ~n83252 & n83265;
  assign n83267 = n83240 & n83260;
  assign n83268 = n83252 & n83267;
  assign n83269 = ~n83266 & ~n83268;
  assign n83270 = n83264 & n83269;
  assign n83271 = n83234 & ~n83270;
  assign n83272 = n83240 & ~n83260;
  assign n83273 = ~n83252 & n83272;
  assign n83274 = n83246 & n83273;
  assign n83275 = ~n83271 & ~n83274;
  assign n83276 = ~n83228 & ~n83275;
  assign n83277 = ~n83228 & ~n83234;
  assign n83278 = n83252 & ~n83260;
  assign n83279 = ~n83246 & n83278;
  assign n83280 = n83252 & n83265;
  assign n83281 = n83246 & n83280;
  assign n83282 = ~n83246 & n83267;
  assign n83283 = ~n83281 & ~n83282;
  assign n83284 = ~n83279 & n83283;
  assign n83285 = n83277 & ~n83284;
  assign n83286 = ~n83276 & ~n83285;
  assign n83287 = ~n83252 & n83261;
  assign n83288 = ~n83261 & ~n83267;
  assign n83289 = n83246 & ~n83288;
  assign n83290 = ~n83287 & ~n83289;
  assign n83291 = ~n83234 & ~n83290;
  assign n83292 = n83252 & n83272;
  assign n83293 = ~n83279 & ~n83292;
  assign n83294 = ~n83281 & n83293;
  assign n83295 = n83234 & ~n83294;
  assign n83296 = ~n83291 & ~n83295;
  assign n83297 = ~n83234 & ~n83246;
  assign n83298 = n83265 & n83297;
  assign n83299 = n83246 & n83287;
  assign n83300 = ~n83252 & n83260;
  assign n83301 = n83240 & n83300;
  assign n83302 = n83246 & n83301;
  assign n83303 = ~n83299 & ~n83302;
  assign n83304 = n83240 & n83253;
  assign n83305 = ~n83260 & n83304;
  assign n83306 = n83303 & ~n83305;
  assign n83307 = ~n83298 & n83306;
  assign n83308 = n83296 & n83307;
  assign n83309 = n83228 & ~n83308;
  assign n83310 = n83234 & ~n83246;
  assign n83311 = n83252 & n83310;
  assign n83312 = n83240 & n83311;
  assign n83313 = ~n83246 & n83266;
  assign n83314 = ~n83312 & ~n83313;
  assign n83315 = ~n83309 & n83314;
  assign n83316 = n83286 & n83315;
  assign n83317 = pi2669 & ~n83316;
  assign n83318 = ~pi2669 & n83314;
  assign n83319 = n83286 & n83318;
  assign n83320 = ~n83309 & n83319;
  assign po2767 = n83317 | n83320;
  assign n83322 = ~n83287 & ~n83292;
  assign n83323 = ~n83234 & ~n83322;
  assign n83324 = n83246 & n83268;
  assign n83325 = ~n83323 & ~n83324;
  assign n83326 = n83246 & n83260;
  assign n83327 = ~n83300 & ~n83326;
  assign n83328 = ~n83262 & n83327;
  assign n83329 = n83234 & ~n83328;
  assign n83330 = n83325 & ~n83329;
  assign n83331 = ~n83228 & ~n83330;
  assign n83332 = ~n83246 & n83301;
  assign n83333 = ~n83234 & n83332;
  assign n83334 = ~n83246 & n83252;
  assign n83335 = ~n83240 & n83334;
  assign n83336 = n83260 & n83335;
  assign n83337 = ~n83234 & n83336;
  assign n83338 = ~n83333 & ~n83337;
  assign n83339 = n83234 & n83305;
  assign n83340 = n83338 & ~n83339;
  assign n83341 = n83234 & ~n83252;
  assign n83342 = n83240 & n83341;
  assign n83343 = ~n83260 & n83342;
  assign n83344 = n83260 & n83334;
  assign n83345 = n83234 & n83344;
  assign n83346 = n83246 & n83292;
  assign n83347 = ~n83234 & n83300;
  assign n83348 = ~n83346 & ~n83347;
  assign n83349 = ~n83299 & n83348;
  assign n83350 = ~n83345 & n83349;
  assign n83351 = ~n83305 & ~n83335;
  assign n83352 = n83350 & n83351;
  assign n83353 = ~n83343 & n83352;
  assign n83354 = n83228 & ~n83353;
  assign n83355 = n83340 & ~n83354;
  assign n83356 = ~n83331 & n83355;
  assign n83357 = ~pi2670 & ~n83356;
  assign n83358 = pi2670 & n83340;
  assign n83359 = ~n83331 & n83358;
  assign n83360 = ~n83354 & n83359;
  assign po2778 = n83357 | n83360;
  assign n83362 = pi5791 & ~pi9040;
  assign n83363 = pi6037 & pi9040;
  assign n83364 = ~n83362 & ~n83363;
  assign n83365 = ~pi2634 & n83364;
  assign n83366 = pi2634 & ~n83364;
  assign n83367 = ~n83365 & ~n83366;
  assign n83368 = pi5812 & pi9040;
  assign n83369 = pi6158 & ~pi9040;
  assign n83370 = ~n83368 & ~n83369;
  assign n83371 = pi2654 & n83370;
  assign n83372 = ~pi2654 & ~n83370;
  assign n83373 = ~n83371 & ~n83372;
  assign n83374 = pi5727 & pi9040;
  assign n83375 = pi5814 & ~pi9040;
  assign n83376 = ~n83374 & ~n83375;
  assign n83377 = pi2625 & n83376;
  assign n83378 = ~pi2625 & ~n83376;
  assign n83379 = ~n83377 & ~n83378;
  assign n83380 = pi5891 & ~pi9040;
  assign n83381 = pi5944 & pi9040;
  assign n83382 = ~n83380 & ~n83381;
  assign n83383 = pi2651 & n83382;
  assign n83384 = ~pi2651 & ~n83382;
  assign n83385 = ~n83383 & ~n83384;
  assign n83386 = pi5747 & ~pi9040;
  assign n83387 = pi5879 & pi9040;
  assign n83388 = ~n83386 & ~n83387;
  assign n83389 = ~pi2645 & ~n83388;
  assign n83390 = pi2645 & n83388;
  assign n83391 = ~n83389 & ~n83390;
  assign n83392 = ~n83385 & n83391;
  assign n83393 = ~n83379 & n83392;
  assign n83394 = ~n83373 & n83393;
  assign n83395 = n83379 & ~n83391;
  assign n83396 = n83385 & n83395;
  assign n83397 = n83373 & n83396;
  assign n83398 = ~n83385 & ~n83391;
  assign n83399 = ~n83379 & n83398;
  assign n83400 = n83373 & n83399;
  assign n83401 = ~n83397 & ~n83400;
  assign n83402 = ~n83394 & n83401;
  assign n83403 = ~n83367 & ~n83402;
  assign n83404 = ~n83373 & n83379;
  assign n83405 = n83391 & n83404;
  assign n83406 = n83385 & n83405;
  assign n83407 = pi5745 & pi9040;
  assign n83408 = pi5727 & ~pi9040;
  assign n83409 = ~n83407 & ~n83408;
  assign n83410 = ~pi2613 & ~n83409;
  assign n83411 = pi2613 & n83409;
  assign n83412 = ~n83410 & ~n83411;
  assign n83413 = ~n83385 & n83404;
  assign n83414 = n83385 & n83391;
  assign n83415 = ~n83379 & n83414;
  assign n83416 = ~n83413 & ~n83415;
  assign n83417 = n83367 & ~n83416;
  assign n83418 = ~n83405 & ~n83417;
  assign n83419 = n83379 & n83414;
  assign n83420 = ~n83379 & ~n83385;
  assign n83421 = ~n83379 & ~n83391;
  assign n83422 = ~n83373 & n83421;
  assign n83423 = n83373 & n83398;
  assign n83424 = ~n83422 & ~n83423;
  assign n83425 = ~n83420 & n83424;
  assign n83426 = ~n83419 & n83425;
  assign n83427 = ~n83367 & ~n83426;
  assign n83428 = n83418 & ~n83427;
  assign n83429 = ~n83397 & n83428;
  assign n83430 = n83412 & ~n83429;
  assign n83431 = ~n83406 & ~n83430;
  assign n83432 = ~n83403 & n83431;
  assign n83433 = n83373 & ~n83379;
  assign n83434 = n83367 & n83433;
  assign n83435 = n83385 & n83434;
  assign n83436 = n83379 & n83392;
  assign n83437 = n83373 & n83436;
  assign n83438 = ~n83367 & n83395;
  assign n83439 = ~n83373 & n83438;
  assign n83440 = ~n83437 & ~n83439;
  assign n83441 = n83379 & ~n83385;
  assign n83442 = n83373 & n83441;
  assign n83443 = n83385 & ~n83391;
  assign n83444 = ~n83379 & n83443;
  assign n83445 = ~n83442 & ~n83444;
  assign n83446 = n83367 & ~n83445;
  assign n83447 = n83367 & n83420;
  assign n83448 = ~n83373 & n83447;
  assign n83449 = ~n83446 & ~n83448;
  assign n83450 = n83440 & n83449;
  assign n83451 = ~n83412 & ~n83450;
  assign n83452 = ~n83435 & ~n83451;
  assign n83453 = n83432 & n83452;
  assign n83454 = pi2671 & n83453;
  assign n83455 = ~n83406 & ~n83435;
  assign n83456 = ~n83451 & n83455;
  assign n83457 = ~n83403 & ~n83430;
  assign n83458 = n83456 & n83457;
  assign n83459 = ~pi2671 & ~n83458;
  assign po2784 = n83454 | n83459;
  assign n83461 = n83240 & n83246;
  assign n83462 = n83252 & n83461;
  assign n83463 = ~n83246 & ~n83260;
  assign n83464 = ~n83335 & ~n83463;
  assign n83465 = ~n83234 & ~n83464;
  assign n83466 = ~n83462 & ~n83465;
  assign n83467 = n83234 & n83267;
  assign n83468 = ~n83246 & n83467;
  assign n83469 = ~n83246 & n83262;
  assign n83470 = ~n83468 & ~n83469;
  assign n83471 = n83466 & n83470;
  assign n83472 = n83228 & ~n83471;
  assign n83473 = ~n83280 & ~n83302;
  assign n83474 = ~n83246 & n83272;
  assign n83475 = n83473 & ~n83474;
  assign n83476 = n83234 & ~n83475;
  assign n83477 = n83267 & n83297;
  assign n83478 = ~n83313 & ~n83477;
  assign n83479 = ~n83476 & n83478;
  assign n83480 = ~n83262 & ~n83274;
  assign n83481 = ~n83234 & ~n83480;
  assign n83482 = n83479 & ~n83481;
  assign n83483 = ~n83228 & ~n83482;
  assign n83484 = ~n83472 & ~n83483;
  assign n83485 = n83246 & n83269;
  assign n83486 = ~n83246 & ~n83261;
  assign n83487 = ~n83485 & ~n83486;
  assign n83488 = ~n83234 & n83487;
  assign n83489 = n83234 & n83246;
  assign n83490 = ~n83280 & n83322;
  assign n83491 = n83489 & ~n83490;
  assign n83492 = ~n83488 & ~n83491;
  assign n83493 = n83484 & n83492;
  assign n83494 = ~pi2679 & ~n83493;
  assign n83495 = pi2679 & n83492;
  assign n83496 = ~n83483 & n83495;
  assign n83497 = ~n83472 & n83496;
  assign po2787 = n83494 | n83497;
  assign n83499 = n83246 & n83278;
  assign n83500 = ~n83268 & ~n83499;
  assign n83501 = ~n83313 & n83500;
  assign n83502 = n83234 & ~n83501;
  assign n83503 = ~n83246 & n83292;
  assign n83504 = ~n83252 & ~n83260;
  assign n83505 = ~n83265 & ~n83504;
  assign n83506 = n83246 & ~n83505;
  assign n83507 = ~n83503 & ~n83506;
  assign n83508 = ~n83332 & n83507;
  assign n83509 = ~n83234 & ~n83508;
  assign n83510 = ~n83502 & ~n83509;
  assign n83511 = n83228 & ~n83510;
  assign n83512 = ~n83260 & n83310;
  assign n83513 = ~n83344 & ~n83499;
  assign n83514 = ~n83234 & ~n83513;
  assign n83515 = ~n83298 & ~n83514;
  assign n83516 = ~n83302 & ~n83336;
  assign n83517 = n83300 & n83489;
  assign n83518 = ~n83343 & ~n83517;
  assign n83519 = n83516 & n83518;
  assign n83520 = n83515 & n83519;
  assign n83521 = ~n83512 & n83520;
  assign n83522 = ~n83228 & ~n83521;
  assign n83523 = ~n83234 & n83287;
  assign n83524 = ~n83246 & n83523;
  assign n83525 = ~n83337 & ~n83524;
  assign n83526 = ~n83339 & n83525;
  assign n83527 = n83246 & n83267;
  assign n83528 = ~n83469 & ~n83527;
  assign n83529 = n83234 & ~n83528;
  assign n83530 = n83526 & ~n83529;
  assign n83531 = ~n83522 & n83530;
  assign n83532 = ~n83511 & n83531;
  assign n83533 = ~pi2677 & n83532;
  assign n83534 = pi2677 & ~n83532;
  assign po2788 = n83533 | n83534;
  assign n83536 = pi5934 & ~pi9040;
  assign n83537 = pi5781 & pi9040;
  assign n83538 = ~n83536 & ~n83537;
  assign n83539 = pi2653 & n83538;
  assign n83540 = ~pi2653 & ~n83538;
  assign n83541 = ~n83539 & ~n83540;
  assign n83542 = pi5804 & ~pi9040;
  assign n83543 = pi5871 & pi9040;
  assign n83544 = ~n83542 & ~n83543;
  assign n83545 = ~pi2610 & ~n83544;
  assign n83546 = pi2610 & n83544;
  assign n83547 = ~n83545 & ~n83546;
  assign n83548 = pi5732 & ~pi9040;
  assign n83549 = pi5862 & pi9040;
  assign n83550 = ~n83548 & ~n83549;
  assign n83551 = pi2639 & n83550;
  assign n83552 = ~pi2639 & ~n83550;
  assign n83553 = ~n83551 & ~n83552;
  assign n83554 = pi5804 & pi9040;
  assign n83555 = pi5862 & ~pi9040;
  assign n83556 = ~n83554 & ~n83555;
  assign n83557 = ~pi2649 & n83556;
  assign n83558 = pi2649 & ~n83556;
  assign n83559 = ~n83557 & ~n83558;
  assign n83560 = n83553 & ~n83559;
  assign n83561 = n83547 & n83560;
  assign n83562 = n83553 & n83559;
  assign n83563 = ~n83547 & n83562;
  assign n83564 = ~n83561 & ~n83563;
  assign n83565 = ~n83541 & ~n83564;
  assign n83566 = pi5725 & pi9040;
  assign n83567 = pi5871 & ~pi9040;
  assign n83568 = ~n83566 & ~n83567;
  assign n83569 = pi2638 & n83568;
  assign n83570 = ~pi2638 & ~n83568;
  assign n83571 = ~n83569 & ~n83570;
  assign n83572 = pi5811 & ~pi9040;
  assign n83573 = pi5873 & pi9040;
  assign n83574 = ~n83572 & ~n83573;
  assign n83575 = pi2629 & n83574;
  assign n83576 = ~pi2629 & ~n83574;
  assign n83577 = ~n83575 & ~n83576;
  assign n83578 = ~n83559 & ~n83577;
  assign n83579 = ~n83553 & n83578;
  assign n83580 = ~n83547 & n83579;
  assign n83581 = n83559 & n83577;
  assign n83582 = ~n83541 & ~n83547;
  assign n83583 = n83581 & n83582;
  assign n83584 = ~n83553 & ~n83559;
  assign n83585 = n83541 & ~n83547;
  assign n83586 = n83584 & n83585;
  assign n83587 = n83553 & n83578;
  assign n83588 = n83547 & ~n83553;
  assign n83589 = ~n83577 & n83588;
  assign n83590 = n83559 & n83589;
  assign n83591 = ~n83587 & ~n83590;
  assign n83592 = ~n83559 & n83577;
  assign n83593 = n83547 & n83592;
  assign n83594 = n83591 & ~n83593;
  assign n83595 = ~n83541 & ~n83594;
  assign n83596 = ~n83586 & ~n83595;
  assign n83597 = ~n83583 & n83596;
  assign n83598 = ~n83580 & n83597;
  assign n83599 = n83553 & n83592;
  assign n83600 = n83547 & n83599;
  assign n83601 = n83553 & n83581;
  assign n83602 = ~n83547 & n83601;
  assign n83603 = ~n83600 & ~n83602;
  assign n83604 = n83598 & n83603;
  assign n83605 = ~n83571 & ~n83604;
  assign n83606 = ~n83553 & ~n83577;
  assign n83607 = n83541 & n83606;
  assign n83608 = ~n83547 & n83607;
  assign n83609 = n83559 & ~n83577;
  assign n83610 = n83553 & n83609;
  assign n83611 = n83547 & n83610;
  assign n83612 = n83581 & n83588;
  assign n83613 = ~n83611 & ~n83612;
  assign n83614 = ~n83579 & n83613;
  assign n83615 = n83541 & ~n83614;
  assign n83616 = ~n83608 & ~n83615;
  assign n83617 = ~n83547 & ~n83553;
  assign n83618 = n83577 & n83617;
  assign n83619 = ~n83559 & n83618;
  assign n83620 = ~n83601 & ~n83619;
  assign n83621 = ~n83541 & ~n83620;
  assign n83622 = ~n83577 & n83617;
  assign n83623 = n83559 & n83622;
  assign n83624 = ~n83612 & ~n83623;
  assign n83625 = ~n83559 & n83588;
  assign n83626 = ~n83547 & n83599;
  assign n83627 = ~n83625 & ~n83626;
  assign n83628 = n83541 & ~n83627;
  assign n83629 = n83624 & ~n83628;
  assign n83630 = ~n83621 & n83629;
  assign n83631 = n83571 & ~n83630;
  assign n83632 = n83616 & ~n83631;
  assign n83633 = ~n83605 & n83632;
  assign n83634 = ~n83565 & n83633;
  assign n83635 = ~pi2656 & ~n83634;
  assign n83636 = pi2656 & n83634;
  assign po2789 = n83635 | n83636;
  assign n83638 = pi5746 & ~pi9040;
  assign n83639 = pi6002 & pi9040;
  assign n83640 = ~n83638 & ~n83639;
  assign n83641 = ~pi2655 & ~n83640;
  assign n83642 = pi2655 & n83640;
  assign n83643 = ~n83641 & ~n83642;
  assign n83644 = pi5884 & ~pi9040;
  assign n83645 = pi5741 & pi9040;
  assign n83646 = ~n83644 & ~n83645;
  assign n83647 = ~pi2644 & n83646;
  assign n83648 = pi2644 & ~n83646;
  assign n83649 = ~n83647 & ~n83648;
  assign n83650 = pi5951 & ~pi9040;
  assign n83651 = pi5800 & pi9040;
  assign n83652 = ~n83650 & ~n83651;
  assign n83653 = pi2643 & n83652;
  assign n83654 = ~pi2643 & ~n83652;
  assign n83655 = ~n83653 & ~n83654;
  assign n83656 = pi5881 & pi9040;
  assign n83657 = pi5800 & ~pi9040;
  assign n83658 = ~n83656 & ~n83657;
  assign n83659 = ~pi2625 & ~n83658;
  assign n83660 = pi2625 & n83658;
  assign n83661 = ~n83659 & ~n83660;
  assign n83662 = pi5799 & ~pi9040;
  assign n83663 = pi6146 & pi9040;
  assign n83664 = ~n83662 & ~n83663;
  assign n83665 = ~pi2637 & n83664;
  assign n83666 = pi2637 & ~n83664;
  assign n83667 = ~n83665 & ~n83666;
  assign n83668 = ~n83661 & n83667;
  assign n83669 = ~n83655 & n83668;
  assign n83670 = n83649 & n83669;
  assign n83671 = ~n83661 & ~n83667;
  assign n83672 = ~n83655 & n83671;
  assign n83673 = ~n83649 & n83672;
  assign n83674 = ~n83670 & ~n83673;
  assign n83675 = n83643 & ~n83674;
  assign n83676 = pi6028 & ~pi9040;
  assign n83677 = pi5874 & pi9040;
  assign n83678 = ~n83676 & ~n83677;
  assign n83679 = ~pi2651 & ~n83678;
  assign n83680 = pi2651 & n83678;
  assign n83681 = ~n83679 & ~n83680;
  assign n83682 = n83649 & n83655;
  assign n83683 = n83661 & n83682;
  assign n83684 = n83667 & n83683;
  assign n83685 = n83655 & n83671;
  assign n83686 = n83643 & n83685;
  assign n83687 = ~n83684 & ~n83686;
  assign n83688 = n83649 & ~n83667;
  assign n83689 = ~n83655 & n83688;
  assign n83690 = n83667 & n83682;
  assign n83691 = ~n83689 & ~n83690;
  assign n83692 = ~n83643 & ~n83691;
  assign n83693 = ~n83643 & ~n83649;
  assign n83694 = n83668 & n83693;
  assign n83695 = ~n83655 & n83694;
  assign n83696 = n83661 & ~n83667;
  assign n83697 = n83655 & n83696;
  assign n83698 = ~n83649 & n83697;
  assign n83699 = n83643 & ~n83655;
  assign n83700 = n83661 & n83699;
  assign n83701 = n83667 & n83700;
  assign n83702 = ~n83698 & ~n83701;
  assign n83703 = ~n83695 & n83702;
  assign n83704 = ~n83692 & n83703;
  assign n83705 = n83687 & n83704;
  assign n83706 = n83681 & ~n83705;
  assign n83707 = ~n83643 & n83684;
  assign n83708 = n83643 & n83649;
  assign n83709 = n83671 & n83708;
  assign n83710 = n83655 & n83709;
  assign n83711 = ~n83707 & ~n83710;
  assign n83712 = ~n83706 & n83711;
  assign n83713 = ~n83675 & n83712;
  assign n83714 = n83643 & ~n83649;
  assign n83715 = n83655 & n83667;
  assign n83716 = n83714 & n83715;
  assign n83717 = n83643 & n83669;
  assign n83718 = ~n83716 & ~n83717;
  assign n83719 = n83643 & n83697;
  assign n83720 = ~n83655 & n83696;
  assign n83721 = n83649 & n83720;
  assign n83722 = ~n83719 & ~n83721;
  assign n83723 = n83655 & n83668;
  assign n83724 = ~n83649 & n83723;
  assign n83725 = ~n83670 & ~n83724;
  assign n83726 = ~n83649 & n83671;
  assign n83727 = ~n83655 & n83661;
  assign n83728 = ~n83726 & ~n83727;
  assign n83729 = ~n83643 & ~n83728;
  assign n83730 = n83725 & ~n83729;
  assign n83731 = n83722 & n83730;
  assign n83732 = n83718 & n83731;
  assign n83733 = ~n83681 & ~n83732;
  assign n83734 = n83713 & ~n83733;
  assign n83735 = ~pi2663 & ~n83734;
  assign n83736 = pi2663 & n83713;
  assign n83737 = ~n83733 & n83736;
  assign po2790 = n83735 | n83737;
  assign n83739 = pi5944 & ~pi9040;
  assign n83740 = pi6158 & pi9040;
  assign n83741 = ~n83739 & ~n83740;
  assign n83742 = pi2630 & n83741;
  assign n83743 = ~pi2630 & ~n83741;
  assign n83744 = ~n83742 & ~n83743;
  assign n83745 = pi5791 & pi9040;
  assign n83746 = pi5745 & ~pi9040;
  assign n83747 = ~n83745 & ~n83746;
  assign n83748 = ~pi2629 & n83747;
  assign n83749 = pi2629 & ~n83747;
  assign n83750 = ~n83748 & ~n83749;
  assign n83751 = pi5747 & pi9040;
  assign n83752 = pi6037 & ~pi9040;
  assign n83753 = ~n83751 & ~n83752;
  assign n83754 = ~pi2626 & n83753;
  assign n83755 = pi2626 & ~n83753;
  assign n83756 = ~n83754 & ~n83755;
  assign n83757 = pi5891 & pi9040;
  assign n83758 = pi5849 & ~pi9040;
  assign n83759 = ~n83757 & ~n83758;
  assign n83760 = ~pi2638 & ~n83759;
  assign n83761 = pi2638 & n83759;
  assign n83762 = ~n83760 & ~n83761;
  assign n83763 = ~n83756 & n83762;
  assign n83764 = n83750 & n83763;
  assign n83765 = pi5932 & pi9040;
  assign n83766 = pi5879 & ~pi9040;
  assign n83767 = ~n83765 & ~n83766;
  assign n83768 = pi2650 & n83767;
  assign n83769 = ~pi2650 & ~n83767;
  assign n83770 = ~n83768 & ~n83769;
  assign n83771 = n83764 & ~n83770;
  assign n83772 = n83756 & ~n83762;
  assign n83773 = n83750 & n83772;
  assign n83774 = ~n83770 & n83773;
  assign n83775 = ~n83771 & ~n83774;
  assign n83776 = ~n83750 & n83770;
  assign n83777 = n83772 & n83776;
  assign n83778 = ~n83756 & ~n83762;
  assign n83779 = n83750 & n83778;
  assign n83780 = n83770 & n83779;
  assign n83781 = ~n83777 & ~n83780;
  assign n83782 = n83775 & n83781;
  assign n83783 = n83744 & ~n83782;
  assign n83784 = pi5814 & pi9040;
  assign n83785 = pi5725 & ~pi9040;
  assign n83786 = ~n83784 & ~n83785;
  assign n83787 = ~pi2647 & ~n83786;
  assign n83788 = pi2647 & n83786;
  assign n83789 = ~n83787 & ~n83788;
  assign n83790 = n83750 & n83770;
  assign n83791 = n83762 & n83790;
  assign n83792 = n83756 & n83791;
  assign n83793 = ~n83779 & ~n83792;
  assign n83794 = n83744 & ~n83793;
  assign n83795 = ~n83744 & n83762;
  assign n83796 = ~n83770 & n83795;
  assign n83797 = ~n83750 & ~n83756;
  assign n83798 = n83770 & n83772;
  assign n83799 = ~n83797 & ~n83798;
  assign n83800 = ~n83744 & ~n83799;
  assign n83801 = ~n83796 & ~n83800;
  assign n83802 = n83756 & n83762;
  assign n83803 = ~n83750 & n83802;
  assign n83804 = ~n83770 & n83803;
  assign n83805 = n83801 & ~n83804;
  assign n83806 = n83762 & n83797;
  assign n83807 = n83770 & n83806;
  assign n83808 = n83805 & ~n83807;
  assign n83809 = ~n83794 & n83808;
  assign n83810 = ~n83789 & ~n83809;
  assign n83811 = n83750 & n83762;
  assign n83812 = ~n83744 & n83770;
  assign n83813 = n83789 & n83812;
  assign n83814 = n83811 & n83813;
  assign n83815 = n83750 & ~n83770;
  assign n83816 = ~n83762 & n83815;
  assign n83817 = ~n83744 & ~n83816;
  assign n83818 = n83756 & n83776;
  assign n83819 = ~n83763 & ~n83811;
  assign n83820 = ~n83770 & ~n83819;
  assign n83821 = ~n83750 & n83772;
  assign n83822 = n83744 & ~n83821;
  assign n83823 = ~n83820 & n83822;
  assign n83824 = ~n83818 & n83823;
  assign n83825 = ~n83817 & ~n83824;
  assign n83826 = ~n83762 & n83776;
  assign n83827 = ~n83756 & n83826;
  assign n83828 = ~n83825 & ~n83827;
  assign n83829 = n83789 & ~n83828;
  assign n83830 = ~n83814 & ~n83829;
  assign n83831 = ~n83810 & n83830;
  assign n83832 = ~n83783 & n83831;
  assign n83833 = ~n83744 & n83804;
  assign n83834 = n83832 & ~n83833;
  assign n83835 = pi2658 & ~n83834;
  assign n83836 = ~pi2658 & ~n83833;
  assign n83837 = n83832 & n83836;
  assign po2791 = n83835 | n83837;
  assign n83839 = n83661 & n83667;
  assign n83840 = n83655 & n83839;
  assign n83841 = ~n83649 & n83840;
  assign n83842 = ~n83649 & n83696;
  assign n83843 = ~n83655 & n83839;
  assign n83844 = n83649 & n83843;
  assign n83845 = ~n83842 & ~n83844;
  assign n83846 = ~n83643 & ~n83845;
  assign n83847 = ~n83841 & ~n83846;
  assign n83848 = n83643 & n83839;
  assign n83849 = ~n83649 & n83848;
  assign n83850 = ~n83717 & ~n83849;
  assign n83851 = n83847 & n83850;
  assign n83852 = ~n83649 & n83685;
  assign n83853 = n83649 & n83723;
  assign n83854 = ~n83852 & ~n83853;
  assign n83855 = n83851 & n83854;
  assign n83856 = n83681 & ~n83855;
  assign n83857 = ~n83643 & ~n83681;
  assign n83858 = ~n83655 & ~n83661;
  assign n83859 = ~n83649 & ~n83655;
  assign n83860 = n83667 & n83859;
  assign n83861 = ~n83858 & ~n83860;
  assign n83862 = n83857 & ~n83861;
  assign n83863 = ~n83684 & ~n83689;
  assign n83864 = n83655 & n83714;
  assign n83865 = ~n83839 & n83864;
  assign n83866 = ~n83686 & ~n83865;
  assign n83867 = n83863 & n83866;
  assign n83868 = ~n83681 & ~n83867;
  assign n83869 = ~n83643 & n83672;
  assign n83870 = n83649 & n83869;
  assign n83871 = n83649 & n83697;
  assign n83872 = ~n83853 & ~n83871;
  assign n83873 = ~n83643 & ~n83872;
  assign n83874 = ~n83870 & ~n83873;
  assign n83875 = n83643 & n83684;
  assign n83876 = n83874 & ~n83875;
  assign n83877 = ~n83868 & n83876;
  assign n83878 = ~n83862 & n83877;
  assign n83879 = ~n83856 & n83878;
  assign n83880 = n83708 & n83720;
  assign n83881 = n83879 & ~n83880;
  assign n83882 = ~pi2660 & ~n83881;
  assign n83883 = pi2660 & ~n83880;
  assign n83884 = n83878 & n83883;
  assign n83885 = ~n83856 & n83884;
  assign po2793 = n83882 | n83885;
  assign n83887 = n83547 & n83579;
  assign n83888 = ~n83560 & ~n83623;
  assign n83889 = n83541 & ~n83888;
  assign n83890 = ~n83887 & ~n83889;
  assign n83891 = ~n83619 & n83890;
  assign n83892 = ~n83541 & n83612;
  assign n83893 = ~n83602 & ~n83892;
  assign n83894 = ~n83611 & n83893;
  assign n83895 = n83891 & n83894;
  assign n83896 = n83571 & ~n83895;
  assign n83897 = ~n83553 & n83592;
  assign n83898 = n83547 & n83897;
  assign n83899 = ~n83590 & ~n83898;
  assign n83900 = ~n83547 & n83610;
  assign n83901 = ~n83580 & ~n83900;
  assign n83902 = n83553 & n83577;
  assign n83903 = n83547 & ~n83559;
  assign n83904 = ~n83902 & ~n83903;
  assign n83905 = ~n83606 & n83904;
  assign n83906 = ~n83541 & ~n83905;
  assign n83907 = ~n83553 & n83581;
  assign n83908 = n83541 & n83907;
  assign n83909 = n83547 & n83601;
  assign n83910 = ~n83908 & ~n83909;
  assign n83911 = ~n83906 & n83910;
  assign n83912 = n83901 & n83911;
  assign n83913 = n83899 & n83912;
  assign n83914 = ~n83571 & ~n83913;
  assign n83915 = ~n83896 & ~n83914;
  assign n83916 = pi2657 & ~n83915;
  assign n83917 = ~pi2657 & ~n83896;
  assign n83918 = ~n83914 & n83917;
  assign po2794 = n83916 | n83918;
  assign n83920 = ~n83710 & ~n83716;
  assign n83921 = ~n83649 & n83843;
  assign n83922 = ~n83698 & ~n83921;
  assign n83923 = ~n83670 & n83922;
  assign n83924 = ~n83643 & ~n83923;
  assign n83925 = ~n83672 & ~n83684;
  assign n83926 = ~n83726 & n83925;
  assign n83927 = ~n83643 & ~n83926;
  assign n83928 = ~n83880 & n83922;
  assign n83929 = n83643 & n83723;
  assign n83930 = n83928 & ~n83929;
  assign n83931 = ~n83927 & n83930;
  assign n83932 = n83681 & ~n83931;
  assign n83933 = ~n83667 & n83682;
  assign n83934 = ~n83724 & ~n83933;
  assign n83935 = ~n83643 & n83696;
  assign n83936 = n83649 & n83935;
  assign n83937 = ~n83643 & n83669;
  assign n83938 = ~n83936 & ~n83937;
  assign n83939 = n83649 & n83848;
  assign n83940 = ~n83667 & n83859;
  assign n83941 = ~n83672 & ~n83940;
  assign n83942 = n83643 & ~n83941;
  assign n83943 = ~n83939 & ~n83942;
  assign n83944 = n83938 & n83943;
  assign n83945 = ~n83670 & n83944;
  assign n83946 = n83934 & n83945;
  assign n83947 = ~n83681 & ~n83946;
  assign n83948 = ~n83932 & ~n83947;
  assign n83949 = ~n83924 & n83948;
  assign n83950 = n83920 & n83949;
  assign n83951 = pi2664 & ~n83950;
  assign n83952 = ~pi2664 & n83950;
  assign po2795 = n83951 | n83952;
  assign n83954 = ~n83547 & n83592;
  assign n83955 = ~n83900 & ~n83954;
  assign n83956 = n83541 & n83955;
  assign n83957 = n83547 & n83562;
  assign n83958 = ~n83578 & ~n83581;
  assign n83959 = n83553 & ~n83958;
  assign n83960 = n83559 & n83617;
  assign n83961 = n83547 & n83578;
  assign n83962 = ~n83960 & ~n83961;
  assign n83963 = ~n83541 & n83962;
  assign n83964 = ~n83959 & n83963;
  assign n83965 = ~n83957 & n83964;
  assign n83966 = ~n83956 & ~n83965;
  assign n83967 = n83547 & n83959;
  assign n83968 = ~n83898 & ~n83967;
  assign n83969 = ~n83966 & n83968;
  assign n83970 = n83571 & ~n83969;
  assign n83971 = n83541 & ~n83958;
  assign n83972 = ~n83547 & n83971;
  assign n83973 = ~n83599 & ~n83609;
  assign n83974 = n83547 & ~n83973;
  assign n83975 = n83541 & n83974;
  assign n83976 = ~n83553 & n83971;
  assign n83977 = ~n83975 & ~n83976;
  assign n83978 = ~n83972 & n83977;
  assign n83979 = ~n83571 & ~n83978;
  assign n83980 = ~n83970 & ~n83979;
  assign n83981 = ~n83541 & ~n83955;
  assign n83982 = ~n83590 & ~n83981;
  assign n83983 = ~n83571 & ~n83982;
  assign n83984 = n83541 & n83590;
  assign n83985 = ~n83541 & ~n83968;
  assign n83986 = ~n83984 & ~n83985;
  assign n83987 = ~n83983 & n83986;
  assign n83988 = n83980 & n83987;
  assign n83989 = pi2666 & ~n83988;
  assign n83990 = ~pi2666 & n83987;
  assign n83991 = ~n83979 & n83990;
  assign n83992 = ~n83970 & n83991;
  assign po2796 = n83989 | n83992;
  assign n83994 = pi5743 & ~pi9040;
  assign n83995 = pi5933 & pi9040;
  assign n83996 = ~n83994 & ~n83995;
  assign n83997 = ~pi2632 & ~n83996;
  assign n83998 = pi2632 & n83996;
  assign n83999 = ~n83997 & ~n83998;
  assign n84000 = pi5723 & pi9040;
  assign n84001 = pi5807 & ~pi9040;
  assign n84002 = ~n84000 & ~n84001;
  assign n84003 = ~pi2626 & ~n84002;
  assign n84004 = pi2626 & n84002;
  assign n84005 = ~n84003 & ~n84004;
  assign n84006 = pi5797 & ~pi9040;
  assign n84007 = pi6016 & pi9040;
  assign n84008 = ~n84006 & ~n84007;
  assign n84009 = ~pi2647 & ~n84008;
  assign n84010 = pi2647 & n84008;
  assign n84011 = ~n84009 & ~n84010;
  assign n84012 = pi5839 & pi9040;
  assign n84013 = pi6036 & ~pi9040;
  assign n84014 = ~n84012 & ~n84013;
  assign n84015 = ~pi2624 & n84014;
  assign n84016 = pi2624 & ~n84014;
  assign n84017 = ~n84015 & ~n84016;
  assign n84018 = ~n84011 & ~n84017;
  assign n84019 = pi5883 & pi9040;
  assign n84020 = pi6146 & ~pi9040;
  assign n84021 = ~n84019 & ~n84020;
  assign n84022 = ~pi2633 & n84021;
  assign n84023 = pi2633 & ~n84021;
  assign n84024 = ~n84022 & ~n84023;
  assign n84025 = pi6045 & pi9040;
  assign n84026 = pi5933 & ~pi9040;
  assign n84027 = ~n84025 & ~n84026;
  assign n84028 = ~pi2648 & n84027;
  assign n84029 = pi2648 & ~n84027;
  assign n84030 = ~n84028 & ~n84029;
  assign n84031 = ~n84024 & ~n84030;
  assign n84032 = n84018 & n84031;
  assign n84033 = n84005 & n84032;
  assign n84034 = n84024 & ~n84030;
  assign n84035 = n84011 & ~n84017;
  assign n84036 = n84034 & n84035;
  assign n84037 = n84011 & n84017;
  assign n84038 = n84005 & n84037;
  assign n84039 = ~n84030 & n84038;
  assign n84040 = ~n84024 & n84039;
  assign n84041 = n84005 & n84024;
  assign n84042 = n84017 & n84041;
  assign n84043 = ~n84011 & n84042;
  assign n84044 = ~n84040 & ~n84043;
  assign n84045 = ~n84036 & n84044;
  assign n84046 = ~n84033 & n84045;
  assign n84047 = ~n84005 & n84024;
  assign n84048 = ~n84017 & n84047;
  assign n84049 = n84011 & n84048;
  assign n84050 = n84046 & ~n84049;
  assign n84051 = ~n83999 & ~n84050;
  assign n84052 = n84005 & n84011;
  assign n84053 = ~n84017 & n84052;
  assign n84054 = ~n84024 & n84053;
  assign n84055 = ~n84042 & ~n84054;
  assign n84056 = ~n84005 & n84018;
  assign n84057 = ~n84024 & n84056;
  assign n84058 = n84055 & ~n84057;
  assign n84059 = n84030 & ~n84058;
  assign n84060 = ~n84005 & n84017;
  assign n84061 = n84011 & n84060;
  assign n84062 = n84030 & n84061;
  assign n84063 = ~n84024 & n84062;
  assign n84064 = ~n84011 & n84041;
  assign n84065 = ~n84011 & n84017;
  assign n84066 = n84024 & n84065;
  assign n84067 = ~n84064 & ~n84066;
  assign n84068 = n84030 & ~n84067;
  assign n84069 = ~n84063 & ~n84068;
  assign n84070 = ~n83999 & ~n84069;
  assign n84071 = ~n84059 & ~n84070;
  assign n84072 = ~n84051 & n84071;
  assign n84073 = ~n84005 & ~n84024;
  assign n84074 = ~n84030 & n84073;
  assign n84075 = n84065 & n84074;
  assign n84076 = ~n84005 & n84011;
  assign n84077 = n84034 & n84076;
  assign n84078 = n84024 & n84061;
  assign n84079 = n84005 & n84030;
  assign n84080 = n84011 & n84079;
  assign n84081 = ~n84011 & ~n84024;
  assign n84082 = ~n84005 & n84081;
  assign n84083 = ~n84080 & ~n84082;
  assign n84084 = ~n84078 & n84083;
  assign n84085 = ~n84056 & n84084;
  assign n84086 = n84018 & ~n84030;
  assign n84087 = n84024 & n84086;
  assign n84088 = ~n84024 & n84065;
  assign n84089 = ~n84005 & ~n84017;
  assign n84090 = ~n84088 & ~n84089;
  assign n84091 = ~n84030 & ~n84090;
  assign n84092 = ~n84087 & ~n84091;
  assign n84093 = n84085 & n84092;
  assign n84094 = n83999 & ~n84093;
  assign n84095 = ~n84077 & ~n84094;
  assign n84096 = ~n84075 & n84095;
  assign n84097 = n84072 & n84096;
  assign n84098 = pi2661 & n84097;
  assign n84099 = ~pi2661 & ~n84097;
  assign po2799 = n84098 | n84099;
  assign n84101 = ~n83852 & ~n83860;
  assign n84102 = n83681 & ~n84101;
  assign n84103 = ~n83683 & ~n83690;
  assign n84104 = ~n83840 & n84103;
  assign n84105 = ~n83643 & ~n84104;
  assign n84106 = n83681 & n84105;
  assign n84107 = ~n84102 & ~n84106;
  assign n84108 = n83685 & n83693;
  assign n84109 = ~n83695 & ~n84108;
  assign n84110 = ~n83689 & ~n83727;
  assign n84111 = n83643 & ~n84110;
  assign n84112 = n83681 & n84111;
  assign n84113 = n84109 & ~n84112;
  assign n84114 = n83649 & n83685;
  assign n84115 = n83649 & n83668;
  assign n84116 = ~n83673 & ~n84115;
  assign n84117 = n83643 & ~n84116;
  assign n84118 = ~n83684 & ~n83698;
  assign n84119 = n83649 & n83671;
  assign n84120 = ~n83720 & ~n84119;
  assign n84121 = ~n83643 & ~n84120;
  assign n84122 = n84118 & ~n84121;
  assign n84123 = ~n84117 & n84122;
  assign n84124 = ~n84114 & n84123;
  assign n84125 = ~n83681 & ~n84124;
  assign n84126 = ~n83724 & n83922;
  assign n84127 = n83643 & ~n84126;
  assign n84128 = ~n84125 & ~n84127;
  assign n84129 = n84113 & n84128;
  assign n84130 = n84107 & n84129;
  assign n84131 = ~pi2678 & ~n84130;
  assign n84132 = pi2678 & n84113;
  assign n84133 = n84107 & n84132;
  assign n84134 = n84128 & n84133;
  assign po2800 = n84131 | n84134;
  assign n84136 = n83367 & ~n83373;
  assign n84137 = n83385 & n84136;
  assign n84138 = n83379 & n83398;
  assign n84139 = n83373 & n84138;
  assign n84140 = n83392 & n83433;
  assign n84141 = ~n84139 & ~n84140;
  assign n84142 = ~n83373 & ~n83379;
  assign n84143 = ~n83391 & n84142;
  assign n84144 = ~n83385 & n84143;
  assign n84145 = ~n83415 & ~n84144;
  assign n84146 = ~n83367 & ~n84145;
  assign n84147 = n84141 & ~n84146;
  assign n84148 = ~n84137 & n84147;
  assign n84149 = n83412 & ~n84148;
  assign n84150 = n83373 & n83444;
  assign n84151 = n83367 & n84150;
  assign n84152 = ~n83367 & ~n83373;
  assign n84153 = n83444 & n84152;
  assign n84154 = ~n83413 & ~n84153;
  assign n84155 = ~n83415 & ~n83436;
  assign n84156 = ~n83373 & n83392;
  assign n84157 = n84155 & ~n84156;
  assign n84158 = n83367 & ~n84157;
  assign n84159 = ~n83367 & n83419;
  assign n84160 = n83401 & ~n84159;
  assign n84161 = ~n84158 & n84160;
  assign n84162 = n84154 & n84161;
  assign n84163 = ~n83412 & ~n84162;
  assign n84164 = ~n84151 & ~n84163;
  assign n84165 = ~n84149 & n84164;
  assign n84166 = n83436 & n84152;
  assign n84167 = n83373 & n83438;
  assign n84168 = ~n84166 & ~n84167;
  assign n84169 = ~n83367 & n84140;
  assign n84170 = n84168 & ~n84169;
  assign n84171 = n84165 & n84170;
  assign n84172 = ~pi2673 & ~n84171;
  assign n84173 = pi2673 & n84170;
  assign n84174 = n84164 & n84173;
  assign n84175 = ~n84149 & n84174;
  assign po2801 = n84172 | n84175;
  assign n84177 = n84024 & n84038;
  assign n84178 = n84024 & n84056;
  assign n84179 = ~n84177 & ~n84178;
  assign n84180 = n84030 & ~n84179;
  assign n84181 = ~n84024 & n84030;
  assign n84182 = n84053 & n84181;
  assign n84183 = ~n84180 & ~n84182;
  assign n84184 = ~n84077 & n84183;
  assign n84185 = ~n84024 & n84061;
  assign n84186 = ~n84056 & ~n84185;
  assign n84187 = n84005 & n84065;
  assign n84188 = n84186 & ~n84187;
  assign n84189 = n83999 & ~n84188;
  assign n84190 = n84030 & n84189;
  assign n84191 = n84005 & ~n84030;
  assign n84192 = n84017 & n84191;
  assign n84193 = ~n84011 & n84192;
  assign n84194 = n84024 & n84193;
  assign n84195 = n84005 & n84018;
  assign n84196 = ~n84030 & n84195;
  assign n84197 = ~n84049 & ~n84075;
  assign n84198 = ~n84040 & n84197;
  assign n84199 = ~n84196 & n84198;
  assign n84200 = n83999 & ~n84199;
  assign n84201 = ~n84194 & ~n84200;
  assign n84202 = n84005 & ~n84024;
  assign n84203 = ~n84017 & n84202;
  assign n84204 = ~n84024 & n84086;
  assign n84205 = ~n84193 & ~n84204;
  assign n84206 = ~n84203 & n84205;
  assign n84207 = n84017 & n84047;
  assign n84208 = ~n84024 & n84035;
  assign n84209 = ~n84052 & ~n84208;
  assign n84210 = n84030 & ~n84209;
  assign n84211 = ~n84207 & ~n84210;
  assign n84212 = n84206 & n84211;
  assign n84213 = ~n83999 & ~n84212;
  assign n84214 = n84201 & ~n84213;
  assign n84215 = ~n84190 & n84214;
  assign n84216 = n84184 & n84215;
  assign n84217 = pi2667 & ~n84216;
  assign n84218 = ~pi2667 & n84184;
  assign n84219 = n84215 & n84218;
  assign po2802 = n84217 | n84219;
  assign n84221 = n83547 & n83907;
  assign n84222 = n83541 & n84221;
  assign n84223 = n83617 & ~n83958;
  assign n84224 = ~n83610 & ~n84223;
  assign n84225 = ~n83898 & n84224;
  assign n84226 = ~n83541 & ~n84225;
  assign n84227 = n83547 & n83587;
  assign n84228 = ~n84226 & ~n84227;
  assign n84229 = ~n83553 & n83609;
  assign n84230 = ~n83547 & n83902;
  assign n84231 = ~n84229 & ~n84230;
  assign n84232 = ~n83961 & n84231;
  assign n84233 = n83541 & ~n84232;
  assign n84234 = n84228 & ~n84233;
  assign n84235 = n83571 & ~n84234;
  assign n84236 = ~n84222 & ~n84235;
  assign n84237 = ~n83547 & n83578;
  assign n84238 = ~n83897 & ~n84237;
  assign n84239 = n83541 & ~n84238;
  assign n84240 = ~n83611 & ~n84239;
  assign n84241 = ~n83600 & ~n84221;
  assign n84242 = n83547 & n83606;
  assign n84243 = ~n83902 & ~n84242;
  assign n84244 = ~n84229 & n84243;
  assign n84245 = ~n83541 & ~n84244;
  assign n84246 = ~n83547 & n83587;
  assign n84247 = ~n84245 & ~n84246;
  assign n84248 = n84241 & n84247;
  assign n84249 = n84240 & n84248;
  assign n84250 = ~n83571 & ~n84249;
  assign n84251 = ~n83626 & ~n83957;
  assign n84252 = ~n83541 & ~n84251;
  assign n84253 = ~n84250 & ~n84252;
  assign n84254 = n84236 & n84253;
  assign n84255 = pi2665 & n84254;
  assign n84256 = ~pi2665 & ~n84254;
  assign po2805 = n84255 | n84256;
  assign n84258 = pi5723 & ~pi9040;
  assign n84259 = pi5951 & pi9040;
  assign n84260 = ~n84258 & ~n84259;
  assign n84261 = pi2616 & n84260;
  assign n84262 = ~pi2616 & ~n84260;
  assign n84263 = ~n84261 & ~n84262;
  assign n84264 = pi5884 & pi9040;
  assign n84265 = pi5735 & ~pi9040;
  assign n84266 = ~n84264 & ~n84265;
  assign n84267 = ~pi2617 & n84266;
  assign n84268 = pi2617 & ~n84266;
  assign n84269 = ~n84267 & ~n84268;
  assign n84270 = pi6045 & ~pi9040;
  assign n84271 = pi5797 & pi9040;
  assign n84272 = ~n84270 & ~n84271;
  assign n84273 = ~pi2636 & ~n84272;
  assign n84274 = pi2636 & n84272;
  assign n84275 = ~n84273 & ~n84274;
  assign n84276 = pi5803 & pi9040;
  assign n84277 = pi6033 & ~pi9040;
  assign n84278 = ~n84276 & ~n84277;
  assign n84279 = ~pi2628 & n84278;
  assign n84280 = pi2628 & ~n84278;
  assign n84281 = ~n84279 & ~n84280;
  assign n84282 = pi5874 & ~pi9040;
  assign n84283 = pi5844 & pi9040;
  assign n84284 = ~n84282 & ~n84283;
  assign n84285 = ~pi2643 & ~n84284;
  assign n84286 = pi2643 & n84284;
  assign n84287 = ~n84285 & ~n84286;
  assign n84288 = n84281 & n84287;
  assign n84289 = n84275 & n84288;
  assign n84290 = ~n84269 & n84289;
  assign n84291 = ~n84263 & n84290;
  assign n84292 = ~n84281 & ~n84287;
  assign n84293 = ~n84263 & ~n84269;
  assign n84294 = n84292 & n84293;
  assign n84295 = ~n84275 & n84294;
  assign n84296 = ~n84291 & ~n84295;
  assign n84297 = ~n84275 & n84288;
  assign n84298 = ~n84263 & n84269;
  assign n84299 = n84297 & n84298;
  assign n84300 = ~n84275 & n84292;
  assign n84301 = ~n84263 & n84300;
  assign n84302 = ~n84299 & ~n84301;
  assign n84303 = n84275 & ~n84281;
  assign n84304 = n84263 & n84303;
  assign n84305 = n84263 & n84288;
  assign n84306 = ~n84304 & ~n84305;
  assign n84307 = ~n84269 & ~n84306;
  assign n84308 = ~n84281 & n84287;
  assign n84309 = n84281 & ~n84287;
  assign n84310 = ~n84308 & ~n84309;
  assign n84311 = ~n84263 & ~n84275;
  assign n84312 = n84269 & ~n84311;
  assign n84313 = ~n84310 & n84312;
  assign n84314 = ~n84263 & ~n84288;
  assign n84315 = ~n84269 & n84314;
  assign n84316 = ~n84275 & n84315;
  assign n84317 = ~n84313 & ~n84316;
  assign n84318 = ~n84307 & n84317;
  assign n84319 = n84302 & n84318;
  assign n84320 = pi5801 & pi9040;
  assign n84321 = pi5806 & ~pi9040;
  assign n84322 = ~n84320 & ~n84321;
  assign n84323 = pi2637 & n84322;
  assign n84324 = ~pi2637 & ~n84322;
  assign n84325 = ~n84323 & ~n84324;
  assign n84326 = ~n84319 & n84325;
  assign n84327 = n84296 & ~n84326;
  assign n84328 = n84275 & n84308;
  assign n84329 = n84269 & n84328;
  assign n84330 = n84263 & n84329;
  assign n84331 = n84269 & ~n84325;
  assign n84332 = n84275 & n84292;
  assign n84333 = ~n84305 & ~n84332;
  assign n84334 = ~n84310 & n84311;
  assign n84335 = n84333 & ~n84334;
  assign n84336 = n84331 & ~n84335;
  assign n84337 = n84263 & n84300;
  assign n84338 = n84263 & ~n84281;
  assign n84339 = ~n84275 & n84338;
  assign n84340 = n84263 & n84309;
  assign n84341 = ~n84339 & ~n84340;
  assign n84342 = ~n84263 & n84288;
  assign n84343 = n84275 & n84309;
  assign n84344 = ~n84342 & ~n84343;
  assign n84345 = n84341 & n84344;
  assign n84346 = ~n84269 & ~n84345;
  assign n84347 = ~n84337 & ~n84346;
  assign n84348 = ~n84325 & ~n84347;
  assign n84349 = ~n84336 & ~n84348;
  assign n84350 = ~n84330 & n84349;
  assign n84351 = n84327 & n84350;
  assign n84352 = pi2688 & ~n84351;
  assign n84353 = ~pi2688 & n84327;
  assign n84354 = n84350 & n84353;
  assign po2806 = n84352 | n84354;
  assign n84356 = ~n84340 & ~n84342;
  assign n84357 = ~n84269 & ~n84356;
  assign n84358 = ~n84295 & ~n84357;
  assign n84359 = n84325 & ~n84358;
  assign n84360 = ~n84275 & ~n84281;
  assign n84361 = ~n84308 & ~n84360;
  assign n84362 = ~n84263 & ~n84361;
  assign n84363 = ~n84289 & ~n84362;
  assign n84364 = n84269 & ~n84363;
  assign n84365 = ~n84334 & ~n84364;
  assign n84366 = n84263 & n84297;
  assign n84367 = ~n84263 & n84275;
  assign n84368 = ~n84287 & n84367;
  assign n84369 = n84263 & ~n84361;
  assign n84370 = ~n84368 & ~n84369;
  assign n84371 = ~n84269 & ~n84370;
  assign n84372 = ~n84366 & ~n84371;
  assign n84373 = n84365 & n84372;
  assign n84374 = ~n84325 & ~n84373;
  assign n84375 = n84263 & n84275;
  assign n84376 = ~n84308 & n84375;
  assign n84377 = n84325 & n84376;
  assign n84378 = n84263 & ~n84275;
  assign n84379 = n84308 & n84378;
  assign n84380 = ~n84269 & n84379;
  assign n84381 = n84263 & n84269;
  assign n84382 = n84275 & n84381;
  assign n84383 = ~n84287 & n84382;
  assign n84384 = ~n84380 & ~n84383;
  assign n84385 = ~n84377 & n84384;
  assign n84386 = ~n84338 & ~n84343;
  assign n84387 = n84269 & n84325;
  assign n84388 = ~n84386 & n84387;
  assign n84389 = n84385 & ~n84388;
  assign n84390 = ~n84374 & n84389;
  assign n84391 = ~n84359 & n84390;
  assign n84392 = pi2685 & ~n84391;
  assign n84393 = ~pi2685 & n84391;
  assign po2807 = n84392 | n84393;
  assign n84395 = pi5883 & ~pi9040;
  assign n84396 = pi5743 & pi9040;
  assign n84397 = ~n84395 & ~n84396;
  assign n84398 = pi2642 & n84397;
  assign n84399 = ~pi2642 & ~n84397;
  assign n84400 = ~n84398 & ~n84399;
  assign n84401 = pi5806 & pi9040;
  assign n84402 = pi5844 & ~pi9040;
  assign n84403 = ~n84401 & ~n84402;
  assign n84404 = ~pi2632 & ~n84403;
  assign n84405 = pi2632 & n84403;
  assign n84406 = ~n84404 & ~n84405;
  assign n84407 = pi6036 & pi9040;
  assign n84408 = pi5877 & ~pi9040;
  assign n84409 = ~n84407 & ~n84408;
  assign n84410 = pi2636 & n84409;
  assign n84411 = ~pi2636 & ~n84409;
  assign n84412 = ~n84410 & ~n84411;
  assign n84413 = n84406 & ~n84412;
  assign n84414 = pi6002 & ~pi9040;
  assign n84415 = pi5877 & pi9040;
  assign n84416 = ~n84414 & ~n84415;
  assign n84417 = ~pi2646 & ~n84416;
  assign n84418 = pi2646 & n84416;
  assign n84419 = ~n84417 & ~n84418;
  assign n84420 = pi5839 & ~pi9040;
  assign n84421 = pi6033 & pi9040;
  assign n84422 = ~n84420 & ~n84421;
  assign n84423 = pi2624 & n84422;
  assign n84424 = ~pi2624 & ~n84422;
  assign n84425 = ~n84423 & ~n84424;
  assign n84426 = n84419 & n84425;
  assign n84427 = n84413 & n84426;
  assign n84428 = n84419 & ~n84425;
  assign n84429 = ~n84406 & n84428;
  assign n84430 = ~n84427 & ~n84429;
  assign n84431 = ~n84400 & ~n84430;
  assign n84432 = pi5801 & ~pi9040;
  assign n84433 = pi5799 & pi9040;
  assign n84434 = ~n84432 & ~n84433;
  assign n84435 = ~pi2628 & ~n84434;
  assign n84436 = pi2628 & n84434;
  assign n84437 = ~n84435 & ~n84436;
  assign n84438 = n84400 & ~n84419;
  assign n84439 = n84406 & n84438;
  assign n84440 = n84413 & ~n84425;
  assign n84441 = n84406 & n84412;
  assign n84442 = n84425 & n84441;
  assign n84443 = ~n84440 & ~n84442;
  assign n84444 = ~n84406 & ~n84412;
  assign n84445 = n84425 & n84444;
  assign n84446 = n84419 & n84445;
  assign n84447 = n84443 & ~n84446;
  assign n84448 = n84400 & ~n84447;
  assign n84449 = ~n84439 & ~n84448;
  assign n84450 = ~n84406 & n84412;
  assign n84451 = ~n84425 & n84450;
  assign n84452 = n84419 & n84451;
  assign n84453 = n84449 & ~n84452;
  assign n84454 = ~n84419 & n84444;
  assign n84455 = n84425 & n84450;
  assign n84456 = ~n84454 & ~n84455;
  assign n84457 = ~n84400 & ~n84456;
  assign n84458 = ~n84425 & n84441;
  assign n84459 = ~n84419 & n84458;
  assign n84460 = ~n84457 & ~n84459;
  assign n84461 = n84453 & n84460;
  assign n84462 = n84437 & ~n84461;
  assign n84463 = ~n84431 & ~n84462;
  assign n84464 = n84400 & ~n84437;
  assign n84465 = ~n84456 & n84464;
  assign n84466 = ~n84425 & n84444;
  assign n84467 = ~n84458 & ~n84466;
  assign n84468 = n84419 & ~n84467;
  assign n84469 = ~n84427 & ~n84468;
  assign n84470 = ~n84437 & ~n84469;
  assign n84471 = ~n84465 & ~n84470;
  assign n84472 = ~n84400 & ~n84437;
  assign n84473 = n84413 & ~n84419;
  assign n84474 = ~n84451 & ~n84473;
  assign n84475 = n84406 & n84425;
  assign n84476 = n84474 & ~n84475;
  assign n84477 = n84472 & ~n84476;
  assign n84478 = n84471 & ~n84477;
  assign n84479 = n84463 & n84478;
  assign n84480 = ~pi2659 & ~n84479;
  assign n84481 = pi2659 & n84471;
  assign n84482 = n84463 & n84481;
  assign n84483 = ~n84477 & n84482;
  assign po2808 = n84480 | n84483;
  assign n84485 = ~n83373 & n84138;
  assign n84486 = ~n83393 & ~n83406;
  assign n84487 = n83373 & n83395;
  assign n84488 = ~n83373 & n83444;
  assign n84489 = ~n84487 & ~n84488;
  assign n84490 = n84486 & n84489;
  assign n84491 = n83367 & ~n84490;
  assign n84492 = n83373 & n83414;
  assign n84493 = ~n83413 & ~n84492;
  assign n84494 = ~n83399 & n84493;
  assign n84495 = ~n83367 & ~n84494;
  assign n84496 = n83391 & n83433;
  assign n84497 = n83385 & n84496;
  assign n84498 = ~n84495 & ~n84497;
  assign n84499 = ~n84491 & n84498;
  assign n84500 = ~n84485 & n84499;
  assign n84501 = ~n83412 & ~n84500;
  assign n84502 = n83367 & n83373;
  assign n84503 = n83419 & n84502;
  assign n84504 = n83367 & n83399;
  assign n84505 = n83367 & n83436;
  assign n84506 = ~n84504 & ~n84505;
  assign n84507 = ~n83373 & ~n84506;
  assign n84508 = ~n84503 & ~n84507;
  assign n84509 = n83373 & n83392;
  assign n84510 = ~n83373 & n83414;
  assign n84511 = ~n84509 & ~n84510;
  assign n84512 = ~n83396 & n84511;
  assign n84513 = ~n83393 & n84512;
  assign n84514 = ~n83367 & ~n84513;
  assign n84515 = ~n83373 & n83415;
  assign n84516 = ~n84514 & ~n84515;
  assign n84517 = ~n83373 & n83396;
  assign n84518 = ~n84150 & ~n84517;
  assign n84519 = n84516 & n84518;
  assign n84520 = n84508 & n84519;
  assign n84521 = n83412 & ~n84520;
  assign n84522 = n83367 & ~n84141;
  assign n84523 = ~n84521 & ~n84522;
  assign n84524 = ~n83400 & ~n84517;
  assign n84525 = ~n83367 & ~n84524;
  assign n84526 = n84523 & ~n84525;
  assign n84527 = ~n84501 & n84526;
  assign n84528 = pi2681 & ~n84527;
  assign n84529 = ~pi2681 & n84527;
  assign po2809 = n84528 | n84529;
  assign n84531 = n84005 & ~n84011;
  assign n84532 = ~n84049 & ~n84531;
  assign n84533 = ~n84081 & n84532;
  assign n84534 = ~n84030 & ~n84533;
  assign n84535 = n84011 & n84181;
  assign n84536 = ~n84177 & ~n84203;
  assign n84537 = ~n84005 & ~n84011;
  assign n84538 = n84024 & n84030;
  assign n84539 = n84537 & n84538;
  assign n84540 = n84536 & ~n84539;
  assign n84541 = ~n84535 & n84540;
  assign n84542 = ~n84534 & n84541;
  assign n84543 = n83999 & ~n84542;
  assign n84544 = n84024 & n84195;
  assign n84545 = ~n84024 & n84187;
  assign n84546 = ~n84544 & ~n84545;
  assign n84547 = ~n84030 & ~n84546;
  assign n84548 = ~n84543 & ~n84547;
  assign n84549 = ~n84024 & n84038;
  assign n84550 = ~n84053 & ~n84061;
  assign n84551 = ~n84030 & ~n84550;
  assign n84552 = ~n84549 & ~n84551;
  assign n84553 = ~n84057 & n84552;
  assign n84554 = ~n83999 & ~n84553;
  assign n84555 = ~n84035 & ~n84065;
  assign n84556 = ~n84005 & ~n84555;
  assign n84557 = ~n84066 & ~n84556;
  assign n84558 = n84030 & ~n84557;
  assign n84559 = ~n83999 & n84558;
  assign n84560 = ~n84554 & ~n84559;
  assign n84561 = n84548 & n84560;
  assign n84562 = pi2662 & ~n84561;
  assign n84563 = ~pi2662 & n84548;
  assign n84564 = n84560 & n84563;
  assign po2810 = n84562 | n84564;
  assign n84566 = ~n84275 & n84308;
  assign n84567 = ~n84289 & ~n84566;
  assign n84568 = ~n84269 & ~n84567;
  assign n84569 = ~n84263 & n84309;
  assign n84570 = ~n84328 & ~n84569;
  assign n84571 = ~n84297 & n84570;
  assign n84572 = n84269 & ~n84571;
  assign n84573 = ~n84568 & ~n84572;
  assign n84574 = ~n84269 & n84332;
  assign n84575 = ~n84275 & n84569;
  assign n84576 = ~n84574 & ~n84575;
  assign n84577 = n84573 & n84576;
  assign n84578 = ~n84325 & ~n84577;
  assign n84579 = n84263 & n84289;
  assign n84580 = ~n84263 & n84292;
  assign n84581 = ~n84340 & ~n84580;
  assign n84582 = n84269 & ~n84581;
  assign n84583 = ~n84579 & ~n84582;
  assign n84584 = ~n84269 & n84275;
  assign n84585 = ~n84287 & n84584;
  assign n84586 = n84281 & n84585;
  assign n84587 = ~n84300 & ~n84328;
  assign n84588 = ~n84586 & n84587;
  assign n84589 = ~n84297 & n84588;
  assign n84590 = ~n84263 & ~n84589;
  assign n84591 = n84583 & ~n84590;
  assign n84592 = n84325 & ~n84591;
  assign n84593 = ~n84578 & ~n84592;
  assign n84594 = n84263 & n84332;
  assign n84595 = ~n84275 & n84340;
  assign n84596 = ~n84594 & ~n84595;
  assign n84597 = ~n84269 & ~n84596;
  assign n84598 = n84269 & n84360;
  assign n84599 = n84263 & n84598;
  assign n84600 = ~n84597 & ~n84599;
  assign n84601 = n84593 & n84600;
  assign n84602 = ~pi2696 & ~n84601;
  assign n84603 = pi2696 & ~n84597;
  assign n84604 = n84593 & n84603;
  assign n84605 = ~n84599 & n84604;
  assign po2811 = n84602 | n84605;
  assign n84607 = ~n84400 & n84419;
  assign n84608 = ~n84444 & ~n84458;
  assign n84609 = n84607 & ~n84608;
  assign n84610 = ~n84400 & ~n84425;
  assign n84611 = n84444 & n84610;
  assign n84612 = ~n84609 & ~n84611;
  assign n84613 = n84437 & ~n84612;
  assign n84614 = ~n84419 & n84442;
  assign n84615 = ~n84419 & n84425;
  assign n84616 = ~n84475 & ~n84615;
  assign n84617 = n84400 & ~n84616;
  assign n84618 = ~n84419 & ~n84425;
  assign n84619 = ~n84412 & n84618;
  assign n84620 = n84406 & n84619;
  assign n84621 = ~n84617 & ~n84620;
  assign n84622 = ~n84614 & n84621;
  assign n84623 = n84437 & ~n84622;
  assign n84624 = ~n84613 & ~n84623;
  assign n84625 = n84412 & n84426;
  assign n84626 = ~n84406 & n84625;
  assign n84627 = ~n84419 & n84451;
  assign n84628 = ~n84626 & ~n84627;
  assign n84629 = ~n84400 & ~n84628;
  assign n84630 = ~n84412 & n84428;
  assign n84631 = ~n84406 & n84630;
  assign n84632 = ~n84419 & n84475;
  assign n84633 = ~n84631 & ~n84632;
  assign n84634 = n84400 & ~n84633;
  assign n84635 = ~n84413 & ~n84475;
  assign n84636 = n84419 & ~n84635;
  assign n84637 = ~n84451 & ~n84636;
  assign n84638 = ~n84400 & ~n84637;
  assign n84639 = n84412 & ~n84419;
  assign n84640 = n84610 & n84639;
  assign n84641 = ~n84412 & n84425;
  assign n84642 = ~n84451 & ~n84641;
  assign n84643 = ~n84419 & ~n84642;
  assign n84644 = n84400 & n84419;
  assign n84645 = n84441 & n84644;
  assign n84646 = ~n84425 & n84645;
  assign n84647 = ~n84643 & ~n84646;
  assign n84648 = ~n84640 & n84647;
  assign n84649 = ~n84638 & n84648;
  assign n84650 = ~n84626 & n84649;
  assign n84651 = ~n84437 & ~n84650;
  assign n84652 = ~n84634 & ~n84651;
  assign n84653 = ~n84629 & n84652;
  assign n84654 = n84624 & n84653;
  assign n84655 = pi2676 & n84654;
  assign n84656 = ~pi2676 & ~n84654;
  assign po2812 = n84655 | n84656;
  assign n84658 = n84287 & n84367;
  assign n84659 = n84587 & ~n84658;
  assign n84660 = n84387 & ~n84659;
  assign n84661 = n84263 & n84325;
  assign n84662 = n84343 & n84661;
  assign n84663 = ~n84275 & n84287;
  assign n84664 = ~n84305 & ~n84663;
  assign n84665 = ~n84269 & ~n84664;
  assign n84666 = ~n84574 & ~n84665;
  assign n84667 = n84325 & ~n84666;
  assign n84668 = ~n84662 & ~n84667;
  assign n84669 = n84287 & n84378;
  assign n84670 = ~n84575 & ~n84669;
  assign n84671 = ~n84269 & ~n84670;
  assign n84672 = n84668 & ~n84671;
  assign n84673 = n84288 & n84381;
  assign n84674 = n84275 & n84673;
  assign n84675 = ~n84310 & n84378;
  assign n84676 = ~n84594 & ~n84675;
  assign n84677 = ~n84310 & n84367;
  assign n84678 = ~n84301 & ~n84677;
  assign n84679 = n84676 & n84678;
  assign n84680 = ~n84299 & n84679;
  assign n84681 = ~n84674 & n84680;
  assign n84682 = n84275 & n84293;
  assign n84683 = n84281 & n84682;
  assign n84684 = n84681 & ~n84683;
  assign n84685 = ~n84325 & ~n84684;
  assign n84686 = n84672 & ~n84685;
  assign n84687 = ~n84660 & n84686;
  assign n84688 = ~pi2682 & ~n84687;
  assign n84689 = pi2682 & n84672;
  assign n84690 = ~n84660 & n84689;
  assign n84691 = ~n84685 & n84690;
  assign po2813 = n84688 | n84691;
  assign n84693 = ~n84419 & n84445;
  assign n84694 = ~n84640 & ~n84693;
  assign n84695 = ~n84458 & ~n84630;
  assign n84696 = ~n84400 & ~n84695;
  assign n84697 = n84419 & n84450;
  assign n84698 = ~n84412 & ~n84419;
  assign n84699 = ~n84425 & n84698;
  assign n84700 = ~n84697 & ~n84699;
  assign n84701 = n84400 & ~n84700;
  assign n84702 = ~n84696 & ~n84701;
  assign n84703 = ~n84427 & n84702;
  assign n84704 = n84694 & n84703;
  assign n84705 = ~n84614 & ~n84626;
  assign n84706 = n84704 & n84705;
  assign n84707 = n84437 & ~n84706;
  assign n84708 = n84413 & n84615;
  assign n84709 = n84467 & ~n84708;
  assign n84710 = n84400 & ~n84709;
  assign n84711 = ~n84419 & n84455;
  assign n84712 = ~n84710 & ~n84711;
  assign n84713 = n84406 & n84428;
  assign n84714 = n84419 & n84441;
  assign n84715 = ~n84713 & ~n84714;
  assign n84716 = n84400 & ~n84715;
  assign n84717 = n84400 & n84450;
  assign n84718 = ~n84419 & n84717;
  assign n84719 = ~n84716 & ~n84718;
  assign n84720 = n84712 & n84719;
  assign n84721 = ~n84437 & ~n84720;
  assign n84722 = ~n84445 & ~n84452;
  assign n84723 = ~n84620 & n84722;
  assign n84724 = n84472 & ~n84723;
  assign n84725 = ~n84721 & ~n84724;
  assign n84726 = ~n84427 & ~n84614;
  assign n84727 = ~n84400 & ~n84726;
  assign n84728 = n84725 & ~n84727;
  assign n84729 = ~n84707 & n84728;
  assign n84730 = ~pi2680 & n84729;
  assign n84731 = pi2680 & ~n84729;
  assign po2814 = n84730 | n84731;
  assign n84733 = ~n83770 & n83806;
  assign n84734 = n83770 & n83811;
  assign n84735 = ~n83803 & ~n84734;
  assign n84736 = n83744 & ~n84735;
  assign n84737 = ~n84733 & ~n84736;
  assign n84738 = ~n83744 & ~n83770;
  assign n84739 = n83762 & n84738;
  assign n84740 = ~n83756 & n84739;
  assign n84741 = n83778 & n83812;
  assign n84742 = ~n84740 & ~n84741;
  assign n84743 = ~n83744 & n83821;
  assign n84744 = n84742 & ~n84743;
  assign n84745 = ~n83774 & ~n83792;
  assign n84746 = ~n83826 & n84745;
  assign n84747 = n84744 & n84746;
  assign n84748 = n84737 & n84747;
  assign n84749 = ~n83789 & ~n84748;
  assign n84750 = n83744 & n83816;
  assign n84751 = ~n83756 & n83815;
  assign n84752 = ~n83750 & n83778;
  assign n84753 = ~n84751 & ~n84752;
  assign n84754 = ~n83750 & n83762;
  assign n84755 = n83770 & n84754;
  assign n84756 = n84753 & ~n84755;
  assign n84757 = n83744 & ~n84756;
  assign n84758 = ~n83770 & n83802;
  assign n84759 = ~n83756 & n83791;
  assign n84760 = ~n84758 & ~n84759;
  assign n84761 = ~n83744 & ~n84760;
  assign n84762 = ~n83770 & n83779;
  assign n84763 = ~n83773 & ~n83803;
  assign n84764 = n83770 & ~n84763;
  assign n84765 = ~n84762 & ~n84764;
  assign n84766 = ~n84761 & n84765;
  assign n84767 = ~n84757 & n84766;
  assign n84768 = ~n84750 & n84767;
  assign n84769 = ~n83789 & ~n84750;
  assign n84770 = ~n84768 & ~n84769;
  assign n84771 = ~n83744 & n84733;
  assign n84772 = ~n84770 & ~n84771;
  assign n84773 = ~n84749 & n84772;
  assign n84774 = ~pi2675 & ~n84773;
  assign n84775 = pi2675 & ~n84770;
  assign n84776 = ~n84749 & n84775;
  assign n84777 = ~n84771 & n84776;
  assign po2815 = n84774 | n84777;
  assign n84779 = ~n84144 & ~n84517;
  assign n84780 = ~n84497 & n84779;
  assign n84781 = n83367 & ~n84780;
  assign n84782 = ~n84153 & ~n84169;
  assign n84783 = ~n84150 & ~n84505;
  assign n84784 = ~n84138 & ~n84510;
  assign n84785 = ~n83367 & ~n84784;
  assign n84786 = ~n83406 & ~n84785;
  assign n84787 = n84783 & n84786;
  assign n84788 = n83412 & ~n84787;
  assign n84789 = ~n83379 & n83391;
  assign n84790 = ~n83420 & ~n84789;
  assign n84791 = n83373 & ~n84790;
  assign n84792 = ~n83396 & ~n84156;
  assign n84793 = ~n83367 & ~n84792;
  assign n84794 = n83373 & n83391;
  assign n84795 = ~n83415 & ~n84794;
  assign n84796 = ~n83398 & n84795;
  assign n84797 = n83367 & ~n84796;
  assign n84798 = ~n84793 & ~n84797;
  assign n84799 = ~n84791 & n84798;
  assign n84800 = ~n83412 & ~n84799;
  assign n84801 = ~n84788 & ~n84800;
  assign n84802 = n84782 & n84801;
  assign n84803 = ~n84781 & n84802;
  assign n84804 = ~pi2689 & ~n84803;
  assign n84805 = pi2689 & n84782;
  assign n84806 = ~n84781 & n84805;
  assign n84807 = n84801 & n84806;
  assign po2816 = n84804 | n84807;
  assign n84809 = ~n84024 & n84556;
  assign n84810 = ~n84060 & ~n84195;
  assign n84811 = n84030 & ~n84810;
  assign n84812 = ~n84809 & ~n84811;
  assign n84813 = n84017 & n84202;
  assign n84814 = ~n84089 & ~n84813;
  assign n84815 = ~n84187 & n84814;
  assign n84816 = ~n84030 & ~n84815;
  assign n84817 = n84812 & ~n84816;
  assign n84818 = n84024 & n84053;
  assign n84819 = n84817 & ~n84818;
  assign n84820 = ~n83999 & ~n84819;
  assign n84821 = ~n84056 & ~n84061;
  assign n84822 = ~n84053 & ~n84187;
  assign n84823 = n84821 & n84822;
  assign n84824 = ~n84024 & ~n84823;
  assign n84825 = n84034 & ~n84810;
  assign n84826 = ~n84824 & ~n84825;
  assign n84827 = ~n84177 & n84826;
  assign n84828 = n83999 & ~n84827;
  assign n84829 = ~n84820 & ~n84828;
  assign n84830 = ~n84024 & n84195;
  assign n84831 = ~n84818 & ~n84830;
  assign n84832 = n84030 & ~n84831;
  assign n84833 = n84829 & ~n84832;
  assign n84834 = pi2672 & ~n84833;
  assign n84835 = ~pi2672 & ~n84832;
  assign n84836 = ~n84828 & n84835;
  assign n84837 = ~n84820 & n84836;
  assign po2817 = n84834 | n84837;
  assign n84839 = ~n83771 & ~n83777;
  assign n84840 = ~n83744 & ~n84839;
  assign n84841 = ~n83833 & ~n84840;
  assign n84842 = n83750 & n83756;
  assign n84843 = n83744 & n84842;
  assign n84844 = n83770 & n84843;
  assign n84845 = n83770 & n83802;
  assign n84846 = ~n84842 & ~n84845;
  assign n84847 = ~n83750 & ~n83770;
  assign n84848 = ~n83756 & n84847;
  assign n84849 = n84846 & ~n84848;
  assign n84850 = n83744 & ~n84849;
  assign n84851 = ~n83780 & ~n84850;
  assign n84852 = ~n83789 & ~n84851;
  assign n84853 = ~n83744 & n83763;
  assign n84854 = n83770 & n84853;
  assign n84855 = ~n84743 & ~n84854;
  assign n84856 = ~n83789 & ~n84855;
  assign n84857 = ~n84852 & ~n84856;
  assign n84858 = ~n84844 & n84857;
  assign n84859 = ~n83803 & ~n83816;
  assign n84860 = ~n84752 & n84859;
  assign n84861 = ~n83744 & ~n84860;
  assign n84862 = ~n83770 & n83821;
  assign n84863 = ~n83806 & ~n84862;
  assign n84864 = n83744 & ~n84863;
  assign n84865 = ~n84861 & ~n84864;
  assign n84866 = ~n84751 & n84865;
  assign n84867 = ~n83792 & ~n83827;
  assign n84868 = n84866 & n84867;
  assign n84869 = n83789 & ~n84868;
  assign n84870 = n84858 & ~n84869;
  assign n84871 = n84841 & n84870;
  assign n84872 = ~pi2693 & ~n84871;
  assign n84873 = pi2693 & n84858;
  assign n84874 = n84841 & n84873;
  assign n84875 = ~n84869 & n84874;
  assign po2819 = n84872 | n84875;
  assign n84877 = ~n83827 & ~n84762;
  assign n84878 = n83744 & ~n84877;
  assign n84879 = ~n83774 & ~n83777;
  assign n84880 = ~n83770 & n84752;
  assign n84881 = ~n84734 & ~n84880;
  assign n84882 = n84879 & n84881;
  assign n84883 = ~n83744 & ~n84882;
  assign n84884 = ~n83789 & n83811;
  assign n84885 = ~n83744 & n84884;
  assign n84886 = n83756 & n84847;
  assign n84887 = ~n84754 & ~n84886;
  assign n84888 = ~n83779 & n84887;
  assign n84889 = n83744 & ~n84888;
  assign n84890 = n83750 & n83802;
  assign n84891 = ~n83770 & n84890;
  assign n84892 = ~n84889 & ~n84891;
  assign n84893 = ~n83789 & ~n84892;
  assign n84894 = ~n84885 & ~n84893;
  assign n84895 = n83750 & ~n83756;
  assign n84896 = ~n83744 & n84895;
  assign n84897 = n83770 & n84896;
  assign n84898 = ~n83770 & n84754;
  assign n84899 = ~n83777 & ~n84898;
  assign n84900 = ~n84759 & n84899;
  assign n84901 = ~n84897 & n84900;
  assign n84902 = n83744 & n83773;
  assign n84903 = n84901 & ~n84902;
  assign n84904 = n83789 & ~n84903;
  assign n84905 = n84894 & ~n84904;
  assign n84906 = ~n84883 & n84905;
  assign n84907 = ~n84878 & n84906;
  assign n84908 = pi2698 & n84907;
  assign n84909 = ~pi2698 & ~n84907;
  assign po2820 = n84908 | n84909;
  assign n84911 = ~n84419 & n84441;
  assign n84912 = ~n84440 & ~n84911;
  assign n84913 = ~n84400 & ~n84912;
  assign n84914 = n84400 & ~n84642;
  assign n84915 = ~n84631 & ~n84914;
  assign n84916 = ~n84913 & n84915;
  assign n84917 = n84437 & ~n84916;
  assign n84918 = ~n84400 & n84455;
  assign n84919 = ~n84917 & ~n84918;
  assign n84920 = ~n84693 & ~n84714;
  assign n84921 = n84400 & ~n84920;
  assign n84922 = n84400 & n84442;
  assign n84923 = n84419 & n84458;
  assign n84924 = n84425 & n84607;
  assign n84925 = ~n84618 & ~n84924;
  assign n84926 = ~n84406 & ~n84925;
  assign n84927 = ~n84699 & ~n84926;
  assign n84928 = ~n84427 & n84927;
  assign n84929 = ~n84923 & n84928;
  assign n84930 = ~n84922 & n84929;
  assign n84931 = ~n84437 & ~n84930;
  assign n84932 = ~n84921 & ~n84931;
  assign n84933 = n84919 & n84932;
  assign n84934 = pi2687 & ~n84933;
  assign n84935 = ~pi2687 & n84933;
  assign po2821 = n84934 | n84935;
  assign n84937 = pi6079 & pi9040;
  assign n84938 = pi6265 & ~pi9040;
  assign n84939 = ~n84937 & ~n84938;
  assign n84940 = ~pi2717 & ~n84939;
  assign n84941 = pi2717 & n84939;
  assign n84942 = ~n84940 & ~n84941;
  assign n84943 = pi6121 & ~pi9040;
  assign n84944 = pi6086 & pi9040;
  assign n84945 = ~n84943 & ~n84944;
  assign n84946 = ~pi2711 & n84945;
  assign n84947 = pi2711 & ~n84945;
  assign n84948 = ~n84946 & ~n84947;
  assign n84949 = pi6275 & ~pi9040;
  assign n84950 = pi5952 & pi9040;
  assign n84951 = ~n84949 & ~n84950;
  assign n84952 = ~pi2710 & ~n84951;
  assign n84953 = pi2710 & n84951;
  assign n84954 = ~n84952 & ~n84953;
  assign n84955 = pi6029 & ~pi9040;
  assign n84956 = pi6266 & pi9040;
  assign n84957 = ~n84955 & ~n84956;
  assign n84958 = ~pi2683 & ~n84957;
  assign n84959 = pi2683 & n84957;
  assign n84960 = ~n84958 & ~n84959;
  assign n84961 = pi6072 & pi9040;
  assign n84962 = pi6046 & ~pi9040;
  assign n84963 = ~n84961 & ~n84962;
  assign n84964 = ~pi2695 & n84963;
  assign n84965 = pi2695 & ~n84963;
  assign n84966 = ~n84964 & ~n84965;
  assign n84967 = n84960 & n84966;
  assign n84968 = n84954 & n84967;
  assign n84969 = ~n84948 & n84968;
  assign n84970 = ~n84960 & n84966;
  assign n84971 = n84954 & n84970;
  assign n84972 = n84948 & n84971;
  assign n84973 = ~n84969 & ~n84972;
  assign n84974 = ~n84960 & ~n84966;
  assign n84975 = n84954 & n84974;
  assign n84976 = ~n84948 & n84975;
  assign n84977 = pi6068 & ~pi9040;
  assign n84978 = pi6074 & pi9040;
  assign n84979 = ~n84977 & ~n84978;
  assign n84980 = ~pi2714 & ~n84979;
  assign n84981 = pi2714 & n84979;
  assign n84982 = ~n84980 & ~n84981;
  assign n84983 = n84960 & ~n84966;
  assign n84984 = ~n84948 & n84983;
  assign n84985 = ~n84954 & n84974;
  assign n84986 = n84948 & n84985;
  assign n84987 = ~n84984 & ~n84986;
  assign n84988 = ~n84982 & ~n84987;
  assign n84989 = ~n84976 & ~n84988;
  assign n84990 = ~n84954 & n84970;
  assign n84991 = n84982 & n84990;
  assign n84992 = n84974 & n84982;
  assign n84993 = ~n84948 & n84992;
  assign n84994 = ~n84991 & ~n84993;
  assign n84995 = n84989 & n84994;
  assign n84996 = n84973 & n84995;
  assign n84997 = n84942 & ~n84996;
  assign n84998 = ~n84942 & ~n84982;
  assign n84999 = ~n84948 & ~n84954;
  assign n85000 = ~n84960 & n84999;
  assign n85001 = ~n84954 & n84966;
  assign n85002 = ~n85000 & ~n85001;
  assign n85003 = n84998 & ~n85002;
  assign n85004 = n84948 & n84954;
  assign n85005 = ~n84966 & n85004;
  assign n85006 = ~n84960 & n85005;
  assign n85007 = n84948 & n84960;
  assign n85008 = ~n84954 & n85007;
  assign n85009 = ~n85006 & ~n85008;
  assign n85010 = ~n84948 & n84982;
  assign n85011 = n84954 & n85010;
  assign n85012 = ~n84974 & n85011;
  assign n85013 = n84968 & n84982;
  assign n85014 = ~n85012 & ~n85013;
  assign n85015 = n85009 & n85014;
  assign n85016 = ~n84942 & ~n85015;
  assign n85017 = ~n84954 & n84967;
  assign n85018 = ~n84982 & n85017;
  assign n85019 = n84948 & n85018;
  assign n85020 = n84954 & n84983;
  assign n85021 = n84948 & n85020;
  assign n85022 = ~n84972 & ~n85021;
  assign n85023 = ~n84982 & ~n85022;
  assign n85024 = ~n85019 & ~n85023;
  assign n85025 = n84982 & n85006;
  assign n85026 = n85024 & ~n85025;
  assign n85027 = ~n85016 & n85026;
  assign n85028 = ~n85003 & n85027;
  assign n85029 = ~n84997 & n85028;
  assign n85030 = ~n84954 & n84983;
  assign n85031 = n84948 & n84982;
  assign n85032 = n85030 & n85031;
  assign n85033 = n85029 & ~n85032;
  assign n85034 = ~pi2729 & ~n85033;
  assign n85035 = pi2729 & ~n85032;
  assign n85036 = n85028 & n85035;
  assign n85037 = ~n84997 & n85036;
  assign po2840 = n85034 | n85037;
  assign n85039 = n84948 & n84990;
  assign n85040 = n84966 & n84999;
  assign n85041 = n84960 & n85040;
  assign n85042 = ~n85039 & ~n85041;
  assign n85043 = n84982 & ~n85042;
  assign n85044 = ~n85006 & ~n85013;
  assign n85045 = ~n84960 & n85004;
  assign n85046 = ~n85008 & ~n85045;
  assign n85047 = ~n84982 & ~n85046;
  assign n85048 = ~n84948 & ~n84982;
  assign n85049 = n84970 & n85048;
  assign n85050 = ~n84954 & n85049;
  assign n85051 = ~n84948 & n85020;
  assign n85052 = ~n84954 & n84982;
  assign n85053 = ~n84966 & n85052;
  assign n85054 = ~n84960 & n85053;
  assign n85055 = ~n85051 & ~n85054;
  assign n85056 = ~n85050 & n85055;
  assign n85057 = ~n85047 & n85056;
  assign n85058 = n85044 & n85057;
  assign n85059 = n84942 & ~n85058;
  assign n85060 = ~n84982 & n85006;
  assign n85061 = n84948 & n85013;
  assign n85062 = ~n85060 & ~n85061;
  assign n85063 = ~n85059 & n85062;
  assign n85064 = ~n85043 & n85063;
  assign n85065 = n84954 & ~n84960;
  assign n85066 = n85010 & n85065;
  assign n85067 = ~n84991 & ~n85066;
  assign n85068 = n84982 & n85020;
  assign n85069 = n84948 & n85030;
  assign n85070 = ~n85068 & ~n85069;
  assign n85071 = ~n84948 & n84971;
  assign n85072 = ~n85039 & ~n85071;
  assign n85073 = ~n84948 & n84967;
  assign n85074 = ~n84954 & ~n84966;
  assign n85075 = ~n85073 & ~n85074;
  assign n85076 = ~n84982 & ~n85075;
  assign n85077 = n85072 & ~n85076;
  assign n85078 = n85070 & n85077;
  assign n85079 = n85067 & n85078;
  assign n85080 = ~n84942 & ~n85079;
  assign n85081 = n85064 & ~n85080;
  assign n85082 = ~pi2731 & ~n85081;
  assign n85083 = pi2731 & ~n85080;
  assign n85084 = n85064 & n85083;
  assign po2843 = n85082 | n85084;
  assign n85086 = ~n85061 & ~n85066;
  assign n85087 = n84948 & n84992;
  assign n85088 = n84960 & n84999;
  assign n85089 = ~n85017 & ~n85088;
  assign n85090 = n84982 & ~n85089;
  assign n85091 = ~n85087 & ~n85090;
  assign n85092 = ~n84982 & n84983;
  assign n85093 = n84948 & n85092;
  assign n85094 = ~n84982 & n84990;
  assign n85095 = ~n85093 & ~n85094;
  assign n85096 = n85091 & n85095;
  assign n85097 = n84960 & n85004;
  assign n85098 = ~n85039 & ~n85097;
  assign n85099 = ~n85071 & n85098;
  assign n85100 = n85096 & n85099;
  assign n85101 = ~n84942 & ~n85100;
  assign n85102 = ~n85006 & ~n85017;
  assign n85103 = ~n85073 & n85102;
  assign n85104 = ~n84982 & ~n85103;
  assign n85105 = ~n84948 & n84985;
  assign n85106 = ~n85051 & ~n85105;
  assign n85107 = ~n85032 & n85106;
  assign n85108 = n84971 & n84982;
  assign n85109 = n85107 & ~n85108;
  assign n85110 = ~n85104 & n85109;
  assign n85111 = n84942 & ~n85110;
  assign n85112 = ~n85039 & n85106;
  assign n85113 = ~n84982 & ~n85112;
  assign n85114 = ~n85111 & ~n85113;
  assign n85115 = ~n85101 & n85114;
  assign n85116 = n85086 & n85115;
  assign n85117 = pi2747 & ~n85116;
  assign n85118 = ~pi2747 & n85116;
  assign po2846 = n85117 | n85118;
  assign n85120 = pi6039 & pi9040;
  assign n85121 = pi6204 & ~pi9040;
  assign n85122 = ~n85120 & ~n85121;
  assign n85123 = ~pi2716 & ~n85122;
  assign n85124 = pi2716 & n85122;
  assign n85125 = ~n85123 & ~n85124;
  assign n85126 = pi6017 & ~pi9040;
  assign n85127 = pi5964 & pi9040;
  assign n85128 = ~n85126 & ~n85127;
  assign n85129 = pi2702 & n85128;
  assign n85130 = ~pi2702 & ~n85128;
  assign n85131 = ~n85129 & ~n85130;
  assign n85132 = pi5963 & ~pi9040;
  assign n85133 = pi6094 & pi9040;
  assign n85134 = ~n85132 & ~n85133;
  assign n85135 = pi2668 & n85134;
  assign n85136 = ~pi2668 & ~n85134;
  assign n85137 = ~n85135 & ~n85136;
  assign n85138 = pi6166 & ~pi9040;
  assign n85139 = pi6043 & pi9040;
  assign n85140 = ~n85138 & ~n85139;
  assign n85141 = ~pi2709 & ~n85140;
  assign n85142 = pi2709 & n85140;
  assign n85143 = ~n85141 & ~n85142;
  assign n85144 = pi6025 & pi9040;
  assign n85145 = pi6167 & ~pi9040;
  assign n85146 = ~n85144 & ~n85145;
  assign n85147 = ~pi2692 & n85146;
  assign n85148 = pi2692 & ~n85146;
  assign n85149 = ~n85147 & ~n85148;
  assign n85150 = n85143 & n85149;
  assign n85151 = n85137 & n85150;
  assign n85152 = pi6089 & ~pi9040;
  assign n85153 = pi6165 & pi9040;
  assign n85154 = ~n85152 & ~n85153;
  assign n85155 = ~pi2700 & ~n85154;
  assign n85156 = pi2700 & n85154;
  assign n85157 = ~n85155 & ~n85156;
  assign n85158 = ~n85149 & n85157;
  assign n85159 = n85143 & n85158;
  assign n85160 = ~n85151 & ~n85159;
  assign n85161 = ~n85149 & ~n85157;
  assign n85162 = ~n85143 & n85161;
  assign n85163 = ~n85137 & n85162;
  assign n85164 = n85160 & ~n85163;
  assign n85165 = n85131 & ~n85164;
  assign n85166 = ~n85143 & ~n85149;
  assign n85167 = n85157 & n85166;
  assign n85168 = ~n85137 & n85167;
  assign n85169 = n85149 & n85157;
  assign n85170 = n85143 & n85169;
  assign n85171 = ~n85137 & n85170;
  assign n85172 = ~n85143 & n85149;
  assign n85173 = ~n85161 & ~n85172;
  assign n85174 = n85137 & ~n85173;
  assign n85175 = ~n85171 & ~n85174;
  assign n85176 = ~n85168 & n85175;
  assign n85177 = ~n85131 & ~n85176;
  assign n85178 = ~n85165 & ~n85177;
  assign n85179 = n85125 & ~n85178;
  assign n85180 = n85131 & ~n85137;
  assign n85181 = n85149 & n85180;
  assign n85182 = ~n85131 & ~n85137;
  assign n85183 = n85161 & n85182;
  assign n85184 = ~n85137 & n85143;
  assign n85185 = ~n85149 & n85184;
  assign n85186 = ~n85151 & ~n85185;
  assign n85187 = ~n85131 & ~n85186;
  assign n85188 = ~n85183 & ~n85187;
  assign n85189 = n85143 & n85161;
  assign n85190 = ~n85137 & n85189;
  assign n85191 = n85137 & n85167;
  assign n85192 = ~n85190 & ~n85191;
  assign n85193 = n85131 & n85137;
  assign n85194 = n85166 & n85193;
  assign n85195 = ~n85143 & n85169;
  assign n85196 = n85131 & n85195;
  assign n85197 = ~n85194 & ~n85196;
  assign n85198 = n85192 & n85197;
  assign n85199 = n85188 & n85198;
  assign n85200 = ~n85181 & n85199;
  assign n85201 = ~n85125 & ~n85200;
  assign n85202 = n85149 & ~n85157;
  assign n85203 = ~n85143 & n85202;
  assign n85204 = ~n85131 & n85203;
  assign n85205 = ~n85137 & n85204;
  assign n85206 = ~n85131 & n85190;
  assign n85207 = ~n85205 & ~n85206;
  assign n85208 = ~n85137 & ~n85143;
  assign n85209 = n85157 & n85208;
  assign n85210 = n85149 & n85209;
  assign n85211 = n85131 & n85210;
  assign n85212 = n85207 & ~n85211;
  assign n85213 = n85150 & ~n85157;
  assign n85214 = ~n85137 & n85213;
  assign n85215 = n85137 & n85158;
  assign n85216 = ~n85214 & ~n85215;
  assign n85217 = n85131 & ~n85216;
  assign n85218 = n85212 & ~n85217;
  assign n85219 = ~n85201 & n85218;
  assign n85220 = ~n85179 & n85219;
  assign n85221 = ~pi2726 & ~n85220;
  assign n85222 = pi2726 & n85220;
  assign po2847 = n85221 | n85222;
  assign n85224 = pi6093 & ~pi9040;
  assign n85225 = pi6145 & pi9040;
  assign n85226 = ~n85224 & ~n85225;
  assign n85227 = pi2690 & n85226;
  assign n85228 = ~pi2690 & ~n85226;
  assign n85229 = ~n85227 & ~n85228;
  assign n85230 = pi6073 & pi9040;
  assign n85231 = pi6179 & ~pi9040;
  assign n85232 = ~n85230 & ~n85231;
  assign n85233 = ~pi2701 & n85232;
  assign n85234 = pi2701 & ~n85232;
  assign n85235 = ~n85233 & ~n85234;
  assign n85236 = pi6040 & ~pi9040;
  assign n85237 = pi6017 & pi9040;
  assign n85238 = ~n85236 & ~n85237;
  assign n85239 = ~pi2694 & n85238;
  assign n85240 = pi2694 & ~n85238;
  assign n85241 = ~n85239 & ~n85240;
  assign n85242 = pi6010 & pi9040;
  assign n85243 = pi6039 & ~pi9040;
  assign n85244 = ~n85242 & ~n85243;
  assign n85245 = ~pi2708 & n85244;
  assign n85246 = pi2708 & ~n85244;
  assign n85247 = ~n85245 & ~n85246;
  assign n85248 = ~n85241 & ~n85247;
  assign n85249 = n85235 & n85248;
  assign n85250 = pi6007 & pi9040;
  assign n85251 = pi6094 & ~pi9040;
  assign n85252 = ~n85250 & ~n85251;
  assign n85253 = pi2718 & n85252;
  assign n85254 = ~pi2718 & ~n85252;
  assign n85255 = ~n85253 & ~n85254;
  assign n85256 = n85249 & ~n85255;
  assign n85257 = n85241 & n85247;
  assign n85258 = n85235 & n85257;
  assign n85259 = ~n85255 & n85258;
  assign n85260 = ~n85256 & ~n85259;
  assign n85261 = ~n85235 & n85257;
  assign n85262 = n85255 & n85261;
  assign n85263 = n85241 & ~n85247;
  assign n85264 = n85235 & n85263;
  assign n85265 = n85255 & n85264;
  assign n85266 = ~n85262 & ~n85265;
  assign n85267 = n85260 & n85266;
  assign n85268 = n85229 & ~n85267;
  assign n85269 = ~n85241 & n85247;
  assign n85270 = n85235 & n85269;
  assign n85271 = n85255 & n85270;
  assign n85272 = ~n85264 & ~n85271;
  assign n85273 = n85229 & ~n85272;
  assign n85274 = ~n85229 & ~n85241;
  assign n85275 = ~n85255 & n85274;
  assign n85276 = ~n85235 & ~n85247;
  assign n85277 = n85255 & n85257;
  assign n85278 = ~n85276 & ~n85277;
  assign n85279 = ~n85229 & ~n85278;
  assign n85280 = ~n85275 & ~n85279;
  assign n85281 = ~n85235 & n85269;
  assign n85282 = ~n85255 & n85281;
  assign n85283 = n85280 & ~n85282;
  assign n85284 = ~n85241 & n85255;
  assign n85285 = ~n85235 & n85284;
  assign n85286 = ~n85247 & n85285;
  assign n85287 = n85283 & ~n85286;
  assign n85288 = ~n85273 & n85287;
  assign n85289 = pi6048 & pi9040;
  assign n85290 = pi6025 & ~pi9040;
  assign n85291 = ~n85289 & ~n85290;
  assign n85292 = ~pi2699 & ~n85291;
  assign n85293 = pi2699 & n85291;
  assign n85294 = ~n85292 & ~n85293;
  assign n85295 = ~n85288 & ~n85294;
  assign n85296 = n85235 & ~n85241;
  assign n85297 = ~n85229 & n85255;
  assign n85298 = n85294 & n85297;
  assign n85299 = n85296 & n85298;
  assign n85300 = n85235 & ~n85255;
  assign n85301 = n85241 & n85300;
  assign n85302 = ~n85229 & ~n85301;
  assign n85303 = ~n85235 & n85255;
  assign n85304 = n85247 & n85303;
  assign n85305 = ~n85248 & ~n85296;
  assign n85306 = ~n85255 & ~n85305;
  assign n85307 = ~n85261 & ~n85306;
  assign n85308 = n85229 & n85307;
  assign n85309 = ~n85304 & n85308;
  assign n85310 = ~n85302 & ~n85309;
  assign n85311 = n85241 & n85303;
  assign n85312 = ~n85247 & n85311;
  assign n85313 = ~n85310 & ~n85312;
  assign n85314 = n85294 & ~n85313;
  assign n85315 = ~n85299 & ~n85314;
  assign n85316 = ~n85295 & n85315;
  assign n85317 = ~n85268 & n85316;
  assign n85318 = ~n85229 & n85282;
  assign n85319 = n85317 & ~n85318;
  assign n85320 = pi2721 & ~n85319;
  assign n85321 = ~pi2721 & ~n85318;
  assign n85322 = n85316 & n85321;
  assign n85323 = ~n85268 & n85322;
  assign po2854 = n85320 | n85323;
  assign n85325 = pi5965 & ~pi9040;
  assign n85326 = pi6032 & pi9040;
  assign n85327 = ~n85325 & ~n85326;
  assign n85328 = pi2719 & n85327;
  assign n85329 = ~pi2719 & ~n85327;
  assign n85330 = ~n85328 & ~n85329;
  assign n85331 = pi6183 & ~pi9040;
  assign n85332 = pi6029 & pi9040;
  assign n85333 = ~n85331 & ~n85332;
  assign n85334 = ~pi2708 & ~n85333;
  assign n85335 = pi2708 & n85333;
  assign n85336 = ~n85334 & ~n85335;
  assign n85337 = pi5956 & ~pi9040;
  assign n85338 = pi6265 & pi9040;
  assign n85339 = ~n85337 & ~n85338;
  assign n85340 = ~pi2699 & n85339;
  assign n85341 = pi2699 & ~n85339;
  assign n85342 = ~n85340 & ~n85341;
  assign n85343 = n85336 & n85342;
  assign n85344 = pi6139 & ~pi9040;
  assign n85345 = pi6044 & pi9040;
  assign n85346 = ~n85344 & ~n85345;
  assign n85347 = ~pi2674 & n85346;
  assign n85348 = pi2674 & ~n85346;
  assign n85349 = ~n85347 & ~n85348;
  assign n85350 = ~n85342 & ~n85349;
  assign n85351 = pi6142 & pi9040;
  assign n85352 = pi6241 & ~pi9040;
  assign n85353 = ~n85351 & ~n85352;
  assign n85354 = pi2707 & n85353;
  assign n85355 = ~pi2707 & ~n85353;
  assign n85356 = ~n85354 & ~n85355;
  assign n85357 = ~n85336 & ~n85356;
  assign n85358 = n85350 & n85357;
  assign n85359 = ~n85343 & ~n85358;
  assign n85360 = n85342 & n85356;
  assign n85361 = n85359 & ~n85360;
  assign n85362 = n85330 & ~n85361;
  assign n85363 = ~n85330 & n85356;
  assign n85364 = ~n85342 & n85363;
  assign n85365 = n85336 & n85356;
  assign n85366 = ~n85349 & n85365;
  assign n85367 = ~n85342 & n85349;
  assign n85368 = n85336 & n85367;
  assign n85369 = ~n85356 & n85368;
  assign n85370 = ~n85366 & ~n85369;
  assign n85371 = ~n85336 & n85342;
  assign n85372 = ~n85330 & ~n85356;
  assign n85373 = n85371 & n85372;
  assign n85374 = n85370 & ~n85373;
  assign n85375 = ~n85364 & n85374;
  assign n85376 = ~n85362 & n85375;
  assign n85377 = pi6047 & pi9040;
  assign n85378 = pi6072 & ~pi9040;
  assign n85379 = ~n85377 & ~n85378;
  assign n85380 = ~pi2713 & ~n85379;
  assign n85381 = pi2713 & n85379;
  assign n85382 = ~n85380 & ~n85381;
  assign n85383 = ~n85376 & n85382;
  assign n85384 = n85342 & ~n85349;
  assign n85385 = n85336 & n85384;
  assign n85386 = ~n85356 & n85385;
  assign n85387 = n85342 & n85349;
  assign n85388 = n85336 & n85387;
  assign n85389 = n85356 & n85388;
  assign n85390 = ~n85386 & ~n85389;
  assign n85391 = n85330 & ~n85390;
  assign n85392 = ~n85383 & ~n85391;
  assign n85393 = n85356 & n85368;
  assign n85394 = n85336 & ~n85342;
  assign n85395 = ~n85349 & n85394;
  assign n85396 = ~n85336 & n85349;
  assign n85397 = ~n85342 & n85396;
  assign n85398 = ~n85395 & ~n85397;
  assign n85399 = n85330 & ~n85398;
  assign n85400 = ~n85393 & ~n85399;
  assign n85401 = ~n85336 & n85384;
  assign n85402 = n85356 & n85401;
  assign n85403 = n85400 & ~n85402;
  assign n85404 = ~n85382 & ~n85403;
  assign n85405 = ~n85350 & ~n85387;
  assign n85406 = ~n85336 & ~n85405;
  assign n85407 = ~n85356 & n85387;
  assign n85408 = ~n85406 & ~n85407;
  assign n85409 = ~n85330 & ~n85408;
  assign n85410 = ~n85382 & n85409;
  assign n85411 = ~n85404 & ~n85410;
  assign n85412 = n85392 & n85411;
  assign n85413 = pi2735 & ~n85412;
  assign n85414 = ~pi2735 & n85392;
  assign n85415 = n85411 & n85414;
  assign po2855 = n85413 | n85415;
  assign n85417 = ~n84969 & ~n85000;
  assign n85418 = n84942 & ~n85417;
  assign n85419 = ~n85005 & ~n85045;
  assign n85420 = ~n84975 & n85419;
  assign n85421 = ~n84982 & ~n85420;
  assign n85422 = n84942 & n85421;
  assign n85423 = ~n85418 & ~n85422;
  assign n85424 = n84968 & n85048;
  assign n85425 = ~n85050 & ~n85424;
  assign n85426 = ~n85008 & ~n85074;
  assign n85427 = n84982 & ~n85426;
  assign n85428 = n84942 & n85427;
  assign n85429 = n85425 & ~n85428;
  assign n85430 = n84966 & n85004;
  assign n85431 = n84960 & n85430;
  assign n85432 = n84948 & n84970;
  assign n85433 = ~n85041 & ~n85432;
  assign n85434 = n84982 & ~n85433;
  assign n85435 = ~n85006 & ~n85051;
  assign n85436 = n84948 & n84967;
  assign n85437 = ~n85030 & ~n85436;
  assign n85438 = ~n84982 & ~n85437;
  assign n85439 = n85435 & ~n85438;
  assign n85440 = ~n85434 & n85439;
  assign n85441 = ~n85431 & n85440;
  assign n85442 = ~n84942 & ~n85441;
  assign n85443 = ~n85071 & n85106;
  assign n85444 = n84982 & ~n85443;
  assign n85445 = ~n85442 & ~n85444;
  assign n85446 = n85429 & n85445;
  assign n85447 = n85423 & n85446;
  assign n85448 = ~pi2750 & ~n85447;
  assign n85449 = pi2750 & n85429;
  assign n85450 = n85423 & n85449;
  assign n85451 = n85445 & n85450;
  assign po2856 = n85448 | n85451;
  assign n85453 = pi6040 & pi9040;
  assign n85454 = pi6165 & ~pi9040;
  assign n85455 = ~n85453 & ~n85454;
  assign n85456 = ~pi2692 & ~n85455;
  assign n85457 = pi2692 & n85455;
  assign n85458 = ~n85456 & ~n85457;
  assign n85459 = pi6010 & ~pi9040;
  assign n85460 = pi6167 & pi9040;
  assign n85461 = ~n85459 & ~n85460;
  assign n85462 = pi2715 & n85461;
  assign n85463 = ~pi2715 & ~n85461;
  assign n85464 = ~n85462 & ~n85463;
  assign n85465 = pi6030 & ~pi9040;
  assign n85466 = pi6093 & pi9040;
  assign n85467 = ~n85465 & ~n85466;
  assign n85468 = pi2697 & n85467;
  assign n85469 = ~pi2697 & ~n85467;
  assign n85470 = ~n85468 & ~n85469;
  assign n85471 = ~n85464 & ~n85470;
  assign n85472 = pi6073 & ~pi9040;
  assign n85473 = pi6166 & pi9040;
  assign n85474 = ~n85472 & ~n85473;
  assign n85475 = ~pi2717 & n85474;
  assign n85476 = pi2717 & ~n85474;
  assign n85477 = ~n85475 & ~n85476;
  assign n85478 = n85471 & ~n85477;
  assign n85479 = pi5963 & pi9040;
  assign n85480 = pi6124 & ~pi9040;
  assign n85481 = ~n85479 & ~n85480;
  assign n85482 = pi2695 & n85481;
  assign n85483 = ~pi2695 & ~n85481;
  assign n85484 = ~n85482 & ~n85483;
  assign n85485 = pi6075 & ~pi9040;
  assign n85486 = pi6034 & pi9040;
  assign n85487 = ~n85485 & ~n85486;
  assign n85488 = pi2709 & n85487;
  assign n85489 = ~pi2709 & ~n85487;
  assign n85490 = ~n85488 & ~n85489;
  assign n85491 = n85477 & ~n85490;
  assign n85492 = n85484 & n85491;
  assign n85493 = n85464 & n85492;
  assign n85494 = n85477 & n85490;
  assign n85495 = ~n85484 & n85494;
  assign n85496 = n85464 & n85495;
  assign n85497 = ~n85493 & ~n85496;
  assign n85498 = ~n85477 & n85490;
  assign n85499 = ~n85484 & n85498;
  assign n85500 = ~n85464 & ~n85484;
  assign n85501 = ~n85490 & n85500;
  assign n85502 = n85477 & n85501;
  assign n85503 = ~n85499 & ~n85502;
  assign n85504 = n85470 & ~n85503;
  assign n85505 = n85497 & ~n85504;
  assign n85506 = ~n85478 & n85505;
  assign n85507 = n85458 & ~n85506;
  assign n85508 = ~n85477 & ~n85490;
  assign n85509 = ~n85484 & n85508;
  assign n85510 = n85464 & n85509;
  assign n85511 = ~n85470 & n85510;
  assign n85512 = ~n85464 & n85470;
  assign n85513 = n85509 & n85512;
  assign n85514 = ~n85464 & n85484;
  assign n85515 = n85477 & n85514;
  assign n85516 = ~n85513 & ~n85515;
  assign n85517 = n85484 & n85494;
  assign n85518 = ~n85499 & ~n85517;
  assign n85519 = ~n85464 & n85494;
  assign n85520 = n85518 & ~n85519;
  assign n85521 = ~n85470 & ~n85520;
  assign n85522 = n85484 & ~n85490;
  assign n85523 = ~n85477 & n85522;
  assign n85524 = n85464 & n85523;
  assign n85525 = ~n85484 & n85491;
  assign n85526 = n85464 & n85525;
  assign n85527 = ~n85524 & ~n85526;
  assign n85528 = n85484 & n85498;
  assign n85529 = n85470 & n85528;
  assign n85530 = n85527 & ~n85529;
  assign n85531 = ~n85521 & n85530;
  assign n85532 = n85516 & n85531;
  assign n85533 = ~n85458 & ~n85532;
  assign n85534 = ~n85511 & ~n85533;
  assign n85535 = ~n85507 & n85534;
  assign n85536 = n85512 & n85517;
  assign n85537 = n85470 & n85522;
  assign n85538 = n85464 & n85537;
  assign n85539 = ~n85536 & ~n85538;
  assign n85540 = n85470 & n85496;
  assign n85541 = n85539 & ~n85540;
  assign n85542 = n85535 & n85541;
  assign n85543 = ~pi2725 & ~n85542;
  assign n85544 = pi2725 & n85541;
  assign n85545 = n85534 & n85544;
  assign n85546 = ~n85507 & n85545;
  assign po2858 = n85543 | n85546;
  assign n85548 = ~n85125 & ~n85131;
  assign n85549 = ~n85137 & n85150;
  assign n85550 = n85137 & n85143;
  assign n85551 = n85161 & n85550;
  assign n85552 = ~n85137 & n85158;
  assign n85553 = ~n85551 & ~n85552;
  assign n85554 = ~n85549 & n85553;
  assign n85555 = n85548 & ~n85554;
  assign n85556 = ~n85157 & n85208;
  assign n85557 = n85137 & n85213;
  assign n85558 = ~n85556 & ~n85557;
  assign n85559 = ~n85159 & ~n85162;
  assign n85560 = n85558 & n85559;
  assign n85561 = n85131 & ~n85560;
  assign n85562 = n85137 & ~n85143;
  assign n85563 = n85157 & n85562;
  assign n85564 = n85149 & n85563;
  assign n85565 = ~n85561 & ~n85564;
  assign n85566 = ~n85125 & ~n85565;
  assign n85567 = ~n85555 & ~n85566;
  assign n85568 = n85143 & n85180;
  assign n85569 = n85157 & n85568;
  assign n85570 = ~n85163 & ~n85569;
  assign n85571 = ~n85158 & ~n85202;
  assign n85572 = n85137 & ~n85571;
  assign n85573 = ~n85203 & ~n85572;
  assign n85574 = ~n85131 & ~n85573;
  assign n85575 = ~n85170 & ~n85549;
  assign n85576 = ~n85551 & n85575;
  assign n85577 = n85131 & ~n85576;
  assign n85578 = ~n85574 & ~n85577;
  assign n85579 = n85137 & n85203;
  assign n85580 = ~n85191 & ~n85579;
  assign n85581 = ~n85210 & n85580;
  assign n85582 = ~n85183 & n85581;
  assign n85583 = n85578 & n85582;
  assign n85584 = n85125 & ~n85583;
  assign n85585 = n85570 & ~n85584;
  assign n85586 = n85567 & n85585;
  assign n85587 = pi2720 & ~n85586;
  assign n85588 = ~pi2720 & n85586;
  assign po2859 = n85587 | n85588;
  assign n85590 = n85330 & n85356;
  assign n85591 = n85384 & n85590;
  assign n85592 = n85336 & n85591;
  assign n85593 = n85330 & ~n85356;
  assign n85594 = n85350 & n85593;
  assign n85595 = n85336 & ~n85356;
  assign n85596 = n85349 & n85595;
  assign n85597 = n85342 & n85596;
  assign n85598 = n85330 & n85368;
  assign n85599 = n85356 & n85598;
  assign n85600 = ~n85597 & ~n85599;
  assign n85601 = ~n85594 & n85600;
  assign n85602 = ~n85592 & n85601;
  assign n85603 = ~n85358 & n85602;
  assign n85604 = ~n85382 & ~n85603;
  assign n85605 = ~n85330 & n85397;
  assign n85606 = n85356 & n85605;
  assign n85607 = n85342 & n85595;
  assign n85608 = ~n85407 & ~n85607;
  assign n85609 = ~n85330 & ~n85608;
  assign n85610 = ~n85606 & ~n85609;
  assign n85611 = ~n85382 & ~n85610;
  assign n85612 = n85356 & n85395;
  assign n85613 = ~n85596 & ~n85612;
  assign n85614 = ~n85402 & n85613;
  assign n85615 = ~n85330 & ~n85614;
  assign n85616 = ~n85611 & ~n85615;
  assign n85617 = ~n85604 & n85616;
  assign n85618 = ~n85336 & n85356;
  assign n85619 = n85330 & n85618;
  assign n85620 = n85387 & n85619;
  assign n85621 = ~n85336 & n85593;
  assign n85622 = ~n85342 & n85621;
  assign n85623 = ~n85356 & n85397;
  assign n85624 = ~n85330 & n85336;
  assign n85625 = ~n85342 & n85624;
  assign n85626 = ~n85336 & n85360;
  assign n85627 = ~n85625 & ~n85626;
  assign n85628 = ~n85623 & n85627;
  assign n85629 = ~n85401 & n85628;
  assign n85630 = n85330 & n85384;
  assign n85631 = ~n85356 & n85630;
  assign n85632 = n85356 & n85387;
  assign n85633 = ~n85336 & ~n85349;
  assign n85634 = ~n85632 & ~n85633;
  assign n85635 = n85330 & ~n85634;
  assign n85636 = ~n85631 & ~n85635;
  assign n85637 = n85629 & n85636;
  assign n85638 = n85382 & ~n85637;
  assign n85639 = ~n85622 & ~n85638;
  assign n85640 = ~n85620 & n85639;
  assign n85641 = n85617 & n85640;
  assign n85642 = pi2732 & n85641;
  assign n85643 = ~pi2732 & ~n85641;
  assign po2860 = n85642 | n85643;
  assign n85645 = pi6204 & pi9040;
  assign n85646 = pi6170 & ~pi9040;
  assign n85647 = ~n85645 & ~n85646;
  assign n85648 = pi2694 & n85647;
  assign n85649 = ~pi2694 & ~n85647;
  assign n85650 = ~n85648 & ~n85649;
  assign n85651 = pi6088 & pi9040;
  assign n85652 = pi5964 & ~pi9040;
  assign n85653 = ~n85651 & ~n85652;
  assign n85654 = ~pi2716 & ~n85653;
  assign n85655 = pi2716 & n85653;
  assign n85656 = ~n85654 & ~n85655;
  assign n85657 = pi5950 & ~pi9040;
  assign n85658 = pi6124 & pi9040;
  assign n85659 = ~n85657 & ~n85658;
  assign n85660 = ~pi2701 & n85659;
  assign n85661 = pi2701 & ~n85659;
  assign n85662 = ~n85660 & ~n85661;
  assign n85663 = pi6043 & ~pi9040;
  assign n85664 = pi6173 & pi9040;
  assign n85665 = ~n85663 & ~n85664;
  assign n85666 = pi2684 & n85665;
  assign n85667 = ~pi2684 & ~n85665;
  assign n85668 = ~n85666 & ~n85667;
  assign n85669 = pi6048 & ~pi9040;
  assign n85670 = pi6075 & pi9040;
  assign n85671 = ~n85669 & ~n85670;
  assign n85672 = pi2704 & n85671;
  assign n85673 = ~pi2704 & ~n85671;
  assign n85674 = ~n85672 & ~n85673;
  assign n85675 = ~n85668 & ~n85674;
  assign n85676 = ~n85662 & n85675;
  assign n85677 = ~n85656 & n85676;
  assign n85678 = pi6007 & ~pi9040;
  assign n85679 = pi6089 & pi9040;
  assign n85680 = ~n85678 & ~n85679;
  assign n85681 = ~pi2700 & n85680;
  assign n85682 = pi2700 & ~n85680;
  assign n85683 = ~n85681 & ~n85682;
  assign n85684 = n85656 & n85662;
  assign n85685 = ~n85683 & n85684;
  assign n85686 = n85668 & n85683;
  assign n85687 = n85662 & n85686;
  assign n85688 = ~n85656 & n85687;
  assign n85689 = ~n85685 & ~n85688;
  assign n85690 = n85656 & ~n85662;
  assign n85691 = n85668 & n85690;
  assign n85692 = n85689 & ~n85691;
  assign n85693 = ~n85674 & ~n85692;
  assign n85694 = n85656 & n85683;
  assign n85695 = ~n85668 & n85674;
  assign n85696 = n85694 & n85695;
  assign n85697 = n85683 & n85684;
  assign n85698 = ~n85668 & n85697;
  assign n85699 = ~n85696 & ~n85698;
  assign n85700 = ~n85693 & n85699;
  assign n85701 = ~n85677 & n85700;
  assign n85702 = ~n85656 & ~n85662;
  assign n85703 = ~n85683 & n85702;
  assign n85704 = ~n85668 & n85703;
  assign n85705 = ~n85683 & n85690;
  assign n85706 = n85668 & n85705;
  assign n85707 = ~n85704 & ~n85706;
  assign n85708 = n85701 & n85707;
  assign n85709 = ~n85650 & ~n85708;
  assign n85710 = n85683 & n85690;
  assign n85711 = ~n85668 & n85710;
  assign n85712 = ~n85703 & ~n85711;
  assign n85713 = ~n85674 & ~n85712;
  assign n85714 = n85686 & n85702;
  assign n85715 = ~n85668 & n85683;
  assign n85716 = n85662 & n85715;
  assign n85717 = ~n85656 & n85716;
  assign n85718 = ~n85714 & ~n85717;
  assign n85719 = n85656 & n85686;
  assign n85720 = ~n85668 & n85705;
  assign n85721 = ~n85719 & ~n85720;
  assign n85722 = n85674 & ~n85721;
  assign n85723 = n85718 & ~n85722;
  assign n85724 = ~n85713 & n85723;
  assign n85725 = n85650 & ~n85724;
  assign n85726 = n85656 & ~n85683;
  assign n85727 = n85668 & n85726;
  assign n85728 = ~n85656 & ~n85683;
  assign n85729 = ~n85668 & n85728;
  assign n85730 = ~n85727 & ~n85729;
  assign n85731 = ~n85674 & ~n85730;
  assign n85732 = ~n85656 & n85662;
  assign n85733 = ~n85683 & n85732;
  assign n85734 = n85668 & n85733;
  assign n85735 = ~n85714 & ~n85734;
  assign n85736 = ~n85697 & n85735;
  assign n85737 = n85674 & ~n85736;
  assign n85738 = ~n85731 & ~n85737;
  assign n85739 = n85662 & n85683;
  assign n85740 = n85674 & n85739;
  assign n85741 = ~n85668 & n85740;
  assign n85742 = n85738 & ~n85741;
  assign n85743 = ~n85725 & n85742;
  assign n85744 = ~n85709 & n85743;
  assign n85745 = ~pi2728 & ~n85744;
  assign n85746 = pi2728 & n85744;
  assign po2861 = n85745 | n85746;
  assign n85748 = n85131 & n85158;
  assign n85749 = ~n85137 & n85748;
  assign n85750 = ~n85214 & ~n85749;
  assign n85751 = n85157 & n85550;
  assign n85752 = ~n85157 & n85184;
  assign n85753 = ~n85137 & n85149;
  assign n85754 = ~n85752 & ~n85753;
  assign n85755 = ~n85131 & ~n85754;
  assign n85756 = ~n85751 & ~n85755;
  assign n85757 = n85750 & n85756;
  assign n85758 = n85125 & ~n85757;
  assign n85759 = ~n85189 & ~n85191;
  assign n85760 = ~n85137 & n85169;
  assign n85761 = n85759 & ~n85760;
  assign n85762 = n85131 & ~n85761;
  assign n85763 = n85158 & n85182;
  assign n85764 = ~n85163 & ~n85763;
  assign n85765 = ~n85762 & n85764;
  assign n85766 = ~n85213 & ~n85564;
  assign n85767 = ~n85131 & ~n85766;
  assign n85768 = n85765 & ~n85767;
  assign n85769 = ~n85125 & ~n85768;
  assign n85770 = ~n85758 & ~n85769;
  assign n85771 = ~n85137 & n85202;
  assign n85772 = n85137 & ~n85559;
  assign n85773 = ~n85771 & ~n85772;
  assign n85774 = ~n85131 & ~n85773;
  assign n85775 = ~n85170 & ~n85203;
  assign n85776 = ~n85189 & n85775;
  assign n85777 = n85193 & ~n85776;
  assign n85778 = ~n85774 & ~n85777;
  assign n85779 = n85770 & n85778;
  assign n85780 = ~pi2722 & ~n85779;
  assign n85781 = pi2722 & n85778;
  assign n85782 = ~n85769 & n85781;
  assign n85783 = ~n85758 & n85782;
  assign po2862 = n85780 | n85783;
  assign n85785 = pi6068 & pi9040;
  assign n85786 = pi6171 & ~pi9040;
  assign n85787 = ~n85785 & ~n85786;
  assign n85788 = pi2705 & n85787;
  assign n85789 = ~pi2705 & ~n85787;
  assign n85790 = ~n85788 & ~n85789;
  assign n85791 = pi5956 & pi9040;
  assign n85792 = pi6266 & ~pi9040;
  assign n85793 = ~n85791 & ~n85792;
  assign n85794 = pi2712 & n85793;
  assign n85795 = ~pi2712 & ~n85793;
  assign n85796 = ~n85794 & ~n85795;
  assign n85797 = pi5952 & ~pi9040;
  assign n85798 = pi6139 & pi9040;
  assign n85799 = ~n85797 & ~n85798;
  assign n85800 = pi2686 & n85799;
  assign n85801 = ~pi2686 & ~n85799;
  assign n85802 = ~n85800 & ~n85801;
  assign n85803 = n85796 & ~n85802;
  assign n85804 = pi6256 & pi9040;
  assign n85805 = pi6142 & ~pi9040;
  assign n85806 = ~n85804 & ~n85805;
  assign n85807 = pi2703 & n85806;
  assign n85808 = ~pi2703 & ~n85806;
  assign n85809 = ~n85807 & ~n85808;
  assign n85810 = pi6046 & pi9040;
  assign n85811 = pi5991 & ~pi9040;
  assign n85812 = ~n85810 & ~n85811;
  assign n85813 = ~pi2713 & ~n85812;
  assign n85814 = pi2713 & n85812;
  assign n85815 = ~n85813 & ~n85814;
  assign n85816 = ~n85809 & ~n85815;
  assign n85817 = pi6047 & ~pi9040;
  assign n85818 = pi6121 & pi9040;
  assign n85819 = ~n85817 & ~n85818;
  assign n85820 = pi2674 & n85819;
  assign n85821 = ~pi2674 & ~n85819;
  assign n85822 = ~n85820 & ~n85821;
  assign n85823 = n85809 & n85815;
  assign n85824 = ~n85822 & n85823;
  assign n85825 = ~n85816 & ~n85824;
  assign n85826 = n85803 & ~n85825;
  assign n85827 = ~n85802 & ~n85822;
  assign n85828 = n85816 & n85827;
  assign n85829 = ~n85826 & ~n85828;
  assign n85830 = n85790 & ~n85829;
  assign n85831 = ~pi2674 & n85819;
  assign n85832 = pi2674 & ~n85819;
  assign n85833 = ~n85831 & ~n85832;
  assign n85834 = n85823 & ~n85833;
  assign n85835 = ~n85796 & n85834;
  assign n85836 = n85815 & ~n85833;
  assign n85837 = ~n85796 & ~n85833;
  assign n85838 = ~n85836 & ~n85837;
  assign n85839 = n85802 & ~n85838;
  assign n85840 = ~n85796 & ~n85822;
  assign n85841 = ~n85809 & n85840;
  assign n85842 = n85815 & n85841;
  assign n85843 = ~n85839 & ~n85842;
  assign n85844 = ~n85835 & n85843;
  assign n85845 = n85790 & ~n85844;
  assign n85846 = ~n85830 & ~n85845;
  assign n85847 = n85796 & ~n85833;
  assign n85848 = n85809 & n85847;
  assign n85849 = ~n85815 & n85848;
  assign n85850 = n85809 & ~n85815;
  assign n85851 = n85833 & n85850;
  assign n85852 = ~n85796 & n85851;
  assign n85853 = ~n85849 & ~n85852;
  assign n85854 = ~n85802 & ~n85853;
  assign n85855 = ~n85809 & n85815;
  assign n85856 = ~n85836 & ~n85855;
  assign n85857 = n85796 & ~n85856;
  assign n85858 = ~n85851 & ~n85857;
  assign n85859 = ~n85802 & ~n85858;
  assign n85860 = ~n85796 & n85809;
  assign n85861 = ~n85802 & n85833;
  assign n85862 = n85860 & n85861;
  assign n85863 = ~n85809 & n85822;
  assign n85864 = ~n85851 & ~n85863;
  assign n85865 = ~n85796 & ~n85864;
  assign n85866 = n85796 & n85802;
  assign n85867 = n85823 & n85866;
  assign n85868 = ~n85822 & n85867;
  assign n85869 = ~n85865 & ~n85868;
  assign n85870 = ~n85862 & n85869;
  assign n85871 = ~n85859 & n85870;
  assign n85872 = ~n85849 & n85871;
  assign n85873 = ~n85790 & ~n85872;
  assign n85874 = n85816 & n85833;
  assign n85875 = n85796 & n85874;
  assign n85876 = ~n85796 & n85836;
  assign n85877 = ~n85875 & ~n85876;
  assign n85878 = n85802 & ~n85877;
  assign n85879 = ~n85873 & ~n85878;
  assign n85880 = ~n85854 & n85879;
  assign n85881 = n85846 & n85880;
  assign n85882 = pi2745 & n85881;
  assign n85883 = ~pi2745 & ~n85881;
  assign po2863 = n85882 | n85883;
  assign n85885 = ~n85131 & ~n85775;
  assign n85886 = n85137 & n85159;
  assign n85887 = ~n85885 & ~n85886;
  assign n85888 = n85137 & ~n85149;
  assign n85889 = ~n85166 & ~n85888;
  assign n85890 = ~n85213 & n85889;
  assign n85891 = n85131 & ~n85890;
  assign n85892 = n85887 & ~n85891;
  assign n85893 = ~n85125 & ~n85892;
  assign n85894 = ~n85131 & n85168;
  assign n85895 = ~n85206 & ~n85894;
  assign n85896 = ~n85211 & n85895;
  assign n85897 = n85131 & n85185;
  assign n85898 = ~n85196 & ~n85897;
  assign n85899 = n85137 & n85170;
  assign n85900 = ~n85131 & n85166;
  assign n85901 = ~n85899 & ~n85900;
  assign n85902 = ~n85579 & n85901;
  assign n85903 = ~n85210 & n85902;
  assign n85904 = n85898 & n85903;
  assign n85905 = ~n85752 & n85904;
  assign n85906 = n85125 & ~n85905;
  assign n85907 = n85896 & ~n85906;
  assign n85908 = ~n85893 & n85907;
  assign n85909 = ~pi2723 & ~n85908;
  assign n85910 = pi2723 & n85896;
  assign n85911 = ~n85893 & n85910;
  assign n85912 = ~n85906 & n85911;
  assign po2864 = n85909 | n85912;
  assign n85914 = n85356 & n85406;
  assign n85915 = ~n85385 & ~n85396;
  assign n85916 = ~n85330 & ~n85915;
  assign n85917 = ~n85914 & ~n85916;
  assign n85918 = n85349 & n85365;
  assign n85919 = ~n85633 & ~n85918;
  assign n85920 = ~n85388 & n85919;
  assign n85921 = n85330 & ~n85920;
  assign n85922 = n85917 & ~n85921;
  assign n85923 = ~n85356 & n85395;
  assign n85924 = n85922 & ~n85923;
  assign n85925 = ~n85382 & ~n85924;
  assign n85926 = n85593 & ~n85915;
  assign n85927 = ~n85397 & ~n85401;
  assign n85928 = ~n85388 & ~n85395;
  assign n85929 = n85927 & n85928;
  assign n85930 = n85356 & ~n85929;
  assign n85931 = ~n85926 & ~n85930;
  assign n85932 = ~n85369 & n85931;
  assign n85933 = n85382 & ~n85932;
  assign n85934 = ~n85925 & ~n85933;
  assign n85935 = n85356 & n85385;
  assign n85936 = ~n85923 & ~n85935;
  assign n85937 = ~n85330 & ~n85936;
  assign n85938 = n85934 & ~n85937;
  assign n85939 = pi2734 & ~n85938;
  assign n85940 = ~pi2734 & ~n85937;
  assign n85941 = ~n85933 & n85940;
  assign n85942 = ~n85925 & n85941;
  assign po2866 = n85939 | n85942;
  assign n85944 = n85668 & n85697;
  assign n85945 = ~n85717 & ~n85726;
  assign n85946 = n85674 & ~n85945;
  assign n85947 = ~n85944 & ~n85946;
  assign n85948 = ~n85711 & n85947;
  assign n85949 = ~n85674 & n85714;
  assign n85950 = ~n85704 & ~n85949;
  assign n85951 = ~n85734 & n85950;
  assign n85952 = n85948 & n85951;
  assign n85953 = n85650 & ~n85952;
  assign n85954 = n85668 & n85710;
  assign n85955 = ~n85688 & ~n85954;
  assign n85956 = n85683 & n85702;
  assign n85957 = n85674 & n85956;
  assign n85958 = n85668 & n85703;
  assign n85959 = ~n85957 & ~n85958;
  assign n85960 = ~n85662 & ~n85683;
  assign n85961 = n85656 & n85668;
  assign n85962 = ~n85960 & ~n85961;
  assign n85963 = ~n85739 & n85962;
  assign n85964 = ~n85674 & ~n85963;
  assign n85965 = ~n85668 & n85733;
  assign n85966 = ~n85698 & ~n85965;
  assign n85967 = ~n85964 & n85966;
  assign n85968 = n85959 & n85967;
  assign n85969 = n85955 & n85968;
  assign n85970 = ~n85650 & ~n85969;
  assign n85971 = ~n85953 & ~n85970;
  assign n85972 = pi2724 & ~n85971;
  assign n85973 = ~pi2724 & ~n85953;
  assign n85974 = ~n85970 & n85973;
  assign po2867 = n85972 | n85974;
  assign n85976 = ~n85796 & n85816;
  assign n85977 = ~n85833 & n85850;
  assign n85978 = ~n85976 & ~n85977;
  assign n85979 = ~n85790 & n85802;
  assign n85980 = ~n85978 & n85979;
  assign n85981 = n85847 & n85855;
  assign n85982 = ~n85824 & ~n85874;
  assign n85983 = n85796 & ~n85982;
  assign n85984 = ~n85981 & ~n85983;
  assign n85985 = ~n85790 & ~n85984;
  assign n85986 = ~n85980 & ~n85985;
  assign n85987 = ~n85796 & n85802;
  assign n85988 = n85815 & n85987;
  assign n85989 = ~n85822 & n85855;
  assign n85990 = ~n85834 & ~n85989;
  assign n85991 = n85816 & n85822;
  assign n85992 = n85796 & n85991;
  assign n85993 = n85990 & ~n85992;
  assign n85994 = n85802 & ~n85993;
  assign n85995 = ~n85988 & ~n85994;
  assign n85996 = ~n85802 & ~n85978;
  assign n85997 = n85995 & ~n85996;
  assign n85998 = n85796 & n85851;
  assign n85999 = ~n85796 & n85824;
  assign n86000 = ~n85998 & ~n85999;
  assign n86001 = n85997 & n86000;
  assign n86002 = n85790 & ~n86001;
  assign n86003 = n85796 & ~n85822;
  assign n86004 = ~n85815 & n86003;
  assign n86005 = ~n85981 & ~n86004;
  assign n86006 = ~n85802 & ~n86005;
  assign n86007 = ~n86002 & ~n86006;
  assign n86008 = ~n85790 & ~n85802;
  assign n86009 = ~n85796 & n85855;
  assign n86010 = ~n85851 & ~n86009;
  assign n86011 = ~n85836 & n86010;
  assign n86012 = n86008 & ~n86011;
  assign n86013 = n86007 & ~n86012;
  assign n86014 = n85986 & n86013;
  assign n86015 = ~pi2730 & ~n86014;
  assign n86016 = pi2730 & n85986;
  assign n86017 = n86007 & n86016;
  assign n86018 = ~n86012 & n86017;
  assign po2868 = n86015 | n86018;
  assign n86020 = n85490 & n85514;
  assign n86021 = ~n85499 & ~n85515;
  assign n86022 = ~n85470 & ~n86021;
  assign n86023 = ~n86020 & ~n86022;
  assign n86024 = ~n85484 & ~n85490;
  assign n86025 = ~n85464 & n86024;
  assign n86026 = n85464 & n85491;
  assign n86027 = ~n86025 & ~n86026;
  assign n86028 = n85477 & ~n85484;
  assign n86029 = n86027 & ~n86028;
  assign n86030 = ~n85528 & n86029;
  assign n86031 = n85470 & ~n86030;
  assign n86032 = n86023 & ~n86031;
  assign n86033 = ~n85524 & n86032;
  assign n86034 = n85458 & ~n86033;
  assign n86035 = ~n85464 & n85495;
  assign n86036 = n85527 & ~n86035;
  assign n86037 = n85470 & ~n86036;
  assign n86038 = ~n86034 & ~n86037;
  assign n86039 = n85484 & n85512;
  assign n86040 = ~n85490 & n86039;
  assign n86041 = n85464 & n85517;
  assign n86042 = ~n86040 & ~n86041;
  assign n86043 = n85477 & n85484;
  assign n86044 = n85464 & n86043;
  assign n86045 = ~n85509 & ~n86044;
  assign n86046 = ~n85470 & ~n86045;
  assign n86047 = ~n85470 & n85477;
  assign n86048 = ~n85484 & n86047;
  assign n86049 = ~n85464 & n86048;
  assign n86050 = ~n86046 & ~n86049;
  assign n86051 = n86042 & n86050;
  assign n86052 = ~n85458 & ~n86051;
  assign n86053 = ~n85477 & ~n85484;
  assign n86054 = ~n85470 & n86053;
  assign n86055 = n85464 & n86054;
  assign n86056 = ~n85464 & n85528;
  assign n86057 = ~n86055 & ~n86056;
  assign n86058 = ~n86052 & n86057;
  assign n86059 = n86038 & n86058;
  assign n86060 = ~pi2727 & ~n86059;
  assign n86061 = ~n86034 & ~n86056;
  assign n86062 = ~n86037 & n86061;
  assign n86063 = ~n86052 & ~n86055;
  assign n86064 = n86062 & n86063;
  assign n86065 = pi2727 & n86064;
  assign po2869 = n86060 | n86065;
  assign n86067 = ~n85356 & n85401;
  assign n86068 = ~n85369 & ~n86067;
  assign n86069 = ~n85330 & ~n86068;
  assign n86070 = n85363 & n85395;
  assign n86071 = ~n86069 & ~n86070;
  assign n86072 = ~n85622 & n86071;
  assign n86073 = n85356 & n85397;
  assign n86074 = ~n85401 & ~n86073;
  assign n86075 = ~n85388 & n86074;
  assign n86076 = ~n85330 & ~n86075;
  assign n86077 = n85382 & n86076;
  assign n86078 = n85330 & n85385;
  assign n86079 = ~n85358 & ~n85620;
  assign n86080 = ~n85599 & n86079;
  assign n86081 = ~n86078 & n86080;
  assign n86082 = n85382 & ~n86081;
  assign n86083 = n85330 & n85336;
  assign n86084 = n85349 & n86083;
  assign n86085 = n85342 & n86084;
  assign n86086 = n85356 & n85630;
  assign n86087 = ~n86085 & ~n86086;
  assign n86088 = ~n85366 & n86087;
  assign n86089 = n85349 & n85357;
  assign n86090 = n85350 & n85356;
  assign n86091 = ~n85394 & ~n86090;
  assign n86092 = ~n85330 & ~n86091;
  assign n86093 = ~n86089 & ~n86092;
  assign n86094 = n86088 & n86093;
  assign n86095 = ~n85382 & ~n86094;
  assign n86096 = ~n85356 & n86085;
  assign n86097 = ~n86095 & ~n86096;
  assign n86098 = ~n86082 & n86097;
  assign n86099 = ~n86077 & n86098;
  assign n86100 = n86072 & n86099;
  assign n86101 = pi2743 & ~n86100;
  assign n86102 = ~pi2743 & n86072;
  assign n86103 = n86099 & n86102;
  assign po2870 = n86101 | n86103;
  assign n86105 = ~n85668 & n85690;
  assign n86106 = ~n85965 & ~n86105;
  assign n86107 = n85674 & n86106;
  assign n86108 = n85668 & n85684;
  assign n86109 = ~n85674 & ~n86108;
  assign n86110 = ~n85684 & ~n85702;
  assign n86111 = ~n85683 & ~n86110;
  assign n86112 = n85668 & n85728;
  assign n86113 = ~n86111 & ~n86112;
  assign n86114 = ~n85656 & n85715;
  assign n86115 = n86113 & ~n86114;
  assign n86116 = n86109 & n86115;
  assign n86117 = ~n86107 & ~n86116;
  assign n86118 = n85668 & n86111;
  assign n86119 = ~n85954 & ~n86118;
  assign n86120 = ~n86117 & n86119;
  assign n86121 = n85650 & ~n86120;
  assign n86122 = n85674 & ~n86110;
  assign n86123 = ~n85668 & n86122;
  assign n86124 = ~n85705 & ~n85732;
  assign n86125 = n85668 & ~n86124;
  assign n86126 = n85674 & n86125;
  assign n86127 = n85683 & n86122;
  assign n86128 = ~n86126 & ~n86127;
  assign n86129 = ~n86123 & n86128;
  assign n86130 = ~n85650 & ~n86129;
  assign n86131 = ~n86121 & ~n86130;
  assign n86132 = n85674 & n85688;
  assign n86133 = ~n85674 & ~n86119;
  assign n86134 = ~n86132 & ~n86133;
  assign n86135 = ~n85674 & ~n86106;
  assign n86136 = ~n85688 & ~n86135;
  assign n86137 = ~n85650 & ~n86136;
  assign n86138 = n86134 & ~n86137;
  assign n86139 = n86131 & n86138;
  assign n86140 = pi2736 & ~n86139;
  assign n86141 = ~pi2736 & n86138;
  assign n86142 = ~n86130 & n86141;
  assign n86143 = ~n86121 & n86142;
  assign po2872 = n86140 | n86143;
  assign n86145 = ~n85809 & n86003;
  assign n86146 = ~n85824 & ~n86145;
  assign n86147 = ~n85802 & ~n86146;
  assign n86148 = n85796 & n85850;
  assign n86149 = ~n85796 & n85833;
  assign n86150 = ~n85809 & n86149;
  assign n86151 = ~n86148 & ~n86150;
  assign n86152 = n85802 & ~n86151;
  assign n86153 = ~n85796 & n85991;
  assign n86154 = ~n85862 & ~n86153;
  assign n86155 = ~n85981 & n86154;
  assign n86156 = ~n86152 & n86155;
  assign n86157 = ~n86147 & n86156;
  assign n86158 = ~n85835 & ~n85849;
  assign n86159 = n86157 & n86158;
  assign n86160 = n85790 & ~n86159;
  assign n86161 = n85837 & n85855;
  assign n86162 = n85982 & ~n86161;
  assign n86163 = n85802 & ~n86162;
  assign n86164 = ~n85796 & n85977;
  assign n86165 = ~n86163 & ~n86164;
  assign n86166 = n85815 & n86003;
  assign n86167 = n85796 & n85823;
  assign n86168 = ~n86166 & ~n86167;
  assign n86169 = n85802 & ~n86168;
  assign n86170 = n85802 & n85850;
  assign n86171 = ~n85796 & n86170;
  assign n86172 = ~n86169 & ~n86171;
  assign n86173 = n86165 & n86172;
  assign n86174 = ~n85790 & ~n86173;
  assign n86175 = ~n85991 & ~n85998;
  assign n86176 = ~n85842 & n86175;
  assign n86177 = n86008 & ~n86176;
  assign n86178 = ~n86174 & ~n86177;
  assign n86179 = ~n85835 & ~n85981;
  assign n86180 = ~n85802 & ~n86179;
  assign n86181 = n86178 & ~n86180;
  assign n86182 = ~n86160 & n86181;
  assign n86183 = ~pi2756 & n86182;
  assign n86184 = pi2756 & ~n86182;
  assign po2873 = n86183 | n86184;
  assign n86186 = ~n85464 & n85492;
  assign n86187 = ~n85495 & ~n86056;
  assign n86188 = n85464 & n85522;
  assign n86189 = ~n85464 & n85509;
  assign n86190 = ~n86188 & ~n86189;
  assign n86191 = n86187 & n86190;
  assign n86192 = ~n85470 & ~n86191;
  assign n86193 = n85464 & n85498;
  assign n86194 = ~n85515 & ~n86193;
  assign n86195 = ~n85525 & n86194;
  assign n86196 = n85470 & ~n86195;
  assign n86197 = n85464 & ~n85484;
  assign n86198 = n85490 & n86197;
  assign n86199 = ~n85477 & n86198;
  assign n86200 = ~n86196 & ~n86199;
  assign n86201 = ~n86192 & n86200;
  assign n86202 = ~n86186 & n86201;
  assign n86203 = ~n85458 & ~n86202;
  assign n86204 = n85464 & ~n85470;
  assign n86205 = n85528 & n86204;
  assign n86206 = ~n85470 & n85525;
  assign n86207 = ~n85470 & n85517;
  assign n86208 = ~n86206 & ~n86207;
  assign n86209 = ~n85464 & ~n86208;
  assign n86210 = ~n86205 & ~n86209;
  assign n86211 = n85464 & n85494;
  assign n86212 = ~n85464 & n85498;
  assign n86213 = ~n86211 & ~n86212;
  assign n86214 = ~n85523 & n86213;
  assign n86215 = ~n85495 & n86214;
  assign n86216 = n85470 & ~n86215;
  assign n86217 = ~n85464 & n85499;
  assign n86218 = ~n86216 & ~n86217;
  assign n86219 = ~n85464 & n85523;
  assign n86220 = ~n85510 & ~n86219;
  assign n86221 = n86218 & n86220;
  assign n86222 = n86210 & n86221;
  assign n86223 = n85458 & ~n86222;
  assign n86224 = ~n85470 & ~n85497;
  assign n86225 = ~n86223 & ~n86224;
  assign n86226 = ~n85526 & ~n86219;
  assign n86227 = n85470 & ~n86226;
  assign n86228 = n86225 & ~n86227;
  assign n86229 = ~n86203 & n86228;
  assign n86230 = pi2744 & ~n86229;
  assign n86231 = ~pi2744 & n86229;
  assign po2874 = n86230 | n86231;
  assign n86233 = ~n85241 & n85276;
  assign n86234 = ~n85255 & n86233;
  assign n86235 = n85255 & n85296;
  assign n86236 = ~n85281 & ~n86235;
  assign n86237 = n85229 & ~n86236;
  assign n86238 = ~n86234 & ~n86237;
  assign n86239 = ~n85229 & ~n85255;
  assign n86240 = ~n85241 & n86239;
  assign n86241 = ~n85247 & n86240;
  assign n86242 = n85241 & n85297;
  assign n86243 = ~n85247 & n86242;
  assign n86244 = ~n86241 & ~n86243;
  assign n86245 = ~n85229 & ~n85235;
  assign n86246 = n85257 & n86245;
  assign n86247 = n86244 & ~n86246;
  assign n86248 = ~n85259 & ~n85271;
  assign n86249 = ~n85311 & n86248;
  assign n86250 = n86247 & n86249;
  assign n86251 = n86238 & n86250;
  assign n86252 = ~n85294 & ~n86251;
  assign n86253 = ~n85258 & ~n85281;
  assign n86254 = n85255 & ~n86253;
  assign n86255 = ~n85247 & n85300;
  assign n86256 = ~n85235 & n85263;
  assign n86257 = ~n86255 & ~n86256;
  assign n86258 = ~n85235 & ~n85241;
  assign n86259 = n85255 & n86258;
  assign n86260 = n86257 & ~n86259;
  assign n86261 = n85229 & ~n86260;
  assign n86262 = ~n85255 & n85269;
  assign n86263 = n85249 & n85255;
  assign n86264 = ~n86262 & ~n86263;
  assign n86265 = ~n85229 & ~n86264;
  assign n86266 = ~n85255 & n85264;
  assign n86267 = ~n86265 & ~n86266;
  assign n86268 = ~n86261 & n86267;
  assign n86269 = ~n86254 & n86268;
  assign n86270 = n85294 & ~n86269;
  assign n86271 = n85229 & n85301;
  assign n86272 = ~n86270 & ~n86271;
  assign n86273 = ~n85229 & n86234;
  assign n86274 = n86272 & ~n86273;
  assign n86275 = ~n86252 & n86274;
  assign n86276 = ~pi2737 & ~n86275;
  assign n86277 = pi2737 & n86272;
  assign n86278 = ~n86252 & n86277;
  assign n86279 = ~n86273 & n86278;
  assign po2875 = n86276 | n86279;
  assign n86281 = pi6074 & ~pi9040;
  assign n86282 = pi6042 & pi9040;
  assign n86283 = ~n86281 & ~n86282;
  assign n86284 = pi2703 & n86283;
  assign n86285 = ~pi2703 & ~n86283;
  assign n86286 = ~n86284 & ~n86285;
  assign n86287 = pi6144 & ~pi9040;
  assign n86288 = pi6275 & pi9040;
  assign n86289 = ~n86287 & ~n86288;
  assign n86290 = ~pi2710 & ~n86289;
  assign n86291 = pi2710 & n86289;
  assign n86292 = ~n86290 & ~n86291;
  assign n86293 = pi5960 & pi9040;
  assign n86294 = pi6032 & ~pi9040;
  assign n86295 = ~n86293 & ~n86294;
  assign n86296 = ~pi2705 & n86295;
  assign n86297 = pi2705 & ~n86295;
  assign n86298 = ~n86296 & ~n86297;
  assign n86299 = n86292 & ~n86298;
  assign n86300 = n86286 & n86299;
  assign n86301 = ~n86292 & ~n86298;
  assign n86302 = ~n86286 & n86301;
  assign n86303 = ~n86300 & ~n86302;
  assign n86304 = pi6079 & ~pi9040;
  assign n86305 = pi6241 & pi9040;
  assign n86306 = ~n86304 & ~n86305;
  assign n86307 = ~pi2691 & n86306;
  assign n86308 = pi2691 & ~n86306;
  assign n86309 = ~n86307 & ~n86308;
  assign n86310 = n86286 & n86309;
  assign n86311 = n86292 & n86310;
  assign n86312 = n86303 & ~n86311;
  assign n86313 = pi6044 & ~pi9040;
  assign n86314 = pi5991 & pi9040;
  assign n86315 = ~n86313 & ~n86314;
  assign n86316 = ~pi2706 & n86315;
  assign n86317 = pi2706 & ~n86315;
  assign n86318 = ~n86316 & ~n86317;
  assign n86319 = pi6172 & pi9040;
  assign n86320 = pi6086 & ~pi9040;
  assign n86321 = ~n86319 & ~n86320;
  assign n86322 = ~pi2683 & ~n86321;
  assign n86323 = pi2683 & n86321;
  assign n86324 = ~n86322 & ~n86323;
  assign n86325 = n86318 & n86324;
  assign n86326 = ~n86312 & n86325;
  assign n86327 = ~n86292 & n86298;
  assign n86328 = n86286 & n86327;
  assign n86329 = ~n86309 & n86324;
  assign n86330 = n86328 & n86329;
  assign n86331 = n86286 & ~n86318;
  assign n86332 = ~n86292 & n86331;
  assign n86333 = ~n86298 & n86332;
  assign n86334 = n86292 & n86298;
  assign n86335 = ~n86309 & n86334;
  assign n86336 = ~n86286 & n86292;
  assign n86337 = ~n86335 & ~n86336;
  assign n86338 = ~n86318 & ~n86337;
  assign n86339 = ~n86333 & ~n86338;
  assign n86340 = n86324 & ~n86339;
  assign n86341 = ~n86330 & ~n86340;
  assign n86342 = ~n86286 & n86309;
  assign n86343 = ~n86292 & n86342;
  assign n86344 = n86298 & n86343;
  assign n86345 = ~n86286 & ~n86309;
  assign n86346 = n86292 & n86345;
  assign n86347 = ~n86344 & ~n86346;
  assign n86348 = ~n86318 & ~n86347;
  assign n86349 = n86341 & ~n86348;
  assign n86350 = ~n86309 & n86318;
  assign n86351 = n86334 & n86350;
  assign n86352 = n86286 & n86351;
  assign n86353 = ~n86299 & ~n86327;
  assign n86354 = n86310 & ~n86353;
  assign n86355 = ~n86298 & n86343;
  assign n86356 = ~n86354 & ~n86355;
  assign n86357 = ~n86286 & n86334;
  assign n86358 = n86309 & n86318;
  assign n86359 = n86357 & n86358;
  assign n86360 = n86345 & ~n86353;
  assign n86361 = n86286 & n86301;
  assign n86362 = ~n86309 & n86361;
  assign n86363 = ~n86360 & ~n86362;
  assign n86364 = ~n86359 & n86363;
  assign n86365 = n86356 & n86364;
  assign n86366 = ~n86352 & n86365;
  assign n86367 = n86309 & ~n86318;
  assign n86368 = n86286 & n86367;
  assign n86369 = n86298 & n86368;
  assign n86370 = n86366 & ~n86369;
  assign n86371 = ~n86324 & ~n86370;
  assign n86372 = n86349 & ~n86371;
  assign n86373 = ~n86326 & n86372;
  assign n86374 = ~pi2742 & ~n86373;
  assign n86375 = pi2742 & n86349;
  assign n86376 = ~n86326 & n86375;
  assign n86377 = ~n86371 & n86376;
  assign po2876 = n86374 | n86377;
  assign n86379 = n85668 & n85956;
  assign n86380 = n85674 & n86379;
  assign n86381 = n85715 & ~n86110;
  assign n86382 = ~n85733 & ~n86381;
  assign n86383 = ~n85954 & n86382;
  assign n86384 = ~n85674 & ~n86383;
  assign n86385 = n85668 & n85685;
  assign n86386 = ~n86384 & ~n86385;
  assign n86387 = n85683 & n85732;
  assign n86388 = ~n85668 & n85960;
  assign n86389 = ~n86387 & ~n86388;
  assign n86390 = ~n86108 & n86389;
  assign n86391 = n85674 & ~n86390;
  assign n86392 = n86386 & ~n86391;
  assign n86393 = n85650 & ~n86392;
  assign n86394 = ~n86380 & ~n86393;
  assign n86395 = ~n85668 & n85684;
  assign n86396 = ~n85710 & ~n86395;
  assign n86397 = n85674 & ~n86396;
  assign n86398 = ~n85734 & ~n86397;
  assign n86399 = ~n85706 & ~n86379;
  assign n86400 = n85668 & n85739;
  assign n86401 = ~n85960 & ~n86400;
  assign n86402 = ~n86387 & n86401;
  assign n86403 = ~n85674 & ~n86402;
  assign n86404 = ~n85668 & n85685;
  assign n86405 = ~n86403 & ~n86404;
  assign n86406 = n86399 & n86405;
  assign n86407 = n86398 & n86406;
  assign n86408 = ~n85650 & ~n86407;
  assign n86409 = ~n85720 & ~n86112;
  assign n86410 = ~n85674 & ~n86409;
  assign n86411 = ~n86408 & ~n86410;
  assign n86412 = n86394 & n86411;
  assign n86413 = pi2749 & n86412;
  assign n86414 = ~pi2749 & ~n86412;
  assign po2877 = n86413 | n86414;
  assign n86416 = ~n85502 & ~n86219;
  assign n86417 = ~n86199 & n86416;
  assign n86418 = ~n85470 & ~n86417;
  assign n86419 = ~n85513 & ~n85540;
  assign n86420 = ~n85510 & ~n86207;
  assign n86421 = ~n85492 & ~n86212;
  assign n86422 = n85470 & ~n86421;
  assign n86423 = ~n86056 & ~n86422;
  assign n86424 = n86420 & n86423;
  assign n86425 = n85458 & ~n86424;
  assign n86426 = ~n85484 & n85490;
  assign n86427 = ~n86028 & ~n86426;
  assign n86428 = n85464 & ~n86427;
  assign n86429 = ~n85519 & ~n85523;
  assign n86430 = n85470 & ~n86429;
  assign n86431 = n85464 & n85490;
  assign n86432 = ~n85499 & ~n86431;
  assign n86433 = ~n85491 & n86432;
  assign n86434 = ~n85470 & ~n86433;
  assign n86435 = ~n86430 & ~n86434;
  assign n86436 = ~n86428 & n86435;
  assign n86437 = ~n85458 & ~n86436;
  assign n86438 = ~n86425 & ~n86437;
  assign n86439 = n86419 & n86438;
  assign n86440 = ~n86418 & n86439;
  assign n86441 = ~pi2751 & ~n86440;
  assign n86442 = pi2751 & n86419;
  assign n86443 = ~n86418 & n86442;
  assign n86444 = n86438 & n86443;
  assign po2878 = n86441 | n86444;
  assign n86446 = n86286 & n86334;
  assign n86447 = ~n86318 & n86446;
  assign n86448 = n86309 & n86447;
  assign n86449 = ~n86318 & n86355;
  assign n86450 = ~n86448 & ~n86449;
  assign n86451 = n86286 & ~n86298;
  assign n86452 = ~n86309 & n86451;
  assign n86453 = ~n86335 & ~n86452;
  assign n86454 = ~n86318 & ~n86453;
  assign n86455 = ~n86334 & n86367;
  assign n86456 = ~n86286 & n86455;
  assign n86457 = ~n86454 & ~n86456;
  assign n86458 = n86318 & ~n86342;
  assign n86459 = ~n86353 & n86458;
  assign n86460 = ~n86359 & ~n86459;
  assign n86461 = ~n86355 & n86460;
  assign n86462 = n86457 & n86461;
  assign n86463 = n86324 & ~n86462;
  assign n86464 = n86450 & ~n86463;
  assign n86465 = n86300 & n86318;
  assign n86466 = ~n86309 & n86465;
  assign n86467 = n86318 & ~n86324;
  assign n86468 = ~n86335 & ~n86361;
  assign n86469 = n86342 & ~n86353;
  assign n86470 = n86468 & ~n86469;
  assign n86471 = n86467 & ~n86470;
  assign n86472 = n86302 & ~n86309;
  assign n86473 = ~n86298 & ~n86309;
  assign n86474 = ~n86286 & n86473;
  assign n86475 = ~n86309 & n86327;
  assign n86476 = ~n86474 & ~n86475;
  assign n86477 = n86309 & n86334;
  assign n86478 = ~n86328 & ~n86477;
  assign n86479 = n86476 & n86478;
  assign n86480 = ~n86318 & ~n86479;
  assign n86481 = ~n86472 & ~n86480;
  assign n86482 = ~n86324 & ~n86481;
  assign n86483 = ~n86471 & ~n86482;
  assign n86484 = ~n86466 & n86483;
  assign n86485 = n86464 & n86484;
  assign n86486 = pi2733 & ~n86485;
  assign n86487 = ~pi2733 & n86464;
  assign n86488 = n86484 & n86487;
  assign po2879 = n86486 | n86488;
  assign n86490 = ~n86475 & ~n86477;
  assign n86491 = ~n86318 & ~n86490;
  assign n86492 = ~n86449 & ~n86491;
  assign n86493 = n86324 & ~n86492;
  assign n86494 = ~n86286 & ~n86298;
  assign n86495 = ~n86299 & ~n86494;
  assign n86496 = n86309 & ~n86495;
  assign n86497 = ~n86446 & ~n86496;
  assign n86498 = n86318 & ~n86497;
  assign n86499 = ~n86469 & ~n86498;
  assign n86500 = ~n86309 & n86357;
  assign n86501 = ~n86292 & n86310;
  assign n86502 = ~n86309 & ~n86495;
  assign n86503 = ~n86501 & ~n86502;
  assign n86504 = ~n86318 & ~n86503;
  assign n86505 = ~n86500 & ~n86504;
  assign n86506 = n86499 & n86505;
  assign n86507 = ~n86324 & ~n86506;
  assign n86508 = n86286 & ~n86309;
  assign n86509 = ~n86299 & n86508;
  assign n86510 = n86324 & n86509;
  assign n86511 = n86299 & n86345;
  assign n86512 = ~n86318 & n86511;
  assign n86513 = n86286 & ~n86292;
  assign n86514 = n86350 & n86513;
  assign n86515 = ~n86512 & ~n86514;
  assign n86516 = ~n86510 & n86515;
  assign n86517 = ~n86328 & ~n86473;
  assign n86518 = n86325 & ~n86517;
  assign n86519 = n86516 & ~n86518;
  assign n86520 = ~n86507 & n86519;
  assign n86521 = ~n86493 & n86520;
  assign n86522 = pi2740 & ~n86521;
  assign n86523 = ~pi2740 & n86521;
  assign po2880 = n86522 | n86523;
  assign n86525 = ~n86333 & ~n86344;
  assign n86526 = ~n86286 & n86299;
  assign n86527 = ~n86446 & ~n86526;
  assign n86528 = ~n86318 & ~n86527;
  assign n86529 = n86525 & ~n86528;
  assign n86530 = n86309 & n86327;
  assign n86531 = ~n86300 & ~n86530;
  assign n86532 = ~n86357 & n86531;
  assign n86533 = n86318 & ~n86532;
  assign n86534 = n86529 & ~n86533;
  assign n86535 = ~n86324 & ~n86534;
  assign n86536 = ~n86309 & n86446;
  assign n86537 = n86301 & n86309;
  assign n86538 = ~n86475 & ~n86537;
  assign n86539 = n86318 & ~n86538;
  assign n86540 = ~n86536 & ~n86539;
  assign n86541 = ~n86318 & n86328;
  assign n86542 = n86303 & ~n86541;
  assign n86543 = ~n86357 & n86542;
  assign n86544 = n86309 & ~n86543;
  assign n86545 = n86540 & ~n86544;
  assign n86546 = n86324 & ~n86545;
  assign n86547 = ~n86535 & ~n86546;
  assign n86548 = ~n86286 & n86475;
  assign n86549 = ~n86362 & ~n86548;
  assign n86550 = ~n86318 & ~n86549;
  assign n86551 = n86318 & n86494;
  assign n86552 = ~n86309 & n86551;
  assign n86553 = ~n86550 & ~n86552;
  assign n86554 = n86547 & n86553;
  assign n86555 = ~pi2746 & ~n86554;
  assign n86556 = pi2746 & ~n86550;
  assign n86557 = n86547 & n86556;
  assign n86558 = ~n86552 & n86557;
  assign po2881 = n86555 | n86558;
  assign n86560 = ~n85256 & ~n85262;
  assign n86561 = ~n85229 & ~n86560;
  assign n86562 = ~n85318 & ~n86561;
  assign n86563 = n85235 & n85247;
  assign n86564 = n85229 & n86563;
  assign n86565 = n85255 & n86564;
  assign n86566 = n85255 & n85269;
  assign n86567 = ~n86563 & ~n86566;
  assign n86568 = ~n85235 & ~n85255;
  assign n86569 = ~n85247 & n86568;
  assign n86570 = n86567 & ~n86569;
  assign n86571 = n85229 & ~n86570;
  assign n86572 = ~n85265 & ~n86571;
  assign n86573 = ~n85294 & ~n86572;
  assign n86574 = ~n85229 & n85248;
  assign n86575 = n85255 & n86574;
  assign n86576 = ~n86246 & ~n86575;
  assign n86577 = ~n85294 & ~n86576;
  assign n86578 = ~n86573 & ~n86577;
  assign n86579 = ~n86565 & n86578;
  assign n86580 = ~n85281 & ~n85301;
  assign n86581 = ~n86256 & n86580;
  assign n86582 = ~n85229 & ~n86581;
  assign n86583 = ~n85255 & n85261;
  assign n86584 = ~n86233 & ~n86583;
  assign n86585 = n85229 & ~n86584;
  assign n86586 = ~n86582 & ~n86585;
  assign n86587 = ~n86255 & n86586;
  assign n86588 = ~n85271 & ~n85312;
  assign n86589 = n86587 & n86588;
  assign n86590 = n85294 & ~n86589;
  assign n86591 = n86579 & ~n86590;
  assign n86592 = n86562 & n86591;
  assign n86593 = ~pi2752 & ~n86592;
  assign n86594 = pi2752 & n86579;
  assign n86595 = n86562 & n86594;
  assign n86596 = ~n86590 & n86595;
  assign po2883 = n86593 | n86596;
  assign n86598 = ~n85796 & n85823;
  assign n86599 = ~n85989 & ~n86598;
  assign n86600 = ~n85802 & ~n86599;
  assign n86601 = n85802 & ~n85864;
  assign n86602 = ~n85875 & ~n86601;
  assign n86603 = ~n86600 & n86602;
  assign n86604 = n85790 & ~n86603;
  assign n86605 = ~n85802 & n85977;
  assign n86606 = ~n86604 & ~n86605;
  assign n86607 = ~n86153 & ~n86167;
  assign n86608 = n85802 & ~n86607;
  assign n86609 = n85802 & n85834;
  assign n86610 = n85809 & n86003;
  assign n86611 = n85815 & n86610;
  assign n86612 = ~n85802 & n85847;
  assign n86613 = ~n86149 & ~n86612;
  assign n86614 = ~n85815 & ~n86613;
  assign n86615 = ~n86150 & ~n86614;
  assign n86616 = ~n85981 & n86615;
  assign n86617 = ~n86611 & n86616;
  assign n86618 = ~n86609 & n86617;
  assign n86619 = ~n85790 & ~n86618;
  assign n86620 = ~n86608 & ~n86619;
  assign n86621 = n86606 & n86620;
  assign n86622 = pi2763 & ~n86621;
  assign n86623 = ~pi2763 & n86621;
  assign po2884 = n86622 | n86623;
  assign n86625 = ~n85312 & ~n86266;
  assign n86626 = n85229 & ~n86625;
  assign n86627 = ~n85294 & n85296;
  assign n86628 = ~n85229 & n86627;
  assign n86629 = n85247 & n86568;
  assign n86630 = ~n86258 & ~n86629;
  assign n86631 = ~n85264 & n86630;
  assign n86632 = n85229 & ~n86631;
  assign n86633 = ~n85255 & n85270;
  assign n86634 = ~n86632 & ~n86633;
  assign n86635 = ~n85294 & ~n86634;
  assign n86636 = ~n86628 & ~n86635;
  assign n86637 = ~n85259 & ~n85262;
  assign n86638 = ~n85255 & n86256;
  assign n86639 = ~n86235 & ~n86638;
  assign n86640 = n86637 & n86639;
  assign n86641 = ~n85229 & ~n86640;
  assign n86642 = n85235 & ~n85247;
  assign n86643 = ~n85229 & n86642;
  assign n86644 = n85255 & n86643;
  assign n86645 = ~n85255 & n86258;
  assign n86646 = ~n85262 & ~n86645;
  assign n86647 = ~n86263 & n86646;
  assign n86648 = ~n86644 & n86647;
  assign n86649 = n85229 & n85258;
  assign n86650 = n86648 & ~n86649;
  assign n86651 = n85294 & ~n86650;
  assign n86652 = ~n86641 & ~n86651;
  assign n86653 = n86636 & n86652;
  assign n86654 = ~n86626 & n86653;
  assign n86655 = pi2774 & n86654;
  assign n86656 = ~pi2774 & ~n86654;
  assign po2885 = n86655 | n86656;
  assign n86658 = pi6387 & ~pi9040;
  assign n86659 = ~pi6383 & pi9040;
  assign n86660 = ~n86658 & ~n86659;
  assign n86661 = pi2765 & n86660;
  assign n86662 = ~pi2765 & ~n86660;
  assign n86663 = ~n86661 & ~n86662;
  assign n86664 = pi6393 & ~pi9040;
  assign n86665 = pi6228 & pi9040;
  assign n86666 = ~n86664 & ~n86665;
  assign n86667 = ~pi2760 & n86666;
  assign n86668 = pi2760 & ~n86666;
  assign n86669 = ~n86667 & ~n86668;
  assign n86670 = pi6258 & pi9040;
  assign n86671 = pi6379 & ~pi9040;
  assign n86672 = ~n86670 & ~n86671;
  assign n86673 = pi2738 & n86672;
  assign n86674 = ~pi2738 & ~n86672;
  assign n86675 = ~n86673 & ~n86674;
  assign n86676 = n86669 & n86675;
  assign n86677 = pi6279 & pi9040;
  assign n86678 = pi6399 & ~pi9040;
  assign n86679 = ~n86677 & ~n86678;
  assign n86680 = ~pi2758 & ~n86679;
  assign n86681 = pi2758 & n86679;
  assign n86682 = ~n86680 & ~n86681;
  assign n86683 = pi6248 & pi9040;
  assign n86684 = pi6301 & ~pi9040;
  assign n86685 = ~n86683 & ~n86684;
  assign n86686 = pi2767 & n86685;
  assign n86687 = ~pi2767 & ~n86685;
  assign n86688 = ~n86686 & ~n86687;
  assign n86689 = ~n86682 & ~n86688;
  assign n86690 = n86676 & n86689;
  assign n86691 = pi6242 & pi9040;
  assign n86692 = pi6384 & ~pi9040;
  assign n86693 = ~n86691 & ~n86692;
  assign n86694 = ~pi2754 & n86693;
  assign n86695 = pi2754 & ~n86693;
  assign n86696 = ~n86694 & ~n86695;
  assign n86697 = ~n86669 & ~n86675;
  assign n86698 = ~n86696 & n86697;
  assign n86699 = n86682 & n86696;
  assign n86700 = ~n86675 & n86699;
  assign n86701 = n86669 & n86700;
  assign n86702 = ~n86698 & ~n86701;
  assign n86703 = ~n86669 & n86675;
  assign n86704 = n86682 & n86703;
  assign n86705 = n86702 & ~n86704;
  assign n86706 = ~n86688 & ~n86705;
  assign n86707 = ~n86669 & n86696;
  assign n86708 = ~n86682 & n86688;
  assign n86709 = n86707 & n86708;
  assign n86710 = n86696 & n86697;
  assign n86711 = ~n86682 & n86710;
  assign n86712 = ~n86709 & ~n86711;
  assign n86713 = ~n86706 & n86712;
  assign n86714 = ~n86690 & n86713;
  assign n86715 = n86676 & ~n86696;
  assign n86716 = ~n86682 & n86715;
  assign n86717 = ~n86696 & n86703;
  assign n86718 = n86682 & n86717;
  assign n86719 = ~n86716 & ~n86718;
  assign n86720 = n86714 & n86719;
  assign n86721 = ~n86663 & ~n86720;
  assign n86722 = ~n86682 & n86707;
  assign n86723 = n86675 & n86722;
  assign n86724 = ~n86715 & ~n86723;
  assign n86725 = ~n86688 & ~n86724;
  assign n86726 = n86676 & n86699;
  assign n86727 = ~n86682 & n86696;
  assign n86728 = ~n86675 & n86727;
  assign n86729 = n86669 & n86728;
  assign n86730 = ~n86726 & ~n86729;
  assign n86731 = ~n86669 & n86699;
  assign n86732 = ~n86682 & n86717;
  assign n86733 = ~n86731 & ~n86732;
  assign n86734 = n86688 & ~n86733;
  assign n86735 = n86730 & ~n86734;
  assign n86736 = ~n86725 & n86735;
  assign n86737 = n86663 & ~n86736;
  assign n86738 = ~n86669 & ~n86696;
  assign n86739 = n86682 & n86738;
  assign n86740 = n86669 & ~n86696;
  assign n86741 = ~n86682 & n86740;
  assign n86742 = ~n86739 & ~n86741;
  assign n86743 = ~n86688 & ~n86742;
  assign n86744 = n86669 & ~n86675;
  assign n86745 = ~n86696 & n86744;
  assign n86746 = n86682 & n86745;
  assign n86747 = ~n86726 & ~n86746;
  assign n86748 = ~n86710 & n86747;
  assign n86749 = n86688 & ~n86748;
  assign n86750 = ~n86743 & ~n86749;
  assign n86751 = ~n86675 & n86696;
  assign n86752 = n86688 & n86751;
  assign n86753 = ~n86682 & n86752;
  assign n86754 = n86750 & ~n86753;
  assign n86755 = ~n86737 & n86754;
  assign n86756 = ~n86721 & n86755;
  assign n86757 = ~pi2790 & ~n86756;
  assign n86758 = pi2790 & n86756;
  assign po2898 = n86757 | n86758;
  assign n86760 = pi6366 & pi9040;
  assign n86761 = pi6365 & ~pi9040;
  assign n86762 = ~n86760 & ~n86761;
  assign n86763 = ~pi2766 & ~n86762;
  assign n86764 = pi2766 & n86762;
  assign n86765 = ~n86763 & ~n86764;
  assign n86766 = pi6242 & ~pi9040;
  assign n86767 = pi6385 & pi9040;
  assign n86768 = ~n86766 & ~n86767;
  assign n86769 = ~pi2776 & ~n86768;
  assign n86770 = pi2776 & n86768;
  assign n86771 = ~n86769 & ~n86770;
  assign n86772 = pi6231 & ~pi9040;
  assign n86773 = pi6240 & pi9040;
  assign n86774 = ~n86772 & ~n86773;
  assign n86775 = pi2780 & n86774;
  assign n86776 = ~pi2780 & ~n86774;
  assign n86777 = ~n86775 & ~n86776;
  assign n86778 = pi6181 & pi9040;
  assign n86779 = pi6188 & ~pi9040;
  assign n86780 = ~n86778 & ~n86779;
  assign n86781 = ~pi2765 & n86780;
  assign n86782 = pi2765 & ~n86780;
  assign n86783 = ~n86781 & ~n86782;
  assign n86784 = ~n86777 & n86783;
  assign n86785 = pi6302 & ~pi9040;
  assign n86786 = pi6407 & pi9040;
  assign n86787 = ~n86785 & ~n86786;
  assign n86788 = ~pi2738 & n86787;
  assign n86789 = pi2738 & ~n86787;
  assign n86790 = ~n86788 & ~n86789;
  assign n86791 = n86784 & ~n86790;
  assign n86792 = n86771 & n86791;
  assign n86793 = n86771 & n86790;
  assign n86794 = n86783 & n86793;
  assign n86795 = n86777 & n86794;
  assign n86796 = ~n86792 & ~n86795;
  assign n86797 = n86777 & ~n86783;
  assign n86798 = n86790 & n86797;
  assign n86799 = ~n86771 & n86798;
  assign n86800 = n86784 & n86790;
  assign n86801 = ~n86771 & n86800;
  assign n86802 = ~n86799 & ~n86801;
  assign n86803 = n86796 & n86802;
  assign n86804 = n86765 & ~n86803;
  assign n86805 = ~n86777 & ~n86783;
  assign n86806 = n86790 & n86805;
  assign n86807 = n86771 & n86806;
  assign n86808 = n86777 & n86783;
  assign n86809 = n86790 & n86808;
  assign n86810 = ~n86807 & ~n86809;
  assign n86811 = n86765 & ~n86810;
  assign n86812 = ~n86765 & ~n86783;
  assign n86813 = ~n86771 & n86812;
  assign n86814 = n86777 & ~n86790;
  assign n86815 = n86771 & n86784;
  assign n86816 = ~n86814 & ~n86815;
  assign n86817 = ~n86765 & ~n86816;
  assign n86818 = ~n86813 & ~n86817;
  assign n86819 = ~n86790 & n86805;
  assign n86820 = ~n86771 & n86819;
  assign n86821 = n86818 & ~n86820;
  assign n86822 = n86771 & ~n86783;
  assign n86823 = ~n86790 & n86822;
  assign n86824 = n86777 & n86823;
  assign n86825 = n86821 & ~n86824;
  assign n86826 = ~n86811 & n86825;
  assign n86827 = pi6248 & ~pi9040;
  assign n86828 = pi6243 & pi9040;
  assign n86829 = ~n86827 & ~n86828;
  assign n86830 = ~pi2779 & ~n86829;
  assign n86831 = pi2779 & n86829;
  assign n86832 = ~n86830 & ~n86831;
  assign n86833 = ~n86826 & ~n86832;
  assign n86834 = ~n86783 & n86790;
  assign n86835 = ~n86765 & n86771;
  assign n86836 = n86832 & n86835;
  assign n86837 = n86834 & n86836;
  assign n86838 = ~n86771 & n86790;
  assign n86839 = n86783 & n86838;
  assign n86840 = ~n86765 & ~n86839;
  assign n86841 = ~n86797 & ~n86834;
  assign n86842 = ~n86771 & ~n86841;
  assign n86843 = n86771 & ~n86790;
  assign n86844 = ~n86777 & n86843;
  assign n86845 = ~n86791 & ~n86844;
  assign n86846 = ~n86842 & n86845;
  assign n86847 = n86765 & n86846;
  assign n86848 = ~n86840 & ~n86847;
  assign n86849 = n86783 & n86843;
  assign n86850 = n86777 & n86849;
  assign n86851 = ~n86848 & ~n86850;
  assign n86852 = n86832 & ~n86851;
  assign n86853 = ~n86837 & ~n86852;
  assign n86854 = ~n86833 & n86853;
  assign n86855 = ~n86804 & n86854;
  assign n86856 = ~n86765 & n86820;
  assign n86857 = n86855 & ~n86856;
  assign n86858 = pi2791 & ~n86857;
  assign n86859 = ~pi2791 & ~n86856;
  assign n86860 = n86854 & n86859;
  assign n86861 = ~n86804 & n86860;
  assign po2904 = n86858 | n86861;
  assign n86863 = n86682 & n86710;
  assign n86864 = ~n86729 & ~n86738;
  assign n86865 = n86688 & ~n86864;
  assign n86866 = ~n86723 & ~n86865;
  assign n86867 = ~n86863 & n86866;
  assign n86868 = ~n86688 & n86726;
  assign n86869 = ~n86716 & ~n86868;
  assign n86870 = ~n86746 & n86869;
  assign n86871 = n86867 & n86870;
  assign n86872 = n86663 & ~n86871;
  assign n86873 = n86696 & n86703;
  assign n86874 = n86682 & n86873;
  assign n86875 = ~n86701 & ~n86874;
  assign n86876 = ~n86682 & n86745;
  assign n86877 = ~n86711 & ~n86876;
  assign n86878 = n86675 & ~n86696;
  assign n86879 = ~n86669 & n86682;
  assign n86880 = ~n86878 & ~n86879;
  assign n86881 = ~n86751 & n86880;
  assign n86882 = ~n86688 & ~n86881;
  assign n86883 = n86676 & n86696;
  assign n86884 = n86688 & n86883;
  assign n86885 = n86682 & n86715;
  assign n86886 = ~n86884 & ~n86885;
  assign n86887 = ~n86882 & n86886;
  assign n86888 = n86877 & n86887;
  assign n86889 = n86875 & n86888;
  assign n86890 = ~n86663 & ~n86889;
  assign n86891 = ~n86872 & ~n86890;
  assign n86892 = pi2798 & ~n86891;
  assign n86893 = ~pi2798 & ~n86872;
  assign n86894 = ~n86890 & n86893;
  assign po2913 = n86892 | n86894;
  assign n86896 = pi6247 & ~pi9040;
  assign n86897 = pi6470 & pi9040;
  assign n86898 = ~n86896 & ~n86897;
  assign n86899 = ~pi2777 & ~n86898;
  assign n86900 = pi2777 & n86898;
  assign n86901 = ~n86899 & ~n86900;
  assign n86902 = pi6320 & pi9040;
  assign n86903 = pi6274 & ~pi9040;
  assign n86904 = ~n86902 & ~n86903;
  assign n86905 = ~pi2773 & n86904;
  assign n86906 = pi2773 & ~n86904;
  assign n86907 = ~n86905 & ~n86906;
  assign n86908 = pi6537 & pi9040;
  assign n86909 = pi6227 & ~pi9040;
  assign n86910 = ~n86908 & ~n86909;
  assign n86911 = ~pi2781 & ~n86910;
  assign n86912 = pi2781 & n86910;
  assign n86913 = ~n86911 & ~n86912;
  assign n86914 = pi6262 & pi9040;
  assign n86915 = pi6538 & ~pi9040;
  assign n86916 = ~n86914 & ~n86915;
  assign n86917 = ~pi2757 & ~n86916;
  assign n86918 = pi2757 & n86916;
  assign n86919 = ~n86917 & ~n86918;
  assign n86920 = pi6177 & ~pi9040;
  assign n86921 = pi6283 & pi9040;
  assign n86922 = ~n86920 & ~n86921;
  assign n86923 = ~pi2762 & ~n86922;
  assign n86924 = pi2762 & n86922;
  assign n86925 = ~n86923 & ~n86924;
  assign n86926 = ~n86919 & n86925;
  assign n86927 = n86913 & n86926;
  assign n86928 = ~n86907 & n86927;
  assign n86929 = pi6276 & pi9040;
  assign n86930 = pi6303 & ~pi9040;
  assign n86931 = ~n86929 & ~n86930;
  assign n86932 = ~pi2782 & ~n86931;
  assign n86933 = pi2782 & n86931;
  assign n86934 = ~n86932 & ~n86933;
  assign n86935 = n86919 & n86925;
  assign n86936 = ~n86907 & n86935;
  assign n86937 = ~n86913 & n86926;
  assign n86938 = n86907 & n86937;
  assign n86939 = ~n86936 & ~n86938;
  assign n86940 = ~n86934 & ~n86939;
  assign n86941 = ~n86928 & ~n86940;
  assign n86942 = ~n86919 & ~n86925;
  assign n86943 = ~n86913 & n86942;
  assign n86944 = n86934 & n86943;
  assign n86945 = n86926 & n86934;
  assign n86946 = ~n86907 & n86945;
  assign n86947 = ~n86944 & ~n86946;
  assign n86948 = n86941 & n86947;
  assign n86949 = n86919 & ~n86925;
  assign n86950 = n86913 & n86949;
  assign n86951 = ~n86907 & n86950;
  assign n86952 = n86913 & n86942;
  assign n86953 = n86907 & n86952;
  assign n86954 = ~n86951 & ~n86953;
  assign n86955 = n86948 & n86954;
  assign n86956 = n86901 & ~n86955;
  assign n86957 = ~n86901 & ~n86934;
  assign n86958 = ~n86907 & ~n86913;
  assign n86959 = ~n86919 & n86958;
  assign n86960 = ~n86913 & ~n86925;
  assign n86961 = ~n86959 & ~n86960;
  assign n86962 = n86957 & ~n86961;
  assign n86963 = n86907 & n86913;
  assign n86964 = n86925 & n86963;
  assign n86965 = ~n86919 & n86964;
  assign n86966 = n86907 & n86919;
  assign n86967 = ~n86913 & n86966;
  assign n86968 = ~n86965 & ~n86967;
  assign n86969 = ~n86907 & n86934;
  assign n86970 = n86913 & n86969;
  assign n86971 = ~n86926 & n86970;
  assign n86972 = n86934 & n86950;
  assign n86973 = ~n86971 & ~n86972;
  assign n86974 = n86968 & n86973;
  assign n86975 = ~n86901 & ~n86974;
  assign n86976 = ~n86913 & n86949;
  assign n86977 = ~n86934 & n86976;
  assign n86978 = n86907 & n86977;
  assign n86979 = n86913 & n86935;
  assign n86980 = n86907 & n86979;
  assign n86981 = ~n86953 & ~n86980;
  assign n86982 = ~n86934 & ~n86981;
  assign n86983 = ~n86978 & ~n86982;
  assign n86984 = n86934 & n86965;
  assign n86985 = n86983 & ~n86984;
  assign n86986 = ~n86975 & n86985;
  assign n86987 = ~n86962 & n86986;
  assign n86988 = ~n86956 & n86987;
  assign n86989 = ~n86913 & n86935;
  assign n86990 = n86907 & n86934;
  assign n86991 = n86989 & n86990;
  assign n86992 = n86988 & ~n86991;
  assign n86993 = ~pi2787 & ~n86992;
  assign n86994 = ~n86956 & ~n86991;
  assign n86995 = n86987 & n86994;
  assign n86996 = pi2787 & n86995;
  assign po2914 = n86993 | n86996;
  assign n86998 = ~n86682 & n86703;
  assign n86999 = ~n86876 & ~n86998;
  assign n87000 = n86688 & n86999;
  assign n87001 = ~n86676 & ~n86697;
  assign n87002 = ~n86696 & ~n87001;
  assign n87003 = n86682 & n86740;
  assign n87004 = n86669 & n86727;
  assign n87005 = n86682 & n86697;
  assign n87006 = ~n87004 & ~n87005;
  assign n87007 = ~n87003 & n87006;
  assign n87008 = ~n87002 & n87007;
  assign n87009 = ~n86688 & n87008;
  assign n87010 = ~n87000 & ~n87009;
  assign n87011 = n86682 & n87002;
  assign n87012 = ~n86874 & ~n87011;
  assign n87013 = ~n87010 & n87012;
  assign n87014 = n86663 & ~n87013;
  assign n87015 = n86688 & ~n87001;
  assign n87016 = ~n86682 & n87015;
  assign n87017 = ~n86717 & ~n86744;
  assign n87018 = n86682 & ~n87017;
  assign n87019 = n86688 & n87018;
  assign n87020 = n86696 & n87015;
  assign n87021 = ~n87019 & ~n87020;
  assign n87022 = ~n87016 & n87021;
  assign n87023 = ~n86663 & ~n87022;
  assign n87024 = ~n87014 & ~n87023;
  assign n87025 = n86688 & n86701;
  assign n87026 = ~n86688 & ~n87012;
  assign n87027 = ~n87025 & ~n87026;
  assign n87028 = ~n86688 & ~n86999;
  assign n87029 = ~n86701 & ~n87028;
  assign n87030 = ~n86663 & ~n87029;
  assign n87031 = n87027 & ~n87030;
  assign n87032 = n87024 & n87031;
  assign n87033 = pi2806 & ~n87032;
  assign n87034 = ~n87014 & n87031;
  assign n87035 = ~n87023 & n87034;
  assign n87036 = ~pi2806 & n87035;
  assign po2916 = n87033 | n87036;
  assign n87038 = pi6255 & pi9040;
  assign n87039 = pi6310 & ~pi9040;
  assign n87040 = ~n87038 & ~n87039;
  assign n87041 = ~pi2778 & ~n87040;
  assign n87042 = pi2778 & n87040;
  assign n87043 = ~n87041 & ~n87042;
  assign n87044 = pi6392 & pi9040;
  assign n87045 = pi6269 & ~pi9040;
  assign n87046 = ~n87044 & ~n87045;
  assign n87047 = pi2741 & n87046;
  assign n87048 = ~pi2741 & ~n87046;
  assign n87049 = ~n87047 & ~n87048;
  assign n87050 = pi6469 & pi9040;
  assign n87051 = pi6262 & ~pi9040;
  assign n87052 = ~n87050 & ~n87051;
  assign n87053 = pi2780 & n87052;
  assign n87054 = ~pi2780 & ~n87052;
  assign n87055 = ~n87053 & ~n87054;
  assign n87056 = pi6373 & ~pi9040;
  assign n87057 = pi6472 & pi9040;
  assign n87058 = ~n87056 & ~n87057;
  assign n87059 = ~pi2775 & n87058;
  assign n87060 = pi2775 & ~n87058;
  assign n87061 = ~n87059 & ~n87060;
  assign n87062 = n87055 & n87061;
  assign n87063 = ~n87049 & n87062;
  assign n87064 = pi6245 & pi9040;
  assign n87065 = pi6470 & ~pi9040;
  assign n87066 = ~n87064 & ~n87065;
  assign n87067 = ~pi2779 & ~n87066;
  assign n87068 = pi2779 & n87066;
  assign n87069 = ~n87067 & ~n87068;
  assign n87070 = n87055 & n87069;
  assign n87071 = n87049 & n87070;
  assign n87072 = ~n87061 & n87071;
  assign n87073 = ~n87063 & ~n87072;
  assign n87074 = n87049 & ~n87069;
  assign n87075 = ~n87055 & n87074;
  assign n87076 = ~n87061 & n87075;
  assign n87077 = n87073 & ~n87076;
  assign n87078 = ~n87043 & ~n87077;
  assign n87079 = pi6246 & ~pi9040;
  assign n87080 = pi6177 & pi9040;
  assign n87081 = ~n87079 & ~n87080;
  assign n87082 = ~pi2753 & ~n87081;
  assign n87083 = pi2753 & n87081;
  assign n87084 = ~n87082 & ~n87083;
  assign n87085 = n87043 & ~n87061;
  assign n87086 = n87074 & n87085;
  assign n87087 = n87055 & n87086;
  assign n87088 = n87043 & n87061;
  assign n87089 = n87049 & n87069;
  assign n87090 = n87088 & n87089;
  assign n87091 = n87063 & ~n87069;
  assign n87092 = ~n87049 & n87069;
  assign n87093 = n87055 & n87092;
  assign n87094 = n87043 & n87093;
  assign n87095 = ~n87061 & n87094;
  assign n87096 = ~n87091 & ~n87095;
  assign n87097 = ~n87090 & n87096;
  assign n87098 = ~n87087 & n87097;
  assign n87099 = n87061 & n87089;
  assign n87100 = ~n87055 & n87099;
  assign n87101 = n87098 & ~n87100;
  assign n87102 = ~n87084 & ~n87101;
  assign n87103 = ~n87049 & ~n87055;
  assign n87104 = n87069 & n87103;
  assign n87105 = ~n87043 & n87104;
  assign n87106 = ~n87061 & n87105;
  assign n87107 = n87062 & ~n87069;
  assign n87108 = ~n87049 & ~n87069;
  assign n87109 = n87061 & n87108;
  assign n87110 = ~n87107 & ~n87109;
  assign n87111 = ~n87043 & ~n87110;
  assign n87112 = ~n87106 & ~n87111;
  assign n87113 = ~n87084 & ~n87112;
  assign n87114 = ~n87102 & ~n87113;
  assign n87115 = ~n87078 & n87114;
  assign n87116 = ~n87055 & ~n87061;
  assign n87117 = n87043 & n87116;
  assign n87118 = n87108 & n87117;
  assign n87119 = ~n87055 & n87069;
  assign n87120 = n87088 & n87119;
  assign n87121 = n87061 & n87104;
  assign n87122 = ~n87043 & n87055;
  assign n87123 = n87069 & n87122;
  assign n87124 = ~n87061 & ~n87069;
  assign n87125 = ~n87055 & n87124;
  assign n87126 = ~n87123 & ~n87125;
  assign n87127 = ~n87121 & n87126;
  assign n87128 = ~n87075 & n87127;
  assign n87129 = n87043 & n87074;
  assign n87130 = n87061 & n87129;
  assign n87131 = ~n87061 & n87108;
  assign n87132 = n87049 & ~n87055;
  assign n87133 = ~n87131 & ~n87132;
  assign n87134 = n87043 & ~n87133;
  assign n87135 = ~n87130 & ~n87134;
  assign n87136 = n87128 & n87135;
  assign n87137 = n87084 & ~n87136;
  assign n87138 = ~n87120 & ~n87137;
  assign n87139 = ~n87118 & n87138;
  assign n87140 = n87115 & n87139;
  assign n87141 = pi2795 & n87140;
  assign n87142 = ~pi2795 & ~n87140;
  assign po2920 = n87141 | n87142;
  assign n87144 = n86907 & n86972;
  assign n87145 = n86913 & ~n86919;
  assign n87146 = n86969 & n87145;
  assign n87147 = ~n87144 & ~n87146;
  assign n87148 = n86907 & n86943;
  assign n87149 = ~n86907 & n86937;
  assign n87150 = ~n86907 & n86913;
  assign n87151 = n86925 & n87150;
  assign n87152 = n86919 & n87151;
  assign n87153 = ~n87149 & ~n87152;
  assign n87154 = ~n87148 & n87153;
  assign n87155 = ~n86934 & ~n87154;
  assign n87156 = n86907 & n86945;
  assign n87157 = n86919 & n86958;
  assign n87158 = ~n86976 & ~n87157;
  assign n87159 = n86934 & ~n87158;
  assign n87160 = ~n87156 & ~n87159;
  assign n87161 = ~n86934 & n86935;
  assign n87162 = n86907 & n87161;
  assign n87163 = ~n86934 & n86943;
  assign n87164 = ~n87162 & ~n87163;
  assign n87165 = n87160 & n87164;
  assign n87166 = n86913 & ~n86925;
  assign n87167 = ~n86907 & n87166;
  assign n87168 = ~n86919 & n87167;
  assign n87169 = n86919 & n86963;
  assign n87170 = ~n87148 & ~n87169;
  assign n87171 = ~n87168 & n87170;
  assign n87172 = n87165 & n87171;
  assign n87173 = ~n86901 & ~n87172;
  assign n87174 = n86934 & n86952;
  assign n87175 = ~n86991 & n87153;
  assign n87176 = ~n86965 & ~n86976;
  assign n87177 = ~n86907 & n86949;
  assign n87178 = n87176 & ~n87177;
  assign n87179 = ~n86934 & ~n87178;
  assign n87180 = n87175 & ~n87179;
  assign n87181 = ~n87174 & n87180;
  assign n87182 = n86901 & ~n87181;
  assign n87183 = ~n87173 & ~n87182;
  assign n87184 = ~n87155 & n87183;
  assign n87185 = n87147 & n87184;
  assign n87186 = pi2803 & ~n87185;
  assign n87187 = ~pi2803 & n87185;
  assign po2921 = n87186 | n87187;
  assign n87189 = ~n86925 & n86958;
  assign n87190 = n86919 & n87189;
  assign n87191 = ~n87148 & ~n87190;
  assign n87192 = n86934 & ~n87191;
  assign n87193 = ~n86934 & n86965;
  assign n87194 = ~n86965 & ~n86972;
  assign n87195 = ~n86919 & n86963;
  assign n87196 = ~n86967 & ~n87195;
  assign n87197 = ~n86934 & ~n87196;
  assign n87198 = ~n86907 & ~n86934;
  assign n87199 = n86942 & n87198;
  assign n87200 = ~n86913 & n87199;
  assign n87201 = ~n86913 & n86934;
  assign n87202 = n86925 & n87201;
  assign n87203 = ~n86919 & n87202;
  assign n87204 = ~n87152 & ~n87203;
  assign n87205 = ~n87200 & n87204;
  assign n87206 = ~n87197 & n87205;
  assign n87207 = n87194 & n87206;
  assign n87208 = n86901 & ~n87207;
  assign n87209 = ~n87144 & ~n87208;
  assign n87210 = ~n87193 & n87209;
  assign n87211 = ~n87192 & n87210;
  assign n87212 = ~n86944 & ~n87146;
  assign n87213 = n86934 & n86979;
  assign n87214 = n86907 & n86989;
  assign n87215 = ~n87213 & ~n87214;
  assign n87216 = ~n87148 & ~n87168;
  assign n87217 = ~n86913 & n86925;
  assign n87218 = ~n87177 & ~n87217;
  assign n87219 = ~n86934 & ~n87218;
  assign n87220 = n87216 & ~n87219;
  assign n87221 = n87215 & n87220;
  assign n87222 = n87212 & n87221;
  assign n87223 = ~n86901 & ~n87222;
  assign n87224 = n87211 & ~n87223;
  assign n87225 = ~pi2785 & ~n87224;
  assign n87226 = pi2785 & n87211;
  assign n87227 = ~n87223 & n87226;
  assign po2922 = n87225 | n87227;
  assign n87229 = pi6227 & pi9040;
  assign n87230 = pi6392 & ~pi9040;
  assign n87231 = ~n87229 & ~n87230;
  assign n87232 = pi2768 & n87231;
  assign n87233 = ~pi2768 & ~n87231;
  assign n87234 = ~n87232 & ~n87233;
  assign n87235 = pi6474 & ~pi9040;
  assign n87236 = pi6373 & pi9040;
  assign n87237 = ~n87235 & ~n87236;
  assign n87238 = pi2769 & n87237;
  assign n87239 = ~pi2769 & ~n87237;
  assign n87240 = ~n87238 & ~n87239;
  assign n87241 = pi6283 & ~pi9040;
  assign n87242 = pi6244 & pi9040;
  assign n87243 = ~n87241 & ~n87242;
  assign n87244 = ~pi2753 & n87243;
  assign n87245 = pi2753 & ~n87243;
  assign n87246 = ~n87244 & ~n87245;
  assign n87247 = ~n87240 & ~n87246;
  assign n87248 = pi6245 & ~pi9040;
  assign n87249 = pi6538 & pi9040;
  assign n87250 = ~n87248 & ~n87249;
  assign n87251 = ~pi2772 & ~n87250;
  assign n87252 = pi2772 & n87250;
  assign n87253 = ~n87251 & ~n87252;
  assign n87254 = pi6246 & pi9040;
  assign n87255 = pi6320 & ~pi9040;
  assign n87256 = ~n87254 & ~n87255;
  assign n87257 = ~pi2741 & n87256;
  assign n87258 = pi2741 & ~n87256;
  assign n87259 = ~n87257 & ~n87258;
  assign n87260 = n87253 & ~n87259;
  assign n87261 = n87247 & n87260;
  assign n87262 = n87253 & n87259;
  assign n87263 = n87246 & n87262;
  assign n87264 = ~n87261 & ~n87263;
  assign n87265 = ~n87234 & ~n87264;
  assign n87266 = pi6267 & pi9040;
  assign n87267 = pi6276 & ~pi9040;
  assign n87268 = ~n87266 & ~n87267;
  assign n87269 = ~pi2759 & ~n87268;
  assign n87270 = pi2759 & n87268;
  assign n87271 = ~n87269 & ~n87270;
  assign n87272 = n87234 & ~n87253;
  assign n87273 = ~n87246 & n87272;
  assign n87274 = n87247 & n87259;
  assign n87275 = n87240 & ~n87246;
  assign n87276 = ~n87259 & n87275;
  assign n87277 = ~n87274 & ~n87276;
  assign n87278 = ~n87240 & n87246;
  assign n87279 = ~n87259 & n87278;
  assign n87280 = n87253 & n87279;
  assign n87281 = n87277 & ~n87280;
  assign n87282 = n87234 & ~n87281;
  assign n87283 = ~n87273 & ~n87282;
  assign n87284 = n87240 & n87246;
  assign n87285 = n87259 & n87284;
  assign n87286 = n87253 & n87285;
  assign n87287 = n87283 & ~n87286;
  assign n87288 = ~n87253 & n87278;
  assign n87289 = ~n87259 & n87284;
  assign n87290 = ~n87288 & ~n87289;
  assign n87291 = ~n87234 & ~n87290;
  assign n87292 = n87259 & n87275;
  assign n87293 = ~n87253 & n87292;
  assign n87294 = ~n87291 & ~n87293;
  assign n87295 = n87287 & n87294;
  assign n87296 = n87271 & ~n87295;
  assign n87297 = ~n87265 & ~n87296;
  assign n87298 = n87234 & ~n87271;
  assign n87299 = ~n87290 & n87298;
  assign n87300 = n87259 & n87278;
  assign n87301 = ~n87292 & ~n87300;
  assign n87302 = n87253 & ~n87301;
  assign n87303 = ~n87261 & ~n87302;
  assign n87304 = ~n87271 & ~n87303;
  assign n87305 = ~n87299 & ~n87304;
  assign n87306 = ~n87234 & ~n87271;
  assign n87307 = n87247 & ~n87253;
  assign n87308 = ~n87285 & ~n87307;
  assign n87309 = ~n87246 & ~n87259;
  assign n87310 = n87308 & ~n87309;
  assign n87311 = n87306 & ~n87310;
  assign n87312 = n87305 & ~n87311;
  assign n87313 = n87297 & n87312;
  assign n87314 = ~pi2789 & ~n87313;
  assign n87315 = pi2789 & n87305;
  assign n87316 = n87297 & n87315;
  assign n87317 = ~n87311 & n87316;
  assign po2924 = n87314 | n87317;
  assign n87319 = n87055 & ~n87069;
  assign n87320 = ~n87100 & ~n87319;
  assign n87321 = ~n87124 & n87320;
  assign n87322 = n87043 & ~n87321;
  assign n87323 = ~n87043 & ~n87061;
  assign n87324 = n87069 & n87323;
  assign n87325 = n87055 & ~n87061;
  assign n87326 = n87049 & n87325;
  assign n87327 = n87061 & n87093;
  assign n87328 = ~n87326 & ~n87327;
  assign n87329 = ~n87055 & ~n87069;
  assign n87330 = ~n87043 & n87061;
  assign n87331 = n87329 & n87330;
  assign n87332 = n87328 & ~n87331;
  assign n87333 = ~n87324 & n87332;
  assign n87334 = ~n87322 & n87333;
  assign n87335 = n87084 & ~n87334;
  assign n87336 = n87055 & n87074;
  assign n87337 = n87061 & n87336;
  assign n87338 = ~n87049 & n87319;
  assign n87339 = ~n87061 & n87338;
  assign n87340 = ~n87337 & ~n87339;
  assign n87341 = n87043 & ~n87340;
  assign n87342 = ~n87335 & ~n87341;
  assign n87343 = ~n87061 & n87093;
  assign n87344 = ~n87071 & ~n87104;
  assign n87345 = n87043 & ~n87344;
  assign n87346 = ~n87343 & ~n87345;
  assign n87347 = ~n87076 & n87346;
  assign n87348 = ~n87084 & ~n87347;
  assign n87349 = ~n87089 & ~n87108;
  assign n87350 = ~n87055 & ~n87349;
  assign n87351 = ~n87109 & ~n87350;
  assign n87352 = ~n87043 & ~n87351;
  assign n87353 = ~n87084 & n87352;
  assign n87354 = ~n87348 & ~n87353;
  assign n87355 = n87342 & n87354;
  assign n87356 = pi2794 & ~n87355;
  assign n87357 = ~pi2794 & n87342;
  assign n87358 = n87354 & n87357;
  assign po2925 = n87356 | n87358;
  assign n87360 = pi6240 & ~pi9040;
  assign n87361 = pi6387 & pi9040;
  assign n87362 = ~n87360 & ~n87361;
  assign n87363 = ~pi2760 & ~n87362;
  assign n87364 = pi2760 & n87362;
  assign n87365 = ~n87363 & ~n87364;
  assign n87366 = pi6188 & pi9040;
  assign n87367 = pi6228 & ~pi9040;
  assign n87368 = ~n87366 & ~n87367;
  assign n87369 = pi2771 & n87368;
  assign n87370 = ~pi2771 & ~n87368;
  assign n87371 = ~n87369 & ~n87370;
  assign n87372 = pi6398 & pi9040;
  assign n87373 = pi6279 & ~pi9040;
  assign n87374 = ~n87372 & ~n87373;
  assign n87375 = pi2761 & n87374;
  assign n87376 = ~pi2761 & ~n87374;
  assign n87377 = ~n87375 & ~n87376;
  assign n87378 = pi6384 & pi9040;
  assign n87379 = pi6381 & ~pi9040;
  assign n87380 = ~n87378 & ~n87379;
  assign n87381 = ~pi2754 & n87380;
  assign n87382 = pi2754 & ~n87380;
  assign n87383 = ~n87381 & ~n87382;
  assign n87384 = pi6243 & ~pi9040;
  assign n87385 = pi6400 & pi9040;
  assign n87386 = ~n87384 & ~n87385;
  assign n87387 = pi2764 & n87386;
  assign n87388 = ~pi2764 & ~n87386;
  assign n87389 = ~n87387 & ~n87388;
  assign n87390 = ~n87383 & ~n87389;
  assign n87391 = n87377 & n87390;
  assign n87392 = n87383 & ~n87389;
  assign n87393 = ~n87377 & n87392;
  assign n87394 = ~n87391 & ~n87393;
  assign n87395 = ~n87371 & ~n87394;
  assign n87396 = pi6234 & pi9040;
  assign n87397 = pi6385 & ~pi9040;
  assign n87398 = ~n87396 & ~n87397;
  assign n87399 = pi2755 & n87398;
  assign n87400 = ~pi2755 & ~n87398;
  assign n87401 = ~n87399 & ~n87400;
  assign n87402 = ~n87383 & n87389;
  assign n87403 = n87377 & n87402;
  assign n87404 = n87401 & n87403;
  assign n87405 = ~n87395 & ~n87404;
  assign n87406 = ~n87377 & n87389;
  assign n87407 = n87389 & n87401;
  assign n87408 = ~n87406 & ~n87407;
  assign n87409 = n87377 & n87392;
  assign n87410 = n87408 & ~n87409;
  assign n87411 = n87371 & ~n87410;
  assign n87412 = n87405 & ~n87411;
  assign n87413 = ~n87365 & ~n87412;
  assign n87414 = ~n87377 & ~n87401;
  assign n87415 = ~n87383 & n87414;
  assign n87416 = ~n87389 & n87415;
  assign n87417 = n87371 & n87416;
  assign n87418 = ~n87383 & n87406;
  assign n87419 = ~n87401 & n87418;
  assign n87420 = ~n87371 & n87419;
  assign n87421 = n87383 & n87389;
  assign n87422 = n87377 & n87421;
  assign n87423 = ~n87401 & n87422;
  assign n87424 = ~n87371 & n87423;
  assign n87425 = ~n87420 & ~n87424;
  assign n87426 = ~n87417 & n87425;
  assign n87427 = n87371 & ~n87377;
  assign n87428 = ~n87383 & n87427;
  assign n87429 = ~n87389 & n87428;
  assign n87430 = n87377 & ~n87401;
  assign n87431 = n87383 & n87430;
  assign n87432 = ~n87416 & ~n87431;
  assign n87433 = n87389 & n87430;
  assign n87434 = n87371 & n87433;
  assign n87435 = n87391 & n87401;
  assign n87436 = ~n87371 & n87406;
  assign n87437 = ~n87435 & ~n87436;
  assign n87438 = n87393 & n87401;
  assign n87439 = n87437 & ~n87438;
  assign n87440 = ~n87434 & n87439;
  assign n87441 = n87432 & n87440;
  assign n87442 = ~n87429 & n87441;
  assign n87443 = n87365 & ~n87442;
  assign n87444 = n87426 & ~n87443;
  assign n87445 = ~n87413 & n87444;
  assign n87446 = ~pi2807 & ~n87445;
  assign n87447 = pi2807 & n87426;
  assign n87448 = ~n87413 & n87447;
  assign n87449 = ~n87443 & n87448;
  assign po2927 = n87446 | n87449;
  assign n87451 = ~n86682 & n86697;
  assign n87452 = ~n86873 & ~n87451;
  assign n87453 = n86688 & ~n87452;
  assign n87454 = ~n86746 & ~n87453;
  assign n87455 = n86682 & n86883;
  assign n87456 = ~n86718 & ~n87455;
  assign n87457 = ~n86682 & n86698;
  assign n87458 = n86682 & n86751;
  assign n87459 = ~n86878 & ~n87458;
  assign n87460 = n86696 & n86744;
  assign n87461 = n87459 & ~n87460;
  assign n87462 = ~n86688 & ~n87461;
  assign n87463 = ~n87457 & ~n87462;
  assign n87464 = n87456 & n87463;
  assign n87465 = n87454 & n87464;
  assign n87466 = ~n86663 & ~n87465;
  assign n87467 = ~n86732 & ~n87003;
  assign n87468 = ~n86688 & ~n87467;
  assign n87469 = ~n87466 & ~n87468;
  assign n87470 = n86688 & n87455;
  assign n87471 = n86727 & ~n87001;
  assign n87472 = ~n86745 & ~n87471;
  assign n87473 = ~n86874 & n87472;
  assign n87474 = ~n86688 & ~n87473;
  assign n87475 = n86682 & n86698;
  assign n87476 = ~n87474 & ~n87475;
  assign n87477 = ~n86682 & n86878;
  assign n87478 = ~n87460 & ~n87477;
  assign n87479 = ~n87005 & n87478;
  assign n87480 = n86688 & ~n87479;
  assign n87481 = n87476 & ~n87480;
  assign n87482 = n86663 & ~n87481;
  assign n87483 = ~n87470 & ~n87482;
  assign n87484 = n87469 & n87483;
  assign n87485 = pi2815 & n87484;
  assign n87486 = ~pi2815 & ~n87484;
  assign po2929 = n87485 | n87486;
  assign n87488 = pi6181 & ~pi9040;
  assign n87489 = pi6381 & pi9040;
  assign n87490 = ~n87488 & ~n87489;
  assign n87491 = ~pi2764 & ~n87490;
  assign n87492 = pi2764 & n87490;
  assign n87493 = ~n87491 & ~n87492;
  assign n87494 = pi6231 & pi9040;
  assign n87495 = pi6400 & ~pi9040;
  assign n87496 = ~n87494 & ~n87495;
  assign n87497 = pi2783 & n87496;
  assign n87498 = ~pi2783 & ~n87496;
  assign n87499 = ~n87497 & ~n87498;
  assign n87500 = pi6302 & pi9040;
  assign n87501 = pi6398 & ~pi9040;
  assign n87502 = ~n87500 & ~n87501;
  assign n87503 = ~pi2777 & ~n87502;
  assign n87504 = pi2777 & n87502;
  assign n87505 = ~n87503 & ~n87504;
  assign n87506 = pi6379 & pi9040;
  assign n87507 = pi6234 & ~pi9040;
  assign n87508 = ~n87506 & ~n87507;
  assign n87509 = ~pi2762 & ~n87508;
  assign n87510 = pi2762 & n87508;
  assign n87511 = ~n87509 & ~n87510;
  assign n87512 = pi6301 & pi9040;
  assign n87513 = pi6273 & ~pi9040;
  assign n87514 = ~n87512 & ~n87513;
  assign n87515 = pi2761 & n87514;
  assign n87516 = ~pi2761 & ~n87514;
  assign n87517 = ~n87515 & ~n87516;
  assign n87518 = n87511 & ~n87517;
  assign n87519 = n87505 & n87518;
  assign n87520 = n87499 & n87519;
  assign n87521 = ~n87499 & n87511;
  assign n87522 = n87517 & n87521;
  assign n87523 = pi6264 & pi9040;
  assign n87524 = pi6366 & ~pi9040;
  assign n87525 = ~n87523 & ~n87524;
  assign n87526 = ~pi2748 & n87525;
  assign n87527 = pi2748 & ~n87525;
  assign n87528 = ~n87526 & ~n87527;
  assign n87529 = ~n87505 & n87521;
  assign n87530 = n87505 & n87517;
  assign n87531 = ~n87511 & n87530;
  assign n87532 = ~n87529 & ~n87531;
  assign n87533 = n87528 & ~n87532;
  assign n87534 = ~n87522 & ~n87533;
  assign n87535 = n87511 & n87530;
  assign n87536 = ~n87511 & ~n87517;
  assign n87537 = ~n87499 & n87536;
  assign n87538 = ~n87505 & ~n87517;
  assign n87539 = n87499 & n87538;
  assign n87540 = ~n87537 & ~n87539;
  assign n87541 = ~n87505 & ~n87511;
  assign n87542 = n87540 & ~n87541;
  assign n87543 = ~n87535 & n87542;
  assign n87544 = ~n87528 & ~n87543;
  assign n87545 = n87534 & ~n87544;
  assign n87546 = ~n87520 & n87545;
  assign n87547 = n87493 & ~n87546;
  assign n87548 = ~n87505 & n87517;
  assign n87549 = ~n87511 & n87548;
  assign n87550 = ~n87499 & n87549;
  assign n87551 = ~n87511 & n87538;
  assign n87552 = n87499 & n87551;
  assign n87553 = ~n87520 & ~n87552;
  assign n87554 = ~n87550 & n87553;
  assign n87555 = ~n87528 & ~n87554;
  assign n87556 = ~n87547 & ~n87555;
  assign n87557 = ~n87499 & n87535;
  assign n87558 = ~n87511 & n87528;
  assign n87559 = n87505 & n87558;
  assign n87560 = n87499 & n87559;
  assign n87561 = n87511 & n87548;
  assign n87562 = n87499 & n87561;
  assign n87563 = n87518 & ~n87528;
  assign n87564 = ~n87499 & n87563;
  assign n87565 = ~n87562 & ~n87564;
  assign n87566 = ~n87505 & n87511;
  assign n87567 = n87499 & n87566;
  assign n87568 = n87505 & ~n87517;
  assign n87569 = ~n87511 & n87568;
  assign n87570 = ~n87567 & ~n87569;
  assign n87571 = n87528 & ~n87570;
  assign n87572 = ~n87505 & n87528;
  assign n87573 = ~n87511 & n87572;
  assign n87574 = ~n87499 & n87573;
  assign n87575 = ~n87571 & ~n87574;
  assign n87576 = n87565 & n87575;
  assign n87577 = ~n87493 & ~n87576;
  assign n87578 = ~n87560 & ~n87577;
  assign n87579 = ~n87557 & n87578;
  assign n87580 = n87556 & n87579;
  assign n87581 = ~pi2784 & ~n87580;
  assign n87582 = ~n87547 & ~n87557;
  assign n87583 = ~n87555 & n87582;
  assign n87584 = n87578 & n87583;
  assign n87585 = pi2784 & n87584;
  assign po2930 = n87581 | n87585;
  assign n87587 = ~n87365 & ~n87371;
  assign n87588 = n87377 & ~n87389;
  assign n87589 = ~n87401 & n87588;
  assign n87590 = n87401 & n87422;
  assign n87591 = ~n87401 & n87402;
  assign n87592 = ~n87590 & ~n87591;
  assign n87593 = ~n87589 & n87592;
  assign n87594 = n87587 & ~n87593;
  assign n87595 = n87383 & n87414;
  assign n87596 = n87401 & n87409;
  assign n87597 = ~n87595 & ~n87596;
  assign n87598 = ~n87377 & n87421;
  assign n87599 = ~n87403 & ~n87598;
  assign n87600 = n87597 & n87599;
  assign n87601 = n87371 & ~n87600;
  assign n87602 = ~n87377 & n87390;
  assign n87603 = n87401 & n87602;
  assign n87604 = ~n87601 & ~n87603;
  assign n87605 = ~n87365 & ~n87604;
  assign n87606 = ~n87594 & ~n87605;
  assign n87607 = n87371 & ~n87401;
  assign n87608 = n87377 & n87607;
  assign n87609 = ~n87383 & n87608;
  assign n87610 = ~n87401 & n87598;
  assign n87611 = ~n87609 & ~n87610;
  assign n87612 = ~n87392 & ~n87402;
  assign n87613 = n87401 & ~n87612;
  assign n87614 = ~n87393 & ~n87613;
  assign n87615 = ~n87371 & ~n87614;
  assign n87616 = ~n87391 & ~n87589;
  assign n87617 = ~n87590 & n87616;
  assign n87618 = n87371 & ~n87617;
  assign n87619 = ~n87615 & ~n87618;
  assign n87620 = ~n87371 & ~n87401;
  assign n87621 = n87421 & n87620;
  assign n87622 = n87401 & n87418;
  assign n87623 = ~n87438 & ~n87622;
  assign n87624 = ~n87416 & n87623;
  assign n87625 = ~n87621 & n87624;
  assign n87626 = n87619 & n87625;
  assign n87627 = n87365 & ~n87626;
  assign n87628 = n87611 & ~n87627;
  assign n87629 = n87606 & n87628;
  assign n87630 = pi2793 & ~n87629;
  assign n87631 = ~pi2793 & n87611;
  assign n87632 = n87606 & n87631;
  assign n87633 = ~n87627 & n87632;
  assign po2931 = n87630 | n87633;
  assign n87635 = n87061 & n87075;
  assign n87636 = ~n87327 & ~n87635;
  assign n87637 = ~n87043 & ~n87636;
  assign n87638 = n87071 & n87323;
  assign n87639 = ~n87637 & ~n87638;
  assign n87640 = ~n87120 & n87639;
  assign n87641 = ~n87061 & n87104;
  assign n87642 = ~n87075 & ~n87641;
  assign n87643 = ~n87338 & n87642;
  assign n87644 = ~n87043 & ~n87643;
  assign n87645 = n87084 & n87644;
  assign n87646 = n87043 & n87055;
  assign n87647 = ~n87049 & n87646;
  assign n87648 = ~n87069 & n87647;
  assign n87649 = n87061 & n87648;
  assign n87650 = n87043 & n87336;
  assign n87651 = ~n87100 & ~n87118;
  assign n87652 = ~n87095 & n87651;
  assign n87653 = ~n87650 & n87652;
  assign n87654 = n87084 & ~n87653;
  assign n87655 = ~n87061 & n87129;
  assign n87656 = ~n87648 & ~n87655;
  assign n87657 = ~n87326 & n87656;
  assign n87658 = ~n87055 & n87061;
  assign n87659 = ~n87049 & n87658;
  assign n87660 = ~n87061 & n87089;
  assign n87661 = ~n87070 & ~n87660;
  assign n87662 = ~n87043 & ~n87661;
  assign n87663 = ~n87659 & ~n87662;
  assign n87664 = n87657 & n87663;
  assign n87665 = ~n87084 & ~n87664;
  assign n87666 = ~n87654 & ~n87665;
  assign n87667 = ~n87649 & n87666;
  assign n87668 = ~n87645 & n87667;
  assign n87669 = n87640 & n87668;
  assign n87670 = pi2799 & ~n87669;
  assign n87671 = ~pi2799 & n87640;
  assign n87672 = n87668 & n87671;
  assign po2932 = n87670 | n87672;
  assign n87674 = ~n87061 & n87350;
  assign n87675 = ~n87103 & ~n87336;
  assign n87676 = ~n87043 & ~n87675;
  assign n87677 = ~n87674 & ~n87676;
  assign n87678 = ~n87049 & n87325;
  assign n87679 = ~n87132 & ~n87678;
  assign n87680 = ~n87338 & n87679;
  assign n87681 = n87043 & ~n87680;
  assign n87682 = n87677 & ~n87681;
  assign n87683 = n87061 & n87071;
  assign n87684 = n87682 & ~n87683;
  assign n87685 = ~n87084 & ~n87684;
  assign n87686 = n87088 & ~n87675;
  assign n87687 = ~n87075 & ~n87104;
  assign n87688 = ~n87071 & ~n87338;
  assign n87689 = n87687 & n87688;
  assign n87690 = ~n87061 & ~n87689;
  assign n87691 = ~n87686 & ~n87690;
  assign n87692 = ~n87327 & n87691;
  assign n87693 = n87084 & ~n87692;
  assign n87694 = ~n87685 & ~n87693;
  assign n87695 = ~n87061 & n87336;
  assign n87696 = ~n87683 & ~n87695;
  assign n87697 = ~n87043 & ~n87696;
  assign n87698 = n87694 & ~n87697;
  assign n87699 = pi2788 & ~n87698;
  assign n87700 = ~pi2788 & ~n87697;
  assign n87701 = ~n87693 & n87700;
  assign n87702 = ~n87685 & n87701;
  assign po2933 = n87699 | n87702;
  assign n87704 = ~n86792 & ~n86799;
  assign n87705 = ~n86765 & ~n87704;
  assign n87706 = ~n86856 & ~n87705;
  assign n87707 = ~n86777 & n86790;
  assign n87708 = n86765 & n87707;
  assign n87709 = n86771 & n87708;
  assign n87710 = n86771 & n86805;
  assign n87711 = ~n87707 & ~n87710;
  assign n87712 = ~n86771 & ~n86790;
  assign n87713 = n86777 & n87712;
  assign n87714 = n87711 & ~n87713;
  assign n87715 = n86765 & ~n87714;
  assign n87716 = ~n86795 & ~n87715;
  assign n87717 = ~n86832 & ~n87716;
  assign n87718 = ~n86765 & n86797;
  assign n87719 = n86771 & n87718;
  assign n87720 = ~n86765 & n86791;
  assign n87721 = ~n87719 & ~n87720;
  assign n87722 = ~n86832 & ~n87721;
  assign n87723 = ~n87717 & ~n87722;
  assign n87724 = ~n87709 & n87723;
  assign n87725 = n86777 & n86838;
  assign n87726 = ~n86819 & ~n86839;
  assign n87727 = ~n86790 & n86808;
  assign n87728 = n87726 & ~n87727;
  assign n87729 = ~n86765 & ~n87728;
  assign n87730 = ~n86771 & n86791;
  assign n87731 = ~n86783 & n86814;
  assign n87732 = ~n87730 & ~n87731;
  assign n87733 = n86765 & ~n87732;
  assign n87734 = ~n87729 & ~n87733;
  assign n87735 = ~n87725 & n87734;
  assign n87736 = ~n86807 & ~n86850;
  assign n87737 = n87735 & n87736;
  assign n87738 = n86832 & ~n87737;
  assign n87739 = n87724 & ~n87738;
  assign n87740 = n87706 & n87739;
  assign n87741 = ~pi2829 & ~n87740;
  assign n87742 = pi2829 & n87724;
  assign n87743 = n87706 & n87742;
  assign n87744 = ~n87738 & n87743;
  assign po2934 = n87741 | n87744;
  assign n87746 = ~n87499 & n87528;
  assign n87747 = n87505 & n87746;
  assign n87748 = n87511 & n87538;
  assign n87749 = n87499 & n87748;
  assign n87750 = n87499 & n87549;
  assign n87751 = ~n87749 & ~n87750;
  assign n87752 = ~n87499 & ~n87511;
  assign n87753 = ~n87517 & n87752;
  assign n87754 = ~n87505 & n87753;
  assign n87755 = ~n87531 & ~n87754;
  assign n87756 = ~n87528 & ~n87755;
  assign n87757 = n87751 & ~n87756;
  assign n87758 = ~n87747 & n87757;
  assign n87759 = n87493 & ~n87758;
  assign n87760 = n87499 & n87569;
  assign n87761 = n87528 & n87760;
  assign n87762 = ~n87499 & ~n87528;
  assign n87763 = n87569 & n87762;
  assign n87764 = ~n87529 & ~n87763;
  assign n87765 = ~n87531 & ~n87561;
  assign n87766 = ~n87499 & n87548;
  assign n87767 = n87765 & ~n87766;
  assign n87768 = n87528 & ~n87767;
  assign n87769 = ~n87528 & n87535;
  assign n87770 = n87553 & ~n87769;
  assign n87771 = ~n87768 & n87770;
  assign n87772 = n87764 & n87771;
  assign n87773 = ~n87493 & ~n87772;
  assign n87774 = ~n87761 & ~n87773;
  assign n87775 = ~n87759 & n87774;
  assign n87776 = n87561 & n87762;
  assign n87777 = n87499 & n87563;
  assign n87778 = ~n87776 & ~n87777;
  assign n87779 = ~n87528 & n87750;
  assign n87780 = n87778 & ~n87779;
  assign n87781 = n87775 & n87780;
  assign n87782 = ~pi2786 & ~n87781;
  assign n87783 = pi2786 & n87780;
  assign n87784 = n87774 & n87783;
  assign n87785 = ~n87759 & n87784;
  assign po2935 = n87782 | n87785;
  assign n87787 = n87401 & n87588;
  assign n87788 = ~n87403 & ~n87787;
  assign n87789 = ~n87610 & n87788;
  assign n87790 = n87371 & ~n87789;
  assign n87791 = ~n87377 & ~n87389;
  assign n87792 = ~n87421 & ~n87791;
  assign n87793 = n87401 & ~n87792;
  assign n87794 = n87391 & ~n87401;
  assign n87795 = ~n87793 & ~n87794;
  assign n87796 = ~n87419 & n87795;
  assign n87797 = ~n87371 & ~n87796;
  assign n87798 = ~n87790 & ~n87797;
  assign n87799 = n87365 & ~n87798;
  assign n87800 = ~n87389 & n87607;
  assign n87801 = ~n87433 & ~n87787;
  assign n87802 = ~n87371 & ~n87801;
  assign n87803 = ~n87621 & ~n87802;
  assign n87804 = ~n87423 & ~n87622;
  assign n87805 = n87371 & n87401;
  assign n87806 = n87406 & n87805;
  assign n87807 = ~n87429 & ~n87806;
  assign n87808 = n87804 & n87807;
  assign n87809 = n87803 & n87808;
  assign n87810 = ~n87800 & n87809;
  assign n87811 = ~n87365 & ~n87810;
  assign n87812 = ~n87371 & n87393;
  assign n87813 = ~n87401 & n87812;
  assign n87814 = ~n87424 & ~n87813;
  assign n87815 = ~n87417 & n87814;
  assign n87816 = ~n87389 & n87431;
  assign n87817 = n87401 & n87402;
  assign n87818 = ~n87816 & ~n87817;
  assign n87819 = n87371 & ~n87818;
  assign n87820 = n87815 & ~n87819;
  assign n87821 = ~n87811 & n87820;
  assign n87822 = ~n87799 & n87821;
  assign n87823 = ~pi2804 & n87822;
  assign n87824 = pi2804 & ~n87822;
  assign po2936 = n87823 | n87824;
  assign n87826 = ~n87234 & n87253;
  assign n87827 = ~n87278 & ~n87292;
  assign n87828 = n87826 & ~n87827;
  assign n87829 = ~n87234 & n87259;
  assign n87830 = n87278 & n87829;
  assign n87831 = ~n87828 & ~n87830;
  assign n87832 = n87271 & ~n87831;
  assign n87833 = ~n87253 & n87276;
  assign n87834 = ~n87253 & ~n87259;
  assign n87835 = ~n87309 & ~n87834;
  assign n87836 = n87234 & ~n87835;
  assign n87837 = ~n87253 & n87259;
  assign n87838 = ~n87240 & n87837;
  assign n87839 = ~n87246 & n87838;
  assign n87840 = ~n87836 & ~n87839;
  assign n87841 = ~n87833 & n87840;
  assign n87842 = n87271 & ~n87841;
  assign n87843 = ~n87832 & ~n87842;
  assign n87844 = n87240 & n87260;
  assign n87845 = n87246 & n87844;
  assign n87846 = ~n87253 & n87285;
  assign n87847 = ~n87845 & ~n87846;
  assign n87848 = ~n87234 & ~n87847;
  assign n87849 = n87253 & n87300;
  assign n87850 = ~n87253 & n87309;
  assign n87851 = ~n87849 & ~n87850;
  assign n87852 = n87234 & ~n87851;
  assign n87853 = ~n87247 & ~n87309;
  assign n87854 = n87253 & ~n87853;
  assign n87855 = ~n87285 & ~n87854;
  assign n87856 = ~n87234 & ~n87855;
  assign n87857 = n87240 & ~n87253;
  assign n87858 = n87829 & n87857;
  assign n87859 = ~n87240 & ~n87259;
  assign n87860 = ~n87285 & ~n87859;
  assign n87861 = ~n87253 & ~n87860;
  assign n87862 = n87234 & n87253;
  assign n87863 = n87275 & n87862;
  assign n87864 = n87259 & n87863;
  assign n87865 = ~n87861 & ~n87864;
  assign n87866 = ~n87858 & n87865;
  assign n87867 = ~n87856 & n87866;
  assign n87868 = ~n87845 & n87867;
  assign n87869 = ~n87271 & ~n87868;
  assign n87870 = ~n87852 & ~n87869;
  assign n87871 = ~n87848 & n87870;
  assign n87872 = n87843 & n87871;
  assign n87873 = pi2792 & n87872;
  assign n87874 = ~pi2792 & ~n87872;
  assign po2937 = n87873 | n87874;
  assign n87876 = ~n86951 & ~n86959;
  assign n87877 = n86901 & ~n87876;
  assign n87878 = ~n86964 & ~n87195;
  assign n87879 = ~n86927 & n87878;
  assign n87880 = ~n86934 & ~n87879;
  assign n87881 = n86901 & n87880;
  assign n87882 = ~n87877 & ~n87881;
  assign n87883 = n86950 & n87198;
  assign n87884 = ~n87200 & ~n87883;
  assign n87885 = ~n86967 & ~n87217;
  assign n87886 = n86934 & ~n87885;
  assign n87887 = n86901 & n87886;
  assign n87888 = n87884 & ~n87887;
  assign n87889 = n86907 & n86950;
  assign n87890 = n86907 & n86942;
  assign n87891 = ~n87190 & ~n87890;
  assign n87892 = n86934 & ~n87891;
  assign n87893 = ~n86965 & ~n87152;
  assign n87894 = n86907 & n86949;
  assign n87895 = ~n86989 & ~n87894;
  assign n87896 = ~n86934 & ~n87895;
  assign n87897 = n87893 & ~n87896;
  assign n87898 = ~n87892 & n87897;
  assign n87899 = ~n87889 & n87898;
  assign n87900 = ~n86901 & ~n87899;
  assign n87901 = n87153 & ~n87168;
  assign n87902 = n86934 & ~n87901;
  assign n87903 = ~n87900 & ~n87902;
  assign n87904 = n87888 & n87903;
  assign n87905 = n87882 & n87904;
  assign n87906 = ~pi2801 & ~n87905;
  assign n87907 = pi2801 & n87888;
  assign n87908 = n87882 & n87907;
  assign n87909 = n87903 & n87908;
  assign po2938 = n87906 | n87909;
  assign n87911 = ~n86771 & n87731;
  assign n87912 = n86771 & n86834;
  assign n87913 = ~n86819 & ~n87912;
  assign n87914 = n86765 & ~n87913;
  assign n87915 = ~n87911 & ~n87914;
  assign n87916 = ~n86765 & ~n86771;
  assign n87917 = ~n86783 & n87916;
  assign n87918 = n86777 & n87917;
  assign n87919 = n86808 & n86835;
  assign n87920 = ~n87918 & ~n87919;
  assign n87921 = ~n87720 & n87920;
  assign n87922 = ~n86801 & ~n86807;
  assign n87923 = ~n86849 & n87922;
  assign n87924 = n87921 & n87923;
  assign n87925 = n87915 & n87924;
  assign n87926 = ~n86832 & ~n87925;
  assign n87927 = ~n86800 & ~n86819;
  assign n87928 = n86771 & ~n87927;
  assign n87929 = ~n87725 & ~n87727;
  assign n87930 = ~n86783 & ~n86790;
  assign n87931 = n86771 & n87930;
  assign n87932 = n87929 & ~n87931;
  assign n87933 = n86765 & ~n87932;
  assign n87934 = ~n86771 & n86805;
  assign n87935 = n86771 & n86798;
  assign n87936 = ~n87934 & ~n87935;
  assign n87937 = ~n86765 & ~n87936;
  assign n87938 = ~n86771 & n86809;
  assign n87939 = ~n87937 & ~n87938;
  assign n87940 = ~n87933 & n87939;
  assign n87941 = ~n87928 & n87940;
  assign n87942 = n86832 & ~n87941;
  assign n87943 = n86765 & n86839;
  assign n87944 = ~n87942 & ~n87943;
  assign n87945 = ~n86765 & n87911;
  assign n87946 = n87944 & ~n87945;
  assign n87947 = ~n87926 & n87946;
  assign n87948 = ~pi2814 & ~n87947;
  assign n87949 = pi2814 & n87944;
  assign n87950 = ~n87926 & n87949;
  assign n87951 = ~n87945 & n87950;
  assign po2939 = n87948 | n87951;
  assign n87953 = ~n87240 & n87262;
  assign n87954 = ~n87292 & ~n87953;
  assign n87955 = ~n87234 & ~n87954;
  assign n87956 = n87253 & n87284;
  assign n87957 = ~n87838 & ~n87956;
  assign n87958 = n87234 & ~n87957;
  assign n87959 = ~n87253 & n87279;
  assign n87960 = ~n87858 & ~n87959;
  assign n87961 = ~n87261 & n87960;
  assign n87962 = ~n87958 & n87961;
  assign n87963 = ~n87955 & n87962;
  assign n87964 = ~n87833 & ~n87845;
  assign n87965 = n87963 & n87964;
  assign n87966 = n87271 & ~n87965;
  assign n87967 = n87247 & n87834;
  assign n87968 = n87301 & ~n87967;
  assign n87969 = n87234 & ~n87968;
  assign n87970 = ~n87253 & n87289;
  assign n87971 = ~n87969 & ~n87970;
  assign n87972 = ~n87246 & n87262;
  assign n87973 = n87253 & n87275;
  assign n87974 = ~n87972 & ~n87973;
  assign n87975 = n87234 & ~n87974;
  assign n87976 = n87234 & n87284;
  assign n87977 = ~n87253 & n87976;
  assign n87978 = ~n87975 & ~n87977;
  assign n87979 = n87971 & n87978;
  assign n87980 = ~n87271 & ~n87979;
  assign n87981 = ~n87279 & ~n87286;
  assign n87982 = ~n87839 & n87981;
  assign n87983 = n87306 & ~n87982;
  assign n87984 = ~n87980 & ~n87983;
  assign n87985 = ~n87261 & ~n87833;
  assign n87986 = ~n87234 & ~n87985;
  assign n87987 = n87984 & ~n87986;
  assign n87988 = ~n87966 & n87987;
  assign n87989 = ~pi2796 & n87988;
  assign n87990 = pi2796 & ~n87988;
  assign po2940 = n87989 | n87990;
  assign n87992 = ~n87499 & n87748;
  assign n87993 = ~n87549 & ~n87557;
  assign n87994 = n87499 & n87518;
  assign n87995 = ~n87499 & n87569;
  assign n87996 = ~n87994 & ~n87995;
  assign n87997 = n87993 & n87996;
  assign n87998 = n87528 & ~n87997;
  assign n87999 = n87499 & n87530;
  assign n88000 = ~n87529 & ~n87999;
  assign n88001 = ~n87551 & n88000;
  assign n88002 = ~n87528 & ~n88001;
  assign n88003 = n87499 & ~n87511;
  assign n88004 = n87517 & n88003;
  assign n88005 = n87505 & n88004;
  assign n88006 = ~n88002 & ~n88005;
  assign n88007 = ~n87998 & n88006;
  assign n88008 = ~n87992 & n88007;
  assign n88009 = ~n87493 & ~n88008;
  assign n88010 = n87499 & n87528;
  assign n88011 = n87535 & n88010;
  assign n88012 = n87528 & n87551;
  assign n88013 = n87528 & n87561;
  assign n88014 = ~n88012 & ~n88013;
  assign n88015 = ~n87499 & ~n88014;
  assign n88016 = ~n88011 & ~n88015;
  assign n88017 = ~n87499 & n87519;
  assign n88018 = ~n87760 & ~n88017;
  assign n88019 = n87499 & n87548;
  assign n88020 = ~n87499 & n87530;
  assign n88021 = ~n88019 & ~n88020;
  assign n88022 = ~n87519 & n88021;
  assign n88023 = ~n87549 & n88022;
  assign n88024 = ~n87528 & ~n88023;
  assign n88025 = ~n87499 & n87531;
  assign n88026 = ~n88024 & ~n88025;
  assign n88027 = n88018 & n88026;
  assign n88028 = n88016 & n88027;
  assign n88029 = n87493 & ~n88028;
  assign n88030 = n87528 & ~n87751;
  assign n88031 = ~n88029 & ~n88030;
  assign n88032 = ~n87552 & ~n88017;
  assign n88033 = ~n87528 & ~n88032;
  assign n88034 = n88031 & ~n88033;
  assign n88035 = ~n88009 & n88034;
  assign n88036 = pi2797 & ~n88035;
  assign n88037 = ~pi2797 & n88035;
  assign po2941 = n88036 | n88037;
  assign n88039 = pi6377 & pi9040;
  assign n88040 = pi6537 & ~pi9040;
  assign n88041 = ~n88039 & ~n88040;
  assign n88042 = ~pi2781 & ~n88041;
  assign n88043 = pi2781 & n88041;
  assign n88044 = ~n88042 & ~n88043;
  assign n88045 = pi6247 & pi9040;
  assign n88046 = pi6472 & ~pi9040;
  assign n88047 = ~n88045 & ~n88046;
  assign n88048 = pi2770 & n88047;
  assign n88049 = ~pi2770 & ~n88047;
  assign n88050 = ~n88048 & ~n88049;
  assign n88051 = pi6303 & pi9040;
  assign n88052 = pi6305 & ~pi9040;
  assign n88053 = ~n88051 & ~n88052;
  assign n88054 = ~pi2769 & n88053;
  assign n88055 = pi2769 & ~n88053;
  assign n88056 = ~n88054 & ~n88055;
  assign n88057 = ~n88050 & ~n88056;
  assign n88058 = n88044 & n88057;
  assign n88059 = pi6232 & ~pi9040;
  assign n88060 = pi6310 & pi9040;
  assign n88061 = ~n88059 & ~n88060;
  assign n88062 = ~pi2759 & n88061;
  assign n88063 = pi2759 & ~n88061;
  assign n88064 = ~n88062 & ~n88063;
  assign n88065 = n88044 & ~n88064;
  assign n88066 = ~n88056 & n88065;
  assign n88067 = ~n88044 & ~n88064;
  assign n88068 = n88056 & n88067;
  assign n88069 = ~n88066 & ~n88068;
  assign n88070 = ~n88058 & n88069;
  assign n88071 = pi6269 & pi9040;
  assign n88072 = pi6244 & ~pi9040;
  assign n88073 = ~n88071 & ~n88072;
  assign n88074 = ~pi2739 & ~n88073;
  assign n88075 = pi2739 & n88073;
  assign n88076 = ~n88074 & ~n88075;
  assign n88077 = pi6299 & ~pi9040;
  assign n88078 = pi6274 & pi9040;
  assign n88079 = ~n88077 & ~n88078;
  assign n88080 = ~pi2757 & ~n88079;
  assign n88081 = pi2757 & n88079;
  assign n88082 = ~n88080 & ~n88081;
  assign n88083 = ~n88076 & n88082;
  assign n88084 = ~n88070 & n88083;
  assign n88085 = ~n88044 & n88064;
  assign n88086 = ~n88056 & n88085;
  assign n88087 = n88050 & n88082;
  assign n88088 = n88086 & n88087;
  assign n88089 = ~n88056 & n88067;
  assign n88090 = n88076 & n88089;
  assign n88091 = n88044 & n88064;
  assign n88092 = n88050 & n88091;
  assign n88093 = n88044 & n88056;
  assign n88094 = ~n88092 & ~n88093;
  assign n88095 = n88076 & ~n88094;
  assign n88096 = ~n88090 & ~n88095;
  assign n88097 = n88082 & ~n88096;
  assign n88098 = ~n88088 & ~n88097;
  assign n88099 = n88050 & n88056;
  assign n88100 = n88044 & n88099;
  assign n88101 = ~n88050 & n88056;
  assign n88102 = ~n88044 & n88101;
  assign n88103 = n88064 & n88102;
  assign n88104 = ~n88100 & ~n88103;
  assign n88105 = n88076 & ~n88104;
  assign n88106 = n88098 & ~n88105;
  assign n88107 = n88050 & ~n88076;
  assign n88108 = n88091 & n88107;
  assign n88109 = ~n88056 & n88108;
  assign n88110 = ~n88065 & ~n88085;
  assign n88111 = n88057 & ~n88110;
  assign n88112 = ~n88064 & n88102;
  assign n88113 = ~n88111 & ~n88112;
  assign n88114 = n88099 & ~n88110;
  assign n88115 = n88050 & ~n88056;
  assign n88116 = ~n88044 & n88115;
  assign n88117 = ~n88064 & n88116;
  assign n88118 = ~n88114 & ~n88117;
  assign n88119 = n88056 & n88091;
  assign n88120 = ~n88050 & ~n88076;
  assign n88121 = n88119 & n88120;
  assign n88122 = n88118 & ~n88121;
  assign n88123 = n88113 & n88122;
  assign n88124 = ~n88109 & n88123;
  assign n88125 = ~n88050 & n88076;
  assign n88126 = ~n88056 & n88125;
  assign n88127 = n88064 & n88126;
  assign n88128 = n88124 & ~n88127;
  assign n88129 = ~n88082 & ~n88128;
  assign n88130 = n88106 & ~n88129;
  assign n88131 = ~n88084 & n88130;
  assign n88132 = ~pi2809 & ~n88131;
  assign n88133 = pi2809 & n88106;
  assign n88134 = ~n88084 & n88133;
  assign n88135 = ~n88129 & n88134;
  assign po2942 = n88132 | n88135;
  assign n88137 = n87371 & n87402;
  assign n88138 = ~n87401 & n88137;
  assign n88139 = ~n87816 & ~n88138;
  assign n88140 = ~n87383 & n87401;
  assign n88141 = n87377 & n88140;
  assign n88142 = ~n87389 & ~n87401;
  assign n88143 = ~n87431 & ~n88142;
  assign n88144 = ~n87371 & ~n88143;
  assign n88145 = ~n88141 & ~n88144;
  assign n88146 = n88139 & n88145;
  assign n88147 = n87365 & ~n88146;
  assign n88148 = ~n87422 & ~n87622;
  assign n88149 = n87390 & ~n87401;
  assign n88150 = n88148 & ~n88149;
  assign n88151 = n87371 & ~n88150;
  assign n88152 = n87402 & n87620;
  assign n88153 = ~n87610 & ~n88152;
  assign n88154 = ~n88151 & n88153;
  assign n88155 = ~n87409 & ~n87603;
  assign n88156 = ~n87371 & ~n88155;
  assign n88157 = n88154 & ~n88156;
  assign n88158 = ~n87365 & ~n88157;
  assign n88159 = ~n88147 & ~n88158;
  assign n88160 = n87392 & ~n87401;
  assign n88161 = n87401 & ~n87599;
  assign n88162 = ~n88160 & ~n88161;
  assign n88163 = ~n87371 & ~n88162;
  assign n88164 = n87394 & ~n87422;
  assign n88165 = n87805 & ~n88164;
  assign n88166 = ~n88163 & ~n88165;
  assign n88167 = n88159 & n88166;
  assign n88168 = ~pi2800 & ~n88167;
  assign n88169 = pi2800 & n88166;
  assign n88170 = ~n88158 & n88169;
  assign n88171 = ~n88147 & n88170;
  assign po2943 = n88168 | n88171;
  assign n88173 = ~n86850 & ~n87938;
  assign n88174 = n86765 & ~n88173;
  assign n88175 = ~n86832 & n86834;
  assign n88176 = ~n86765 & n88175;
  assign n88177 = ~n86777 & n87712;
  assign n88178 = ~n87930 & ~n88177;
  assign n88179 = ~n86809 & n88178;
  assign n88180 = n86765 & ~n88179;
  assign n88181 = ~n86771 & n86806;
  assign n88182 = ~n88180 & ~n88181;
  assign n88183 = ~n86832 & ~n88182;
  assign n88184 = ~n88176 & ~n88183;
  assign n88185 = ~n86792 & ~n86801;
  assign n88186 = ~n86771 & n87727;
  assign n88187 = ~n87912 & ~n88186;
  assign n88188 = n88185 & n88187;
  assign n88189 = ~n86765 & ~n88188;
  assign n88190 = n86777 & n86790;
  assign n88191 = ~n86765 & n88190;
  assign n88192 = n86771 & n88191;
  assign n88193 = ~n86771 & n87930;
  assign n88194 = ~n86792 & ~n88193;
  assign n88195 = ~n87935 & n88194;
  assign n88196 = ~n88192 & n88195;
  assign n88197 = n86765 & n86800;
  assign n88198 = n88196 & ~n88197;
  assign n88199 = n86832 & ~n88198;
  assign n88200 = ~n88189 & ~n88199;
  assign n88201 = n88184 & n88200;
  assign n88202 = ~n88174 & n88201;
  assign n88203 = pi2843 & n88202;
  assign n88204 = ~pi2843 & ~n88202;
  assign po2944 = n88203 | n88204;
  assign n88206 = ~n87253 & n87275;
  assign n88207 = ~n87274 & ~n88206;
  assign n88208 = ~n87234 & ~n88207;
  assign n88209 = n87234 & ~n87860;
  assign n88210 = ~n87849 & ~n88209;
  assign n88211 = ~n88208 & n88210;
  assign n88212 = n87271 & ~n88211;
  assign n88213 = ~n87234 & n87289;
  assign n88214 = ~n88212 & ~n88213;
  assign n88215 = ~n87959 & ~n87973;
  assign n88216 = n87234 & ~n88215;
  assign n88217 = n87234 & n87276;
  assign n88218 = n87240 & n87262;
  assign n88219 = ~n87246 & n88218;
  assign n88220 = ~n87234 & n87260;
  assign n88221 = ~n87837 & ~n88220;
  assign n88222 = n87246 & ~n88221;
  assign n88223 = ~n87838 & ~n88222;
  assign n88224 = ~n87261 & n88223;
  assign n88225 = ~n88219 & n88224;
  assign n88226 = ~n88217 & n88225;
  assign n88227 = ~n87271 & ~n88226;
  assign n88228 = ~n88216 & ~n88227;
  assign n88229 = n88214 & n88228;
  assign n88230 = pi2810 & ~n88229;
  assign n88231 = ~pi2810 & n88229;
  assign po2945 = n88230 | n88231;
  assign n88233 = ~n88056 & n88091;
  assign n88234 = n88076 & n88233;
  assign n88235 = ~n88050 & n88234;
  assign n88236 = n88076 & n88112;
  assign n88237 = ~n88235 & ~n88236;
  assign n88238 = ~n88112 & ~n88121;
  assign n88239 = ~n88056 & ~n88064;
  assign n88240 = n88050 & n88239;
  assign n88241 = ~n88092 & ~n88240;
  assign n88242 = n88076 & ~n88241;
  assign n88243 = ~n88076 & ~n88101;
  assign n88244 = ~n88110 & n88243;
  assign n88245 = ~n88050 & ~n88091;
  assign n88246 = n88076 & n88245;
  assign n88247 = n88056 & n88246;
  assign n88248 = ~n88244 & ~n88247;
  assign n88249 = ~n88242 & n88248;
  assign n88250 = n88238 & n88249;
  assign n88251 = n88082 & ~n88250;
  assign n88252 = n88237 & ~n88251;
  assign n88253 = n88066 & ~n88076;
  assign n88254 = n88050 & n88253;
  assign n88255 = ~n88076 & ~n88082;
  assign n88256 = ~n88089 & ~n88092;
  assign n88257 = n88101 & ~n88110;
  assign n88258 = n88256 & ~n88257;
  assign n88259 = n88255 & ~n88258;
  assign n88260 = n88050 & n88068;
  assign n88261 = n88050 & ~n88064;
  assign n88262 = n88056 & n88261;
  assign n88263 = n88050 & n88085;
  assign n88264 = ~n88262 & ~n88263;
  assign n88265 = ~n88050 & n88091;
  assign n88266 = ~n88086 & ~n88265;
  assign n88267 = n88264 & n88266;
  assign n88268 = n88076 & ~n88267;
  assign n88269 = ~n88260 & ~n88268;
  assign n88270 = ~n88082 & ~n88269;
  assign n88271 = ~n88259 & ~n88270;
  assign n88272 = ~n88254 & n88271;
  assign n88273 = n88252 & n88272;
  assign n88274 = pi2805 & ~n88273;
  assign n88275 = ~pi2805 & n88252;
  assign n88276 = n88272 & n88275;
  assign po2946 = n88274 | n88276;
  assign n88278 = n88056 & n88065;
  assign n88279 = ~n88233 & ~n88278;
  assign n88280 = n88076 & ~n88279;
  assign n88281 = ~n88050 & n88085;
  assign n88282 = ~n88066 & ~n88281;
  assign n88283 = ~n88119 & n88282;
  assign n88284 = ~n88076 & ~n88283;
  assign n88285 = ~n88280 & ~n88284;
  assign n88286 = ~n88090 & ~n88103;
  assign n88287 = n88285 & n88286;
  assign n88288 = ~n88082 & ~n88287;
  assign n88289 = n88050 & n88233;
  assign n88290 = ~n88050 & n88067;
  assign n88291 = ~n88263 & ~n88290;
  assign n88292 = ~n88076 & ~n88291;
  assign n88293 = ~n88289 & ~n88292;
  assign n88294 = n88076 & n88086;
  assign n88295 = n88069 & ~n88294;
  assign n88296 = ~n88119 & n88295;
  assign n88297 = ~n88050 & ~n88296;
  assign n88298 = n88293 & ~n88297;
  assign n88299 = n88082 & ~n88298;
  assign n88300 = ~n88288 & ~n88299;
  assign n88301 = n88056 & n88263;
  assign n88302 = ~n88117 & ~n88301;
  assign n88303 = n88076 & ~n88302;
  assign n88304 = n88056 & ~n88064;
  assign n88305 = ~n88076 & n88304;
  assign n88306 = n88050 & n88305;
  assign n88307 = ~n88303 & ~n88306;
  assign n88308 = n88300 & n88307;
  assign n88309 = ~pi2816 & ~n88308;
  assign n88310 = pi2816 & ~n88303;
  assign n88311 = n88300 & n88310;
  assign n88312 = ~n88306 & n88311;
  assign po2947 = n88309 | n88312;
  assign n88314 = ~n88263 & ~n88265;
  assign n88315 = n88076 & ~n88314;
  assign n88316 = ~n88236 & ~n88315;
  assign n88317 = n88082 & ~n88316;
  assign n88318 = ~n88065 & ~n88304;
  assign n88319 = ~n88050 & ~n88318;
  assign n88320 = ~n88233 & ~n88319;
  assign n88321 = ~n88076 & ~n88320;
  assign n88322 = ~n88257 & ~n88321;
  assign n88323 = n88050 & n88119;
  assign n88324 = ~n88044 & n88057;
  assign n88325 = n88050 & ~n88318;
  assign n88326 = ~n88324 & ~n88325;
  assign n88327 = n88076 & ~n88326;
  assign n88328 = ~n88323 & ~n88327;
  assign n88329 = n88322 & n88328;
  assign n88330 = ~n88082 & ~n88329;
  assign n88331 = ~n88065 & n88115;
  assign n88332 = n88082 & n88331;
  assign n88333 = n88065 & n88099;
  assign n88334 = n88076 & n88333;
  assign n88335 = ~n88056 & n88107;
  assign n88336 = ~n88044 & n88335;
  assign n88337 = ~n88334 & ~n88336;
  assign n88338 = ~n88332 & n88337;
  assign n88339 = ~n88086 & ~n88261;
  assign n88340 = n88083 & ~n88339;
  assign n88341 = n88338 & ~n88340;
  assign n88342 = ~n88330 & n88341;
  assign n88343 = ~n88317 & n88342;
  assign n88344 = pi2811 & ~n88343;
  assign n88345 = ~pi2811 & n88343;
  assign po2948 = n88344 | n88345;
  assign n88347 = ~n87754 & ~n88017;
  assign n88348 = ~n88005 & n88347;
  assign n88349 = n87528 & ~n88348;
  assign n88350 = ~n87763 & ~n87779;
  assign n88351 = ~n87760 & ~n88013;
  assign n88352 = ~n87748 & ~n88020;
  assign n88353 = ~n87528 & ~n88352;
  assign n88354 = ~n87557 & ~n88353;
  assign n88355 = n88351 & n88354;
  assign n88356 = n87493 & ~n88355;
  assign n88357 = ~n87511 & n87517;
  assign n88358 = ~n87541 & ~n88357;
  assign n88359 = n87499 & ~n88358;
  assign n88360 = ~n87519 & ~n87766;
  assign n88361 = ~n87528 & ~n88360;
  assign n88362 = n87499 & n87517;
  assign n88363 = ~n87531 & ~n88362;
  assign n88364 = ~n87538 & n88363;
  assign n88365 = n87528 & ~n88364;
  assign n88366 = ~n88361 & ~n88365;
  assign n88367 = ~n88359 & n88366;
  assign n88368 = ~n87493 & ~n88367;
  assign n88369 = ~n88356 & ~n88368;
  assign n88370 = n88350 & n88369;
  assign n88371 = ~n88349 & n88370;
  assign n88372 = ~pi2808 & ~n88371;
  assign n88373 = pi2808 & n88350;
  assign n88374 = ~n88349 & n88373;
  assign n88375 = n88369 & n88374;
  assign po2949 = n88372 | n88375;
  assign n88377 = pi6485 & ~pi9040;
  assign n88378 = pi6599 & pi9040;
  assign n88379 = ~n88377 & ~n88378;
  assign n88380 = ~pi2802 & n88379;
  assign n88381 = pi2802 & ~n88379;
  assign n88382 = ~n88380 & ~n88381;
  assign n88383 = pi6491 & ~pi9040;
  assign n88384 = pi6637 & pi9040;
  assign n88385 = ~n88383 & ~n88384;
  assign n88386 = ~pi2844 & ~n88385;
  assign n88387 = pi2844 & n88385;
  assign n88388 = ~n88386 & ~n88387;
  assign n88389 = pi6610 & ~pi9040;
  assign n88390 = pi6416 & pi9040;
  assign n88391 = ~n88389 & ~n88390;
  assign n88392 = pi2820 & n88391;
  assign n88393 = ~pi2820 & ~n88391;
  assign n88394 = ~n88392 & ~n88393;
  assign n88395 = pi6598 & pi9040;
  assign n88396 = pi6637 & ~pi9040;
  assign n88397 = ~n88395 & ~n88396;
  assign n88398 = ~pi2835 & ~n88397;
  assign n88399 = pi2835 & n88397;
  assign n88400 = ~n88398 & ~n88399;
  assign n88401 = ~n88394 & n88400;
  assign n88402 = n88388 & n88401;
  assign n88403 = ~n88382 & n88402;
  assign n88404 = pi6494 & ~pi9040;
  assign n88405 = pi6404 & pi9040;
  assign n88406 = ~n88404 & ~n88405;
  assign n88407 = ~pi2818 & ~n88406;
  assign n88408 = pi2818 & n88406;
  assign n88409 = ~n88407 & ~n88408;
  assign n88410 = ~n88388 & ~n88394;
  assign n88411 = n88382 & n88410;
  assign n88412 = n88409 & n88411;
  assign n88413 = ~n88403 & ~n88412;
  assign n88414 = pi6614 & ~pi9040;
  assign n88415 = pi6459 & pi9040;
  assign n88416 = ~n88414 & ~n88415;
  assign n88417 = ~pi2839 & ~n88416;
  assign n88418 = pi2839 & n88416;
  assign n88419 = ~n88417 & ~n88418;
  assign n88420 = ~n88400 & ~n88419;
  assign n88421 = ~n88382 & n88409;
  assign n88422 = ~n88394 & n88421;
  assign n88423 = n88382 & n88409;
  assign n88424 = n88388 & n88423;
  assign n88425 = n88394 & n88424;
  assign n88426 = ~n88422 & ~n88425;
  assign n88427 = n88388 & ~n88409;
  assign n88428 = ~n88394 & n88427;
  assign n88429 = n88426 & ~n88428;
  assign n88430 = n88420 & ~n88429;
  assign n88431 = ~n88388 & n88423;
  assign n88432 = n88388 & n88421;
  assign n88433 = ~n88431 & ~n88432;
  assign n88434 = n88382 & n88427;
  assign n88435 = n88394 & n88434;
  assign n88436 = ~n88411 & ~n88435;
  assign n88437 = n88433 & n88436;
  assign n88438 = n88400 & ~n88437;
  assign n88439 = ~n88382 & ~n88409;
  assign n88440 = ~n88388 & n88439;
  assign n88441 = n88394 & n88440;
  assign n88442 = ~n88438 & ~n88441;
  assign n88443 = ~n88419 & ~n88442;
  assign n88444 = ~n88430 & ~n88443;
  assign n88445 = n88382 & ~n88409;
  assign n88446 = ~n88388 & n88445;
  assign n88447 = ~n88421 & ~n88445;
  assign n88448 = n88394 & ~n88447;
  assign n88449 = ~n88446 & ~n88448;
  assign n88450 = ~n88400 & ~n88449;
  assign n88451 = n88388 & n88439;
  assign n88452 = ~n88428 & ~n88451;
  assign n88453 = ~n88425 & n88452;
  assign n88454 = n88400 & ~n88453;
  assign n88455 = ~n88450 & ~n88454;
  assign n88456 = ~n88394 & ~n88400;
  assign n88457 = n88423 & n88456;
  assign n88458 = n88394 & n88446;
  assign n88459 = ~n88388 & n88409;
  assign n88460 = ~n88382 & n88459;
  assign n88461 = n88394 & n88460;
  assign n88462 = ~n88458 & ~n88461;
  assign n88463 = ~n88382 & n88410;
  assign n88464 = ~n88409 & n88463;
  assign n88465 = n88462 & ~n88464;
  assign n88466 = ~n88457 & n88465;
  assign n88467 = n88455 & n88466;
  assign n88468 = n88419 & ~n88467;
  assign n88469 = n88444 & ~n88468;
  assign n88470 = n88413 & n88469;
  assign n88471 = pi2861 & ~n88470;
  assign n88472 = ~pi2861 & n88413;
  assign n88473 = n88444 & n88472;
  assign n88474 = ~n88468 & n88473;
  assign po2968 = n88471 | n88474;
  assign n88476 = n88394 & n88427;
  assign n88477 = ~n88432 & ~n88476;
  assign n88478 = ~n88412 & n88477;
  assign n88479 = n88400 & ~n88478;
  assign n88480 = ~n88394 & n88460;
  assign n88481 = ~n88394 & n88451;
  assign n88482 = ~n88388 & ~n88409;
  assign n88483 = ~n88423 & ~n88482;
  assign n88484 = n88394 & ~n88483;
  assign n88485 = ~n88481 & ~n88484;
  assign n88486 = ~n88480 & n88485;
  assign n88487 = ~n88400 & ~n88486;
  assign n88488 = ~n88479 & ~n88487;
  assign n88489 = n88419 & ~n88488;
  assign n88490 = ~n88400 & n88446;
  assign n88491 = ~n88394 & n88490;
  assign n88492 = ~n88394 & n88424;
  assign n88493 = ~n88400 & n88492;
  assign n88494 = ~n88491 & ~n88493;
  assign n88495 = n88400 & n88464;
  assign n88496 = n88494 & ~n88495;
  assign n88497 = n88401 & ~n88409;
  assign n88498 = ~n88394 & n88409;
  assign n88499 = n88388 & n88498;
  assign n88500 = ~n88476 & ~n88499;
  assign n88501 = ~n88400 & ~n88500;
  assign n88502 = ~n88457 & ~n88501;
  assign n88503 = ~n88461 & ~n88492;
  assign n88504 = n88394 & n88400;
  assign n88505 = n88459 & n88504;
  assign n88506 = n88400 & n88440;
  assign n88507 = ~n88505 & ~n88506;
  assign n88508 = n88503 & n88507;
  assign n88509 = n88502 & n88508;
  assign n88510 = ~n88497 & n88509;
  assign n88511 = ~n88419 & ~n88510;
  assign n88512 = ~n88394 & n88434;
  assign n88513 = n88394 & n88421;
  assign n88514 = ~n88512 & ~n88513;
  assign n88515 = n88400 & ~n88514;
  assign n88516 = ~n88511 & ~n88515;
  assign n88517 = n88496 & n88516;
  assign n88518 = ~n88489 & n88517;
  assign n88519 = ~pi2857 & ~n88518;
  assign n88520 = pi2857 & n88518;
  assign po2969 = n88519 | n88520;
  assign n88522 = pi6627 & pi9040;
  assign n88523 = pi6619 & ~pi9040;
  assign n88524 = ~n88522 & ~n88523;
  assign n88525 = ~pi2821 & ~n88524;
  assign n88526 = pi2821 & n88524;
  assign n88527 = ~n88525 & ~n88526;
  assign n88528 = pi6500 & ~pi9040;
  assign n88529 = pi6481 & pi9040;
  assign n88530 = ~n88528 & ~n88529;
  assign n88531 = ~pi2827 & ~n88530;
  assign n88532 = pi2827 & n88530;
  assign n88533 = ~n88531 & ~n88532;
  assign n88534 = pi6468 & ~pi9040;
  assign n88535 = pi6555 & pi9040;
  assign n88536 = ~n88534 & ~n88535;
  assign n88537 = ~pi2830 & n88536;
  assign n88538 = pi2830 & ~n88536;
  assign n88539 = ~n88537 & ~n88538;
  assign n88540 = pi6604 & ~pi9040;
  assign n88541 = pi6610 & pi9040;
  assign n88542 = ~n88540 & ~n88541;
  assign n88543 = ~pi2813 & ~n88542;
  assign n88544 = pi2813 & n88542;
  assign n88545 = ~n88543 & ~n88544;
  assign n88546 = ~n88539 & n88545;
  assign n88547 = ~n88533 & n88546;
  assign n88548 = pi6598 & ~pi9040;
  assign n88549 = pi6577 & pi9040;
  assign n88550 = ~n88548 & ~n88549;
  assign n88551 = pi2842 & n88550;
  assign n88552 = ~pi2842 & ~n88550;
  assign n88553 = ~n88551 & ~n88552;
  assign n88554 = n88547 & ~n88553;
  assign n88555 = n88539 & ~n88545;
  assign n88556 = ~n88533 & n88555;
  assign n88557 = ~n88553 & n88556;
  assign n88558 = ~n88554 & ~n88557;
  assign n88559 = n88533 & n88555;
  assign n88560 = n88553 & n88559;
  assign n88561 = ~n88539 & ~n88545;
  assign n88562 = ~n88533 & n88561;
  assign n88563 = n88553 & n88562;
  assign n88564 = ~n88560 & ~n88563;
  assign n88565 = n88558 & n88564;
  assign n88566 = n88527 & ~n88565;
  assign n88567 = ~n88533 & n88553;
  assign n88568 = n88545 & n88567;
  assign n88569 = n88539 & n88568;
  assign n88570 = ~n88562 & ~n88569;
  assign n88571 = n88527 & ~n88570;
  assign n88572 = ~n88527 & n88545;
  assign n88573 = ~n88553 & n88572;
  assign n88574 = n88533 & ~n88539;
  assign n88575 = n88553 & n88555;
  assign n88576 = ~n88574 & ~n88575;
  assign n88577 = ~n88527 & ~n88576;
  assign n88578 = ~n88573 & ~n88577;
  assign n88579 = n88539 & n88545;
  assign n88580 = n88533 & n88579;
  assign n88581 = ~n88553 & n88580;
  assign n88582 = n88578 & ~n88581;
  assign n88583 = n88545 & n88574;
  assign n88584 = n88553 & n88583;
  assign n88585 = n88582 & ~n88584;
  assign n88586 = ~n88571 & n88585;
  assign n88587 = pi6419 & pi9040;
  assign n88588 = pi6542 & ~pi9040;
  assign n88589 = ~n88587 & ~n88588;
  assign n88590 = ~pi2846 & ~n88589;
  assign n88591 = pi2846 & n88589;
  assign n88592 = ~n88590 & ~n88591;
  assign n88593 = ~n88586 & ~n88592;
  assign n88594 = ~n88533 & n88545;
  assign n88595 = ~n88527 & n88553;
  assign n88596 = n88592 & n88595;
  assign n88597 = n88594 & n88596;
  assign n88598 = ~n88533 & ~n88553;
  assign n88599 = ~n88545 & n88598;
  assign n88600 = ~n88527 & ~n88599;
  assign n88601 = n88533 & n88553;
  assign n88602 = n88539 & n88601;
  assign n88603 = ~n88546 & ~n88594;
  assign n88604 = ~n88553 & ~n88603;
  assign n88605 = n88527 & ~n88559;
  assign n88606 = ~n88604 & n88605;
  assign n88607 = ~n88602 & n88606;
  assign n88608 = ~n88600 & ~n88607;
  assign n88609 = n88533 & n88561;
  assign n88610 = n88553 & n88609;
  assign n88611 = ~n88608 & ~n88610;
  assign n88612 = n88592 & ~n88611;
  assign n88613 = ~n88597 & ~n88612;
  assign n88614 = ~n88593 & n88613;
  assign n88615 = ~n88566 & n88614;
  assign n88616 = ~n88527 & n88581;
  assign n88617 = n88615 & ~n88616;
  assign n88618 = pi2852 & ~n88617;
  assign n88619 = n88614 & ~n88616;
  assign n88620 = ~pi2852 & n88619;
  assign n88621 = ~n88566 & n88620;
  assign po2971 = n88618 | n88621;
  assign n88623 = ~n88446 & ~n88451;
  assign n88624 = ~n88400 & ~n88623;
  assign n88625 = n88394 & n88432;
  assign n88626 = ~n88624 & ~n88625;
  assign n88627 = n88394 & n88409;
  assign n88628 = ~n88459 & ~n88627;
  assign n88629 = ~n88434 & n88628;
  assign n88630 = n88400 & ~n88629;
  assign n88631 = n88626 & ~n88630;
  assign n88632 = ~n88419 & ~n88631;
  assign n88633 = ~n88400 & n88480;
  assign n88634 = ~n88493 & ~n88633;
  assign n88635 = ~n88495 & n88634;
  assign n88636 = n88388 & ~n88394;
  assign n88637 = n88382 & n88636;
  assign n88638 = ~n88464 & ~n88637;
  assign n88639 = n88400 & n88499;
  assign n88640 = n88394 & n88451;
  assign n88641 = ~n88400 & n88459;
  assign n88642 = ~n88640 & ~n88641;
  assign n88643 = ~n88458 & n88642;
  assign n88644 = ~n88639 & n88643;
  assign n88645 = n88638 & n88644;
  assign n88646 = ~n88506 & n88645;
  assign n88647 = n88419 & ~n88646;
  assign n88648 = n88635 & ~n88647;
  assign n88649 = ~n88632 & n88648;
  assign n88650 = ~pi2870 & ~n88649;
  assign n88651 = pi2870 & n88635;
  assign n88652 = ~n88632 & n88651;
  assign n88653 = ~n88647 & n88652;
  assign po2978 = n88650 | n88653;
  assign n88655 = n88400 & n88421;
  assign n88656 = ~n88394 & n88655;
  assign n88657 = ~n88512 & ~n88656;
  assign n88658 = ~n88382 & n88394;
  assign n88659 = n88388 & n88658;
  assign n88660 = ~n88394 & ~n88409;
  assign n88661 = ~n88637 & ~n88660;
  assign n88662 = ~n88400 & ~n88661;
  assign n88663 = ~n88659 & ~n88662;
  assign n88664 = n88657 & n88663;
  assign n88665 = n88419 & ~n88664;
  assign n88666 = ~n88424 & ~n88461;
  assign n88667 = ~n88394 & n88439;
  assign n88668 = n88666 & ~n88667;
  assign n88669 = n88400 & ~n88668;
  assign n88670 = n88421 & n88456;
  assign n88671 = ~n88412 & ~n88670;
  assign n88672 = ~n88669 & n88671;
  assign n88673 = ~n88434 & ~n88441;
  assign n88674 = ~n88400 & ~n88673;
  assign n88675 = n88672 & ~n88674;
  assign n88676 = ~n88419 & ~n88675;
  assign n88677 = ~n88665 & ~n88676;
  assign n88678 = ~n88394 & n88445;
  assign n88679 = n88394 & ~n88433;
  assign n88680 = ~n88678 & ~n88679;
  assign n88681 = ~n88400 & ~n88680;
  assign n88682 = ~n88424 & n88623;
  assign n88683 = n88504 & ~n88682;
  assign n88684 = ~n88681 & ~n88683;
  assign n88685 = n88677 & n88684;
  assign n88686 = ~pi2869 & ~n88685;
  assign n88687 = ~n88676 & n88684;
  assign n88688 = pi2869 & n88687;
  assign n88689 = ~n88665 & n88688;
  assign po2983 = n88686 | n88689;
  assign n88691 = pi6465 & pi9040;
  assign n88692 = pi6481 & ~pi9040;
  assign n88693 = ~n88691 & ~n88692;
  assign n88694 = pi2818 & n88693;
  assign n88695 = ~pi2818 & ~n88693;
  assign n88696 = ~n88694 & ~n88695;
  assign n88697 = pi6484 & ~pi9040;
  assign n88698 = pi6619 & pi9040;
  assign n88699 = ~n88697 & ~n88698;
  assign n88700 = pi2841 & n88699;
  assign n88701 = ~pi2841 & ~n88699;
  assign n88702 = ~n88700 & ~n88701;
  assign n88703 = pi6604 & pi9040;
  assign n88704 = pi6627 & ~pi9040;
  assign n88705 = ~n88703 & ~n88704;
  assign n88706 = ~pi2845 & n88705;
  assign n88707 = pi2845 & ~n88705;
  assign n88708 = ~n88706 & ~n88707;
  assign n88709 = pi6465 & ~pi9040;
  assign n88710 = pi6542 & pi9040;
  assign n88711 = ~n88709 & ~n88710;
  assign n88712 = ~pi2826 & ~n88711;
  assign n88713 = pi2826 & n88711;
  assign n88714 = ~n88712 & ~n88713;
  assign n88715 = pi6468 & pi9040;
  assign n88716 = pi6577 & ~pi9040;
  assign n88717 = ~n88715 & ~n88716;
  assign n88718 = ~pi2844 & ~n88717;
  assign n88719 = pi2844 & n88717;
  assign n88720 = ~n88718 & ~n88719;
  assign n88721 = n88714 & ~n88720;
  assign n88722 = ~n88708 & n88721;
  assign n88723 = n88702 & n88722;
  assign n88724 = pi6500 & pi9040;
  assign n88725 = pi6555 & ~pi9040;
  assign n88726 = ~n88724 & ~n88725;
  assign n88727 = pi2828 & n88726;
  assign n88728 = ~pi2828 & ~n88726;
  assign n88729 = ~n88727 & ~n88728;
  assign n88730 = ~n88708 & n88720;
  assign n88731 = n88714 & n88730;
  assign n88732 = n88708 & ~n88714;
  assign n88733 = ~n88714 & ~n88720;
  assign n88734 = ~n88702 & n88733;
  assign n88735 = n88708 & ~n88720;
  assign n88736 = n88702 & n88735;
  assign n88737 = ~n88734 & ~n88736;
  assign n88738 = ~n88732 & n88737;
  assign n88739 = ~n88731 & n88738;
  assign n88740 = n88729 & ~n88739;
  assign n88741 = ~n88702 & n88714;
  assign n88742 = n88720 & n88741;
  assign n88743 = n88708 & n88741;
  assign n88744 = ~n88714 & n88730;
  assign n88745 = ~n88743 & ~n88744;
  assign n88746 = ~n88729 & ~n88745;
  assign n88747 = ~n88742 & ~n88746;
  assign n88748 = ~n88740 & n88747;
  assign n88749 = ~n88723 & n88748;
  assign n88750 = n88696 & ~n88749;
  assign n88751 = n88708 & n88720;
  assign n88752 = ~n88714 & n88751;
  assign n88753 = ~n88702 & n88752;
  assign n88754 = ~n88714 & n88735;
  assign n88755 = n88702 & n88754;
  assign n88756 = ~n88723 & ~n88755;
  assign n88757 = ~n88753 & n88756;
  assign n88758 = n88729 & ~n88757;
  assign n88759 = ~n88750 & ~n88758;
  assign n88760 = ~n88708 & n88742;
  assign n88761 = ~n88708 & ~n88714;
  assign n88762 = ~n88729 & n88761;
  assign n88763 = n88702 & n88762;
  assign n88764 = ~n88702 & n88729;
  assign n88765 = n88714 & n88764;
  assign n88766 = ~n88720 & n88765;
  assign n88767 = n88714 & n88751;
  assign n88768 = n88702 & n88767;
  assign n88769 = ~n88766 & ~n88768;
  assign n88770 = n88708 & n88714;
  assign n88771 = n88702 & n88770;
  assign n88772 = ~n88708 & ~n88720;
  assign n88773 = ~n88714 & n88772;
  assign n88774 = ~n88771 & ~n88773;
  assign n88775 = ~n88729 & ~n88774;
  assign n88776 = ~n88729 & n88732;
  assign n88777 = ~n88702 & n88776;
  assign n88778 = ~n88775 & ~n88777;
  assign n88779 = n88769 & n88778;
  assign n88780 = ~n88696 & ~n88779;
  assign n88781 = ~n88763 & ~n88780;
  assign n88782 = ~n88760 & n88781;
  assign n88783 = n88759 & n88782;
  assign n88784 = ~pi2851 & ~n88783;
  assign n88785 = ~n88750 & ~n88760;
  assign n88786 = ~n88758 & n88785;
  assign n88787 = n88781 & n88786;
  assign n88788 = pi2851 & n88787;
  assign po2984 = n88784 | n88788;
  assign n88790 = pi6613 & pi9040;
  assign n88791 = pi6419 & ~pi9040;
  assign n88792 = ~n88790 & ~n88791;
  assign n88793 = ~pi2813 & ~n88792;
  assign n88794 = pi2813 & n88792;
  assign n88795 = ~n88793 & ~n88794;
  assign n88796 = pi6541 & ~pi9040;
  assign n88797 = pi6480 & pi9040;
  assign n88798 = ~n88796 & ~n88797;
  assign n88799 = ~pi2839 & ~n88798;
  assign n88800 = pi2839 & n88798;
  assign n88801 = ~n88799 & ~n88800;
  assign n88802 = pi6494 & pi9040;
  assign n88803 = pi6599 & ~pi9040;
  assign n88804 = ~n88802 & ~n88803;
  assign n88805 = ~pi2827 & ~n88804;
  assign n88806 = pi2827 & n88804;
  assign n88807 = ~n88805 & ~n88806;
  assign n88808 = ~n88801 & n88807;
  assign n88809 = pi6541 & pi9040;
  assign n88810 = pi6613 & ~pi9040;
  assign n88811 = ~n88809 & ~n88810;
  assign n88812 = ~pi2817 & ~n88811;
  assign n88813 = pi2817 & n88811;
  assign n88814 = ~n88812 & ~n88813;
  assign n88815 = pi6614 & pi9040;
  assign n88816 = pi6416 & ~pi9040;
  assign n88817 = ~n88815 & ~n88816;
  assign n88818 = pi2840 & n88817;
  assign n88819 = ~pi2840 & ~n88817;
  assign n88820 = ~n88818 & ~n88819;
  assign n88821 = ~n88814 & ~n88820;
  assign n88822 = n88808 & n88821;
  assign n88823 = pi6408 & pi9040;
  assign n88824 = pi6480 & ~pi9040;
  assign n88825 = ~n88823 & ~n88824;
  assign n88826 = ~pi2802 & n88825;
  assign n88827 = pi2802 & ~n88825;
  assign n88828 = ~n88826 & ~n88827;
  assign n88829 = n88801 & ~n88807;
  assign n88830 = ~n88828 & n88829;
  assign n88831 = n88814 & n88828;
  assign n88832 = ~n88807 & n88831;
  assign n88833 = ~n88801 & n88832;
  assign n88834 = ~n88830 & ~n88833;
  assign n88835 = n88801 & n88807;
  assign n88836 = n88814 & n88835;
  assign n88837 = n88834 & ~n88836;
  assign n88838 = ~n88820 & ~n88837;
  assign n88839 = n88801 & n88828;
  assign n88840 = ~n88814 & n88820;
  assign n88841 = n88839 & n88840;
  assign n88842 = n88828 & n88829;
  assign n88843 = ~n88814 & n88842;
  assign n88844 = ~n88841 & ~n88843;
  assign n88845 = ~n88838 & n88844;
  assign n88846 = ~n88822 & n88845;
  assign n88847 = n88808 & ~n88828;
  assign n88848 = ~n88814 & n88847;
  assign n88849 = ~n88828 & n88835;
  assign n88850 = n88814 & n88849;
  assign n88851 = ~n88848 & ~n88850;
  assign n88852 = n88846 & n88851;
  assign n88853 = ~n88795 & ~n88852;
  assign n88854 = ~n88814 & n88828;
  assign n88855 = n88807 & n88854;
  assign n88856 = n88801 & n88855;
  assign n88857 = ~n88847 & ~n88856;
  assign n88858 = ~n88820 & ~n88857;
  assign n88859 = n88808 & n88831;
  assign n88860 = ~n88807 & n88828;
  assign n88861 = ~n88814 & n88860;
  assign n88862 = ~n88801 & n88861;
  assign n88863 = ~n88859 & ~n88862;
  assign n88864 = n88801 & n88831;
  assign n88865 = ~n88814 & n88849;
  assign n88866 = ~n88864 & ~n88865;
  assign n88867 = n88820 & ~n88866;
  assign n88868 = n88863 & ~n88867;
  assign n88869 = ~n88858 & n88868;
  assign n88870 = n88795 & ~n88869;
  assign n88871 = n88801 & ~n88828;
  assign n88872 = n88814 & n88871;
  assign n88873 = ~n88801 & ~n88828;
  assign n88874 = ~n88814 & n88873;
  assign n88875 = ~n88872 & ~n88874;
  assign n88876 = ~n88820 & ~n88875;
  assign n88877 = ~n88801 & ~n88807;
  assign n88878 = ~n88828 & n88877;
  assign n88879 = n88814 & n88878;
  assign n88880 = ~n88859 & ~n88879;
  assign n88881 = ~n88842 & n88880;
  assign n88882 = n88820 & ~n88881;
  assign n88883 = ~n88876 & ~n88882;
  assign n88884 = n88820 & n88860;
  assign n88885 = ~n88814 & n88884;
  assign n88886 = n88883 & ~n88885;
  assign n88887 = ~n88870 & n88886;
  assign n88888 = ~n88853 & n88887;
  assign n88889 = ~pi2848 & ~n88888;
  assign n88890 = pi2848 & n88888;
  assign po2985 = n88889 | n88890;
  assign n88892 = n88814 & n88842;
  assign n88893 = ~n88862 & ~n88871;
  assign n88894 = n88820 & ~n88893;
  assign n88895 = ~n88892 & ~n88894;
  assign n88896 = ~n88856 & n88895;
  assign n88897 = ~n88820 & n88859;
  assign n88898 = ~n88848 & ~n88897;
  assign n88899 = ~n88879 & n88898;
  assign n88900 = n88896 & n88899;
  assign n88901 = n88795 & ~n88900;
  assign n88902 = n88807 & n88831;
  assign n88903 = n88801 & n88902;
  assign n88904 = ~n88833 & ~n88903;
  assign n88905 = ~n88814 & n88878;
  assign n88906 = ~n88843 & ~n88905;
  assign n88907 = n88808 & n88828;
  assign n88908 = n88820 & n88907;
  assign n88909 = n88814 & n88847;
  assign n88910 = ~n88908 & ~n88909;
  assign n88911 = n88807 & ~n88828;
  assign n88912 = n88801 & n88814;
  assign n88913 = ~n88911 & ~n88912;
  assign n88914 = ~n88860 & n88913;
  assign n88915 = ~n88820 & ~n88914;
  assign n88916 = n88910 & ~n88915;
  assign n88917 = n88906 & n88916;
  assign n88918 = n88904 & n88917;
  assign n88919 = ~n88795 & ~n88918;
  assign n88920 = ~n88901 & ~n88919;
  assign n88921 = pi2849 & ~n88920;
  assign n88922 = ~pi2849 & ~n88901;
  assign n88923 = ~n88919 & n88922;
  assign po2987 = n88921 | n88923;
  assign n88925 = pi6624 & pi9040;
  assign n88926 = pi6506 & ~pi9040;
  assign n88927 = ~n88925 & ~n88926;
  assign n88928 = ~pi2845 & ~n88927;
  assign n88929 = pi2845 & n88927;
  assign n88930 = ~n88928 & ~n88929;
  assign n88931 = pi6464 & pi9040;
  assign n88932 = pi6463 & ~pi9040;
  assign n88933 = ~n88931 & ~n88932;
  assign n88934 = ~pi2825 & n88933;
  assign n88935 = pi2825 & ~n88933;
  assign n88936 = ~n88934 & ~n88935;
  assign n88937 = pi6707 & pi9040;
  assign n88938 = pi6501 & ~pi9040;
  assign n88939 = ~n88937 & ~n88938;
  assign n88940 = ~pi2824 & n88939;
  assign n88941 = pi2824 & ~n88939;
  assign n88942 = ~n88940 & ~n88941;
  assign n88943 = pi6681 & ~pi9040;
  assign n88944 = pi6504 & pi9040;
  assign n88945 = ~n88943 & ~n88944;
  assign n88946 = ~pi2831 & n88945;
  assign n88947 = pi2831 & ~n88945;
  assign n88948 = ~n88946 & ~n88947;
  assign n88949 = pi6551 & ~pi9040;
  assign n88950 = pi6501 & pi9040;
  assign n88951 = ~n88949 & ~n88950;
  assign n88952 = ~pi2826 & n88951;
  assign n88953 = pi2826 & ~n88951;
  assign n88954 = ~n88952 & ~n88953;
  assign n88955 = ~n88948 & n88954;
  assign n88956 = ~n88942 & n88955;
  assign n88957 = ~n88936 & n88956;
  assign n88958 = pi2831 & n88945;
  assign n88959 = ~pi2831 & ~n88945;
  assign n88960 = ~n88958 & ~n88959;
  assign n88961 = n88954 & ~n88960;
  assign n88962 = ~n88942 & n88961;
  assign n88963 = n88936 & n88962;
  assign n88964 = ~n88957 & ~n88963;
  assign n88965 = ~n88954 & ~n88960;
  assign n88966 = ~n88942 & n88965;
  assign n88967 = ~n88936 & n88966;
  assign n88968 = pi6409 & pi9040;
  assign n88969 = pi6680 & ~pi9040;
  assign n88970 = ~n88968 & ~n88969;
  assign n88971 = ~pi2847 & ~n88970;
  assign n88972 = pi2847 & n88970;
  assign n88973 = ~n88971 & ~n88972;
  assign n88974 = ~n88948 & ~n88954;
  assign n88975 = ~n88936 & n88974;
  assign n88976 = n88942 & n88965;
  assign n88977 = n88936 & n88976;
  assign n88978 = ~n88975 & ~n88977;
  assign n88979 = ~n88973 & ~n88978;
  assign n88980 = ~n88967 & ~n88979;
  assign n88981 = n88942 & n88961;
  assign n88982 = n88973 & n88981;
  assign n88983 = n88965 & n88973;
  assign n88984 = ~n88936 & n88983;
  assign n88985 = ~n88982 & ~n88984;
  assign n88986 = n88980 & n88985;
  assign n88987 = n88964 & n88986;
  assign n88988 = n88930 & ~n88987;
  assign n88989 = ~n88930 & ~n88973;
  assign n88990 = ~n88936 & n88942;
  assign n88991 = n88948 & n88990;
  assign n88992 = n88942 & n88954;
  assign n88993 = ~n88991 & ~n88992;
  assign n88994 = n88989 & ~n88993;
  assign n88995 = n88936 & ~n88942;
  assign n88996 = ~n88954 & n88995;
  assign n88997 = ~n88960 & n88996;
  assign n88998 = n88936 & ~n88948;
  assign n88999 = n88942 & n88998;
  assign n89000 = ~n88997 & ~n88999;
  assign n89001 = ~n88936 & n88973;
  assign n89002 = ~n88942 & n89001;
  assign n89003 = ~n88965 & n89002;
  assign n89004 = n88956 & n88973;
  assign n89005 = ~n89003 & ~n89004;
  assign n89006 = n89000 & n89005;
  assign n89007 = ~n88930 & ~n89006;
  assign n89008 = n88942 & n88955;
  assign n89009 = ~n88973 & n89008;
  assign n89010 = n88936 & n89009;
  assign n89011 = ~n88942 & n88974;
  assign n89012 = n88936 & n89011;
  assign n89013 = ~n88963 & ~n89012;
  assign n89014 = ~n88973 & ~n89013;
  assign n89015 = ~n89010 & ~n89014;
  assign n89016 = n88973 & n88997;
  assign n89017 = n89015 & ~n89016;
  assign n89018 = ~n89007 & n89017;
  assign n89019 = ~n88994 & n89018;
  assign n89020 = ~n88988 & n89019;
  assign n89021 = n88942 & n88974;
  assign n89022 = n88936 & n88973;
  assign n89023 = n89021 & n89022;
  assign n89024 = n89020 & ~n89023;
  assign n89025 = ~pi2858 & ~n89024;
  assign n89026 = pi2858 & ~n89023;
  assign n89027 = n89020 & n89026;
  assign po2988 = n89025 | n89027;
  assign n89029 = ~n88702 & ~n88729;
  assign n89030 = ~n88708 & n89029;
  assign n89031 = n88714 & n88735;
  assign n89032 = n88702 & n89031;
  assign n89033 = n88702 & n88752;
  assign n89034 = ~n89032 & ~n89033;
  assign n89035 = ~n88702 & n88754;
  assign n89036 = ~n88744 & ~n89035;
  assign n89037 = n88729 & ~n89036;
  assign n89038 = n89034 & ~n89037;
  assign n89039 = ~n89030 & n89038;
  assign n89040 = n88696 & ~n89039;
  assign n89041 = n88702 & n88773;
  assign n89042 = ~n88729 & n89041;
  assign n89043 = n88764 & n88773;
  assign n89044 = ~n88743 & ~n89043;
  assign n89045 = ~n88744 & ~n88767;
  assign n89046 = ~n88702 & n88751;
  assign n89047 = n89045 & ~n89046;
  assign n89048 = ~n88729 & ~n89047;
  assign n89049 = n88729 & n88731;
  assign n89050 = n88756 & ~n89049;
  assign n89051 = ~n89048 & n89050;
  assign n89052 = n89044 & n89051;
  assign n89053 = ~n88696 & ~n89052;
  assign n89054 = ~n89042 & ~n89053;
  assign n89055 = ~n89040 & n89054;
  assign n89056 = n88764 & n88767;
  assign n89057 = n88721 & n88729;
  assign n89058 = n88702 & n89057;
  assign n89059 = ~n89056 & ~n89058;
  assign n89060 = n88729 & n89033;
  assign n89061 = n89059 & ~n89060;
  assign n89062 = n89055 & n89061;
  assign n89063 = ~pi2855 & ~n89062;
  assign n89064 = pi2855 & n89061;
  assign n89065 = n89054 & n89064;
  assign n89066 = ~n89040 & n89065;
  assign po2989 = n89063 | n89066;
  assign n89068 = pi6460 & pi9040;
  assign n89069 = pi6707 & ~pi9040;
  assign n89070 = ~n89068 & ~n89069;
  assign n89071 = ~pi2833 & n89070;
  assign n89072 = pi2833 & ~n89070;
  assign n89073 = ~n89071 & ~n89072;
  assign n89074 = pi6464 & ~pi9040;
  assign n89075 = pi6483 & pi9040;
  assign n89076 = ~n89074 & ~n89075;
  assign n89077 = pi2819 & n89076;
  assign n89078 = ~pi2819 & ~n89076;
  assign n89079 = ~n89077 & ~n89078;
  assign n89080 = pi6495 & pi9040;
  assign n89081 = pi6499 & ~pi9040;
  assign n89082 = ~n89080 & ~n89081;
  assign n89083 = pi2832 & n89082;
  assign n89084 = ~pi2832 & ~n89082;
  assign n89085 = ~n89083 & ~n89084;
  assign n89086 = pi6498 & ~pi9040;
  assign n89087 = pi6508 & pi9040;
  assign n89088 = ~n89086 & ~n89087;
  assign n89089 = ~pi2812 & n89088;
  assign n89090 = pi2812 & ~n89088;
  assign n89091 = ~n89089 & ~n89090;
  assign n89092 = pi6506 & pi9040;
  assign n89093 = pi6602 & ~pi9040;
  assign n89094 = ~n89092 & ~n89093;
  assign n89095 = ~pi2824 & n89094;
  assign n89096 = pi2824 & ~n89094;
  assign n89097 = ~n89095 & ~n89096;
  assign n89098 = n89091 & ~n89097;
  assign n89099 = n89085 & n89098;
  assign n89100 = n89079 & n89099;
  assign n89101 = n89073 & n89100;
  assign n89102 = ~n89091 & n89097;
  assign n89103 = n89073 & n89079;
  assign n89104 = n89102 & n89103;
  assign n89105 = ~n89085 & n89104;
  assign n89106 = ~n89101 & ~n89105;
  assign n89107 = ~n89085 & n89098;
  assign n89108 = n89073 & ~n89079;
  assign n89109 = n89107 & n89108;
  assign n89110 = n89073 & ~n89085;
  assign n89111 = n89097 & n89110;
  assign n89112 = ~n89091 & n89111;
  assign n89113 = ~n89109 & ~n89112;
  assign n89114 = n89085 & ~n89091;
  assign n89115 = ~n89073 & n89114;
  assign n89116 = ~n89073 & n89098;
  assign n89117 = ~n89115 & ~n89116;
  assign n89118 = n89079 & ~n89117;
  assign n89119 = ~n89091 & ~n89097;
  assign n89120 = n89091 & n89097;
  assign n89121 = ~n89119 & ~n89120;
  assign n89122 = ~n89079 & ~n89110;
  assign n89123 = ~n89121 & n89122;
  assign n89124 = n89073 & ~n89098;
  assign n89125 = n89079 & n89124;
  assign n89126 = ~n89085 & n89125;
  assign n89127 = ~n89123 & ~n89126;
  assign n89128 = ~n89118 & n89127;
  assign n89129 = n89113 & n89128;
  assign n89130 = pi6461 & pi9040;
  assign n89131 = pi6502 & ~pi9040;
  assign n89132 = ~n89130 & ~n89131;
  assign n89133 = ~pi2831 & ~n89132;
  assign n89134 = pi2831 & n89132;
  assign n89135 = ~n89133 & ~n89134;
  assign n89136 = ~n89129 & n89135;
  assign n89137 = n89106 & ~n89136;
  assign n89138 = n89085 & n89119;
  assign n89139 = ~n89079 & n89138;
  assign n89140 = ~n89073 & n89139;
  assign n89141 = ~n89079 & ~n89135;
  assign n89142 = n89085 & n89102;
  assign n89143 = ~n89116 & ~n89142;
  assign n89144 = n89110 & ~n89121;
  assign n89145 = n89143 & ~n89144;
  assign n89146 = n89141 & ~n89145;
  assign n89147 = ~n89085 & n89102;
  assign n89148 = ~n89073 & n89147;
  assign n89149 = ~n89073 & ~n89091;
  assign n89150 = ~n89085 & n89149;
  assign n89151 = ~n89073 & n89120;
  assign n89152 = ~n89150 & ~n89151;
  assign n89153 = n89073 & n89098;
  assign n89154 = n89085 & n89120;
  assign n89155 = ~n89153 & ~n89154;
  assign n89156 = n89152 & n89155;
  assign n89157 = n89079 & ~n89156;
  assign n89158 = ~n89148 & ~n89157;
  assign n89159 = ~n89135 & ~n89158;
  assign n89160 = ~n89146 & ~n89159;
  assign n89161 = ~n89140 & n89160;
  assign n89162 = n89137 & n89161;
  assign n89163 = pi2866 & ~n89162;
  assign n89164 = ~pi2866 & n89137;
  assign n89165 = n89161 & n89164;
  assign po2990 = n89163 | n89165;
  assign n89167 = ~n88553 & n88583;
  assign n89168 = n88553 & n88594;
  assign n89169 = ~n88580 & ~n89168;
  assign n89170 = n88527 & ~n89169;
  assign n89171 = ~n89167 & ~n89170;
  assign n89172 = ~n88527 & ~n88553;
  assign n89173 = n88545 & n89172;
  assign n89174 = ~n88539 & n89173;
  assign n89175 = n88561 & n88595;
  assign n89176 = ~n89174 & ~n89175;
  assign n89177 = ~n88527 & n88533;
  assign n89178 = n88555 & n89177;
  assign n89179 = n89176 & ~n89178;
  assign n89180 = ~n88557 & ~n88569;
  assign n89181 = ~n88545 & n88601;
  assign n89182 = n89180 & ~n89181;
  assign n89183 = n89179 & n89182;
  assign n89184 = n89171 & n89183;
  assign n89185 = ~n88592 & ~n89184;
  assign n89186 = ~n88556 & ~n88580;
  assign n89187 = n88553 & ~n89186;
  assign n89188 = ~n88539 & n88598;
  assign n89189 = ~n88609 & ~n89188;
  assign n89190 = n88533 & n88545;
  assign n89191 = n88553 & n89190;
  assign n89192 = n89189 & ~n89191;
  assign n89193 = n88527 & ~n89192;
  assign n89194 = ~n88553 & n88579;
  assign n89195 = ~n88539 & n88568;
  assign n89196 = ~n89194 & ~n89195;
  assign n89197 = ~n88527 & ~n89196;
  assign n89198 = ~n88553 & n88562;
  assign n89199 = ~n89197 & ~n89198;
  assign n89200 = ~n89193 & n89199;
  assign n89201 = ~n89187 & n89200;
  assign n89202 = n88592 & ~n89201;
  assign n89203 = n88527 & n88599;
  assign n89204 = ~n89202 & ~n89203;
  assign n89205 = n88574 & n89172;
  assign n89206 = n88545 & n89205;
  assign n89207 = n89204 & ~n89206;
  assign n89208 = ~n89185 & n89207;
  assign n89209 = ~pi2874 & ~n89208;
  assign n89210 = pi2874 & n89204;
  assign n89211 = ~n89185 & n89210;
  assign n89212 = ~n89206 & n89211;
  assign po2991 = n89209 | n89212;
  assign n89214 = pi6495 & ~pi9040;
  assign n89215 = pi6503 & pi9040;
  assign n89216 = ~n89214 & ~n89215;
  assign n89217 = pi2836 & n89216;
  assign n89218 = ~pi2836 & ~n89216;
  assign n89219 = ~n89217 & ~n89218;
  assign n89220 = pi6499 & pi9040;
  assign n89221 = pi6698 & ~pi9040;
  assign n89222 = ~n89220 & ~n89221;
  assign n89223 = ~pi2846 & ~n89222;
  assign n89224 = pi2846 & n89222;
  assign n89225 = ~n89223 & ~n89224;
  assign n89226 = pi6460 & ~pi9040;
  assign n89227 = pi6514 & pi9040;
  assign n89228 = ~n89226 & ~n89227;
  assign n89229 = ~pi2830 & ~n89228;
  assign n89230 = pi2830 & n89228;
  assign n89231 = ~n89229 & ~n89230;
  assign n89232 = ~n89225 & n89231;
  assign n89233 = pi6507 & ~pi9040;
  assign n89234 = pi6745 & pi9040;
  assign n89235 = ~n89233 & ~n89234;
  assign n89236 = ~pi2822 & ~n89235;
  assign n89237 = pi2822 & n89235;
  assign n89238 = ~n89236 & ~n89237;
  assign n89239 = n89225 & n89238;
  assign n89240 = pi6603 & ~pi9040;
  assign n89241 = pi6681 & pi9040;
  assign n89242 = ~n89240 & ~n89241;
  assign n89243 = ~pi2823 & n89242;
  assign n89244 = pi2823 & ~n89242;
  assign n89245 = ~n89243 & ~n89244;
  assign n89246 = ~n89231 & n89245;
  assign n89247 = n89239 & n89246;
  assign n89248 = ~n89232 & ~n89247;
  assign n89249 = ~n89225 & ~n89245;
  assign n89250 = n89248 & ~n89249;
  assign n89251 = n89219 & ~n89250;
  assign n89252 = ~n89219 & ~n89245;
  assign n89253 = n89225 & n89252;
  assign n89254 = ~n89225 & ~n89231;
  assign n89255 = ~n89219 & n89245;
  assign n89256 = n89254 & n89255;
  assign n89257 = n89231 & ~n89245;
  assign n89258 = n89238 & n89257;
  assign n89259 = n89225 & ~n89238;
  assign n89260 = n89231 & n89259;
  assign n89261 = n89245 & n89260;
  assign n89262 = ~n89258 & ~n89261;
  assign n89263 = ~n89256 & n89262;
  assign n89264 = ~n89253 & n89263;
  assign n89265 = ~n89251 & n89264;
  assign n89266 = pi6405 & pi9040;
  assign n89267 = pi6503 & ~pi9040;
  assign n89268 = ~n89266 & ~n89267;
  assign n89269 = pi2834 & n89268;
  assign n89270 = ~pi2834 & ~n89268;
  assign n89271 = ~n89269 & ~n89270;
  assign n89272 = ~n89265 & n89271;
  assign n89273 = ~n89225 & n89238;
  assign n89274 = n89231 & n89273;
  assign n89275 = n89245 & n89274;
  assign n89276 = n89232 & ~n89238;
  assign n89277 = ~n89245 & n89276;
  assign n89278 = ~n89275 & ~n89277;
  assign n89279 = n89219 & ~n89278;
  assign n89280 = ~n89272 & ~n89279;
  assign n89281 = ~n89245 & n89260;
  assign n89282 = n89225 & n89231;
  assign n89283 = n89238 & n89282;
  assign n89284 = ~n89231 & ~n89238;
  assign n89285 = n89225 & n89284;
  assign n89286 = ~n89283 & ~n89285;
  assign n89287 = n89219 & ~n89286;
  assign n89288 = ~n89281 & ~n89287;
  assign n89289 = ~n89231 & n89273;
  assign n89290 = ~n89245 & n89289;
  assign n89291 = n89288 & ~n89290;
  assign n89292 = ~n89271 & ~n89291;
  assign n89293 = ~n89225 & ~n89238;
  assign n89294 = ~n89239 & ~n89293;
  assign n89295 = ~n89231 & ~n89294;
  assign n89296 = n89245 & n89293;
  assign n89297 = ~n89295 & ~n89296;
  assign n89298 = ~n89219 & ~n89297;
  assign n89299 = ~n89271 & n89298;
  assign n89300 = ~n89292 & ~n89299;
  assign n89301 = n89280 & n89300;
  assign n89302 = pi2854 & ~n89301;
  assign n89303 = ~pi2854 & n89280;
  assign n89304 = n89300 & n89303;
  assign po2992 = n89302 | n89304;
  assign n89306 = n88936 & n88981;
  assign n89307 = n88954 & n88990;
  assign n89308 = ~n88948 & n89307;
  assign n89309 = ~n89306 & ~n89308;
  assign n89310 = n88973 & ~n89309;
  assign n89311 = ~n88973 & n88997;
  assign n89312 = ~n88997 & ~n89004;
  assign n89313 = ~n88960 & n88995;
  assign n89314 = ~n88999 & ~n89313;
  assign n89315 = ~n88973 & ~n89314;
  assign n89316 = ~n88936 & ~n88973;
  assign n89317 = n88961 & n89316;
  assign n89318 = n88942 & n89317;
  assign n89319 = ~n88936 & ~n88942;
  assign n89320 = ~n88954 & n89319;
  assign n89321 = ~n88948 & n89320;
  assign n89322 = n88973 & n88976;
  assign n89323 = ~n89321 & ~n89322;
  assign n89324 = ~n89318 & n89323;
  assign n89325 = ~n89315 & n89324;
  assign n89326 = n89312 & n89325;
  assign n89327 = n88930 & ~n89326;
  assign n89328 = n88955 & n89022;
  assign n89329 = ~n88942 & n89328;
  assign n89330 = ~n89327 & ~n89329;
  assign n89331 = ~n89311 & n89330;
  assign n89332 = ~n89310 & n89331;
  assign n89333 = ~n88942 & ~n88960;
  assign n89334 = n89001 & n89333;
  assign n89335 = ~n88982 & ~n89334;
  assign n89336 = n88973 & n89011;
  assign n89337 = n88936 & n89021;
  assign n89338 = ~n89336 & ~n89337;
  assign n89339 = ~n88936 & n88962;
  assign n89340 = ~n89306 & ~n89339;
  assign n89341 = ~n88936 & n88955;
  assign n89342 = n88942 & ~n88954;
  assign n89343 = ~n89341 & ~n89342;
  assign n89344 = ~n88973 & ~n89343;
  assign n89345 = n89340 & ~n89344;
  assign n89346 = n89338 & n89345;
  assign n89347 = n89335 & n89346;
  assign n89348 = ~n88930 & ~n89347;
  assign n89349 = n89332 & ~n89348;
  assign n89350 = ~pi2860 & ~n89349;
  assign n89351 = pi2860 & n89332;
  assign n89352 = ~n89348 & n89351;
  assign po2994 = n89350 | n89352;
  assign n89354 = pi6603 & pi9040;
  assign n89355 = pi6405 & ~pi9040;
  assign n89356 = ~n89354 & ~n89355;
  assign n89357 = pi2838 & n89356;
  assign n89358 = ~pi2838 & ~n89356;
  assign n89359 = ~n89357 & ~n89358;
  assign n89360 = pi6461 & ~pi9040;
  assign n89361 = pi6602 & pi9040;
  assign n89362 = ~n89360 & ~n89361;
  assign n89363 = ~pi2834 & ~n89362;
  assign n89364 = pi2834 & n89362;
  assign n89365 = ~n89363 & ~n89364;
  assign n89366 = pi6745 & ~pi9040;
  assign n89367 = pi6421 & pi9040;
  assign n89368 = ~n89366 & ~n89367;
  assign n89369 = pi2832 & n89368;
  assign n89370 = ~pi2832 & ~n89368;
  assign n89371 = ~n89369 & ~n89370;
  assign n89372 = n89365 & ~n89371;
  assign n89373 = pi6680 & pi9040;
  assign n89374 = pi6421 & ~pi9040;
  assign n89375 = ~n89373 & ~n89374;
  assign n89376 = pi2837 & n89375;
  assign n89377 = ~pi2837 & ~n89375;
  assign n89378 = ~n89376 & ~n89377;
  assign n89379 = pi6507 & pi9040;
  assign n89380 = pi6508 & ~pi9040;
  assign n89381 = ~n89379 & ~n89380;
  assign n89382 = ~pi2822 & n89381;
  assign n89383 = pi2822 & ~n89381;
  assign n89384 = ~n89382 & ~n89383;
  assign n89385 = n89378 & ~n89384;
  assign n89386 = n89372 & n89385;
  assign n89387 = n89378 & n89384;
  assign n89388 = ~n89365 & n89387;
  assign n89389 = ~n89386 & ~n89388;
  assign n89390 = ~n89359 & ~n89389;
  assign n89391 = pi6502 & pi9040;
  assign n89392 = pi6504 & ~pi9040;
  assign n89393 = ~n89391 & ~n89392;
  assign n89394 = ~pi2812 & ~n89393;
  assign n89395 = pi2812 & n89393;
  assign n89396 = ~n89394 & ~n89395;
  assign n89397 = n89359 & ~n89378;
  assign n89398 = n89365 & n89397;
  assign n89399 = n89372 & n89384;
  assign n89400 = n89365 & n89371;
  assign n89401 = ~n89384 & n89400;
  assign n89402 = ~n89399 & ~n89401;
  assign n89403 = ~n89365 & ~n89371;
  assign n89404 = ~n89384 & n89403;
  assign n89405 = n89378 & n89404;
  assign n89406 = n89402 & ~n89405;
  assign n89407 = n89359 & ~n89406;
  assign n89408 = ~n89398 & ~n89407;
  assign n89409 = ~n89365 & n89371;
  assign n89410 = n89384 & n89409;
  assign n89411 = n89378 & n89410;
  assign n89412 = n89408 & ~n89411;
  assign n89413 = ~n89378 & n89403;
  assign n89414 = ~n89384 & n89409;
  assign n89415 = ~n89413 & ~n89414;
  assign n89416 = ~n89359 & ~n89415;
  assign n89417 = n89384 & n89400;
  assign n89418 = ~n89378 & n89417;
  assign n89419 = ~n89416 & ~n89418;
  assign n89420 = n89412 & n89419;
  assign n89421 = n89396 & ~n89420;
  assign n89422 = ~n89390 & ~n89421;
  assign n89423 = n89359 & ~n89396;
  assign n89424 = ~n89415 & n89423;
  assign n89425 = n89384 & n89403;
  assign n89426 = ~n89417 & ~n89425;
  assign n89427 = n89378 & ~n89426;
  assign n89428 = ~n89386 & ~n89427;
  assign n89429 = ~n89396 & ~n89428;
  assign n89430 = ~n89424 & ~n89429;
  assign n89431 = ~n89359 & ~n89396;
  assign n89432 = n89372 & ~n89378;
  assign n89433 = ~n89410 & ~n89432;
  assign n89434 = n89365 & ~n89384;
  assign n89435 = n89433 & ~n89434;
  assign n89436 = n89431 & ~n89435;
  assign n89437 = n89430 & ~n89436;
  assign n89438 = n89422 & n89437;
  assign n89439 = ~pi2853 & ~n89438;
  assign n89440 = pi2853 & n89430;
  assign n89441 = n89422 & n89440;
  assign n89442 = ~n89436 & n89441;
  assign po2995 = n89439 | n89442;
  assign n89444 = n89219 & ~n89245;
  assign n89445 = n89273 & n89444;
  assign n89446 = n89231 & n89445;
  assign n89447 = n89219 & n89245;
  assign n89448 = n89239 & n89447;
  assign n89449 = n89231 & n89245;
  assign n89450 = ~n89238 & n89449;
  assign n89451 = ~n89225 & n89450;
  assign n89452 = n89219 & n89260;
  assign n89453 = ~n89245 & n89452;
  assign n89454 = ~n89451 & ~n89453;
  assign n89455 = ~n89448 & n89454;
  assign n89456 = ~n89446 & n89455;
  assign n89457 = ~n89247 & n89456;
  assign n89458 = ~n89271 & ~n89457;
  assign n89459 = ~n89245 & n89283;
  assign n89460 = ~n89450 & ~n89459;
  assign n89461 = ~n89290 & n89460;
  assign n89462 = ~n89219 & ~n89461;
  assign n89463 = ~n89219 & n89285;
  assign n89464 = ~n89245 & n89463;
  assign n89465 = ~n89225 & n89449;
  assign n89466 = ~n89296 & ~n89465;
  assign n89467 = ~n89219 & ~n89466;
  assign n89468 = ~n89464 & ~n89467;
  assign n89469 = ~n89271 & ~n89468;
  assign n89470 = ~n89462 & ~n89469;
  assign n89471 = ~n89458 & n89470;
  assign n89472 = ~n89231 & ~n89245;
  assign n89473 = n89219 & n89472;
  assign n89474 = n89293 & n89473;
  assign n89475 = ~n89231 & n89447;
  assign n89476 = n89225 & n89475;
  assign n89477 = n89245 & n89285;
  assign n89478 = ~n89219 & n89231;
  assign n89479 = n89225 & n89478;
  assign n89480 = ~n89231 & n89249;
  assign n89481 = ~n89479 & ~n89480;
  assign n89482 = ~n89477 & n89481;
  assign n89483 = ~n89289 & n89482;
  assign n89484 = n89219 & n89273;
  assign n89485 = n89245 & n89484;
  assign n89486 = ~n89245 & n89293;
  assign n89487 = ~n89231 & n89238;
  assign n89488 = ~n89486 & ~n89487;
  assign n89489 = n89219 & ~n89488;
  assign n89490 = ~n89485 & ~n89489;
  assign n89491 = n89483 & n89490;
  assign n89492 = n89271 & ~n89491;
  assign n89493 = ~n89476 & ~n89492;
  assign n89494 = ~n89474 & n89493;
  assign n89495 = n89471 & n89494;
  assign n89496 = pi2850 & n89495;
  assign n89497 = ~pi2850 & ~n89495;
  assign po2996 = n89496 | n89497;
  assign n89499 = ~n88554 & ~n88560;
  assign n89500 = ~n88527 & ~n89499;
  assign n89501 = ~n88616 & ~n89500;
  assign n89502 = ~n88533 & n88539;
  assign n89503 = n88527 & n89502;
  assign n89504 = n88553 & n89503;
  assign n89505 = n88553 & n88579;
  assign n89506 = ~n89502 & ~n89505;
  assign n89507 = n88533 & ~n88553;
  assign n89508 = ~n88539 & n89507;
  assign n89509 = n89506 & ~n89508;
  assign n89510 = n88527 & ~n89509;
  assign n89511 = ~n88563 & ~n89510;
  assign n89512 = ~n88592 & ~n89511;
  assign n89513 = ~n88527 & n88546;
  assign n89514 = n88553 & n89513;
  assign n89515 = ~n89178 & ~n89514;
  assign n89516 = ~n88592 & ~n89515;
  assign n89517 = ~n89512 & ~n89516;
  assign n89518 = ~n89504 & n89517;
  assign n89519 = ~n88580 & ~n88599;
  assign n89520 = ~n88609 & n89519;
  assign n89521 = ~n88527 & ~n89520;
  assign n89522 = ~n88553 & n88559;
  assign n89523 = ~n88583 & ~n89522;
  assign n89524 = n88527 & ~n89523;
  assign n89525 = ~n89521 & ~n89524;
  assign n89526 = ~n89188 & n89525;
  assign n89527 = ~n88569 & ~n88610;
  assign n89528 = n89526 & n89527;
  assign n89529 = n88592 & ~n89528;
  assign n89530 = n89518 & ~n89529;
  assign n89531 = n89501 & n89530;
  assign n89532 = ~pi2893 & ~n89531;
  assign n89533 = pi2893 & n89518;
  assign n89534 = n89501 & n89533;
  assign n89535 = ~n89529 & n89534;
  assign po2997 = n89532 | n89535;
  assign n89537 = ~n88814 & n88835;
  assign n89538 = ~n88905 & ~n89537;
  assign n89539 = n88820 & n89538;
  assign n89540 = ~n88808 & ~n88829;
  assign n89541 = ~n88828 & ~n89540;
  assign n89542 = n88814 & n88873;
  assign n89543 = ~n88801 & n88854;
  assign n89544 = n88814 & n88829;
  assign n89545 = ~n89543 & ~n89544;
  assign n89546 = ~n89542 & n89545;
  assign n89547 = ~n89541 & n89546;
  assign n89548 = ~n88820 & n89547;
  assign n89549 = ~n89539 & ~n89548;
  assign n89550 = n88814 & n89541;
  assign n89551 = ~n88903 & ~n89550;
  assign n89552 = ~n89549 & n89551;
  assign n89553 = n88795 & ~n89552;
  assign n89554 = n88820 & ~n89540;
  assign n89555 = ~n88814 & n89554;
  assign n89556 = ~n88849 & ~n88877;
  assign n89557 = n88814 & ~n89556;
  assign n89558 = n88820 & n89557;
  assign n89559 = n88828 & n89554;
  assign n89560 = ~n89558 & ~n89559;
  assign n89561 = ~n89555 & n89560;
  assign n89562 = ~n88795 & ~n89561;
  assign n89563 = ~n89553 & ~n89562;
  assign n89564 = ~n88820 & ~n89538;
  assign n89565 = ~n88833 & ~n89564;
  assign n89566 = ~n88795 & ~n89565;
  assign n89567 = n88820 & n88833;
  assign n89568 = ~n88820 & ~n89551;
  assign n89569 = ~n89567 & ~n89568;
  assign n89570 = ~n89566 & n89569;
  assign n89571 = n89563 & n89570;
  assign n89572 = pi2856 & ~n89571;
  assign n89573 = ~pi2856 & n89570;
  assign n89574 = ~n89562 & n89573;
  assign n89575 = ~n89553 & n89574;
  assign po2998 = n89572 | n89575;
  assign n89577 = ~n89245 & n89295;
  assign n89578 = ~n89274 & ~n89284;
  assign n89579 = ~n89219 & ~n89578;
  assign n89580 = ~n89577 & ~n89579;
  assign n89581 = ~n89238 & n89257;
  assign n89582 = ~n89487 & ~n89581;
  assign n89583 = ~n89276 & n89582;
  assign n89584 = n89219 & ~n89583;
  assign n89585 = n89580 & ~n89584;
  assign n89586 = n89245 & n89283;
  assign n89587 = n89585 & ~n89586;
  assign n89588 = ~n89271 & ~n89587;
  assign n89589 = n89447 & ~n89578;
  assign n89590 = ~n89285 & ~n89289;
  assign n89591 = ~n89276 & ~n89283;
  assign n89592 = n89590 & n89591;
  assign n89593 = ~n89245 & ~n89592;
  assign n89594 = ~n89589 & ~n89593;
  assign n89595 = ~n89261 & n89594;
  assign n89596 = n89271 & ~n89595;
  assign n89597 = ~n89588 & ~n89596;
  assign n89598 = ~n89245 & n89274;
  assign n89599 = ~n89586 & ~n89598;
  assign n89600 = ~n89219 & ~n89599;
  assign n89601 = n89597 & ~n89600;
  assign n89602 = pi2865 & ~n89601;
  assign n89603 = ~pi2865 & ~n89600;
  assign n89604 = ~n89596 & n89603;
  assign n89605 = ~n89588 & n89604;
  assign po2999 = n89602 | n89605;
  assign n89607 = ~n89329 & ~n89334;
  assign n89608 = ~n88997 & ~n89008;
  assign n89609 = ~n89341 & n89608;
  assign n89610 = ~n88973 & ~n89609;
  assign n89611 = ~n88936 & n88976;
  assign n89612 = ~n89321 & ~n89611;
  assign n89613 = ~n89023 & n89612;
  assign n89614 = n88962 & n88973;
  assign n89615 = n89613 & ~n89614;
  assign n89616 = ~n89610 & n89615;
  assign n89617 = n88930 & ~n89616;
  assign n89618 = n88936 & n88983;
  assign n89619 = n88960 & n88990;
  assign n89620 = ~n89008 & ~n89619;
  assign n89621 = n88973 & ~n89620;
  assign n89622 = ~n89618 & ~n89621;
  assign n89623 = ~n88973 & n88974;
  assign n89624 = n88936 & n89623;
  assign n89625 = ~n88973 & n88981;
  assign n89626 = ~n89624 & ~n89625;
  assign n89627 = n89622 & n89626;
  assign n89628 = n88960 & n88995;
  assign n89629 = ~n89306 & ~n89628;
  assign n89630 = ~n89339 & n89629;
  assign n89631 = n89627 & n89630;
  assign n89632 = ~n88930 & ~n89631;
  assign n89633 = ~n89306 & n89612;
  assign n89634 = ~n88973 & ~n89633;
  assign n89635 = ~n89632 & ~n89634;
  assign n89636 = ~n89617 & n89635;
  assign n89637 = n89607 & n89636;
  assign n89638 = pi2875 & ~n89637;
  assign n89639 = ~pi2875 & n89637;
  assign po3000 = n89638 | n89639;
  assign n89641 = n89245 & n89289;
  assign n89642 = ~n89261 & ~n89641;
  assign n89643 = ~n89219 & ~n89642;
  assign n89644 = n89252 & n89283;
  assign n89645 = ~n89643 & ~n89644;
  assign n89646 = ~n89476 & n89645;
  assign n89647 = n89219 & n89231;
  assign n89648 = ~n89238 & n89647;
  assign n89649 = ~n89225 & n89648;
  assign n89650 = n89245 & n89649;
  assign n89651 = ~n89245 & n89285;
  assign n89652 = ~n89289 & ~n89651;
  assign n89653 = ~n89276 & n89652;
  assign n89654 = ~n89219 & ~n89653;
  assign n89655 = n89271 & n89654;
  assign n89656 = n89219 & n89274;
  assign n89657 = ~n89247 & ~n89474;
  assign n89658 = ~n89453 & n89657;
  assign n89659 = ~n89656 & n89658;
  assign n89660 = n89271 & ~n89659;
  assign n89661 = ~n89245 & n89484;
  assign n89662 = ~n89649 & ~n89661;
  assign n89663 = ~n89258 & n89662;
  assign n89664 = ~n89238 & n89246;
  assign n89665 = n89239 & ~n89245;
  assign n89666 = ~n89282 & ~n89665;
  assign n89667 = ~n89219 & ~n89666;
  assign n89668 = ~n89664 & ~n89667;
  assign n89669 = n89663 & n89668;
  assign n89670 = ~n89271 & ~n89669;
  assign n89671 = ~n89660 & ~n89670;
  assign n89672 = ~n89655 & n89671;
  assign n89673 = ~n89650 & n89672;
  assign n89674 = n89646 & n89673;
  assign n89675 = pi2864 & ~n89674;
  assign n89676 = ~pi2864 & n89646;
  assign n89677 = n89673 & n89676;
  assign po3001 = n89675 | n89677;
  assign n89679 = ~n89138 & ~n89147;
  assign n89680 = n89073 & n89085;
  assign n89681 = ~n89097 & n89680;
  assign n89682 = n89679 & ~n89681;
  assign n89683 = ~n89079 & n89135;
  assign n89684 = ~n89682 & n89683;
  assign n89685 = ~n89073 & n89135;
  assign n89686 = n89154 & n89685;
  assign n89687 = n89079 & n89142;
  assign n89688 = ~n89085 & ~n89097;
  assign n89689 = ~n89116 & ~n89688;
  assign n89690 = n89079 & ~n89689;
  assign n89691 = ~n89687 & ~n89690;
  assign n89692 = n89135 & ~n89691;
  assign n89693 = ~n89686 & ~n89692;
  assign n89694 = n89091 & n89111;
  assign n89695 = ~n89073 & ~n89085;
  assign n89696 = ~n89097 & n89695;
  assign n89697 = ~n89694 & ~n89696;
  assign n89698 = n89079 & ~n89697;
  assign n89699 = n89693 & ~n89698;
  assign n89700 = ~n89073 & ~n89079;
  assign n89701 = n89098 & n89700;
  assign n89702 = n89085 & n89701;
  assign n89703 = ~n89121 & n89680;
  assign n89704 = ~n89112 & ~n89703;
  assign n89705 = ~n89121 & n89695;
  assign n89706 = ~n89073 & n89142;
  assign n89707 = ~n89705 & ~n89706;
  assign n89708 = ~n89109 & n89707;
  assign n89709 = n89704 & n89708;
  assign n89710 = ~n89702 & n89709;
  assign n89711 = n89085 & n89103;
  assign n89712 = n89091 & n89711;
  assign n89713 = n89710 & ~n89712;
  assign n89714 = ~n89135 & ~n89713;
  assign n89715 = n89699 & ~n89714;
  assign n89716 = ~n89684 & n89715;
  assign n89717 = ~pi2876 & ~n89716;
  assign n89718 = pi2876 & n89699;
  assign n89719 = ~n89684 & n89718;
  assign n89720 = ~n89714 & n89719;
  assign po3002 = n89717 | n89720;
  assign n89722 = ~n88702 & n89031;
  assign n89723 = n88702 & n88721;
  assign n89724 = ~n88702 & n88773;
  assign n89725 = ~n89723 & ~n89724;
  assign n89726 = ~n88752 & ~n88760;
  assign n89727 = n89725 & n89726;
  assign n89728 = ~n88729 & ~n89727;
  assign n89729 = n88702 & n88730;
  assign n89730 = ~n88743 & ~n89729;
  assign n89731 = ~n88754 & n89730;
  assign n89732 = n88729 & ~n89731;
  assign n89733 = n88702 & ~n88714;
  assign n89734 = n88720 & n89733;
  assign n89735 = ~n88708 & n89734;
  assign n89736 = ~n89732 & ~n89735;
  assign n89737 = ~n89728 & n89736;
  assign n89738 = ~n89722 & n89737;
  assign n89739 = ~n88696 & ~n89738;
  assign n89740 = n88702 & ~n88729;
  assign n89741 = n88731 & n89740;
  assign n89742 = ~n88729 & n88754;
  assign n89743 = ~n88729 & n88767;
  assign n89744 = ~n89742 & ~n89743;
  assign n89745 = ~n88702 & ~n89744;
  assign n89746 = ~n89741 & ~n89745;
  assign n89747 = n88702 & n88751;
  assign n89748 = ~n88702 & n88730;
  assign n89749 = ~n89747 & ~n89748;
  assign n89750 = ~n88722 & n89749;
  assign n89751 = ~n88752 & n89750;
  assign n89752 = n88729 & ~n89751;
  assign n89753 = ~n88702 & n88744;
  assign n89754 = ~n89752 & ~n89753;
  assign n89755 = ~n88702 & n88722;
  assign n89756 = ~n89041 & ~n89755;
  assign n89757 = n89754 & n89756;
  assign n89758 = n89746 & n89757;
  assign n89759 = n88696 & ~n89758;
  assign n89760 = ~n88729 & ~n89034;
  assign n89761 = ~n89759 & ~n89760;
  assign n89762 = ~n88755 & ~n89755;
  assign n89763 = n88729 & ~n89762;
  assign n89764 = n89761 & ~n89763;
  assign n89765 = ~n89739 & n89764;
  assign n89766 = pi2862 & ~n89765;
  assign n89767 = ~pi2862 & n89765;
  assign po3003 = n89766 | n89767;
  assign n89769 = ~n89359 & ~n89377;
  assign n89770 = ~n89376 & n89769;
  assign n89771 = ~n89403 & ~n89417;
  assign n89772 = n89770 & ~n89771;
  assign n89773 = ~n89359 & n89384;
  assign n89774 = n89403 & n89773;
  assign n89775 = ~n89772 & ~n89774;
  assign n89776 = n89396 & ~n89775;
  assign n89777 = ~n89378 & n89401;
  assign n89778 = ~n89378 & ~n89384;
  assign n89779 = ~n89434 & ~n89778;
  assign n89780 = n89359 & ~n89779;
  assign n89781 = ~n89378 & n89384;
  assign n89782 = ~n89371 & n89781;
  assign n89783 = n89365 & n89782;
  assign n89784 = ~n89780 & ~n89783;
  assign n89785 = ~n89777 & n89784;
  assign n89786 = n89396 & ~n89785;
  assign n89787 = ~n89776 & ~n89786;
  assign n89788 = n89371 & n89385;
  assign n89789 = ~n89365 & n89788;
  assign n89790 = ~n89378 & n89410;
  assign n89791 = ~n89789 & ~n89790;
  assign n89792 = ~n89359 & ~n89791;
  assign n89793 = ~n89371 & n89387;
  assign n89794 = ~n89365 & n89793;
  assign n89795 = ~n89378 & n89434;
  assign n89796 = ~n89794 & ~n89795;
  assign n89797 = n89359 & ~n89796;
  assign n89798 = ~n89372 & ~n89434;
  assign n89799 = n89378 & ~n89798;
  assign n89800 = ~n89410 & ~n89799;
  assign n89801 = ~n89359 & ~n89800;
  assign n89802 = n89371 & ~n89378;
  assign n89803 = n89773 & n89802;
  assign n89804 = ~n89371 & ~n89384;
  assign n89805 = ~n89410 & ~n89804;
  assign n89806 = ~n89378 & ~n89805;
  assign n89807 = n89359 & n89378;
  assign n89808 = n89400 & n89807;
  assign n89809 = n89384 & n89808;
  assign n89810 = ~n89806 & ~n89809;
  assign n89811 = ~n89803 & n89810;
  assign n89812 = ~n89801 & n89811;
  assign n89813 = ~n89789 & n89812;
  assign n89814 = ~n89396 & ~n89813;
  assign n89815 = ~n89797 & ~n89814;
  assign n89816 = ~n89792 & n89815;
  assign n89817 = n89787 & n89816;
  assign n89818 = pi2863 & n89817;
  assign n89819 = ~pi2863 & ~n89817;
  assign po3005 = n89818 | n89819;
  assign n89821 = ~n89151 & ~n89153;
  assign n89822 = n89079 & ~n89821;
  assign n89823 = ~n89105 & ~n89822;
  assign n89824 = n89135 & ~n89823;
  assign n89825 = ~n89085 & ~n89091;
  assign n89826 = ~n89119 & ~n89825;
  assign n89827 = n89073 & ~n89826;
  assign n89828 = ~n89099 & ~n89827;
  assign n89829 = ~n89079 & ~n89828;
  assign n89830 = ~n89144 & ~n89829;
  assign n89831 = ~n89073 & n89107;
  assign n89832 = n89097 & n89680;
  assign n89833 = ~n89073 & ~n89826;
  assign n89834 = ~n89832 & ~n89833;
  assign n89835 = n89079 & ~n89834;
  assign n89836 = ~n89831 & ~n89835;
  assign n89837 = n89830 & n89836;
  assign n89838 = ~n89135 & ~n89837;
  assign n89839 = ~n89073 & n89085;
  assign n89840 = ~n89119 & n89839;
  assign n89841 = n89135 & n89840;
  assign n89842 = n89119 & n89695;
  assign n89843 = n89079 & n89842;
  assign n89844 = n89085 & n89097;
  assign n89845 = n89700 & n89844;
  assign n89846 = ~n89843 & ~n89845;
  assign n89847 = ~n89841 & n89846;
  assign n89848 = ~n89149 & ~n89154;
  assign n89849 = n89683 & ~n89848;
  assign n89850 = n89847 & ~n89849;
  assign n89851 = ~n89838 & n89850;
  assign n89852 = ~n89824 & n89851;
  assign n89853 = pi2884 & ~n89852;
  assign n89854 = ~pi2884 & n89852;
  assign po3006 = n89853 | n89854;
  assign n89856 = ~n89085 & n89119;
  assign n89857 = ~n89099 & ~n89856;
  assign n89858 = n89079 & ~n89857;
  assign n89859 = n89073 & n89120;
  assign n89860 = ~n89138 & ~n89859;
  assign n89861 = ~n89107 & n89860;
  assign n89862 = ~n89079 & ~n89861;
  assign n89863 = ~n89858 & ~n89862;
  assign n89864 = ~n89687 & ~n89694;
  assign n89865 = n89863 & n89864;
  assign n89866 = ~n89135 & ~n89865;
  assign n89867 = ~n89073 & n89099;
  assign n89868 = n89073 & n89102;
  assign n89869 = ~n89151 & ~n89868;
  assign n89870 = ~n89079 & ~n89869;
  assign n89871 = ~n89867 & ~n89870;
  assign n89872 = n89079 & n89085;
  assign n89873 = n89097 & n89872;
  assign n89874 = n89091 & n89873;
  assign n89875 = n89679 & ~n89874;
  assign n89876 = ~n89107 & n89875;
  assign n89877 = n89073 & ~n89876;
  assign n89878 = n89871 & ~n89877;
  assign n89879 = n89135 & ~n89878;
  assign n89880 = ~n89866 & ~n89879;
  assign n89881 = ~n89085 & n89151;
  assign n89882 = ~n89706 & ~n89881;
  assign n89883 = n89079 & ~n89882;
  assign n89884 = n89700 & n89825;
  assign n89885 = ~n89883 & ~n89884;
  assign n89886 = n89880 & n89885;
  assign n89887 = ~pi2883 & ~n89886;
  assign n89888 = n89880 & ~n89883;
  assign n89889 = pi2883 & n89888;
  assign n89890 = ~n89884 & n89889;
  assign po3007 = n89887 | n89890;
  assign n89892 = ~n89035 & ~n89755;
  assign n89893 = ~n89735 & n89892;
  assign n89894 = ~n88729 & ~n89893;
  assign n89895 = ~n89041 & ~n89743;
  assign n89896 = ~n89031 & ~n89748;
  assign n89897 = n88729 & ~n89896;
  assign n89898 = ~n88760 & ~n89897;
  assign n89899 = n89895 & n89898;
  assign n89900 = n88696 & ~n89899;
  assign n89901 = ~n88714 & n88720;
  assign n89902 = ~n88732 & ~n89901;
  assign n89903 = n88702 & ~n89902;
  assign n89904 = ~n88722 & ~n89046;
  assign n89905 = n88729 & ~n89904;
  assign n89906 = n88702 & n88720;
  assign n89907 = ~n88744 & ~n89906;
  assign n89908 = ~n88735 & n89907;
  assign n89909 = ~n88729 & ~n89908;
  assign n89910 = ~n89905 & ~n89909;
  assign n89911 = ~n89903 & n89910;
  assign n89912 = ~n88696 & ~n89911;
  assign n89913 = ~n89900 & ~n89912;
  assign n89914 = ~n89043 & ~n89060;
  assign n89915 = n89913 & n89914;
  assign n89916 = ~n89894 & n89915;
  assign n89917 = ~pi2871 & ~n89916;
  assign n89918 = pi2871 & n89914;
  assign n89919 = ~n89894 & n89918;
  assign n89920 = n89913 & n89919;
  assign po3008 = n89917 | n89920;
  assign n89922 = n88814 & n88907;
  assign n89923 = n88820 & n89922;
  assign n89924 = n88854 & ~n89540;
  assign n89925 = ~n88878 & ~n88903;
  assign n89926 = ~n89924 & n89925;
  assign n89927 = ~n88820 & ~n89926;
  assign n89928 = n88814 & n88830;
  assign n89929 = ~n89927 & ~n89928;
  assign n89930 = n88828 & n88877;
  assign n89931 = ~n88814 & n88911;
  assign n89932 = ~n89930 & ~n89931;
  assign n89933 = ~n89544 & n89932;
  assign n89934 = n88820 & ~n89933;
  assign n89935 = n89929 & ~n89934;
  assign n89936 = n88795 & ~n89935;
  assign n89937 = ~n89923 & ~n89936;
  assign n89938 = ~n88814 & n88829;
  assign n89939 = n88828 & n88835;
  assign n89940 = ~n89938 & ~n89939;
  assign n89941 = n88820 & ~n89940;
  assign n89942 = ~n88879 & ~n89941;
  assign n89943 = ~n88850 & ~n89922;
  assign n89944 = n88814 & n88860;
  assign n89945 = ~n88911 & ~n89944;
  assign n89946 = ~n89930 & n89945;
  assign n89947 = ~n88820 & ~n89946;
  assign n89948 = ~n88814 & n88830;
  assign n89949 = ~n89947 & ~n89948;
  assign n89950 = n89943 & n89949;
  assign n89951 = n89942 & n89950;
  assign n89952 = ~n88795 & ~n89951;
  assign n89953 = ~n88865 & ~n89542;
  assign n89954 = ~n88820 & ~n89953;
  assign n89955 = ~n89952 & ~n89954;
  assign n89956 = n89937 & n89955;
  assign n89957 = pi2859 & n89956;
  assign n89958 = ~pi2859 & ~n89956;
  assign po3009 = n89957 | n89958;
  assign n89960 = ~n88957 & ~n88991;
  assign n89961 = n88930 & ~n89960;
  assign n89962 = ~n88996 & ~n89313;
  assign n89963 = ~n88966 & n89962;
  assign n89964 = ~n88973 & ~n89963;
  assign n89965 = n88930 & n89964;
  assign n89966 = ~n89961 & ~n89965;
  assign n89967 = n88956 & n89316;
  assign n89968 = ~n89318 & ~n89967;
  assign n89969 = ~n88999 & ~n89342;
  assign n89970 = n88973 & ~n89969;
  assign n89971 = n88930 & n89970;
  assign n89972 = n89968 & ~n89971;
  assign n89973 = ~n88997 & ~n89321;
  assign n89974 = n88936 & n88961;
  assign n89975 = ~n89308 & ~n89974;
  assign n89976 = n88973 & ~n89975;
  assign n89977 = n88936 & n88956;
  assign n89978 = n88936 & n88955;
  assign n89979 = ~n89021 & ~n89978;
  assign n89980 = ~n88973 & ~n89979;
  assign n89981 = ~n89977 & ~n89980;
  assign n89982 = ~n89976 & n89981;
  assign n89983 = n89973 & n89982;
  assign n89984 = ~n88930 & ~n89983;
  assign n89985 = ~n89339 & n89612;
  assign n89986 = n88973 & ~n89985;
  assign n89987 = ~n89984 & ~n89986;
  assign n89988 = n89972 & n89987;
  assign n89989 = n89966 & n89988;
  assign n89990 = ~pi2877 & ~n89989;
  assign n89991 = pi2877 & n89972;
  assign n89992 = n89966 & n89991;
  assign n89993 = n89987 & n89992;
  assign po3010 = n89990 | n89993;
  assign n89995 = ~n89378 & n89404;
  assign n89996 = ~n89803 & ~n89995;
  assign n89997 = ~n89417 & ~n89793;
  assign n89998 = ~n89359 & ~n89997;
  assign n89999 = n89378 & n89409;
  assign n90000 = ~n89782 & ~n89999;
  assign n90001 = n89359 & ~n90000;
  assign n90002 = ~n89998 & ~n90001;
  assign n90003 = ~n89386 & n90002;
  assign n90004 = n89996 & n90003;
  assign n90005 = ~n89777 & ~n89789;
  assign n90006 = n90004 & n90005;
  assign n90007 = n89396 & ~n90006;
  assign n90008 = n89372 & n89778;
  assign n90009 = n89426 & ~n90008;
  assign n90010 = n89359 & ~n90009;
  assign n90011 = ~n89378 & n89414;
  assign n90012 = ~n90010 & ~n90011;
  assign n90013 = n89365 & n89387;
  assign n90014 = n89378 & n89400;
  assign n90015 = ~n90013 & ~n90014;
  assign n90016 = n89359 & ~n90015;
  assign n90017 = n89359 & n89409;
  assign n90018 = ~n89378 & n90017;
  assign n90019 = ~n90016 & ~n90018;
  assign n90020 = n90012 & n90019;
  assign n90021 = ~n89396 & ~n90020;
  assign n90022 = ~n89404 & ~n89411;
  assign n90023 = ~n89783 & n90022;
  assign n90024 = n89431 & ~n90023;
  assign n90025 = ~n90021 & ~n90024;
  assign n90026 = ~n89386 & ~n89777;
  assign n90027 = ~n89359 & ~n90026;
  assign n90028 = n90025 & ~n90027;
  assign n90029 = ~n90007 & n90028;
  assign n90030 = ~pi2867 & n90029;
  assign n90031 = pi2867 & ~n90029;
  assign po3011 = n90030 | n90031;
  assign n90033 = ~n88610 & ~n89198;
  assign n90034 = n88527 & ~n90033;
  assign n90035 = ~n88557 & ~n88560;
  assign n90036 = ~n88553 & n88609;
  assign n90037 = ~n89168 & ~n90036;
  assign n90038 = n90035 & n90037;
  assign n90039 = ~n88527 & ~n90038;
  assign n90040 = ~n88592 & n88594;
  assign n90041 = ~n88527 & n90040;
  assign n90042 = n88539 & n89507;
  assign n90043 = ~n89190 & ~n90042;
  assign n90044 = ~n88562 & n90043;
  assign n90045 = n88527 & ~n90044;
  assign n90046 = ~n88533 & n88579;
  assign n90047 = ~n88553 & n90046;
  assign n90048 = ~n90045 & ~n90047;
  assign n90049 = ~n88592 & ~n90048;
  assign n90050 = ~n90041 & ~n90049;
  assign n90051 = ~n88533 & ~n88539;
  assign n90052 = ~n88527 & n90051;
  assign n90053 = n88553 & n90052;
  assign n90054 = ~n88553 & n89190;
  assign n90055 = ~n88560 & ~n90054;
  assign n90056 = ~n89195 & n90055;
  assign n90057 = ~n90053 & n90056;
  assign n90058 = n88527 & n88556;
  assign n90059 = n90057 & ~n90058;
  assign n90060 = n88592 & ~n90059;
  assign n90061 = n90050 & ~n90060;
  assign n90062 = ~n90039 & n90061;
  assign n90063 = ~n90034 & n90062;
  assign n90064 = pi2898 & n90063;
  assign n90065 = ~pi2898 & ~n90063;
  assign po3012 = n90064 | n90065;
  assign n90067 = ~n89378 & n89400;
  assign n90068 = ~n89399 & ~n90067;
  assign n90069 = ~n89359 & ~n90068;
  assign n90070 = n89359 & ~n89805;
  assign n90071 = ~n89794 & ~n90070;
  assign n90072 = ~n90069 & n90071;
  assign n90073 = n89396 & ~n90072;
  assign n90074 = ~n89359 & n89414;
  assign n90075 = ~n90073 & ~n90074;
  assign n90076 = ~n89995 & ~n90014;
  assign n90077 = n89359 & ~n90076;
  assign n90078 = n89359 & n89401;
  assign n90079 = n89378 & n89417;
  assign n90080 = ~n89384 & n89770;
  assign n90081 = ~n89781 & ~n90080;
  assign n90082 = ~n89365 & ~n90081;
  assign n90083 = ~n89782 & ~n90082;
  assign n90084 = ~n89386 & n90083;
  assign n90085 = ~n90079 & n90084;
  assign n90086 = ~n90078 & n90085;
  assign n90087 = ~n89396 & ~n90086;
  assign n90088 = ~n90077 & ~n90087;
  assign n90089 = n90075 & n90088;
  assign n90090 = pi2889 & ~n90089;
  assign n90091 = ~pi2889 & n90089;
  assign po3013 = n90090 | n90091;
  assign n90093 = pi6663 & pi9040;
  assign n90094 = pi6811 & ~pi9040;
  assign n90095 = ~n90093 & ~n90094;
  assign n90096 = ~pi2901 & ~n90095;
  assign n90097 = pi2901 & n90095;
  assign n90098 = ~n90096 & ~n90097;
  assign n90099 = pi6671 & pi9040;
  assign n90100 = pi6732 & ~pi9040;
  assign n90101 = ~n90099 & ~n90100;
  assign n90102 = ~pi2911 & n90101;
  assign n90103 = pi2911 & ~n90101;
  assign n90104 = ~n90102 & ~n90103;
  assign n90105 = pi6806 & ~pi9040;
  assign n90106 = pi6684 & pi9040;
  assign n90107 = ~n90105 & ~n90106;
  assign n90108 = ~pi2908 & ~n90107;
  assign n90109 = pi2908 & n90107;
  assign n90110 = ~n90108 & ~n90109;
  assign n90111 = pi6668 & pi9040;
  assign n90112 = pi6794 & ~pi9040;
  assign n90113 = ~n90111 & ~n90112;
  assign n90114 = ~pi2881 & ~n90113;
  assign n90115 = pi2881 & n90113;
  assign n90116 = ~n90114 & ~n90115;
  assign n90117 = pi6676 & pi9040;
  assign n90118 = pi6839 & ~pi9040;
  assign n90119 = ~n90117 & ~n90118;
  assign n90120 = ~pi2905 & ~n90119;
  assign n90121 = pi2905 & n90119;
  assign n90122 = ~n90120 & ~n90121;
  assign n90123 = n90116 & ~n90122;
  assign n90124 = n90110 & n90123;
  assign n90125 = ~n90104 & n90124;
  assign n90126 = n90104 & n90116;
  assign n90127 = n90122 & n90126;
  assign n90128 = pi6737 & pi9040;
  assign n90129 = pi6655 & ~pi9040;
  assign n90130 = ~n90128 & ~n90129;
  assign n90131 = ~pi2900 & n90130;
  assign n90132 = pi2900 & ~n90130;
  assign n90133 = ~n90131 & ~n90132;
  assign n90134 = ~n90110 & n90126;
  assign n90135 = n90110 & n90122;
  assign n90136 = ~n90116 & n90135;
  assign n90137 = ~n90134 & ~n90136;
  assign n90138 = n90133 & ~n90137;
  assign n90139 = ~n90127 & ~n90138;
  assign n90140 = n90116 & n90135;
  assign n90141 = ~n90110 & ~n90116;
  assign n90142 = ~n90116 & ~n90122;
  assign n90143 = n90104 & n90142;
  assign n90144 = ~n90110 & ~n90122;
  assign n90145 = ~n90104 & n90144;
  assign n90146 = ~n90143 & ~n90145;
  assign n90147 = ~n90141 & n90146;
  assign n90148 = ~n90140 & n90147;
  assign n90149 = ~n90133 & ~n90148;
  assign n90150 = n90139 & ~n90149;
  assign n90151 = ~n90125 & n90150;
  assign n90152 = n90098 & ~n90151;
  assign n90153 = ~n90110 & n90122;
  assign n90154 = ~n90116 & n90153;
  assign n90155 = n90104 & n90154;
  assign n90156 = ~n90104 & ~n90116;
  assign n90157 = ~n90122 & n90156;
  assign n90158 = ~n90110 & n90157;
  assign n90159 = ~n90125 & ~n90158;
  assign n90160 = ~n90155 & n90159;
  assign n90161 = ~n90133 & ~n90160;
  assign n90162 = ~n90152 & ~n90161;
  assign n90163 = n90104 & n90140;
  assign n90164 = n90110 & ~n90116;
  assign n90165 = n90133 & n90164;
  assign n90166 = ~n90104 & n90165;
  assign n90167 = n90116 & n90153;
  assign n90168 = ~n90104 & n90167;
  assign n90169 = n90123 & ~n90133;
  assign n90170 = n90104 & n90169;
  assign n90171 = ~n90168 & ~n90170;
  assign n90172 = ~n90110 & n90116;
  assign n90173 = ~n90104 & n90172;
  assign n90174 = n90110 & ~n90122;
  assign n90175 = ~n90116 & n90174;
  assign n90176 = ~n90173 & ~n90175;
  assign n90177 = n90133 & ~n90176;
  assign n90178 = n90133 & n90141;
  assign n90179 = n90104 & n90178;
  assign n90180 = ~n90177 & ~n90179;
  assign n90181 = n90171 & n90180;
  assign n90182 = ~n90098 & ~n90181;
  assign n90183 = ~n90166 & ~n90182;
  assign n90184 = ~n90163 & n90183;
  assign n90185 = n90162 & n90184;
  assign n90186 = ~pi2921 & ~n90185;
  assign n90187 = ~n90152 & ~n90163;
  assign n90188 = ~n90161 & n90187;
  assign n90189 = n90183 & n90188;
  assign n90190 = pi2921 & n90189;
  assign po3032 = n90186 | n90190;
  assign n90192 = n90104 & n90133;
  assign n90193 = n90110 & n90192;
  assign n90194 = n90116 & n90144;
  assign n90195 = ~n90104 & n90194;
  assign n90196 = ~n90104 & n90154;
  assign n90197 = ~n90195 & ~n90196;
  assign n90198 = n90104 & ~n90116;
  assign n90199 = ~n90122 & n90198;
  assign n90200 = ~n90110 & n90199;
  assign n90201 = ~n90136 & ~n90200;
  assign n90202 = ~n90133 & ~n90201;
  assign n90203 = n90197 & ~n90202;
  assign n90204 = ~n90193 & n90203;
  assign n90205 = n90098 & ~n90204;
  assign n90206 = ~n90104 & n90175;
  assign n90207 = n90133 & n90206;
  assign n90208 = n90104 & ~n90133;
  assign n90209 = n90175 & n90208;
  assign n90210 = ~n90134 & ~n90209;
  assign n90211 = ~n90136 & ~n90167;
  assign n90212 = n90104 & n90153;
  assign n90213 = n90211 & ~n90212;
  assign n90214 = n90133 & ~n90213;
  assign n90215 = ~n90133 & n90140;
  assign n90216 = n90159 & ~n90215;
  assign n90217 = ~n90214 & n90216;
  assign n90218 = n90210 & n90217;
  assign n90219 = ~n90098 & ~n90218;
  assign n90220 = ~n90207 & ~n90219;
  assign n90221 = ~n90205 & n90220;
  assign n90222 = n90167 & n90208;
  assign n90223 = ~n90104 & n90169;
  assign n90224 = ~n90222 & ~n90223;
  assign n90225 = ~n90133 & n90196;
  assign n90226 = n90224 & ~n90225;
  assign n90227 = n90221 & n90226;
  assign n90228 = ~pi2926 & ~n90227;
  assign n90229 = pi2926 & n90226;
  assign n90230 = n90220 & n90229;
  assign n90231 = ~n90205 & n90230;
  assign po3042 = n90228 | n90231;
  assign n90233 = pi6738 & pi9040;
  assign n90234 = pi6765 & ~pi9040;
  assign n90235 = ~n90233 & ~n90234;
  assign n90236 = ~pi2903 & ~n90235;
  assign n90237 = pi2903 & n90235;
  assign n90238 = ~n90236 & ~n90237;
  assign n90239 = pi6987 & pi9040;
  assign n90240 = pi6736 & ~pi9040;
  assign n90241 = ~n90239 & ~n90240;
  assign n90242 = ~pi2897 & ~n90241;
  assign n90243 = pi2897 & n90241;
  assign n90244 = ~n90242 & ~n90243;
  assign n90245 = pi6667 & pi9040;
  assign n90246 = pi6809 & ~pi9040;
  assign n90247 = ~n90245 & ~n90246;
  assign n90248 = ~pi2895 & n90247;
  assign n90249 = pi2895 & ~n90247;
  assign n90250 = ~n90248 & ~n90249;
  assign n90251 = ~n90244 & n90250;
  assign n90252 = ~n90238 & n90251;
  assign n90253 = pi6727 & pi9040;
  assign n90254 = pi6722 & ~pi9040;
  assign n90255 = ~n90253 & ~n90254;
  assign n90256 = pi2872 & n90255;
  assign n90257 = ~pi2872 & ~n90255;
  assign n90258 = ~n90256 & ~n90257;
  assign n90259 = ~n90244 & ~n90250;
  assign n90260 = n90258 & n90259;
  assign n90261 = ~n90252 & ~n90260;
  assign n90262 = pi6674 & ~pi9040;
  assign n90263 = pi6765 & pi9040;
  assign n90264 = ~n90262 & ~n90263;
  assign n90265 = pi2878 & n90264;
  assign n90266 = ~pi2878 & ~n90264;
  assign n90267 = ~n90265 & ~n90266;
  assign n90268 = pi6735 & pi9040;
  assign n90269 = pi6766 & ~pi9040;
  assign n90270 = ~n90268 & ~n90269;
  assign n90271 = ~pi2890 & ~n90270;
  assign n90272 = pi2890 & n90270;
  assign n90273 = ~n90271 & ~n90272;
  assign n90274 = n90267 & ~n90273;
  assign n90275 = ~n90261 & n90274;
  assign n90276 = n90244 & n90250;
  assign n90277 = n90238 & n90258;
  assign n90278 = n90276 & n90277;
  assign n90279 = n90244 & ~n90250;
  assign n90280 = ~n90258 & n90279;
  assign n90281 = n90251 & ~n90258;
  assign n90282 = ~n90280 & ~n90281;
  assign n90283 = n90238 & ~n90282;
  assign n90284 = ~n90278 & ~n90283;
  assign n90285 = ~n90273 & ~n90284;
  assign n90286 = ~n90275 & ~n90285;
  assign n90287 = n90238 & ~n90258;
  assign n90288 = ~n90244 & n90287;
  assign n90289 = ~n90278 & ~n90288;
  assign n90290 = ~n90267 & ~n90289;
  assign n90291 = ~n90238 & n90267;
  assign n90292 = n90244 & n90291;
  assign n90293 = ~n90258 & n90276;
  assign n90294 = n90258 & n90279;
  assign n90295 = ~n90293 & ~n90294;
  assign n90296 = n90251 & n90258;
  assign n90297 = n90238 & n90296;
  assign n90298 = n90295 & ~n90297;
  assign n90299 = n90267 & ~n90298;
  assign n90300 = ~n90292 & ~n90299;
  assign n90301 = ~n90258 & n90259;
  assign n90302 = n90238 & n90301;
  assign n90303 = n90300 & ~n90302;
  assign n90304 = ~n90261 & ~n90267;
  assign n90305 = ~n90238 & n90280;
  assign n90306 = ~n90304 & ~n90305;
  assign n90307 = n90303 & n90306;
  assign n90308 = n90273 & ~n90307;
  assign n90309 = ~n90290 & ~n90308;
  assign n90310 = ~n90267 & ~n90273;
  assign n90311 = ~n90238 & n90276;
  assign n90312 = ~n90301 & ~n90311;
  assign n90313 = n90244 & n90258;
  assign n90314 = n90312 & ~n90313;
  assign n90315 = n90310 & ~n90314;
  assign n90316 = n90309 & ~n90315;
  assign n90317 = n90286 & n90316;
  assign n90318 = ~pi2918 & ~n90317;
  assign n90319 = pi2918 & n90286;
  assign n90320 = n90309 & n90319;
  assign n90321 = ~n90315 & n90320;
  assign po3043 = n90318 | n90321;
  assign n90323 = pi6807 & pi9040;
  assign n90324 = pi6721 & ~pi9040;
  assign n90325 = ~n90323 & ~n90324;
  assign n90326 = ~pi2908 & ~n90325;
  assign n90327 = pi2908 & n90325;
  assign n90328 = ~n90326 & ~n90327;
  assign n90329 = pi6661 & ~pi9040;
  assign n90330 = pi6634 & pi9040;
  assign n90331 = ~n90329 & ~n90330;
  assign n90332 = ~pi2886 & n90331;
  assign n90333 = pi2886 & ~n90331;
  assign n90334 = ~n90332 & ~n90333;
  assign n90335 = pi6730 & ~pi9040;
  assign n90336 = pi6896 & pi9040;
  assign n90337 = ~n90335 & ~n90336;
  assign n90338 = ~pi2899 & ~n90337;
  assign n90339 = pi2899 & n90337;
  assign n90340 = ~n90338 & ~n90339;
  assign n90341 = pi6774 & pi9040;
  assign n90342 = pi6896 & ~pi9040;
  assign n90343 = ~n90341 & ~n90342;
  assign n90344 = ~pi2880 & n90343;
  assign n90345 = pi2880 & ~n90343;
  assign n90346 = ~n90344 & ~n90345;
  assign n90347 = pi6632 & pi9040;
  assign n90348 = pi6735 & ~pi9040;
  assign n90349 = ~n90347 & ~n90348;
  assign n90350 = ~pi2881 & ~n90349;
  assign n90351 = pi2881 & n90349;
  assign n90352 = ~n90350 & ~n90351;
  assign n90353 = n90346 & n90352;
  assign n90354 = n90340 & n90353;
  assign n90355 = ~n90334 & n90354;
  assign n90356 = pi6658 & pi9040;
  assign n90357 = pi6853 & ~pi9040;
  assign n90358 = ~n90356 & ~n90357;
  assign n90359 = ~pi2909 & ~n90358;
  assign n90360 = pi2909 & n90358;
  assign n90361 = ~n90359 & ~n90360;
  assign n90362 = ~n90346 & n90352;
  assign n90363 = ~n90334 & n90362;
  assign n90364 = ~n90340 & n90353;
  assign n90365 = n90334 & n90364;
  assign n90366 = ~n90363 & ~n90365;
  assign n90367 = ~n90361 & ~n90366;
  assign n90368 = ~n90355 & ~n90367;
  assign n90369 = n90346 & ~n90352;
  assign n90370 = ~n90340 & n90369;
  assign n90371 = n90361 & n90370;
  assign n90372 = n90353 & n90361;
  assign n90373 = ~n90334 & n90372;
  assign n90374 = ~n90371 & ~n90373;
  assign n90375 = n90368 & n90374;
  assign n90376 = ~n90346 & ~n90352;
  assign n90377 = n90340 & n90376;
  assign n90378 = ~n90334 & n90377;
  assign n90379 = n90340 & n90369;
  assign n90380 = n90334 & n90379;
  assign n90381 = ~n90378 & ~n90380;
  assign n90382 = n90375 & n90381;
  assign n90383 = n90328 & ~n90382;
  assign n90384 = ~n90328 & ~n90361;
  assign n90385 = ~n90334 & ~n90340;
  assign n90386 = n90346 & n90385;
  assign n90387 = ~n90340 & ~n90352;
  assign n90388 = ~n90386 & ~n90387;
  assign n90389 = n90384 & ~n90388;
  assign n90390 = n90334 & n90340;
  assign n90391 = n90352 & n90390;
  assign n90392 = n90346 & n90391;
  assign n90393 = n90361 & n90392;
  assign n90394 = ~n90340 & n90376;
  assign n90395 = ~n90361 & n90394;
  assign n90396 = n90334 & n90395;
  assign n90397 = ~n90393 & ~n90396;
  assign n90398 = n90340 & n90362;
  assign n90399 = n90334 & n90398;
  assign n90400 = ~n90380 & ~n90399;
  assign n90401 = ~n90361 & ~n90400;
  assign n90402 = n90334 & ~n90346;
  assign n90403 = ~n90340 & n90402;
  assign n90404 = ~n90392 & ~n90403;
  assign n90405 = ~n90334 & n90361;
  assign n90406 = n90340 & n90405;
  assign n90407 = ~n90353 & n90406;
  assign n90408 = n90361 & n90377;
  assign n90409 = ~n90407 & ~n90408;
  assign n90410 = n90404 & n90409;
  assign n90411 = ~n90328 & ~n90410;
  assign n90412 = ~n90401 & ~n90411;
  assign n90413 = n90397 & n90412;
  assign n90414 = ~n90389 & n90413;
  assign n90415 = ~n90383 & n90414;
  assign n90416 = ~n90340 & n90362;
  assign n90417 = n90334 & n90361;
  assign n90418 = n90416 & n90417;
  assign n90419 = n90415 & ~n90418;
  assign n90420 = ~pi2929 & ~n90419;
  assign n90421 = pi2929 & ~n90418;
  assign n90422 = n90414 & n90421;
  assign n90423 = ~n90383 & n90422;
  assign po3047 = n90420 | n90423;
  assign n90425 = n90334 & ~n90340;
  assign n90426 = ~n90352 & n90425;
  assign n90427 = n90346 & n90426;
  assign n90428 = ~n90334 & n90394;
  assign n90429 = ~n90427 & ~n90428;
  assign n90430 = n90361 & ~n90429;
  assign n90431 = ~n90361 & n90392;
  assign n90432 = ~n90392 & ~n90408;
  assign n90433 = n90346 & n90390;
  assign n90434 = ~n90403 & ~n90433;
  assign n90435 = ~n90361 & ~n90434;
  assign n90436 = ~n90334 & ~n90361;
  assign n90437 = n90369 & n90436;
  assign n90438 = ~n90340 & n90437;
  assign n90439 = ~n90340 & n90361;
  assign n90440 = n90352 & n90439;
  assign n90441 = n90346 & n90440;
  assign n90442 = ~n90334 & n90340;
  assign n90443 = n90352 & n90442;
  assign n90444 = ~n90346 & n90443;
  assign n90445 = ~n90441 & ~n90444;
  assign n90446 = ~n90438 & n90445;
  assign n90447 = ~n90435 & n90446;
  assign n90448 = n90432 & n90447;
  assign n90449 = n90328 & ~n90448;
  assign n90450 = n90334 & n90408;
  assign n90451 = ~n90449 & ~n90450;
  assign n90452 = ~n90431 & n90451;
  assign n90453 = ~n90430 & n90452;
  assign n90454 = n90340 & n90346;
  assign n90455 = n90405 & n90454;
  assign n90456 = ~n90371 & ~n90455;
  assign n90457 = n90361 & n90398;
  assign n90458 = n90334 & n90416;
  assign n90459 = ~n90457 & ~n90458;
  assign n90460 = ~n90334 & n90376;
  assign n90461 = ~n90340 & n90352;
  assign n90462 = ~n90460 & ~n90461;
  assign n90463 = ~n90361 & ~n90462;
  assign n90464 = ~n90334 & n90379;
  assign n90465 = ~n90427 & ~n90464;
  assign n90466 = ~n90463 & n90465;
  assign n90467 = n90459 & n90466;
  assign n90468 = n90456 & n90467;
  assign n90469 = ~n90328 & ~n90468;
  assign n90470 = n90453 & ~n90469;
  assign n90471 = ~pi2923 & ~n90470;
  assign n90472 = pi2923 & n90453;
  assign n90473 = ~n90469 & n90472;
  assign po3048 = n90471 | n90473;
  assign n90475 = pi6668 & ~pi9040;
  assign n90476 = pi6672 & pi9040;
  assign n90477 = ~n90475 & ~n90476;
  assign n90478 = ~pi2904 & ~n90477;
  assign n90479 = pi2904 & n90477;
  assign n90480 = ~n90478 & ~n90479;
  assign n90481 = pi6769 & ~pi9040;
  assign n90482 = pi6660 & pi9040;
  assign n90483 = ~n90481 & ~n90482;
  assign n90484 = pi2894 & ~n90483;
  assign n90485 = ~pi2894 & n90483;
  assign n90486 = ~n90484 & ~n90485;
  assign n90487 = pi6726 & pi9040;
  assign n90488 = pi6670 & ~pi9040;
  assign n90489 = ~n90487 & ~n90488;
  assign n90490 = ~pi2868 & ~n90489;
  assign n90491 = pi2868 & n90489;
  assign n90492 = ~n90490 & ~n90491;
  assign n90493 = pi6801 & ~pi9040;
  assign n90494 = pi6739 & pi9040;
  assign n90495 = ~n90493 & ~n90494;
  assign n90496 = ~pi2879 & n90495;
  assign n90497 = pi2879 & ~n90495;
  assign n90498 = ~n90496 & ~n90497;
  assign n90499 = pi6671 & ~pi9040;
  assign n90500 = pi6662 & pi9040;
  assign n90501 = ~n90499 & ~n90500;
  assign n90502 = ~pi2905 & ~n90501;
  assign n90503 = pi2905 & n90501;
  assign n90504 = ~n90502 & ~n90503;
  assign n90505 = pi6828 & pi9040;
  assign n90506 = pi6699 & ~pi9040;
  assign n90507 = ~n90505 & ~n90506;
  assign n90508 = ~pi2901 & ~n90507;
  assign n90509 = pi2901 & n90507;
  assign n90510 = ~n90508 & ~n90509;
  assign n90511 = ~n90504 & n90510;
  assign n90512 = ~n90498 & n90511;
  assign n90513 = ~n90492 & n90512;
  assign n90514 = ~n90498 & ~n90510;
  assign n90515 = n90504 & n90514;
  assign n90516 = ~n90492 & ~n90515;
  assign n90517 = n90498 & n90510;
  assign n90518 = ~n90504 & ~n90510;
  assign n90519 = ~n90517 & ~n90518;
  assign n90520 = n90492 & n90519;
  assign n90521 = ~n90516 & ~n90520;
  assign n90522 = ~n90513 & ~n90521;
  assign n90523 = n90486 & ~n90522;
  assign n90524 = n90504 & ~n90510;
  assign n90525 = n90492 & n90524;
  assign n90526 = ~n90498 & n90510;
  assign n90527 = n90504 & n90526;
  assign n90528 = ~n90525 & ~n90527;
  assign n90529 = ~n90492 & ~n90504;
  assign n90530 = n90498 & n90529;
  assign n90531 = n90510 & n90530;
  assign n90532 = n90528 & ~n90531;
  assign n90533 = ~n90486 & ~n90532;
  assign n90534 = ~n90523 & ~n90533;
  assign n90535 = n90480 & ~n90534;
  assign n90536 = ~n90486 & ~n90492;
  assign n90537 = ~n90510 & n90536;
  assign n90538 = n90486 & n90517;
  assign n90539 = ~n90492 & n90538;
  assign n90540 = ~n90492 & n90510;
  assign n90541 = n90504 & n90540;
  assign n90542 = ~n90525 & ~n90541;
  assign n90543 = n90486 & ~n90542;
  assign n90544 = ~n90539 & ~n90543;
  assign n90545 = n90504 & n90517;
  assign n90546 = ~n90492 & n90545;
  assign n90547 = n90492 & n90512;
  assign n90548 = ~n90546 & ~n90547;
  assign n90549 = ~n90486 & n90492;
  assign n90550 = n90511 & n90549;
  assign n90551 = ~n90486 & ~n90504;
  assign n90552 = ~n90498 & n90551;
  assign n90553 = ~n90510 & n90552;
  assign n90554 = ~n90550 & ~n90553;
  assign n90555 = n90548 & n90554;
  assign n90556 = n90544 & n90555;
  assign n90557 = ~n90537 & n90556;
  assign n90558 = ~n90480 & ~n90557;
  assign n90559 = n90486 & n90546;
  assign n90560 = n90498 & ~n90510;
  assign n90561 = ~n90504 & n90560;
  assign n90562 = n90486 & n90561;
  assign n90563 = ~n90492 & n90562;
  assign n90564 = ~n90559 & ~n90563;
  assign n90565 = ~n90498 & n90518;
  assign n90566 = ~n90492 & n90565;
  assign n90567 = ~n90486 & n90566;
  assign n90568 = n90564 & ~n90567;
  assign n90569 = ~n90492 & n90504;
  assign n90570 = n90498 & n90569;
  assign n90571 = ~n90510 & n90570;
  assign n90572 = n90492 & n90526;
  assign n90573 = ~n90571 & ~n90572;
  assign n90574 = ~n90486 & ~n90573;
  assign n90575 = n90568 & ~n90574;
  assign n90576 = ~n90558 & n90575;
  assign n90577 = ~n90535 & n90576;
  assign n90578 = ~pi2920 & n90577;
  assign n90579 = pi2920 & ~n90577;
  assign po3049 = n90578 | n90579;
  assign n90581 = pi6740 & pi9040;
  assign n90582 = pi6669 & ~pi9040;
  assign n90583 = ~n90581 & ~n90582;
  assign n90584 = ~pi2888 & ~n90583;
  assign n90585 = pi2888 & n90583;
  assign n90586 = ~n90584 & ~n90585;
  assign n90587 = pi6800 & pi9040;
  assign n90588 = pi6734 & ~pi9040;
  assign n90589 = ~n90587 & ~n90588;
  assign n90590 = ~pi2904 & ~n90589;
  assign n90591 = pi2904 & n90589;
  assign n90592 = ~n90590 & ~n90591;
  assign n90593 = pi6669 & pi9040;
  assign n90594 = pi6800 & ~pi9040;
  assign n90595 = ~n90593 & ~n90594;
  assign n90596 = ~pi2887 & n90595;
  assign n90597 = pi2887 & ~n90595;
  assign n90598 = ~n90596 & ~n90597;
  assign n90599 = ~n90592 & ~n90598;
  assign n90600 = pi6801 & pi9040;
  assign n90601 = pi6828 & ~pi9040;
  assign n90602 = ~n90600 & ~n90601;
  assign n90603 = ~pi2885 & ~n90602;
  assign n90604 = pi2885 & n90602;
  assign n90605 = ~n90603 & ~n90604;
  assign n90606 = pi6663 & ~pi9040;
  assign n90607 = pi6655 & pi9040;
  assign n90608 = ~n90606 & ~n90607;
  assign n90609 = pi2902 & n90608;
  assign n90610 = ~pi2902 & ~n90608;
  assign n90611 = ~n90609 & ~n90610;
  assign n90612 = ~n90605 & ~n90611;
  assign n90613 = n90599 & n90612;
  assign n90614 = pi6699 & pi9040;
  assign n90615 = pi6662 & ~pi9040;
  assign n90616 = ~n90614 & ~n90615;
  assign n90617 = ~pi2879 & n90616;
  assign n90618 = pi2879 & ~n90616;
  assign n90619 = ~n90617 & ~n90618;
  assign n90620 = n90592 & n90598;
  assign n90621 = ~n90619 & n90620;
  assign n90622 = n90605 & n90619;
  assign n90623 = n90598 & n90622;
  assign n90624 = ~n90592 & n90623;
  assign n90625 = ~n90621 & ~n90624;
  assign n90626 = n90592 & ~n90598;
  assign n90627 = n90605 & n90626;
  assign n90628 = n90625 & ~n90627;
  assign n90629 = ~n90611 & ~n90628;
  assign n90630 = n90592 & n90619;
  assign n90631 = ~n90605 & n90611;
  assign n90632 = n90630 & n90631;
  assign n90633 = ~n90605 & n90619;
  assign n90634 = n90598 & n90633;
  assign n90635 = n90592 & n90634;
  assign n90636 = ~n90632 & ~n90635;
  assign n90637 = ~n90629 & n90636;
  assign n90638 = ~n90613 & n90637;
  assign n90639 = n90599 & ~n90619;
  assign n90640 = ~n90605 & n90639;
  assign n90641 = ~n90619 & n90626;
  assign n90642 = n90605 & n90641;
  assign n90643 = ~n90640 & ~n90642;
  assign n90644 = n90638 & n90643;
  assign n90645 = ~n90586 & ~n90644;
  assign n90646 = n90619 & n90626;
  assign n90647 = ~n90605 & n90646;
  assign n90648 = ~n90639 & ~n90647;
  assign n90649 = ~n90611 & ~n90648;
  assign n90650 = n90599 & n90622;
  assign n90651 = ~n90592 & n90619;
  assign n90652 = n90598 & n90651;
  assign n90653 = ~n90605 & n90652;
  assign n90654 = ~n90650 & ~n90653;
  assign n90655 = n90592 & n90622;
  assign n90656 = ~n90605 & n90641;
  assign n90657 = ~n90655 & ~n90656;
  assign n90658 = n90611 & ~n90657;
  assign n90659 = n90654 & ~n90658;
  assign n90660 = ~n90649 & n90659;
  assign n90661 = n90586 & ~n90660;
  assign n90662 = n90592 & ~n90619;
  assign n90663 = n90605 & n90662;
  assign n90664 = ~n90592 & ~n90619;
  assign n90665 = ~n90605 & n90664;
  assign n90666 = ~n90663 & ~n90665;
  assign n90667 = ~n90611 & ~n90666;
  assign n90668 = ~n90592 & n90598;
  assign n90669 = ~n90619 & n90668;
  assign n90670 = n90605 & n90669;
  assign n90671 = ~n90650 & ~n90670;
  assign n90672 = n90619 & n90620;
  assign n90673 = n90671 & ~n90672;
  assign n90674 = n90611 & ~n90673;
  assign n90675 = ~n90667 & ~n90674;
  assign n90676 = n90598 & n90619;
  assign n90677 = n90611 & n90676;
  assign n90678 = ~n90605 & n90677;
  assign n90679 = n90675 & ~n90678;
  assign n90680 = ~n90661 & n90679;
  assign n90681 = ~n90645 & n90680;
  assign n90682 = ~pi2914 & ~n90681;
  assign n90683 = pi2914 & n90681;
  assign po3050 = n90682 | n90683;
  assign n90685 = pi6809 & pi9040;
  assign n90686 = pi6658 & ~pi9040;
  assign n90687 = ~n90685 & ~n90686;
  assign n90688 = ~pi2897 & ~n90687;
  assign n90689 = pi2897 & n90687;
  assign n90690 = ~n90688 & ~n90689;
  assign n90691 = pi6763 & pi9040;
  assign n90692 = pi6664 & ~pi9040;
  assign n90693 = ~n90691 & ~n90692;
  assign n90694 = ~pi2907 & ~n90693;
  assign n90695 = pi2907 & n90693;
  assign n90696 = ~n90694 & ~n90695;
  assign n90697 = pi6866 & ~pi9040;
  assign n90698 = pi6731 & pi9040;
  assign n90699 = ~n90697 & ~n90698;
  assign n90700 = ~pi2891 & ~n90699;
  assign n90701 = pi2891 & n90699;
  assign n90702 = ~n90700 & ~n90701;
  assign n90703 = pi6866 & pi9040;
  assign n90704 = pi6673 & ~pi9040;
  assign n90705 = ~n90703 & ~n90704;
  assign n90706 = ~pi2872 & ~n90705;
  assign n90707 = pi2872 & n90705;
  assign n90708 = ~n90706 & ~n90707;
  assign n90709 = ~n90702 & n90708;
  assign n90710 = pi6632 & ~pi9040;
  assign n90711 = pi6853 & pi9040;
  assign n90712 = ~n90710 & ~n90711;
  assign n90713 = ~pi2892 & n90712;
  assign n90714 = pi2892 & ~n90712;
  assign n90715 = ~n90713 & ~n90714;
  assign n90716 = pi6673 & pi9040;
  assign n90717 = pi6738 & ~pi9040;
  assign n90718 = ~n90716 & ~n90717;
  assign n90719 = pi2896 & n90718;
  assign n90720 = ~pi2896 & ~n90718;
  assign n90721 = ~n90719 & ~n90720;
  assign n90722 = ~n90715 & n90721;
  assign n90723 = n90709 & n90722;
  assign n90724 = n90696 & n90723;
  assign n90725 = n90715 & n90721;
  assign n90726 = n90708 & n90725;
  assign n90727 = n90702 & n90726;
  assign n90728 = n90696 & n90715;
  assign n90729 = ~n90708 & n90728;
  assign n90730 = ~n90702 & n90729;
  assign n90731 = n90702 & ~n90708;
  assign n90732 = n90696 & n90731;
  assign n90733 = n90721 & n90732;
  assign n90734 = ~n90715 & n90733;
  assign n90735 = ~n90730 & ~n90734;
  assign n90736 = ~n90727 & n90735;
  assign n90737 = ~n90724 & n90736;
  assign n90738 = n90702 & n90708;
  assign n90739 = ~n90696 & n90715;
  assign n90740 = n90738 & n90739;
  assign n90741 = n90737 & ~n90740;
  assign n90742 = ~n90690 & ~n90741;
  assign n90743 = n90696 & n90702;
  assign n90744 = n90708 & n90743;
  assign n90745 = ~n90715 & n90744;
  assign n90746 = ~n90729 & ~n90745;
  assign n90747 = ~n90696 & n90709;
  assign n90748 = ~n90715 & n90747;
  assign n90749 = n90746 & ~n90748;
  assign n90750 = ~n90721 & ~n90749;
  assign n90751 = ~n90696 & ~n90708;
  assign n90752 = n90702 & n90751;
  assign n90753 = ~n90721 & n90752;
  assign n90754 = ~n90715 & n90753;
  assign n90755 = ~n90702 & n90728;
  assign n90756 = ~n90702 & ~n90708;
  assign n90757 = n90715 & n90756;
  assign n90758 = ~n90755 & ~n90757;
  assign n90759 = ~n90721 & ~n90758;
  assign n90760 = ~n90754 & ~n90759;
  assign n90761 = ~n90690 & ~n90760;
  assign n90762 = ~n90750 & ~n90761;
  assign n90763 = ~n90742 & n90762;
  assign n90764 = ~n90696 & ~n90715;
  assign n90765 = n90721 & n90764;
  assign n90766 = n90756 & n90765;
  assign n90767 = ~n90696 & n90702;
  assign n90768 = n90725 & n90767;
  assign n90769 = n90715 & n90752;
  assign n90770 = n90696 & ~n90721;
  assign n90771 = n90702 & n90770;
  assign n90772 = ~n90702 & ~n90715;
  assign n90773 = ~n90696 & n90772;
  assign n90774 = ~n90771 & ~n90773;
  assign n90775 = ~n90769 & n90774;
  assign n90776 = ~n90747 & n90775;
  assign n90777 = n90709 & n90721;
  assign n90778 = n90715 & n90777;
  assign n90779 = ~n90715 & n90756;
  assign n90780 = ~n90696 & n90708;
  assign n90781 = ~n90779 & ~n90780;
  assign n90782 = n90721 & ~n90781;
  assign n90783 = ~n90778 & ~n90782;
  assign n90784 = n90776 & n90783;
  assign n90785 = n90690 & ~n90784;
  assign n90786 = ~n90768 & ~n90785;
  assign n90787 = ~n90766 & n90786;
  assign n90788 = n90763 & n90787;
  assign n90789 = pi2924 & n90788;
  assign n90790 = ~pi2924 & ~n90788;
  assign po3051 = n90789 | n90790;
  assign n90792 = pi6676 & ~pi9040;
  assign n90793 = pi6769 & pi9040;
  assign n90794 = ~n90792 & ~n90793;
  assign n90795 = ~pi2882 & n90794;
  assign n90796 = pi2882 & ~n90794;
  assign n90797 = ~n90795 & ~n90796;
  assign n90798 = pi6672 & ~pi9040;
  assign n90799 = pi6670 & pi9040;
  assign n90800 = ~n90798 & ~n90799;
  assign n90801 = ~pi2887 & n90800;
  assign n90802 = pi2887 & ~n90800;
  assign n90803 = ~n90801 & ~n90802;
  assign n90804 = pi6806 & pi9040;
  assign n90805 = pi6726 & ~pi9040;
  assign n90806 = ~n90804 & ~n90805;
  assign n90807 = ~pi2907 & n90806;
  assign n90808 = pi2907 & ~n90806;
  assign n90809 = ~n90807 & ~n90808;
  assign n90810 = pi6737 & ~pi9040;
  assign n90811 = pi6839 & pi9040;
  assign n90812 = ~n90810 & ~n90811;
  assign n90813 = ~pi2888 & n90812;
  assign n90814 = pi2888 & ~n90812;
  assign n90815 = ~n90813 & ~n90814;
  assign n90816 = ~n90809 & ~n90815;
  assign n90817 = n90803 & n90816;
  assign n90818 = pi6732 & pi9040;
  assign n90819 = pi6684 & ~pi9040;
  assign n90820 = ~n90818 & ~n90819;
  assign n90821 = pi2910 & n90820;
  assign n90822 = ~pi2910 & ~n90820;
  assign n90823 = ~n90821 & ~n90822;
  assign n90824 = n90817 & ~n90823;
  assign n90825 = n90809 & n90815;
  assign n90826 = n90803 & n90825;
  assign n90827 = ~n90823 & n90826;
  assign n90828 = ~n90824 & ~n90827;
  assign n90829 = ~n90803 & n90825;
  assign n90830 = n90823 & n90829;
  assign n90831 = ~n90809 & n90815;
  assign n90832 = n90803 & n90831;
  assign n90833 = n90823 & n90832;
  assign n90834 = ~n90830 & ~n90833;
  assign n90835 = n90828 & n90834;
  assign n90836 = ~n90797 & ~n90835;
  assign n90837 = n90809 & ~n90815;
  assign n90838 = n90803 & n90837;
  assign n90839 = n90823 & n90838;
  assign n90840 = ~n90832 & ~n90839;
  assign n90841 = ~n90797 & ~n90840;
  assign n90842 = n90797 & ~n90815;
  assign n90843 = ~n90823 & n90842;
  assign n90844 = ~n90803 & ~n90809;
  assign n90845 = n90823 & n90825;
  assign n90846 = ~n90844 & ~n90845;
  assign n90847 = n90797 & ~n90846;
  assign n90848 = ~n90843 & ~n90847;
  assign n90849 = ~n90803 & ~n90823;
  assign n90850 = n90837 & n90849;
  assign n90851 = n90848 & ~n90850;
  assign n90852 = ~n90815 & n90844;
  assign n90853 = n90823 & n90852;
  assign n90854 = n90851 & ~n90853;
  assign n90855 = ~n90841 & n90854;
  assign n90856 = pi6739 & ~pi9040;
  assign n90857 = pi6706 & pi9040;
  assign n90858 = ~n90856 & ~n90857;
  assign n90859 = ~pi2891 & ~n90858;
  assign n90860 = pi2891 & n90858;
  assign n90861 = ~n90859 & ~n90860;
  assign n90862 = ~n90855 & ~n90861;
  assign n90863 = n90803 & ~n90815;
  assign n90864 = n90797 & n90823;
  assign n90865 = n90861 & n90864;
  assign n90866 = n90863 & n90865;
  assign n90867 = n90803 & ~n90823;
  assign n90868 = n90815 & n90867;
  assign n90869 = n90797 & ~n90868;
  assign n90870 = ~n90803 & n90823;
  assign n90871 = n90809 & n90870;
  assign n90872 = ~n90816 & ~n90863;
  assign n90873 = ~n90823 & ~n90872;
  assign n90874 = ~n90797 & ~n90829;
  assign n90875 = ~n90873 & n90874;
  assign n90876 = ~n90871 & n90875;
  assign n90877 = ~n90869 & ~n90876;
  assign n90878 = n90815 & n90870;
  assign n90879 = ~n90809 & n90878;
  assign n90880 = ~n90877 & ~n90879;
  assign n90881 = n90861 & ~n90880;
  assign n90882 = ~n90866 & ~n90881;
  assign n90883 = ~n90862 & n90882;
  assign n90884 = ~n90836 & n90883;
  assign n90885 = n90797 & n90850;
  assign n90886 = n90884 & ~n90885;
  assign n90887 = pi2912 & ~n90886;
  assign n90888 = ~pi2912 & ~n90885;
  assign n90889 = n90883 & n90888;
  assign n90890 = ~n90836 & n90889;
  assign po3052 = n90887 | n90890;
  assign n90892 = n90238 & ~n90267;
  assign n90893 = ~n90251 & ~n90280;
  assign n90894 = n90892 & ~n90893;
  assign n90895 = ~n90258 & ~n90267;
  assign n90896 = n90251 & n90895;
  assign n90897 = ~n90894 & ~n90896;
  assign n90898 = n90273 & ~n90897;
  assign n90899 = ~n90238 & n90258;
  assign n90900 = ~n90250 & n90899;
  assign n90901 = n90244 & n90900;
  assign n90902 = ~n90313 & ~n90899;
  assign n90903 = n90267 & ~n90902;
  assign n90904 = ~n90238 & ~n90258;
  assign n90905 = n90250 & n90904;
  assign n90906 = n90244 & n90905;
  assign n90907 = ~n90903 & ~n90906;
  assign n90908 = ~n90901 & n90907;
  assign n90909 = n90273 & ~n90908;
  assign n90910 = ~n90898 & ~n90909;
  assign n90911 = ~n90244 & n90258;
  assign n90912 = ~n90250 & n90911;
  assign n90913 = n90238 & n90912;
  assign n90914 = ~n90238 & n90301;
  assign n90915 = ~n90913 & ~n90914;
  assign n90916 = ~n90267 & ~n90915;
  assign n90917 = n90238 & n90281;
  assign n90918 = ~n90238 & n90313;
  assign n90919 = ~n90917 & ~n90918;
  assign n90920 = n90267 & ~n90919;
  assign n90921 = ~n90276 & ~n90313;
  assign n90922 = n90238 & ~n90921;
  assign n90923 = ~n90301 & ~n90922;
  assign n90924 = ~n90267 & ~n90923;
  assign n90925 = ~n90238 & ~n90250;
  assign n90926 = n90895 & n90925;
  assign n90927 = n90250 & n90258;
  assign n90928 = ~n90301 & ~n90927;
  assign n90929 = ~n90238 & ~n90928;
  assign n90930 = n90238 & n90267;
  assign n90931 = n90279 & n90930;
  assign n90932 = ~n90258 & n90931;
  assign n90933 = ~n90929 & ~n90932;
  assign n90934 = ~n90926 & n90933;
  assign n90935 = ~n90924 & n90934;
  assign n90936 = ~n90913 & n90935;
  assign n90937 = ~n90273 & ~n90936;
  assign n90938 = ~n90920 & ~n90937;
  assign n90939 = ~n90916 & n90938;
  assign n90940 = n90910 & n90939;
  assign n90941 = pi2934 & n90940;
  assign n90942 = ~pi2934 & ~n90940;
  assign po3053 = n90941 | n90942;
  assign n90944 = n90250 & n90287;
  assign n90945 = ~n90280 & ~n90944;
  assign n90946 = ~n90267 & ~n90945;
  assign n90947 = n90238 & n90259;
  assign n90948 = ~n90238 & n90250;
  assign n90949 = ~n90258 & n90948;
  assign n90950 = ~n90947 & ~n90949;
  assign n90951 = n90267 & ~n90950;
  assign n90952 = ~n90238 & n90296;
  assign n90953 = ~n90926 & ~n90952;
  assign n90954 = ~n90278 & n90953;
  assign n90955 = ~n90951 & n90954;
  assign n90956 = ~n90946 & n90955;
  assign n90957 = ~n90901 & ~n90913;
  assign n90958 = n90956 & n90957;
  assign n90959 = n90273 & ~n90958;
  assign n90960 = n90276 & n90899;
  assign n90961 = n90282 & ~n90960;
  assign n90962 = n90267 & ~n90961;
  assign n90963 = ~n90238 & n90260;
  assign n90964 = ~n90962 & ~n90963;
  assign n90965 = n90244 & n90287;
  assign n90966 = n90238 & n90279;
  assign n90967 = ~n90965 & ~n90966;
  assign n90968 = n90267 & ~n90967;
  assign n90969 = n90259 & n90267;
  assign n90970 = ~n90238 & n90969;
  assign n90971 = ~n90968 & ~n90970;
  assign n90972 = n90964 & n90971;
  assign n90973 = ~n90273 & ~n90972;
  assign n90974 = ~n90296 & ~n90302;
  assign n90975 = ~n90906 & n90974;
  assign n90976 = n90310 & ~n90975;
  assign n90977 = ~n90973 & ~n90976;
  assign n90978 = ~n90278 & ~n90901;
  assign n90979 = ~n90267 & ~n90978;
  assign n90980 = n90977 & ~n90979;
  assign n90981 = ~n90959 & n90980;
  assign n90982 = ~pi2951 & n90981;
  assign n90983 = pi2951 & ~n90981;
  assign po3054 = n90982 | n90983;
  assign n90985 = n90104 & n90194;
  assign n90986 = ~n90154 & ~n90163;
  assign n90987 = ~n90104 & n90123;
  assign n90988 = n90104 & n90175;
  assign n90989 = ~n90987 & ~n90988;
  assign n90990 = n90986 & n90989;
  assign n90991 = n90133 & ~n90990;
  assign n90992 = ~n90116 & n90144;
  assign n90993 = ~n90104 & n90135;
  assign n90994 = ~n90134 & ~n90993;
  assign n90995 = ~n90992 & n90994;
  assign n90996 = ~n90133 & ~n90995;
  assign n90997 = n90122 & n90156;
  assign n90998 = n90110 & n90997;
  assign n90999 = ~n90996 & ~n90998;
  assign n91000 = ~n90991 & n90999;
  assign n91001 = ~n90985 & n91000;
  assign n91002 = ~n90098 & ~n91001;
  assign n91003 = n90133 & n90140;
  assign n91004 = ~n90104 & n91003;
  assign n91005 = n90133 & n90992;
  assign n91006 = n90133 & n90167;
  assign n91007 = ~n91005 & ~n91006;
  assign n91008 = n90104 & ~n91007;
  assign n91009 = ~n91004 & ~n91008;
  assign n91010 = n90104 & n90124;
  assign n91011 = ~n90206 & ~n91010;
  assign n91012 = ~n90104 & n90153;
  assign n91013 = n90104 & n90135;
  assign n91014 = ~n91012 & ~n91013;
  assign n91015 = ~n90124 & n91014;
  assign n91016 = ~n90154 & n91015;
  assign n91017 = ~n90133 & ~n91016;
  assign n91018 = n90104 & n90136;
  assign n91019 = ~n91017 & ~n91018;
  assign n91020 = n91011 & n91019;
  assign n91021 = n91009 & n91020;
  assign n91022 = n90098 & ~n91021;
  assign n91023 = n90133 & ~n90197;
  assign n91024 = ~n91022 & ~n91023;
  assign n91025 = ~n90158 & ~n91010;
  assign n91026 = ~n90133 & ~n91025;
  assign n91027 = n91024 & ~n91026;
  assign n91028 = ~n91002 & n91027;
  assign n91029 = pi2935 & ~n91028;
  assign n91030 = ~pi2935 & n91028;
  assign po3055 = n91029 | n91030;
  assign n91032 = n90696 & ~n90702;
  assign n91033 = ~n90740 & ~n91032;
  assign n91034 = ~n90772 & n91033;
  assign n91035 = n90721 & ~n91034;
  assign n91036 = ~n90715 & ~n90721;
  assign n91037 = n90702 & n91036;
  assign n91038 = ~n90696 & ~n90702;
  assign n91039 = n90715 & ~n90721;
  assign n91040 = n91038 & n91039;
  assign n91041 = n90696 & ~n90715;
  assign n91042 = n90708 & n91041;
  assign n91043 = n90715 & n90732;
  assign n91044 = ~n91042 & ~n91043;
  assign n91045 = ~n91040 & n91044;
  assign n91046 = ~n91037 & n91045;
  assign n91047 = ~n91035 & n91046;
  assign n91048 = n90690 & ~n91047;
  assign n91049 = n90696 & n90709;
  assign n91050 = n90715 & n91049;
  assign n91051 = n90696 & n90756;
  assign n91052 = ~n90715 & n91051;
  assign n91053 = ~n91050 & ~n91052;
  assign n91054 = n90721 & ~n91053;
  assign n91055 = ~n91048 & ~n91054;
  assign n91056 = ~n90715 & n90732;
  assign n91057 = ~n90744 & ~n90752;
  assign n91058 = n90721 & ~n91057;
  assign n91059 = ~n91056 & ~n91058;
  assign n91060 = ~n90748 & n91059;
  assign n91061 = ~n90690 & ~n91060;
  assign n91062 = ~n90738 & ~n90756;
  assign n91063 = ~n90696 & ~n91062;
  assign n91064 = ~n90757 & ~n91063;
  assign n91065 = ~n90721 & ~n91064;
  assign n91066 = ~n90690 & n91065;
  assign n91067 = ~n91061 & ~n91066;
  assign n91068 = n91055 & n91067;
  assign n91069 = pi2925 & ~n91068;
  assign n91070 = ~pi2925 & n91055;
  assign n91071 = n91067 & n91070;
  assign po3056 = n91069 | n91071;
  assign n91073 = ~n90480 & n90486;
  assign n91074 = ~n90492 & n90524;
  assign n91075 = n90492 & n90545;
  assign n91076 = ~n90492 & n90526;
  assign n91077 = ~n91075 & ~n91076;
  assign n91078 = ~n91074 & n91077;
  assign n91079 = n91073 & ~n91078;
  assign n91080 = n90504 & n90560;
  assign n91081 = n90492 & n91080;
  assign n91082 = ~n90530 & ~n91081;
  assign n91083 = ~n90504 & n90517;
  assign n91084 = ~n90527 & ~n91083;
  assign n91085 = n91082 & n91084;
  assign n91086 = ~n90486 & ~n91085;
  assign n91087 = ~n90504 & n90514;
  assign n91088 = n90492 & n91087;
  assign n91089 = ~n91086 & ~n91088;
  assign n91090 = ~n90480 & ~n91089;
  assign n91091 = ~n91079 & ~n91090;
  assign n91092 = n90504 & n90536;
  assign n91093 = ~n90498 & n91092;
  assign n91094 = ~n90531 & ~n91093;
  assign n91095 = ~n90526 & ~n90560;
  assign n91096 = n90492 & ~n91095;
  assign n91097 = ~n90561 & ~n91096;
  assign n91098 = n90486 & ~n91097;
  assign n91099 = ~n90515 & ~n91074;
  assign n91100 = ~n91075 & n91099;
  assign n91101 = ~n90486 & ~n91100;
  assign n91102 = ~n91098 & ~n91101;
  assign n91103 = n90492 & n90561;
  assign n91104 = ~n90547 & ~n91103;
  assign n91105 = ~n90566 & n91104;
  assign n91106 = ~n90539 & n91105;
  assign n91107 = n91102 & n91106;
  assign n91108 = n90480 & ~n91107;
  assign n91109 = n91094 & ~n91108;
  assign n91110 = n91091 & n91109;
  assign n91111 = pi2913 & ~n91110;
  assign n91112 = ~pi2913 & n91094;
  assign n91113 = n91091 & n91112;
  assign n91114 = ~n91108 & n91113;
  assign po3057 = n91111 | n91114;
  assign n91116 = ~n90515 & ~n90561;
  assign n91117 = n90486 & ~n91116;
  assign n91118 = n90492 & n90527;
  assign n91119 = ~n91117 & ~n91118;
  assign n91120 = n90492 & n90510;
  assign n91121 = ~n90511 & ~n91120;
  assign n91122 = ~n91080 & n91121;
  assign n91123 = ~n90486 & ~n91122;
  assign n91124 = n91119 & ~n91123;
  assign n91125 = ~n90480 & ~n91124;
  assign n91126 = ~n90566 & ~n90570;
  assign n91127 = ~n90486 & n90541;
  assign n91128 = n90492 & n90515;
  assign n91129 = n90486 & n90511;
  assign n91130 = ~n91128 & ~n91129;
  assign n91131 = ~n91103 & n91130;
  assign n91132 = ~n91127 & n91131;
  assign n91133 = n91126 & n91132;
  assign n91134 = ~n90553 & n91133;
  assign n91135 = n90480 & ~n91134;
  assign n91136 = n90486 & n90513;
  assign n91137 = ~n90559 & ~n91136;
  assign n91138 = ~n90567 & n91137;
  assign n91139 = ~n91135 & n91138;
  assign n91140 = ~n91125 & n91139;
  assign n91141 = ~pi2916 & ~n91140;
  assign n91142 = pi2916 & n91138;
  assign n91143 = ~n91125 & n91142;
  assign n91144 = ~n91135 & n91143;
  assign po3058 = n91141 | n91144;
  assign n91146 = ~n90378 & ~n90386;
  assign n91147 = n90328 & ~n91146;
  assign n91148 = ~n90391 & ~n90433;
  assign n91149 = ~n90354 & n91148;
  assign n91150 = ~n90361 & ~n91149;
  assign n91151 = n90328 & n91150;
  assign n91152 = ~n91147 & ~n91151;
  assign n91153 = n90377 & n90436;
  assign n91154 = ~n90438 & ~n91153;
  assign n91155 = ~n90403 & ~n90461;
  assign n91156 = n90361 & ~n91155;
  assign n91157 = n90328 & n91156;
  assign n91158 = n91154 & ~n91157;
  assign n91159 = ~n90392 & ~n90444;
  assign n91160 = n90334 & n90369;
  assign n91161 = ~n90428 & ~n91160;
  assign n91162 = n90361 & ~n91161;
  assign n91163 = n90334 & n90377;
  assign n91164 = n90334 & n90376;
  assign n91165 = ~n90416 & ~n91164;
  assign n91166 = ~n90361 & ~n91165;
  assign n91167 = ~n91163 & ~n91166;
  assign n91168 = ~n91162 & n91167;
  assign n91169 = n91159 & n91168;
  assign n91170 = ~n90328 & ~n91169;
  assign n91171 = ~n90334 & n90364;
  assign n91172 = ~n90444 & ~n91171;
  assign n91173 = ~n90464 & n91172;
  assign n91174 = n90361 & ~n91173;
  assign n91175 = ~n91170 & ~n91174;
  assign n91176 = n91158 & n91175;
  assign n91177 = n91152 & n91176;
  assign n91178 = ~pi2950 & ~n91177;
  assign n91179 = pi2950 & n91158;
  assign n91180 = n91152 & n91179;
  assign n91181 = n91175 & n91180;
  assign po3060 = n91178 | n91181;
  assign n91183 = n90605 & n90672;
  assign n91184 = ~n90653 & ~n90662;
  assign n91185 = n90611 & ~n91184;
  assign n91186 = ~n91183 & ~n91185;
  assign n91187 = ~n90647 & n91186;
  assign n91188 = ~n90611 & n90650;
  assign n91189 = ~n90640 & ~n91188;
  assign n91190 = ~n90670 & n91189;
  assign n91191 = n91187 & n91190;
  assign n91192 = n90586 & ~n91191;
  assign n91193 = n90605 & n90646;
  assign n91194 = ~n90624 & ~n91193;
  assign n91195 = n90599 & n90619;
  assign n91196 = n90611 & n91195;
  assign n91197 = n90605 & n90639;
  assign n91198 = ~n91196 & ~n91197;
  assign n91199 = ~n90598 & ~n90619;
  assign n91200 = n90592 & n90605;
  assign n91201 = ~n91199 & ~n91200;
  assign n91202 = ~n90676 & n91201;
  assign n91203 = ~n90611 & ~n91202;
  assign n91204 = ~n90605 & n90669;
  assign n91205 = ~n90635 & ~n91204;
  assign n91206 = ~n91203 & n91205;
  assign n91207 = n91198 & n91206;
  assign n91208 = n91194 & n91207;
  assign n91209 = ~n90586 & ~n91208;
  assign n91210 = ~n91192 & ~n91209;
  assign n91211 = pi2915 & ~n91210;
  assign n91212 = ~pi2915 & ~n91192;
  assign n91213 = ~n91209 & n91212;
  assign po3061 = n91211 | n91213;
  assign n91215 = ~n90751 & ~n91049;
  assign n91216 = n90725 & ~n91215;
  assign n91217 = ~n90747 & ~n90752;
  assign n91218 = ~n90744 & ~n91051;
  assign n91219 = n91217 & n91218;
  assign n91220 = ~n90715 & ~n91219;
  assign n91221 = ~n91216 & ~n91220;
  assign n91222 = ~n91043 & n91221;
  assign n91223 = n90690 & ~n91222;
  assign n91224 = ~n90715 & n91049;
  assign n91225 = n90715 & n90744;
  assign n91226 = ~n91224 & ~n91225;
  assign n91227 = ~n90721 & ~n91226;
  assign n91228 = ~n90715 & ~n91062;
  assign n91229 = ~n90696 & n91228;
  assign n91230 = ~n90708 & n91041;
  assign n91231 = ~n90780 & ~n91230;
  assign n91232 = ~n91051 & n91231;
  assign n91233 = n90721 & ~n91232;
  assign n91234 = ~n90721 & ~n91215;
  assign n91235 = ~n91233 & ~n91234;
  assign n91236 = ~n91229 & n91235;
  assign n91237 = ~n91225 & n91236;
  assign n91238 = ~n90690 & ~n91237;
  assign n91239 = ~n91227 & ~n91238;
  assign n91240 = ~n91223 & n91239;
  assign n91241 = ~pi2917 & ~n91240;
  assign n91242 = pi2917 & ~n91227;
  assign n91243 = ~n91223 & n91242;
  assign n91244 = ~n91238 & n91243;
  assign po3062 = n91241 | n91244;
  assign n91246 = ~n90450 & ~n90455;
  assign n91247 = ~n90392 & ~n90394;
  assign n91248 = ~n90460 & n91247;
  assign n91249 = ~n90361 & ~n91248;
  assign n91250 = ~n90418 & n91172;
  assign n91251 = n90361 & n90379;
  assign n91252 = n91250 & ~n91251;
  assign n91253 = ~n91249 & n91252;
  assign n91254 = n90328 & ~n91253;
  assign n91255 = n90334 & n90372;
  assign n91256 = ~n90346 & n90385;
  assign n91257 = ~n90394 & ~n91256;
  assign n91258 = n90361 & ~n91257;
  assign n91259 = ~n91255 & ~n91258;
  assign n91260 = ~n90361 & n90362;
  assign n91261 = n90334 & n91260;
  assign n91262 = ~n90361 & n90370;
  assign n91263 = ~n91261 & ~n91262;
  assign n91264 = n91259 & n91263;
  assign n91265 = ~n90346 & n90390;
  assign n91266 = ~n90427 & ~n91265;
  assign n91267 = ~n90464 & n91266;
  assign n91268 = n91264 & n91267;
  assign n91269 = ~n90328 & ~n91268;
  assign n91270 = ~n90427 & n91172;
  assign n91271 = ~n90361 & ~n91270;
  assign n91272 = ~n91269 & ~n91271;
  assign n91273 = ~n91254 & n91272;
  assign n91274 = n91246 & n91273;
  assign n91275 = pi2939 & ~n91274;
  assign n91276 = ~pi2939 & n91274;
  assign po3063 = n91275 | n91276;
  assign n91278 = ~n90486 & n90526;
  assign n91279 = ~n90492 & n91278;
  assign n91280 = ~n90571 & ~n91279;
  assign n91281 = n90492 & ~n90498;
  assign n91282 = n90504 & n91281;
  assign n91283 = ~n90492 & ~n90510;
  assign n91284 = ~n90570 & ~n91283;
  assign n91285 = n90486 & ~n91284;
  assign n91286 = ~n91282 & ~n91285;
  assign n91287 = n91280 & n91286;
  assign n91288 = n90480 & ~n91287;
  assign n91289 = ~n90545 & ~n90547;
  assign n91290 = ~n90492 & n90514;
  assign n91291 = n91289 & ~n91290;
  assign n91292 = ~n90486 & ~n91291;
  assign n91293 = n90486 & ~n90492;
  assign n91294 = n90526 & n91293;
  assign n91295 = ~n90531 & ~n91294;
  assign n91296 = ~n91292 & n91295;
  assign n91297 = ~n91080 & ~n91088;
  assign n91298 = n90486 & ~n91297;
  assign n91299 = n91296 & ~n91298;
  assign n91300 = ~n90480 & ~n91299;
  assign n91301 = ~n91288 & ~n91300;
  assign n91302 = n90492 & n91084;
  assign n91303 = ~n90492 & ~n90560;
  assign n91304 = ~n91302 & ~n91303;
  assign n91305 = n90486 & n91304;
  assign n91306 = ~n90545 & n91116;
  assign n91307 = n90549 & ~n91306;
  assign n91308 = ~n91305 & ~n91307;
  assign n91309 = n91301 & n91308;
  assign n91310 = ~pi2919 & ~n91309;
  assign n91311 = pi2919 & n91308;
  assign n91312 = ~n91300 & n91311;
  assign n91313 = ~n91288 & n91312;
  assign po3064 = n91310 | n91313;
  assign n91315 = n90715 & n90747;
  assign n91316 = ~n91043 & ~n91315;
  assign n91317 = ~n90721 & ~n91316;
  assign n91318 = n90744 & n91036;
  assign n91319 = ~n91317 & ~n91318;
  assign n91320 = ~n90768 & n91319;
  assign n91321 = ~n90715 & n90752;
  assign n91322 = ~n90747 & ~n91321;
  assign n91323 = ~n91051 & n91322;
  assign n91324 = ~n90721 & ~n91323;
  assign n91325 = n90690 & n91324;
  assign n91326 = n90721 & n91049;
  assign n91327 = ~n90740 & ~n90766;
  assign n91328 = ~n90734 & n91327;
  assign n91329 = ~n91326 & n91328;
  assign n91330 = n90690 & ~n91329;
  assign n91331 = n90696 & n90721;
  assign n91332 = ~n90708 & n91331;
  assign n91333 = ~n90702 & n91332;
  assign n91334 = n90715 & n91333;
  assign n91335 = ~n90715 & n90777;
  assign n91336 = ~n91333 & ~n91335;
  assign n91337 = ~n91042 & n91336;
  assign n91338 = ~n90708 & n90739;
  assign n91339 = ~n90715 & n90738;
  assign n91340 = ~n90743 & ~n91339;
  assign n91341 = ~n90721 & ~n91340;
  assign n91342 = ~n91338 & ~n91341;
  assign n91343 = n91337 & n91342;
  assign n91344 = ~n90690 & ~n91343;
  assign n91345 = ~n91334 & ~n91344;
  assign n91346 = ~n91330 & n91345;
  assign n91347 = ~n91325 & n91346;
  assign n91348 = n91320 & n91347;
  assign n91349 = pi2932 & ~n91348;
  assign n91350 = ~pi2932 & n91320;
  assign n91351 = n91347 & n91350;
  assign po3065 = n91349 | n91351;
  assign n91353 = ~n90200 & ~n91010;
  assign n91354 = ~n90998 & n91353;
  assign n91355 = n90133 & ~n91354;
  assign n91356 = ~n90209 & ~n90225;
  assign n91357 = ~n90206 & ~n91006;
  assign n91358 = ~n90194 & ~n91013;
  assign n91359 = ~n90133 & ~n91358;
  assign n91360 = ~n90163 & ~n91359;
  assign n91361 = n91357 & n91360;
  assign n91362 = n90098 & ~n91361;
  assign n91363 = ~n90116 & n90122;
  assign n91364 = ~n90141 & ~n91363;
  assign n91365 = ~n90104 & ~n91364;
  assign n91366 = ~n90124 & ~n90212;
  assign n91367 = ~n90133 & ~n91366;
  assign n91368 = ~n90104 & n90122;
  assign n91369 = ~n90136 & ~n91368;
  assign n91370 = ~n90144 & n91369;
  assign n91371 = n90133 & ~n91370;
  assign n91372 = ~n91367 & ~n91371;
  assign n91373 = ~n91365 & n91372;
  assign n91374 = ~n90098 & ~n91373;
  assign n91375 = ~n91362 & ~n91374;
  assign n91376 = n91356 & n91375;
  assign n91377 = ~n91355 & n91376;
  assign n91378 = ~pi2955 & ~n91377;
  assign n91379 = pi2955 & n91356;
  assign n91380 = ~n91355 & n91379;
  assign n91381 = n91375 & n91380;
  assign po3066 = n91378 | n91381;
  assign n91383 = pi6664 & pi9040;
  assign n91384 = pi6634 & ~pi9040;
  assign n91385 = ~n91383 & ~n91384;
  assign n91386 = ~pi2899 & n91385;
  assign n91387 = pi2899 & ~n91385;
  assign n91388 = ~n91386 & ~n91387;
  assign n91389 = pi6987 & ~pi9040;
  assign n91390 = pi6766 & pi9040;
  assign n91391 = ~n91389 & ~n91390;
  assign n91392 = ~pi2906 & n91391;
  assign n91393 = pi2906 & ~n91391;
  assign n91394 = ~n91392 & ~n91393;
  assign n91395 = pi6667 & ~pi9040;
  assign n91396 = pi6722 & pi9040;
  assign n91397 = ~n91395 & ~n91396;
  assign n91398 = ~pi2895 & n91397;
  assign n91399 = pi2895 & ~n91397;
  assign n91400 = ~n91398 & ~n91399;
  assign n91401 = n91394 & ~n91400;
  assign n91402 = ~n91388 & n91401;
  assign n91403 = pi6799 & pi9040;
  assign n91404 = pi6731 & ~pi9040;
  assign n91405 = ~n91403 & ~n91404;
  assign n91406 = ~pi2890 & n91405;
  assign n91407 = pi2890 & ~n91405;
  assign n91408 = ~n91406 & ~n91407;
  assign n91409 = n91388 & ~n91408;
  assign n91410 = n91400 & n91409;
  assign n91411 = ~n91388 & ~n91408;
  assign n91412 = ~n91400 & n91411;
  assign n91413 = ~n91410 & ~n91412;
  assign n91414 = ~n91402 & n91413;
  assign n91415 = pi6721 & pi9040;
  assign n91416 = pi6799 & ~pi9040;
  assign n91417 = ~n91415 & ~n91416;
  assign n91418 = ~pi2873 & n91417;
  assign n91419 = pi2873 & ~n91417;
  assign n91420 = ~n91418 & ~n91419;
  assign n91421 = pi6730 & pi9040;
  assign n91422 = pi6763 & ~pi9040;
  assign n91423 = ~n91421 & ~n91422;
  assign n91424 = pi2880 & n91423;
  assign n91425 = ~pi2880 & ~n91423;
  assign n91426 = ~n91424 & ~n91425;
  assign n91427 = n91420 & n91426;
  assign n91428 = ~n91414 & n91427;
  assign n91429 = n91388 & n91408;
  assign n91430 = ~n91400 & n91429;
  assign n91431 = ~n91394 & n91426;
  assign n91432 = n91430 & n91431;
  assign n91433 = ~n91400 & n91409;
  assign n91434 = ~n91420 & n91433;
  assign n91435 = ~n91388 & n91408;
  assign n91436 = ~n91394 & n91435;
  assign n91437 = ~n91388 & n91400;
  assign n91438 = ~n91436 & ~n91437;
  assign n91439 = ~n91420 & ~n91438;
  assign n91440 = ~n91434 & ~n91439;
  assign n91441 = n91426 & ~n91440;
  assign n91442 = ~n91432 & ~n91441;
  assign n91443 = ~n91394 & n91400;
  assign n91444 = ~n91388 & n91443;
  assign n91445 = n91394 & n91400;
  assign n91446 = n91388 & n91445;
  assign n91447 = n91408 & n91446;
  assign n91448 = ~n91444 & ~n91447;
  assign n91449 = ~n91420 & ~n91448;
  assign n91450 = n91442 & ~n91449;
  assign n91451 = ~n91394 & n91420;
  assign n91452 = n91435 & n91451;
  assign n91453 = ~n91400 & n91452;
  assign n91454 = ~n91411 & ~n91429;
  assign n91455 = n91401 & ~n91454;
  assign n91456 = n91394 & n91410;
  assign n91457 = ~n91455 & ~n91456;
  assign n91458 = n91400 & n91435;
  assign n91459 = n91394 & n91420;
  assign n91460 = n91458 & n91459;
  assign n91461 = n91443 & ~n91454;
  assign n91462 = ~n91394 & ~n91400;
  assign n91463 = n91388 & n91462;
  assign n91464 = ~n91408 & n91463;
  assign n91465 = ~n91461 & ~n91464;
  assign n91466 = ~n91460 & n91465;
  assign n91467 = n91457 & n91466;
  assign n91468 = ~n91453 & n91467;
  assign n91469 = n91394 & ~n91420;
  assign n91470 = ~n91400 & n91469;
  assign n91471 = n91408 & n91470;
  assign n91472 = n91468 & ~n91471;
  assign n91473 = ~n91426 & ~n91472;
  assign n91474 = n91450 & ~n91473;
  assign n91475 = ~n91428 & n91474;
  assign n91476 = ~pi2942 & ~n91475;
  assign n91477 = pi2942 & n91450;
  assign n91478 = ~n91428 & n91477;
  assign n91479 = ~n91473 & n91478;
  assign po3067 = n91476 | n91479;
  assign n91481 = ~n90605 & n90626;
  assign n91482 = ~n91204 & ~n91481;
  assign n91483 = n90611 & n91482;
  assign n91484 = n90605 & n90664;
  assign n91485 = ~n90599 & ~n90620;
  assign n91486 = ~n90619 & ~n91485;
  assign n91487 = ~n90592 & n90633;
  assign n91488 = n90605 & n90620;
  assign n91489 = ~n91487 & ~n91488;
  assign n91490 = ~n90611 & n91489;
  assign n91491 = ~n91486 & n91490;
  assign n91492 = ~n91484 & n91491;
  assign n91493 = ~n91483 & ~n91492;
  assign n91494 = n90605 & n91486;
  assign n91495 = ~n91193 & ~n91494;
  assign n91496 = ~n91493 & n91495;
  assign n91497 = n90586 & ~n91496;
  assign n91498 = n90611 & ~n91485;
  assign n91499 = ~n90605 & n91498;
  assign n91500 = ~n90641 & ~n90668;
  assign n91501 = n90605 & ~n91500;
  assign n91502 = n90611 & n91501;
  assign n91503 = n90619 & n91498;
  assign n91504 = ~n91502 & ~n91503;
  assign n91505 = ~n91499 & n91504;
  assign n91506 = ~n90586 & ~n91505;
  assign n91507 = ~n91497 & ~n91506;
  assign n91508 = n90611 & n90624;
  assign n91509 = ~n90611 & ~n91495;
  assign n91510 = ~n91508 & ~n91509;
  assign n91511 = ~n90611 & ~n91482;
  assign n91512 = ~n90624 & ~n91511;
  assign n91513 = ~n90586 & ~n91512;
  assign n91514 = n91510 & ~n91513;
  assign n91515 = n91507 & n91514;
  assign n91516 = pi2928 & ~n91515;
  assign n91517 = ~n91497 & n91514;
  assign n91518 = ~n91506 & n91517;
  assign n91519 = ~pi2928 & n91518;
  assign po3068 = n91516 | n91519;
  assign n91521 = ~n91400 & n91435;
  assign n91522 = ~n91420 & n91521;
  assign n91523 = n91394 & n91522;
  assign n91524 = n91409 & n91469;
  assign n91525 = n91400 & n91524;
  assign n91526 = ~n91523 & ~n91525;
  assign n91527 = ~n91456 & ~n91460;
  assign n91528 = ~n91400 & ~n91408;
  assign n91529 = ~n91394 & n91528;
  assign n91530 = ~n91436 & ~n91529;
  assign n91531 = ~n91420 & ~n91530;
  assign n91532 = n91420 & ~n91445;
  assign n91533 = ~n91454 & n91532;
  assign n91534 = n91394 & ~n91435;
  assign n91535 = ~n91420 & n91534;
  assign n91536 = n91400 & n91535;
  assign n91537 = ~n91533 & ~n91536;
  assign n91538 = ~n91531 & n91537;
  assign n91539 = n91527 & n91538;
  assign n91540 = n91426 & ~n91539;
  assign n91541 = n91526 & ~n91540;
  assign n91542 = n91412 & n91420;
  assign n91543 = ~n91394 & n91542;
  assign n91544 = ~n91433 & ~n91436;
  assign n91545 = n91445 & ~n91454;
  assign n91546 = n91544 & ~n91545;
  assign n91547 = n91420 & ~n91426;
  assign n91548 = ~n91546 & n91547;
  assign n91549 = ~n91543 & ~n91548;
  assign n91550 = ~n91394 & n91410;
  assign n91551 = ~n91394 & ~n91408;
  assign n91552 = n91400 & n91551;
  assign n91553 = ~n91394 & n91429;
  assign n91554 = ~n91552 & ~n91553;
  assign n91555 = n91394 & n91435;
  assign n91556 = ~n91430 & ~n91555;
  assign n91557 = n91554 & n91556;
  assign n91558 = ~n91420 & ~n91557;
  assign n91559 = ~n91550 & ~n91558;
  assign n91560 = ~n91426 & ~n91559;
  assign n91561 = n91549 & ~n91560;
  assign n91562 = n91541 & n91561;
  assign n91563 = pi2940 & ~n91562;
  assign n91564 = ~pi2940 & n91541;
  assign n91565 = n91561 & n91564;
  assign po3069 = n91563 | n91565;
  assign n91567 = ~n90824 & ~n90830;
  assign n91568 = n90797 & ~n91567;
  assign n91569 = ~n90885 & ~n91568;
  assign n91570 = n90803 & n90809;
  assign n91571 = ~n90797 & n91570;
  assign n91572 = n90823 & n91571;
  assign n91573 = n90823 & n90837;
  assign n91574 = ~n91570 & ~n91573;
  assign n91575 = ~n90809 & n90849;
  assign n91576 = n91574 & ~n91575;
  assign n91577 = ~n90797 & ~n91576;
  assign n91578 = ~n90833 & ~n91577;
  assign n91579 = ~n90861 & ~n91578;
  assign n91580 = n90797 & n90816;
  assign n91581 = n90823 & n91580;
  assign n91582 = n90797 & n90829;
  assign n91583 = ~n91581 & ~n91582;
  assign n91584 = ~n90861 & ~n91583;
  assign n91585 = ~n91579 & ~n91584;
  assign n91586 = ~n91572 & n91585;
  assign n91587 = ~n90809 & n90867;
  assign n91588 = ~n90803 & n90837;
  assign n91589 = ~n90868 & ~n91588;
  assign n91590 = ~n90803 & n90831;
  assign n91591 = n91589 & ~n91590;
  assign n91592 = n90797 & ~n91591;
  assign n91593 = ~n90823 & n90829;
  assign n91594 = ~n90852 & ~n91593;
  assign n91595 = ~n90797 & ~n91594;
  assign n91596 = ~n91592 & ~n91595;
  assign n91597 = ~n91587 & n91596;
  assign n91598 = ~n90839 & ~n90879;
  assign n91599 = n91597 & n91598;
  assign n91600 = n90861 & ~n91599;
  assign n91601 = n91586 & ~n91600;
  assign n91602 = n91569 & n91601;
  assign n91603 = ~pi2933 & ~n91602;
  assign n91604 = pi2933 & n91586;
  assign n91605 = n91569 & n91604;
  assign n91606 = ~n91600 & n91605;
  assign po3070 = n91603 | n91606;
  assign n91608 = ~n90238 & n90279;
  assign n91609 = ~n90293 & ~n91608;
  assign n91610 = ~n90267 & ~n91609;
  assign n91611 = n90267 & ~n90928;
  assign n91612 = ~n90917 & ~n91611;
  assign n91613 = ~n91610 & n91612;
  assign n91614 = n90273 & ~n91613;
  assign n91615 = n90260 & ~n90267;
  assign n91616 = ~n91614 & ~n91615;
  assign n91617 = ~n90952 & ~n90966;
  assign n91618 = n90267 & ~n91617;
  assign n91619 = n90267 & n90294;
  assign n91620 = n90238 & n90280;
  assign n91621 = ~n90267 & n90277;
  assign n91622 = ~n90904 & ~n91621;
  assign n91623 = ~n90244 & ~n91622;
  assign n91624 = ~n90949 & ~n91623;
  assign n91625 = ~n90278 & n91624;
  assign n91626 = ~n91620 & n91625;
  assign n91627 = ~n91619 & n91626;
  assign n91628 = ~n90273 & ~n91627;
  assign n91629 = ~n91618 & ~n91628;
  assign n91630 = n91616 & n91629;
  assign n91631 = pi2958 & ~n91630;
  assign n91632 = ~pi2958 & n91630;
  assign po3071 = n91631 | n91632;
  assign n91634 = ~n91553 & ~n91555;
  assign n91635 = ~n91420 & ~n91634;
  assign n91636 = ~n91525 & ~n91635;
  assign n91637 = n91426 & ~n91636;
  assign n91638 = ~n91411 & n91462;
  assign n91639 = n91426 & n91638;
  assign n91640 = n91411 & n91443;
  assign n91641 = ~n91420 & n91640;
  assign n91642 = ~n91400 & n91451;
  assign n91643 = n91388 & n91642;
  assign n91644 = ~n91641 & ~n91643;
  assign n91645 = ~n91639 & n91644;
  assign n91646 = n91400 & ~n91408;
  assign n91647 = ~n91411 & ~n91646;
  assign n91648 = n91394 & ~n91647;
  assign n91649 = ~n91521 & ~n91648;
  assign n91650 = n91420 & ~n91649;
  assign n91651 = ~n91545 & ~n91650;
  assign n91652 = ~n91394 & n91458;
  assign n91653 = n91388 & n91401;
  assign n91654 = ~n91394 & ~n91647;
  assign n91655 = ~n91653 & ~n91654;
  assign n91656 = ~n91420 & ~n91655;
  assign n91657 = ~n91652 & ~n91656;
  assign n91658 = n91651 & n91657;
  assign n91659 = ~n91426 & ~n91658;
  assign n91660 = ~n91430 & ~n91551;
  assign n91661 = n91427 & ~n91660;
  assign n91662 = ~n91659 & ~n91661;
  assign n91663 = n91645 & n91662;
  assign n91664 = ~n91637 & n91663;
  assign n91665 = pi2943 & ~n91664;
  assign n91666 = ~pi2943 & n91664;
  assign po3072 = n91665 | n91666;
  assign n91668 = n90797 & ~n90823;
  assign n91669 = ~n90815 & n91668;
  assign n91670 = ~n90809 & n91669;
  assign n91671 = n90831 & n90864;
  assign n91672 = ~n91670 & ~n91671;
  assign n91673 = n90823 & n90863;
  assign n91674 = ~n91588 & ~n91673;
  assign n91675 = ~n90797 & ~n91674;
  assign n91676 = n91672 & ~n91675;
  assign n91677 = ~n90839 & ~n90878;
  assign n91678 = ~n91582 & n91677;
  assign n91679 = ~n90823 & n90852;
  assign n91680 = ~n90827 & ~n91679;
  assign n91681 = n91678 & n91680;
  assign n91682 = n91676 & n91681;
  assign n91683 = ~n90861 & ~n91682;
  assign n91684 = ~n90826 & ~n91588;
  assign n91685 = n90823 & ~n91684;
  assign n91686 = ~n91587 & ~n91590;
  assign n91687 = ~n90803 & ~n90815;
  assign n91688 = n90823 & n91687;
  assign n91689 = n91686 & ~n91688;
  assign n91690 = ~n90797 & ~n91689;
  assign n91691 = ~n90823 & n90837;
  assign n91692 = n90803 & n90823;
  assign n91693 = ~n90815 & n91692;
  assign n91694 = ~n90809 & n91693;
  assign n91695 = ~n91691 & ~n91694;
  assign n91696 = n90797 & ~n91695;
  assign n91697 = ~n90823 & n90832;
  assign n91698 = ~n91696 & ~n91697;
  assign n91699 = ~n91690 & n91698;
  assign n91700 = ~n91685 & n91699;
  assign n91701 = n90861 & ~n91700;
  assign n91702 = ~n90797 & n90868;
  assign n91703 = ~n91701 & ~n91702;
  assign n91704 = n90844 & n91668;
  assign n91705 = ~n90815 & n91704;
  assign n91706 = n91703 & ~n91705;
  assign n91707 = ~n91683 & n91706;
  assign n91708 = ~pi2922 & ~n91707;
  assign n91709 = pi2922 & n91703;
  assign n91710 = ~n91683 & n91709;
  assign n91711 = ~n91705 & n91710;
  assign po3074 = n91708 | n91711;
  assign n91713 = n91400 & n91411;
  assign n91714 = ~n91521 & ~n91713;
  assign n91715 = ~n91420 & ~n91714;
  assign n91716 = n91394 & n91429;
  assign n91717 = ~n91412 & ~n91716;
  assign n91718 = ~n91458 & n91717;
  assign n91719 = n91420 & ~n91718;
  assign n91720 = ~n91715 & ~n91719;
  assign n91721 = ~n91434 & ~n91447;
  assign n91722 = n91720 & n91721;
  assign n91723 = ~n91426 & ~n91722;
  assign n91724 = ~n91394 & n91521;
  assign n91725 = n91394 & n91409;
  assign n91726 = ~n91553 & ~n91725;
  assign n91727 = n91420 & ~n91726;
  assign n91728 = ~n91724 & ~n91727;
  assign n91729 = ~n91400 & ~n91420;
  assign n91730 = n91388 & n91729;
  assign n91731 = n91408 & n91730;
  assign n91732 = n91413 & ~n91731;
  assign n91733 = ~n91458 & n91732;
  assign n91734 = n91394 & ~n91733;
  assign n91735 = n91728 & ~n91734;
  assign n91736 = n91426 & ~n91735;
  assign n91737 = ~n91723 & ~n91736;
  assign n91738 = n91400 & n91553;
  assign n91739 = ~n91464 & ~n91738;
  assign n91740 = ~n91420 & ~n91739;
  assign n91741 = n91451 & n91646;
  assign n91742 = ~n91740 & ~n91741;
  assign n91743 = n91737 & n91742;
  assign n91744 = ~pi2927 & ~n91743;
  assign n91745 = pi2927 & ~n91740;
  assign n91746 = n91737 & n91745;
  assign n91747 = ~n91741 & n91746;
  assign po3075 = n91744 | n91747;
  assign n91749 = n90605 & n91195;
  assign n91750 = n90611 & n91749;
  assign n91751 = n90633 & ~n91485;
  assign n91752 = ~n90669 & ~n91751;
  assign n91753 = ~n91193 & n91752;
  assign n91754 = ~n90611 & ~n91753;
  assign n91755 = n90605 & n90621;
  assign n91756 = ~n91754 & ~n91755;
  assign n91757 = n90619 & n90668;
  assign n91758 = ~n90605 & n91199;
  assign n91759 = ~n91757 & ~n91758;
  assign n91760 = ~n91488 & n91759;
  assign n91761 = n90611 & ~n91760;
  assign n91762 = n91756 & ~n91761;
  assign n91763 = n90586 & ~n91762;
  assign n91764 = ~n91750 & ~n91763;
  assign n91765 = ~n90605 & n90620;
  assign n91766 = ~n90646 & ~n91765;
  assign n91767 = n90611 & ~n91766;
  assign n91768 = ~n90670 & ~n91767;
  assign n91769 = ~n90642 & ~n91749;
  assign n91770 = n90605 & n90676;
  assign n91771 = ~n91199 & ~n91770;
  assign n91772 = ~n91757 & n91771;
  assign n91773 = ~n90611 & ~n91772;
  assign n91774 = ~n90605 & n90621;
  assign n91775 = ~n91773 & ~n91774;
  assign n91776 = n91769 & n91775;
  assign n91777 = n91768 & n91776;
  assign n91778 = ~n90586 & ~n91777;
  assign n91779 = ~n90656 & ~n91484;
  assign n91780 = ~n90611 & ~n91779;
  assign n91781 = ~n91778 & ~n91780;
  assign n91782 = n91764 & n91781;
  assign n91783 = pi2931 & n91782;
  assign n91784 = ~pi2931 & ~n91782;
  assign po3076 = n91783 | n91784;
  assign n91786 = ~n90879 & ~n91697;
  assign n91787 = ~n90797 & ~n91786;
  assign n91788 = ~n90861 & n90863;
  assign n91789 = n90797 & n91788;
  assign n91790 = n90809 & n90849;
  assign n91791 = ~n91687 & ~n91790;
  assign n91792 = ~n90832 & n91791;
  assign n91793 = ~n90797 & ~n91792;
  assign n91794 = ~n90823 & n90838;
  assign n91795 = ~n91793 & ~n91794;
  assign n91796 = ~n90861 & ~n91795;
  assign n91797 = ~n91789 & ~n91796;
  assign n91798 = ~n90827 & ~n90830;
  assign n91799 = ~n90823 & n91590;
  assign n91800 = ~n91673 & ~n91799;
  assign n91801 = n91798 & n91800;
  assign n91802 = n90797 & ~n91801;
  assign n91803 = n90803 & ~n90809;
  assign n91804 = n90797 & n91803;
  assign n91805 = n90823 & n91804;
  assign n91806 = ~n90823 & n91687;
  assign n91807 = ~n90830 & ~n91806;
  assign n91808 = ~n91694 & n91807;
  assign n91809 = ~n91805 & n91808;
  assign n91810 = ~n90797 & n90826;
  assign n91811 = n91809 & ~n91810;
  assign n91812 = n90861 & ~n91811;
  assign n91813 = ~n91802 & ~n91812;
  assign n91814 = n91797 & n91813;
  assign n91815 = ~n91787 & n91814;
  assign n91816 = pi2948 & n91815;
  assign n91817 = ~pi2948 & ~n91815;
  assign po3077 = n91816 | n91817;
  assign n91819 = ~pi6868 & pi9040;
  assign n91820 = pi6999 & ~pi9040;
  assign n91821 = ~n91819 & ~n91820;
  assign n91822 = ~pi2961 & ~n91821;
  assign n91823 = pi2961 & n91821;
  assign n91824 = ~n91822 & ~n91823;
  assign n91825 = pi6879 & ~pi9040;
  assign n91826 = pi7018 & pi9040;
  assign n91827 = ~n91825 & ~n91826;
  assign n91828 = ~pi2970 & n91827;
  assign n91829 = pi2970 & ~n91827;
  assign n91830 = ~n91828 & ~n91829;
  assign n91831 = pi6936 & pi9040;
  assign n91832 = pi6913 & ~pi9040;
  assign n91833 = ~n91831 & ~n91832;
  assign n91834 = ~pi2936 & ~n91833;
  assign n91835 = pi2936 & n91833;
  assign n91836 = ~n91834 & ~n91835;
  assign n91837 = n91830 & n91836;
  assign n91838 = pi6909 & pi9040;
  assign n91839 = pi6864 & ~pi9040;
  assign n91840 = ~n91838 & ~n91839;
  assign n91841 = pi2956 & n91840;
  assign n91842 = ~pi2956 & ~n91840;
  assign n91843 = ~n91841 & ~n91842;
  assign n91844 = pi6884 & ~pi9040;
  assign n91845 = pi7080 & pi9040;
  assign n91846 = ~n91844 & ~n91845;
  assign n91847 = pi2949 & n91846;
  assign n91848 = ~pi2949 & ~n91846;
  assign n91849 = ~n91847 & ~n91848;
  assign n91850 = ~n91843 & ~n91849;
  assign n91851 = n91837 & n91850;
  assign n91852 = pi6999 & pi9040;
  assign n91853 = pi7028 & ~pi9040;
  assign n91854 = ~n91852 & ~n91853;
  assign n91855 = ~pi2953 & n91854;
  assign n91856 = pi2953 & ~n91854;
  assign n91857 = ~n91855 & ~n91856;
  assign n91858 = ~n91830 & ~n91836;
  assign n91859 = ~n91857 & n91858;
  assign n91860 = n91843 & n91857;
  assign n91861 = ~n91836 & n91860;
  assign n91862 = n91830 & n91861;
  assign n91863 = ~n91859 & ~n91862;
  assign n91864 = ~n91830 & n91836;
  assign n91865 = n91843 & n91864;
  assign n91866 = n91863 & ~n91865;
  assign n91867 = ~n91849 & ~n91866;
  assign n91868 = ~n91830 & n91857;
  assign n91869 = ~n91843 & n91849;
  assign n91870 = n91868 & n91869;
  assign n91871 = n91857 & n91858;
  assign n91872 = ~n91843 & n91871;
  assign n91873 = ~n91870 & ~n91872;
  assign n91874 = ~n91867 & n91873;
  assign n91875 = ~n91851 & n91874;
  assign n91876 = ~n91857 & n91864;
  assign n91877 = n91843 & n91876;
  assign n91878 = n91837 & ~n91857;
  assign n91879 = ~n91843 & n91878;
  assign n91880 = ~n91877 & ~n91879;
  assign n91881 = n91875 & n91880;
  assign n91882 = ~n91824 & ~n91881;
  assign n91883 = n91836 & n91868;
  assign n91884 = ~n91843 & n91883;
  assign n91885 = ~n91878 & ~n91884;
  assign n91886 = ~n91849 & ~n91885;
  assign n91887 = n91837 & n91860;
  assign n91888 = ~n91843 & n91857;
  assign n91889 = ~n91836 & n91888;
  assign n91890 = n91830 & n91889;
  assign n91891 = ~n91887 & ~n91890;
  assign n91892 = ~n91830 & n91860;
  assign n91893 = ~n91843 & n91876;
  assign n91894 = ~n91892 & ~n91893;
  assign n91895 = n91849 & ~n91894;
  assign n91896 = n91891 & ~n91895;
  assign n91897 = ~n91886 & n91896;
  assign n91898 = n91824 & ~n91897;
  assign n91899 = ~n91830 & ~n91857;
  assign n91900 = n91843 & n91899;
  assign n91901 = n91830 & ~n91857;
  assign n91902 = ~n91843 & n91901;
  assign n91903 = ~n91900 & ~n91902;
  assign n91904 = ~n91849 & ~n91903;
  assign n91905 = n91830 & ~n91836;
  assign n91906 = ~n91857 & n91905;
  assign n91907 = n91843 & n91906;
  assign n91908 = ~n91887 & ~n91907;
  assign n91909 = ~n91871 & n91908;
  assign n91910 = n91849 & ~n91909;
  assign n91911 = ~n91904 & ~n91910;
  assign n91912 = ~n91836 & n91857;
  assign n91913 = n91849 & n91912;
  assign n91914 = ~n91843 & n91913;
  assign n91915 = n91911 & ~n91914;
  assign n91916 = ~n91898 & n91915;
  assign n91917 = ~n91882 & n91916;
  assign n91918 = ~pi3189 & ~n91917;
  assign n91919 = pi3189 & n91917;
  assign po3098 = n91918 | n91919;
  assign n91921 = pi6895 & ~pi9040;
  assign n91922 = pi7028 & pi9040;
  assign n91923 = ~n91921 & ~n91922;
  assign n91924 = pi2945 & n91923;
  assign n91925 = ~pi2945 & ~n91923;
  assign n91926 = ~n91924 & ~n91925;
  assign n91927 = pi7020 & pi9040;
  assign n91928 = pi6860 & ~pi9040;
  assign n91929 = ~n91927 & ~n91928;
  assign n91930 = ~pi2936 & n91929;
  assign n91931 = pi2936 & ~n91929;
  assign n91932 = ~n91930 & ~n91931;
  assign n91933 = pi7011 & pi9040;
  assign n91934 = pi6889 & ~pi9040;
  assign n91935 = ~n91933 & ~n91934;
  assign n91936 = ~pi2972 & n91935;
  assign n91937 = pi2972 & ~n91935;
  assign n91938 = ~n91936 & ~n91937;
  assign n91939 = pi6872 & ~pi9040;
  assign n91940 = pi6989 & pi9040;
  assign n91941 = ~n91939 & ~n91940;
  assign n91942 = ~pi2961 & n91941;
  assign n91943 = pi2961 & ~n91941;
  assign n91944 = ~n91942 & ~n91943;
  assign n91945 = ~n91938 & ~n91944;
  assign n91946 = n91932 & n91945;
  assign n91947 = pi7063 & ~pi9040;
  assign n91948 = pi6874 & pi9040;
  assign n91949 = ~n91947 & ~n91948;
  assign n91950 = ~pi2969 & ~n91949;
  assign n91951 = pi2969 & n91949;
  assign n91952 = ~n91950 & ~n91951;
  assign n91953 = n91946 & ~n91952;
  assign n91954 = n91938 & n91944;
  assign n91955 = n91932 & n91954;
  assign n91956 = ~n91952 & n91955;
  assign n91957 = ~n91953 & ~n91956;
  assign n91958 = ~n91932 & n91954;
  assign n91959 = n91952 & n91958;
  assign n91960 = ~n91938 & n91944;
  assign n91961 = n91932 & n91960;
  assign n91962 = n91952 & n91961;
  assign n91963 = ~n91959 & ~n91962;
  assign n91964 = n91957 & n91963;
  assign n91965 = n91926 & ~n91964;
  assign n91966 = n91938 & ~n91944;
  assign n91967 = n91932 & n91966;
  assign n91968 = n91952 & n91967;
  assign n91969 = ~n91961 & ~n91968;
  assign n91970 = n91926 & ~n91969;
  assign n91971 = ~n91926 & ~n91944;
  assign n91972 = ~n91952 & n91971;
  assign n91973 = ~n91932 & ~n91938;
  assign n91974 = n91952 & n91954;
  assign n91975 = ~n91973 & ~n91974;
  assign n91976 = ~n91926 & ~n91975;
  assign n91977 = ~n91972 & ~n91976;
  assign n91978 = ~n91932 & n91966;
  assign n91979 = ~n91952 & n91978;
  assign n91980 = n91977 & ~n91979;
  assign n91981 = ~n91944 & n91952;
  assign n91982 = ~n91932 & n91981;
  assign n91983 = ~n91938 & n91982;
  assign n91984 = n91980 & ~n91983;
  assign n91985 = ~n91970 & n91984;
  assign n91986 = pi6860 & pi9040;
  assign n91987 = pi7018 & ~pi9040;
  assign n91988 = ~n91986 & ~n91987;
  assign n91989 = pi2967 & n91988;
  assign n91990 = ~pi2967 & ~n91988;
  assign n91991 = ~n91989 & ~n91990;
  assign n91992 = ~n91985 & ~n91991;
  assign n91993 = n91932 & ~n91944;
  assign n91994 = ~n91926 & n91952;
  assign n91995 = n91991 & n91994;
  assign n91996 = n91993 & n91995;
  assign n91997 = n91932 & ~n91952;
  assign n91998 = n91944 & n91997;
  assign n91999 = ~n91926 & ~n91998;
  assign n92000 = ~n91932 & n91952;
  assign n92001 = n91938 & n92000;
  assign n92002 = ~n91945 & ~n91993;
  assign n92003 = ~n91952 & ~n92002;
  assign n92004 = ~n91958 & ~n92003;
  assign n92005 = n91926 & n92004;
  assign n92006 = ~n92001 & n92005;
  assign n92007 = ~n91999 & ~n92006;
  assign n92008 = n91944 & n92000;
  assign n92009 = ~n91938 & n92008;
  assign n92010 = ~n92007 & ~n92009;
  assign n92011 = n91991 & ~n92010;
  assign n92012 = ~n91996 & ~n92011;
  assign n92013 = ~n91992 & n92012;
  assign n92014 = ~n91965 & n92013;
  assign n92015 = ~n91926 & n91979;
  assign n92016 = n92014 & ~n92015;
  assign n92017 = pi3191 & ~n92016;
  assign n92018 = ~pi3191 & ~n92015;
  assign n92019 = n92013 & n92018;
  assign n92020 = ~n91965 & n92019;
  assign po3102 = n92017 | n92020;
  assign n92022 = pi6927 & ~pi9040;
  assign n92023 = pi6872 & pi9040;
  assign n92024 = ~n92022 & ~n92023;
  assign n92025 = ~pi2970 & ~n92024;
  assign n92026 = pi2970 & n92024;
  assign n92027 = ~n92025 & ~n92026;
  assign n92028 = pi6870 & pi9040;
  assign n92029 = pi7011 & ~pi9040;
  assign n92030 = ~n92028 & ~n92029;
  assign n92031 = pi2957 & n92030;
  assign n92032 = ~pi2957 & ~n92030;
  assign n92033 = ~n92031 & ~n92032;
  assign n92034 = pi6895 & pi9040;
  assign n92035 = pi6922 & ~pi9040;
  assign n92036 = ~n92034 & ~n92035;
  assign n92037 = pi2938 & n92036;
  assign n92038 = ~pi2938 & ~n92036;
  assign n92039 = ~n92037 & ~n92038;
  assign n92040 = pi6913 & pi9040;
  assign n92041 = pi6915 & ~pi9040;
  assign n92042 = ~n92040 & ~n92041;
  assign n92043 = ~pi2954 & ~n92042;
  assign n92044 = pi2954 & n92042;
  assign n92045 = ~n92043 & ~n92044;
  assign n92046 = pi6870 & ~pi9040;
  assign n92047 = pi7016 & pi9040;
  assign n92048 = ~n92046 & ~n92047;
  assign n92049 = ~pi2962 & n92048;
  assign n92050 = pi2962 & ~n92048;
  assign n92051 = ~n92049 & ~n92050;
  assign n92052 = n92045 & n92051;
  assign n92053 = n92039 & n92052;
  assign n92054 = pi7013 & ~pi9040;
  assign n92055 = pi6927 & pi9040;
  assign n92056 = ~n92054 & ~n92055;
  assign n92057 = ~pi2953 & ~n92056;
  assign n92058 = pi2953 & n92056;
  assign n92059 = ~n92057 & ~n92058;
  assign n92060 = ~n92051 & n92059;
  assign n92061 = n92045 & n92060;
  assign n92062 = ~n92053 & ~n92061;
  assign n92063 = ~n92051 & ~n92059;
  assign n92064 = ~n92045 & n92063;
  assign n92065 = ~n92039 & n92064;
  assign n92066 = n92062 & ~n92065;
  assign n92067 = n92033 & ~n92066;
  assign n92068 = ~n92045 & ~n92051;
  assign n92069 = n92059 & n92068;
  assign n92070 = ~n92039 & n92069;
  assign n92071 = n92051 & n92059;
  assign n92072 = n92045 & n92071;
  assign n92073 = ~n92039 & n92072;
  assign n92074 = ~n92045 & n92051;
  assign n92075 = ~n92063 & ~n92074;
  assign n92076 = n92039 & ~n92075;
  assign n92077 = ~n92073 & ~n92076;
  assign n92078 = ~n92070 & n92077;
  assign n92079 = ~n92033 & ~n92078;
  assign n92080 = ~n92067 & ~n92079;
  assign n92081 = n92027 & ~n92080;
  assign n92082 = n92033 & ~n92039;
  assign n92083 = n92051 & n92082;
  assign n92084 = ~n92033 & ~n92039;
  assign n92085 = n92063 & n92084;
  assign n92086 = ~n92039 & ~n92051;
  assign n92087 = n92045 & n92086;
  assign n92088 = ~n92053 & ~n92087;
  assign n92089 = ~n92033 & ~n92088;
  assign n92090 = ~n92085 & ~n92089;
  assign n92091 = n92045 & n92063;
  assign n92092 = ~n92039 & n92091;
  assign n92093 = n92039 & n92069;
  assign n92094 = ~n92092 & ~n92093;
  assign n92095 = n92033 & n92039;
  assign n92096 = n92068 & n92095;
  assign n92097 = ~n92045 & n92071;
  assign n92098 = n92033 & n92097;
  assign n92099 = ~n92096 & ~n92098;
  assign n92100 = n92094 & n92099;
  assign n92101 = n92090 & n92100;
  assign n92102 = ~n92083 & n92101;
  assign n92103 = ~n92027 & ~n92102;
  assign n92104 = n92051 & ~n92059;
  assign n92105 = ~n92045 & n92104;
  assign n92106 = ~n92033 & n92105;
  assign n92107 = ~n92039 & n92106;
  assign n92108 = ~n92033 & n92092;
  assign n92109 = ~n92107 & ~n92108;
  assign n92110 = ~n92039 & ~n92045;
  assign n92111 = n92059 & n92110;
  assign n92112 = n92051 & n92111;
  assign n92113 = n92033 & n92112;
  assign n92114 = n92109 & ~n92113;
  assign n92115 = n92052 & ~n92059;
  assign n92116 = ~n92039 & n92115;
  assign n92117 = n92039 & n92060;
  assign n92118 = ~n92116 & ~n92117;
  assign n92119 = n92033 & ~n92118;
  assign n92120 = n92114 & ~n92119;
  assign n92121 = ~n92103 & n92120;
  assign n92122 = ~n92081 & n92121;
  assign n92123 = ~pi3192 & ~n92122;
  assign n92124 = pi3192 & n92122;
  assign po3103 = n92123 | n92124;
  assign n92126 = ~n91843 & n91864;
  assign n92127 = ~n91843 & n91906;
  assign n92128 = ~n92126 & ~n92127;
  assign n92129 = n91849 & n92128;
  assign n92130 = n91843 & n91901;
  assign n92131 = ~n91837 & ~n91858;
  assign n92132 = ~n91857 & ~n92131;
  assign n92133 = n91830 & n91888;
  assign n92134 = n91843 & n91858;
  assign n92135 = ~n92133 & ~n92134;
  assign n92136 = ~n91849 & n92135;
  assign n92137 = ~n92132 & n92136;
  assign n92138 = ~n92130 & n92137;
  assign n92139 = ~n92129 & ~n92138;
  assign n92140 = n91843 & n92132;
  assign n92141 = n91857 & n91864;
  assign n92142 = n91843 & n92141;
  assign n92143 = ~n92140 & ~n92142;
  assign n92144 = ~n92139 & n92143;
  assign n92145 = n91824 & ~n92144;
  assign n92146 = n91849 & ~n92131;
  assign n92147 = ~n91843 & n92146;
  assign n92148 = ~n91876 & ~n91905;
  assign n92149 = n91843 & ~n92148;
  assign n92150 = n91849 & n92149;
  assign n92151 = n91857 & n92146;
  assign n92152 = ~n92150 & ~n92151;
  assign n92153 = ~n92147 & n92152;
  assign n92154 = ~n91824 & ~n92153;
  assign n92155 = ~n92145 & ~n92154;
  assign n92156 = n91849 & n91862;
  assign n92157 = ~n91849 & ~n92143;
  assign n92158 = ~n92156 & ~n92157;
  assign n92159 = ~n91849 & ~n92128;
  assign n92160 = ~n91862 & ~n92159;
  assign n92161 = ~n91824 & ~n92160;
  assign n92162 = n92158 & ~n92161;
  assign n92163 = n92155 & n92162;
  assign n92164 = pi3242 & ~n92163;
  assign n92165 = ~pi3242 & n92162;
  assign n92166 = ~n92154 & n92165;
  assign n92167 = ~n92145 & n92166;
  assign po3108 = n92164 | n92167;
  assign n92169 = pi7063 & pi9040;
  assign n92170 = pi6878 & ~pi9040;
  assign n92171 = ~n92169 & ~n92170;
  assign n92172 = pi2941 & n92171;
  assign n92173 = ~pi2941 & ~n92171;
  assign n92174 = ~n92172 & ~n92173;
  assign n92175 = pi6879 & pi9040;
  assign n92176 = pi6989 & ~pi9040;
  assign n92177 = ~n92175 & ~n92176;
  assign n92178 = pi2975 & n92177;
  assign n92179 = ~pi2975 & ~n92177;
  assign n92180 = ~n92178 & ~n92179;
  assign n92181 = pi6878 & pi9040;
  assign n92182 = pi6909 & ~pi9040;
  assign n92183 = ~n92181 & ~n92182;
  assign n92184 = pi2947 & n92183;
  assign n92185 = ~pi2947 & ~n92183;
  assign n92186 = ~n92184 & ~n92185;
  assign n92187 = pi7048 & pi9040;
  assign n92188 = pi7080 & ~pi9040;
  assign n92189 = ~n92187 & ~n92188;
  assign n92190 = pi2966 & n92189;
  assign n92191 = ~pi2966 & ~n92189;
  assign n92192 = ~n92190 & ~n92191;
  assign n92193 = pi7020 & ~pi9040;
  assign n92194 = pi6915 & pi9040;
  assign n92195 = ~n92193 & ~n92194;
  assign n92196 = pi2954 & n92195;
  assign n92197 = ~pi2954 & ~n92195;
  assign n92198 = ~n92196 & ~n92197;
  assign n92199 = ~n92192 & n92198;
  assign n92200 = ~n92186 & n92199;
  assign n92201 = ~n92180 & n92200;
  assign n92202 = n92186 & ~n92198;
  assign n92203 = n92192 & n92202;
  assign n92204 = n92180 & n92203;
  assign n92205 = ~n92192 & ~n92198;
  assign n92206 = ~n92186 & n92205;
  assign n92207 = n92180 & n92206;
  assign n92208 = ~n92204 & ~n92207;
  assign n92209 = ~n92201 & n92208;
  assign n92210 = n92174 & ~n92209;
  assign n92211 = ~n92180 & n92186;
  assign n92212 = n92198 & n92211;
  assign n92213 = n92192 & n92212;
  assign n92214 = pi6889 & pi9040;
  assign n92215 = ~pi6868 & ~pi9040;
  assign n92216 = ~n92214 & ~n92215;
  assign n92217 = ~pi2962 & ~n92216;
  assign n92218 = pi2962 & n92216;
  assign n92219 = ~n92217 & ~n92218;
  assign n92220 = ~n92192 & n92211;
  assign n92221 = n92192 & n92198;
  assign n92222 = ~n92186 & n92221;
  assign n92223 = ~n92220 & ~n92222;
  assign n92224 = ~n92174 & ~n92223;
  assign n92225 = ~n92212 & ~n92224;
  assign n92226 = n92186 & n92221;
  assign n92227 = ~n92186 & ~n92198;
  assign n92228 = ~n92180 & n92227;
  assign n92229 = n92180 & n92205;
  assign n92230 = ~n92228 & ~n92229;
  assign n92231 = ~n92186 & ~n92192;
  assign n92232 = n92230 & ~n92231;
  assign n92233 = ~n92226 & n92232;
  assign n92234 = n92174 & ~n92233;
  assign n92235 = n92225 & ~n92234;
  assign n92236 = ~n92204 & n92235;
  assign n92237 = n92219 & ~n92236;
  assign n92238 = ~n92213 & ~n92237;
  assign n92239 = ~n92210 & n92238;
  assign n92240 = ~n92186 & n92192;
  assign n92241 = ~n92174 & n92240;
  assign n92242 = n92180 & n92241;
  assign n92243 = n92174 & ~n92180;
  assign n92244 = n92186 & n92243;
  assign n92245 = ~n92198 & n92244;
  assign n92246 = n92186 & n92199;
  assign n92247 = n92180 & n92246;
  assign n92248 = ~n92245 & ~n92247;
  assign n92249 = n92186 & ~n92192;
  assign n92250 = n92180 & n92249;
  assign n92251 = n92192 & ~n92198;
  assign n92252 = ~n92186 & n92251;
  assign n92253 = ~n92250 & ~n92252;
  assign n92254 = ~n92174 & ~n92253;
  assign n92255 = ~n92174 & ~n92192;
  assign n92256 = ~n92186 & n92255;
  assign n92257 = ~n92180 & n92256;
  assign n92258 = ~n92254 & ~n92257;
  assign n92259 = n92248 & n92258;
  assign n92260 = ~n92219 & ~n92259;
  assign n92261 = ~n92242 & ~n92260;
  assign n92262 = n92239 & n92261;
  assign n92263 = pi3186 & n92262;
  assign n92264 = ~n92213 & ~n92242;
  assign n92265 = ~n92260 & n92264;
  assign n92266 = ~n92210 & ~n92237;
  assign n92267 = n92265 & n92266;
  assign n92268 = ~pi3186 & ~n92267;
  assign po3109 = n92263 | n92268;
  assign n92270 = n91843 & n91871;
  assign n92271 = ~n91890 & ~n91899;
  assign n92272 = n91849 & ~n92271;
  assign n92273 = ~n92270 & ~n92272;
  assign n92274 = ~n91884 & n92273;
  assign n92275 = ~n91849 & n91887;
  assign n92276 = ~n91879 & ~n92275;
  assign n92277 = ~n91907 & n92276;
  assign n92278 = n92274 & n92277;
  assign n92279 = n91824 & ~n92278;
  assign n92280 = ~n91862 & ~n92142;
  assign n92281 = ~n91872 & ~n92127;
  assign n92282 = n91837 & n91857;
  assign n92283 = n91849 & n92282;
  assign n92284 = n91843 & n91878;
  assign n92285 = ~n92283 & ~n92284;
  assign n92286 = n91836 & ~n91857;
  assign n92287 = ~n91830 & n91843;
  assign n92288 = ~n92286 & ~n92287;
  assign n92289 = ~n91912 & n92288;
  assign n92290 = ~n91849 & ~n92289;
  assign n92291 = n92285 & ~n92290;
  assign n92292 = n92281 & n92291;
  assign n92293 = n92280 & n92292;
  assign n92294 = ~n91824 & ~n92293;
  assign n92295 = ~n92279 & ~n92294;
  assign n92296 = pi3185 & ~n92295;
  assign n92297 = ~pi3185 & ~n92294;
  assign n92298 = ~n92279 & n92297;
  assign po3110 = n92296 | n92298;
  assign n92300 = pi7098 & pi9040;
  assign n92301 = pi6861 & ~pi9040;
  assign n92302 = ~n92300 & ~n92301;
  assign n92303 = ~pi2946 & ~n92302;
  assign n92304 = pi2946 & n92302;
  assign n92305 = ~n92303 & ~n92304;
  assign n92306 = pi7000 & pi9040;
  assign n92307 = pi7073 & ~pi9040;
  assign n92308 = ~n92306 & ~n92307;
  assign n92309 = pi2974 & n92308;
  assign n92310 = ~pi2974 & ~n92308;
  assign n92311 = ~n92309 & ~n92310;
  assign n92312 = pi6997 & ~pi9040;
  assign n92313 = pi6977 & pi9040;
  assign n92314 = ~n92312 & ~n92313;
  assign n92315 = pi2972 & n92314;
  assign n92316 = ~pi2972 & ~n92314;
  assign n92317 = ~n92315 & ~n92316;
  assign n92318 = pi7098 & ~pi9040;
  assign n92319 = pi6995 & pi9040;
  assign n92320 = ~n92318 & ~n92319;
  assign n92321 = ~pi2967 & n92320;
  assign n92322 = pi2967 & ~n92320;
  assign n92323 = ~n92321 & ~n92322;
  assign n92324 = n92317 & n92323;
  assign n92325 = pi7073 & pi9040;
  assign n92326 = pi6963 & ~pi9040;
  assign n92327 = ~n92325 & ~n92326;
  assign n92328 = pi2968 & n92327;
  assign n92329 = ~pi2968 & ~n92327;
  assign n92330 = ~n92328 & ~n92329;
  assign n92331 = pi6964 & ~pi9040;
  assign n92332 = pi7167 & pi9040;
  assign n92333 = ~n92331 & ~n92332;
  assign n92334 = ~pi2930 & n92333;
  assign n92335 = pi2930 & ~n92333;
  assign n92336 = ~n92334 & ~n92335;
  assign n92337 = ~n92323 & ~n92336;
  assign n92338 = ~n92330 & n92337;
  assign n92339 = ~n92317 & n92338;
  assign n92340 = ~n92324 & ~n92339;
  assign n92341 = n92323 & n92330;
  assign n92342 = n92340 & ~n92341;
  assign n92343 = n92311 & ~n92342;
  assign n92344 = ~n92311 & n92330;
  assign n92345 = ~n92323 & n92344;
  assign n92346 = n92317 & n92330;
  assign n92347 = ~n92336 & n92346;
  assign n92348 = ~n92323 & n92336;
  assign n92349 = n92317 & n92348;
  assign n92350 = ~n92330 & n92349;
  assign n92351 = ~n92347 & ~n92350;
  assign n92352 = ~n92317 & n92323;
  assign n92353 = ~n92311 & ~n92330;
  assign n92354 = n92352 & n92353;
  assign n92355 = n92351 & ~n92354;
  assign n92356 = ~n92345 & n92355;
  assign n92357 = ~n92343 & n92356;
  assign n92358 = n92305 & ~n92357;
  assign n92359 = n92323 & ~n92336;
  assign n92360 = n92317 & n92359;
  assign n92361 = ~n92330 & n92360;
  assign n92362 = n92323 & n92336;
  assign n92363 = n92317 & n92362;
  assign n92364 = n92330 & n92363;
  assign n92365 = ~n92361 & ~n92364;
  assign n92366 = n92311 & ~n92365;
  assign n92367 = ~n92358 & ~n92366;
  assign n92368 = n92330 & n92349;
  assign n92369 = n92317 & ~n92323;
  assign n92370 = ~n92336 & n92369;
  assign n92371 = ~n92317 & n92336;
  assign n92372 = ~n92323 & n92371;
  assign n92373 = ~n92370 & ~n92372;
  assign n92374 = n92311 & ~n92373;
  assign n92375 = ~n92368 & ~n92374;
  assign n92376 = ~n92317 & n92359;
  assign n92377 = n92330 & n92376;
  assign n92378 = n92375 & ~n92377;
  assign n92379 = ~n92305 & ~n92378;
  assign n92380 = ~n92337 & ~n92362;
  assign n92381 = ~n92317 & ~n92380;
  assign n92382 = ~n92330 & n92362;
  assign n92383 = ~n92381 & ~n92382;
  assign n92384 = ~n92311 & ~n92383;
  assign n92385 = ~n92305 & n92384;
  assign n92386 = ~n92379 & ~n92385;
  assign n92387 = n92367 & n92386;
  assign n92388 = ~pi3244 & n92387;
  assign n92389 = pi3244 & ~n92387;
  assign po3111 = n92388 | n92389;
  assign n92391 = n92311 & n92330;
  assign n92392 = n92359 & n92391;
  assign n92393 = n92317 & n92392;
  assign n92394 = n92311 & ~n92330;
  assign n92395 = n92337 & n92394;
  assign n92396 = n92317 & ~n92330;
  assign n92397 = n92336 & n92396;
  assign n92398 = n92323 & n92397;
  assign n92399 = n92311 & n92349;
  assign n92400 = n92330 & n92399;
  assign n92401 = ~n92398 & ~n92400;
  assign n92402 = ~n92395 & n92401;
  assign n92403 = ~n92393 & n92402;
  assign n92404 = ~n92339 & n92403;
  assign n92405 = ~n92305 & ~n92404;
  assign n92406 = ~n92311 & n92372;
  assign n92407 = n92330 & n92406;
  assign n92408 = n92323 & n92396;
  assign n92409 = ~n92382 & ~n92408;
  assign n92410 = ~n92311 & ~n92409;
  assign n92411 = ~n92407 & ~n92410;
  assign n92412 = ~n92305 & ~n92411;
  assign n92413 = n92330 & n92370;
  assign n92414 = ~n92397 & ~n92413;
  assign n92415 = ~n92377 & n92414;
  assign n92416 = ~n92311 & ~n92415;
  assign n92417 = ~n92412 & ~n92416;
  assign n92418 = ~n92405 & n92417;
  assign n92419 = ~n92317 & n92330;
  assign n92420 = n92311 & n92419;
  assign n92421 = n92362 & n92420;
  assign n92422 = ~n92317 & n92394;
  assign n92423 = ~n92323 & n92422;
  assign n92424 = ~n92330 & n92372;
  assign n92425 = ~n92311 & n92317;
  assign n92426 = ~n92323 & n92425;
  assign n92427 = ~n92317 & n92341;
  assign n92428 = ~n92426 & ~n92427;
  assign n92429 = ~n92424 & n92428;
  assign n92430 = ~n92376 & n92429;
  assign n92431 = n92311 & n92359;
  assign n92432 = ~n92330 & n92431;
  assign n92433 = n92330 & n92362;
  assign n92434 = ~n92317 & ~n92336;
  assign n92435 = ~n92433 & ~n92434;
  assign n92436 = n92311 & ~n92435;
  assign n92437 = ~n92432 & ~n92436;
  assign n92438 = n92430 & n92437;
  assign n92439 = n92305 & ~n92438;
  assign n92440 = ~n92423 & ~n92439;
  assign n92441 = ~n92421 & n92440;
  assign n92442 = n92418 & n92441;
  assign n92443 = pi3190 & n92442;
  assign n92444 = ~pi3190 & ~n92442;
  assign po3112 = n92443 | n92444;
  assign n92446 = ~pi6885 & ~pi9040;
  assign n92447 = pi6918 & pi9040;
  assign n92448 = ~n92446 & ~n92447;
  assign n92449 = ~pi2966 & n92448;
  assign n92450 = pi2966 & ~n92448;
  assign n92451 = ~n92449 & ~n92450;
  assign n92452 = pi6995 & ~pi9040;
  assign n92453 = pi7022 & pi9040;
  assign n92454 = ~n92452 & ~n92453;
  assign n92455 = ~pi2964 & n92454;
  assign n92456 = pi2964 & ~n92454;
  assign n92457 = ~n92455 & ~n92456;
  assign n92458 = pi6911 & ~pi9040;
  assign n92459 = pi7025 & pi9040;
  assign n92460 = ~n92458 & ~n92459;
  assign n92461 = pi2973 & n92460;
  assign n92462 = ~pi2973 & ~n92460;
  assign n92463 = ~n92461 & ~n92462;
  assign n92464 = pi7134 & ~pi9040;
  assign n92465 = pi6861 & pi9040;
  assign n92466 = ~n92464 & ~n92465;
  assign n92467 = pi2944 & n92466;
  assign n92468 = ~pi2944 & ~n92466;
  assign n92469 = ~n92467 & ~n92468;
  assign n92470 = pi7010 & pi9040;
  assign n92471 = pi6977 & ~pi9040;
  assign n92472 = ~n92470 & ~n92471;
  assign n92473 = ~pi2947 & n92472;
  assign n92474 = pi2947 & ~n92472;
  assign n92475 = ~n92473 & ~n92474;
  assign n92476 = ~n92469 & ~n92475;
  assign n92477 = n92463 & n92476;
  assign n92478 = ~n92457 & n92477;
  assign n92479 = pi6964 & pi9040;
  assign n92480 = pi7025 & ~pi9040;
  assign n92481 = ~n92479 & ~n92480;
  assign n92482 = ~pi2963 & ~n92481;
  assign n92483 = pi2963 & n92481;
  assign n92484 = ~n92482 & ~n92483;
  assign n92485 = ~pi2944 & n92466;
  assign n92486 = pi2944 & ~n92466;
  assign n92487 = ~n92485 & ~n92486;
  assign n92488 = ~n92475 & ~n92487;
  assign n92489 = ~n92457 & n92488;
  assign n92490 = ~n92463 & n92476;
  assign n92491 = n92457 & n92490;
  assign n92492 = ~n92489 & ~n92491;
  assign n92493 = ~n92484 & ~n92492;
  assign n92494 = ~n92478 & ~n92493;
  assign n92495 = ~n92469 & n92475;
  assign n92496 = ~n92463 & n92495;
  assign n92497 = n92484 & n92496;
  assign n92498 = n92476 & n92484;
  assign n92499 = ~n92457 & n92498;
  assign n92500 = ~n92497 & ~n92499;
  assign n92501 = n92494 & n92500;
  assign n92502 = n92475 & ~n92487;
  assign n92503 = n92463 & n92502;
  assign n92504 = ~n92457 & n92503;
  assign n92505 = n92463 & n92495;
  assign n92506 = n92457 & n92505;
  assign n92507 = ~n92504 & ~n92506;
  assign n92508 = n92501 & n92507;
  assign n92509 = n92451 & ~n92508;
  assign n92510 = ~n92451 & ~n92484;
  assign n92511 = ~n92457 & ~n92463;
  assign n92512 = n92487 & n92511;
  assign n92513 = ~n92463 & n92475;
  assign n92514 = ~n92512 & ~n92513;
  assign n92515 = n92510 & ~n92514;
  assign n92516 = n92457 & n92463;
  assign n92517 = ~n92475 & n92516;
  assign n92518 = ~n92469 & n92517;
  assign n92519 = n92457 & ~n92487;
  assign n92520 = ~n92463 & n92519;
  assign n92521 = ~n92518 & ~n92520;
  assign n92522 = ~n92457 & n92484;
  assign n92523 = n92463 & n92522;
  assign n92524 = ~n92476 & n92523;
  assign n92525 = n92484 & n92503;
  assign n92526 = ~n92524 & ~n92525;
  assign n92527 = n92521 & n92526;
  assign n92528 = ~n92451 & ~n92527;
  assign n92529 = ~n92463 & n92502;
  assign n92530 = ~n92484 & n92529;
  assign n92531 = n92457 & n92530;
  assign n92532 = n92463 & n92488;
  assign n92533 = n92457 & n92532;
  assign n92534 = ~n92506 & ~n92533;
  assign n92535 = ~n92484 & ~n92534;
  assign n92536 = ~n92531 & ~n92535;
  assign n92537 = n92484 & n92518;
  assign n92538 = n92536 & ~n92537;
  assign n92539 = ~n92528 & n92538;
  assign n92540 = ~n92515 & n92539;
  assign n92541 = ~n92509 & n92540;
  assign n92542 = ~n92463 & n92488;
  assign n92543 = n92457 & n92484;
  assign n92544 = n92542 & n92543;
  assign n92545 = n92541 & ~n92544;
  assign n92546 = ~pi3237 & ~n92545;
  assign n92547 = ~n92509 & ~n92544;
  assign n92548 = n92540 & n92547;
  assign n92549 = pi3237 & n92548;
  assign po3115 = n92546 | n92549;
  assign n92551 = n92186 & n92205;
  assign n92552 = ~n92180 & n92551;
  assign n92553 = ~n92200 & ~n92213;
  assign n92554 = n92180 & n92202;
  assign n92555 = ~n92180 & n92252;
  assign n92556 = ~n92554 & ~n92555;
  assign n92557 = n92553 & n92556;
  assign n92558 = ~n92174 & ~n92557;
  assign n92559 = n92180 & n92221;
  assign n92560 = ~n92220 & ~n92559;
  assign n92561 = ~n92206 & n92560;
  assign n92562 = n92174 & ~n92561;
  assign n92563 = n92180 & n92222;
  assign n92564 = ~n92562 & ~n92563;
  assign n92565 = ~n92558 & n92564;
  assign n92566 = ~n92552 & n92565;
  assign n92567 = ~n92219 & ~n92566;
  assign n92568 = ~n92174 & n92180;
  assign n92569 = n92226 & n92568;
  assign n92570 = ~n92174 & n92206;
  assign n92571 = ~n92174 & n92246;
  assign n92572 = ~n92570 & ~n92571;
  assign n92573 = ~n92180 & ~n92572;
  assign n92574 = ~n92569 & ~n92573;
  assign n92575 = ~n92180 & n92203;
  assign n92576 = n92180 & n92252;
  assign n92577 = ~n92575 & ~n92576;
  assign n92578 = n92180 & n92199;
  assign n92579 = ~n92180 & n92221;
  assign n92580 = ~n92578 & ~n92579;
  assign n92581 = ~n92203 & n92580;
  assign n92582 = ~n92200 & n92581;
  assign n92583 = n92174 & ~n92582;
  assign n92584 = ~n92180 & n92222;
  assign n92585 = ~n92583 & ~n92584;
  assign n92586 = n92577 & n92585;
  assign n92587 = n92574 & n92586;
  assign n92588 = n92219 & ~n92587;
  assign n92589 = n92180 & n92551;
  assign n92590 = n92180 & n92200;
  assign n92591 = ~n92589 & ~n92590;
  assign n92592 = ~n92174 & ~n92591;
  assign n92593 = ~n92588 & ~n92592;
  assign n92594 = ~n92207 & ~n92575;
  assign n92595 = n92174 & ~n92594;
  assign n92596 = n92593 & ~n92595;
  assign n92597 = ~n92567 & n92596;
  assign n92598 = pi3261 & ~n92597;
  assign n92599 = ~pi3261 & n92597;
  assign po3116 = n92598 | n92599;
  assign n92601 = ~n92027 & ~n92033;
  assign n92602 = ~n92039 & n92052;
  assign n92603 = n92039 & n92091;
  assign n92604 = ~n92039 & n92060;
  assign n92605 = ~n92603 & ~n92604;
  assign n92606 = ~n92602 & n92605;
  assign n92607 = n92601 & ~n92606;
  assign n92608 = ~n92059 & n92110;
  assign n92609 = n92039 & n92115;
  assign n92610 = ~n92608 & ~n92609;
  assign n92611 = ~n92061 & ~n92064;
  assign n92612 = n92610 & n92611;
  assign n92613 = n92033 & ~n92612;
  assign n92614 = n92039 & n92097;
  assign n92615 = ~n92613 & ~n92614;
  assign n92616 = ~n92027 & ~n92615;
  assign n92617 = ~n92607 & ~n92616;
  assign n92618 = n92045 & n92082;
  assign n92619 = n92059 & n92618;
  assign n92620 = ~n92065 & ~n92619;
  assign n92621 = ~n92060 & ~n92104;
  assign n92622 = n92039 & ~n92621;
  assign n92623 = ~n92105 & ~n92622;
  assign n92624 = ~n92033 & ~n92623;
  assign n92625 = ~n92072 & ~n92602;
  assign n92626 = ~n92603 & n92625;
  assign n92627 = n92033 & ~n92626;
  assign n92628 = ~n92624 & ~n92627;
  assign n92629 = n92039 & ~n92045;
  assign n92630 = ~n92059 & n92629;
  assign n92631 = n92051 & n92630;
  assign n92632 = ~n92093 & ~n92631;
  assign n92633 = ~n92112 & n92632;
  assign n92634 = ~n92085 & n92633;
  assign n92635 = n92628 & n92634;
  assign n92636 = n92027 & ~n92635;
  assign n92637 = n92620 & ~n92636;
  assign n92638 = n92617 & n92637;
  assign n92639 = pi3193 & ~n92638;
  assign n92640 = ~pi3193 & n92620;
  assign n92641 = n92617 & n92640;
  assign n92642 = ~n92636 & n92641;
  assign po3117 = n92639 | n92642;
  assign n92644 = pi7001 & pi9040;
  assign n92645 = pi6905 & ~pi9040;
  assign n92646 = ~n92644 & ~n92645;
  assign n92647 = ~pi2952 & ~n92646;
  assign n92648 = pi2952 & n92646;
  assign n92649 = ~n92647 & ~n92648;
  assign n92650 = pi7134 & pi9040;
  assign n92651 = pi6937 & ~pi9040;
  assign n92652 = ~n92650 & ~n92651;
  assign n92653 = ~pi2946 & ~n92652;
  assign n92654 = pi2946 & n92652;
  assign n92655 = ~n92653 & ~n92654;
  assign n92656 = pi6970 & pi9040;
  assign n92657 = pi6897 & ~pi9040;
  assign n92658 = ~n92656 & ~n92657;
  assign n92659 = pi2960 & n92658;
  assign n92660 = ~pi2960 & ~n92658;
  assign n92661 = ~n92659 & ~n92660;
  assign n92662 = n92655 & ~n92661;
  assign n92663 = pi6991 & pi9040;
  assign n92664 = pi7010 & ~pi9040;
  assign n92665 = ~n92663 & ~n92664;
  assign n92666 = ~pi2971 & ~n92665;
  assign n92667 = pi2971 & n92665;
  assign n92668 = ~n92666 & ~n92667;
  assign n92669 = pi6991 & ~pi9040;
  assign n92670 = pi6885 & pi9040;
  assign n92671 = ~n92669 & ~n92670;
  assign n92672 = ~pi2930 & n92671;
  assign n92673 = pi2930 & ~n92671;
  assign n92674 = ~n92672 & ~n92673;
  assign n92675 = n92668 & ~n92674;
  assign n92676 = n92662 & n92675;
  assign n92677 = ~pi2930 & ~n92671;
  assign n92678 = pi2930 & n92671;
  assign n92679 = ~n92677 & ~n92678;
  assign n92680 = n92655 & n92661;
  assign n92681 = ~n92679 & n92680;
  assign n92682 = ~n92655 & ~n92661;
  assign n92683 = n92674 & n92682;
  assign n92684 = ~n92681 & ~n92683;
  assign n92685 = n92668 & ~n92684;
  assign n92686 = ~n92676 & ~n92685;
  assign n92687 = ~n92649 & ~n92686;
  assign n92688 = ~n92668 & n92682;
  assign n92689 = ~n92655 & n92661;
  assign n92690 = ~n92674 & n92689;
  assign n92691 = ~n92688 & ~n92690;
  assign n92692 = pi7001 & ~pi9040;
  assign n92693 = pi6917 & pi9040;
  assign n92694 = ~n92692 & ~n92693;
  assign n92695 = pi2959 & n92694;
  assign n92696 = ~pi2959 & ~n92694;
  assign n92697 = ~n92695 & ~n92696;
  assign n92698 = ~n92649 & n92697;
  assign n92699 = ~n92691 & n92698;
  assign n92700 = ~n92687 & ~n92699;
  assign n92701 = n92668 & ~n92679;
  assign n92702 = ~n92655 & n92701;
  assign n92703 = ~n92676 & ~n92702;
  assign n92704 = ~n92697 & ~n92703;
  assign n92705 = ~n92668 & n92697;
  assign n92706 = n92655 & n92705;
  assign n92707 = n92662 & ~n92679;
  assign n92708 = ~n92674 & n92680;
  assign n92709 = ~n92707 & ~n92708;
  assign n92710 = n92679 & n92682;
  assign n92711 = n92668 & n92710;
  assign n92712 = n92709 & ~n92711;
  assign n92713 = n92697 & ~n92712;
  assign n92714 = ~n92706 & ~n92713;
  assign n92715 = n92674 & n92689;
  assign n92716 = n92668 & n92715;
  assign n92717 = n92714 & ~n92716;
  assign n92718 = ~n92691 & ~n92697;
  assign n92719 = ~n92668 & n92681;
  assign n92720 = ~n92718 & ~n92719;
  assign n92721 = n92717 & n92720;
  assign n92722 = n92649 & ~n92721;
  assign n92723 = ~n92704 & ~n92722;
  assign n92724 = ~n92649 & ~n92697;
  assign n92725 = n92662 & ~n92668;
  assign n92726 = ~n92715 & ~n92725;
  assign n92727 = n92655 & ~n92674;
  assign n92728 = n92726 & ~n92727;
  assign n92729 = n92724 & ~n92728;
  assign n92730 = n92723 & ~n92729;
  assign n92731 = n92700 & n92730;
  assign n92732 = ~pi3187 & ~n92731;
  assign n92733 = pi3187 & n92700;
  assign n92734 = n92723 & n92733;
  assign n92735 = ~n92729 & n92734;
  assign po3118 = n92732 | n92735;
  assign n92737 = ~n92174 & ~n92180;
  assign n92738 = n92192 & n92737;
  assign n92739 = ~n92180 & ~n92186;
  assign n92740 = ~n92198 & n92739;
  assign n92741 = ~n92192 & n92740;
  assign n92742 = ~n92222 & ~n92741;
  assign n92743 = n92174 & ~n92742;
  assign n92744 = n92591 & ~n92743;
  assign n92745 = ~n92738 & n92744;
  assign n92746 = n92219 & ~n92745;
  assign n92747 = ~n92174 & n92576;
  assign n92748 = n92243 & n92252;
  assign n92749 = ~n92220 & ~n92748;
  assign n92750 = ~n92222 & ~n92246;
  assign n92751 = ~n92180 & n92199;
  assign n92752 = n92750 & ~n92751;
  assign n92753 = ~n92174 & ~n92752;
  assign n92754 = n92174 & n92226;
  assign n92755 = n92208 & ~n92754;
  assign n92756 = ~n92753 & n92755;
  assign n92757 = n92749 & n92756;
  assign n92758 = ~n92219 & ~n92757;
  assign n92759 = ~n92747 & ~n92758;
  assign n92760 = ~n92746 & n92759;
  assign n92761 = n92243 & n92246;
  assign n92762 = n92174 & n92202;
  assign n92763 = n92180 & n92762;
  assign n92764 = ~n92761 & ~n92763;
  assign n92765 = n92174 & n92590;
  assign n92766 = n92764 & ~n92765;
  assign n92767 = n92760 & n92766;
  assign n92768 = ~pi3241 & ~n92767;
  assign n92769 = pi3241 & n92766;
  assign n92770 = n92759 & n92769;
  assign n92771 = ~n92746 & n92770;
  assign po3120 = n92768 | n92771;
  assign n92773 = ~n91843 & n91858;
  assign n92774 = ~n92141 & ~n92773;
  assign n92775 = n91849 & ~n92774;
  assign n92776 = ~n91907 & ~n92775;
  assign n92777 = n91843 & n92282;
  assign n92778 = ~n91877 & ~n92777;
  assign n92779 = n91843 & n91912;
  assign n92780 = ~n92286 & ~n92779;
  assign n92781 = n91857 & n91905;
  assign n92782 = n92780 & ~n92781;
  assign n92783 = ~n91849 & ~n92782;
  assign n92784 = ~n91843 & n91859;
  assign n92785 = ~n92783 & ~n92784;
  assign n92786 = n92778 & n92785;
  assign n92787 = n92776 & n92786;
  assign n92788 = ~n91824 & ~n92787;
  assign n92789 = ~n91893 & ~n92130;
  assign n92790 = ~n91849 & ~n92789;
  assign n92791 = ~n92788 & ~n92790;
  assign n92792 = n91849 & n92777;
  assign n92793 = n91888 & ~n92131;
  assign n92794 = ~n91906 & ~n92142;
  assign n92795 = ~n92793 & n92794;
  assign n92796 = ~n91849 & ~n92795;
  assign n92797 = n91843 & n91859;
  assign n92798 = ~n92796 & ~n92797;
  assign n92799 = ~n91843 & n92286;
  assign n92800 = ~n92781 & ~n92799;
  assign n92801 = ~n92134 & n92800;
  assign n92802 = n91849 & ~n92801;
  assign n92803 = n92798 & ~n92802;
  assign n92804 = n91824 & ~n92803;
  assign n92805 = ~n92792 & ~n92804;
  assign n92806 = n92791 & n92805;
  assign n92807 = pi3249 & n92806;
  assign n92808 = ~pi3249 & ~n92806;
  assign po3121 = n92807 | n92808;
  assign n92810 = n92668 & ~n92697;
  assign n92811 = ~n92681 & ~n92682;
  assign n92812 = n92810 & ~n92811;
  assign n92813 = ~n92679 & ~n92697;
  assign n92814 = n92682 & n92813;
  assign n92815 = ~n92812 & ~n92814;
  assign n92816 = n92649 & ~n92815;
  assign n92817 = ~n92668 & n92708;
  assign n92818 = ~n92668 & ~n92674;
  assign n92819 = ~n92727 & ~n92818;
  assign n92820 = n92697 & ~n92819;
  assign n92821 = ~n92668 & ~n92679;
  assign n92822 = ~n92661 & n92821;
  assign n92823 = n92655 & n92822;
  assign n92824 = ~n92820 & ~n92823;
  assign n92825 = ~n92817 & n92824;
  assign n92826 = n92649 & ~n92825;
  assign n92827 = ~n92816 & ~n92826;
  assign n92828 = n92661 & n92675;
  assign n92829 = ~n92655 & n92828;
  assign n92830 = ~n92668 & n92715;
  assign n92831 = ~n92829 & ~n92830;
  assign n92832 = ~n92697 & ~n92831;
  assign n92833 = n92661 & ~n92668;
  assign n92834 = n92674 & ~n92697;
  assign n92835 = n92833 & n92834;
  assign n92836 = ~n92662 & ~n92727;
  assign n92837 = n92668 & ~n92836;
  assign n92838 = ~n92715 & ~n92837;
  assign n92839 = ~n92697 & ~n92838;
  assign n92840 = ~n92661 & n92679;
  assign n92841 = ~n92715 & ~n92840;
  assign n92842 = ~n92668 & ~n92841;
  assign n92843 = n92668 & n92697;
  assign n92844 = n92680 & n92843;
  assign n92845 = ~n92679 & n92844;
  assign n92846 = ~n92842 & ~n92845;
  assign n92847 = ~n92839 & n92846;
  assign n92848 = ~n92835 & n92847;
  assign n92849 = ~n92829 & n92848;
  assign n92850 = ~n92649 & ~n92849;
  assign n92851 = n92668 & n92683;
  assign n92852 = ~n92668 & n92727;
  assign n92853 = ~n92851 & ~n92852;
  assign n92854 = n92697 & ~n92853;
  assign n92855 = ~n92850 & ~n92854;
  assign n92856 = ~n92832 & n92855;
  assign n92857 = n92827 & n92856;
  assign n92858 = pi3243 & n92857;
  assign n92859 = ~pi3243 & ~n92857;
  assign po3122 = n92858 | n92859;
  assign n92861 = ~n92330 & n92376;
  assign n92862 = ~n92350 & ~n92861;
  assign n92863 = ~n92311 & ~n92862;
  assign n92864 = n92344 & n92370;
  assign n92865 = ~n92863 & ~n92864;
  assign n92866 = ~n92423 & n92865;
  assign n92867 = n92311 & n92317;
  assign n92868 = n92336 & n92867;
  assign n92869 = n92323 & n92868;
  assign n92870 = ~n92330 & n92869;
  assign n92871 = n92311 & n92360;
  assign n92872 = ~n92339 & ~n92421;
  assign n92873 = ~n92400 & n92872;
  assign n92874 = ~n92871 & n92873;
  assign n92875 = n92305 & ~n92874;
  assign n92876 = n92330 & n92372;
  assign n92877 = ~n92376 & ~n92876;
  assign n92878 = ~n92363 & n92877;
  assign n92879 = ~n92311 & ~n92878;
  assign n92880 = n92305 & n92879;
  assign n92881 = n92330 & n92431;
  assign n92882 = ~n92869 & ~n92881;
  assign n92883 = ~n92347 & n92882;
  assign n92884 = ~n92317 & ~n92330;
  assign n92885 = n92336 & n92884;
  assign n92886 = n92330 & n92337;
  assign n92887 = ~n92369 & ~n92886;
  assign n92888 = ~n92311 & ~n92887;
  assign n92889 = ~n92885 & ~n92888;
  assign n92890 = n92883 & n92889;
  assign n92891 = ~n92305 & ~n92890;
  assign n92892 = ~n92880 & ~n92891;
  assign n92893 = ~n92875 & n92892;
  assign n92894 = ~n92870 & n92893;
  assign n92895 = n92866 & n92894;
  assign n92896 = pi3260 & ~n92895;
  assign n92897 = ~pi3260 & n92866;
  assign n92898 = n92894 & n92897;
  assign po3124 = n92896 | n92898;
  assign n92900 = n92330 & n92381;
  assign n92901 = ~n92360 & ~n92371;
  assign n92902 = ~n92311 & ~n92901;
  assign n92903 = ~n92900 & ~n92902;
  assign n92904 = n92336 & n92346;
  assign n92905 = ~n92434 & ~n92904;
  assign n92906 = ~n92363 & n92905;
  assign n92907 = n92311 & ~n92906;
  assign n92908 = n92903 & ~n92907;
  assign n92909 = ~n92330 & n92370;
  assign n92910 = n92908 & ~n92909;
  assign n92911 = ~n92305 & ~n92910;
  assign n92912 = ~n92372 & ~n92376;
  assign n92913 = ~n92363 & ~n92370;
  assign n92914 = n92912 & n92913;
  assign n92915 = n92330 & ~n92914;
  assign n92916 = n92394 & ~n92901;
  assign n92917 = ~n92915 & ~n92916;
  assign n92918 = ~n92350 & n92917;
  assign n92919 = n92305 & ~n92918;
  assign n92920 = ~n92911 & ~n92919;
  assign n92921 = n92330 & n92360;
  assign n92922 = ~n92909 & ~n92921;
  assign n92923 = ~n92311 & ~n92922;
  assign n92924 = n92920 & ~n92923;
  assign n92925 = pi3245 & ~n92924;
  assign n92926 = ~pi3245 & ~n92923;
  assign n92927 = ~n92919 & n92926;
  assign n92928 = ~n92911 & n92927;
  assign po3125 = n92925 | n92928;
  assign n92930 = ~n92575 & ~n92741;
  assign n92931 = ~n92563 & n92930;
  assign n92932 = ~n92174 & ~n92931;
  assign n92933 = ~n92571 & ~n92576;
  assign n92934 = ~n92551 & ~n92579;
  assign n92935 = n92174 & ~n92934;
  assign n92936 = ~n92213 & ~n92935;
  assign n92937 = n92933 & n92936;
  assign n92938 = n92219 & ~n92937;
  assign n92939 = ~n92186 & n92198;
  assign n92940 = ~n92231 & ~n92939;
  assign n92941 = n92180 & ~n92940;
  assign n92942 = ~n92203 & ~n92751;
  assign n92943 = n92174 & ~n92942;
  assign n92944 = n92180 & n92198;
  assign n92945 = ~n92222 & ~n92944;
  assign n92946 = ~n92205 & n92945;
  assign n92947 = ~n92174 & ~n92946;
  assign n92948 = ~n92943 & ~n92947;
  assign n92949 = ~n92941 & n92948;
  assign n92950 = ~n92219 & ~n92949;
  assign n92951 = ~n92938 & ~n92950;
  assign n92952 = ~n92748 & ~n92765;
  assign n92953 = n92951 & n92952;
  assign n92954 = ~n92932 & n92953;
  assign n92955 = ~pi3328 & ~n92954;
  assign n92956 = pi3328 & n92952;
  assign n92957 = ~n92932 & n92956;
  assign n92958 = n92951 & n92957;
  assign po3126 = n92955 | n92958;
  assign n92960 = n92033 & n92060;
  assign n92961 = ~n92039 & n92960;
  assign n92962 = ~n92116 & ~n92961;
  assign n92963 = n92039 & n92059;
  assign n92964 = n92045 & n92963;
  assign n92965 = ~n92039 & n92045;
  assign n92966 = ~n92059 & n92965;
  assign n92967 = ~n92039 & n92051;
  assign n92968 = ~n92966 & ~n92967;
  assign n92969 = ~n92033 & ~n92968;
  assign n92970 = ~n92964 & ~n92969;
  assign n92971 = n92962 & n92970;
  assign n92972 = n92027 & ~n92971;
  assign n92973 = ~n92091 & ~n92093;
  assign n92974 = ~n92039 & n92071;
  assign n92975 = n92973 & ~n92974;
  assign n92976 = n92033 & ~n92975;
  assign n92977 = n92060 & n92084;
  assign n92978 = ~n92065 & ~n92977;
  assign n92979 = ~n92976 & n92978;
  assign n92980 = ~n92115 & ~n92614;
  assign n92981 = ~n92033 & ~n92980;
  assign n92982 = n92979 & ~n92981;
  assign n92983 = ~n92027 & ~n92982;
  assign n92984 = ~n92972 & ~n92983;
  assign n92985 = ~n92039 & n92104;
  assign n92986 = n92039 & ~n92611;
  assign n92987 = ~n92985 & ~n92986;
  assign n92988 = ~n92033 & ~n92987;
  assign n92989 = ~n92072 & ~n92105;
  assign n92990 = ~n92091 & n92989;
  assign n92991 = n92095 & ~n92990;
  assign n92992 = ~n92988 & ~n92991;
  assign n92993 = n92984 & n92992;
  assign n92994 = ~pi3236 & ~n92993;
  assign n92995 = ~n92972 & n92992;
  assign n92996 = ~n92983 & n92995;
  assign n92997 = pi3236 & n92996;
  assign po3127 = n92994 | n92997;
  assign n92999 = ~n92661 & n92701;
  assign n93000 = ~n92681 & ~n92999;
  assign n93001 = ~n92697 & ~n93000;
  assign n93002 = n92668 & n92689;
  assign n93003 = ~n92668 & n92674;
  assign n93004 = ~n92661 & n93003;
  assign n93005 = ~n93002 & ~n93004;
  assign n93006 = n92697 & ~n93005;
  assign n93007 = ~n92668 & n92710;
  assign n93008 = ~n92835 & ~n93007;
  assign n93009 = ~n92676 & n93008;
  assign n93010 = ~n93006 & n93009;
  assign n93011 = ~n93001 & n93010;
  assign n93012 = ~n92817 & ~n92829;
  assign n93013 = n93011 & n93012;
  assign n93014 = n92649 & ~n93013;
  assign n93015 = n92662 & n92818;
  assign n93016 = n92684 & ~n93015;
  assign n93017 = n92697 & ~n93016;
  assign n93018 = ~n92668 & n92690;
  assign n93019 = ~n93017 & ~n93018;
  assign n93020 = n92655 & n92701;
  assign n93021 = n92668 & n92680;
  assign n93022 = ~n93020 & ~n93021;
  assign n93023 = n92697 & ~n93022;
  assign n93024 = n92689 & n92697;
  assign n93025 = ~n92668 & n93024;
  assign n93026 = ~n93023 & ~n93025;
  assign n93027 = n93019 & n93026;
  assign n93028 = ~n92649 & ~n93027;
  assign n93029 = ~n92710 & ~n92716;
  assign n93030 = ~n92823 & n93029;
  assign n93031 = n92724 & ~n93030;
  assign n93032 = ~n93028 & ~n93031;
  assign n93033 = ~n92676 & ~n92817;
  assign n93034 = ~n92697 & ~n93033;
  assign n93035 = n93032 & ~n93034;
  assign n93036 = ~n93014 & n93035;
  assign n93037 = ~pi3262 & n93036;
  assign n93038 = pi3262 & ~n93036;
  assign po3129 = n93037 | n93038;
  assign n93040 = ~n92033 & n92070;
  assign n93041 = ~n92108 & ~n93040;
  assign n93042 = ~n92113 & n93041;
  assign n93043 = ~n92033 & ~n92989;
  assign n93044 = n92039 & n92061;
  assign n93045 = ~n93043 & ~n93044;
  assign n93046 = n92039 & ~n92051;
  assign n93047 = ~n92068 & ~n93046;
  assign n93048 = ~n92115 & n93047;
  assign n93049 = n92033 & ~n93048;
  assign n93050 = n93045 & ~n93049;
  assign n93051 = ~n92027 & ~n93050;
  assign n93052 = n92033 & n92087;
  assign n93053 = ~n92098 & ~n93052;
  assign n93054 = n92039 & n92072;
  assign n93055 = ~n92033 & n92068;
  assign n93056 = ~n93054 & ~n93055;
  assign n93057 = ~n92631 & n93056;
  assign n93058 = ~n92112 & n93057;
  assign n93059 = n93053 & n93058;
  assign n93060 = ~n92966 & n93059;
  assign n93061 = n92027 & ~n93060;
  assign n93062 = ~n93051 & ~n93061;
  assign n93063 = n93042 & n93062;
  assign n93064 = ~pi3231 & ~n93063;
  assign n93065 = pi3231 & n93042;
  assign n93066 = ~n93051 & n93065;
  assign n93067 = ~n93061 & n93066;
  assign po3130 = n93064 | n93067;
  assign n93069 = n92457 & n92496;
  assign n93070 = n92475 & n92511;
  assign n93071 = ~n92487 & n93070;
  assign n93072 = ~n93069 & ~n93071;
  assign n93073 = n92484 & ~n93072;
  assign n93074 = ~n92518 & ~n92525;
  assign n93075 = ~n92469 & n92516;
  assign n93076 = ~n92520 & ~n93075;
  assign n93077 = ~n92484 & ~n93076;
  assign n93078 = ~n92457 & ~n92484;
  assign n93079 = n92495 & n93078;
  assign n93080 = ~n92463 & n93079;
  assign n93081 = ~n92463 & n92484;
  assign n93082 = ~n92475 & n93081;
  assign n93083 = ~n92469 & n93082;
  assign n93084 = ~n92457 & n92463;
  assign n93085 = ~n92475 & n93084;
  assign n93086 = ~n92487 & n93085;
  assign n93087 = ~n93083 & ~n93086;
  assign n93088 = ~n93080 & n93087;
  assign n93089 = ~n93077 & n93088;
  assign n93090 = n93074 & n93089;
  assign n93091 = n92451 & ~n93090;
  assign n93092 = ~n92484 & n92518;
  assign n93093 = n92457 & n92525;
  assign n93094 = ~n93092 & ~n93093;
  assign n93095 = ~n93091 & n93094;
  assign n93096 = ~n93073 & n93095;
  assign n93097 = n92463 & ~n92469;
  assign n93098 = n92522 & n93097;
  assign n93099 = ~n92497 & ~n93098;
  assign n93100 = n92484 & n92532;
  assign n93101 = n92457 & n92542;
  assign n93102 = ~n93100 & ~n93101;
  assign n93103 = ~n92457 & n92505;
  assign n93104 = ~n93069 & ~n93103;
  assign n93105 = ~n92457 & n92502;
  assign n93106 = ~n92463 & ~n92475;
  assign n93107 = ~n93105 & ~n93106;
  assign n93108 = ~n92484 & ~n93107;
  assign n93109 = n93104 & ~n93108;
  assign n93110 = n93102 & n93109;
  assign n93111 = n93099 & n93110;
  assign n93112 = ~n92451 & ~n93111;
  assign n93113 = n93096 & ~n93112;
  assign n93114 = ~pi3173 & ~n93113;
  assign n93115 = pi3173 & n93096;
  assign n93116 = ~n93112 & n93115;
  assign po3131 = n93114 | n93116;
  assign n93118 = ~n91953 & ~n91959;
  assign n93119 = ~n91926 & ~n93118;
  assign n93120 = ~n92015 & ~n93119;
  assign n93121 = n91932 & n91938;
  assign n93122 = n91926 & n93121;
  assign n93123 = n91952 & n93122;
  assign n93124 = n91952 & n91966;
  assign n93125 = ~n93121 & ~n93124;
  assign n93126 = ~n91932 & ~n91952;
  assign n93127 = ~n91938 & n93126;
  assign n93128 = n93125 & ~n93127;
  assign n93129 = n91926 & ~n93128;
  assign n93130 = ~n91962 & ~n93129;
  assign n93131 = ~n91991 & ~n93130;
  assign n93132 = ~n91926 & n91945;
  assign n93133 = n91952 & n93132;
  assign n93134 = ~n91926 & n91958;
  assign n93135 = ~n93133 & ~n93134;
  assign n93136 = ~n91991 & ~n93135;
  assign n93137 = ~n93131 & ~n93136;
  assign n93138 = ~n93123 & n93137;
  assign n93139 = ~n91938 & n91997;
  assign n93140 = ~n91978 & ~n91998;
  assign n93141 = ~n91932 & n91960;
  assign n93142 = n93140 & ~n93141;
  assign n93143 = ~n91926 & ~n93142;
  assign n93144 = ~n91952 & n91958;
  assign n93145 = ~n91932 & n91945;
  assign n93146 = ~n93144 & ~n93145;
  assign n93147 = n91926 & ~n93146;
  assign n93148 = ~n93143 & ~n93147;
  assign n93149 = ~n93139 & n93148;
  assign n93150 = ~n91968 & ~n92009;
  assign n93151 = n93149 & n93150;
  assign n93152 = n91991 & ~n93151;
  assign n93153 = n93138 & ~n93152;
  assign n93154 = n93120 & n93153;
  assign n93155 = ~pi3323 & ~n93154;
  assign n93156 = pi3323 & n93138;
  assign n93157 = n93120 & n93156;
  assign n93158 = ~n93152 & n93157;
  assign po3132 = n93155 | n93158;
  assign n93160 = pi6971 & pi9040;
  assign n93161 = pi6917 & ~pi9040;
  assign n93162 = ~n93160 & ~n93161;
  assign n93163 = ~pi2960 & n93162;
  assign n93164 = pi2960 & ~n93162;
  assign n93165 = ~n93163 & ~n93164;
  assign n93166 = pi6905 & pi9040;
  assign n93167 = pi6867 & ~pi9040;
  assign n93168 = ~n93166 & ~n93167;
  assign n93169 = pi2973 & n93168;
  assign n93170 = ~pi2973 & ~n93168;
  assign n93171 = ~n93169 & ~n93170;
  assign n93172 = pi6867 & pi9040;
  assign n93173 = pi6970 & ~pi9040;
  assign n93174 = ~n93172 & ~n93173;
  assign n93175 = ~pi2952 & n93174;
  assign n93176 = pi2952 & ~n93174;
  assign n93177 = ~n93175 & ~n93176;
  assign n93178 = ~n93171 & ~n93177;
  assign n93179 = n93165 & n93178;
  assign n93180 = n93171 & ~n93177;
  assign n93181 = ~n93165 & n93180;
  assign n93182 = ~n93179 & ~n93181;
  assign n93183 = pi6998 & pi9040;
  assign n93184 = pi7022 & ~pi9040;
  assign n93185 = ~n93183 & ~n93184;
  assign n93186 = pi2965 & n93185;
  assign n93187 = ~pi2965 & ~n93185;
  assign n93188 = ~n93186 & ~n93187;
  assign n93189 = ~n93165 & ~n93188;
  assign n93190 = n93171 & n93189;
  assign n93191 = n93182 & ~n93190;
  assign n93192 = pi6997 & pi9040;
  assign n93193 = pi6971 & ~pi9040;
  assign n93194 = ~n93192 & ~n93193;
  assign n93195 = ~pi2937 & n93194;
  assign n93196 = pi2937 & ~n93194;
  assign n93197 = ~n93195 & ~n93196;
  assign n93198 = ~pi6963 & pi9040;
  assign n93199 = pi6918 & ~pi9040;
  assign n93200 = ~n93198 & ~n93199;
  assign n93201 = ~pi2944 & n93200;
  assign n93202 = pi2944 & ~n93200;
  assign n93203 = ~n93201 & ~n93202;
  assign n93204 = n93197 & n93203;
  assign n93205 = ~n93191 & n93204;
  assign n93206 = ~n93171 & n93177;
  assign n93207 = ~n93165 & n93206;
  assign n93208 = n93188 & n93203;
  assign n93209 = n93207 & n93208;
  assign n93210 = ~n93165 & n93178;
  assign n93211 = ~n93197 & n93210;
  assign n93212 = n93171 & n93177;
  assign n93213 = n93188 & n93212;
  assign n93214 = n93165 & n93171;
  assign n93215 = ~n93213 & ~n93214;
  assign n93216 = ~n93197 & ~n93215;
  assign n93217 = ~n93211 & ~n93216;
  assign n93218 = n93203 & ~n93217;
  assign n93219 = ~n93209 & ~n93218;
  assign n93220 = n93165 & ~n93188;
  assign n93221 = ~n93171 & n93220;
  assign n93222 = n93177 & n93221;
  assign n93223 = n93165 & n93188;
  assign n93224 = n93171 & n93223;
  assign n93225 = ~n93222 & ~n93224;
  assign n93226 = ~n93197 & ~n93225;
  assign n93227 = n93219 & ~n93226;
  assign n93228 = n93188 & n93197;
  assign n93229 = n93212 & n93228;
  assign n93230 = ~n93165 & n93229;
  assign n93231 = ~n93180 & ~n93206;
  assign n93232 = n93189 & ~n93231;
  assign n93233 = n93179 & ~n93188;
  assign n93234 = ~n93232 & ~n93233;
  assign n93235 = n93165 & n93212;
  assign n93236 = ~n93188 & n93197;
  assign n93237 = n93235 & n93236;
  assign n93238 = n93223 & ~n93231;
  assign n93239 = n93188 & n93210;
  assign n93240 = ~n93238 & ~n93239;
  assign n93241 = ~n93237 & n93240;
  assign n93242 = n93234 & n93241;
  assign n93243 = ~n93230 & n93242;
  assign n93244 = ~n93188 & ~n93197;
  assign n93245 = ~n93165 & n93244;
  assign n93246 = n93177 & n93245;
  assign n93247 = n93243 & ~n93246;
  assign n93248 = ~n93203 & ~n93247;
  assign n93249 = n93227 & ~n93248;
  assign n93250 = ~n93205 & n93249;
  assign n93251 = ~pi3264 & ~n93250;
  assign n93252 = pi3264 & n93227;
  assign n93253 = ~n93205 & n93252;
  assign n93254 = ~n93248 & n93253;
  assign po3133 = n93251 | n93254;
  assign n93256 = ~n93165 & n93212;
  assign n93257 = ~n93197 & n93256;
  assign n93258 = ~n93188 & n93257;
  assign n93259 = n93178 & n93244;
  assign n93260 = n93165 & n93259;
  assign n93261 = ~n93258 & ~n93260;
  assign n93262 = ~n93233 & ~n93237;
  assign n93263 = ~n93165 & ~n93177;
  assign n93264 = n93188 & n93263;
  assign n93265 = ~n93213 & ~n93264;
  assign n93266 = ~n93197 & ~n93265;
  assign n93267 = n93197 & ~n93220;
  assign n93268 = ~n93231 & n93267;
  assign n93269 = ~n93212 & n93244;
  assign n93270 = n93165 & n93269;
  assign n93271 = ~n93268 & ~n93270;
  assign n93272 = ~n93266 & n93271;
  assign n93273 = n93262 & n93272;
  assign n93274 = n93203 & ~n93273;
  assign n93275 = n93261 & ~n93274;
  assign n93276 = n93181 & n93197;
  assign n93277 = n93188 & n93276;
  assign n93278 = n93197 & ~n93203;
  assign n93279 = ~n93210 & ~n93213;
  assign n93280 = n93220 & ~n93231;
  assign n93281 = n93279 & ~n93280;
  assign n93282 = n93278 & ~n93281;
  assign n93283 = n93179 & n93188;
  assign n93284 = ~n93177 & n93188;
  assign n93285 = n93165 & n93284;
  assign n93286 = n93188 & n93206;
  assign n93287 = ~n93285 & ~n93286;
  assign n93288 = ~n93188 & n93212;
  assign n93289 = ~n93207 & ~n93288;
  assign n93290 = n93287 & n93289;
  assign n93291 = ~n93197 & ~n93290;
  assign n93292 = ~n93283 & ~n93291;
  assign n93293 = ~n93203 & ~n93292;
  assign n93294 = ~n93282 & ~n93293;
  assign n93295 = ~n93277 & n93294;
  assign n93296 = n93275 & n93295;
  assign n93297 = pi3331 & ~n93296;
  assign n93298 = ~pi3331 & n93275;
  assign n93299 = n93295 & n93298;
  assign po3134 = n93297 | n93299;
  assign n93301 = ~n91952 & n93145;
  assign n93302 = n91932 & n91981;
  assign n93303 = ~n91978 & ~n93302;
  assign n93304 = n91926 & ~n93303;
  assign n93305 = ~n93301 & ~n93304;
  assign n93306 = ~n91926 & ~n91952;
  assign n93307 = ~n91944 & n93306;
  assign n93308 = ~n91938 & n93307;
  assign n93309 = n91960 & n91994;
  assign n93310 = ~n93308 & ~n93309;
  assign n93311 = ~n93134 & n93310;
  assign n93312 = ~n91956 & ~n91968;
  assign n93313 = ~n92008 & n93312;
  assign n93314 = n93311 & n93313;
  assign n93315 = n93305 & n93314;
  assign n93316 = ~n91991 & ~n93315;
  assign n93317 = n91926 & n91998;
  assign n93318 = ~n91955 & ~n91978;
  assign n93319 = n91952 & ~n93318;
  assign n93320 = ~n91952 & n91966;
  assign n93321 = n91946 & n91952;
  assign n93322 = ~n93320 & ~n93321;
  assign n93323 = ~n91926 & ~n93322;
  assign n93324 = ~n93139 & ~n93141;
  assign n93325 = ~n91932 & ~n91944;
  assign n93326 = n91952 & n93325;
  assign n93327 = n93324 & ~n93326;
  assign n93328 = n91926 & ~n93327;
  assign n93329 = ~n91952 & n91961;
  assign n93330 = ~n93328 & ~n93329;
  assign n93331 = ~n93323 & n93330;
  assign n93332 = ~n93319 & n93331;
  assign n93333 = ~n93317 & n93332;
  assign n93334 = ~n91991 & ~n93317;
  assign n93335 = ~n93333 & ~n93334;
  assign n93336 = ~n91926 & n93301;
  assign n93337 = ~n93335 & ~n93336;
  assign n93338 = ~n93316 & n93337;
  assign n93339 = ~pi3271 & ~n93338;
  assign n93340 = pi3271 & ~n93335;
  assign n93341 = ~n93316 & n93340;
  assign n93342 = ~n93336 & n93341;
  assign po3135 = n93339 | n93342;
  assign n93344 = ~n93093 & ~n93098;
  assign n93345 = ~n92457 & n92490;
  assign n93346 = ~n93086 & ~n93345;
  assign n93347 = ~n93069 & n93346;
  assign n93348 = ~n92484 & ~n93347;
  assign n93349 = n92457 & n92498;
  assign n93350 = n92469 & n92511;
  assign n93351 = ~n92529 & ~n93350;
  assign n93352 = n92484 & ~n93351;
  assign n93353 = ~n93349 & ~n93352;
  assign n93354 = ~n92484 & n92488;
  assign n93355 = n92457 & n93354;
  assign n93356 = ~n92484 & n92496;
  assign n93357 = ~n93355 & ~n93356;
  assign n93358 = n93353 & n93357;
  assign n93359 = n92469 & n92516;
  assign n93360 = ~n93069 & ~n93359;
  assign n93361 = ~n93103 & n93360;
  assign n93362 = n93358 & n93361;
  assign n93363 = ~n92451 & ~n93362;
  assign n93364 = n92484 & n92505;
  assign n93365 = ~n92544 & n93346;
  assign n93366 = ~n92518 & ~n92529;
  assign n93367 = ~n93105 & n93366;
  assign n93368 = ~n92484 & ~n93367;
  assign n93369 = n93365 & ~n93368;
  assign n93370 = ~n93364 & n93369;
  assign n93371 = n92451 & ~n93370;
  assign n93372 = ~n93363 & ~n93371;
  assign n93373 = ~n93348 & n93372;
  assign n93374 = n93344 & n93373;
  assign n93375 = pi3247 & ~n93374;
  assign n93376 = ~pi3247 & n93374;
  assign po3136 = n93375 | n93376;
  assign n93378 = ~n92504 & ~n92512;
  assign n93379 = n92451 & ~n93378;
  assign n93380 = ~n92517 & ~n93075;
  assign n93381 = ~n92477 & n93380;
  assign n93382 = ~n92484 & ~n93381;
  assign n93383 = n92451 & n93382;
  assign n93384 = ~n93379 & ~n93383;
  assign n93385 = n92503 & n93078;
  assign n93386 = ~n93080 & ~n93385;
  assign n93387 = ~n92520 & ~n93106;
  assign n93388 = n92484 & ~n93387;
  assign n93389 = n92451 & n93388;
  assign n93390 = n93386 & ~n93389;
  assign n93391 = n92457 & n92503;
  assign n93392 = n92457 & n92495;
  assign n93393 = ~n93071 & ~n93392;
  assign n93394 = n92484 & ~n93393;
  assign n93395 = ~n92518 & ~n93086;
  assign n93396 = n92457 & n92502;
  assign n93397 = ~n92542 & ~n93396;
  assign n93398 = ~n92484 & ~n93397;
  assign n93399 = n93395 & ~n93398;
  assign n93400 = ~n93394 & n93399;
  assign n93401 = ~n93391 & n93400;
  assign n93402 = ~n92451 & ~n93401;
  assign n93403 = ~n93103 & n93346;
  assign n93404 = n92484 & ~n93403;
  assign n93405 = ~n93402 & ~n93404;
  assign n93406 = n93390 & n93405;
  assign n93407 = n93384 & n93406;
  assign n93408 = ~pi3248 & ~n93407;
  assign n93409 = pi3248 & n93390;
  assign n93410 = n93384 & n93409;
  assign n93411 = n93405 & n93410;
  assign po3137 = n93408 | n93411;
  assign n93413 = n93165 & n93286;
  assign n93414 = ~n93239 & ~n93413;
  assign n93415 = ~n93197 & ~n93414;
  assign n93416 = n93165 & n93180;
  assign n93417 = ~n93256 & ~n93416;
  assign n93418 = ~n93197 & ~n93417;
  assign n93419 = ~n93188 & n93206;
  assign n93420 = ~n93181 & ~n93419;
  assign n93421 = ~n93235 & n93420;
  assign n93422 = n93197 & ~n93421;
  assign n93423 = ~n93418 & ~n93422;
  assign n93424 = ~n93211 & ~n93222;
  assign n93425 = n93423 & n93424;
  assign n93426 = ~n93203 & ~n93425;
  assign n93427 = n93188 & n93256;
  assign n93428 = n93178 & ~n93188;
  assign n93429 = ~n93286 & ~n93428;
  assign n93430 = n93197 & ~n93429;
  assign n93431 = ~n93427 & ~n93430;
  assign n93432 = ~n93197 & n93207;
  assign n93433 = n93182 & ~n93432;
  assign n93434 = ~n93235 & n93433;
  assign n93435 = ~n93188 & ~n93434;
  assign n93436 = n93431 & ~n93435;
  assign n93437 = n93203 & ~n93436;
  assign n93438 = ~n93426 & ~n93437;
  assign n93439 = n93165 & ~n93177;
  assign n93440 = n93197 & n93439;
  assign n93441 = n93188 & n93440;
  assign n93442 = n93438 & ~n93441;
  assign n93443 = ~n93415 & n93442;
  assign n93444 = ~pi3350 & ~n93443;
  assign n93445 = pi3350 & ~n93415;
  assign n93446 = n93438 & n93445;
  assign n93447 = ~n93441 & n93446;
  assign po3138 = n93444 | n93447;
  assign n93449 = ~n92009 & ~n93329;
  assign n93450 = n91926 & ~n93449;
  assign n93451 = ~n91991 & n91993;
  assign n93452 = ~n91926 & n93451;
  assign n93453 = n91938 & n93126;
  assign n93454 = ~n93325 & ~n93453;
  assign n93455 = ~n91961 & n93454;
  assign n93456 = n91926 & ~n93455;
  assign n93457 = ~n91952 & n91967;
  assign n93458 = ~n93456 & ~n93457;
  assign n93459 = ~n91991 & ~n93458;
  assign n93460 = ~n93452 & ~n93459;
  assign n93461 = ~n91956 & ~n91959;
  assign n93462 = ~n91952 & n93141;
  assign n93463 = ~n93302 & ~n93462;
  assign n93464 = n93461 & n93463;
  assign n93465 = ~n91926 & ~n93464;
  assign n93466 = n91932 & ~n91938;
  assign n93467 = ~n91926 & n93466;
  assign n93468 = n91952 & n93467;
  assign n93469 = ~n91952 & n93325;
  assign n93470 = ~n91959 & ~n93469;
  assign n93471 = ~n93321 & n93470;
  assign n93472 = ~n93468 & n93471;
  assign n93473 = n91926 & n91955;
  assign n93474 = n93472 & ~n93473;
  assign n93475 = n91991 & ~n93474;
  assign n93476 = ~n93465 & ~n93475;
  assign n93477 = n93460 & n93476;
  assign n93478 = ~n93450 & n93477;
  assign n93479 = pi3349 & n93478;
  assign n93480 = ~pi3349 & ~n93478;
  assign po3139 = n93479 | n93480;
  assign n93482 = ~n93286 & ~n93288;
  assign n93483 = ~n93197 & ~n93482;
  assign n93484 = ~n93260 & ~n93483;
  assign n93485 = n93203 & ~n93484;
  assign n93486 = ~n93180 & ~n93439;
  assign n93487 = ~n93188 & ~n93486;
  assign n93488 = ~n93256 & ~n93487;
  assign n93489 = n93197 & ~n93488;
  assign n93490 = ~n93280 & ~n93489;
  assign n93491 = n93188 & n93235;
  assign n93492 = ~n93171 & n93189;
  assign n93493 = n93188 & ~n93486;
  assign n93494 = ~n93492 & ~n93493;
  assign n93495 = ~n93197 & ~n93494;
  assign n93496 = ~n93491 & ~n93495;
  assign n93497 = n93490 & n93496;
  assign n93498 = ~n93203 & ~n93497;
  assign n93499 = ~n93165 & n93203;
  assign n93500 = ~n93180 & n93499;
  assign n93501 = n93188 & n93500;
  assign n93502 = n93180 & n93223;
  assign n93503 = ~n93197 & n93502;
  assign n93504 = ~n93165 & ~n93171;
  assign n93505 = n93228 & n93504;
  assign n93506 = ~n93503 & ~n93505;
  assign n93507 = ~n93501 & n93506;
  assign n93508 = ~n93207 & ~n93284;
  assign n93509 = n93204 & ~n93508;
  assign n93510 = n93507 & ~n93509;
  assign n93511 = ~n93498 & n93510;
  assign n93512 = ~n93485 & n93511;
  assign n93513 = pi3329 & ~n93512;
  assign n93514 = ~pi3329 & n93512;
  assign po3140 = n93513 | n93514;
  assign n93516 = ~n92668 & n92680;
  assign n93517 = ~n92707 & ~n93516;
  assign n93518 = ~n92697 & ~n93517;
  assign n93519 = n92697 & ~n92841;
  assign n93520 = ~n92851 & ~n93519;
  assign n93521 = ~n93518 & n93520;
  assign n93522 = n92649 & ~n93521;
  assign n93523 = n92690 & ~n92697;
  assign n93524 = ~n93522 & ~n93523;
  assign n93525 = ~n93007 & ~n93021;
  assign n93526 = n92697 & ~n93525;
  assign n93527 = n92697 & n92708;
  assign n93528 = n92661 & n92701;
  assign n93529 = n92655 & n93528;
  assign n93530 = n92675 & ~n92697;
  assign n93531 = ~n93003 & ~n93530;
  assign n93532 = ~n92655 & ~n93531;
  assign n93533 = ~n93004 & ~n93532;
  assign n93534 = ~n92676 & n93533;
  assign n93535 = ~n93529 & n93534;
  assign n93536 = ~n93527 & n93535;
  assign n93537 = ~n92649 & ~n93536;
  assign n93538 = ~n93526 & ~n93537;
  assign n93539 = n93524 & n93538;
  assign n93540 = pi3273 & ~n93539;
  assign n93541 = ~pi3273 & n93539;
  assign po3141 = n93540 | n93541;
  assign n93543 = pi7150 & ~pi9040;
  assign n93544 = pi7141 & pi9040;
  assign n93545 = ~n93543 & ~n93544;
  assign n93546 = pi3269 & n93545;
  assign n93547 = ~pi3269 & ~n93545;
  assign n93548 = ~n93546 & ~n93547;
  assign n93549 = pi7148 & ~pi9040;
  assign n93550 = pi7248 & pi9040;
  assign n93551 = ~n93549 & ~n93550;
  assign n93552 = ~pi3272 & n93551;
  assign n93553 = pi3272 & ~n93551;
  assign n93554 = ~n93552 & ~n93553;
  assign n93555 = pi7143 & ~pi9040;
  assign n93556 = pi7177 & pi9040;
  assign n93557 = ~n93555 & ~n93556;
  assign n93558 = ~pi3325 & n93557;
  assign n93559 = pi3325 & ~n93557;
  assign n93560 = ~n93558 & ~n93559;
  assign n93561 = pi7117 & ~pi9040;
  assign n93562 = pi7135 & pi9040;
  assign n93563 = ~n93561 & ~n93562;
  assign n93564 = ~pi3267 & ~n93563;
  assign n93565 = pi3267 & n93563;
  assign n93566 = ~n93564 & ~n93565;
  assign n93567 = ~n93560 & n93566;
  assign n93568 = n93554 & n93567;
  assign n93569 = pi7156 & ~pi9040;
  assign n93570 = pi7153 & pi9040;
  assign n93571 = ~n93569 & ~n93570;
  assign n93572 = pi3403 & n93571;
  assign n93573 = ~pi3403 & ~n93571;
  assign n93574 = ~n93572 & ~n93573;
  assign n93575 = n93568 & ~n93574;
  assign n93576 = n93560 & ~n93566;
  assign n93577 = n93554 & n93576;
  assign n93578 = ~n93574 & n93577;
  assign n93579 = ~n93575 & ~n93578;
  assign n93580 = ~n93554 & n93576;
  assign n93581 = n93574 & n93580;
  assign n93582 = ~n93560 & ~n93566;
  assign n93583 = n93554 & n93582;
  assign n93584 = n93574 & n93583;
  assign n93585 = ~n93581 & ~n93584;
  assign n93586 = n93579 & n93585;
  assign n93587 = n93548 & ~n93586;
  assign n93588 = n93560 & n93566;
  assign n93589 = n93554 & n93588;
  assign n93590 = n93574 & n93589;
  assign n93591 = ~n93583 & ~n93590;
  assign n93592 = n93548 & ~n93591;
  assign n93593 = ~n93548 & n93566;
  assign n93594 = ~n93574 & n93593;
  assign n93595 = ~n93554 & ~n93560;
  assign n93596 = n93574 & n93576;
  assign n93597 = ~n93595 & ~n93596;
  assign n93598 = ~n93548 & ~n93597;
  assign n93599 = ~n93594 & ~n93598;
  assign n93600 = ~n93554 & n93588;
  assign n93601 = ~n93574 & n93600;
  assign n93602 = n93599 & ~n93601;
  assign n93603 = n93566 & n93595;
  assign n93604 = n93574 & n93603;
  assign n93605 = n93602 & ~n93604;
  assign n93606 = ~n93592 & n93605;
  assign n93607 = pi7117 & pi9040;
  assign n93608 = pi7294 & ~pi9040;
  assign n93609 = ~n93607 & ~n93608;
  assign n93610 = ~pi3347 & ~n93609;
  assign n93611 = pi3347 & n93609;
  assign n93612 = ~n93610 & ~n93611;
  assign n93613 = ~n93606 & ~n93612;
  assign n93614 = n93554 & n93566;
  assign n93615 = ~n93548 & n93574;
  assign n93616 = n93612 & n93615;
  assign n93617 = n93614 & n93616;
  assign n93618 = n93554 & ~n93574;
  assign n93619 = ~n93566 & n93618;
  assign n93620 = ~n93548 & ~n93619;
  assign n93621 = ~n93554 & n93574;
  assign n93622 = n93560 & n93621;
  assign n93623 = ~n93567 & ~n93614;
  assign n93624 = ~n93574 & ~n93623;
  assign n93625 = n93548 & ~n93580;
  assign n93626 = ~n93624 & n93625;
  assign n93627 = ~n93622 & n93626;
  assign n93628 = ~n93620 & ~n93627;
  assign n93629 = ~n93566 & n93621;
  assign n93630 = ~n93560 & n93629;
  assign n93631 = ~n93628 & ~n93630;
  assign n93632 = n93612 & ~n93631;
  assign n93633 = ~n93617 & ~n93632;
  assign n93634 = ~n93613 & n93633;
  assign n93635 = ~n93587 & n93634;
  assign n93636 = ~n93548 & n93601;
  assign n93637 = n93635 & ~n93636;
  assign n93638 = pi3762 & ~n93637;
  assign n93639 = ~pi3762 & ~n93636;
  assign n93640 = n93634 & n93639;
  assign n93641 = ~n93587 & n93640;
  assign po3160 = n93638 | n93641;
  assign n93643 = pi7285 & ~pi9040;
  assign n93644 = pi7101 & pi9040;
  assign n93645 = ~n93643 & ~n93644;
  assign n93646 = ~pi3348 & ~n93645;
  assign n93647 = pi3348 & n93645;
  assign n93648 = ~n93646 & ~n93647;
  assign n93649 = pi7164 & ~pi9040;
  assign n93650 = pi7156 & pi9040;
  assign n93651 = ~n93649 & ~n93650;
  assign n93652 = ~pi3404 & ~n93651;
  assign n93653 = pi3404 & n93651;
  assign n93654 = ~n93652 & ~n93653;
  assign n93655 = ~n93648 & ~n93654;
  assign n93656 = pi7137 & pi9040;
  assign n93657 = pi7232 & ~pi9040;
  assign n93658 = ~n93656 & ~n93657;
  assign n93659 = pi3268 & n93658;
  assign n93660 = ~pi3268 & ~n93658;
  assign n93661 = ~n93659 & ~n93660;
  assign n93662 = pi7137 & ~pi9040;
  assign n93663 = pi7294 & pi9040;
  assign n93664 = ~n93662 & ~n93663;
  assign n93665 = ~pi3357 & ~n93664;
  assign n93666 = pi3357 & n93664;
  assign n93667 = ~n93665 & ~n93666;
  assign n93668 = pi7161 & ~pi9040;
  assign n93669 = pi7136 & pi9040;
  assign n93670 = ~n93668 & ~n93669;
  assign n93671 = pi3270 & n93670;
  assign n93672 = ~pi3270 & ~n93670;
  assign n93673 = ~n93671 & ~n93672;
  assign n93674 = n93667 & ~n93673;
  assign n93675 = ~n93661 & n93674;
  assign n93676 = pi7146 & pi9040;
  assign n93677 = pi7142 & ~pi9040;
  assign n93678 = ~n93676 & ~n93677;
  assign n93679 = pi3310 & n93678;
  assign n93680 = ~pi3310 & ~n93678;
  assign n93681 = ~n93679 & ~n93680;
  assign n93682 = n93673 & ~n93681;
  assign n93683 = n93667 & n93682;
  assign n93684 = n93661 & n93683;
  assign n93685 = n93673 & n93681;
  assign n93686 = ~n93661 & n93685;
  assign n93687 = ~n93684 & ~n93686;
  assign n93688 = ~n93675 & n93687;
  assign n93689 = n93655 & ~n93688;
  assign n93690 = ~n93661 & ~n93667;
  assign n93691 = ~n93681 & n93690;
  assign n93692 = ~n93673 & ~n93681;
  assign n93693 = n93667 & n93692;
  assign n93694 = n93661 & n93693;
  assign n93695 = ~n93691 & ~n93694;
  assign n93696 = ~n93667 & n93682;
  assign n93697 = n93667 & n93685;
  assign n93698 = ~n93696 & ~n93697;
  assign n93699 = n93695 & n93698;
  assign n93700 = n93648 & ~n93699;
  assign n93701 = ~n93673 & n93681;
  assign n93702 = ~n93667 & n93701;
  assign n93703 = n93661 & n93702;
  assign n93704 = ~n93700 & ~n93703;
  assign n93705 = ~n93654 & ~n93704;
  assign n93706 = ~n93689 & ~n93705;
  assign n93707 = n93648 & ~n93661;
  assign n93708 = n93667 & n93707;
  assign n93709 = n93681 & n93708;
  assign n93710 = ~n93661 & n93696;
  assign n93711 = ~n93709 & ~n93710;
  assign n93712 = ~n93685 & ~n93692;
  assign n93713 = n93661 & ~n93712;
  assign n93714 = ~n93667 & n93692;
  assign n93715 = ~n93713 & ~n93714;
  assign n93716 = ~n93648 & ~n93715;
  assign n93717 = n93667 & n93701;
  assign n93718 = ~n93675 & ~n93717;
  assign n93719 = ~n93684 & n93718;
  assign n93720 = n93648 & ~n93719;
  assign n93721 = ~n93716 & ~n93720;
  assign n93722 = ~n93648 & ~n93661;
  assign n93723 = n93682 & n93722;
  assign n93724 = n93661 & ~n93667;
  assign n93725 = ~n93681 & n93724;
  assign n93726 = ~n93673 & n93725;
  assign n93727 = ~n93667 & n93673;
  assign n93728 = n93681 & n93727;
  assign n93729 = n93661 & n93728;
  assign n93730 = ~n93726 & ~n93729;
  assign n93731 = ~n93661 & n93702;
  assign n93732 = n93730 & ~n93731;
  assign n93733 = ~n93723 & n93732;
  assign n93734 = n93721 & n93733;
  assign n93735 = n93654 & ~n93734;
  assign n93736 = n93711 & ~n93735;
  assign n93737 = n93706 & n93736;
  assign n93738 = pi3763 & ~n93737;
  assign n93739 = ~pi3763 & n93711;
  assign n93740 = n93706 & n93739;
  assign n93741 = ~n93735 & n93740;
  assign po3166 = n93738 | n93741;
  assign n93743 = n93661 & n93674;
  assign n93744 = ~n93697 & ~n93743;
  assign n93745 = ~n93710 & n93744;
  assign n93746 = n93648 & ~n93745;
  assign n93747 = ~n93661 & n93728;
  assign n93748 = ~n93661 & n93717;
  assign n93749 = ~n93667 & ~n93673;
  assign n93750 = ~n93682 & ~n93749;
  assign n93751 = n93661 & ~n93750;
  assign n93752 = ~n93748 & ~n93751;
  assign n93753 = ~n93747 & n93752;
  assign n93754 = ~n93648 & ~n93753;
  assign n93755 = ~n93746 & ~n93754;
  assign n93756 = n93654 & ~n93755;
  assign n93757 = ~n93648 & n93714;
  assign n93758 = ~n93661 & n93757;
  assign n93759 = ~n93661 & n93683;
  assign n93760 = ~n93648 & n93759;
  assign n93761 = ~n93758 & ~n93760;
  assign n93762 = n93648 & n93731;
  assign n93763 = n93761 & ~n93762;
  assign n93764 = ~n93673 & n93707;
  assign n93765 = ~n93661 & n93673;
  assign n93766 = n93667 & n93765;
  assign n93767 = ~n93743 & ~n93766;
  assign n93768 = ~n93648 & ~n93767;
  assign n93769 = ~n93723 & ~n93768;
  assign n93770 = ~n93729 & ~n93759;
  assign n93771 = n93648 & ~n93667;
  assign n93772 = n93701 & n93771;
  assign n93773 = n93648 & n93661;
  assign n93774 = n93727 & n93773;
  assign n93775 = ~n93772 & ~n93774;
  assign n93776 = n93770 & n93775;
  assign n93777 = n93769 & n93776;
  assign n93778 = ~n93764 & n93777;
  assign n93779 = ~n93654 & ~n93778;
  assign n93780 = ~n93661 & n93667;
  assign n93781 = ~n93681 & n93780;
  assign n93782 = ~n93673 & n93781;
  assign n93783 = n93661 & n93685;
  assign n93784 = ~n93782 & ~n93783;
  assign n93785 = n93648 & ~n93784;
  assign n93786 = ~n93779 & ~n93785;
  assign n93787 = n93763 & n93786;
  assign n93788 = ~n93756 & n93787;
  assign n93789 = ~pi3783 & ~n93788;
  assign n93790 = pi3783 & n93788;
  assign po3167 = n93789 | n93790;
  assign n93792 = pi7232 & pi9040;
  assign n93793 = pi7101 & ~pi9040;
  assign n93794 = ~n93792 & ~n93793;
  assign n93795 = ~pi3267 & ~n93794;
  assign n93796 = pi3267 & n93794;
  assign n93797 = ~n93795 & ~n93796;
  assign n93798 = pi7159 & ~pi9040;
  assign n93799 = pi7164 & pi9040;
  assign n93800 = ~n93798 & ~n93799;
  assign n93801 = ~pi3404 & n93800;
  assign n93802 = pi3404 & ~n93800;
  assign n93803 = ~n93801 & ~n93802;
  assign n93804 = pi7148 & pi9040;
  assign n93805 = pi7141 & ~pi9040;
  assign n93806 = ~n93804 & ~n93805;
  assign n93807 = pi3272 & n93806;
  assign n93808 = ~pi3272 & ~n93806;
  assign n93809 = ~n93807 & ~n93808;
  assign n93810 = n93803 & n93809;
  assign n93811 = pi7153 & ~pi9040;
  assign n93812 = pi7250 & pi9040;
  assign n93813 = ~n93811 & ~n93812;
  assign n93814 = ~pi3309 & ~n93813;
  assign n93815 = pi3309 & n93813;
  assign n93816 = ~n93814 & ~n93815;
  assign n93817 = pi7285 & pi9040;
  assign n93818 = pi7250 & ~pi9040;
  assign n93819 = ~n93817 & ~n93818;
  assign n93820 = pi3358 & n93819;
  assign n93821 = ~pi3358 & ~n93819;
  assign n93822 = ~n93820 & ~n93821;
  assign n93823 = ~n93816 & ~n93822;
  assign n93824 = n93810 & n93823;
  assign n93825 = pi7158 & pi9040;
  assign n93826 = pi7177 & ~pi9040;
  assign n93827 = ~n93825 & ~n93826;
  assign n93828 = ~pi3310 & n93827;
  assign n93829 = pi3310 & ~n93827;
  assign n93830 = ~n93828 & ~n93829;
  assign n93831 = ~n93803 & ~n93809;
  assign n93832 = ~n93830 & n93831;
  assign n93833 = n93816 & n93830;
  assign n93834 = ~n93809 & n93833;
  assign n93835 = n93803 & n93834;
  assign n93836 = ~n93832 & ~n93835;
  assign n93837 = ~n93803 & n93809;
  assign n93838 = n93816 & n93837;
  assign n93839 = n93836 & ~n93838;
  assign n93840 = ~n93822 & ~n93839;
  assign n93841 = ~n93803 & n93830;
  assign n93842 = ~n93816 & n93822;
  assign n93843 = n93841 & n93842;
  assign n93844 = n93830 & n93831;
  assign n93845 = ~n93816 & n93844;
  assign n93846 = ~n93843 & ~n93845;
  assign n93847 = ~n93840 & n93846;
  assign n93848 = ~n93824 & n93847;
  assign n93849 = ~n93830 & n93837;
  assign n93850 = n93816 & n93849;
  assign n93851 = n93810 & ~n93830;
  assign n93852 = ~n93816 & n93851;
  assign n93853 = ~n93850 & ~n93852;
  assign n93854 = n93848 & n93853;
  assign n93855 = ~n93797 & ~n93854;
  assign n93856 = ~n93816 & n93830;
  assign n93857 = n93809 & n93856;
  assign n93858 = ~n93803 & n93857;
  assign n93859 = ~n93851 & ~n93858;
  assign n93860 = ~n93822 & ~n93859;
  assign n93861 = ~n93803 & n93833;
  assign n93862 = ~n93816 & n93849;
  assign n93863 = ~n93861 & ~n93862;
  assign n93864 = n93822 & ~n93863;
  assign n93865 = n93810 & n93833;
  assign n93866 = ~n93809 & n93856;
  assign n93867 = n93803 & n93866;
  assign n93868 = ~n93865 & ~n93867;
  assign n93869 = ~n93864 & n93868;
  assign n93870 = ~n93860 & n93869;
  assign n93871 = n93797 & ~n93870;
  assign n93872 = ~n93803 & ~n93830;
  assign n93873 = n93816 & n93872;
  assign n93874 = n93803 & ~n93830;
  assign n93875 = ~n93816 & n93874;
  assign n93876 = ~n93873 & ~n93875;
  assign n93877 = ~n93822 & ~n93876;
  assign n93878 = n93803 & ~n93809;
  assign n93879 = ~n93830 & n93878;
  assign n93880 = n93816 & n93879;
  assign n93881 = ~n93865 & ~n93880;
  assign n93882 = ~n93844 & n93881;
  assign n93883 = n93822 & ~n93882;
  assign n93884 = ~n93877 & ~n93883;
  assign n93885 = ~n93809 & n93830;
  assign n93886 = n93822 & n93885;
  assign n93887 = ~n93816 & n93886;
  assign n93888 = n93884 & ~n93887;
  assign n93889 = ~n93871 & n93888;
  assign n93890 = ~n93855 & n93889;
  assign n93891 = ~pi3710 & ~n93890;
  assign n93892 = pi3710 & n93890;
  assign po3168 = n93891 | n93892;
  assign n93894 = ~n93714 & ~n93717;
  assign n93895 = ~n93648 & ~n93894;
  assign n93896 = n93661 & n93697;
  assign n93897 = ~n93895 & ~n93896;
  assign n93898 = n93661 & n93673;
  assign n93899 = ~n93727 & ~n93898;
  assign n93900 = ~n93693 & n93899;
  assign n93901 = n93648 & ~n93900;
  assign n93902 = n93897 & ~n93901;
  assign n93903 = ~n93654 & ~n93902;
  assign n93904 = ~n93648 & n93747;
  assign n93905 = ~n93760 & ~n93904;
  assign n93906 = ~n93762 & n93905;
  assign n93907 = ~n93731 & ~n93781;
  assign n93908 = n93648 & n93766;
  assign n93909 = n93661 & n93717;
  assign n93910 = ~n93648 & n93727;
  assign n93911 = ~n93909 & ~n93910;
  assign n93912 = ~n93726 & n93911;
  assign n93913 = ~n93908 & n93912;
  assign n93914 = n93907 & n93913;
  assign n93915 = ~n93772 & n93914;
  assign n93916 = n93654 & ~n93915;
  assign n93917 = n93906 & ~n93916;
  assign n93918 = ~n93903 & n93917;
  assign n93919 = ~pi3781 & ~n93918;
  assign n93920 = pi3781 & n93906;
  assign n93921 = ~n93903 & n93920;
  assign n93922 = ~n93916 & n93921;
  assign po3171 = n93919 | n93922;
  assign n93924 = n93816 & n93844;
  assign n93925 = ~n93867 & ~n93872;
  assign n93926 = n93822 & ~n93925;
  assign n93927 = ~n93924 & ~n93926;
  assign n93928 = ~n93858 & n93927;
  assign n93929 = ~n93822 & n93865;
  assign n93930 = ~n93852 & ~n93929;
  assign n93931 = ~n93880 & n93930;
  assign n93932 = n93928 & n93931;
  assign n93933 = n93797 & ~n93932;
  assign n93934 = ~n93816 & n93879;
  assign n93935 = n93809 & ~n93830;
  assign n93936 = ~n93803 & n93816;
  assign n93937 = ~n93935 & ~n93936;
  assign n93938 = ~n93885 & n93937;
  assign n93939 = ~n93822 & ~n93938;
  assign n93940 = ~n93934 & ~n93939;
  assign n93941 = n93816 & n93851;
  assign n93942 = n93830 & n93837;
  assign n93943 = n93816 & n93942;
  assign n93944 = ~n93835 & ~n93943;
  assign n93945 = n93810 & n93830;
  assign n93946 = n93822 & n93945;
  assign n93947 = n93944 & ~n93946;
  assign n93948 = ~n93941 & n93947;
  assign n93949 = ~n93845 & n93948;
  assign n93950 = n93940 & n93949;
  assign n93951 = ~n93797 & ~n93950;
  assign n93952 = ~n93933 & ~n93951;
  assign n93953 = pi3761 & ~n93952;
  assign n93954 = ~pi3761 & ~n93933;
  assign n93955 = ~n93951 & n93954;
  assign po3174 = n93953 | n93955;
  assign n93957 = pi7155 & ~pi9040;
  assign n93958 = pi7293 & pi9040;
  assign n93959 = ~n93957 & ~n93958;
  assign n93960 = ~pi3324 & ~n93959;
  assign n93961 = pi3324 & n93959;
  assign n93962 = ~n93960 & ~n93961;
  assign n93963 = pi7224 & ~pi9040;
  assign n93964 = pi7218 & pi9040;
  assign n93965 = ~n93963 & ~n93964;
  assign n93966 = ~pi3325 & ~n93965;
  assign n93967 = pi3325 & n93965;
  assign n93968 = ~n93966 & ~n93967;
  assign n93969 = pi7169 & pi9040;
  assign n93970 = pi7292 & ~pi9040;
  assign n93971 = ~n93969 & ~n93970;
  assign n93972 = ~pi3347 & ~n93971;
  assign n93973 = pi3347 & n93971;
  assign n93974 = ~n93972 & ~n93973;
  assign n93975 = pi7272 & pi9040;
  assign n93976 = pi7147 & ~pi9040;
  assign n93977 = ~n93975 & ~n93976;
  assign n93978 = ~pi3266 & ~n93977;
  assign n93979 = pi3266 & n93977;
  assign n93980 = ~n93978 & ~n93979;
  assign n93981 = ~n93974 & n93980;
  assign n93982 = pi7233 & ~pi9040;
  assign n93983 = pi7157 & pi9040;
  assign n93984 = ~n93982 & ~n93983;
  assign n93985 = ~pi3332 & n93984;
  assign n93986 = pi3332 & ~n93984;
  assign n93987 = ~n93985 & ~n93986;
  assign n93988 = pi7118 & pi9040;
  assign n93989 = pi7235 & ~pi9040;
  assign n93990 = ~n93988 & ~n93989;
  assign n93991 = pi3405 & n93990;
  assign n93992 = ~pi3405 & ~n93990;
  assign n93993 = ~n93991 & ~n93992;
  assign n93994 = ~n93987 & n93993;
  assign n93995 = n93981 & n93994;
  assign n93996 = n93968 & n93995;
  assign n93997 = n93987 & n93993;
  assign n93998 = n93974 & n93980;
  assign n93999 = n93997 & n93998;
  assign n94000 = n93968 & n93987;
  assign n94001 = ~n93980 & n94000;
  assign n94002 = ~n93974 & n94001;
  assign n94003 = n93974 & ~n93980;
  assign n94004 = n93968 & n94003;
  assign n94005 = n93993 & n94004;
  assign n94006 = ~n93987 & n94005;
  assign n94007 = ~n94002 & ~n94006;
  assign n94008 = ~n93999 & n94007;
  assign n94009 = ~n93996 & n94008;
  assign n94010 = ~n93968 & n93987;
  assign n94011 = n93998 & n94010;
  assign n94012 = n94009 & ~n94011;
  assign n94013 = ~n93962 & ~n94012;
  assign n94014 = n93968 & n93974;
  assign n94015 = n93980 & n94014;
  assign n94016 = ~n93987 & n94015;
  assign n94017 = ~n94001 & ~n94016;
  assign n94018 = ~n93968 & n93981;
  assign n94019 = ~n93987 & n94018;
  assign n94020 = n94017 & ~n94019;
  assign n94021 = ~n93993 & ~n94020;
  assign n94022 = ~n93968 & ~n93980;
  assign n94023 = n93974 & n94022;
  assign n94024 = ~n93993 & n94023;
  assign n94025 = ~n93987 & n94024;
  assign n94026 = ~n93974 & n94000;
  assign n94027 = ~n93974 & ~n93980;
  assign n94028 = n93987 & n94027;
  assign n94029 = ~n94026 & ~n94028;
  assign n94030 = ~n93993 & ~n94029;
  assign n94031 = ~n94025 & ~n94030;
  assign n94032 = ~n93962 & ~n94031;
  assign n94033 = ~n94021 & ~n94032;
  assign n94034 = ~n94013 & n94033;
  assign n94035 = ~n93968 & ~n93987;
  assign n94036 = n93993 & n94035;
  assign n94037 = n94027 & n94036;
  assign n94038 = ~n93968 & n93974;
  assign n94039 = n93997 & n94038;
  assign n94040 = n93987 & n94023;
  assign n94041 = n93968 & ~n93993;
  assign n94042 = n93974 & n94041;
  assign n94043 = ~n93974 & ~n93987;
  assign n94044 = ~n93968 & n94043;
  assign n94045 = ~n94042 & ~n94044;
  assign n94046 = ~n94040 & n94045;
  assign n94047 = ~n94018 & n94046;
  assign n94048 = n93981 & n93993;
  assign n94049 = n93987 & n94048;
  assign n94050 = ~n93987 & n94027;
  assign n94051 = ~n93968 & n93980;
  assign n94052 = ~n94050 & ~n94051;
  assign n94053 = n93993 & ~n94052;
  assign n94054 = ~n94049 & ~n94053;
  assign n94055 = n94047 & n94054;
  assign n94056 = n93962 & ~n94055;
  assign n94057 = ~n94039 & ~n94056;
  assign n94058 = ~n94037 & n94057;
  assign n94059 = n94034 & n94058;
  assign n94060 = pi3759 & n94059;
  assign n94061 = ~pi3759 & ~n94059;
  assign po3175 = n94060 | n94061;
  assign n94063 = n93648 & n93685;
  assign n94064 = ~n93661 & n94063;
  assign n94065 = ~n93782 & ~n94064;
  assign n94066 = n93661 & n93681;
  assign n94067 = n93667 & n94066;
  assign n94068 = ~n93661 & ~n93673;
  assign n94069 = ~n93781 & ~n94068;
  assign n94070 = ~n93648 & ~n94069;
  assign n94071 = ~n94067 & ~n94070;
  assign n94072 = n94065 & n94071;
  assign n94073 = n93654 & ~n94072;
  assign n94074 = ~n93683 & ~n93729;
  assign n94075 = ~n93661 & n93701;
  assign n94076 = n94074 & ~n94075;
  assign n94077 = n93648 & ~n94076;
  assign n94078 = n93685 & n93722;
  assign n94079 = ~n93710 & ~n94078;
  assign n94080 = ~n94077 & n94079;
  assign n94081 = ~n93693 & ~n93703;
  assign n94082 = ~n93648 & ~n94081;
  assign n94083 = n94080 & ~n94082;
  assign n94084 = ~n93654 & ~n94083;
  assign n94085 = ~n94073 & ~n94084;
  assign n94086 = ~n93661 & n93692;
  assign n94087 = n93661 & ~n93698;
  assign n94088 = ~n94086 & ~n94087;
  assign n94089 = ~n93648 & ~n94088;
  assign n94090 = ~n93683 & n93894;
  assign n94091 = n93773 & ~n94090;
  assign n94092 = ~n94089 & ~n94091;
  assign n94093 = n94085 & n94092;
  assign n94094 = ~pi3778 & ~n94093;
  assign n94095 = pi3778 & n94092;
  assign n94096 = ~n94084 & n94095;
  assign n94097 = ~n94073 & n94096;
  assign po3176 = n94094 | n94097;
  assign n94099 = n93968 & ~n93974;
  assign n94100 = ~n94011 & ~n94099;
  assign n94101 = ~n94043 & n94100;
  assign n94102 = n93993 & ~n94101;
  assign n94103 = ~n93987 & ~n93993;
  assign n94104 = n93974 & n94103;
  assign n94105 = n93968 & ~n93987;
  assign n94106 = n93980 & n94105;
  assign n94107 = n93987 & n94004;
  assign n94108 = ~n94106 & ~n94107;
  assign n94109 = ~n93968 & ~n93974;
  assign n94110 = n93987 & ~n93993;
  assign n94111 = n94109 & n94110;
  assign n94112 = n94108 & ~n94111;
  assign n94113 = ~n94104 & n94112;
  assign n94114 = ~n94102 & n94113;
  assign n94115 = n93962 & ~n94114;
  assign n94116 = n93968 & n93981;
  assign n94117 = n93987 & n94116;
  assign n94118 = ~n93980 & n94099;
  assign n94119 = ~n93987 & n94118;
  assign n94120 = ~n94117 & ~n94119;
  assign n94121 = n93993 & ~n94120;
  assign n94122 = ~n94115 & ~n94121;
  assign n94123 = ~n93987 & n94004;
  assign n94124 = ~n94015 & ~n94023;
  assign n94125 = n93993 & ~n94124;
  assign n94126 = ~n94123 & ~n94125;
  assign n94127 = ~n94019 & n94126;
  assign n94128 = ~n93962 & ~n94127;
  assign n94129 = ~n93998 & ~n94027;
  assign n94130 = ~n93968 & ~n94129;
  assign n94131 = ~n94028 & ~n94130;
  assign n94132 = ~n93993 & ~n94131;
  assign n94133 = ~n93962 & n94132;
  assign n94134 = ~n94128 & ~n94133;
  assign n94135 = n94122 & n94134;
  assign n94136 = pi3776 & ~n94135;
  assign n94137 = ~pi3776 & n94122;
  assign n94138 = n94134 & n94137;
  assign po3177 = n94136 | n94138;
  assign n94140 = ~n93575 & ~n93581;
  assign n94141 = ~n93548 & ~n94140;
  assign n94142 = ~n93636 & ~n94141;
  assign n94143 = n93554 & n93560;
  assign n94144 = n93548 & n94143;
  assign n94145 = n93574 & n94144;
  assign n94146 = n93574 & n93588;
  assign n94147 = ~n94143 & ~n94146;
  assign n94148 = ~n93554 & ~n93574;
  assign n94149 = ~n93560 & n94148;
  assign n94150 = n94147 & ~n94149;
  assign n94151 = n93548 & ~n94150;
  assign n94152 = ~n93584 & ~n94151;
  assign n94153 = ~n93612 & ~n94152;
  assign n94154 = ~n93548 & n93567;
  assign n94155 = n93574 & n94154;
  assign n94156 = ~n93548 & n93580;
  assign n94157 = ~n94155 & ~n94156;
  assign n94158 = ~n93612 & ~n94157;
  assign n94159 = ~n94153 & ~n94158;
  assign n94160 = ~n94145 & n94159;
  assign n94161 = ~n93560 & n93618;
  assign n94162 = ~n93600 & ~n93619;
  assign n94163 = ~n93554 & n93582;
  assign n94164 = n94162 & ~n94163;
  assign n94165 = ~n93548 & ~n94164;
  assign n94166 = n93576 & n94148;
  assign n94167 = ~n93603 & ~n94166;
  assign n94168 = n93548 & ~n94167;
  assign n94169 = ~n94165 & ~n94168;
  assign n94170 = ~n94161 & n94169;
  assign n94171 = ~n93590 & ~n93630;
  assign n94172 = n94170 & n94171;
  assign n94173 = n93612 & ~n94172;
  assign n94174 = n94160 & ~n94173;
  assign n94175 = n94142 & n94174;
  assign n94176 = ~pi3849 & ~n94175;
  assign n94177 = pi3849 & n94160;
  assign n94178 = n94142 & n94177;
  assign n94179 = ~n94173 & n94178;
  assign po3179 = n94176 | n94179;
  assign n94181 = pi7136 & ~pi9040;
  assign n94182 = pi7150 & pi9040;
  assign n94183 = ~n94181 & ~n94182;
  assign n94184 = ~pi3270 & ~n94183;
  assign n94185 = pi3270 & n94183;
  assign n94186 = ~n94184 & ~n94185;
  assign n94187 = pi7142 & pi9040;
  assign n94188 = pi7248 & ~pi9040;
  assign n94189 = ~n94187 & ~n94188;
  assign n94190 = pi3360 & n94189;
  assign n94191 = ~pi3360 & ~n94189;
  assign n94192 = ~n94190 & ~n94191;
  assign n94193 = pi7146 & ~pi9040;
  assign n94194 = pi7144 & pi9040;
  assign n94195 = ~n94193 & ~n94194;
  assign n94196 = ~pi3314 & n94195;
  assign n94197 = pi3314 & ~n94195;
  assign n94198 = ~n94196 & ~n94197;
  assign n94199 = ~n94192 & n94198;
  assign n94200 = pi7161 & pi9040;
  assign n94201 = pi7154 & ~pi9040;
  assign n94202 = ~n94200 & ~n94201;
  assign n94203 = ~pi3422 & n94202;
  assign n94204 = pi3422 & ~n94202;
  assign n94205 = ~n94203 & ~n94204;
  assign n94206 = n94199 & ~n94205;
  assign n94207 = pi7246 & ~pi9040;
  assign n94208 = pi7154 & pi9040;
  assign n94209 = ~n94207 & ~n94208;
  assign n94210 = pi3326 & n94209;
  assign n94211 = ~pi3326 & ~n94209;
  assign n94212 = ~n94210 & ~n94211;
  assign n94213 = pi7159 & pi9040;
  assign n94214 = pi7165 & ~pi9040;
  assign n94215 = ~n94213 & ~n94214;
  assign n94216 = pi3357 & n94215;
  assign n94217 = ~pi3357 & ~n94215;
  assign n94218 = ~n94216 & ~n94217;
  assign n94219 = n94205 & ~n94218;
  assign n94220 = n94212 & n94219;
  assign n94221 = n94192 & n94220;
  assign n94222 = n94205 & n94218;
  assign n94223 = ~n94212 & n94222;
  assign n94224 = n94192 & n94223;
  assign n94225 = ~n94221 & ~n94224;
  assign n94226 = ~n94205 & n94218;
  assign n94227 = ~n94212 & n94226;
  assign n94228 = ~n94212 & n94219;
  assign n94229 = ~n94192 & n94228;
  assign n94230 = ~n94227 & ~n94229;
  assign n94231 = ~n94198 & ~n94230;
  assign n94232 = n94225 & ~n94231;
  assign n94233 = ~n94206 & n94232;
  assign n94234 = n94186 & ~n94233;
  assign n94235 = ~n94205 & ~n94218;
  assign n94236 = ~n94212 & n94235;
  assign n94237 = n94192 & n94236;
  assign n94238 = n94198 & n94237;
  assign n94239 = ~n94192 & ~n94198;
  assign n94240 = n94236 & n94239;
  assign n94241 = ~n94192 & n94212;
  assign n94242 = n94205 & n94241;
  assign n94243 = ~n94240 & ~n94242;
  assign n94244 = n94212 & n94222;
  assign n94245 = ~n94227 & ~n94244;
  assign n94246 = ~n94192 & n94222;
  assign n94247 = n94245 & ~n94246;
  assign n94248 = n94198 & ~n94247;
  assign n94249 = n94212 & ~n94218;
  assign n94250 = ~n94205 & n94249;
  assign n94251 = n94192 & n94250;
  assign n94252 = n94192 & ~n94212;
  assign n94253 = ~n94218 & n94252;
  assign n94254 = n94205 & n94253;
  assign n94255 = ~n94251 & ~n94254;
  assign n94256 = n94212 & n94226;
  assign n94257 = ~n94198 & n94256;
  assign n94258 = n94255 & ~n94257;
  assign n94259 = ~n94248 & n94258;
  assign n94260 = n94243 & n94259;
  assign n94261 = ~n94186 & ~n94260;
  assign n94262 = ~n94238 & ~n94261;
  assign n94263 = ~n94234 & n94262;
  assign n94264 = n94239 & n94244;
  assign n94265 = ~n94198 & n94249;
  assign n94266 = n94192 & n94265;
  assign n94267 = ~n94264 & ~n94266;
  assign n94268 = ~n94198 & n94224;
  assign n94269 = n94267 & ~n94268;
  assign n94270 = n94263 & n94269;
  assign n94271 = ~pi3800 & ~n94270;
  assign n94272 = pi3800 & n94269;
  assign n94273 = n94262 & n94272;
  assign n94274 = ~n94234 & n94273;
  assign po3182 = n94271 | n94274;
  assign n94276 = n94205 & ~n94212;
  assign n94277 = ~n94212 & ~n94218;
  assign n94278 = ~n94192 & n94277;
  assign n94279 = n94192 & n94219;
  assign n94280 = ~n94278 & ~n94279;
  assign n94281 = ~n94276 & n94280;
  assign n94282 = ~n94256 & n94281;
  assign n94283 = ~n94198 & ~n94282;
  assign n94284 = n94218 & n94241;
  assign n94285 = ~n94227 & ~n94242;
  assign n94286 = n94198 & ~n94285;
  assign n94287 = ~n94284 & ~n94286;
  assign n94288 = ~n94283 & n94287;
  assign n94289 = ~n94251 & n94288;
  assign n94290 = n94186 & ~n94289;
  assign n94291 = ~n94192 & ~n94212;
  assign n94292 = n94222 & n94291;
  assign n94293 = n94255 & ~n94292;
  assign n94294 = ~n94198 & ~n94293;
  assign n94295 = ~n94290 & ~n94294;
  assign n94296 = ~n94205 & n94284;
  assign n94297 = n94198 & n94252;
  assign n94298 = ~n94205 & n94297;
  assign n94299 = n94192 & n94244;
  assign n94300 = ~n94192 & n94265;
  assign n94301 = ~n94299 & ~n94300;
  assign n94302 = n94205 & n94212;
  assign n94303 = n94192 & n94302;
  assign n94304 = ~n94236 & ~n94303;
  assign n94305 = n94198 & ~n94304;
  assign n94306 = n94198 & n94276;
  assign n94307 = ~n94192 & n94306;
  assign n94308 = ~n94305 & ~n94307;
  assign n94309 = n94301 & n94308;
  assign n94310 = ~n94186 & ~n94309;
  assign n94311 = ~n94298 & ~n94310;
  assign n94312 = ~n94296 & n94311;
  assign n94313 = n94295 & n94312;
  assign n94314 = ~pi3843 & ~n94313;
  assign n94315 = ~n94290 & ~n94296;
  assign n94316 = ~n94294 & n94315;
  assign n94317 = n94311 & n94316;
  assign n94318 = pi3843 & n94317;
  assign po3183 = n94314 | n94318;
  assign n94320 = ~n93574 & n93603;
  assign n94321 = n93574 & n93614;
  assign n94322 = ~n93600 & ~n94321;
  assign n94323 = n93548 & ~n94322;
  assign n94324 = ~n94320 & ~n94323;
  assign n94325 = ~n93548 & ~n93574;
  assign n94326 = n93566 & n94325;
  assign n94327 = ~n93560 & n94326;
  assign n94328 = ~n93566 & n93615;
  assign n94329 = ~n93560 & n94328;
  assign n94330 = ~n94327 & ~n94329;
  assign n94331 = ~n94156 & n94330;
  assign n94332 = ~n93578 & ~n93590;
  assign n94333 = ~n93629 & n94332;
  assign n94334 = n94331 & n94333;
  assign n94335 = n94324 & n94334;
  assign n94336 = ~n93612 & ~n94335;
  assign n94337 = ~n93577 & ~n93600;
  assign n94338 = n93574 & ~n94337;
  assign n94339 = ~n93574 & n93588;
  assign n94340 = n93554 & n93574;
  assign n94341 = n93566 & n94340;
  assign n94342 = ~n93560 & n94341;
  assign n94343 = ~n94339 & ~n94342;
  assign n94344 = ~n93548 & ~n94343;
  assign n94345 = ~n94161 & ~n94163;
  assign n94346 = ~n93554 & n93566;
  assign n94347 = n93574 & n94346;
  assign n94348 = n94345 & ~n94347;
  assign n94349 = n93548 & ~n94348;
  assign n94350 = ~n93574 & n93583;
  assign n94351 = ~n94349 & ~n94350;
  assign n94352 = ~n94344 & n94351;
  assign n94353 = ~n94338 & n94352;
  assign n94354 = n93612 & ~n94353;
  assign n94355 = n93548 & n93619;
  assign n94356 = ~n94354 & ~n94355;
  assign n94357 = ~n93548 & n94320;
  assign n94358 = n94356 & ~n94357;
  assign n94359 = ~n94336 & n94358;
  assign n94360 = ~pi3809 & ~n94359;
  assign n94361 = pi3809 & n94356;
  assign n94362 = ~n94336 & n94361;
  assign n94363 = ~n94357 & n94362;
  assign po3184 = n94360 | n94363;
  assign n94365 = pi7118 & ~pi9040;
  assign n94366 = pi7138 & pi9040;
  assign n94367 = ~n94365 & ~n94366;
  assign n94368 = ~pi3422 & ~n94367;
  assign n94369 = pi3422 & n94367;
  assign n94370 = ~n94368 & ~n94369;
  assign n94371 = pi7423 & pi9040;
  assign n94372 = pi7234 & ~pi9040;
  assign n94373 = ~n94371 & ~n94372;
  assign n94374 = ~pi3353 & n94373;
  assign n94375 = pi3353 & ~n94373;
  assign n94376 = ~n94374 & ~n94375;
  assign n94377 = pi7230 & ~pi9040;
  assign n94378 = pi7235 & pi9040;
  assign n94379 = ~n94377 & ~n94378;
  assign n94380 = pi3351 & n94379;
  assign n94381 = ~pi3351 & ~n94379;
  assign n94382 = ~n94380 & ~n94381;
  assign n94383 = pi7423 & ~pi9040;
  assign n94384 = pi7147 & pi9040;
  assign n94385 = ~n94383 & ~n94384;
  assign n94386 = pi3311 & n94385;
  assign n94387 = ~pi3311 & ~n94385;
  assign n94388 = ~n94386 & ~n94387;
  assign n94389 = pi7138 & ~pi9040;
  assign n94390 = pi7229 & pi9040;
  assign n94391 = ~n94389 & ~n94390;
  assign n94392 = ~pi3326 & n94391;
  assign n94393 = pi3326 & ~n94391;
  assign n94394 = ~n94392 & ~n94393;
  assign n94395 = ~n94388 & ~n94394;
  assign n94396 = n94382 & n94395;
  assign n94397 = ~n94376 & n94396;
  assign n94398 = pi7145 & pi9040;
  assign n94399 = pi7426 & ~pi9040;
  assign n94400 = ~n94398 & ~n94399;
  assign n94401 = ~pi3387 & ~n94400;
  assign n94402 = pi3387 & n94400;
  assign n94403 = ~n94401 & ~n94402;
  assign n94404 = ~pi3311 & n94385;
  assign n94405 = pi3311 & ~n94385;
  assign n94406 = ~n94404 & ~n94405;
  assign n94407 = ~n94394 & ~n94406;
  assign n94408 = ~n94376 & n94407;
  assign n94409 = ~n94382 & n94395;
  assign n94410 = n94376 & n94409;
  assign n94411 = ~n94408 & ~n94410;
  assign n94412 = ~n94403 & ~n94411;
  assign n94413 = ~n94397 & ~n94412;
  assign n94414 = ~n94388 & n94394;
  assign n94415 = ~n94382 & n94414;
  assign n94416 = n94403 & n94415;
  assign n94417 = n94395 & n94403;
  assign n94418 = ~n94376 & n94417;
  assign n94419 = ~n94416 & ~n94418;
  assign n94420 = n94413 & n94419;
  assign n94421 = n94394 & ~n94406;
  assign n94422 = n94382 & n94421;
  assign n94423 = ~n94376 & n94422;
  assign n94424 = n94382 & n94414;
  assign n94425 = n94376 & n94424;
  assign n94426 = ~n94423 & ~n94425;
  assign n94427 = n94420 & n94426;
  assign n94428 = n94370 & ~n94427;
  assign n94429 = ~n94370 & ~n94403;
  assign n94430 = ~n94376 & ~n94382;
  assign n94431 = n94406 & n94430;
  assign n94432 = ~n94382 & n94394;
  assign n94433 = ~n94431 & ~n94432;
  assign n94434 = n94429 & ~n94433;
  assign n94435 = n94382 & ~n94388;
  assign n94436 = ~n94394 & n94435;
  assign n94437 = n94376 & n94436;
  assign n94438 = n94376 & ~n94406;
  assign n94439 = ~n94382 & n94438;
  assign n94440 = ~n94437 & ~n94439;
  assign n94441 = ~n94376 & n94403;
  assign n94442 = ~n94395 & n94441;
  assign n94443 = n94382 & n94442;
  assign n94444 = n94403 & n94422;
  assign n94445 = ~n94443 & ~n94444;
  assign n94446 = n94440 & n94445;
  assign n94447 = ~n94370 & ~n94446;
  assign n94448 = ~n94382 & n94421;
  assign n94449 = ~n94403 & n94448;
  assign n94450 = n94376 & n94449;
  assign n94451 = n94382 & n94407;
  assign n94452 = n94376 & n94451;
  assign n94453 = ~n94425 & ~n94452;
  assign n94454 = ~n94403 & ~n94453;
  assign n94455 = ~n94450 & ~n94454;
  assign n94456 = n94403 & n94437;
  assign n94457 = n94455 & ~n94456;
  assign n94458 = ~n94447 & n94457;
  assign n94459 = ~n94434 & n94458;
  assign n94460 = ~n94428 & n94459;
  assign n94461 = ~n94382 & n94407;
  assign n94462 = n94376 & n94403;
  assign n94463 = n94461 & n94462;
  assign n94464 = n94460 & ~n94463;
  assign n94465 = ~pi3764 & ~n94464;
  assign n94466 = ~n94428 & ~n94463;
  assign n94467 = n94459 & n94466;
  assign n94468 = pi3764 & n94467;
  assign po3186 = n94465 | n94468;
  assign n94470 = n93987 & n94018;
  assign n94471 = ~n94107 & ~n94470;
  assign n94472 = ~n93993 & ~n94471;
  assign n94473 = n94015 & n94103;
  assign n94474 = ~n94472 & ~n94473;
  assign n94475 = ~n94039 & n94474;
  assign n94476 = ~n93987 & n94023;
  assign n94477 = ~n94018 & ~n94476;
  assign n94478 = ~n94118 & n94477;
  assign n94479 = ~n93993 & ~n94478;
  assign n94480 = n93962 & n94479;
  assign n94481 = n93968 & n93993;
  assign n94482 = ~n93980 & n94481;
  assign n94483 = ~n93974 & n94482;
  assign n94484 = n93987 & n94483;
  assign n94485 = n93993 & n94116;
  assign n94486 = ~n94011 & ~n94037;
  assign n94487 = ~n94006 & n94486;
  assign n94488 = ~n94485 & n94487;
  assign n94489 = n93962 & ~n94488;
  assign n94490 = ~n93987 & n94048;
  assign n94491 = ~n94483 & ~n94490;
  assign n94492 = ~n94106 & n94491;
  assign n94493 = ~n93980 & n94010;
  assign n94494 = ~n93987 & n93998;
  assign n94495 = ~n94014 & ~n94494;
  assign n94496 = ~n93993 & ~n94495;
  assign n94497 = ~n94493 & ~n94496;
  assign n94498 = n94492 & n94497;
  assign n94499 = ~n93962 & ~n94498;
  assign n94500 = ~n94489 & ~n94499;
  assign n94501 = ~n94484 & n94500;
  assign n94502 = ~n94480 & n94501;
  assign n94503 = n94475 & n94502;
  assign n94504 = pi3824 & ~n94503;
  assign n94505 = ~pi3824 & n94475;
  assign n94506 = n94502 & n94505;
  assign po3187 = n94504 | n94506;
  assign n94508 = ~n93810 & ~n93831;
  assign n94509 = n93822 & ~n94508;
  assign n94510 = ~n93816 & n94509;
  assign n94511 = ~n93849 & ~n93878;
  assign n94512 = n93816 & ~n94511;
  assign n94513 = n93822 & n94512;
  assign n94514 = n93830 & n94509;
  assign n94515 = ~n94513 & ~n94514;
  assign n94516 = ~n94510 & n94515;
  assign n94517 = ~n93797 & ~n94516;
  assign n94518 = ~n93816 & n93837;
  assign n94519 = ~n93934 & ~n94518;
  assign n94520 = n93822 & n94519;
  assign n94521 = ~n93830 & ~n94508;
  assign n94522 = n93803 & n93856;
  assign n94523 = n93816 & n93831;
  assign n94524 = ~n94522 & ~n94523;
  assign n94525 = n93816 & n93874;
  assign n94526 = n94524 & ~n94525;
  assign n94527 = ~n94521 & n94526;
  assign n94528 = ~n93822 & n94527;
  assign n94529 = ~n94520 & ~n94528;
  assign n94530 = n93816 & n94521;
  assign n94531 = ~n93943 & ~n94530;
  assign n94532 = ~n94529 & n94531;
  assign n94533 = n93797 & ~n94532;
  assign n94534 = ~n94517 & ~n94533;
  assign n94535 = n93822 & n93835;
  assign n94536 = ~n93822 & ~n94531;
  assign n94537 = ~n94535 & ~n94536;
  assign n94538 = ~n93822 & ~n94519;
  assign n94539 = ~n93835 & ~n94538;
  assign n94540 = ~n93797 & ~n94539;
  assign n94541 = n94537 & ~n94540;
  assign n94542 = n94534 & n94541;
  assign n94543 = pi3771 & ~n94542;
  assign n94544 = ~pi3771 & n94541;
  assign n94545 = ~n94517 & n94544;
  assign n94546 = ~n94533 & n94545;
  assign po3189 = n94543 | n94546;
  assign n94548 = ~n93987 & n94130;
  assign n94549 = ~n94022 & ~n94116;
  assign n94550 = ~n93993 & ~n94549;
  assign n94551 = ~n94548 & ~n94550;
  assign n94552 = ~n93980 & n94105;
  assign n94553 = ~n94051 & ~n94552;
  assign n94554 = ~n94118 & n94553;
  assign n94555 = n93993 & ~n94554;
  assign n94556 = n94551 & ~n94555;
  assign n94557 = n93987 & n94015;
  assign n94558 = n94556 & ~n94557;
  assign n94559 = ~n93962 & ~n94558;
  assign n94560 = n93997 & ~n94549;
  assign n94561 = ~n94018 & ~n94023;
  assign n94562 = ~n94015 & ~n94118;
  assign n94563 = n94561 & n94562;
  assign n94564 = ~n93987 & ~n94563;
  assign n94565 = ~n94560 & ~n94564;
  assign n94566 = ~n94107 & n94565;
  assign n94567 = n93962 & ~n94566;
  assign n94568 = ~n94559 & ~n94567;
  assign n94569 = ~n93987 & n94116;
  assign n94570 = ~n94557 & ~n94569;
  assign n94571 = ~n93993 & ~n94570;
  assign n94572 = n94568 & ~n94571;
  assign n94573 = pi3810 & ~n94572;
  assign n94574 = ~pi3810 & ~n94571;
  assign n94575 = ~n94567 & n94574;
  assign n94576 = ~n94559 & n94575;
  assign po3190 = n94573 | n94576;
  assign n94578 = pi7140 & pi9040;
  assign n94579 = pi7218 & ~pi9040;
  assign n94580 = ~n94578 & ~n94579;
  assign n94581 = pi3327 & n94580;
  assign n94582 = ~pi3327 & ~n94580;
  assign n94583 = ~n94581 & ~n94582;
  assign n94584 = pi7169 & ~pi9040;
  assign n94585 = pi7426 & pi9040;
  assign n94586 = ~n94584 & ~n94585;
  assign n94587 = pi3324 & n94586;
  assign n94588 = ~pi3324 & ~n94586;
  assign n94589 = ~n94587 & ~n94588;
  assign n94590 = pi7151 & ~pi9040;
  assign n94591 = pi7234 & pi9040;
  assign n94592 = ~n94590 & ~n94591;
  assign n94593 = pi3356 & n94592;
  assign n94594 = ~pi3356 & ~n94592;
  assign n94595 = ~n94593 & ~n94594;
  assign n94596 = n94589 & ~n94595;
  assign n94597 = pi7166 & ~pi9040;
  assign n94598 = pi7228 & pi9040;
  assign n94599 = ~n94597 & ~n94598;
  assign n94600 = ~pi3359 & ~n94599;
  assign n94601 = pi3359 & n94599;
  assign n94602 = ~n94600 & ~n94601;
  assign n94603 = pi7224 & pi9040;
  assign n94604 = pi7157 & ~pi9040;
  assign n94605 = ~n94603 & ~n94604;
  assign n94606 = ~pi3266 & ~n94605;
  assign n94607 = pi3266 & n94605;
  assign n94608 = ~n94606 & ~n94607;
  assign n94609 = n94602 & n94608;
  assign n94610 = n94596 & n94609;
  assign n94611 = n94602 & ~n94608;
  assign n94612 = ~n94589 & n94611;
  assign n94613 = ~n94610 & ~n94612;
  assign n94614 = ~n94583 & ~n94613;
  assign n94615 = pi7151 & pi9040;
  assign n94616 = pi7160 & ~pi9040;
  assign n94617 = ~n94615 & ~n94616;
  assign n94618 = ~pi3346 & ~n94617;
  assign n94619 = pi3346 & n94617;
  assign n94620 = ~n94618 & ~n94619;
  assign n94621 = n94583 & ~n94602;
  assign n94622 = n94589 & n94621;
  assign n94623 = n94596 & ~n94608;
  assign n94624 = n94589 & n94595;
  assign n94625 = n94608 & n94624;
  assign n94626 = ~n94623 & ~n94625;
  assign n94627 = ~n94589 & ~n94595;
  assign n94628 = n94608 & n94627;
  assign n94629 = n94602 & n94628;
  assign n94630 = n94626 & ~n94629;
  assign n94631 = n94583 & ~n94630;
  assign n94632 = ~n94622 & ~n94631;
  assign n94633 = ~n94589 & n94595;
  assign n94634 = ~n94608 & n94633;
  assign n94635 = n94602 & n94634;
  assign n94636 = n94632 & ~n94635;
  assign n94637 = ~n94602 & n94627;
  assign n94638 = n94608 & n94633;
  assign n94639 = ~n94637 & ~n94638;
  assign n94640 = ~n94583 & ~n94639;
  assign n94641 = ~n94608 & n94624;
  assign n94642 = ~n94602 & n94641;
  assign n94643 = ~n94640 & ~n94642;
  assign n94644 = n94636 & n94643;
  assign n94645 = n94620 & ~n94644;
  assign n94646 = ~n94614 & ~n94645;
  assign n94647 = n94583 & ~n94620;
  assign n94648 = ~n94639 & n94647;
  assign n94649 = ~n94608 & n94627;
  assign n94650 = ~n94641 & ~n94649;
  assign n94651 = n94602 & ~n94650;
  assign n94652 = ~n94610 & ~n94651;
  assign n94653 = ~n94620 & ~n94652;
  assign n94654 = ~n94648 & ~n94653;
  assign n94655 = ~n94583 & ~n94620;
  assign n94656 = n94596 & ~n94602;
  assign n94657 = ~n94634 & ~n94656;
  assign n94658 = n94589 & n94608;
  assign n94659 = n94657 & ~n94658;
  assign n94660 = n94655 & ~n94659;
  assign n94661 = n94654 & ~n94660;
  assign n94662 = n94646 & n94661;
  assign n94663 = ~pi3779 & ~n94662;
  assign n94664 = pi3779 & n94654;
  assign n94665 = n94646 & n94664;
  assign n94666 = ~n94660 & n94665;
  assign po3191 = n94663 | n94666;
  assign n94668 = n94376 & n94415;
  assign n94669 = n94394 & n94430;
  assign n94670 = ~n94406 & n94669;
  assign n94671 = ~n94668 & ~n94670;
  assign n94672 = n94403 & ~n94671;
  assign n94673 = ~n94403 & n94437;
  assign n94674 = ~n94437 & ~n94444;
  assign n94675 = ~n94376 & n94382;
  assign n94676 = ~n94394 & n94675;
  assign n94677 = ~n94406 & n94676;
  assign n94678 = ~n94376 & ~n94403;
  assign n94679 = n94414 & n94678;
  assign n94680 = ~n94382 & n94679;
  assign n94681 = n94376 & n94382;
  assign n94682 = ~n94388 & n94681;
  assign n94683 = ~n94439 & ~n94682;
  assign n94684 = ~n94403 & ~n94683;
  assign n94685 = ~n94382 & n94403;
  assign n94686 = ~n94394 & n94685;
  assign n94687 = ~n94388 & n94686;
  assign n94688 = ~n94684 & ~n94687;
  assign n94689 = ~n94680 & n94688;
  assign n94690 = ~n94677 & n94689;
  assign n94691 = n94674 & n94690;
  assign n94692 = n94370 & ~n94691;
  assign n94693 = n94376 & n94444;
  assign n94694 = ~n94692 & ~n94693;
  assign n94695 = ~n94673 & n94694;
  assign n94696 = ~n94672 & n94695;
  assign n94697 = n94435 & n94441;
  assign n94698 = ~n94416 & ~n94697;
  assign n94699 = n94403 & n94451;
  assign n94700 = n94376 & n94461;
  assign n94701 = ~n94699 & ~n94700;
  assign n94702 = ~n94376 & n94424;
  assign n94703 = ~n94668 & ~n94702;
  assign n94704 = ~n94376 & n94421;
  assign n94705 = ~n94382 & ~n94394;
  assign n94706 = ~n94704 & ~n94705;
  assign n94707 = ~n94403 & ~n94706;
  assign n94708 = n94703 & ~n94707;
  assign n94709 = n94701 & n94708;
  assign n94710 = n94698 & n94709;
  assign n94711 = ~n94370 & ~n94710;
  assign n94712 = n94696 & ~n94711;
  assign n94713 = ~pi3760 & ~n94712;
  assign n94714 = pi3760 & n94696;
  assign n94715 = ~n94711 & n94714;
  assign po3192 = n94713 | n94715;
  assign n94717 = ~n93630 & ~n94350;
  assign n94718 = n93548 & ~n94717;
  assign n94719 = ~n93612 & n93614;
  assign n94720 = ~n93548 & n94719;
  assign n94721 = n93560 & n94148;
  assign n94722 = ~n94346 & ~n94721;
  assign n94723 = ~n93583 & n94722;
  assign n94724 = n93548 & ~n94723;
  assign n94725 = ~n93574 & n93589;
  assign n94726 = ~n94724 & ~n94725;
  assign n94727 = ~n93612 & ~n94726;
  assign n94728 = ~n94720 & ~n94727;
  assign n94729 = ~n93578 & ~n93581;
  assign n94730 = ~n93574 & n94163;
  assign n94731 = ~n94321 & ~n94730;
  assign n94732 = n94729 & n94731;
  assign n94733 = ~n93548 & ~n94732;
  assign n94734 = n93554 & ~n93560;
  assign n94735 = ~n93548 & n94734;
  assign n94736 = n93574 & n94735;
  assign n94737 = ~n93574 & n94346;
  assign n94738 = ~n93581 & ~n94737;
  assign n94739 = ~n94342 & n94738;
  assign n94740 = ~n94736 & n94739;
  assign n94741 = n93548 & n93577;
  assign n94742 = n94740 & ~n94741;
  assign n94743 = n93612 & ~n94742;
  assign n94744 = ~n94733 & ~n94743;
  assign n94745 = n94728 & n94744;
  assign n94746 = ~n94718 & n94745;
  assign n94747 = pi3867 & n94746;
  assign n94748 = ~pi3867 & ~n94746;
  assign po3193 = n94747 | n94748;
  assign n94750 = ~n94192 & n94220;
  assign n94751 = ~n94223 & ~n94296;
  assign n94752 = n94192 & n94249;
  assign n94753 = ~n94192 & n94236;
  assign n94754 = ~n94752 & ~n94753;
  assign n94755 = n94751 & n94754;
  assign n94756 = n94198 & ~n94755;
  assign n94757 = n94192 & n94226;
  assign n94758 = ~n94242 & ~n94757;
  assign n94759 = ~n94228 & n94758;
  assign n94760 = ~n94198 & ~n94759;
  assign n94761 = n94218 & n94252;
  assign n94762 = ~n94205 & n94761;
  assign n94763 = ~n94760 & ~n94762;
  assign n94764 = ~n94756 & n94763;
  assign n94765 = ~n94750 & n94764;
  assign n94766 = ~n94186 & ~n94765;
  assign n94767 = n94192 & n94198;
  assign n94768 = n94256 & n94767;
  assign n94769 = n94198 & n94228;
  assign n94770 = n94198 & n94244;
  assign n94771 = ~n94769 & ~n94770;
  assign n94772 = ~n94192 & ~n94771;
  assign n94773 = ~n94768 & ~n94772;
  assign n94774 = ~n94192 & n94250;
  assign n94775 = ~n94237 & ~n94774;
  assign n94776 = ~n94192 & n94226;
  assign n94777 = n94192 & n94222;
  assign n94778 = ~n94776 & ~n94777;
  assign n94779 = ~n94250 & n94778;
  assign n94780 = ~n94223 & n94779;
  assign n94781 = ~n94198 & ~n94780;
  assign n94782 = ~n94192 & n94227;
  assign n94783 = ~n94781 & ~n94782;
  assign n94784 = n94775 & n94783;
  assign n94785 = n94773 & n94784;
  assign n94786 = n94186 & ~n94785;
  assign n94787 = n94198 & ~n94225;
  assign n94788 = ~n94786 & ~n94787;
  assign n94789 = ~n94254 & ~n94774;
  assign n94790 = ~n94198 & ~n94789;
  assign n94791 = n94788 & ~n94790;
  assign n94792 = ~n94766 & n94791;
  assign n94793 = pi3864 & ~n94792;
  assign n94794 = ~pi3864 & n94792;
  assign po3194 = n94793 | n94794;
  assign n94796 = ~n94693 & ~n94697;
  assign n94797 = ~n94437 & ~n94448;
  assign n94798 = ~n94704 & n94797;
  assign n94799 = ~n94403 & ~n94798;
  assign n94800 = ~n94376 & n94409;
  assign n94801 = ~n94677 & ~n94800;
  assign n94802 = ~n94463 & n94801;
  assign n94803 = n94403 & n94424;
  assign n94804 = n94802 & ~n94803;
  assign n94805 = ~n94799 & n94804;
  assign n94806 = n94370 & ~n94805;
  assign n94807 = n94376 & n94417;
  assign n94808 = n94388 & n94430;
  assign n94809 = ~n94448 & ~n94808;
  assign n94810 = n94403 & ~n94809;
  assign n94811 = ~n94807 & ~n94810;
  assign n94812 = ~n94403 & n94407;
  assign n94813 = n94376 & n94812;
  assign n94814 = ~n94403 & n94415;
  assign n94815 = ~n94813 & ~n94814;
  assign n94816 = n94811 & n94815;
  assign n94817 = n94388 & n94681;
  assign n94818 = ~n94668 & ~n94817;
  assign n94819 = ~n94702 & n94818;
  assign n94820 = n94816 & n94819;
  assign n94821 = ~n94370 & ~n94820;
  assign n94822 = ~n94668 & n94801;
  assign n94823 = ~n94403 & ~n94822;
  assign n94824 = ~n94821 & ~n94823;
  assign n94825 = ~n94806 & n94824;
  assign n94826 = n94796 & n94825;
  assign n94827 = pi3767 & ~n94826;
  assign n94828 = ~pi3767 & n94826;
  assign po3195 = n94827 | n94828;
  assign n94830 = pi7155 & pi9040;
  assign n94831 = pi7162 & ~pi9040;
  assign n94832 = ~n94830 & ~n94831;
  assign n94833 = pi3330 & n94832;
  assign n94834 = ~pi3330 & ~n94832;
  assign n94835 = ~n94833 & ~n94834;
  assign n94836 = pi7160 & pi9040;
  assign n94837 = pi7228 & ~pi9040;
  assign n94838 = ~n94836 & ~n94837;
  assign n94839 = pi3265 & n94838;
  assign n94840 = ~pi3265 & ~n94838;
  assign n94841 = ~n94839 & ~n94840;
  assign n94842 = pi7140 & ~pi9040;
  assign n94843 = pi7162 & pi9040;
  assign n94844 = ~n94842 & ~n94843;
  assign n94845 = pi3346 & n94844;
  assign n94846 = ~pi3346 & ~n94844;
  assign n94847 = ~n94845 & ~n94846;
  assign n94848 = pi7236 & pi9040;
  assign n94849 = pi7229 & ~pi9040;
  assign n94850 = ~n94848 & ~n94849;
  assign n94851 = pi3356 & n94850;
  assign n94852 = ~pi3356 & ~n94850;
  assign n94853 = ~n94851 & ~n94852;
  assign n94854 = n94847 & ~n94853;
  assign n94855 = ~n94841 & n94854;
  assign n94856 = n94835 & n94855;
  assign n94857 = pi7085 & ~pi9040;
  assign n94858 = pi7166 & pi9040;
  assign n94859 = ~n94857 & ~n94858;
  assign n94860 = pi3311 & ~n94859;
  assign n94861 = ~pi3311 & n94859;
  assign n94862 = ~n94860 & ~n94861;
  assign n94863 = pi7236 & ~pi9040;
  assign n94864 = pi7231 & pi9040;
  assign n94865 = ~n94863 & ~n94864;
  assign n94866 = ~pi3351 & n94865;
  assign n94867 = pi3351 & ~n94865;
  assign n94868 = ~n94866 & ~n94867;
  assign n94869 = n94847 & ~n94868;
  assign n94870 = n94853 & n94869;
  assign n94871 = ~n94847 & ~n94868;
  assign n94872 = ~n94853 & n94871;
  assign n94873 = ~n94847 & n94868;
  assign n94874 = ~n94835 & n94873;
  assign n94875 = ~n94872 & ~n94874;
  assign n94876 = ~n94870 & n94875;
  assign n94877 = ~n94841 & ~n94876;
  assign n94878 = n94853 & n94871;
  assign n94879 = ~n94853 & n94869;
  assign n94880 = ~n94878 & ~n94879;
  assign n94881 = n94841 & ~n94880;
  assign n94882 = ~n94877 & ~n94881;
  assign n94883 = n94847 & n94868;
  assign n94884 = n94853 & n94883;
  assign n94885 = n94841 & n94884;
  assign n94886 = ~n94853 & n94874;
  assign n94887 = ~n94885 & ~n94886;
  assign n94888 = n94882 & n94887;
  assign n94889 = n94862 & ~n94888;
  assign n94890 = n94835 & n94878;
  assign n94891 = ~n94835 & n94883;
  assign n94892 = n94835 & n94873;
  assign n94893 = ~n94891 & ~n94892;
  assign n94894 = ~n94841 & ~n94893;
  assign n94895 = ~n94890 & ~n94894;
  assign n94896 = n94853 & n94873;
  assign n94897 = n94841 & n94896;
  assign n94898 = ~n94853 & n94883;
  assign n94899 = ~n94870 & ~n94898;
  assign n94900 = ~n94897 & n94899;
  assign n94901 = ~n94872 & n94900;
  assign n94902 = ~n94835 & ~n94901;
  assign n94903 = n94895 & ~n94902;
  assign n94904 = ~n94862 & ~n94903;
  assign n94905 = ~n94889 & ~n94904;
  assign n94906 = ~n94856 & n94905;
  assign n94907 = n94835 & n94853;
  assign n94908 = n94868 & n94907;
  assign n94909 = n94847 & n94908;
  assign n94910 = ~n94853 & n94892;
  assign n94911 = ~n94909 & ~n94910;
  assign n94912 = n94841 & ~n94911;
  assign n94913 = n94906 & ~n94912;
  assign n94914 = ~pi3789 & ~n94913;
  assign n94915 = pi3789 & ~n94912;
  assign n94916 = n94905 & n94915;
  assign n94917 = ~n94856 & n94916;
  assign po3196 = n94914 | n94917;
  assign n94919 = n93816 & n93945;
  assign n94920 = n93822 & n94919;
  assign n94921 = n93856 & ~n94508;
  assign n94922 = ~n93879 & ~n93943;
  assign n94923 = ~n94921 & n94922;
  assign n94924 = ~n93822 & ~n94923;
  assign n94925 = n93816 & n93832;
  assign n94926 = ~n94924 & ~n94925;
  assign n94927 = n93830 & n93878;
  assign n94928 = ~n93816 & n93935;
  assign n94929 = ~n94927 & ~n94928;
  assign n94930 = ~n94523 & n94929;
  assign n94931 = n93822 & ~n94930;
  assign n94932 = n94926 & ~n94931;
  assign n94933 = n93797 & ~n94932;
  assign n94934 = ~n94920 & ~n94933;
  assign n94935 = ~n93816 & n93831;
  assign n94936 = ~n93942 & ~n94935;
  assign n94937 = n93822 & ~n94936;
  assign n94938 = ~n93880 & ~n94937;
  assign n94939 = ~n93850 & ~n94919;
  assign n94940 = ~n93816 & n93832;
  assign n94941 = n93816 & n93885;
  assign n94942 = ~n93935 & ~n94941;
  assign n94943 = ~n94927 & n94942;
  assign n94944 = ~n93822 & ~n94943;
  assign n94945 = ~n94940 & ~n94944;
  assign n94946 = n94939 & n94945;
  assign n94947 = n94938 & n94946;
  assign n94948 = ~n93797 & ~n94947;
  assign n94949 = ~n93862 & ~n94525;
  assign n94950 = ~n93822 & ~n94949;
  assign n94951 = ~n94948 & ~n94950;
  assign n94952 = n94934 & n94951;
  assign n94953 = pi3770 & n94952;
  assign n94954 = ~pi3770 & ~n94952;
  assign po3197 = n94953 | n94954;
  assign n94956 = ~n94583 & n94602;
  assign n94957 = ~n94627 & ~n94641;
  assign n94958 = n94956 & ~n94957;
  assign n94959 = ~n94583 & ~n94608;
  assign n94960 = n94627 & n94959;
  assign n94961 = ~n94958 & ~n94960;
  assign n94962 = n94620 & ~n94961;
  assign n94963 = ~n94602 & n94625;
  assign n94964 = ~n94602 & n94608;
  assign n94965 = ~n94658 & ~n94964;
  assign n94966 = n94583 & ~n94965;
  assign n94967 = ~n94602 & ~n94608;
  assign n94968 = ~n94595 & n94967;
  assign n94969 = n94589 & n94968;
  assign n94970 = ~n94966 & ~n94969;
  assign n94971 = ~n94963 & n94970;
  assign n94972 = n94620 & ~n94971;
  assign n94973 = ~n94962 & ~n94972;
  assign n94974 = n94595 & n94609;
  assign n94975 = ~n94589 & n94974;
  assign n94976 = ~n94602 & n94634;
  assign n94977 = ~n94975 & ~n94976;
  assign n94978 = ~n94583 & ~n94977;
  assign n94979 = n94602 & n94649;
  assign n94980 = ~n94602 & n94658;
  assign n94981 = ~n94979 & ~n94980;
  assign n94982 = n94583 & ~n94981;
  assign n94983 = ~n94596 & ~n94658;
  assign n94984 = n94602 & ~n94983;
  assign n94985 = ~n94634 & ~n94984;
  assign n94986 = ~n94583 & ~n94985;
  assign n94987 = n94595 & ~n94602;
  assign n94988 = n94959 & n94987;
  assign n94989 = ~n94595 & n94608;
  assign n94990 = ~n94634 & ~n94989;
  assign n94991 = ~n94602 & ~n94990;
  assign n94992 = n94583 & n94602;
  assign n94993 = n94624 & n94992;
  assign n94994 = ~n94608 & n94993;
  assign n94995 = ~n94991 & ~n94994;
  assign n94996 = ~n94988 & n94995;
  assign n94997 = ~n94986 & n94996;
  assign n94998 = ~n94975 & n94997;
  assign n94999 = ~n94620 & ~n94998;
  assign n95000 = ~n94982 & ~n94999;
  assign n95001 = ~n94978 & n95000;
  assign n95002 = n94973 & n95001;
  assign n95003 = pi3847 & n95002;
  assign n95004 = ~pi3847 & ~n95002;
  assign po3198 = n95003 | n95004;
  assign n95006 = ~n94835 & n94871;
  assign n95007 = ~n94892 & ~n95006;
  assign n95008 = n94841 & ~n95007;
  assign n95009 = ~n94835 & n94841;
  assign n95010 = n94883 & n95009;
  assign n95011 = ~n94853 & n95010;
  assign n95012 = ~n95008 & ~n95011;
  assign n95013 = ~n94862 & ~n95012;
  assign n95014 = ~n94835 & ~n94853;
  assign n95015 = ~n94869 & ~n94873;
  assign n95016 = n95014 & ~n95015;
  assign n95017 = ~n94854 & ~n94869;
  assign n95018 = ~n94835 & ~n95017;
  assign n95019 = ~n94878 & ~n95018;
  assign n95020 = ~n94841 & ~n95019;
  assign n95021 = ~n95016 & ~n95020;
  assign n95022 = n94835 & n94872;
  assign n95023 = ~n94835 & n94853;
  assign n95024 = n94868 & n95023;
  assign n95025 = n94835 & ~n95017;
  assign n95026 = ~n95024 & ~n95025;
  assign n95027 = n94841 & ~n95026;
  assign n95028 = ~n95022 & ~n95027;
  assign n95029 = n95021 & n95028;
  assign n95030 = n94862 & ~n95029;
  assign n95031 = ~n94869 & n94907;
  assign n95032 = ~n94862 & n95031;
  assign n95033 = n94835 & ~n94853;
  assign n95034 = n94869 & n95033;
  assign n95035 = n94841 & n95034;
  assign n95036 = n94835 & ~n94841;
  assign n95037 = n94853 & n95036;
  assign n95038 = n94868 & n95037;
  assign n95039 = ~n95035 & ~n95038;
  assign n95040 = ~n95032 & n95039;
  assign n95041 = n94835 & n94847;
  assign n95042 = ~n94896 & ~n95041;
  assign n95043 = ~n94841 & ~n94862;
  assign n95044 = ~n95042 & n95043;
  assign n95045 = n95040 & ~n95044;
  assign n95046 = ~n95030 & n95045;
  assign n95047 = ~n95013 & n95046;
  assign n95048 = pi3780 & ~n95047;
  assign n95049 = ~pi3780 & n95047;
  assign po3199 = n95048 | n95049;
  assign n95051 = n94841 & n94878;
  assign n95052 = ~n94835 & n95051;
  assign n95053 = ~n95011 & ~n95052;
  assign n95054 = ~n94841 & n94872;
  assign n95055 = ~n94835 & n95054;
  assign n95056 = ~n94835 & n94898;
  assign n95057 = ~n95055 & ~n95056;
  assign n95058 = n94847 & n94853;
  assign n95059 = n94835 & n95058;
  assign n95060 = n94835 & n94871;
  assign n95061 = ~n95059 & ~n95060;
  assign n95062 = n94841 & ~n95061;
  assign n95063 = ~n94841 & ~n95014;
  assign n95064 = ~n95015 & n95063;
  assign n95065 = ~n94871 & n95009;
  assign n95066 = ~n94853 & n95065;
  assign n95067 = ~n95064 & ~n95066;
  assign n95068 = ~n95062 & n95067;
  assign n95069 = n95057 & n95068;
  assign n95070 = ~n94862 & ~n95069;
  assign n95071 = n95053 & ~n95070;
  assign n95072 = ~n94841 & n94870;
  assign n95073 = n94835 & n95072;
  assign n95074 = ~n94841 & n94862;
  assign n95075 = ~n94884 & ~n95060;
  assign n95076 = ~n95016 & n95075;
  assign n95077 = n95074 & ~n95076;
  assign n95078 = n94835 & n94898;
  assign n95079 = ~n94853 & n95041;
  assign n95080 = ~n94892 & ~n95079;
  assign n95081 = ~n94896 & ~n95006;
  assign n95082 = n95080 & n95081;
  assign n95083 = n94841 & ~n95082;
  assign n95084 = ~n95078 & ~n95083;
  assign n95085 = n94862 & ~n95084;
  assign n95086 = ~n95077 & ~n95085;
  assign n95087 = ~n95073 & n95086;
  assign n95088 = n95071 & n95087;
  assign n95089 = pi3844 & ~n95088;
  assign n95090 = ~pi3844 & n95071;
  assign n95091 = n95087 & n95090;
  assign po3200 = n95089 | n95091;
  assign n95093 = ~n94868 & n95023;
  assign n95094 = n94899 & ~n95093;
  assign n95095 = n95043 & ~n95094;
  assign n95096 = ~n94862 & n94896;
  assign n95097 = n94835 & n95096;
  assign n95098 = ~n94853 & ~n94868;
  assign n95099 = ~n95060 & ~n95098;
  assign n95100 = n94841 & ~n95099;
  assign n95101 = ~n94885 & ~n95100;
  assign n95102 = ~n94862 & ~n95101;
  assign n95103 = ~n95097 & ~n95102;
  assign n95104 = ~n94868 & n95033;
  assign n95105 = ~n94886 & ~n95104;
  assign n95106 = n94841 & ~n95105;
  assign n95107 = n95103 & ~n95106;
  assign n95108 = n94871 & n95036;
  assign n95109 = n94853 & n95108;
  assign n95110 = ~n95015 & n95033;
  assign n95111 = ~n95109 & ~n95110;
  assign n95112 = ~n94909 & n95111;
  assign n95113 = ~n95015 & n95023;
  assign n95114 = ~n95056 & ~n95113;
  assign n95115 = n94853 & n95009;
  assign n95116 = ~n94847 & n95115;
  assign n95117 = ~n95055 & ~n95116;
  assign n95118 = n95114 & n95117;
  assign n95119 = n95112 & n95118;
  assign n95120 = n94862 & ~n95119;
  assign n95121 = n95107 & ~n95120;
  assign n95122 = ~n95095 & n95121;
  assign n95123 = ~pi3857 & ~n95122;
  assign n95124 = pi3857 & n95107;
  assign n95125 = ~n95095 & n95124;
  assign n95126 = ~n95120 & n95125;
  assign po3201 = n95123 | n95126;
  assign n95128 = ~n94423 & ~n94431;
  assign n95129 = n94370 & ~n95128;
  assign n95130 = ~n94394 & n94681;
  assign n95131 = ~n94682 & ~n95130;
  assign n95132 = ~n94396 & n95131;
  assign n95133 = ~n94403 & ~n95132;
  assign n95134 = n94370 & n95133;
  assign n95135 = ~n95129 & ~n95134;
  assign n95136 = n94422 & n94678;
  assign n95137 = ~n94680 & ~n95136;
  assign n95138 = ~n94439 & ~n94705;
  assign n95139 = n94403 & ~n95138;
  assign n95140 = n94370 & n95139;
  assign n95141 = n95137 & ~n95140;
  assign n95142 = n94376 & n94422;
  assign n95143 = n94376 & n94414;
  assign n95144 = ~n94670 & ~n95143;
  assign n95145 = n94403 & ~n95144;
  assign n95146 = ~n94437 & ~n94677;
  assign n95147 = n94376 & n94421;
  assign n95148 = ~n94461 & ~n95147;
  assign n95149 = ~n94403 & ~n95148;
  assign n95150 = n95146 & ~n95149;
  assign n95151 = ~n95145 & n95150;
  assign n95152 = ~n95142 & n95151;
  assign n95153 = ~n94370 & ~n95152;
  assign n95154 = ~n94702 & n94801;
  assign n95155 = n94403 & ~n95154;
  assign n95156 = ~n95153 & ~n95155;
  assign n95157 = n95141 & n95156;
  assign n95158 = n95135 & n95157;
  assign n95159 = ~pi3841 & ~n95158;
  assign n95160 = pi3841 & n95141;
  assign n95161 = n95135 & n95160;
  assign n95162 = n95156 & n95161;
  assign po3202 = n95159 | n95162;
  assign n95164 = ~n94595 & n94611;
  assign n95165 = ~n94641 & ~n95164;
  assign n95166 = ~n94583 & ~n95165;
  assign n95167 = ~n94589 & n94602;
  assign n95168 = n94595 & n95167;
  assign n95169 = ~n94968 & ~n95168;
  assign n95170 = n94583 & ~n95169;
  assign n95171 = ~n94602 & n94628;
  assign n95172 = ~n94988 & ~n95171;
  assign n95173 = ~n94610 & n95172;
  assign n95174 = ~n95170 & n95173;
  assign n95175 = ~n95166 & n95174;
  assign n95176 = ~n94963 & ~n94975;
  assign n95177 = n95175 & n95176;
  assign n95178 = n94620 & ~n95177;
  assign n95179 = n94596 & n94964;
  assign n95180 = n94650 & ~n95179;
  assign n95181 = n94583 & ~n95180;
  assign n95182 = ~n94602 & n94638;
  assign n95183 = ~n95181 & ~n95182;
  assign n95184 = n94589 & n94611;
  assign n95185 = n94602 & n94624;
  assign n95186 = ~n95184 & ~n95185;
  assign n95187 = n94583 & ~n95186;
  assign n95188 = n94583 & n94633;
  assign n95189 = ~n94602 & n95188;
  assign n95190 = ~n95187 & ~n95189;
  assign n95191 = n95183 & n95190;
  assign n95192 = ~n94620 & ~n95191;
  assign n95193 = ~n94628 & ~n94635;
  assign n95194 = ~n94969 & n95193;
  assign n95195 = n94655 & ~n95194;
  assign n95196 = ~n95192 & ~n95195;
  assign n95197 = ~n94610 & ~n94963;
  assign n95198 = ~n94583 & ~n95197;
  assign n95199 = n95196 & ~n95198;
  assign n95200 = ~n95178 & n95199;
  assign n95201 = ~pi3856 & n95200;
  assign n95202 = pi3856 & ~n95200;
  assign po3203 = n95201 | n95202;
  assign n95204 = ~n94229 & ~n94774;
  assign n95205 = ~n94762 & n95204;
  assign n95206 = n94198 & ~n95205;
  assign n95207 = ~n94240 & ~n94268;
  assign n95208 = ~n94237 & ~n94770;
  assign n95209 = ~n94220 & ~n94776;
  assign n95210 = ~n94198 & ~n95209;
  assign n95211 = ~n94296 & ~n95210;
  assign n95212 = n95208 & n95211;
  assign n95213 = n94186 & ~n95212;
  assign n95214 = ~n94212 & n94218;
  assign n95215 = ~n94276 & ~n95214;
  assign n95216 = n94192 & ~n95215;
  assign n95217 = ~n94246 & ~n94250;
  assign n95218 = ~n94198 & ~n95217;
  assign n95219 = n94192 & n94218;
  assign n95220 = ~n94227 & ~n95219;
  assign n95221 = ~n94219 & n95220;
  assign n95222 = n94198 & ~n95221;
  assign n95223 = ~n95218 & ~n95222;
  assign n95224 = ~n95216 & n95223;
  assign n95225 = ~n94186 & ~n95224;
  assign n95226 = ~n95213 & ~n95225;
  assign n95227 = n95207 & n95226;
  assign n95228 = ~n95206 & n95227;
  assign n95229 = ~pi3921 & ~n95228;
  assign n95230 = pi3921 & n95207;
  assign n95231 = ~n95206 & n95230;
  assign n95232 = n95226 & n95231;
  assign po3204 = n95229 | n95232;
  assign n95234 = ~n94602 & n94624;
  assign n95235 = ~n94623 & ~n95234;
  assign n95236 = ~n94583 & ~n95235;
  assign n95237 = n94583 & ~n94990;
  assign n95238 = ~n94979 & ~n95237;
  assign n95239 = ~n95236 & n95238;
  assign n95240 = n94620 & ~n95239;
  assign n95241 = ~n94583 & n94638;
  assign n95242 = ~n95240 & ~n95241;
  assign n95243 = ~n95171 & ~n95185;
  assign n95244 = n94583 & ~n95243;
  assign n95245 = n94583 & n94625;
  assign n95246 = n94602 & n94641;
  assign n95247 = ~n94583 & n94609;
  assign n95248 = ~n94967 & ~n95247;
  assign n95249 = ~n94589 & ~n95248;
  assign n95250 = ~n94968 & ~n95249;
  assign n95251 = ~n94610 & n95250;
  assign n95252 = ~n95246 & n95251;
  assign n95253 = ~n95245 & n95252;
  assign n95254 = ~n94620 & ~n95253;
  assign n95255 = ~n95244 & ~n95254;
  assign n95256 = n95242 & n95255;
  assign n95257 = pi3917 & ~n95256;
  assign n95258 = ~pi3917 & n95256;
  assign po3205 = n95257 | n95258;
  assign n95260 = pi7534 & ~pi9040;
  assign n95261 = pi7449 & pi9040;
  assign n95262 = ~n95260 & ~n95261;
  assign n95263 = ~pi3936 & ~n95262;
  assign n95264 = pi3936 & n95262;
  assign n95265 = ~n95263 & ~n95264;
  assign n95266 = pi7454 & pi9040;
  assign n95267 = pi7425 & ~pi9040;
  assign n95268 = ~n95266 & ~n95267;
  assign n95269 = ~pi3895 & ~n95268;
  assign n95270 = pi3895 & n95268;
  assign n95271 = ~n95269 & ~n95270;
  assign n95272 = pi7431 & ~pi9040;
  assign n95273 = pi7386 & pi9040;
  assign n95274 = ~n95272 & ~n95273;
  assign n95275 = pi3782 & n95274;
  assign n95276 = ~pi3782 & ~n95274;
  assign n95277 = ~n95275 & ~n95276;
  assign n95278 = pi7431 & pi9040;
  assign n95279 = pi7568 & ~pi9040;
  assign n95280 = ~n95278 & ~n95279;
  assign n95281 = ~pi3866 & ~n95280;
  assign n95282 = pi3866 & n95280;
  assign n95283 = ~n95281 & ~n95282;
  assign n95284 = pi7385 & ~pi9040;
  assign n95285 = pi7534 & pi9040;
  assign n95286 = ~n95284 & ~n95285;
  assign n95287 = pi3912 & n95286;
  assign n95288 = ~pi3912 & ~n95286;
  assign n95289 = ~n95287 & ~n95288;
  assign n95290 = ~n95283 & n95289;
  assign n95291 = n95277 & n95290;
  assign n95292 = pi7461 & ~pi9040;
  assign n95293 = pi7453 & pi9040;
  assign n95294 = ~n95292 & ~n95293;
  assign n95295 = ~pi3929 & ~n95294;
  assign n95296 = pi3929 & n95294;
  assign n95297 = ~n95295 & ~n95296;
  assign n95298 = n95283 & n95297;
  assign n95299 = n95289 & n95298;
  assign n95300 = ~n95291 & ~n95299;
  assign n95301 = n95283 & ~n95297;
  assign n95302 = ~n95289 & n95301;
  assign n95303 = ~n95277 & n95302;
  assign n95304 = n95300 & ~n95303;
  assign n95305 = n95271 & ~n95304;
  assign n95306 = n95283 & ~n95289;
  assign n95307 = n95297 & n95306;
  assign n95308 = ~n95277 & n95307;
  assign n95309 = ~n95283 & n95297;
  assign n95310 = n95289 & n95309;
  assign n95311 = ~n95277 & n95310;
  assign n95312 = ~n95283 & ~n95289;
  assign n95313 = ~n95301 & ~n95312;
  assign n95314 = n95277 & ~n95313;
  assign n95315 = ~n95311 & ~n95314;
  assign n95316 = ~n95308 & n95315;
  assign n95317 = ~n95271 & ~n95316;
  assign n95318 = ~n95305 & ~n95317;
  assign n95319 = n95265 & ~n95318;
  assign n95320 = n95271 & ~n95277;
  assign n95321 = ~n95283 & n95320;
  assign n95322 = ~n95271 & ~n95277;
  assign n95323 = n95301 & n95322;
  assign n95324 = ~n95277 & n95283;
  assign n95325 = n95289 & n95324;
  assign n95326 = ~n95291 & ~n95325;
  assign n95327 = ~n95271 & ~n95326;
  assign n95328 = ~n95323 & ~n95327;
  assign n95329 = n95271 & n95277;
  assign n95330 = n95306 & n95329;
  assign n95331 = ~n95289 & n95309;
  assign n95332 = n95271 & n95331;
  assign n95333 = ~n95330 & ~n95332;
  assign n95334 = n95289 & n95301;
  assign n95335 = ~n95277 & n95334;
  assign n95336 = n95277 & n95307;
  assign n95337 = ~n95335 & ~n95336;
  assign n95338 = n95333 & n95337;
  assign n95339 = n95328 & n95338;
  assign n95340 = ~n95321 & n95339;
  assign n95341 = ~n95265 & ~n95340;
  assign n95342 = ~n95271 & n95335;
  assign n95343 = ~n95283 & ~n95297;
  assign n95344 = ~n95289 & n95343;
  assign n95345 = ~n95271 & n95344;
  assign n95346 = ~n95277 & n95345;
  assign n95347 = ~n95342 & ~n95346;
  assign n95348 = ~n95277 & ~n95289;
  assign n95349 = n95297 & n95348;
  assign n95350 = ~n95283 & n95349;
  assign n95351 = n95271 & n95350;
  assign n95352 = n95347 & ~n95351;
  assign n95353 = n95289 & n95343;
  assign n95354 = ~n95277 & n95353;
  assign n95355 = n95277 & n95298;
  assign n95356 = ~n95354 & ~n95355;
  assign n95357 = n95271 & ~n95356;
  assign n95358 = n95352 & ~n95357;
  assign n95359 = ~n95341 & n95358;
  assign n95360 = ~n95319 & n95359;
  assign n95361 = ~pi5202 & ~n95360;
  assign n95362 = pi5202 & n95360;
  assign po3495 = n95361 | n95362;
  assign n95364 = pi7412 & pi9040;
  assign n95365 = pi7369 & ~pi9040;
  assign n95366 = ~n95364 & ~n95365;
  assign n95367 = pi3839 & n95366;
  assign n95368 = ~pi3839 & ~n95366;
  assign n95369 = ~n95367 & ~n95368;
  assign n95370 = pi7444 & ~pi9040;
  assign n95371 = pi7417 & pi9040;
  assign n95372 = ~n95370 & ~n95371;
  assign n95373 = ~pi3845 & n95372;
  assign n95374 = pi3845 & ~n95372;
  assign n95375 = ~n95373 & ~n95374;
  assign n95376 = pi7450 & ~pi9040;
  assign n95377 = pi7518 & pi9040;
  assign n95378 = ~n95376 & ~n95377;
  assign n95379 = ~pi3931 & n95378;
  assign n95380 = pi3931 & ~n95378;
  assign n95381 = ~n95379 & ~n95380;
  assign n95382 = pi7424 & pi9040;
  assign n95383 = pi7410 & ~pi9040;
  assign n95384 = ~n95382 & ~n95383;
  assign n95385 = pi3892 & n95384;
  assign n95386 = ~pi3892 & ~n95384;
  assign n95387 = ~n95385 & ~n95386;
  assign n95388 = ~n95381 & n95387;
  assign n95389 = n95375 & n95388;
  assign n95390 = pi7383 & ~pi9040;
  assign n95391 = pi7413 & pi9040;
  assign n95392 = ~n95390 & ~n95391;
  assign n95393 = ~pi3862 & ~n95392;
  assign n95394 = pi3862 & n95392;
  assign n95395 = ~n95393 & ~n95394;
  assign n95396 = n95389 & ~n95395;
  assign n95397 = n95381 & ~n95387;
  assign n95398 = n95375 & n95397;
  assign n95399 = ~n95395 & n95398;
  assign n95400 = ~n95396 & ~n95399;
  assign n95401 = ~n95375 & n95395;
  assign n95402 = n95397 & n95401;
  assign n95403 = ~n95381 & ~n95387;
  assign n95404 = n95375 & n95403;
  assign n95405 = n95395 & n95404;
  assign n95406 = ~n95402 & ~n95405;
  assign n95407 = n95400 & n95406;
  assign n95408 = n95369 & ~n95407;
  assign n95409 = n95381 & n95387;
  assign n95410 = n95375 & n95409;
  assign n95411 = n95395 & n95410;
  assign n95412 = ~n95404 & ~n95411;
  assign n95413 = n95369 & ~n95412;
  assign n95414 = ~n95369 & n95387;
  assign n95415 = ~n95395 & n95414;
  assign n95416 = ~n95375 & ~n95381;
  assign n95417 = n95395 & n95397;
  assign n95418 = ~n95416 & ~n95417;
  assign n95419 = ~n95369 & ~n95418;
  assign n95420 = ~n95415 & ~n95419;
  assign n95421 = ~n95375 & n95409;
  assign n95422 = ~n95395 & n95421;
  assign n95423 = n95420 & ~n95422;
  assign n95424 = n95387 & n95416;
  assign n95425 = n95395 & n95424;
  assign n95426 = n95423 & ~n95425;
  assign n95427 = ~n95413 & n95426;
  assign n95428 = pi7383 & pi9040;
  assign n95429 = pi7412 & ~pi9040;
  assign n95430 = ~n95428 & ~n95429;
  assign n95431 = ~pi3863 & ~n95430;
  assign n95432 = pi3863 & n95430;
  assign n95433 = ~n95431 & ~n95432;
  assign n95434 = ~n95427 & ~n95433;
  assign n95435 = n95375 & n95387;
  assign n95436 = ~n95369 & n95395;
  assign n95437 = n95433 & n95436;
  assign n95438 = n95435 & n95437;
  assign n95439 = n95375 & ~n95395;
  assign n95440 = ~n95387 & n95439;
  assign n95441 = ~n95369 & ~n95440;
  assign n95442 = n95381 & n95401;
  assign n95443 = ~n95388 & ~n95435;
  assign n95444 = ~n95395 & ~n95443;
  assign n95445 = ~n95375 & n95397;
  assign n95446 = ~n95444 & ~n95445;
  assign n95447 = ~n95442 & n95446;
  assign n95448 = n95369 & n95447;
  assign n95449 = ~n95441 & ~n95448;
  assign n95450 = ~n95387 & n95401;
  assign n95451 = ~n95381 & n95450;
  assign n95452 = ~n95449 & ~n95451;
  assign n95453 = n95433 & ~n95452;
  assign n95454 = ~n95438 & ~n95453;
  assign n95455 = ~n95434 & n95454;
  assign n95456 = ~n95408 & n95455;
  assign n95457 = ~n95369 & ~n95395;
  assign n95458 = n95409 & n95457;
  assign n95459 = ~n95375 & n95458;
  assign n95460 = n95456 & ~n95459;
  assign n95461 = pi5217 & ~n95460;
  assign n95462 = n95455 & ~n95459;
  assign n95463 = ~pi5217 & n95462;
  assign n95464 = ~n95408 & n95463;
  assign po3496 = n95461 | n95464;
  assign n95466 = pi7522 & pi9040;
  assign n95467 = pi7439 & ~pi9040;
  assign n95468 = ~n95466 & ~n95467;
  assign n95469 = pi3851 & n95468;
  assign n95470 = ~pi3851 & ~n95468;
  assign n95471 = ~n95469 & ~n95470;
  assign n95472 = pi7421 & ~pi9040;
  assign n95473 = pi7591 & pi9040;
  assign n95474 = ~n95472 & ~n95473;
  assign n95475 = ~pi3865 & ~n95474;
  assign n95476 = pi3865 & n95474;
  assign n95477 = ~n95475 & ~n95476;
  assign n95478 = pi7421 & pi9040;
  assign n95479 = pi7521 & ~pi9040;
  assign n95480 = ~n95478 & ~n95479;
  assign n95481 = ~pi3930 & n95480;
  assign n95482 = pi3930 & ~n95480;
  assign n95483 = ~n95481 & ~n95482;
  assign n95484 = n95477 & n95483;
  assign n95485 = pi7466 & pi9040;
  assign n95486 = pi7422 & ~pi9040;
  assign n95487 = ~n95485 & ~n95486;
  assign n95488 = ~pi3958 & n95487;
  assign n95489 = pi3958 & ~n95487;
  assign n95490 = ~n95488 & ~n95489;
  assign n95491 = pi7511 & pi9040;
  assign n95492 = pi7446 & ~pi9040;
  assign n95493 = ~n95491 & ~n95492;
  assign n95494 = ~pi3842 & ~n95493;
  assign n95495 = pi3842 & n95493;
  assign n95496 = ~n95494 & ~n95495;
  assign n95497 = ~n95490 & n95496;
  assign n95498 = n95484 & n95497;
  assign n95499 = ~n95490 & ~n95496;
  assign n95500 = ~n95477 & n95499;
  assign n95501 = ~n95498 & ~n95500;
  assign n95502 = ~n95471 & ~n95501;
  assign n95503 = pi7434 & pi9040;
  assign n95504 = pi7511 & ~pi9040;
  assign n95505 = ~n95503 & ~n95504;
  assign n95506 = ~pi3940 & ~n95505;
  assign n95507 = pi3940 & n95505;
  assign n95508 = ~n95506 & ~n95507;
  assign n95509 = n95471 & n95490;
  assign n95510 = n95477 & n95509;
  assign n95511 = n95484 & ~n95496;
  assign n95512 = n95477 & ~n95483;
  assign n95513 = n95496 & n95512;
  assign n95514 = ~n95511 & ~n95513;
  assign n95515 = ~n95477 & n95483;
  assign n95516 = n95496 & n95515;
  assign n95517 = ~n95490 & n95516;
  assign n95518 = n95514 & ~n95517;
  assign n95519 = n95471 & ~n95518;
  assign n95520 = ~n95510 & ~n95519;
  assign n95521 = ~n95477 & ~n95483;
  assign n95522 = ~n95496 & n95521;
  assign n95523 = ~n95490 & n95522;
  assign n95524 = n95520 & ~n95523;
  assign n95525 = n95490 & n95515;
  assign n95526 = ~n95477 & n95496;
  assign n95527 = ~n95483 & n95526;
  assign n95528 = ~n95525 & ~n95527;
  assign n95529 = ~n95471 & ~n95528;
  assign n95530 = ~n95496 & n95512;
  assign n95531 = n95490 & n95530;
  assign n95532 = ~n95529 & ~n95531;
  assign n95533 = n95524 & n95532;
  assign n95534 = n95508 & ~n95533;
  assign n95535 = ~n95502 & ~n95534;
  assign n95536 = n95471 & ~n95508;
  assign n95537 = ~n95528 & n95536;
  assign n95538 = ~n95496 & n95515;
  assign n95539 = ~n95530 & ~n95538;
  assign n95540 = ~n95490 & ~n95539;
  assign n95541 = ~n95498 & ~n95540;
  assign n95542 = ~n95508 & ~n95541;
  assign n95543 = ~n95537 & ~n95542;
  assign n95544 = ~n95471 & ~n95508;
  assign n95545 = n95484 & n95490;
  assign n95546 = ~n95522 & ~n95545;
  assign n95547 = n95477 & n95496;
  assign n95548 = n95546 & ~n95547;
  assign n95549 = n95544 & ~n95548;
  assign n95550 = n95543 & ~n95549;
  assign n95551 = n95535 & n95550;
  assign n95552 = ~pi5280 & ~n95551;
  assign n95553 = pi5280 & n95543;
  assign n95554 = n95535 & n95553;
  assign n95555 = ~n95549 & n95554;
  assign po3497 = n95552 | n95555;
  assign n95557 = pi7429 & pi9040;
  assign n95558 = pi7411 & ~pi9040;
  assign n95559 = ~n95557 & ~n95558;
  assign n95560 = ~pi3892 & ~n95559;
  assign n95561 = pi3892 & n95559;
  assign n95562 = ~n95560 & ~n95561;
  assign n95563 = pi7462 & pi9040;
  assign n95564 = pi7386 & ~pi9040;
  assign n95565 = ~n95563 & ~n95564;
  assign n95566 = ~pi3936 & n95565;
  assign n95567 = pi3936 & ~n95565;
  assign n95568 = ~n95566 & ~n95567;
  assign n95569 = pi7410 & pi9040;
  assign n95570 = pi7518 & ~pi9040;
  assign n95571 = ~n95569 & ~n95570;
  assign n95572 = ~pi3845 & n95571;
  assign n95573 = pi3845 & ~n95571;
  assign n95574 = ~n95572 & ~n95573;
  assign n95575 = n95568 & ~n95574;
  assign n95576 = pi7450 & pi9040;
  assign n95577 = pi7424 & ~pi9040;
  assign n95578 = ~n95576 & ~n95577;
  assign n95579 = ~pi3853 & n95578;
  assign n95580 = pi3853 & ~n95578;
  assign n95581 = ~n95579 & ~n95580;
  assign n95582 = pi7409 & pi9040;
  assign n95583 = pi7433 & ~pi9040;
  assign n95584 = ~n95582 & ~n95583;
  assign n95585 = ~pi3875 & ~n95584;
  assign n95586 = pi3875 & n95584;
  assign n95587 = ~n95585 & ~n95586;
  assign n95588 = n95581 & ~n95587;
  assign n95589 = n95575 & n95588;
  assign n95590 = pi7409 & ~pi9040;
  assign n95591 = pi7444 & pi9040;
  assign n95592 = ~n95590 & ~n95591;
  assign n95593 = ~pi3929 & ~n95592;
  assign n95594 = pi3929 & n95592;
  assign n95595 = ~n95593 & ~n95594;
  assign n95596 = ~n95568 & n95574;
  assign n95597 = n95595 & n95596;
  assign n95598 = ~n95581 & ~n95595;
  assign n95599 = n95574 & n95598;
  assign n95600 = n95568 & n95599;
  assign n95601 = ~n95597 & ~n95600;
  assign n95602 = ~n95568 & ~n95574;
  assign n95603 = ~n95581 & n95602;
  assign n95604 = n95601 & ~n95603;
  assign n95605 = ~n95587 & ~n95604;
  assign n95606 = ~n95568 & ~n95595;
  assign n95607 = n95581 & n95587;
  assign n95608 = n95606 & n95607;
  assign n95609 = ~n95595 & n95596;
  assign n95610 = n95581 & n95609;
  assign n95611 = ~n95608 & ~n95610;
  assign n95612 = ~n95605 & n95611;
  assign n95613 = ~n95589 & n95612;
  assign n95614 = n95595 & n95602;
  assign n95615 = ~n95581 & n95614;
  assign n95616 = n95575 & n95595;
  assign n95617 = n95581 & n95616;
  assign n95618 = ~n95615 & ~n95617;
  assign n95619 = n95613 & n95618;
  assign n95620 = ~n95562 & ~n95619;
  assign n95621 = n95581 & ~n95595;
  assign n95622 = ~n95574 & n95621;
  assign n95623 = ~n95568 & n95622;
  assign n95624 = ~n95616 & ~n95623;
  assign n95625 = ~n95587 & ~n95624;
  assign n95626 = n95575 & ~n95595;
  assign n95627 = ~n95581 & n95626;
  assign n95628 = n95574 & n95621;
  assign n95629 = n95568 & n95628;
  assign n95630 = ~n95627 & ~n95629;
  assign n95631 = ~n95568 & n95598;
  assign n95632 = n95581 & n95595;
  assign n95633 = ~n95574 & n95632;
  assign n95634 = ~n95568 & n95633;
  assign n95635 = ~n95631 & ~n95634;
  assign n95636 = n95587 & ~n95635;
  assign n95637 = n95630 & ~n95636;
  assign n95638 = ~n95625 & n95637;
  assign n95639 = n95562 & ~n95638;
  assign n95640 = ~n95568 & n95595;
  assign n95641 = ~n95581 & n95640;
  assign n95642 = n95568 & n95595;
  assign n95643 = n95581 & n95642;
  assign n95644 = ~n95641 & ~n95643;
  assign n95645 = ~n95587 & ~n95644;
  assign n95646 = n95568 & n95574;
  assign n95647 = n95595 & n95646;
  assign n95648 = ~n95581 & n95647;
  assign n95649 = ~n95609 & ~n95648;
  assign n95650 = ~n95627 & n95649;
  assign n95651 = n95587 & ~n95650;
  assign n95652 = ~n95645 & ~n95651;
  assign n95653 = n95574 & ~n95595;
  assign n95654 = n95587 & n95653;
  assign n95655 = n95581 & n95654;
  assign n95656 = n95652 & ~n95655;
  assign n95657 = ~n95639 & n95656;
  assign n95658 = ~n95620 & n95657;
  assign n95659 = ~pi5307 & ~n95658;
  assign n95660 = pi5307 & n95658;
  assign po3498 = n95659 | n95660;
  assign n95662 = pi7436 & pi9040;
  assign n95663 = pi7414 & ~pi9040;
  assign n95664 = ~n95662 & ~n95663;
  assign n95665 = pi3935 & n95664;
  assign n95666 = ~pi3935 & ~n95664;
  assign n95667 = ~n95665 & ~n95666;
  assign n95668 = pi7415 & pi9040;
  assign n95669 = pi7434 & ~pi9040;
  assign n95670 = ~n95668 & ~n95669;
  assign n95671 = pi3863 & n95670;
  assign n95672 = ~pi3863 & ~n95670;
  assign n95673 = ~n95671 & ~n95672;
  assign n95674 = pi7521 & pi9040;
  assign n95675 = pi7440 & ~pi9040;
  assign n95676 = ~n95674 & ~n95675;
  assign n95677 = ~pi3931 & n95676;
  assign n95678 = pi3931 & ~n95676;
  assign n95679 = ~n95677 & ~n95678;
  assign n95680 = pi7379 & ~pi9040;
  assign n95681 = pi7396 & pi9040;
  assign n95682 = ~n95680 & ~n95681;
  assign n95683 = ~pi3842 & n95682;
  assign n95684 = pi3842 & ~n95682;
  assign n95685 = ~n95683 & ~n95684;
  assign n95686 = n95679 & n95685;
  assign n95687 = n95673 & n95686;
  assign n95688 = ~n95667 & n95687;
  assign n95689 = pi7440 & pi9040;
  assign n95690 = pi7591 & ~pi9040;
  assign n95691 = ~n95689 & ~n95690;
  assign n95692 = ~pi3989 & n95691;
  assign n95693 = pi3989 & ~n95691;
  assign n95694 = ~n95692 & ~n95693;
  assign n95695 = n95673 & ~n95679;
  assign n95696 = n95694 & n95695;
  assign n95697 = n95667 & ~n95673;
  assign n95698 = n95679 & n95697;
  assign n95699 = ~n95696 & ~n95698;
  assign n95700 = ~n95673 & ~n95685;
  assign n95701 = n95679 & n95700;
  assign n95702 = n95699 & ~n95701;
  assign n95703 = ~n95688 & n95702;
  assign n95704 = ~n95694 & n95700;
  assign n95705 = ~n95667 & n95704;
  assign n95706 = ~n95673 & n95685;
  assign n95707 = n95667 & n95706;
  assign n95708 = n95679 & ~n95685;
  assign n95709 = ~n95707 & ~n95708;
  assign n95710 = ~n95694 & ~n95709;
  assign n95711 = ~n95705 & ~n95710;
  assign n95712 = n95703 & n95711;
  assign n95713 = pi7575 & pi9040;
  assign n95714 = pi7430 & ~pi9040;
  assign n95715 = ~n95713 & ~n95714;
  assign n95716 = ~pi3865 & ~n95715;
  assign n95717 = pi3865 & n95715;
  assign n95718 = ~n95716 & ~n95717;
  assign n95719 = ~n95712 & n95718;
  assign n95720 = n95667 & n95694;
  assign n95721 = n95687 & n95720;
  assign n95722 = ~n95667 & ~n95679;
  assign n95723 = ~n95673 & n95722;
  assign n95724 = ~n95667 & ~n95673;
  assign n95725 = n95685 & n95724;
  assign n95726 = ~n95723 & ~n95725;
  assign n95727 = n95694 & ~n95726;
  assign n95728 = ~n95721 & ~n95727;
  assign n95729 = ~n95718 & ~n95728;
  assign n95730 = n95667 & n95679;
  assign n95731 = ~n95694 & n95730;
  assign n95732 = n95706 & n95731;
  assign n95733 = n95667 & ~n95694;
  assign n95734 = n95700 & n95733;
  assign n95735 = ~n95679 & n95734;
  assign n95736 = n95673 & ~n95685;
  assign n95737 = ~n95667 & ~n95694;
  assign n95738 = n95736 & n95737;
  assign n95739 = n95685 & n95722;
  assign n95740 = ~n95673 & n95739;
  assign n95741 = n95673 & n95685;
  assign n95742 = ~n95679 & n95741;
  assign n95743 = ~n95694 & n95742;
  assign n95744 = n95667 & n95743;
  assign n95745 = ~n95740 & ~n95744;
  assign n95746 = ~n95738 & n95745;
  assign n95747 = ~n95735 & n95746;
  assign n95748 = ~n95667 & n95736;
  assign n95749 = n95679 & n95748;
  assign n95750 = n95747 & ~n95749;
  assign n95751 = ~n95718 & ~n95750;
  assign n95752 = ~n95685 & n95695;
  assign n95753 = n95667 & n95752;
  assign n95754 = ~n95739 & ~n95753;
  assign n95755 = n95667 & n95701;
  assign n95756 = n95754 & ~n95755;
  assign n95757 = n95694 & ~n95756;
  assign n95758 = ~n95751 & ~n95757;
  assign n95759 = ~n95732 & n95758;
  assign n95760 = ~n95729 & n95759;
  assign n95761 = ~n95719 & n95760;
  assign n95762 = n95673 & n95679;
  assign n95763 = n95737 & n95762;
  assign n95764 = n95761 & ~n95763;
  assign n95765 = ~pi5238 & ~n95764;
  assign n95766 = pi5238 & ~n95763;
  assign n95767 = n95760 & n95766;
  assign n95768 = ~n95719 & n95767;
  assign po3499 = n95765 | n95768;
  assign n95770 = pi7537 & ~pi9040;
  assign n95771 = pi7397 & pi9040;
  assign n95772 = ~n95770 & ~n95771;
  assign n95773 = ~pi3939 & ~n95772;
  assign n95774 = pi3939 & n95772;
  assign n95775 = ~n95773 & ~n95774;
  assign n95776 = pi7537 & pi9040;
  assign n95777 = pi7522 & ~pi9040;
  assign n95778 = ~n95776 & ~n95777;
  assign n95779 = pi3960 & n95778;
  assign n95780 = ~pi3960 & ~n95778;
  assign n95781 = ~n95779 & ~n95780;
  assign n95782 = pi7446 & pi9040;
  assign n95783 = pi7415 & ~pi9040;
  assign n95784 = ~n95782 & ~n95783;
  assign n95785 = ~pi3943 & ~n95784;
  assign n95786 = pi3943 & n95784;
  assign n95787 = ~n95785 & ~n95786;
  assign n95788 = pi7456 & ~pi9040;
  assign n95789 = pi7460 & pi9040;
  assign n95790 = ~n95788 & ~n95789;
  assign n95791 = ~pi3915 & n95790;
  assign n95792 = pi3915 & ~n95790;
  assign n95793 = ~n95791 & ~n95792;
  assign n95794 = pi7519 & pi9040;
  assign n95795 = pi7528 & ~pi9040;
  assign n95796 = ~n95794 & ~n95795;
  assign n95797 = ~pi3840 & n95796;
  assign n95798 = pi3840 & ~n95796;
  assign n95799 = ~n95797 & ~n95798;
  assign n95800 = n95793 & n95799;
  assign n95801 = ~n95787 & n95800;
  assign n95802 = ~n95781 & n95801;
  assign n95803 = n95793 & ~n95799;
  assign n95804 = ~n95787 & n95803;
  assign n95805 = n95781 & n95804;
  assign n95806 = ~n95802 & ~n95805;
  assign n95807 = n95775 & ~n95806;
  assign n95808 = pi7439 & pi9040;
  assign n95809 = pi7397 & ~pi9040;
  assign n95810 = ~n95808 & ~n95809;
  assign n95811 = ~pi3870 & ~n95810;
  assign n95812 = pi3870 & n95810;
  assign n95813 = ~n95811 & ~n95812;
  assign n95814 = ~n95781 & n95787;
  assign n95815 = ~n95793 & n95814;
  assign n95816 = n95799 & n95815;
  assign n95817 = n95787 & n95803;
  assign n95818 = n95775 & n95817;
  assign n95819 = ~n95816 & ~n95818;
  assign n95820 = ~n95781 & ~n95799;
  assign n95821 = ~n95787 & n95820;
  assign n95822 = n95799 & n95814;
  assign n95823 = ~n95821 & ~n95822;
  assign n95824 = ~n95775 & ~n95823;
  assign n95825 = ~n95775 & n95781;
  assign n95826 = n95800 & n95825;
  assign n95827 = ~n95787 & n95826;
  assign n95828 = n95775 & ~n95787;
  assign n95829 = ~n95793 & n95828;
  assign n95830 = n95799 & n95829;
  assign n95831 = ~n95793 & ~n95799;
  assign n95832 = n95787 & n95831;
  assign n95833 = n95781 & n95832;
  assign n95834 = ~n95830 & ~n95833;
  assign n95835 = ~n95827 & n95834;
  assign n95836 = ~n95824 & n95835;
  assign n95837 = n95819 & n95836;
  assign n95838 = n95813 & ~n95837;
  assign n95839 = ~n95775 & n95816;
  assign n95840 = ~n95781 & n95818;
  assign n95841 = ~n95839 & ~n95840;
  assign n95842 = ~n95838 & n95841;
  assign n95843 = ~n95807 & n95842;
  assign n95844 = n95775 & n95781;
  assign n95845 = n95787 & n95799;
  assign n95846 = n95844 & n95845;
  assign n95847 = n95775 & n95801;
  assign n95848 = ~n95846 & ~n95847;
  assign n95849 = n95775 & n95832;
  assign n95850 = ~n95787 & n95831;
  assign n95851 = ~n95781 & n95850;
  assign n95852 = ~n95849 & ~n95851;
  assign n95853 = n95781 & n95787;
  assign n95854 = n95793 & n95853;
  assign n95855 = n95799 & n95854;
  assign n95856 = ~n95802 & ~n95855;
  assign n95857 = n95781 & n95803;
  assign n95858 = ~n95787 & ~n95793;
  assign n95859 = ~n95857 & ~n95858;
  assign n95860 = ~n95775 & ~n95859;
  assign n95861 = n95856 & ~n95860;
  assign n95862 = n95852 & n95861;
  assign n95863 = n95848 & n95862;
  assign n95864 = ~n95813 & ~n95863;
  assign n95865 = n95843 & ~n95864;
  assign n95866 = ~pi5216 & ~n95865;
  assign n95867 = pi5216 & n95843;
  assign n95868 = ~n95864 & n95867;
  assign po3500 = n95866 | n95868;
  assign n95870 = ~n95265 & ~n95271;
  assign n95871 = ~n95277 & n95290;
  assign n95872 = n95277 & n95334;
  assign n95873 = ~n95277 & n95298;
  assign n95874 = ~n95872 & ~n95873;
  assign n95875 = ~n95871 & n95874;
  assign n95876 = n95870 & ~n95875;
  assign n95877 = ~n95297 & n95348;
  assign n95878 = n95277 & n95353;
  assign n95879 = ~n95877 & ~n95878;
  assign n95880 = ~n95299 & ~n95302;
  assign n95881 = n95879 & n95880;
  assign n95882 = n95271 & ~n95881;
  assign n95883 = n95277 & ~n95289;
  assign n95884 = n95297 & n95883;
  assign n95885 = ~n95283 & n95884;
  assign n95886 = ~n95882 & ~n95885;
  assign n95887 = ~n95265 & ~n95886;
  assign n95888 = ~n95876 & ~n95887;
  assign n95889 = n95289 & n95320;
  assign n95890 = n95297 & n95889;
  assign n95891 = ~n95303 & ~n95890;
  assign n95892 = ~n95298 & ~n95343;
  assign n95893 = n95277 & ~n95892;
  assign n95894 = ~n95344 & ~n95893;
  assign n95895 = ~n95271 & ~n95894;
  assign n95896 = ~n95310 & ~n95871;
  assign n95897 = ~n95872 & n95896;
  assign n95898 = n95271 & ~n95897;
  assign n95899 = ~n95895 & ~n95898;
  assign n95900 = n95277 & n95344;
  assign n95901 = ~n95336 & ~n95900;
  assign n95902 = ~n95350 & n95901;
  assign n95903 = ~n95323 & n95902;
  assign n95904 = n95899 & n95903;
  assign n95905 = n95265 & ~n95904;
  assign n95906 = n95891 & ~n95905;
  assign n95907 = n95888 & n95906;
  assign n95908 = pi5191 & ~n95907;
  assign n95909 = ~pi5191 & n95891;
  assign n95910 = n95888 & n95909;
  assign n95911 = ~n95905 & n95910;
  assign po3502 = n95908 | n95911;
  assign n95913 = ~n95793 & n95799;
  assign n95914 = n95787 & n95913;
  assign n95915 = n95781 & n95914;
  assign n95916 = n95781 & n95831;
  assign n95917 = ~n95787 & n95913;
  assign n95918 = ~n95781 & n95917;
  assign n95919 = ~n95916 & ~n95918;
  assign n95920 = ~n95775 & ~n95919;
  assign n95921 = ~n95915 & ~n95920;
  assign n95922 = n95775 & n95913;
  assign n95923 = n95781 & n95922;
  assign n95924 = ~n95847 & ~n95923;
  assign n95925 = n95921 & n95924;
  assign n95926 = n95781 & n95817;
  assign n95927 = n95787 & n95800;
  assign n95928 = ~n95781 & n95927;
  assign n95929 = ~n95926 & ~n95928;
  assign n95930 = n95925 & n95929;
  assign n95931 = n95813 & ~n95930;
  assign n95932 = ~n95775 & ~n95813;
  assign n95933 = n95781 & ~n95787;
  assign n95934 = n95799 & n95933;
  assign n95935 = ~n95787 & n95793;
  assign n95936 = ~n95934 & ~n95935;
  assign n95937 = n95932 & ~n95936;
  assign n95938 = ~n95816 & ~n95821;
  assign n95939 = n95787 & n95844;
  assign n95940 = ~n95913 & n95939;
  assign n95941 = ~n95818 & ~n95940;
  assign n95942 = n95938 & n95941;
  assign n95943 = ~n95813 & ~n95942;
  assign n95944 = ~n95775 & n95804;
  assign n95945 = ~n95781 & n95944;
  assign n95946 = ~n95781 & n95832;
  assign n95947 = ~n95928 & ~n95946;
  assign n95948 = ~n95775 & ~n95947;
  assign n95949 = ~n95945 & ~n95948;
  assign n95950 = n95775 & n95816;
  assign n95951 = n95949 & ~n95950;
  assign n95952 = ~n95943 & n95951;
  assign n95953 = ~n95937 & n95952;
  assign n95954 = ~n95931 & n95953;
  assign n95955 = n95775 & ~n95781;
  assign n95956 = n95850 & n95955;
  assign n95957 = n95954 & ~n95956;
  assign n95958 = ~pi5350 & ~n95957;
  assign n95959 = pi5350 & ~n95956;
  assign n95960 = n95953 & n95959;
  assign n95961 = ~n95931 & n95960;
  assign po3539 = n95958 | n95961;
  assign n95963 = pi7427 & ~pi9040;
  assign n95964 = pi7385 & pi9040;
  assign n95965 = ~n95963 & ~n95964;
  assign n95966 = ~pi3866 & ~n95965;
  assign n95967 = pi3866 & n95965;
  assign n95968 = ~n95966 & ~n95967;
  assign n95969 = pi7376 & pi9040;
  assign n95970 = pi7589 & ~pi9040;
  assign n95971 = ~n95969 & ~n95970;
  assign n95972 = pi3972 & n95971;
  assign n95973 = ~pi3972 & ~n95971;
  assign n95974 = ~n95972 & ~n95973;
  assign n95975 = pi7411 & pi9040;
  assign n95976 = pi7453 & ~pi9040;
  assign n95977 = ~n95975 & ~n95976;
  assign n95978 = ~pi3870 & ~n95977;
  assign n95979 = pi3870 & n95977;
  assign n95980 = ~n95978 & ~n95979;
  assign n95981 = pi7376 & ~pi9040;
  assign n95982 = pi7425 & pi9040;
  assign n95983 = ~n95981 & ~n95982;
  assign n95984 = ~pi3915 & ~n95983;
  assign n95985 = pi3915 & n95983;
  assign n95986 = ~n95984 & ~n95985;
  assign n95987 = pi7461 & pi9040;
  assign n95988 = pi7429 & ~pi9040;
  assign n95989 = ~n95987 & ~n95988;
  assign n95990 = pi3912 & n95989;
  assign n95991 = ~pi3912 & ~n95989;
  assign n95992 = ~n95990 & ~n95991;
  assign n95993 = n95986 & ~n95992;
  assign n95994 = n95980 & n95993;
  assign n95995 = n95974 & n95994;
  assign n95996 = ~pi3912 & n95989;
  assign n95997 = pi3912 & ~n95989;
  assign n95998 = ~n95996 & ~n95997;
  assign n95999 = ~n95974 & n95986;
  assign n96000 = ~n95998 & n95999;
  assign n96001 = pi7568 & pi9040;
  assign n96002 = pi7462 & ~pi9040;
  assign n96003 = ~n96001 & ~n96002;
  assign n96004 = ~pi3861 & n96003;
  assign n96005 = pi3861 & ~n96003;
  assign n96006 = ~n96004 & ~n96005;
  assign n96007 = ~n95980 & n95999;
  assign n96008 = n95980 & ~n95998;
  assign n96009 = ~n95986 & n96008;
  assign n96010 = ~n96007 & ~n96009;
  assign n96011 = n96006 & ~n96010;
  assign n96012 = ~n96000 & ~n96011;
  assign n96013 = n95986 & n96008;
  assign n96014 = ~n95980 & ~n95986;
  assign n96015 = ~n95974 & ~n95986;
  assign n96016 = n95998 & n96015;
  assign n96017 = ~n95980 & ~n95992;
  assign n96018 = n95974 & n96017;
  assign n96019 = ~n96016 & ~n96018;
  assign n96020 = ~n96014 & n96019;
  assign n96021 = ~n96013 & n96020;
  assign n96022 = ~n96006 & ~n96021;
  assign n96023 = n96012 & ~n96022;
  assign n96024 = ~n95995 & n96023;
  assign n96025 = n95968 & ~n96024;
  assign n96026 = ~n95980 & ~n95998;
  assign n96027 = ~n95986 & n96026;
  assign n96028 = ~n95974 & n96027;
  assign n96029 = ~n95986 & n96017;
  assign n96030 = n95974 & n96029;
  assign n96031 = ~n95995 & ~n96030;
  assign n96032 = ~n96028 & n96031;
  assign n96033 = ~n96006 & ~n96032;
  assign n96034 = ~n96025 & ~n96033;
  assign n96035 = n95980 & n96000;
  assign n96036 = n95980 & ~n95986;
  assign n96037 = n96006 & n96036;
  assign n96038 = n95974 & n96037;
  assign n96039 = ~n95974 & ~n96006;
  assign n96040 = n95993 & n96039;
  assign n96041 = n95986 & n96026;
  assign n96042 = n95974 & n96041;
  assign n96043 = ~n96040 & ~n96042;
  assign n96044 = ~n95974 & n96006;
  assign n96045 = n96014 & n96044;
  assign n96046 = ~n95980 & n95986;
  assign n96047 = n95974 & n96046;
  assign n96048 = n95980 & ~n95992;
  assign n96049 = ~n95986 & n96048;
  assign n96050 = ~n96047 & ~n96049;
  assign n96051 = n96006 & ~n96050;
  assign n96052 = ~n96045 & ~n96051;
  assign n96053 = n96043 & n96052;
  assign n96054 = ~n95968 & ~n96053;
  assign n96055 = ~n96038 & ~n96054;
  assign n96056 = ~n96035 & n96055;
  assign n96057 = n96034 & n96056;
  assign n96058 = ~pi5098 & ~n96057;
  assign n96059 = ~n96025 & ~n96035;
  assign n96060 = ~n96033 & n96059;
  assign n96061 = n96055 & n96060;
  assign n96062 = pi5098 & n96061;
  assign po3540 = n96058 | n96062;
  assign n96064 = ~n95629 & ~n95640;
  assign n96065 = n95587 & ~n96064;
  assign n96066 = ~n95581 & n95609;
  assign n96067 = ~n96065 & ~n96066;
  assign n96068 = ~n95623 & n96067;
  assign n96069 = ~n95587 & n95627;
  assign n96070 = ~n95617 & ~n96069;
  assign n96071 = ~n95648 & n96070;
  assign n96072 = n96068 & n96071;
  assign n96073 = n95562 & ~n96072;
  assign n96074 = ~n95595 & n95602;
  assign n96075 = ~n95581 & n96074;
  assign n96076 = ~n95600 & ~n96075;
  assign n96077 = n95587 & n95626;
  assign n96078 = ~n95581 & n95616;
  assign n96079 = ~n96077 & ~n96078;
  assign n96080 = ~n95574 & n95595;
  assign n96081 = ~n95568 & ~n95581;
  assign n96082 = ~n96080 & ~n96081;
  assign n96083 = ~n95653 & n96082;
  assign n96084 = ~n95587 & ~n96083;
  assign n96085 = n95581 & n95647;
  assign n96086 = ~n95610 & ~n96085;
  assign n96087 = ~n96084 & n96086;
  assign n96088 = n96079 & n96087;
  assign n96089 = n96076 & n96088;
  assign n96090 = ~n95562 & ~n96089;
  assign n96091 = ~n96073 & ~n96090;
  assign n96092 = pi5183 & ~n96091;
  assign n96093 = ~pi5183 & ~n96073;
  assign n96094 = ~n96090 & n96093;
  assign po3541 = n96092 | n96094;
  assign n96096 = ~n95310 & ~n95344;
  assign n96097 = ~n95271 & ~n96096;
  assign n96098 = n95277 & n95299;
  assign n96099 = ~n96097 & ~n96098;
  assign n96100 = n95277 & n95283;
  assign n96101 = ~n95306 & ~n96100;
  assign n96102 = ~n95353 & n96101;
  assign n96103 = n95271 & ~n96102;
  assign n96104 = n96099 & ~n96103;
  assign n96105 = ~n95265 & ~n96104;
  assign n96106 = ~n95271 & n95308;
  assign n96107 = ~n95342 & ~n96106;
  assign n96108 = ~n95351 & n96107;
  assign n96109 = ~n95277 & n95289;
  assign n96110 = ~n95297 & n96109;
  assign n96111 = ~n95350 & ~n96110;
  assign n96112 = n95271 & n95325;
  assign n96113 = n95277 & n95310;
  assign n96114 = ~n95271 & n95306;
  assign n96115 = ~n96113 & ~n96114;
  assign n96116 = ~n95900 & n96115;
  assign n96117 = ~n96112 & n96116;
  assign n96118 = n96111 & n96117;
  assign n96119 = ~n95332 & n96118;
  assign n96120 = n95265 & ~n96119;
  assign n96121 = n96108 & ~n96120;
  assign n96122 = ~n96105 & n96121;
  assign n96123 = ~pi5428 & ~n96122;
  assign n96124 = pi5428 & n96108;
  assign n96125 = ~n96105 & n96124;
  assign n96126 = ~n96120 & n96125;
  assign po3544 = n96123 | n96126;
  assign n96128 = n95271 & n95298;
  assign n96129 = ~n95277 & n96128;
  assign n96130 = ~n95354 & ~n96129;
  assign n96131 = n95277 & n95289;
  assign n96132 = n95297 & n96131;
  assign n96133 = ~n95277 & ~n95283;
  assign n96134 = ~n96110 & ~n96133;
  assign n96135 = ~n95271 & ~n96134;
  assign n96136 = ~n96132 & ~n96135;
  assign n96137 = n96130 & n96136;
  assign n96138 = n95265 & ~n96137;
  assign n96139 = ~n95334 & ~n95336;
  assign n96140 = ~n95277 & n95309;
  assign n96141 = n96139 & ~n96140;
  assign n96142 = n95271 & ~n96141;
  assign n96143 = n95298 & n95322;
  assign n96144 = ~n95303 & ~n96143;
  assign n96145 = ~n96142 & n96144;
  assign n96146 = ~n95353 & ~n95885;
  assign n96147 = ~n95271 & ~n96146;
  assign n96148 = n96145 & ~n96147;
  assign n96149 = ~n95265 & ~n96148;
  assign n96150 = ~n96138 & ~n96149;
  assign n96151 = n95277 & n95880;
  assign n96152 = ~n95277 & ~n95343;
  assign n96153 = ~n96151 & ~n96152;
  assign n96154 = ~n95271 & n96153;
  assign n96155 = ~n95334 & n96096;
  assign n96156 = n95329 & ~n96155;
  assign n96157 = ~n96154 & ~n96156;
  assign n96158 = n96150 & n96157;
  assign n96159 = ~pi5426 & ~n96158;
  assign n96160 = ~n96149 & n96157;
  assign n96161 = pi5426 & n96160;
  assign n96162 = ~n96138 & n96161;
  assign po3554 = n96159 | n96162;
  assign n96164 = ~n95926 & ~n95934;
  assign n96165 = n95813 & ~n96164;
  assign n96166 = ~n95815 & ~n95822;
  assign n96167 = ~n95914 & n96166;
  assign n96168 = ~n95775 & ~n96167;
  assign n96169 = n95813 & n96168;
  assign n96170 = ~n96165 & ~n96169;
  assign n96171 = n95817 & n95825;
  assign n96172 = ~n95827 & ~n96171;
  assign n96173 = ~n95821 & ~n95858;
  assign n96174 = n95775 & ~n96173;
  assign n96175 = n95813 & n96174;
  assign n96176 = n96172 & ~n96175;
  assign n96177 = n95793 & n95814;
  assign n96178 = ~n95799 & n96177;
  assign n96179 = ~n95781 & n95800;
  assign n96180 = ~n95805 & ~n96179;
  assign n96181 = n95775 & ~n96180;
  assign n96182 = ~n95816 & ~n95833;
  assign n96183 = ~n95781 & n95803;
  assign n96184 = ~n95850 & ~n96183;
  assign n96185 = ~n95775 & ~n96184;
  assign n96186 = n96182 & ~n96185;
  assign n96187 = ~n96181 & n96186;
  assign n96188 = ~n96178 & n96187;
  assign n96189 = ~n95813 & ~n96188;
  assign n96190 = n95781 & n95917;
  assign n96191 = ~n95833 & ~n96190;
  assign n96192 = ~n95855 & n96191;
  assign n96193 = n95775 & ~n96192;
  assign n96194 = ~n96189 & ~n96193;
  assign n96195 = n96176 & n96194;
  assign n96196 = n96170 & n96195;
  assign n96197 = ~pi5427 & ~n96196;
  assign n96198 = pi5427 & n96176;
  assign n96199 = n96170 & n96198;
  assign n96200 = n96194 & n96199;
  assign po3555 = n96197 | n96200;
  assign n96202 = ~n95673 & ~n95679;
  assign n96203 = ~n95749 & ~n96202;
  assign n96204 = ~n95697 & n96203;
  assign n96205 = ~n95694 & ~n96204;
  assign n96206 = n95673 & n95720;
  assign n96207 = n95667 & ~n95679;
  assign n96208 = ~n95685 & n96207;
  assign n96209 = ~n95667 & n95742;
  assign n96210 = ~n96208 & ~n96209;
  assign n96211 = ~n95673 & n95679;
  assign n96212 = ~n95667 & n95694;
  assign n96213 = n96211 & n96212;
  assign n96214 = n96210 & ~n96213;
  assign n96215 = ~n96206 & n96214;
  assign n96216 = ~n96205 & n96215;
  assign n96217 = n95718 & ~n96216;
  assign n96218 = ~n95679 & n95706;
  assign n96219 = n95667 & n96218;
  assign n96220 = ~n95679 & n95700;
  assign n96221 = ~n95667 & n96220;
  assign n96222 = ~n96219 & ~n96221;
  assign n96223 = ~n95694 & ~n96222;
  assign n96224 = ~n96217 & ~n96223;
  assign n96225 = n95667 & n95742;
  assign n96226 = ~n95687 & ~n95752;
  assign n96227 = ~n95694 & ~n96226;
  assign n96228 = ~n96225 & ~n96227;
  assign n96229 = ~n95755 & n96228;
  assign n96230 = ~n95718 & ~n96229;
  assign n96231 = ~n95706 & ~n95736;
  assign n96232 = n95679 & ~n96231;
  assign n96233 = ~n95725 & ~n96232;
  assign n96234 = n95694 & ~n96233;
  assign n96235 = ~n95718 & n96234;
  assign n96236 = ~n96230 & ~n96235;
  assign n96237 = n96224 & n96236;
  assign n96238 = pi5499 & ~n96237;
  assign n96239 = ~pi5499 & n96224;
  assign n96240 = n96236 & n96239;
  assign po3556 = n96238 | n96240;
  assign n96242 = n95581 & n95602;
  assign n96243 = ~n96085 & ~n96242;
  assign n96244 = n95587 & n96243;
  assign n96245 = ~n95581 & n95642;
  assign n96246 = ~n95575 & ~n95596;
  assign n96247 = n95595 & ~n96246;
  assign n96248 = n95568 & n95621;
  assign n96249 = ~n95581 & n95596;
  assign n96250 = ~n96248 & ~n96249;
  assign n96251 = ~n95587 & n96250;
  assign n96252 = ~n96247 & n96251;
  assign n96253 = ~n96245 & n96252;
  assign n96254 = ~n96244 & ~n96253;
  assign n96255 = ~n95581 & n96247;
  assign n96256 = ~n96075 & ~n96255;
  assign n96257 = ~n96254 & n96256;
  assign n96258 = n95562 & ~n96257;
  assign n96259 = n95587 & ~n96246;
  assign n96260 = n95581 & n96259;
  assign n96261 = ~n95581 & n95646;
  assign n96262 = ~n95615 & ~n96261;
  assign n96263 = n95587 & ~n96262;
  assign n96264 = ~n95595 & n96259;
  assign n96265 = ~n96263 & ~n96264;
  assign n96266 = ~n96260 & n96265;
  assign n96267 = ~n95562 & ~n96266;
  assign n96268 = ~n96258 & ~n96267;
  assign n96269 = ~n95587 & ~n96243;
  assign n96270 = ~n95600 & ~n96269;
  assign n96271 = ~n95562 & ~n96270;
  assign n96272 = n95587 & n95600;
  assign n96273 = ~n95587 & ~n96256;
  assign n96274 = ~n96272 & ~n96273;
  assign n96275 = ~n96271 & n96274;
  assign n96276 = n96268 & n96275;
  assign n96277 = pi5349 & ~n96276;
  assign n96278 = ~pi5349 & n96275;
  assign n96279 = ~n96267 & n96278;
  assign n96280 = ~n96258 & n96279;
  assign po3557 = n96277 | n96280;
  assign n96282 = ~n95840 & ~n95846;
  assign n96283 = ~n95802 & n96191;
  assign n96284 = ~n95775 & ~n96283;
  assign n96285 = n95775 & n95927;
  assign n96286 = ~n95956 & n96191;
  assign n96287 = ~n95804 & ~n95816;
  assign n96288 = ~n95857 & n96287;
  assign n96289 = ~n95775 & ~n96288;
  assign n96290 = n96286 & ~n96289;
  assign n96291 = ~n96285 & n96290;
  assign n96292 = n95813 & ~n96291;
  assign n96293 = ~n95781 & n95922;
  assign n96294 = ~n95799 & n95933;
  assign n96295 = ~n95804 & ~n96294;
  assign n96296 = n95775 & ~n96295;
  assign n96297 = ~n96293 & ~n96296;
  assign n96298 = ~n95775 & n95831;
  assign n96299 = ~n95781 & n96298;
  assign n96300 = ~n95775 & n95801;
  assign n96301 = ~n96299 & ~n96300;
  assign n96302 = n96297 & n96301;
  assign n96303 = ~n95799 & n95814;
  assign n96304 = ~n95802 & ~n96303;
  assign n96305 = ~n95855 & n96304;
  assign n96306 = n96302 & n96305;
  assign n96307 = ~n95813 & ~n96306;
  assign n96308 = ~n96292 & ~n96307;
  assign n96309 = ~n96284 & n96308;
  assign n96310 = n96282 & n96309;
  assign n96311 = pi5352 & ~n96310;
  assign n96312 = ~pi5352 & n96310;
  assign po3560 = n96311 | n96312;
  assign n96314 = ~n95490 & n95538;
  assign n96315 = n95490 & n95547;
  assign n96316 = ~n96314 & ~n96315;
  assign n96317 = n95471 & ~n96316;
  assign n96318 = ~n95490 & n95527;
  assign n96319 = n95490 & n95522;
  assign n96320 = ~n96318 & ~n96319;
  assign n96321 = ~n95471 & ~n96320;
  assign n96322 = ~n95484 & ~n95547;
  assign n96323 = ~n95490 & ~n96322;
  assign n96324 = ~n95522 & ~n96323;
  assign n96325 = ~n95471 & ~n96324;
  assign n96326 = ~n95483 & n95490;
  assign n96327 = ~n95471 & ~n95496;
  assign n96328 = n96326 & n96327;
  assign n96329 = n95483 & n95496;
  assign n96330 = ~n95522 & ~n96329;
  assign n96331 = n95490 & ~n96330;
  assign n96332 = n95471 & ~n95490;
  assign n96333 = n95512 & n96332;
  assign n96334 = ~n95496 & n96333;
  assign n96335 = ~n96331 & ~n96334;
  assign n96336 = ~n96328 & n96335;
  assign n96337 = ~n96325 & n96336;
  assign n96338 = ~n96318 & n96337;
  assign n96339 = ~n95508 & ~n96338;
  assign n96340 = ~n95471 & ~n95490;
  assign n96341 = ~n95515 & ~n95530;
  assign n96342 = n96340 & ~n96341;
  assign n96343 = n95515 & n96327;
  assign n96344 = ~n96342 & ~n96343;
  assign n96345 = n95508 & ~n96344;
  assign n96346 = n95490 & n95513;
  assign n96347 = n95490 & n95496;
  assign n96348 = ~n95547 & ~n96347;
  assign n96349 = n95471 & ~n96348;
  assign n96350 = n95490 & ~n95496;
  assign n96351 = n95483 & n96350;
  assign n96352 = n95477 & n96351;
  assign n96353 = ~n96349 & ~n96352;
  assign n96354 = ~n96346 & n96353;
  assign n96355 = n95508 & ~n96354;
  assign n96356 = ~n96345 & ~n96355;
  assign n96357 = ~n96339 & n96356;
  assign n96358 = ~n96321 & n96357;
  assign n96359 = ~n96317 & n96358;
  assign n96360 = pi5432 & n96359;
  assign n96361 = ~pi5432 & ~n96359;
  assign po3562 = n96360 | n96361;
  assign n96363 = n95980 & n96044;
  assign n96364 = n95986 & n96017;
  assign n96365 = n95974 & n96364;
  assign n96366 = n95974 & n96027;
  assign n96367 = ~n96365 & ~n96366;
  assign n96368 = ~n95992 & n96015;
  assign n96369 = ~n95980 & n96368;
  assign n96370 = ~n96009 & ~n96369;
  assign n96371 = ~n96006 & ~n96370;
  assign n96372 = n96367 & ~n96371;
  assign n96373 = ~n96363 & n96372;
  assign n96374 = n95968 & ~n96373;
  assign n96375 = n95974 & n96049;
  assign n96376 = n96006 & n96375;
  assign n96377 = n96039 & n96049;
  assign n96378 = ~n96007 & ~n96377;
  assign n96379 = ~n96009 & ~n96041;
  assign n96380 = ~n95974 & n96026;
  assign n96381 = n96379 & ~n96380;
  assign n96382 = n96006 & ~n96381;
  assign n96383 = ~n96006 & n96013;
  assign n96384 = n96031 & ~n96383;
  assign n96385 = ~n96382 & n96384;
  assign n96386 = n96378 & n96385;
  assign n96387 = ~n95968 & ~n96386;
  assign n96388 = ~n96376 & ~n96387;
  assign n96389 = ~n96374 & n96388;
  assign n96390 = n96039 & n96041;
  assign n96391 = n95993 & ~n96006;
  assign n96392 = n95974 & n96391;
  assign n96393 = ~n96390 & ~n96392;
  assign n96394 = ~n96006 & n96366;
  assign n96395 = n96393 & ~n96394;
  assign n96396 = n96389 & n96395;
  assign n96397 = ~pi5301 & ~n96396;
  assign n96398 = pi5301 & n96395;
  assign n96399 = n96388 & n96398;
  assign n96400 = ~n96374 & n96399;
  assign po3576 = n96397 | n96400;
  assign n96402 = n95587 & n95627;
  assign n96403 = n95621 & ~n96246;
  assign n96404 = ~n95647 & ~n96403;
  assign n96405 = ~n96075 & n96404;
  assign n96406 = ~n95587 & ~n96405;
  assign n96407 = ~n95581 & n95597;
  assign n96408 = ~n96406 & ~n96407;
  assign n96409 = ~n95595 & n95646;
  assign n96410 = n95581 & n96080;
  assign n96411 = ~n96409 & ~n96410;
  assign n96412 = ~n96249 & n96411;
  assign n96413 = n95587 & ~n96412;
  assign n96414 = n96408 & ~n96413;
  assign n96415 = n95562 & ~n96414;
  assign n96416 = ~n96402 & ~n96415;
  assign n96417 = n95581 & n95596;
  assign n96418 = ~n96074 & ~n96417;
  assign n96419 = n95587 & ~n96418;
  assign n96420 = ~n95648 & ~n96419;
  assign n96421 = ~n95615 & ~n95627;
  assign n96422 = ~n95581 & n95653;
  assign n96423 = ~n96080 & ~n96422;
  assign n96424 = ~n96409 & n96423;
  assign n96425 = ~n95587 & ~n96424;
  assign n96426 = n95581 & n95597;
  assign n96427 = ~n96425 & ~n96426;
  assign n96428 = n96421 & n96427;
  assign n96429 = n96420 & n96428;
  assign n96430 = ~n95562 & ~n96429;
  assign n96431 = ~n95634 & ~n96245;
  assign n96432 = ~n95587 & ~n96431;
  assign n96433 = ~n96430 & ~n96432;
  assign n96434 = n96416 & n96433;
  assign n96435 = pi5356 & n96434;
  assign n96436 = ~pi5356 & ~n96434;
  assign po3577 = n96435 | n96436;
  assign n96438 = ~n95667 & n95701;
  assign n96439 = ~n96209 & ~n96438;
  assign n96440 = n95694 & ~n96439;
  assign n96441 = n95720 & n95752;
  assign n96442 = ~n96440 & ~n96441;
  assign n96443 = ~n95763 & n96442;
  assign n96444 = n95667 & n95687;
  assign n96445 = ~n95701 & ~n96444;
  assign n96446 = ~n96218 & n96445;
  assign n96447 = n95694 & ~n96446;
  assign n96448 = n95718 & n96447;
  assign n96449 = ~n95679 & ~n95694;
  assign n96450 = n95685 & n96449;
  assign n96451 = ~n95673 & n96450;
  assign n96452 = ~n95667 & n96451;
  assign n96453 = n95667 & n95704;
  assign n96454 = ~n96208 & ~n96453;
  assign n96455 = ~n96451 & n96454;
  assign n96456 = ~n95667 & n95679;
  assign n96457 = n95685 & n96456;
  assign n96458 = n95667 & n95736;
  assign n96459 = ~n95695 & ~n96458;
  assign n96460 = n95694 & ~n96459;
  assign n96461 = ~n96457 & ~n96460;
  assign n96462 = n96455 & n96461;
  assign n96463 = ~n95718 & ~n96462;
  assign n96464 = ~n95694 & n96220;
  assign n96465 = ~n95732 & ~n95749;
  assign n96466 = ~n95744 & n96465;
  assign n96467 = ~n96464 & n96466;
  assign n96468 = n95718 & ~n96467;
  assign n96469 = ~n96463 & ~n96468;
  assign n96470 = ~n96452 & n96469;
  assign n96471 = ~n96448 & n96470;
  assign n96472 = n96443 & n96471;
  assign n96473 = pi5689 & ~n96472;
  assign n96474 = ~pi5689 & n96443;
  assign n96475 = n96471 & n96474;
  assign po3578 = n96473 | n96475;
  assign n96477 = ~n95490 & n95521;
  assign n96478 = n95483 & n95490;
  assign n96479 = ~n95496 & n96478;
  assign n96480 = ~n96477 & ~n96479;
  assign n96481 = n95471 & ~n96480;
  assign n96482 = n95483 & n95499;
  assign n96483 = ~n95530 & ~n96482;
  assign n96484 = ~n95471 & ~n96483;
  assign n96485 = n95490 & n95516;
  assign n96486 = ~n96328 & ~n96485;
  assign n96487 = ~n96484 & n96486;
  assign n96488 = ~n96481 & n96487;
  assign n96489 = ~n95498 & n96488;
  assign n96490 = ~n96318 & ~n96346;
  assign n96491 = n96489 & n96490;
  assign n96492 = n95508 & ~n96491;
  assign n96493 = n95484 & n96347;
  assign n96494 = n95539 & ~n96493;
  assign n96495 = n95471 & ~n96494;
  assign n96496 = n95490 & n95527;
  assign n96497 = ~n96495 & ~n96496;
  assign n96498 = n95477 & n95499;
  assign n96499 = ~n95490 & n95512;
  assign n96500 = ~n96498 & ~n96499;
  assign n96501 = n95471 & ~n96500;
  assign n96502 = n95471 & n95521;
  assign n96503 = n95490 & n96502;
  assign n96504 = ~n96501 & ~n96503;
  assign n96505 = n96497 & n96504;
  assign n96506 = ~n95508 & ~n96505;
  assign n96507 = ~n95516 & ~n96352;
  assign n96508 = ~n95523 & n96507;
  assign n96509 = n95544 & ~n96508;
  assign n96510 = ~n96506 & ~n96509;
  assign n96511 = ~n95498 & ~n96346;
  assign n96512 = ~n95471 & ~n96511;
  assign n96513 = n96510 & ~n96512;
  assign n96514 = ~n96492 & n96513;
  assign n96515 = ~pi5551 & n96514;
  assign n96516 = pi5551 & ~n96514;
  assign po3581 = n96515 | n96516;
  assign n96518 = ~n95974 & n96364;
  assign n96519 = ~n96027 & ~n96035;
  assign n96520 = n95974 & n95993;
  assign n96521 = ~n95974 & n96049;
  assign n96522 = ~n96520 & ~n96521;
  assign n96523 = n96519 & n96522;
  assign n96524 = n96006 & ~n96523;
  assign n96525 = n95974 & n96008;
  assign n96526 = ~n96007 & ~n96525;
  assign n96527 = ~n96029 & n96526;
  assign n96528 = ~n96006 & ~n96527;
  assign n96529 = n95974 & ~n95986;
  assign n96530 = ~n95998 & n96529;
  assign n96531 = n95980 & n96530;
  assign n96532 = ~n96528 & ~n96531;
  assign n96533 = ~n96524 & n96532;
  assign n96534 = ~n96518 & n96533;
  assign n96535 = ~n95968 & ~n96534;
  assign n96536 = n95974 & n96006;
  assign n96537 = n96013 & n96536;
  assign n96538 = n96006 & n96029;
  assign n96539 = n96006 & n96041;
  assign n96540 = ~n96538 & ~n96539;
  assign n96541 = ~n95974 & ~n96540;
  assign n96542 = ~n96537 & ~n96541;
  assign n96543 = ~n95974 & n95994;
  assign n96544 = ~n96375 & ~n96543;
  assign n96545 = n95974 & n96026;
  assign n96546 = ~n95974 & n96008;
  assign n96547 = ~n96545 & ~n96546;
  assign n96548 = ~n95994 & n96547;
  assign n96549 = ~n96027 & n96548;
  assign n96550 = ~n96006 & ~n96549;
  assign n96551 = ~n95974 & n96009;
  assign n96552 = ~n96550 & ~n96551;
  assign n96553 = n96544 & n96552;
  assign n96554 = n96542 & n96553;
  assign n96555 = n95968 & ~n96554;
  assign n96556 = n96006 & ~n96367;
  assign n96557 = ~n96555 & ~n96556;
  assign n96558 = ~n96030 & ~n96543;
  assign n96559 = ~n96006 & ~n96558;
  assign n96560 = n96557 & ~n96559;
  assign n96561 = ~n96535 & n96560;
  assign n96562 = pi5300 & ~n96561;
  assign n96563 = ~pi5300 & n96561;
  assign po3583 = n96562 | n96563;
  assign n96565 = ~n95687 & ~n95701;
  assign n96566 = ~n95752 & ~n96218;
  assign n96567 = n96565 & n96566;
  assign n96568 = n95667 & ~n96567;
  assign n96569 = ~n95686 & ~n96220;
  assign n96570 = n95737 & ~n96569;
  assign n96571 = ~n96568 & ~n96570;
  assign n96572 = ~n96209 & n96571;
  assign n96573 = n95718 & ~n96572;
  assign n96574 = n95667 & n96232;
  assign n96575 = n95685 & n96207;
  assign n96576 = ~n95708 & ~n96575;
  assign n96577 = ~n96218 & n96576;
  assign n96578 = ~n95694 & ~n96577;
  assign n96579 = n95694 & ~n96569;
  assign n96580 = ~n96578 & ~n96579;
  assign n96581 = ~n96574 & n96580;
  assign n96582 = ~n95667 & n95752;
  assign n96583 = n96581 & ~n96582;
  assign n96584 = ~n95718 & ~n96583;
  assign n96585 = n95667 & n96220;
  assign n96586 = ~n96582 & ~n96585;
  assign n96587 = n95694 & ~n96586;
  assign n96588 = ~n96584 & ~n96587;
  assign n96589 = ~n96573 & n96588;
  assign n96590 = ~pi5647 & ~n96589;
  assign n96591 = pi5647 & ~n96587;
  assign n96592 = ~n96573 & n96591;
  assign n96593 = ~n96584 & n96592;
  assign po3586 = n96590 | n96593;
  assign n96595 = ~n95395 & n95424;
  assign n96596 = n95395 & n95435;
  assign n96597 = ~n95421 & ~n96596;
  assign n96598 = n95369 & ~n96597;
  assign n96599 = ~n96595 & ~n96598;
  assign n96600 = n95387 & n95457;
  assign n96601 = ~n95381 & n96600;
  assign n96602 = n95403 & n95436;
  assign n96603 = ~n96601 & ~n96602;
  assign n96604 = ~n95369 & n95445;
  assign n96605 = n96603 & ~n96604;
  assign n96606 = ~n95399 & ~n95411;
  assign n96607 = ~n95450 & n96606;
  assign n96608 = n96605 & n96607;
  assign n96609 = n96599 & n96608;
  assign n96610 = ~n95433 & ~n96609;
  assign n96611 = ~n95398 & ~n95421;
  assign n96612 = n95395 & ~n96611;
  assign n96613 = ~n95381 & n95439;
  assign n96614 = ~n95375 & n95403;
  assign n96615 = ~n96613 & ~n96614;
  assign n96616 = ~n95375 & n95387;
  assign n96617 = n95395 & n96616;
  assign n96618 = n96615 & ~n96617;
  assign n96619 = n95369 & ~n96618;
  assign n96620 = ~n95395 & n95409;
  assign n96621 = n95389 & n95395;
  assign n96622 = ~n96620 & ~n96621;
  assign n96623 = ~n95369 & ~n96622;
  assign n96624 = ~n95395 & n95404;
  assign n96625 = ~n96623 & ~n96624;
  assign n96626 = ~n96619 & n96625;
  assign n96627 = ~n96612 & n96626;
  assign n96628 = n95433 & ~n96627;
  assign n96629 = n95369 & n95440;
  assign n96630 = ~n96628 & ~n96629;
  assign n96631 = n95416 & n95457;
  assign n96632 = n95387 & n96631;
  assign n96633 = n96630 & ~n96632;
  assign n96634 = ~n96610 & n96633;
  assign n96635 = ~pi5467 & ~n96634;
  assign n96636 = pi5467 & n96630;
  assign n96637 = ~n96610 & n96636;
  assign n96638 = ~n96632 & n96637;
  assign po3587 = n96635 | n96638;
  assign n96640 = ~n95396 & ~n95402;
  assign n96641 = ~n95369 & ~n96640;
  assign n96642 = ~n95459 & ~n96641;
  assign n96643 = n95375 & n95381;
  assign n96644 = n95369 & n96643;
  assign n96645 = n95395 & n96644;
  assign n96646 = n95395 & n95409;
  assign n96647 = ~n96643 & ~n96646;
  assign n96648 = ~n95375 & ~n95395;
  assign n96649 = ~n95381 & n96648;
  assign n96650 = n96647 & ~n96649;
  assign n96651 = n95369 & ~n96650;
  assign n96652 = ~n95405 & ~n96651;
  assign n96653 = ~n95433 & ~n96652;
  assign n96654 = ~n95369 & n95388;
  assign n96655 = n95395 & n96654;
  assign n96656 = ~n96604 & ~n96655;
  assign n96657 = ~n95433 & ~n96656;
  assign n96658 = ~n96653 & ~n96657;
  assign n96659 = ~n96645 & n96658;
  assign n96660 = ~n95421 & ~n95440;
  assign n96661 = ~n96614 & n96660;
  assign n96662 = ~n95369 & ~n96661;
  assign n96663 = ~n95387 & n96648;
  assign n96664 = n95381 & n96663;
  assign n96665 = ~n95424 & ~n96664;
  assign n96666 = n95369 & ~n96665;
  assign n96667 = ~n96613 & ~n96666;
  assign n96668 = ~n96662 & n96667;
  assign n96669 = ~n95411 & ~n95451;
  assign n96670 = n96668 & n96669;
  assign n96671 = n95433 & ~n96670;
  assign n96672 = n96659 & ~n96671;
  assign n96673 = n96642 & n96672;
  assign n96674 = ~pi5497 & ~n96673;
  assign n96675 = pi5497 & n96659;
  assign n96676 = n96642 & n96675;
  assign n96677 = ~n96671 & n96676;
  assign po3588 = n96674 | n96677;
  assign n96679 = pi7466 & ~pi9040;
  assign n96680 = pi7430 & pi9040;
  assign n96681 = ~n96679 & ~n96680;
  assign n96682 = ~pi3943 & ~n96681;
  assign n96683 = pi3943 & n96681;
  assign n96684 = ~n96682 & ~n96683;
  assign n96685 = pi7379 & pi9040;
  assign n96686 = pi7428 & ~pi9040;
  assign n96687 = ~n96685 & ~n96686;
  assign n96688 = ~pi3852 & n96687;
  assign n96689 = pi3852 & ~n96687;
  assign n96690 = ~n96688 & ~n96689;
  assign n96691 = pi7428 & pi9040;
  assign n96692 = pi7401 & ~pi9040;
  assign n96693 = ~n96691 & ~n96692;
  assign n96694 = ~pi3930 & n96693;
  assign n96695 = pi3930 & ~n96693;
  assign n96696 = ~n96694 & ~n96695;
  assign n96697 = n96690 & ~n96696;
  assign n96698 = n96684 & n96697;
  assign n96699 = pi7528 & pi9040;
  assign n96700 = pi7460 & ~pi9040;
  assign n96701 = ~n96699 & ~n96700;
  assign n96702 = ~pi3940 & n96701;
  assign n96703 = pi3940 & ~n96701;
  assign n96704 = ~n96702 & ~n96703;
  assign n96705 = n96684 & ~n96704;
  assign n96706 = ~n96696 & n96705;
  assign n96707 = ~n96684 & ~n96704;
  assign n96708 = n96696 & n96707;
  assign n96709 = ~n96706 & ~n96708;
  assign n96710 = ~n96698 & n96709;
  assign n96711 = pi7366 & pi9040;
  assign n96712 = pi7436 & ~pi9040;
  assign n96713 = ~n96711 & ~n96712;
  assign n96714 = pi3846 & n96713;
  assign n96715 = ~pi3846 & ~n96713;
  assign n96716 = ~n96714 & ~n96715;
  assign n96717 = pi7396 & ~pi9040;
  assign n96718 = pi7401 & pi9040;
  assign n96719 = ~n96717 & ~n96718;
  assign n96720 = ~pi3840 & ~n96719;
  assign n96721 = pi3840 & n96719;
  assign n96722 = ~n96720 & ~n96721;
  assign n96723 = ~n96716 & n96722;
  assign n96724 = ~n96710 & n96723;
  assign n96725 = ~n96684 & n96704;
  assign n96726 = ~n96696 & n96725;
  assign n96727 = ~n96690 & n96722;
  assign n96728 = n96726 & n96727;
  assign n96729 = ~n96696 & n96707;
  assign n96730 = n96716 & n96729;
  assign n96731 = n96684 & n96704;
  assign n96732 = ~n96690 & n96731;
  assign n96733 = n96684 & n96696;
  assign n96734 = ~n96732 & ~n96733;
  assign n96735 = n96716 & ~n96734;
  assign n96736 = ~n96730 & ~n96735;
  assign n96737 = n96722 & ~n96736;
  assign n96738 = ~n96728 & ~n96737;
  assign n96739 = ~n96690 & n96696;
  assign n96740 = n96684 & n96739;
  assign n96741 = n96690 & n96696;
  assign n96742 = ~n96684 & n96741;
  assign n96743 = n96704 & n96742;
  assign n96744 = ~n96740 & ~n96743;
  assign n96745 = n96716 & ~n96744;
  assign n96746 = n96738 & ~n96745;
  assign n96747 = ~n96690 & ~n96716;
  assign n96748 = n96731 & n96747;
  assign n96749 = ~n96696 & n96748;
  assign n96750 = ~n96705 & ~n96725;
  assign n96751 = n96697 & ~n96750;
  assign n96752 = ~n96704 & n96742;
  assign n96753 = ~n96751 & ~n96752;
  assign n96754 = n96696 & n96731;
  assign n96755 = n96690 & ~n96716;
  assign n96756 = n96754 & n96755;
  assign n96757 = n96739 & ~n96750;
  assign n96758 = ~n96690 & ~n96696;
  assign n96759 = ~n96684 & n96758;
  assign n96760 = ~n96704 & n96759;
  assign n96761 = ~n96757 & ~n96760;
  assign n96762 = ~n96756 & n96761;
  assign n96763 = n96753 & n96762;
  assign n96764 = ~n96749 & n96763;
  assign n96765 = n96690 & n96716;
  assign n96766 = ~n96696 & n96765;
  assign n96767 = n96704 & n96766;
  assign n96768 = n96764 & ~n96767;
  assign n96769 = ~n96722 & ~n96768;
  assign n96770 = n96746 & ~n96769;
  assign n96771 = ~n96724 & n96770;
  assign n96772 = ~pi5433 & ~n96771;
  assign n96773 = pi5433 & n96746;
  assign n96774 = ~n96724 & n96773;
  assign n96775 = ~n96769 & n96774;
  assign po3589 = n96772 | n96775;
  assign n96777 = n95490 & n95512;
  assign n96778 = ~n95511 & ~n96777;
  assign n96779 = ~n95471 & ~n96778;
  assign n96780 = n95471 & ~n96330;
  assign n96781 = ~n96314 & ~n96780;
  assign n96782 = ~n96779 & n96781;
  assign n96783 = n95508 & ~n96782;
  assign n96784 = ~n95471 & n95527;
  assign n96785 = ~n96783 & ~n96784;
  assign n96786 = ~n96485 & ~n96499;
  assign n96787 = n95471 & ~n96786;
  assign n96788 = n95496 & n96340;
  assign n96789 = ~n96350 & ~n96788;
  assign n96790 = ~n95477 & ~n96789;
  assign n96791 = ~n96479 & ~n96790;
  assign n96792 = ~n95498 & n96791;
  assign n96793 = n95471 & n95513;
  assign n96794 = ~n95490 & n95530;
  assign n96795 = ~n96793 & ~n96794;
  assign n96796 = n96792 & n96795;
  assign n96797 = ~n95508 & ~n96796;
  assign n96798 = ~n96787 & ~n96797;
  assign n96799 = n96785 & n96798;
  assign n96800 = pi5603 & ~n96799;
  assign n96801 = ~pi5603 & n96799;
  assign po3590 = n96800 | n96801;
  assign n96803 = ~n95451 & ~n96624;
  assign n96804 = n95369 & ~n96803;
  assign n96805 = ~n95433 & n95435;
  assign n96806 = ~n95369 & n96805;
  assign n96807 = n95381 & n96648;
  assign n96808 = ~n96616 & ~n96807;
  assign n96809 = ~n95404 & n96808;
  assign n96810 = n95369 & ~n96809;
  assign n96811 = ~n95395 & n95410;
  assign n96812 = ~n96810 & ~n96811;
  assign n96813 = ~n95433 & ~n96812;
  assign n96814 = ~n96806 & ~n96813;
  assign n96815 = ~n95399 & ~n95402;
  assign n96816 = ~n95395 & n96614;
  assign n96817 = ~n96596 & ~n96816;
  assign n96818 = n96815 & n96817;
  assign n96819 = ~n95369 & ~n96818;
  assign n96820 = n95375 & n95436;
  assign n96821 = ~n95381 & n96820;
  assign n96822 = ~n95395 & n96616;
  assign n96823 = ~n95402 & ~n96822;
  assign n96824 = ~n96621 & n96823;
  assign n96825 = ~n96821 & n96824;
  assign n96826 = n95369 & n95398;
  assign n96827 = n96825 & ~n96826;
  assign n96828 = n95433 & ~n96827;
  assign n96829 = ~n96819 & ~n96828;
  assign n96830 = n96814 & n96829;
  assign n96831 = ~n96804 & n96830;
  assign n96832 = pi5691 & n96831;
  assign n96833 = ~pi5691 & ~n96831;
  assign po3617 = n96832 | n96833;
  assign n96835 = ~n96690 & n96725;
  assign n96836 = n96690 & n96731;
  assign n96837 = ~n96835 & ~n96836;
  assign n96838 = n96716 & ~n96837;
  assign n96839 = n96716 & n96752;
  assign n96840 = ~n96838 & ~n96839;
  assign n96841 = n96722 & ~n96840;
  assign n96842 = n96741 & ~n96750;
  assign n96843 = ~n96696 & n96731;
  assign n96844 = n96696 & ~n96704;
  assign n96845 = ~n96705 & ~n96844;
  assign n96846 = n96690 & ~n96845;
  assign n96847 = ~n96843 & ~n96846;
  assign n96848 = ~n96716 & ~n96847;
  assign n96849 = ~n96842 & ~n96848;
  assign n96850 = ~n96690 & n96754;
  assign n96851 = ~n96684 & n96697;
  assign n96852 = ~n96690 & ~n96845;
  assign n96853 = ~n96851 & ~n96852;
  assign n96854 = n96716 & ~n96853;
  assign n96855 = ~n96850 & ~n96854;
  assign n96856 = n96849 & n96855;
  assign n96857 = ~n96722 & ~n96856;
  assign n96858 = ~n96696 & n96722;
  assign n96859 = ~n96705 & n96858;
  assign n96860 = ~n96690 & n96859;
  assign n96861 = n96705 & n96739;
  assign n96862 = n96716 & n96861;
  assign n96863 = ~n96696 & n96747;
  assign n96864 = ~n96684 & n96863;
  assign n96865 = ~n96862 & ~n96864;
  assign n96866 = ~n96860 & n96865;
  assign n96867 = ~n96690 & ~n96704;
  assign n96868 = ~n96726 & ~n96867;
  assign n96869 = n96723 & ~n96868;
  assign n96870 = n96866 & ~n96869;
  assign n96871 = ~n96857 & n96870;
  assign n96872 = ~n96841 & n96871;
  assign n96873 = pi5646 & ~n96872;
  assign n96874 = ~pi5646 & n96872;
  assign po3633 = n96873 | n96874;
  assign n96876 = n96716 & n96843;
  assign n96877 = n96690 & n96876;
  assign n96878 = ~n96839 & ~n96877;
  assign n96879 = ~n96752 & ~n96756;
  assign n96880 = ~n96716 & ~n96741;
  assign n96881 = ~n96750 & n96880;
  assign n96882 = ~n96731 & n96765;
  assign n96883 = n96696 & n96882;
  assign n96884 = ~n96696 & ~n96704;
  assign n96885 = ~n96690 & n96884;
  assign n96886 = ~n96732 & ~n96885;
  assign n96887 = n96716 & ~n96886;
  assign n96888 = ~n96883 & ~n96887;
  assign n96889 = ~n96881 & n96888;
  assign n96890 = n96879 & n96889;
  assign n96891 = n96722 & ~n96890;
  assign n96892 = n96878 & ~n96891;
  assign n96893 = n96706 & ~n96716;
  assign n96894 = ~n96690 & n96893;
  assign n96895 = ~n96716 & ~n96722;
  assign n96896 = ~n96729 & ~n96732;
  assign n96897 = ~n96842 & n96896;
  assign n96898 = n96895 & ~n96897;
  assign n96899 = ~n96690 & n96708;
  assign n96900 = n96696 & n96867;
  assign n96901 = ~n96835 & ~n96900;
  assign n96902 = ~n96726 & ~n96836;
  assign n96903 = n96901 & n96902;
  assign n96904 = n96716 & ~n96903;
  assign n96905 = ~n96899 & ~n96904;
  assign n96906 = ~n96722 & ~n96905;
  assign n96907 = ~n96898 & ~n96906;
  assign n96908 = ~n96894 & n96907;
  assign n96909 = n96892 & n96908;
  assign n96910 = pi5599 & ~n96909;
  assign n96911 = ~pi5599 & n96892;
  assign n96912 = n96908 & n96911;
  assign po3634 = n96910 | n96912;
  assign n96914 = ~n96369 & ~n96543;
  assign n96915 = ~n96531 & n96914;
  assign n96916 = n96006 & ~n96915;
  assign n96917 = ~n96377 & ~n96394;
  assign n96918 = ~n96375 & ~n96539;
  assign n96919 = ~n96364 & ~n96546;
  assign n96920 = ~n96006 & ~n96919;
  assign n96921 = ~n96035 & ~n96920;
  assign n96922 = n96918 & n96921;
  assign n96923 = n95968 & ~n96922;
  assign n96924 = ~n95986 & ~n95998;
  assign n96925 = ~n96014 & ~n96924;
  assign n96926 = n95974 & ~n96925;
  assign n96927 = ~n95994 & ~n96380;
  assign n96928 = ~n96006 & ~n96927;
  assign n96929 = n95974 & n95992;
  assign n96930 = ~n96009 & ~n96929;
  assign n96931 = ~n96017 & n96930;
  assign n96932 = n96006 & ~n96931;
  assign n96933 = ~n96928 & ~n96932;
  assign n96934 = ~n96926 & n96933;
  assign n96935 = ~n95968 & ~n96934;
  assign n96936 = ~n96923 & ~n96935;
  assign n96937 = n96917 & n96936;
  assign n96938 = ~n96916 & n96937;
  assign n96939 = ~pi5531 & ~n96938;
  assign n96940 = pi5531 & n96917;
  assign n96941 = ~n96916 & n96940;
  assign n96942 = n96936 & n96941;
  assign po3635 = n96939 | n96942;
  assign n96944 = n96696 & n96835;
  assign n96945 = ~n96760 & ~n96944;
  assign n96946 = n96716 & ~n96945;
  assign n96947 = n96696 & n96705;
  assign n96948 = ~n96843 & ~n96947;
  assign n96949 = n96716 & ~n96948;
  assign n96950 = n96690 & n96725;
  assign n96951 = ~n96706 & ~n96950;
  assign n96952 = ~n96754 & n96951;
  assign n96953 = ~n96716 & ~n96952;
  assign n96954 = ~n96949 & ~n96953;
  assign n96955 = ~n96730 & ~n96743;
  assign n96956 = n96954 & n96955;
  assign n96957 = ~n96722 & ~n96956;
  assign n96958 = ~n96690 & n96843;
  assign n96959 = n96690 & n96707;
  assign n96960 = ~n96835 & ~n96959;
  assign n96961 = ~n96716 & ~n96960;
  assign n96962 = ~n96958 & ~n96961;
  assign n96963 = n96716 & n96726;
  assign n96964 = n96709 & ~n96963;
  assign n96965 = ~n96754 & n96964;
  assign n96966 = n96690 & ~n96965;
  assign n96967 = n96962 & ~n96966;
  assign n96968 = n96722 & ~n96967;
  assign n96969 = ~n96957 & ~n96968;
  assign n96970 = ~n96716 & n96844;
  assign n96971 = ~n96690 & n96970;
  assign n96972 = n96969 & ~n96971;
  assign n96973 = ~n96946 & n96972;
  assign n96974 = ~pi5523 & ~n96973;
  assign n96975 = pi5523 & ~n96946;
  assign n96976 = n96969 & n96975;
  assign n96977 = ~n96971 & n96976;
  assign po3652 = n96974 | n96977;
  assign n96979 = pi7659 & pi9040;
  assign n96980 = pi7666 & ~pi9040;
  assign n96981 = ~n96979 & ~n96980;
  assign n96982 = ~pi5607 & ~n96981;
  assign n96983 = pi5607 & n96981;
  assign n96984 = ~n96982 & ~n96983;
  assign n96985 = pi7675 & ~pi9040;
  assign n96986 = pi7648 & pi9040;
  assign n96987 = ~n96985 & ~n96986;
  assign n96988 = ~pi5658 & n96987;
  assign n96989 = pi5658 & ~n96987;
  assign n96990 = ~n96988 & ~n96989;
  assign n96991 = pi7749 & ~pi9040;
  assign n96992 = pi7739 & pi9040;
  assign n96993 = ~n96991 & ~n96992;
  assign n96994 = pi5684 & n96993;
  assign n96995 = ~pi5684 & ~n96993;
  assign n96996 = ~n96994 & ~n96995;
  assign n96997 = pi7662 & ~pi9040;
  assign n96998 = pi7725 & pi9040;
  assign n96999 = ~n96997 & ~n96998;
  assign n97000 = ~pi5856 & n96999;
  assign n97001 = pi5856 & ~n96999;
  assign n97002 = ~n97000 & ~n97001;
  assign n97003 = pi7720 & pi9040;
  assign n97004 = pi7739 & ~pi9040;
  assign n97005 = ~n97003 & ~n97004;
  assign n97006 = ~pi5431 & ~n97005;
  assign n97007 = pi5431 & n97005;
  assign n97008 = ~n97006 & ~n97007;
  assign n97009 = n97002 & n97008;
  assign n97010 = n96996 & n97009;
  assign n97011 = n96990 & n97010;
  assign n97012 = pi7653 & ~pi9040;
  assign n97013 = pi7745 & pi9040;
  assign n97014 = ~n97012 & ~n97013;
  assign n97015 = pi5512 & n97014;
  assign n97016 = ~pi5512 & ~n97014;
  assign n97017 = ~n97015 & ~n97016;
  assign n97018 = ~n97002 & ~n97008;
  assign n97019 = n97017 & n97018;
  assign n97020 = ~n96990 & ~n97017;
  assign n97021 = ~n97008 & n97020;
  assign n97022 = n97002 & n97021;
  assign n97023 = ~n97019 & ~n97022;
  assign n97024 = ~n97002 & n97008;
  assign n97025 = ~n96990 & n97024;
  assign n97026 = n97023 & ~n97025;
  assign n97027 = n96996 & ~n97026;
  assign n97028 = ~n97002 & ~n97017;
  assign n97029 = n96990 & ~n96996;
  assign n97030 = n97028 & n97029;
  assign n97031 = n96990 & ~n97017;
  assign n97032 = ~n97008 & n97031;
  assign n97033 = ~n97002 & n97032;
  assign n97034 = ~n97030 & ~n97033;
  assign n97035 = ~n97027 & n97034;
  assign n97036 = ~n97011 & n97035;
  assign n97037 = n97009 & n97017;
  assign n97038 = n96990 & n97037;
  assign n97039 = n97017 & n97024;
  assign n97040 = ~n96990 & n97039;
  assign n97041 = ~n97038 & ~n97040;
  assign n97042 = n97036 & n97041;
  assign n97043 = ~n96984 & ~n97042;
  assign n97044 = ~n97017 & n97024;
  assign n97045 = n96990 & n97044;
  assign n97046 = ~n97037 & ~n97045;
  assign n97047 = n96996 & ~n97046;
  assign n97048 = n97009 & ~n97017;
  assign n97049 = ~n96990 & n97048;
  assign n97050 = n97002 & ~n97008;
  assign n97051 = n97031 & n97050;
  assign n97052 = ~n97049 & ~n97051;
  assign n97053 = ~n97002 & n97020;
  assign n97054 = n96990 & n97039;
  assign n97055 = ~n97053 & ~n97054;
  assign n97056 = ~n96996 & ~n97055;
  assign n97057 = n97052 & ~n97056;
  assign n97058 = ~n97047 & n97057;
  assign n97059 = n96984 & ~n97058;
  assign n97060 = ~n97002 & n97017;
  assign n97061 = ~n96990 & n97060;
  assign n97062 = n97002 & n97017;
  assign n97063 = n96990 & n97062;
  assign n97064 = ~n97061 & ~n97063;
  assign n97065 = n96996 & ~n97064;
  assign n97066 = n97017 & n97050;
  assign n97067 = ~n96990 & n97066;
  assign n97068 = ~n97049 & ~n97067;
  assign n97069 = ~n97017 & n97018;
  assign n97070 = n97068 & ~n97069;
  assign n97071 = ~n96996 & ~n97070;
  assign n97072 = ~n97065 & ~n97071;
  assign n97073 = ~n97008 & ~n97017;
  assign n97074 = ~n96996 & n97073;
  assign n97075 = n96990 & n97074;
  assign n97076 = n97072 & ~n97075;
  assign n97077 = ~n97059 & n97076;
  assign n97078 = ~n97043 & n97077;
  assign n97079 = ~pi8568 & ~n97078;
  assign n97080 = pi8568 & n97078;
  assign po4012 = n97079 | n97080;
  assign n97082 = pi7742 & pi9040;
  assign n97083 = pi7741 & ~pi9040;
  assign n97084 = ~n97082 & ~n97083;
  assign n97085 = ~pi5694 & n97084;
  assign n97086 = pi5694 & ~n97084;
  assign n97087 = ~n97085 & ~n97086;
  assign n97088 = pi7811 & ~pi9040;
  assign n97089 = pi7689 & pi9040;
  assign n97090 = ~n97088 & ~n97089;
  assign n97091 = ~pi5693 & n97090;
  assign n97092 = pi5693 & ~n97090;
  assign n97093 = ~n97091 & ~n97092;
  assign n97094 = pi7742 & ~pi9040;
  assign n97095 = pi7811 & pi9040;
  assign n97096 = ~n97094 & ~n97095;
  assign n97097 = ~pi5703 & n97096;
  assign n97098 = pi5703 & ~n97096;
  assign n97099 = ~n97097 & ~n97098;
  assign n97100 = ~n97093 & n97099;
  assign n97101 = n97087 & n97100;
  assign n97102 = pi7661 & pi9040;
  assign n97103 = pi7817 & ~pi9040;
  assign n97104 = ~n97102 & ~n97103;
  assign n97105 = ~pi5841 & n97104;
  assign n97106 = pi5841 & ~n97104;
  assign n97107 = ~n97105 & ~n97106;
  assign n97108 = ~n97087 & ~n97099;
  assign n97109 = n97107 & n97108;
  assign n97110 = ~n97101 & ~n97109;
  assign n97111 = pi7683 & ~pi9040;
  assign n97112 = pi7752 & pi9040;
  assign n97113 = ~n97111 & ~n97112;
  assign n97114 = ~pi5475 & ~n97113;
  assign n97115 = pi5475 & n97113;
  assign n97116 = ~n97114 & ~n97115;
  assign n97117 = n97099 & n97116;
  assign n97118 = n97087 & n97117;
  assign n97119 = ~n97107 & n97117;
  assign n97120 = n97093 & n97119;
  assign n97121 = n97099 & ~n97116;
  assign n97122 = ~n97093 & n97121;
  assign n97123 = n97087 & n97116;
  assign n97124 = ~n97122 & ~n97123;
  assign n97125 = ~n97107 & ~n97124;
  assign n97126 = ~n97120 & ~n97125;
  assign n97127 = n97087 & ~n97116;
  assign n97128 = ~n97099 & n97127;
  assign n97129 = n97093 & n97128;
  assign n97130 = n97126 & ~n97129;
  assign n97131 = ~n97118 & n97130;
  assign n97132 = n97110 & n97131;
  assign n97133 = pi7700 & ~pi9040;
  assign n97134 = pi7650 & pi9040;
  assign n97135 = ~n97133 & ~n97134;
  assign n97136 = ~pi5674 & ~n97135;
  assign n97137 = pi5674 & n97135;
  assign n97138 = ~n97136 & ~n97137;
  assign n97139 = ~n97132 & n97138;
  assign n97140 = ~n97093 & n97107;
  assign n97141 = n97128 & n97140;
  assign n97142 = ~n97087 & n97093;
  assign n97143 = n97099 & n97142;
  assign n97144 = n97093 & n97099;
  assign n97145 = ~n97116 & n97144;
  assign n97146 = ~n97143 & ~n97145;
  assign n97147 = n97107 & ~n97146;
  assign n97148 = ~n97141 & ~n97147;
  assign n97149 = ~n97138 & ~n97148;
  assign n97150 = ~n97093 & ~n97107;
  assign n97151 = n97117 & n97150;
  assign n97152 = ~n97087 & n97151;
  assign n97153 = ~n97099 & n97116;
  assign n97154 = n97093 & ~n97107;
  assign n97155 = n97153 & n97154;
  assign n97156 = ~n97116 & n97142;
  assign n97157 = n97099 & n97156;
  assign n97158 = ~n97099 & ~n97116;
  assign n97159 = ~n97087 & n97158;
  assign n97160 = ~n97107 & n97159;
  assign n97161 = ~n97093 & n97160;
  assign n97162 = ~n97157 & ~n97161;
  assign n97163 = ~n97155 & n97162;
  assign n97164 = ~n97152 & n97163;
  assign n97165 = n97087 & n97093;
  assign n97166 = n97153 & n97165;
  assign n97167 = n97164 & ~n97166;
  assign n97168 = ~n97138 & ~n97167;
  assign n97169 = n97108 & n97116;
  assign n97170 = ~n97093 & n97169;
  assign n97171 = ~n97156 & ~n97170;
  assign n97172 = ~n97093 & n97118;
  assign n97173 = n97171 & ~n97172;
  assign n97174 = n97107 & ~n97173;
  assign n97175 = n97087 & ~n97093;
  assign n97176 = ~n97107 & n97175;
  assign n97177 = n97121 & n97176;
  assign n97178 = ~n97174 & ~n97177;
  assign n97179 = ~n97168 & n97178;
  assign n97180 = ~n97149 & n97179;
  assign n97181 = ~n97139 & n97180;
  assign n97182 = n97087 & ~n97099;
  assign n97183 = n97154 & n97182;
  assign n97184 = n97181 & ~n97183;
  assign n97185 = ~pi8556 & ~n97184;
  assign n97186 = pi8556 & ~n97183;
  assign n97187 = n97180 & n97186;
  assign n97188 = ~n97139 & n97187;
  assign po4069 = n97185 | n97188;
  assign n97190 = ~n96990 & n97069;
  assign n97191 = ~n97051 & ~n97060;
  assign n97192 = ~n96996 & ~n97191;
  assign n97193 = ~n97190 & ~n97192;
  assign n97194 = ~n97045 & n97193;
  assign n97195 = n96996 & n97049;
  assign n97196 = ~n97038 & ~n97195;
  assign n97197 = ~n97067 & n97196;
  assign n97198 = n97194 & n97197;
  assign n97199 = n96984 & ~n97198;
  assign n97200 = n96990 & n97066;
  assign n97201 = ~n96990 & n97044;
  assign n97202 = ~n97022 & ~n97201;
  assign n97203 = ~n96996 & n97048;
  assign n97204 = ~n96990 & n97037;
  assign n97205 = ~n97203 & ~n97204;
  assign n97206 = n97202 & n97205;
  assign n97207 = n97008 & n97017;
  assign n97208 = ~n96990 & ~n97002;
  assign n97209 = ~n97207 & ~n97208;
  assign n97210 = ~n97073 & n97209;
  assign n97211 = n96996 & ~n97210;
  assign n97212 = n97206 & ~n97211;
  assign n97213 = ~n97033 & n97212;
  assign n97214 = ~n97200 & n97213;
  assign n97215 = ~n96984 & ~n97214;
  assign n97216 = ~n97199 & ~n97215;
  assign n97217 = pi8602 & ~n97216;
  assign n97218 = ~pi8602 & ~n97199;
  assign n97219 = ~n97215 & n97218;
  assign po4070 = n97217 | n97219;
  assign n97221 = pi7648 & ~pi9040;
  assign n97222 = pi7813 & pi9040;
  assign n97223 = ~n97221 & ~n97222;
  assign n97224 = pi5465 & n97223;
  assign n97225 = ~pi5465 & ~n97223;
  assign n97226 = ~n97224 & ~n97225;
  assign n97227 = pi7660 & ~pi9040;
  assign n97228 = pi7675 & pi9040;
  assign n97229 = ~n97227 & ~n97228;
  assign n97230 = ~pi5431 & n97229;
  assign n97231 = pi5431 & ~n97229;
  assign n97232 = ~n97230 & ~n97231;
  assign n97233 = pi7821 & ~pi9040;
  assign n97234 = pi7658 & pi9040;
  assign n97235 = ~n97233 & ~n97234;
  assign n97236 = ~pi5694 & n97235;
  assign n97237 = pi5694 & ~n97235;
  assign n97238 = ~n97236 & ~n97237;
  assign n97239 = pi7745 & ~pi9040;
  assign n97240 = pi7679 & pi9040;
  assign n97241 = ~n97239 & ~n97240;
  assign n97242 = pi5607 & n97241;
  assign n97243 = ~pi5607 & ~n97241;
  assign n97244 = ~n97242 & ~n97243;
  assign n97245 = ~n97238 & n97244;
  assign n97246 = n97232 & n97245;
  assign n97247 = pi7720 & ~pi9040;
  assign n97248 = pi7670 & pi9040;
  assign n97249 = ~n97247 & ~n97248;
  assign n97250 = ~pi5895 & ~n97249;
  assign n97251 = pi5895 & n97249;
  assign n97252 = ~n97250 & ~n97251;
  assign n97253 = n97246 & ~n97252;
  assign n97254 = n97232 & ~n97252;
  assign n97255 = ~n97244 & n97254;
  assign n97256 = n97238 & n97255;
  assign n97257 = ~n97253 & ~n97256;
  assign n97258 = n97238 & ~n97244;
  assign n97259 = ~n97232 & n97258;
  assign n97260 = n97252 & n97259;
  assign n97261 = ~n97238 & ~n97244;
  assign n97262 = n97232 & n97261;
  assign n97263 = n97252 & n97262;
  assign n97264 = ~n97260 & ~n97263;
  assign n97265 = n97257 & n97264;
  assign n97266 = n97226 & ~n97265;
  assign n97267 = n97238 & n97244;
  assign n97268 = n97232 & n97267;
  assign n97269 = n97252 & n97268;
  assign n97270 = ~n97262 & ~n97269;
  assign n97271 = n97226 & ~n97270;
  assign n97272 = ~n97232 & n97267;
  assign n97273 = ~n97252 & n97272;
  assign n97274 = ~n97226 & n97244;
  assign n97275 = ~n97252 & n97274;
  assign n97276 = ~n97232 & ~n97238;
  assign n97277 = n97252 & n97258;
  assign n97278 = ~n97276 & ~n97277;
  assign n97279 = ~n97226 & ~n97278;
  assign n97280 = ~n97275 & ~n97279;
  assign n97281 = ~n97273 & n97280;
  assign n97282 = n97244 & n97276;
  assign n97283 = n97252 & n97282;
  assign n97284 = n97281 & ~n97283;
  assign n97285 = ~n97271 & n97284;
  assign n97286 = pi7744 & pi9040;
  assign n97287 = pi7658 & ~pi9040;
  assign n97288 = ~n97286 & ~n97287;
  assign n97289 = ~pi5703 & ~n97288;
  assign n97290 = pi5703 & n97288;
  assign n97291 = ~n97289 & ~n97290;
  assign n97292 = ~n97285 & ~n97291;
  assign n97293 = n97232 & n97244;
  assign n97294 = ~n97226 & n97252;
  assign n97295 = n97291 & n97294;
  assign n97296 = n97293 & n97295;
  assign n97297 = ~n97226 & ~n97255;
  assign n97298 = ~n97232 & n97252;
  assign n97299 = n97238 & n97298;
  assign n97300 = ~n97245 & ~n97293;
  assign n97301 = ~n97252 & ~n97300;
  assign n97302 = ~n97232 & n97238;
  assign n97303 = ~n97244 & n97302;
  assign n97304 = ~n97301 & ~n97303;
  assign n97305 = n97226 & n97304;
  assign n97306 = ~n97299 & n97305;
  assign n97307 = ~n97297 & ~n97306;
  assign n97308 = ~n97232 & n97261;
  assign n97309 = n97252 & n97308;
  assign n97310 = ~n97307 & ~n97309;
  assign n97311 = n97291 & ~n97310;
  assign n97312 = ~n97296 & ~n97311;
  assign n97313 = ~n97292 & n97312;
  assign n97314 = ~n97266 & n97313;
  assign n97315 = ~n97226 & ~n97252;
  assign n97316 = n97267 & n97315;
  assign n97317 = ~n97232 & n97316;
  assign n97318 = n97314 & ~n97317;
  assign n97319 = pi8557 & ~n97318;
  assign n97320 = n97313 & ~n97317;
  assign n97321 = ~pi8557 & n97320;
  assign n97322 = ~n97266 & n97321;
  assign po4072 = n97319 | n97322;
  assign n97324 = pi7660 & pi9040;
  assign n97325 = pi7693 & ~pi9040;
  assign n97326 = ~n97324 & ~n97325;
  assign n97327 = pi5813 & n97326;
  assign n97328 = ~pi5813 & ~n97326;
  assign n97329 = ~n97327 & ~n97328;
  assign n97330 = pi7664 & pi9040;
  assign n97331 = pi7813 & ~pi9040;
  assign n97332 = ~n97330 & ~n97331;
  assign n97333 = ~pi5856 & n97332;
  assign n97334 = pi5856 & ~n97332;
  assign n97335 = ~n97333 & ~n97334;
  assign n97336 = ~n97329 & n97335;
  assign n97337 = pi7727 & pi9040;
  assign n97338 = pi7736 & ~pi9040;
  assign n97339 = ~n97337 & ~n97338;
  assign n97340 = pi5550 & n97339;
  assign n97341 = ~pi5550 & ~n97339;
  assign n97342 = ~n97340 & ~n97341;
  assign n97343 = pi7655 & ~pi9040;
  assign n97344 = pi7663 & pi9040;
  assign n97345 = ~n97343 & ~n97344;
  assign n97346 = ~pi5750 & ~n97345;
  assign n97347 = pi5750 & n97345;
  assign n97348 = ~n97346 & ~n97347;
  assign n97349 = pi7664 & ~pi9040;
  assign n97350 = pi7795 & pi9040;
  assign n97351 = ~n97349 & ~n97350;
  assign n97352 = ~pi5585 & ~n97351;
  assign n97353 = pi5585 & n97351;
  assign n97354 = ~n97352 & ~n97353;
  assign n97355 = n97348 & ~n97354;
  assign n97356 = ~n97342 & n97355;
  assign n97357 = pi7727 & ~pi9040;
  assign n97358 = pi7693 & pi9040;
  assign n97359 = ~n97357 & ~n97358;
  assign n97360 = ~pi5512 & ~n97359;
  assign n97361 = pi5512 & n97359;
  assign n97362 = ~n97360 & ~n97361;
  assign n97363 = n97354 & ~n97362;
  assign n97364 = n97348 & n97363;
  assign n97365 = n97342 & n97364;
  assign n97366 = n97354 & n97362;
  assign n97367 = ~n97342 & n97366;
  assign n97368 = ~n97365 & ~n97367;
  assign n97369 = ~n97356 & n97368;
  assign n97370 = n97336 & ~n97369;
  assign n97371 = ~n97342 & ~n97348;
  assign n97372 = ~n97362 & n97371;
  assign n97373 = ~n97354 & ~n97362;
  assign n97374 = n97348 & n97373;
  assign n97375 = n97342 & n97374;
  assign n97376 = ~n97372 & ~n97375;
  assign n97377 = ~n97348 & n97363;
  assign n97378 = n97348 & n97366;
  assign n97379 = ~n97377 & ~n97378;
  assign n97380 = n97376 & n97379;
  assign n97381 = n97329 & ~n97380;
  assign n97382 = ~n97354 & n97362;
  assign n97383 = ~n97348 & n97382;
  assign n97384 = n97342 & n97383;
  assign n97385 = ~n97381 & ~n97384;
  assign n97386 = n97335 & ~n97385;
  assign n97387 = ~n97370 & ~n97386;
  assign n97388 = n97329 & ~n97342;
  assign n97389 = n97348 & n97388;
  assign n97390 = n97362 & n97389;
  assign n97391 = n97354 & n97372;
  assign n97392 = ~n97390 & ~n97391;
  assign n97393 = ~n97348 & n97373;
  assign n97394 = ~n97366 & ~n97373;
  assign n97395 = n97342 & ~n97394;
  assign n97396 = ~n97393 & ~n97395;
  assign n97397 = ~n97329 & ~n97396;
  assign n97398 = n97348 & n97382;
  assign n97399 = ~n97356 & ~n97398;
  assign n97400 = ~n97365 & n97399;
  assign n97401 = n97329 & ~n97400;
  assign n97402 = ~n97397 & ~n97401;
  assign n97403 = ~n97329 & ~n97342;
  assign n97404 = n97363 & n97403;
  assign n97405 = n97342 & n97393;
  assign n97406 = ~n97348 & n97354;
  assign n97407 = n97362 & n97406;
  assign n97408 = n97342 & n97407;
  assign n97409 = ~n97405 & ~n97408;
  assign n97410 = n97362 & n97371;
  assign n97411 = ~n97354 & n97410;
  assign n97412 = n97409 & ~n97411;
  assign n97413 = ~n97404 & n97412;
  assign n97414 = n97402 & n97413;
  assign n97415 = ~n97335 & ~n97414;
  assign n97416 = n97392 & ~n97415;
  assign n97417 = n97387 & n97416;
  assign n97418 = pi8605 & ~n97417;
  assign n97419 = ~pi8605 & n97392;
  assign n97420 = n97387 & n97419;
  assign n97421 = ~n97415 & n97420;
  assign po4075 = n97418 | n97421;
  assign n97423 = n97342 & n97355;
  assign n97424 = ~n97378 & ~n97423;
  assign n97425 = ~n97391 & n97424;
  assign n97426 = n97329 & ~n97425;
  assign n97427 = ~n97342 & n97407;
  assign n97428 = ~n97342 & n97398;
  assign n97429 = ~n97348 & ~n97354;
  assign n97430 = ~n97363 & ~n97429;
  assign n97431 = n97342 & ~n97430;
  assign n97432 = ~n97428 & ~n97431;
  assign n97433 = ~n97427 & n97432;
  assign n97434 = ~n97329 & ~n97433;
  assign n97435 = ~n97426 & ~n97434;
  assign n97436 = ~n97335 & ~n97435;
  assign n97437 = ~n97354 & n97388;
  assign n97438 = ~n97342 & n97354;
  assign n97439 = n97348 & n97438;
  assign n97440 = ~n97423 & ~n97439;
  assign n97441 = ~n97329 & ~n97440;
  assign n97442 = ~n97404 & ~n97441;
  assign n97443 = ~n97342 & n97364;
  assign n97444 = ~n97408 & ~n97443;
  assign n97445 = n97329 & n97342;
  assign n97446 = n97406 & n97445;
  assign n97447 = n97329 & ~n97348;
  assign n97448 = n97362 & n97447;
  assign n97449 = ~n97354 & n97448;
  assign n97450 = ~n97446 & ~n97449;
  assign n97451 = n97444 & n97450;
  assign n97452 = n97442 & n97451;
  assign n97453 = ~n97437 & n97452;
  assign n97454 = n97335 & ~n97453;
  assign n97455 = ~n97329 & n97443;
  assign n97456 = ~n97329 & n97393;
  assign n97457 = ~n97342 & n97456;
  assign n97458 = ~n97455 & ~n97457;
  assign n97459 = n97329 & n97411;
  assign n97460 = n97458 & ~n97459;
  assign n97461 = ~n97342 & n97374;
  assign n97462 = n97342 & n97366;
  assign n97463 = ~n97461 & ~n97462;
  assign n97464 = n97329 & ~n97463;
  assign n97465 = n97460 & ~n97464;
  assign n97466 = ~n97454 & n97465;
  assign n97467 = ~n97436 & n97466;
  assign n97468 = ~pi8592 & ~n97467;
  assign n97469 = pi8592 & n97467;
  assign po4076 = n97468 | n97469;
  assign n97471 = n96990 & n97024;
  assign n97472 = ~n97200 & ~n97471;
  assign n97473 = ~n96996 & n97472;
  assign n97474 = ~n96990 & n97062;
  assign n97475 = ~n97009 & ~n97018;
  assign n97476 = n97017 & ~n97475;
  assign n97477 = n97002 & n97031;
  assign n97478 = ~n96990 & n97018;
  assign n97479 = ~n97477 & ~n97478;
  assign n97480 = n96996 & n97479;
  assign n97481 = ~n97476 & n97480;
  assign n97482 = ~n97474 & n97481;
  assign n97483 = ~n97473 & ~n97482;
  assign n97484 = ~n96990 & n97476;
  assign n97485 = ~n97201 & ~n97484;
  assign n97486 = ~n97483 & n97485;
  assign n97487 = n96984 & ~n97486;
  assign n97488 = ~n96996 & ~n97475;
  assign n97489 = n96990 & n97488;
  assign n97490 = ~n96990 & n97050;
  assign n97491 = ~n97040 & ~n97490;
  assign n97492 = ~n96996 & ~n97491;
  assign n97493 = ~n97017 & n97488;
  assign n97494 = ~n97492 & ~n97493;
  assign n97495 = ~n97489 & n97494;
  assign n97496 = ~n96984 & ~n97495;
  assign n97497 = ~n97487 & ~n97496;
  assign n97498 = ~n96996 & n97022;
  assign n97499 = n96996 & ~n97485;
  assign n97500 = ~n97498 & ~n97499;
  assign n97501 = n96996 & ~n97472;
  assign n97502 = ~n97022 & ~n97501;
  assign n97503 = ~n96984 & ~n97502;
  assign n97504 = n97500 & ~n97503;
  assign n97505 = n97497 & n97504;
  assign n97506 = pi8550 & ~n97505;
  assign n97507 = ~pi8550 & n97504;
  assign n97508 = ~n97496 & n97507;
  assign n97509 = ~n97487 & n97508;
  assign po4081 = n97506 | n97509;
  assign n97511 = pi7703 & ~pi9040;
  assign n97512 = pi7817 & pi9040;
  assign n97513 = ~n97511 & ~n97512;
  assign n97514 = pi5586 & n97513;
  assign n97515 = ~pi5586 & ~n97513;
  assign n97516 = ~n97514 & ~n97515;
  assign n97517 = pi7846 & ~pi9040;
  assign n97518 = pi7741 & pi9040;
  assign n97519 = ~n97517 & ~n97518;
  assign n97520 = pi5795 & n97519;
  assign n97521 = ~pi5795 & ~n97519;
  assign n97522 = ~n97520 & ~n97521;
  assign n97523 = n97516 & n97522;
  assign n97524 = pi7674 & ~pi9040;
  assign n97525 = pi7721 & pi9040;
  assign n97526 = ~n97524 & ~n97525;
  assign n97527 = pi5805 & n97526;
  assign n97528 = ~pi5805 & ~n97526;
  assign n97529 = ~n97527 & ~n97528;
  assign n97530 = pi7651 & pi9040;
  assign n97531 = pi7733 & ~pi9040;
  assign n97532 = ~n97530 & ~n97531;
  assign n97533 = ~pi5534 & ~n97532;
  assign n97534 = pi5534 & n97532;
  assign n97535 = ~n97533 & ~n97534;
  assign n97536 = n97529 & ~n97535;
  assign n97537 = n97523 & n97536;
  assign n97538 = pi7703 & pi9040;
  assign n97539 = pi7752 & ~pi9040;
  assign n97540 = ~n97538 & ~n97539;
  assign n97541 = ~pi5748 & n97540;
  assign n97542 = pi5748 & ~n97540;
  assign n97543 = ~n97541 & ~n97542;
  assign n97544 = n97535 & n97543;
  assign n97545 = n97529 & n97544;
  assign n97546 = n97522 & n97545;
  assign n97547 = ~n97516 & n97546;
  assign n97548 = ~n97537 & ~n97547;
  assign n97549 = pi7723 & pi9040;
  assign n97550 = pi7651 & ~pi9040;
  assign n97551 = ~n97549 & ~n97550;
  assign n97552 = ~pi5749 & ~n97551;
  assign n97553 = pi5749 & n97551;
  assign n97554 = ~n97552 & ~n97553;
  assign n97555 = ~n97535 & ~n97543;
  assign n97556 = n97522 & n97555;
  assign n97557 = ~n97516 & n97556;
  assign n97558 = ~n97529 & n97544;
  assign n97559 = n97516 & ~n97529;
  assign n97560 = n97535 & n97559;
  assign n97561 = ~n97558 & ~n97560;
  assign n97562 = n97522 & ~n97561;
  assign n97563 = ~n97557 & ~n97562;
  assign n97564 = n97535 & ~n97543;
  assign n97565 = ~n97522 & n97564;
  assign n97566 = ~n97516 & n97565;
  assign n97567 = ~n97535 & n97543;
  assign n97568 = ~n97529 & n97567;
  assign n97569 = ~n97522 & n97568;
  assign n97570 = ~n97566 & ~n97569;
  assign n97571 = n97563 & n97570;
  assign n97572 = n97529 & n97567;
  assign n97573 = n97516 & n97572;
  assign n97574 = ~n97516 & n97568;
  assign n97575 = ~n97516 & n97529;
  assign n97576 = n97535 & n97575;
  assign n97577 = ~n97574 & ~n97576;
  assign n97578 = ~n97573 & n97577;
  assign n97579 = n97571 & n97578;
  assign n97580 = ~n97554 & ~n97579;
  assign n97581 = n97529 & n97564;
  assign n97582 = n97516 & n97581;
  assign n97583 = ~n97529 & n97555;
  assign n97584 = n97516 & n97583;
  assign n97585 = ~n97582 & ~n97584;
  assign n97586 = ~n97574 & n97585;
  assign n97587 = ~n97522 & ~n97586;
  assign n97588 = ~n97543 & n97575;
  assign n97589 = ~n97535 & n97588;
  assign n97590 = ~n97558 & ~n97589;
  assign n97591 = n97516 & n97544;
  assign n97592 = n97590 & ~n97591;
  assign n97593 = ~n97522 & ~n97592;
  assign n97594 = ~n97529 & n97564;
  assign n97595 = ~n97516 & n97522;
  assign n97596 = n97594 & n97595;
  assign n97597 = n97585 & ~n97596;
  assign n97598 = n97522 & n97572;
  assign n97599 = n97597 & ~n97598;
  assign n97600 = ~n97593 & n97599;
  assign n97601 = n97554 & ~n97600;
  assign n97602 = ~n97587 & ~n97601;
  assign n97603 = ~n97580 & n97602;
  assign n97604 = n97548 & n97603;
  assign n97605 = ~pi8554 & n97604;
  assign n97606 = pi8554 & ~n97604;
  assign po4082 = n97605 | n97606;
  assign n97608 = n97529 & n97555;
  assign n97609 = n97516 & n97608;
  assign n97610 = n97516 & n97564;
  assign n97611 = ~n97516 & n97583;
  assign n97612 = ~n97610 & ~n97611;
  assign n97613 = ~n97522 & ~n97612;
  assign n97614 = ~n97609 & ~n97613;
  assign n97615 = n97522 & n97568;
  assign n97616 = n97516 & n97556;
  assign n97617 = ~n97615 & ~n97616;
  assign n97618 = n97614 & n97617;
  assign n97619 = n97516 & n97545;
  assign n97620 = ~n97516 & n97572;
  assign n97621 = ~n97619 & ~n97620;
  assign n97622 = n97618 & n97621;
  assign n97623 = n97554 & ~n97622;
  assign n97624 = ~n97522 & ~n97554;
  assign n97625 = ~n97535 & n97559;
  assign n97626 = ~n97529 & n97543;
  assign n97627 = ~n97625 & ~n97626;
  assign n97628 = n97624 & ~n97627;
  assign n97629 = ~n97516 & n97535;
  assign n97630 = ~n97529 & n97629;
  assign n97631 = ~n97589 & ~n97630;
  assign n97632 = n97523 & n97529;
  assign n97633 = ~n97555 & n97632;
  assign n97634 = ~n97546 & ~n97633;
  assign n97635 = n97631 & n97634;
  assign n97636 = ~n97554 & ~n97635;
  assign n97637 = ~n97522 & n97558;
  assign n97638 = ~n97516 & n97637;
  assign n97639 = ~n97516 & n97581;
  assign n97640 = ~n97620 & ~n97639;
  assign n97641 = ~n97522 & ~n97640;
  assign n97642 = ~n97638 & ~n97641;
  assign n97643 = n97522 & n97589;
  assign n97644 = n97642 & ~n97643;
  assign n97645 = ~n97636 & n97644;
  assign n97646 = ~n97628 & n97645;
  assign n97647 = ~n97623 & n97646;
  assign n97648 = ~n97596 & n97647;
  assign n97649 = ~pi8579 & ~n97648;
  assign n97650 = pi8579 & ~n97596;
  assign n97651 = n97646 & n97650;
  assign n97652 = ~n97623 & n97651;
  assign po4083 = n97649 | n97652;
  assign n97654 = ~n97393 & ~n97398;
  assign n97655 = ~n97329 & ~n97654;
  assign n97656 = n97342 & n97378;
  assign n97657 = ~n97655 & ~n97656;
  assign n97658 = n97342 & n97354;
  assign n97659 = ~n97406 & ~n97658;
  assign n97660 = ~n97374 & n97659;
  assign n97661 = n97329 & ~n97660;
  assign n97662 = n97657 & ~n97661;
  assign n97663 = n97335 & ~n97662;
  assign n97664 = ~n97329 & n97427;
  assign n97665 = ~n97455 & ~n97664;
  assign n97666 = ~n97459 & n97665;
  assign n97667 = ~n97342 & n97348;
  assign n97668 = ~n97362 & n97667;
  assign n97669 = ~n97411 & ~n97668;
  assign n97670 = n97329 & n97439;
  assign n97671 = n97342 & n97398;
  assign n97672 = ~n97329 & n97406;
  assign n97673 = ~n97671 & ~n97672;
  assign n97674 = ~n97405 & n97673;
  assign n97675 = ~n97670 & n97674;
  assign n97676 = n97669 & n97675;
  assign n97677 = ~n97449 & n97676;
  assign n97678 = ~n97335 & ~n97677;
  assign n97679 = n97666 & ~n97678;
  assign n97680 = ~n97663 & n97679;
  assign n97681 = ~pi8633 & ~n97680;
  assign n97682 = ~n97663 & ~n97678;
  assign n97683 = n97666 & n97682;
  assign n97684 = pi8633 & n97683;
  assign po4091 = n97681 | n97684;
  assign n97686 = pi7650 & ~pi9040;
  assign n97687 = pi7686 & pi9040;
  assign n97688 = ~n97686 & ~n97687;
  assign n97689 = ~pi5534 & ~n97688;
  assign n97690 = pi5534 & n97688;
  assign n97691 = ~n97689 & ~n97690;
  assign n97692 = pi7721 & ~pi9040;
  assign n97693 = pi7700 & pi9040;
  assign n97694 = ~n97692 & ~n97693;
  assign n97695 = ~pi5446 & n97694;
  assign n97696 = pi5446 & ~n97694;
  assign n97697 = ~n97695 & ~n97696;
  assign n97698 = pi7803 & ~pi9040;
  assign n97699 = pi7668 & pi9040;
  assign n97700 = ~n97698 & ~n97699;
  assign n97701 = ~pi5650 & n97700;
  assign n97702 = pi5650 & ~n97700;
  assign n97703 = ~n97701 & ~n97702;
  assign n97704 = pi7686 & ~pi9040;
  assign n97705 = pi7846 & pi9040;
  assign n97706 = ~n97704 & ~n97705;
  assign n97707 = ~pi5587 & n97706;
  assign n97708 = pi5587 & ~n97706;
  assign n97709 = ~n97707 & ~n97708;
  assign n97710 = pi7683 & pi9040;
  assign n97711 = pi7689 & ~pi9040;
  assign n97712 = ~n97710 & ~n97711;
  assign n97713 = ~pi5805 & n97712;
  assign n97714 = pi5805 & ~n97712;
  assign n97715 = ~n97713 & ~n97714;
  assign n97716 = n97709 & n97715;
  assign n97717 = ~n97703 & n97716;
  assign n97718 = n97709 & ~n97715;
  assign n97719 = n97703 & n97718;
  assign n97720 = ~n97717 & ~n97719;
  assign n97721 = ~n97697 & ~n97720;
  assign n97722 = pi7677 & ~pi9040;
  assign n97723 = pi7733 & pi9040;
  assign n97724 = ~n97722 & ~n97723;
  assign n97725 = ~pi5798 & n97724;
  assign n97726 = pi5798 & ~n97724;
  assign n97727 = ~n97725 & ~n97726;
  assign n97728 = ~n97709 & n97715;
  assign n97729 = ~n97697 & n97703;
  assign n97730 = n97728 & n97729;
  assign n97731 = n97727 & n97730;
  assign n97732 = ~n97721 & ~n97731;
  assign n97733 = n97691 & ~n97732;
  assign n97734 = ~n97709 & ~n97715;
  assign n97735 = ~n97709 & n97727;
  assign n97736 = ~n97734 & ~n97735;
  assign n97737 = n97703 & ~n97736;
  assign n97738 = n97718 & ~n97727;
  assign n97739 = ~n97737 & ~n97738;
  assign n97740 = n97697 & ~n97739;
  assign n97741 = n97703 & n97727;
  assign n97742 = ~n97716 & ~n97734;
  assign n97743 = n97741 & ~n97742;
  assign n97744 = ~n97740 & ~n97743;
  assign n97745 = n97718 & n97727;
  assign n97746 = ~n97703 & n97745;
  assign n97747 = ~n97703 & ~n97736;
  assign n97748 = n97703 & ~n97727;
  assign n97749 = n97715 & n97748;
  assign n97750 = ~n97747 & ~n97749;
  assign n97751 = ~n97697 & ~n97750;
  assign n97752 = ~n97746 & ~n97751;
  assign n97753 = n97744 & n97752;
  assign n97754 = ~n97691 & ~n97753;
  assign n97755 = ~n97703 & ~n97727;
  assign n97756 = ~n97734 & n97755;
  assign n97757 = n97691 & n97756;
  assign n97758 = ~n97703 & n97727;
  assign n97759 = n97734 & n97758;
  assign n97760 = ~n97697 & n97759;
  assign n97761 = n97697 & ~n97703;
  assign n97762 = ~n97727 & n97761;
  assign n97763 = n97715 & n97762;
  assign n97764 = ~n97760 & ~n97763;
  assign n97765 = ~n97757 & n97764;
  assign n97766 = ~n97703 & ~n97709;
  assign n97767 = n97716 & ~n97727;
  assign n97768 = ~n97766 & ~n97767;
  assign n97769 = n97691 & n97697;
  assign n97770 = ~n97768 & n97769;
  assign n97771 = n97765 & ~n97770;
  assign n97772 = ~n97754 & n97771;
  assign n97773 = ~n97733 & n97772;
  assign n97774 = ~pi8629 & ~n97773;
  assign n97775 = pi8629 & n97773;
  assign po4092 = n97774 | n97775;
  assign n97777 = ~n96996 & n97049;
  assign n97778 = n96990 & n97207;
  assign n97779 = ~n97478 & ~n97778;
  assign n97780 = ~n97017 & n97050;
  assign n97781 = n97779 & ~n97780;
  assign n97782 = ~n96996 & ~n97781;
  assign n97783 = n97031 & ~n97475;
  assign n97784 = ~n97066 & ~n97783;
  assign n97785 = ~n97201 & n97784;
  assign n97786 = n96996 & ~n97785;
  assign n97787 = ~n96990 & n97019;
  assign n97788 = ~n97786 & ~n97787;
  assign n97789 = ~n97782 & n97788;
  assign n97790 = n96984 & ~n97789;
  assign n97791 = ~n97777 & ~n97790;
  assign n97792 = n96990 & n97018;
  assign n97793 = ~n97044 & ~n97792;
  assign n97794 = ~n96996 & ~n97793;
  assign n97795 = ~n97067 & ~n97794;
  assign n97796 = ~n97040 & ~n97049;
  assign n97797 = ~n96990 & n97073;
  assign n97798 = ~n97207 & ~n97797;
  assign n97799 = ~n97780 & n97798;
  assign n97800 = n96996 & ~n97799;
  assign n97801 = n96990 & n97019;
  assign n97802 = ~n97800 & ~n97801;
  assign n97803 = n97796 & n97802;
  assign n97804 = n97795 & n97803;
  assign n97805 = ~n96984 & ~n97804;
  assign n97806 = ~n97054 & ~n97474;
  assign n97807 = n96996 & ~n97806;
  assign n97808 = ~n97805 & ~n97807;
  assign n97809 = n97791 & n97808;
  assign n97810 = pi8561 & n97809;
  assign n97811 = ~pi8561 & ~n97809;
  assign po4093 = n97810 | n97811;
  assign n97813 = n97342 & n97348;
  assign n97814 = n97362 & n97813;
  assign n97815 = ~n97342 & ~n97354;
  assign n97816 = ~n97668 & ~n97815;
  assign n97817 = ~n97329 & ~n97816;
  assign n97818 = n97329 & n97366;
  assign n97819 = ~n97342 & n97818;
  assign n97820 = ~n97461 & ~n97819;
  assign n97821 = ~n97817 & n97820;
  assign n97822 = ~n97814 & n97821;
  assign n97823 = ~n97335 & ~n97822;
  assign n97824 = ~n97374 & ~n97384;
  assign n97825 = ~n97329 & ~n97824;
  assign n97826 = ~n97364 & ~n97408;
  assign n97827 = ~n97342 & n97382;
  assign n97828 = n97826 & ~n97827;
  assign n97829 = n97329 & ~n97828;
  assign n97830 = n97366 & n97403;
  assign n97831 = ~n97391 & ~n97830;
  assign n97832 = ~n97829 & n97831;
  assign n97833 = ~n97825 & n97832;
  assign n97834 = n97335 & ~n97833;
  assign n97835 = ~n97823 & ~n97834;
  assign n97836 = n97342 & n97379;
  assign n97837 = ~n97342 & ~n97373;
  assign n97838 = ~n97836 & ~n97837;
  assign n97839 = ~n97329 & n97838;
  assign n97840 = ~n97364 & n97654;
  assign n97841 = n97445 & ~n97840;
  assign n97842 = ~n97839 & ~n97841;
  assign n97843 = n97835 & n97842;
  assign n97844 = ~pi8570 & ~n97843;
  assign n97845 = pi8570 & n97842;
  assign n97846 = ~n97834 & n97845;
  assign n97847 = ~n97823 & n97846;
  assign po4095 = n97844 | n97847;
  assign n97849 = n97543 & n97559;
  assign n97850 = n97535 & n97849;
  assign n97851 = ~n97574 & ~n97850;
  assign n97852 = n97522 & ~n97851;
  assign n97853 = ~n97546 & ~n97589;
  assign n97854 = ~n97535 & n97575;
  assign n97855 = ~n97630 & ~n97854;
  assign n97856 = ~n97522 & ~n97855;
  assign n97857 = n97516 & ~n97522;
  assign n97858 = n97567 & n97857;
  assign n97859 = ~n97529 & n97858;
  assign n97860 = n97522 & ~n97529;
  assign n97861 = ~n97543 & n97860;
  assign n97862 = ~n97535 & n97861;
  assign n97863 = ~n97582 & ~n97862;
  assign n97864 = ~n97859 & n97863;
  assign n97865 = ~n97856 & n97864;
  assign n97866 = n97853 & n97865;
  assign n97867 = n97554 & ~n97866;
  assign n97868 = ~n97522 & n97589;
  assign n97869 = ~n97547 & ~n97868;
  assign n97870 = ~n97867 & n97869;
  assign n97871 = ~n97852 & n97870;
  assign n97872 = n97522 & n97529;
  assign n97873 = ~n97543 & n97872;
  assign n97874 = n97535 & n97873;
  assign n97875 = ~n97516 & ~n97529;
  assign n97876 = ~n97543 & n97875;
  assign n97877 = n97535 & n97876;
  assign n97878 = ~n97537 & ~n97615;
  assign n97879 = ~n97877 & n97878;
  assign n97880 = ~n97874 & n97879;
  assign n97881 = ~n97529 & ~n97543;
  assign n97882 = ~n97591 & ~n97881;
  assign n97883 = ~n97522 & ~n97882;
  assign n97884 = n97880 & ~n97883;
  assign n97885 = ~n97573 & n97884;
  assign n97886 = ~n97574 & n97885;
  assign n97887 = ~n97554 & ~n97886;
  assign n97888 = n97871 & ~n97887;
  assign n97889 = ~pi8503 & ~n97888;
  assign n97890 = pi8503 & n97871;
  assign n97891 = ~n97887 & n97890;
  assign po4096 = n97889 | n97891;
  assign n97893 = n97697 & n97735;
  assign n97894 = ~n97703 & n97893;
  assign n97895 = ~n97727 & n97734;
  assign n97896 = n97703 & n97716;
  assign n97897 = ~n97745 & ~n97896;
  assign n97898 = ~n97895 & n97897;
  assign n97899 = n97697 & ~n97898;
  assign n97900 = n97727 & n97734;
  assign n97901 = ~n97738 & ~n97900;
  assign n97902 = ~n97697 & ~n97901;
  assign n97903 = ~n97899 & ~n97902;
  assign n97904 = ~n97727 & n97728;
  assign n97905 = ~n97697 & n97904;
  assign n97906 = n97727 & n97896;
  assign n97907 = ~n97905 & ~n97906;
  assign n97908 = n97903 & n97907;
  assign n97909 = ~n97691 & ~n97908;
  assign n97910 = n97703 & n97728;
  assign n97911 = ~n97717 & ~n97910;
  assign n97912 = n97697 & ~n97911;
  assign n97913 = ~n97703 & n97738;
  assign n97914 = ~n97912 & ~n97913;
  assign n97915 = ~n97697 & n97767;
  assign n97916 = n97727 & n97728;
  assign n97917 = ~n97895 & ~n97916;
  assign n97918 = ~n97915 & n97917;
  assign n97919 = ~n97745 & n97918;
  assign n97920 = n97703 & ~n97919;
  assign n97921 = n97914 & ~n97920;
  assign n97922 = n97691 & ~n97921;
  assign n97923 = ~n97909 & ~n97922;
  assign n97924 = ~n97894 & n97923;
  assign n97925 = n97715 & n97755;
  assign n97926 = ~n97709 & n97925;
  assign n97927 = n97717 & n97727;
  assign n97928 = ~n97926 & ~n97927;
  assign n97929 = ~n97697 & ~n97928;
  assign n97930 = n97924 & ~n97929;
  assign n97931 = ~pi8520 & ~n97930;
  assign n97932 = n97923 & ~n97929;
  assign n97933 = pi8520 & n97932;
  assign n97934 = ~n97894 & n97933;
  assign po4100 = n97931 | n97934;
  assign n97936 = ~n97253 & ~n97260;
  assign n97937 = ~n97226 & ~n97936;
  assign n97938 = ~n97317 & ~n97937;
  assign n97939 = n97232 & n97238;
  assign n97940 = n97226 & n97939;
  assign n97941 = n97252 & n97940;
  assign n97942 = n97252 & n97267;
  assign n97943 = ~n97939 & ~n97942;
  assign n97944 = ~n97232 & ~n97252;
  assign n97945 = ~n97238 & n97944;
  assign n97946 = n97943 & ~n97945;
  assign n97947 = n97226 & ~n97946;
  assign n97948 = ~n97263 & ~n97947;
  assign n97949 = ~n97291 & ~n97948;
  assign n97950 = ~n97226 & n97245;
  assign n97951 = n97252 & n97950;
  assign n97952 = ~n97226 & n97303;
  assign n97953 = ~n97951 & ~n97952;
  assign n97954 = ~n97291 & ~n97953;
  assign n97955 = ~n97949 & ~n97954;
  assign n97956 = ~n97941 & n97955;
  assign n97957 = ~n97238 & n97254;
  assign n97958 = ~n97255 & ~n97272;
  assign n97959 = ~n97308 & n97958;
  assign n97960 = ~n97226 & ~n97959;
  assign n97961 = ~n97244 & n97944;
  assign n97962 = n97238 & n97961;
  assign n97963 = ~n97282 & ~n97962;
  assign n97964 = n97226 & ~n97963;
  assign n97965 = ~n97960 & ~n97964;
  assign n97966 = ~n97957 & n97965;
  assign n97967 = ~n97269 & ~n97309;
  assign n97968 = n97966 & n97967;
  assign n97969 = n97291 & ~n97968;
  assign n97970 = n97956 & ~n97969;
  assign n97971 = n97938 & n97970;
  assign n97972 = ~pi8685 & ~n97971;
  assign n97973 = pi8685 & n97956;
  assign n97974 = n97938 & n97973;
  assign n97975 = ~n97969 & n97974;
  assign po4105 = n97972 | n97975;
  assign n97977 = pi7705 & ~pi9040;
  assign n97978 = pi7708 & pi9040;
  assign n97979 = ~n97977 & ~n97978;
  assign n97980 = pi5598 & n97979;
  assign n97981 = ~pi5598 & ~n97979;
  assign n97982 = ~n97980 & ~n97981;
  assign n97983 = pi7684 & ~pi9040;
  assign n97984 = pi7803 & pi9040;
  assign n97985 = ~n97983 & ~n97984;
  assign n97986 = ~pi5690 & n97985;
  assign n97987 = pi5690 & ~n97985;
  assign n97988 = ~n97986 & ~n97987;
  assign n97989 = pi7674 & pi9040;
  assign n97990 = pi7723 & ~pi9040;
  assign n97991 = ~n97989 & ~n97990;
  assign n97992 = pi5798 & n97991;
  assign n97993 = ~pi5798 & ~n97991;
  assign n97994 = ~n97992 & ~n97993;
  assign n97995 = pi7708 & ~pi9040;
  assign n97996 = pi7649 & pi9040;
  assign n97997 = ~n97995 & ~n97996;
  assign n97998 = ~pi5674 & n97997;
  assign n97999 = pi5674 & ~n97997;
  assign n98000 = ~n97998 & ~n97999;
  assign n98001 = pi7698 & pi9040;
  assign n98002 = pi7649 & ~pi9040;
  assign n98003 = ~n98001 & ~n98002;
  assign n98004 = ~pi5475 & n98003;
  assign n98005 = pi5475 & ~n98003;
  assign n98006 = ~n98004 & ~n98005;
  assign n98007 = ~n98000 & ~n98006;
  assign n98008 = ~n97994 & n98007;
  assign n98009 = ~n97988 & n98008;
  assign n98010 = ~n97988 & n98006;
  assign n98011 = n98000 & n98010;
  assign n98012 = ~n98009 & ~n98011;
  assign n98013 = ~n97982 & ~n98012;
  assign n98014 = pi7746 & pi9040;
  assign n98015 = pi7661 & ~pi9040;
  assign n98016 = ~n98014 & ~n98015;
  assign n98017 = ~pi5587 & n98016;
  assign n98018 = pi5587 & ~n98016;
  assign n98019 = ~n98017 & ~n98018;
  assign n98020 = n97982 & n97988;
  assign n98021 = ~n98000 & n98020;
  assign n98022 = ~n97994 & ~n98000;
  assign n98023 = n98006 & n98022;
  assign n98024 = ~pi5798 & n97991;
  assign n98025 = pi5798 & ~n97991;
  assign n98026 = ~n98024 & ~n98025;
  assign n98027 = ~n98000 & ~n98026;
  assign n98028 = ~n98006 & n98027;
  assign n98029 = ~n98023 & ~n98028;
  assign n98030 = ~n97994 & n98000;
  assign n98031 = ~n98006 & n98030;
  assign n98032 = ~n97988 & n98031;
  assign n98033 = n98029 & ~n98032;
  assign n98034 = n97982 & ~n98033;
  assign n98035 = ~n98021 & ~n98034;
  assign n98036 = n98000 & ~n98026;
  assign n98037 = n98006 & n98036;
  assign n98038 = ~n97988 & n98037;
  assign n98039 = n98035 & ~n98038;
  assign n98040 = n97988 & n98030;
  assign n98041 = n98000 & ~n98006;
  assign n98042 = ~n98026 & n98041;
  assign n98043 = ~n98040 & ~n98042;
  assign n98044 = ~n97982 & ~n98043;
  assign n98045 = n98006 & n98027;
  assign n98046 = n97988 & n98045;
  assign n98047 = ~n98044 & ~n98046;
  assign n98048 = n98039 & n98047;
  assign n98049 = ~n98019 & ~n98048;
  assign n98050 = ~n98013 & ~n98049;
  assign n98051 = n97982 & n98019;
  assign n98052 = ~n98043 & n98051;
  assign n98053 = n98006 & n98030;
  assign n98054 = ~n98045 & ~n98053;
  assign n98055 = ~n97988 & ~n98054;
  assign n98056 = ~n98009 & ~n98055;
  assign n98057 = n98019 & ~n98056;
  assign n98058 = ~n98052 & ~n98057;
  assign n98059 = ~n97982 & n98019;
  assign n98060 = n97988 & n98022;
  assign n98061 = ~n98037 & ~n98060;
  assign n98062 = ~n98007 & n98061;
  assign n98063 = n98059 & ~n98062;
  assign n98064 = n98058 & ~n98063;
  assign n98065 = n98050 & n98064;
  assign n98066 = ~pi8549 & ~n98065;
  assign n98067 = pi8549 & n98058;
  assign n98068 = n98050 & n98067;
  assign n98069 = ~n98063 & n98068;
  assign po4122 = n98066 | n98069;
  assign n98071 = n97093 & n97159;
  assign n98072 = n97093 & n97118;
  assign n98073 = ~n98071 & ~n98072;
  assign n98074 = n97107 & ~n98073;
  assign n98075 = n97140 & n97169;
  assign n98076 = ~n98074 & ~n98075;
  assign n98077 = ~n97183 & n98076;
  assign n98078 = ~n97087 & n97117;
  assign n98079 = ~n97107 & n98078;
  assign n98080 = ~n97166 & ~n97177;
  assign n98081 = ~n97161 & n98080;
  assign n98082 = ~n98079 & n98081;
  assign n98083 = n97138 & ~n98082;
  assign n98084 = ~n97087 & n97099;
  assign n98085 = ~n97116 & n98084;
  assign n98086 = ~n97107 & n98085;
  assign n98087 = n97093 & n98086;
  assign n98088 = ~n97093 & n97128;
  assign n98089 = ~n97118 & ~n98088;
  assign n98090 = ~n98085 & n98089;
  assign n98091 = n97107 & ~n98090;
  assign n98092 = n97138 & n98091;
  assign n98093 = ~n97093 & n97119;
  assign n98094 = ~n97087 & ~n97093;
  assign n98095 = n97116 & n98094;
  assign n98096 = ~n98093 & ~n98095;
  assign n98097 = ~n98086 & n98096;
  assign n98098 = ~n97116 & n97165;
  assign n98099 = ~n97093 & n97153;
  assign n98100 = ~n97108 & ~n98099;
  assign n98101 = n97107 & ~n98100;
  assign n98102 = ~n98098 & ~n98101;
  assign n98103 = n98097 & n98102;
  assign n98104 = ~n97138 & ~n98103;
  assign n98105 = ~n98092 & ~n98104;
  assign n98106 = ~n98087 & n98105;
  assign n98107 = ~n98083 & n98106;
  assign n98108 = n98077 & n98107;
  assign n98109 = pi8594 & ~n98108;
  assign n98110 = ~pi8594 & n98077;
  assign n98111 = n98107 & n98110;
  assign po4125 = n98109 | n98111;
  assign n98113 = ~n97252 & n97282;
  assign n98114 = n97252 & n97293;
  assign n98115 = ~n97272 & ~n98114;
  assign n98116 = n97226 & ~n98115;
  assign n98117 = ~n98113 & ~n98116;
  assign n98118 = ~n97226 & n97261;
  assign n98119 = n97252 & n98118;
  assign n98120 = ~n97252 & n97950;
  assign n98121 = ~n98119 & ~n98120;
  assign n98122 = ~n97952 & n98121;
  assign n98123 = ~n97256 & ~n97269;
  assign n98124 = ~n97244 & n97298;
  assign n98125 = n98123 & ~n98124;
  assign n98126 = n98122 & n98125;
  assign n98127 = n98117 & n98126;
  assign n98128 = ~n97291 & ~n98127;
  assign n98129 = n97232 & n97258;
  assign n98130 = ~n97272 & ~n98129;
  assign n98131 = n97252 & ~n98130;
  assign n98132 = ~n97308 & ~n97957;
  assign n98133 = ~n97232 & n97244;
  assign n98134 = n97252 & n98133;
  assign n98135 = n98132 & ~n98134;
  assign n98136 = n97226 & ~n98135;
  assign n98137 = ~n97252 & n97267;
  assign n98138 = n97232 & n97252;
  assign n98139 = n97244 & n98138;
  assign n98140 = ~n97238 & n98139;
  assign n98141 = ~n98137 & ~n98140;
  assign n98142 = ~n97226 & ~n98141;
  assign n98143 = ~n97252 & n97262;
  assign n98144 = ~n98142 & ~n98143;
  assign n98145 = ~n98136 & n98144;
  assign n98146 = ~n98131 & n98145;
  assign n98147 = n97291 & ~n98146;
  assign n98148 = n97226 & n97255;
  assign n98149 = ~n98147 & ~n98148;
  assign n98150 = n97276 & n97315;
  assign n98151 = n97244 & n98150;
  assign n98152 = n98149 & ~n98151;
  assign n98153 = ~n98128 & n98152;
  assign n98154 = ~pi8559 & ~n98153;
  assign n98155 = pi8559 & n98149;
  assign n98156 = ~n98128 & n98155;
  assign n98157 = ~n98151 & n98156;
  assign po4142 = n98154 | n98157;
  assign n98159 = ~n97166 & ~n98084;
  assign n98160 = ~n97100 & n98159;
  assign n98161 = ~n97107 & ~n98160;
  assign n98162 = ~n97099 & n97140;
  assign n98163 = ~n98071 & ~n98095;
  assign n98164 = n97087 & n97099;
  assign n98165 = n97093 & n97107;
  assign n98166 = n98164 & n98165;
  assign n98167 = n98163 & ~n98166;
  assign n98168 = ~n98162 & n98167;
  assign n98169 = ~n98161 & n98168;
  assign n98170 = n97138 & ~n98169;
  assign n98171 = ~n97093 & n98085;
  assign n98172 = n97093 & n98078;
  assign n98173 = ~n98171 & ~n98172;
  assign n98174 = ~n97107 & ~n98173;
  assign n98175 = ~n98170 & ~n98174;
  assign n98176 = ~n97093 & n97159;
  assign n98177 = ~n97128 & ~n97169;
  assign n98178 = ~n97107 & ~n98177;
  assign n98179 = ~n98176 & ~n98178;
  assign n98180 = ~n97172 & n98179;
  assign n98181 = ~n97138 & ~n98180;
  assign n98182 = ~n97121 & ~n97153;
  assign n98183 = n97087 & ~n98182;
  assign n98184 = ~n97145 & ~n98183;
  assign n98185 = n97107 & ~n98184;
  assign n98186 = ~n97138 & n98185;
  assign n98187 = ~n98181 & ~n98186;
  assign n98188 = n98175 & n98187;
  assign n98189 = pi8575 & ~n98188;
  assign n98190 = ~pi8575 & n98175;
  assign n98191 = n98187 & n98190;
  assign po4145 = n98189 | n98191;
  assign n98193 = pi7662 & pi9040;
  assign n98194 = pi7670 & ~pi9040;
  assign n98195 = ~n98193 & ~n98194;
  assign n98196 = pi5585 & n98195;
  assign n98197 = ~pi5585 & ~n98195;
  assign n98198 = ~n98196 & ~n98197;
  assign n98199 = pi7749 & pi9040;
  assign n98200 = pi7659 & ~pi9040;
  assign n98201 = ~n98199 & ~n98200;
  assign n98202 = pi5888 & n98201;
  assign n98203 = ~pi5888 & ~n98201;
  assign n98204 = ~n98202 & ~n98203;
  assign n98205 = pi7725 & ~pi9040;
  assign n98206 = pi7726 & pi9040;
  assign n98207 = ~n98205 & ~n98206;
  assign n98208 = ~pi5749 & ~n98207;
  assign n98209 = pi5749 & n98207;
  assign n98210 = ~n98208 & ~n98209;
  assign n98211 = pi7653 & pi9040;
  assign n98212 = pi7711 & ~pi9040;
  assign n98213 = ~n98211 & ~n98212;
  assign n98214 = ~pi5748 & ~n98213;
  assign n98215 = pi5748 & n98213;
  assign n98216 = ~n98214 & ~n98215;
  assign n98217 = pi7711 & pi9040;
  assign n98218 = pi7795 & ~pi9040;
  assign n98219 = ~n98217 & ~n98218;
  assign n98220 = pi5750 & n98219;
  assign n98221 = ~pi5750 & ~n98219;
  assign n98222 = ~n98220 & ~n98221;
  assign n98223 = n98216 & ~n98222;
  assign n98224 = n98210 & n98223;
  assign n98225 = n98204 & n98224;
  assign n98226 = ~n98204 & n98216;
  assign n98227 = n98222 & n98226;
  assign n98228 = pi7666 & pi9040;
  assign n98229 = pi7663 & ~pi9040;
  assign n98230 = ~n98228 & ~n98229;
  assign n98231 = ~pi5692 & n98230;
  assign n98232 = pi5692 & ~n98230;
  assign n98233 = ~n98231 & ~n98232;
  assign n98234 = ~n98210 & n98226;
  assign n98235 = n98210 & n98222;
  assign n98236 = ~n98216 & n98235;
  assign n98237 = ~n98234 & ~n98236;
  assign n98238 = n98233 & ~n98237;
  assign n98239 = ~n98227 & ~n98238;
  assign n98240 = n98216 & n98235;
  assign n98241 = ~n98210 & ~n98216;
  assign n98242 = ~n98204 & ~n98216;
  assign n98243 = ~n98222 & n98242;
  assign n98244 = ~n98210 & ~n98222;
  assign n98245 = n98204 & n98244;
  assign n98246 = ~n98243 & ~n98245;
  assign n98247 = ~n98241 & n98246;
  assign n98248 = ~n98240 & n98247;
  assign n98249 = ~n98233 & ~n98248;
  assign n98250 = n98239 & ~n98249;
  assign n98251 = ~n98225 & n98250;
  assign n98252 = n98198 & ~n98251;
  assign n98253 = ~n98210 & n98222;
  assign n98254 = ~n98216 & n98253;
  assign n98255 = ~n98204 & n98254;
  assign n98256 = n98204 & ~n98216;
  assign n98257 = ~n98222 & n98256;
  assign n98258 = ~n98210 & n98257;
  assign n98259 = ~n98225 & ~n98258;
  assign n98260 = ~n98255 & n98259;
  assign n98261 = ~n98233 & ~n98260;
  assign n98262 = ~n98252 & ~n98261;
  assign n98263 = ~n98204 & n98240;
  assign n98264 = n98210 & ~n98216;
  assign n98265 = n98233 & n98264;
  assign n98266 = n98204 & n98265;
  assign n98267 = n98223 & ~n98233;
  assign n98268 = ~n98204 & n98267;
  assign n98269 = n98216 & n98253;
  assign n98270 = n98204 & n98269;
  assign n98271 = ~n98268 & ~n98270;
  assign n98272 = ~n98204 & n98233;
  assign n98273 = n98241 & n98272;
  assign n98274 = ~n98210 & n98216;
  assign n98275 = n98204 & n98274;
  assign n98276 = n98210 & ~n98222;
  assign n98277 = ~n98216 & n98276;
  assign n98278 = ~n98275 & ~n98277;
  assign n98279 = n98233 & ~n98278;
  assign n98280 = ~n98273 & ~n98279;
  assign n98281 = n98271 & n98280;
  assign n98282 = ~n98198 & ~n98281;
  assign n98283 = ~n98266 & ~n98282;
  assign n98284 = ~n98263 & n98283;
  assign n98285 = n98262 & n98284;
  assign n98286 = ~pi8547 & ~n98285;
  assign n98287 = ~n98252 & ~n98263;
  assign n98288 = ~n98261 & n98287;
  assign n98289 = n98283 & n98288;
  assign n98290 = pi8547 & n98289;
  assign po4159 = n98286 | n98290;
  assign n98292 = ~n97116 & n98094;
  assign n98293 = ~n97123 & ~n98292;
  assign n98294 = ~n98085 & n98293;
  assign n98295 = ~n97107 & ~n98294;
  assign n98296 = ~n97093 & n98183;
  assign n98297 = ~n97127 & ~n98078;
  assign n98298 = n97107 & ~n98297;
  assign n98299 = ~n98296 & ~n98298;
  assign n98300 = ~n98295 & n98299;
  assign n98301 = n97093 & n97169;
  assign n98302 = n98300 & ~n98301;
  assign n98303 = ~n97138 & ~n98302;
  assign n98304 = n97154 & ~n98297;
  assign n98305 = ~n97118 & ~n97128;
  assign n98306 = ~n97169 & ~n98085;
  assign n98307 = n98305 & n98306;
  assign n98308 = ~n97093 & ~n98307;
  assign n98309 = ~n98304 & ~n98308;
  assign n98310 = ~n98071 & n98309;
  assign n98311 = n97138 & ~n98310;
  assign n98312 = ~n98303 & ~n98311;
  assign n98313 = ~n97093 & n98078;
  assign n98314 = ~n98301 & ~n98313;
  assign n98315 = n97107 & ~n98314;
  assign n98316 = n98312 & ~n98315;
  assign n98317 = pi8615 & ~n98316;
  assign n98318 = ~pi8615 & ~n98315;
  assign n98319 = ~n98311 & n98318;
  assign n98320 = ~n98303 & n98319;
  assign po4160 = n98317 | n98320;
  assign n98322 = ~n97619 & ~n97625;
  assign n98323 = n97554 & ~n98322;
  assign n98324 = ~n97588 & ~n97854;
  assign n98325 = ~n97608 & n98324;
  assign n98326 = ~n97522 & ~n98325;
  assign n98327 = n97554 & n98326;
  assign n98328 = ~n98323 & ~n98327;
  assign n98329 = n97545 & n97857;
  assign n98330 = ~n97859 & ~n98329;
  assign n98331 = ~n97630 & ~n97881;
  assign n98332 = n97522 & ~n98331;
  assign n98333 = n97554 & n98332;
  assign n98334 = n98330 & ~n98333;
  assign n98335 = ~n97516 & n97545;
  assign n98336 = ~n97516 & n97567;
  assign n98337 = ~n97850 & ~n98336;
  assign n98338 = n97522 & ~n98337;
  assign n98339 = ~n97582 & ~n97589;
  assign n98340 = ~n97516 & n97544;
  assign n98341 = ~n97594 & ~n98340;
  assign n98342 = ~n97522 & ~n98341;
  assign n98343 = n98339 & ~n98342;
  assign n98344 = ~n98338 & n98343;
  assign n98345 = ~n98335 & n98344;
  assign n98346 = ~n97554 & ~n98345;
  assign n98347 = ~n97573 & n97585;
  assign n98348 = n97522 & ~n98347;
  assign n98349 = ~n98346 & ~n98348;
  assign n98350 = n98334 & n98349;
  assign n98351 = n98328 & n98350;
  assign n98352 = ~pi8583 & ~n98351;
  assign n98353 = pi8583 & n98334;
  assign n98354 = n98328 & n98353;
  assign n98355 = n98349 & n98354;
  assign po4161 = n98352 | n98355;
  assign n98357 = ~n97988 & n98053;
  assign n98358 = n97988 & n98007;
  assign n98359 = ~n98357 & ~n98358;
  assign n98360 = n97982 & ~n98359;
  assign n98361 = ~n97988 & n98042;
  assign n98362 = n97988 & n98037;
  assign n98363 = ~n98361 & ~n98362;
  assign n98364 = ~n97982 & ~n98363;
  assign n98365 = ~n97982 & ~n97988;
  assign n98366 = ~n98030 & ~n98045;
  assign n98367 = n98365 & ~n98366;
  assign n98368 = ~n97982 & n98030;
  assign n98369 = n98006 & n98368;
  assign n98370 = ~n98367 & ~n98369;
  assign n98371 = ~n98019 & ~n98370;
  assign n98372 = n97988 & ~n98006;
  assign n98373 = n98027 & n98372;
  assign n98374 = ~n98007 & ~n98372;
  assign n98375 = n97982 & ~n98374;
  assign n98376 = n97988 & n98023;
  assign n98377 = ~n98375 & ~n98376;
  assign n98378 = ~n98373 & n98377;
  assign n98379 = ~n98019 & ~n98378;
  assign n98380 = ~n98371 & ~n98379;
  assign n98381 = ~n98007 & ~n98022;
  assign n98382 = ~n97988 & ~n98381;
  assign n98383 = ~n98037 & ~n98382;
  assign n98384 = ~n97982 & ~n98383;
  assign n98385 = n97988 & n97994;
  assign n98386 = ~n97982 & n98006;
  assign n98387 = n98385 & n98386;
  assign n98388 = ~n98006 & n98026;
  assign n98389 = ~n98037 & ~n98388;
  assign n98390 = n97988 & ~n98389;
  assign n98391 = n97982 & ~n97988;
  assign n98392 = n98027 & n98391;
  assign n98393 = n98006 & n98392;
  assign n98394 = ~n98390 & ~n98393;
  assign n98395 = ~n98387 & n98394;
  assign n98396 = ~n98384 & n98395;
  assign n98397 = ~n98361 & n98396;
  assign n98398 = n98019 & ~n98397;
  assign n98399 = n98380 & ~n98398;
  assign n98400 = ~n98364 & n98399;
  assign n98401 = ~n98360 & n98400;
  assign n98402 = pi8600 & n98401;
  assign n98403 = ~pi8600 & ~n98401;
  assign po4165 = n98402 | n98403;
  assign n98405 = n97727 & n97766;
  assign n98406 = ~n97717 & ~n98405;
  assign n98407 = ~n97719 & ~n97767;
  assign n98408 = n98406 & n98407;
  assign n98409 = ~n97697 & ~n98408;
  assign n98410 = ~n97703 & n97916;
  assign n98411 = ~n98409 & ~n98410;
  assign n98412 = ~n97691 & ~n98411;
  assign n98413 = n97697 & n97895;
  assign n98414 = ~n97703 & n98413;
  assign n98415 = ~n97703 & n97718;
  assign n98416 = ~n97743 & ~n98415;
  assign n98417 = ~n97904 & n98416;
  assign n98418 = ~n97691 & n97697;
  assign n98419 = ~n98417 & n98418;
  assign n98420 = ~n98414 & ~n98419;
  assign n98421 = ~n98412 & n98420;
  assign n98422 = ~n97697 & n97738;
  assign n98423 = n97703 & n98422;
  assign n98424 = ~n97731 & ~n98423;
  assign n98425 = n97697 & n97745;
  assign n98426 = n97703 & n98425;
  assign n98427 = n97715 & n97741;
  assign n98428 = ~n97709 & n98427;
  assign n98429 = ~n98426 & ~n98428;
  assign n98430 = ~n97741 & ~n97742;
  assign n98431 = n97697 & n98430;
  assign n98432 = ~n97718 & n97727;
  assign n98433 = n97729 & n98432;
  assign n98434 = ~n97709 & ~n97727;
  assign n98435 = ~n97703 & n98434;
  assign n98436 = ~n98415 & ~n98435;
  assign n98437 = ~n97697 & ~n98436;
  assign n98438 = ~n98433 & ~n98437;
  assign n98439 = ~n98431 & n98438;
  assign n98440 = n98429 & n98439;
  assign n98441 = n97691 & ~n98440;
  assign n98442 = n98424 & ~n98441;
  assign n98443 = ~pi8528 & n98442;
  assign n98444 = n98421 & n98443;
  assign n98445 = n98421 & n98442;
  assign n98446 = pi8528 & ~n98445;
  assign po4166 = n98444 | n98446;
  assign n98448 = ~n97309 & ~n98143;
  assign n98449 = n97226 & ~n98448;
  assign n98450 = ~n97291 & n97293;
  assign n98451 = ~n97226 & n98450;
  assign n98452 = n97238 & n97944;
  assign n98453 = ~n98133 & ~n98452;
  assign n98454 = ~n97262 & n98453;
  assign n98455 = n97226 & ~n98454;
  assign n98456 = ~n97252 & n97268;
  assign n98457 = ~n98455 & ~n98456;
  assign n98458 = ~n97291 & ~n98457;
  assign n98459 = ~n98451 & ~n98458;
  assign n98460 = ~n97256 & ~n97260;
  assign n98461 = ~n97252 & n97308;
  assign n98462 = ~n98114 & ~n98461;
  assign n98463 = n98460 & n98462;
  assign n98464 = ~n97226 & ~n98463;
  assign n98465 = ~n97252 & n98133;
  assign n98466 = n97232 & n97294;
  assign n98467 = ~n97238 & n98466;
  assign n98468 = ~n97260 & ~n98467;
  assign n98469 = ~n98140 & n98468;
  assign n98470 = ~n98465 & n98469;
  assign n98471 = n97226 & n98129;
  assign n98472 = n98470 & ~n98471;
  assign n98473 = n97291 & ~n98472;
  assign n98474 = ~n98464 & ~n98473;
  assign n98475 = n98459 & n98474;
  assign n98476 = ~n98449 & n98475;
  assign n98477 = pi8678 & n98476;
  assign n98478 = ~pi8678 & ~n98476;
  assign po4169 = n98477 | n98478;
  assign n98480 = n98216 & n98244;
  assign n98481 = n98204 & n98480;
  assign n98482 = n98204 & n98254;
  assign n98483 = ~n98481 & ~n98482;
  assign n98484 = ~n98210 & n98243;
  assign n98485 = ~n98236 & ~n98484;
  assign n98486 = ~n98233 & ~n98485;
  assign n98487 = n98483 & ~n98486;
  assign n98488 = n98210 & n98272;
  assign n98489 = n98487 & ~n98488;
  assign n98490 = n98198 & ~n98489;
  assign n98491 = ~n98204 & ~n98233;
  assign n98492 = n98277 & n98491;
  assign n98493 = ~n98234 & ~n98492;
  assign n98494 = n98259 & n98493;
  assign n98495 = ~n98236 & ~n98269;
  assign n98496 = ~n98204 & n98253;
  assign n98497 = n98495 & ~n98496;
  assign n98498 = n98233 & ~n98497;
  assign n98499 = ~n98233 & n98240;
  assign n98500 = ~n98498 & ~n98499;
  assign n98501 = n98494 & n98500;
  assign n98502 = ~n98198 & ~n98501;
  assign n98503 = n98204 & n98277;
  assign n98504 = n98233 & n98503;
  assign n98505 = ~n98502 & ~n98504;
  assign n98506 = ~n98490 & n98505;
  assign n98507 = n98269 & n98491;
  assign n98508 = n98204 & n98267;
  assign n98509 = ~n98507 & ~n98508;
  assign n98510 = ~n98233 & n98482;
  assign n98511 = n98509 & ~n98510;
  assign n98512 = n98506 & n98511;
  assign n98513 = ~pi8548 & ~n98512;
  assign n98514 = pi8548 & n98511;
  assign n98515 = n98505 & n98514;
  assign n98516 = ~n98490 & n98515;
  assign po4170 = n98513 | n98516;
  assign n98518 = n98010 & n98026;
  assign n98519 = ~n98045 & ~n98518;
  assign n98520 = ~n97982 & ~n98519;
  assign n98521 = ~n97988 & n98000;
  assign n98522 = ~n98026 & n98521;
  assign n98523 = n97988 & n98006;
  assign n98524 = ~n97994 & n98523;
  assign n98525 = ~n98522 & ~n98524;
  assign n98526 = n97982 & ~n98525;
  assign n98527 = n97988 & n98031;
  assign n98528 = ~n98387 & ~n98527;
  assign n98529 = ~n98009 & n98528;
  assign n98530 = ~n98526 & n98529;
  assign n98531 = ~n98520 & n98530;
  assign n98532 = ~n98361 & ~n98373;
  assign n98533 = n98531 & n98532;
  assign n98534 = ~n98019 & ~n98533;
  assign n98535 = n98022 & n98372;
  assign n98536 = n98054 & ~n98535;
  assign n98537 = n97982 & ~n98536;
  assign n98538 = n97988 & n98042;
  assign n98539 = ~n98537 & ~n98538;
  assign n98540 = n98020 & n98036;
  assign n98541 = ~n98000 & n98010;
  assign n98542 = ~n97988 & n98027;
  assign n98543 = ~n98541 & ~n98542;
  assign n98544 = n97982 & ~n98543;
  assign n98545 = ~n98540 & ~n98544;
  assign n98546 = n98539 & n98545;
  assign n98547 = n98019 & ~n98546;
  assign n98548 = ~n98031 & ~n98376;
  assign n98549 = ~n98038 & n98548;
  assign n98550 = n98059 & ~n98549;
  assign n98551 = ~n98547 & ~n98550;
  assign n98552 = ~n98009 & ~n98373;
  assign n98553 = ~n97982 & ~n98552;
  assign n98554 = n98551 & ~n98553;
  assign n98555 = ~n98534 & n98554;
  assign n98556 = ~pi8585 & n98555;
  assign n98557 = pi8585 & ~n98555;
  assign po4173 = n98556 | n98557;
  assign n98559 = ~n97715 & n97748;
  assign n98560 = n97917 & ~n98559;
  assign n98561 = n97769 & ~n98560;
  assign n98562 = n97718 & n97761;
  assign n98563 = ~n97727 & n98562;
  assign n98564 = ~n97742 & n97758;
  assign n98565 = ~n98563 & ~n98564;
  assign n98566 = ~n97926 & n98565;
  assign n98567 = ~n97742 & n97748;
  assign n98568 = ~n98428 & ~n98567;
  assign n98569 = ~n97727 & n97729;
  assign n98570 = n97709 & n98569;
  assign n98571 = ~n98426 & ~n98570;
  assign n98572 = n98568 & n98571;
  assign n98573 = n98566 & n98572;
  assign n98574 = ~n97691 & ~n98573;
  assign n98575 = n97691 & n97767;
  assign n98576 = ~n97703 & n98575;
  assign n98577 = ~n97715 & n97727;
  assign n98578 = ~n98415 & ~n98577;
  assign n98579 = ~n97697 & ~n98578;
  assign n98580 = ~n97905 & ~n98579;
  assign n98581 = n97691 & ~n98580;
  assign n98582 = ~n98576 & ~n98581;
  assign n98583 = ~n97715 & n97758;
  assign n98584 = ~n97906 & ~n98583;
  assign n98585 = ~n97697 & ~n98584;
  assign n98586 = n98582 & ~n98585;
  assign n98587 = ~n98574 & n98586;
  assign n98588 = ~n98561 & n98587;
  assign n98589 = ~pi8582 & ~n98588;
  assign n98590 = pi8582 & n98586;
  assign n98591 = ~n98561 & n98590;
  assign n98592 = ~n98574 & n98591;
  assign po4188 = n98589 | n98592;
  assign n98594 = ~n98204 & n98480;
  assign n98595 = ~n98254 & ~n98263;
  assign n98596 = n98204 & n98223;
  assign n98597 = ~n98204 & n98277;
  assign n98598 = ~n98596 & ~n98597;
  assign n98599 = n98595 & n98598;
  assign n98600 = n98233 & ~n98599;
  assign n98601 = ~n98216 & n98244;
  assign n98602 = n98204 & n98235;
  assign n98603 = ~n98234 & ~n98602;
  assign n98604 = ~n98601 & n98603;
  assign n98605 = ~n98233 & ~n98604;
  assign n98606 = n98222 & n98256;
  assign n98607 = n98210 & n98606;
  assign n98608 = ~n98605 & ~n98607;
  assign n98609 = ~n98600 & n98608;
  assign n98610 = ~n98594 & n98609;
  assign n98611 = ~n98198 & ~n98610;
  assign n98612 = n98204 & n98233;
  assign n98613 = n98240 & n98612;
  assign n98614 = n98233 & n98601;
  assign n98615 = n98233 & n98269;
  assign n98616 = ~n98614 & ~n98615;
  assign n98617 = ~n98204 & ~n98616;
  assign n98618 = ~n98613 & ~n98617;
  assign n98619 = ~n98204 & n98224;
  assign n98620 = ~n98503 & ~n98619;
  assign n98621 = n98204 & n98253;
  assign n98622 = ~n98204 & n98235;
  assign n98623 = ~n98621 & ~n98622;
  assign n98624 = ~n98224 & n98623;
  assign n98625 = ~n98254 & n98624;
  assign n98626 = ~n98233 & ~n98625;
  assign n98627 = ~n98204 & n98236;
  assign n98628 = ~n98626 & ~n98627;
  assign n98629 = n98620 & n98628;
  assign n98630 = n98618 & n98629;
  assign n98631 = n98198 & ~n98630;
  assign n98632 = n98233 & ~n98483;
  assign n98633 = ~n98631 & ~n98632;
  assign n98634 = ~n98258 & ~n98619;
  assign n98635 = ~n98233 & ~n98634;
  assign n98636 = n98633 & ~n98635;
  assign n98637 = ~n98611 & n98636;
  assign n98638 = pi8601 & ~n98637;
  assign n98639 = ~pi8601 & n98637;
  assign po4190 = n98638 | n98639;
  assign n98641 = ~n97982 & n98042;
  assign n98642 = n97988 & n98027;
  assign n98643 = ~n98023 & ~n98642;
  assign n98644 = ~n97982 & ~n98643;
  assign n98645 = n97982 & ~n98389;
  assign n98646 = ~n98357 & ~n98645;
  assign n98647 = ~n98644 & n98646;
  assign n98648 = ~n98019 & ~n98647;
  assign n98649 = ~n98641 & ~n98648;
  assign n98650 = n97982 & n98028;
  assign n98651 = ~n97988 & n98045;
  assign n98652 = ~n98006 & n98365;
  assign n98653 = ~n98523 & ~n98652;
  assign n98654 = n98000 & ~n98653;
  assign n98655 = ~n98524 & ~n98654;
  assign n98656 = ~n98009 & n98655;
  assign n98657 = ~n98651 & n98656;
  assign n98658 = ~n98650 & n98657;
  assign n98659 = n98019 & ~n98658;
  assign n98660 = ~n98527 & ~n98542;
  assign n98661 = n97982 & ~n98660;
  assign n98662 = ~n98659 & ~n98661;
  assign n98663 = n98649 & n98662;
  assign n98664 = pi8624 & n98663;
  assign n98665 = ~pi8624 & ~n98663;
  assign po4202 = n98664 | n98665;
  assign n98667 = ~n98484 & ~n98619;
  assign n98668 = ~n98607 & n98667;
  assign n98669 = n98233 & ~n98668;
  assign n98670 = ~n98503 & ~n98615;
  assign n98671 = ~n98480 & ~n98622;
  assign n98672 = ~n98233 & ~n98671;
  assign n98673 = ~n98263 & ~n98672;
  assign n98674 = n98670 & n98673;
  assign n98675 = n98198 & ~n98674;
  assign n98676 = ~n98216 & n98222;
  assign n98677 = ~n98241 & ~n98676;
  assign n98678 = n98204 & ~n98677;
  assign n98679 = ~n98224 & ~n98496;
  assign n98680 = ~n98233 & ~n98679;
  assign n98681 = n98204 & n98222;
  assign n98682 = ~n98236 & ~n98681;
  assign n98683 = ~n98244 & n98682;
  assign n98684 = n98233 & ~n98683;
  assign n98685 = ~n98680 & ~n98684;
  assign n98686 = ~n98678 & n98685;
  assign n98687 = ~n98198 & ~n98686;
  assign n98688 = ~n98675 & ~n98687;
  assign n98689 = ~n98492 & ~n98510;
  assign n98690 = n98688 & n98689;
  assign n98691 = ~n98669 & n98690;
  assign n98692 = ~pi8622 & ~n98691;
  assign n98693 = pi8622 & n98689;
  assign n98694 = ~n98669 & n98693;
  assign n98695 = n98688 & n98694;
  assign po4219 = n98692 | n98695;
  assign n98697 = pi7942 & ~pi9040;
  assign n98698 = pi7978 & pi9040;
  assign n98699 = ~n98697 & ~n98698;
  assign n98700 = pi8748 & n98699;
  assign n98701 = ~pi8748 & ~n98699;
  assign n98702 = ~n98700 & ~n98701;
  assign n98703 = pi7999 & ~pi9040;
  assign n98704 = pi7979 & pi9040;
  assign n98705 = ~n98703 & ~n98704;
  assign n98706 = ~pi8803 & ~n98705;
  assign n98707 = pi8803 & n98705;
  assign n98708 = ~n98706 & ~n98707;
  assign n98709 = pi7954 & ~pi9040;
  assign n98710 = pi8033 & pi9040;
  assign n98711 = ~n98709 & ~n98710;
  assign n98712 = ~pi8738 & ~n98711;
  assign n98713 = pi8738 & n98711;
  assign n98714 = ~n98712 & ~n98713;
  assign n98715 = pi7997 & ~pi9040;
  assign n98716 = pi7940 & pi9040;
  assign n98717 = ~n98715 & ~n98716;
  assign n98718 = ~pi8727 & n98717;
  assign n98719 = pi8727 & ~n98717;
  assign n98720 = ~n98718 & ~n98719;
  assign n98721 = n98714 & n98720;
  assign n98722 = n98708 & n98721;
  assign n98723 = n98702 & n98722;
  assign n98724 = pi8028 & pi9040;
  assign n98725 = pi8004 & ~pi9040;
  assign n98726 = ~n98724 & ~n98725;
  assign n98727 = ~pi8742 & ~n98726;
  assign n98728 = pi8742 & n98726;
  assign n98729 = ~n98727 & ~n98728;
  assign n98730 = ~n98702 & n98729;
  assign n98731 = ~n98708 & n98730;
  assign n98732 = n98720 & n98731;
  assign n98733 = ~n98723 & ~n98732;
  assign n98734 = pi7991 & pi9040;
  assign n98735 = pi7958 & ~pi9040;
  assign n98736 = ~n98734 & ~n98735;
  assign n98737 = ~pi8802 & ~n98736;
  assign n98738 = pi8802 & n98736;
  assign n98739 = ~n98737 & ~n98738;
  assign n98740 = ~n98714 & ~n98739;
  assign n98741 = n98708 & n98730;
  assign n98742 = ~n98720 & n98741;
  assign n98743 = n98708 & ~n98729;
  assign n98744 = n98720 & n98743;
  assign n98745 = n98702 & n98729;
  assign n98746 = n98720 & n98745;
  assign n98747 = ~n98744 & ~n98746;
  assign n98748 = ~n98742 & n98747;
  assign n98749 = n98740 & ~n98748;
  assign n98750 = ~n98708 & n98720;
  assign n98751 = ~n98702 & n98750;
  assign n98752 = ~n98702 & ~n98729;
  assign n98753 = n98708 & n98752;
  assign n98754 = ~n98720 & n98753;
  assign n98755 = ~n98751 & ~n98754;
  assign n98756 = n98708 & n98745;
  assign n98757 = ~n98731 & ~n98756;
  assign n98758 = n98755 & n98757;
  assign n98759 = n98714 & ~n98758;
  assign n98760 = n98702 & ~n98729;
  assign n98761 = ~n98708 & n98760;
  assign n98762 = ~n98720 & n98761;
  assign n98763 = ~n98759 & ~n98762;
  assign n98764 = ~n98739 & ~n98763;
  assign n98765 = ~n98749 & ~n98764;
  assign n98766 = ~n98745 & ~n98752;
  assign n98767 = ~n98720 & ~n98766;
  assign n98768 = ~n98708 & n98752;
  assign n98769 = ~n98767 & ~n98768;
  assign n98770 = ~n98714 & ~n98769;
  assign n98771 = n98708 & n98760;
  assign n98772 = ~n98744 & ~n98771;
  assign n98773 = ~n98742 & n98772;
  assign n98774 = n98714 & ~n98773;
  assign n98775 = ~n98770 & ~n98774;
  assign n98776 = ~n98714 & n98720;
  assign n98777 = n98730 & n98776;
  assign n98778 = ~n98708 & ~n98720;
  assign n98779 = ~n98702 & n98778;
  assign n98780 = ~n98729 & n98779;
  assign n98781 = ~n98708 & n98729;
  assign n98782 = n98702 & n98781;
  assign n98783 = ~n98720 & n98782;
  assign n98784 = ~n98780 & ~n98783;
  assign n98785 = n98720 & n98761;
  assign n98786 = n98784 & ~n98785;
  assign n98787 = ~n98777 & n98786;
  assign n98788 = n98775 & n98787;
  assign n98789 = n98739 & ~n98788;
  assign n98790 = n98765 & ~n98789;
  assign n98791 = n98733 & n98790;
  assign n98792 = pi8696 & ~n98791;
  assign n98793 = ~pi8696 & n98733;
  assign n98794 = n98765 & n98793;
  assign n98795 = ~n98789 & n98794;
  assign po5661 = n98792 | n98795;
  assign n98797 = ~n98720 & n98743;
  assign n98798 = ~n98756 & ~n98797;
  assign n98799 = ~n98732 & n98798;
  assign n98800 = n98714 & ~n98799;
  assign n98801 = n98720 & n98782;
  assign n98802 = n98720 & n98771;
  assign n98803 = ~n98708 & ~n98729;
  assign n98804 = ~n98730 & ~n98803;
  assign n98805 = ~n98720 & ~n98804;
  assign n98806 = ~n98802 & ~n98805;
  assign n98807 = ~n98801 & n98806;
  assign n98808 = ~n98714 & ~n98807;
  assign n98809 = ~n98800 & ~n98808;
  assign n98810 = n98739 & ~n98809;
  assign n98811 = n98721 & ~n98729;
  assign n98812 = n98708 & n98720;
  assign n98813 = n98729 & n98812;
  assign n98814 = ~n98797 & ~n98813;
  assign n98815 = ~n98714 & ~n98814;
  assign n98816 = ~n98777 & ~n98815;
  assign n98817 = ~n98702 & n98812;
  assign n98818 = n98729 & n98817;
  assign n98819 = ~n98783 & ~n98818;
  assign n98820 = n98714 & n98781;
  assign n98821 = ~n98720 & n98820;
  assign n98822 = n98714 & n98761;
  assign n98823 = ~n98821 & ~n98822;
  assign n98824 = n98819 & n98823;
  assign n98825 = n98816 & n98824;
  assign n98826 = ~n98811 & n98825;
  assign n98827 = ~n98739 & ~n98826;
  assign n98828 = ~n98714 & n98768;
  assign n98829 = n98720 & n98828;
  assign n98830 = ~n98714 & n98818;
  assign n98831 = ~n98829 & ~n98830;
  assign n98832 = n98721 & n98760;
  assign n98833 = ~n98708 & n98832;
  assign n98834 = n98831 & ~n98833;
  assign n98835 = n98720 & n98753;
  assign n98836 = ~n98720 & n98745;
  assign n98837 = ~n98835 & ~n98836;
  assign n98838 = n98714 & ~n98837;
  assign n98839 = n98834 & ~n98838;
  assign n98840 = ~n98827 & n98839;
  assign n98841 = ~n98810 & n98840;
  assign n98842 = ~pi8716 & ~n98841;
  assign n98843 = pi8716 & n98841;
  assign po5676 = n98842 | n98843;
  assign n98845 = pi8016 & pi9040;
  assign n98846 = pi7998 & ~pi9040;
  assign n98847 = ~n98845 & ~n98846;
  assign n98848 = ~pi8776 & n98847;
  assign n98849 = pi8776 & ~n98847;
  assign n98850 = ~n98848 & ~n98849;
  assign n98851 = pi7972 & pi9040;
  assign n98852 = pi7974 & ~pi9040;
  assign n98853 = ~n98851 & ~n98852;
  assign n98854 = ~pi8719 & n98853;
  assign n98855 = pi8719 & ~n98853;
  assign n98856 = ~n98854 & ~n98855;
  assign n98857 = pi8034 & ~pi9040;
  assign n98858 = pi7975 & pi9040;
  assign n98859 = ~n98857 & ~n98858;
  assign n98860 = ~pi8715 & n98859;
  assign n98861 = pi8715 & ~n98859;
  assign n98862 = ~n98860 & ~n98861;
  assign n98863 = pi8005 & ~pi9040;
  assign n98864 = pi7952 & pi9040;
  assign n98865 = ~n98863 & ~n98864;
  assign n98866 = ~pi8796 & n98865;
  assign n98867 = pi8796 & ~n98865;
  assign n98868 = ~n98866 & ~n98867;
  assign n98869 = ~n98862 & n98868;
  assign n98870 = n98856 & n98869;
  assign n98871 = pi7935 & ~pi9040;
  assign n98872 = pi7929 & pi9040;
  assign n98873 = ~n98871 & ~n98872;
  assign n98874 = pi8798 & n98873;
  assign n98875 = ~pi8798 & ~n98873;
  assign n98876 = ~n98874 & ~n98875;
  assign n98877 = ~n98856 & ~n98868;
  assign n98878 = ~n98876 & n98877;
  assign n98879 = ~n98870 & ~n98878;
  assign n98880 = pi7931 & pi9040;
  assign n98881 = pi8000 & ~pi9040;
  assign n98882 = ~n98880 & ~n98881;
  assign n98883 = ~pi8761 & ~n98882;
  assign n98884 = pi8761 & n98882;
  assign n98885 = ~n98883 & ~n98884;
  assign n98886 = n98868 & n98885;
  assign n98887 = n98856 & n98886;
  assign n98888 = n98876 & n98886;
  assign n98889 = n98862 & n98888;
  assign n98890 = n98868 & ~n98885;
  assign n98891 = ~n98862 & n98890;
  assign n98892 = n98856 & n98885;
  assign n98893 = ~n98891 & ~n98892;
  assign n98894 = n98876 & ~n98893;
  assign n98895 = ~n98889 & ~n98894;
  assign n98896 = n98856 & ~n98885;
  assign n98897 = ~n98868 & n98896;
  assign n98898 = n98862 & n98897;
  assign n98899 = n98895 & ~n98898;
  assign n98900 = ~n98887 & n98899;
  assign n98901 = n98879 & n98900;
  assign n98902 = ~n98850 & ~n98901;
  assign n98903 = n98856 & ~n98862;
  assign n98904 = n98876 & n98903;
  assign n98905 = n98890 & n98904;
  assign n98906 = ~n98862 & ~n98876;
  assign n98907 = n98897 & n98906;
  assign n98908 = ~n98856 & n98862;
  assign n98909 = n98868 & n98908;
  assign n98910 = n98862 & n98868;
  assign n98911 = ~n98885 & n98910;
  assign n98912 = ~n98909 & ~n98911;
  assign n98913 = ~n98876 & ~n98912;
  assign n98914 = ~n98907 & ~n98913;
  assign n98915 = n98850 & ~n98914;
  assign n98916 = ~n98885 & n98908;
  assign n98917 = n98877 & n98885;
  assign n98918 = ~n98862 & n98917;
  assign n98919 = ~n98916 & ~n98918;
  assign n98920 = ~n98862 & n98887;
  assign n98921 = n98919 & ~n98920;
  assign n98922 = ~n98876 & ~n98921;
  assign n98923 = ~n98862 & n98876;
  assign n98924 = n98886 & n98923;
  assign n98925 = ~n98856 & n98924;
  assign n98926 = ~n98868 & n98885;
  assign n98927 = n98862 & n98876;
  assign n98928 = n98926 & n98927;
  assign n98929 = n98868 & n98916;
  assign n98930 = ~n98868 & ~n98885;
  assign n98931 = ~n98856 & n98930;
  assign n98932 = n98876 & n98931;
  assign n98933 = ~n98862 & n98932;
  assign n98934 = ~n98929 & ~n98933;
  assign n98935 = ~n98928 & n98934;
  assign n98936 = ~n98925 & n98935;
  assign n98937 = n98856 & n98862;
  assign n98938 = n98926 & n98937;
  assign n98939 = n98936 & ~n98938;
  assign n98940 = n98850 & ~n98939;
  assign n98941 = ~n98922 & ~n98940;
  assign n98942 = ~n98915 & n98941;
  assign n98943 = ~n98905 & n98942;
  assign n98944 = ~n98902 & n98943;
  assign n98945 = ~n98868 & n98927;
  assign n98946 = n98856 & n98945;
  assign n98947 = n98944 & ~n98946;
  assign n98948 = ~pi8754 & ~n98947;
  assign n98949 = pi8754 & ~n98946;
  assign n98950 = ~n98902 & n98949;
  assign n98951 = n98943 & n98950;
  assign po5695 = n98948 | n98951;
  assign n98953 = pi8015 & pi9040;
  assign n98954 = pi8013 & ~pi9040;
  assign n98955 = ~n98953 & ~n98954;
  assign n98956 = pi8766 & n98955;
  assign n98957 = ~pi8766 & ~n98955;
  assign n98958 = ~n98956 & ~n98957;
  assign n98959 = pi7965 & ~pi9040;
  assign n98960 = pi8001 & pi9040;
  assign n98961 = ~n98959 & ~n98960;
  assign n98962 = pi8705 & n98961;
  assign n98963 = ~pi8705 & ~n98961;
  assign n98964 = ~n98962 & ~n98963;
  assign n98965 = pi7991 & ~pi9040;
  assign n98966 = pi8003 & pi9040;
  assign n98967 = ~n98965 & ~n98966;
  assign n98968 = pi8719 & n98967;
  assign n98969 = ~pi8719 & ~n98967;
  assign n98970 = ~n98968 & ~n98969;
  assign n98971 = pi7954 & pi9040;
  assign n98972 = pi7968 & ~pi9040;
  assign n98973 = ~n98971 & ~n98972;
  assign n98974 = ~pi8712 & n98973;
  assign n98975 = pi8712 & ~n98973;
  assign n98976 = ~n98974 & ~n98975;
  assign n98977 = n98970 & ~n98976;
  assign n98978 = ~n98964 & n98977;
  assign n98979 = pi7940 & ~pi9040;
  assign n98980 = pi7946 & pi9040;
  assign n98981 = ~n98979 & ~n98980;
  assign n98982 = pi8807 & n98981;
  assign n98983 = ~pi8807 & ~n98981;
  assign n98984 = ~n98982 & ~n98983;
  assign n98985 = n98978 & ~n98984;
  assign n98986 = ~n98970 & n98976;
  assign n98987 = ~n98964 & n98986;
  assign n98988 = ~n98984 & n98987;
  assign n98989 = ~n98985 & ~n98988;
  assign n98990 = n98964 & n98984;
  assign n98991 = n98976 & n98990;
  assign n98992 = ~n98970 & n98991;
  assign n98993 = n98970 & n98976;
  assign n98994 = ~n98964 & n98993;
  assign n98995 = n98984 & n98994;
  assign n98996 = ~n98992 & ~n98995;
  assign n98997 = n98989 & n98996;
  assign n98998 = n98958 & ~n98997;
  assign n98999 = ~n98970 & ~n98976;
  assign n99000 = ~n98964 & n98999;
  assign n99001 = n98984 & n99000;
  assign n99002 = ~n98994 & ~n99001;
  assign n99003 = n98958 & ~n99002;
  assign n99004 = ~n98958 & ~n98976;
  assign n99005 = ~n98984 & n99004;
  assign n99006 = n98964 & n98970;
  assign n99007 = n98984 & n98986;
  assign n99008 = ~n99006 & ~n99007;
  assign n99009 = ~n98958 & ~n99008;
  assign n99010 = ~n99005 & ~n99009;
  assign n99011 = n98964 & n98999;
  assign n99012 = ~n98984 & n99011;
  assign n99013 = n99010 & ~n99012;
  assign n99014 = ~n98976 & n99006;
  assign n99015 = n98984 & n99014;
  assign n99016 = n99013 & ~n99015;
  assign n99017 = ~n99003 & n99016;
  assign n99018 = pi8039 & pi9040;
  assign n99019 = pi8028 & ~pi9040;
  assign n99020 = ~n99018 & ~n99019;
  assign n99021 = ~pi8796 & ~n99020;
  assign n99022 = pi8796 & n99020;
  assign n99023 = ~n99021 & ~n99022;
  assign n99024 = ~n99017 & ~n99023;
  assign n99025 = ~n98964 & ~n98976;
  assign n99026 = ~n98958 & n98984;
  assign n99027 = n99023 & n99026;
  assign n99028 = n99025 & n99027;
  assign n99029 = ~n98964 & ~n98984;
  assign n99030 = n98976 & n99029;
  assign n99031 = ~n98958 & ~n99030;
  assign n99032 = ~n98970 & n98990;
  assign n99033 = ~n98977 & ~n99025;
  assign n99034 = ~n98984 & ~n99033;
  assign n99035 = n98964 & n98986;
  assign n99036 = n98958 & ~n99035;
  assign n99037 = ~n99034 & n99036;
  assign n99038 = ~n99032 & n99037;
  assign n99039 = ~n99031 & ~n99038;
  assign n99040 = n98964 & n98993;
  assign n99041 = n98984 & n99040;
  assign n99042 = ~n99039 & ~n99041;
  assign n99043 = n99023 & ~n99042;
  assign n99044 = ~n99028 & ~n99043;
  assign n99045 = ~n99024 & n99044;
  assign n99046 = ~n98998 & n99045;
  assign n99047 = ~n98958 & ~n98984;
  assign n99048 = n98999 & n99047;
  assign n99049 = n98964 & n99048;
  assign n99050 = n99046 & ~n99049;
  assign n99051 = pi8749 & ~n99050;
  assign n99052 = ~pi8749 & ~n99049;
  assign n99053 = n99045 & n99052;
  assign n99054 = ~n98998 & n99053;
  assign po5705 = n99051 | n99054;
  assign n99056 = pi8001 & ~pi9040;
  assign n99057 = pi7999 & pi9040;
  assign n99058 = ~n99056 & ~n99057;
  assign n99059 = ~pi8752 & ~n99058;
  assign n99060 = pi8752 & n99058;
  assign n99061 = ~n99059 & ~n99060;
  assign n99062 = pi7997 & pi9040;
  assign n99063 = pi7966 & ~pi9040;
  assign n99064 = ~n99062 & ~n99063;
  assign n99065 = ~pi8781 & ~n99064;
  assign n99066 = pi8781 & n99064;
  assign n99067 = ~n99065 & ~n99066;
  assign n99068 = pi8003 & ~pi9040;
  assign n99069 = pi8004 & pi9040;
  assign n99070 = ~n99068 & ~n99069;
  assign n99071 = ~pi8799 & n99070;
  assign n99072 = pi8799 & ~n99070;
  assign n99073 = ~n99071 & ~n99072;
  assign n99074 = pi7961 & ~pi9040;
  assign n99075 = pi8013 & pi9040;
  assign n99076 = ~n99074 & ~n99075;
  assign n99077 = pi8702 & n99076;
  assign n99078 = ~pi8702 & ~n99076;
  assign n99079 = ~n99077 & ~n99078;
  assign n99080 = ~n99073 & ~n99079;
  assign n99081 = ~n99067 & n99080;
  assign n99082 = n99061 & n99081;
  assign n99083 = pi7968 & pi9040;
  assign n99084 = pi7978 & ~pi9040;
  assign n99085 = ~n99083 & ~n99084;
  assign n99086 = ~pi8742 & n99085;
  assign n99087 = pi8742 & ~n99085;
  assign n99088 = ~n99086 & ~n99087;
  assign n99089 = pi7943 & ~pi9040;
  assign n99090 = pi7957 & pi9040;
  assign n99091 = ~n99089 & ~n99090;
  assign n99092 = ~pi8803 & ~n99091;
  assign n99093 = pi8803 & n99091;
  assign n99094 = ~n99092 & ~n99093;
  assign n99095 = n99067 & ~n99094;
  assign n99096 = n99079 & n99095;
  assign n99097 = n99073 & n99096;
  assign n99098 = ~n99061 & n99094;
  assign n99099 = n99067 & n99098;
  assign n99100 = ~n99073 & n99099;
  assign n99101 = ~n99097 & ~n99100;
  assign n99102 = ~n99061 & ~n99067;
  assign n99103 = ~n99079 & n99102;
  assign n99104 = n99073 & n99103;
  assign n99105 = n99067 & ~n99073;
  assign n99106 = ~n99061 & n99105;
  assign n99107 = n99061 & ~n99094;
  assign n99108 = ~n99067 & n99107;
  assign n99109 = ~n99106 & ~n99108;
  assign n99110 = ~n99079 & ~n99109;
  assign n99111 = ~n99104 & ~n99110;
  assign n99112 = n99101 & n99111;
  assign n99113 = n99088 & ~n99112;
  assign n99114 = ~n99067 & n99098;
  assign n99115 = n99073 & n99114;
  assign n99116 = n99061 & n99095;
  assign n99117 = ~n99073 & n99116;
  assign n99118 = ~n99061 & ~n99094;
  assign n99119 = ~n99067 & n99118;
  assign n99120 = ~n99073 & n99119;
  assign n99121 = ~n99117 & ~n99120;
  assign n99122 = ~n99115 & n99121;
  assign n99123 = n99079 & ~n99122;
  assign n99124 = n99061 & n99073;
  assign n99125 = n99067 & n99124;
  assign n99126 = n99094 & n99125;
  assign n99127 = ~n99123 & ~n99126;
  assign n99128 = ~n99113 & n99127;
  assign n99129 = n99067 & n99073;
  assign n99130 = ~n99061 & n99129;
  assign n99131 = n99061 & n99094;
  assign n99132 = ~n99067 & n99131;
  assign n99133 = ~n99130 & ~n99132;
  assign n99134 = ~n99079 & ~n99133;
  assign n99135 = n99094 & n99129;
  assign n99136 = ~n99134 & ~n99135;
  assign n99137 = n99067 & n99131;
  assign n99138 = ~n99067 & n99073;
  assign n99139 = ~n99094 & n99138;
  assign n99140 = ~n99073 & n99118;
  assign n99141 = ~n99139 & ~n99140;
  assign n99142 = ~n99102 & n99141;
  assign n99143 = ~n99137 & n99142;
  assign n99144 = n99079 & ~n99143;
  assign n99145 = n99136 & ~n99144;
  assign n99146 = ~n99117 & n99145;
  assign n99147 = ~n99088 & ~n99146;
  assign n99148 = n99128 & ~n99147;
  assign n99149 = ~n99082 & n99148;
  assign n99150 = ~pi8697 & ~n99149;
  assign n99151 = ~n99126 & ~n99147;
  assign n99152 = ~n99123 & n99151;
  assign n99153 = ~n99113 & n99152;
  assign n99154 = ~n99082 & n99153;
  assign n99155 = pi8697 & n99154;
  assign po5742 = n99150 | n99155;
  assign n99157 = pi7979 & ~pi9040;
  assign n99158 = pi8017 & pi9040;
  assign n99159 = ~n99157 & ~n99158;
  assign n99160 = ~pi8717 & n99159;
  assign n99161 = pi8717 & ~n99159;
  assign n99162 = ~n99160 & ~n99161;
  assign n99163 = pi7946 & ~pi9040;
  assign n99164 = pi7942 & pi9040;
  assign n99165 = ~n99163 & ~n99164;
  assign n99166 = pi8748 & n99165;
  assign n99167 = ~pi8748 & ~n99165;
  assign n99168 = ~n99166 & ~n99167;
  assign n99169 = pi8038 & pi9040;
  assign n99170 = pi8033 & ~pi9040;
  assign n99171 = ~n99169 & ~n99170;
  assign n99172 = pi8802 & n99171;
  assign n99173 = ~pi8802 & ~n99171;
  assign n99174 = ~n99172 & ~n99173;
  assign n99175 = pi8011 & ~pi9040;
  assign n99176 = pi7966 & pi9040;
  assign n99177 = ~n99175 & ~n99176;
  assign n99178 = ~pi8705 & n99177;
  assign n99179 = pi8705 & ~n99177;
  assign n99180 = ~n99178 & ~n99179;
  assign n99181 = n99174 & ~n99180;
  assign n99182 = ~n99168 & n99181;
  assign n99183 = n99162 & n99182;
  assign n99184 = n99174 & n99180;
  assign n99185 = ~n99168 & n99184;
  assign n99186 = ~n99162 & n99185;
  assign n99187 = pi7943 & pi9040;
  assign n99188 = pi8039 & ~pi9040;
  assign n99189 = ~n99187 & ~n99188;
  assign n99190 = pi8710 & ~n99189;
  assign n99191 = ~pi8710 & n99189;
  assign n99192 = ~n99190 & ~n99191;
  assign n99193 = n99162 & ~n99168;
  assign n99194 = n99180 & n99193;
  assign n99195 = ~n99174 & n99194;
  assign n99196 = n99168 & n99174;
  assign n99197 = ~n99195 & ~n99196;
  assign n99198 = ~n99192 & ~n99197;
  assign n99199 = ~n99186 & ~n99198;
  assign n99200 = ~n99183 & n99199;
  assign n99201 = ~n99174 & n99180;
  assign n99202 = n99168 & n99201;
  assign n99203 = ~n99162 & n99202;
  assign n99204 = ~n99174 & ~n99180;
  assign n99205 = n99168 & n99204;
  assign n99206 = n99162 & n99205;
  assign n99207 = ~n99168 & n99204;
  assign n99208 = ~n99162 & n99207;
  assign n99209 = n99192 & n99208;
  assign n99210 = ~n99206 & ~n99209;
  assign n99211 = ~n99203 & n99210;
  assign n99212 = n99200 & n99211;
  assign n99213 = pi7958 & pi9040;
  assign n99214 = pi7937 & ~pi9040;
  assign n99215 = ~n99213 & ~n99214;
  assign n99216 = ~pi8712 & ~n99215;
  assign n99217 = pi8712 & n99215;
  assign n99218 = ~n99216 & ~n99217;
  assign n99219 = ~n99212 & n99218;
  assign n99220 = n99162 & n99202;
  assign n99221 = ~n99192 & n99207;
  assign n99222 = ~n99162 & n99182;
  assign n99223 = ~n99162 & n99205;
  assign n99224 = ~n99162 & ~n99168;
  assign n99225 = n99180 & n99224;
  assign n99226 = ~n99174 & n99225;
  assign n99227 = ~n99223 & ~n99226;
  assign n99228 = ~n99222 & n99227;
  assign n99229 = ~n99221 & n99228;
  assign n99230 = n99168 & ~n99180;
  assign n99231 = ~n99162 & n99174;
  assign n99232 = ~n99230 & ~n99231;
  assign n99233 = ~n99168 & n99180;
  assign n99234 = n99232 & ~n99233;
  assign n99235 = n99192 & ~n99234;
  assign n99236 = n99229 & ~n99235;
  assign n99237 = n99174 & n99194;
  assign n99238 = n99236 & ~n99237;
  assign n99239 = ~n99220 & n99238;
  assign n99240 = ~n99218 & ~n99239;
  assign n99241 = ~n99219 & ~n99240;
  assign n99242 = pi8788 & ~n99241;
  assign n99243 = ~pi8788 & ~n99219;
  assign n99244 = ~n99240 & n99243;
  assign po5764 = n99242 | n99244;
  assign n99246 = n99192 & n99204;
  assign n99247 = n99162 & n99246;
  assign n99248 = n99168 & n99184;
  assign n99249 = ~n99226 & ~n99248;
  assign n99250 = ~n99162 & n99181;
  assign n99251 = n99249 & ~n99250;
  assign n99252 = n99192 & ~n99251;
  assign n99253 = ~n99168 & n99174;
  assign n99254 = n99162 & ~n99192;
  assign n99255 = n99253 & n99254;
  assign n99256 = ~n99237 & ~n99255;
  assign n99257 = ~n99252 & n99256;
  assign n99258 = ~n99247 & n99257;
  assign n99259 = n99168 & n99181;
  assign n99260 = ~n99162 & n99259;
  assign n99261 = ~n99206 & ~n99260;
  assign n99262 = n99258 & n99261;
  assign n99263 = ~n99218 & ~n99262;
  assign n99264 = ~n99183 & ~n99205;
  assign n99265 = n99192 & ~n99264;
  assign n99266 = ~n99195 & ~n99208;
  assign n99267 = n99174 & n99224;
  assign n99268 = n99162 & n99168;
  assign n99269 = ~n99180 & n99268;
  assign n99270 = n99174 & n99269;
  assign n99271 = ~n99267 & ~n99270;
  assign n99272 = ~n99192 & ~n99271;
  assign n99273 = n99266 & ~n99272;
  assign n99274 = ~n99265 & n99273;
  assign n99275 = n99218 & ~n99274;
  assign n99276 = ~n99162 & n99196;
  assign n99277 = n99168 & ~n99174;
  assign n99278 = n99162 & n99277;
  assign n99279 = ~n99276 & ~n99278;
  assign n99280 = n99192 & ~n99279;
  assign n99281 = ~n99203 & ~n99208;
  assign n99282 = ~n99185 & n99281;
  assign n99283 = ~n99192 & ~n99282;
  assign n99284 = ~n99280 & ~n99283;
  assign n99285 = ~n99192 & n99233;
  assign n99286 = n99162 & n99285;
  assign n99287 = n99284 & ~n99286;
  assign n99288 = ~n99275 & n99287;
  assign n99289 = ~n99263 & n99288;
  assign n99290 = ~pi8709 & ~n99289;
  assign n99291 = pi8709 & n99289;
  assign po5780 = n99290 | n99291;
  assign n99293 = pi8036 & ~pi9040;
  assign n99294 = pi7949 & pi9040;
  assign n99295 = ~n99293 & ~n99294;
  assign n99296 = pi8772 & n99295;
  assign n99297 = ~pi8772 & ~n99295;
  assign n99298 = ~n99296 & ~n99297;
  assign n99299 = pi8023 & ~pi9040;
  assign n99300 = pi7959 & pi9040;
  assign n99301 = ~n99299 & ~n99300;
  assign n99302 = pi8778 & n99301;
  assign n99303 = ~pi8778 & ~n99301;
  assign n99304 = ~n99302 & ~n99303;
  assign n99305 = pi8025 & ~pi9040;
  assign n99306 = pi7971 & pi9040;
  assign n99307 = ~n99305 & ~n99306;
  assign n99308 = ~pi8773 & n99307;
  assign n99309 = pi8773 & ~n99307;
  assign n99310 = ~n99308 & ~n99309;
  assign n99311 = pi8010 & pi9040;
  assign n99312 = pi7972 & ~pi9040;
  assign n99313 = ~n99311 & ~n99312;
  assign n99314 = ~pi8775 & ~n99313;
  assign n99315 = pi8775 & n99313;
  assign n99316 = ~n99314 & ~n99315;
  assign n99317 = pi8022 & ~pi9040;
  assign n99318 = pi7998 & pi9040;
  assign n99319 = ~n99317 & ~n99318;
  assign n99320 = pi8781 & n99319;
  assign n99321 = ~pi8781 & ~n99319;
  assign n99322 = ~n99320 & ~n99321;
  assign n99323 = n99316 & ~n99322;
  assign n99324 = n99310 & n99323;
  assign n99325 = n99304 & n99324;
  assign n99326 = ~n99316 & ~n99322;
  assign n99327 = n99310 & n99326;
  assign n99328 = ~n99304 & n99327;
  assign n99329 = ~n99325 & ~n99328;
  assign n99330 = n99298 & ~n99329;
  assign n99331 = ~n99304 & ~n99310;
  assign n99332 = n99322 & n99331;
  assign n99333 = ~n99316 & n99332;
  assign n99334 = ~n99298 & n99333;
  assign n99335 = pi7963 & pi9040;
  assign n99336 = pi7952 & ~pi9040;
  assign n99337 = ~n99335 & ~n99336;
  assign n99338 = ~pi8752 & ~n99337;
  assign n99339 = pi8752 & n99337;
  assign n99340 = ~n99338 & ~n99339;
  assign n99341 = ~n99310 & n99323;
  assign n99342 = n99298 & n99341;
  assign n99343 = ~n99333 & ~n99342;
  assign n99344 = ~n99304 & n99316;
  assign n99345 = n99310 & n99344;
  assign n99346 = ~n99316 & n99331;
  assign n99347 = ~n99345 & ~n99346;
  assign n99348 = ~n99298 & ~n99347;
  assign n99349 = ~n99298 & n99304;
  assign n99350 = n99326 & n99349;
  assign n99351 = n99310 & n99350;
  assign n99352 = n99316 & n99322;
  assign n99353 = ~n99310 & n99352;
  assign n99354 = n99304 & n99353;
  assign n99355 = n99298 & n99310;
  assign n99356 = n99322 & n99355;
  assign n99357 = ~n99316 & n99356;
  assign n99358 = ~n99354 & ~n99357;
  assign n99359 = ~n99351 & n99358;
  assign n99360 = ~n99348 & n99359;
  assign n99361 = n99343 & n99360;
  assign n99362 = n99340 & ~n99361;
  assign n99363 = ~n99304 & n99342;
  assign n99364 = ~n99362 & ~n99363;
  assign n99365 = ~n99334 & n99364;
  assign n99366 = ~n99330 & n99365;
  assign n99367 = n99304 & n99323;
  assign n99368 = n99310 & n99322;
  assign n99369 = ~n99367 & ~n99368;
  assign n99370 = ~n99298 & ~n99369;
  assign n99371 = n99298 & n99304;
  assign n99372 = ~n99310 & ~n99316;
  assign n99373 = n99371 & n99372;
  assign n99374 = n99298 & n99327;
  assign n99375 = ~n99373 & ~n99374;
  assign n99376 = n99310 & n99352;
  assign n99377 = ~n99304 & n99376;
  assign n99378 = n99298 & n99353;
  assign n99379 = ~n99377 & ~n99378;
  assign n99380 = n99375 & n99379;
  assign n99381 = ~n99370 & n99380;
  assign n99382 = n99304 & ~n99310;
  assign n99383 = ~n99322 & n99382;
  assign n99384 = ~n99316 & n99383;
  assign n99385 = n99381 & ~n99384;
  assign n99386 = ~n99328 & n99385;
  assign n99387 = ~n99340 & ~n99386;
  assign n99388 = n99366 & ~n99387;
  assign n99389 = ~pi8695 & ~n99388;
  assign n99390 = pi8695 & n99366;
  assign n99391 = ~n99387 & n99390;
  assign po5815 = n99389 | n99391;
  assign n99393 = n99073 & n99116;
  assign n99394 = ~n99120 & ~n99393;
  assign n99395 = n99079 & ~n99394;
  assign n99396 = ~n99061 & n99067;
  assign n99397 = ~n99094 & n99396;
  assign n99398 = ~n99073 & n99397;
  assign n99399 = ~n99073 & n99114;
  assign n99400 = ~n99398 & ~n99399;
  assign n99401 = ~n99079 & ~n99400;
  assign n99402 = ~n99395 & ~n99401;
  assign n99403 = n99073 & n99397;
  assign n99404 = ~n99114 & ~n99126;
  assign n99405 = ~n99073 & n99095;
  assign n99406 = n99073 & n99108;
  assign n99407 = ~n99405 & ~n99406;
  assign n99408 = n99404 & n99407;
  assign n99409 = ~n99079 & ~n99408;
  assign n99410 = ~n99073 & n99132;
  assign n99411 = ~n99073 & n99131;
  assign n99412 = ~n99130 & ~n99411;
  assign n99413 = ~n99119 & n99412;
  assign n99414 = n99079 & ~n99413;
  assign n99415 = ~n99410 & ~n99414;
  assign n99416 = ~n99409 & n99415;
  assign n99417 = ~n99403 & n99416;
  assign n99418 = n99088 & ~n99417;
  assign n99419 = n99080 & n99137;
  assign n99420 = ~n99079 & n99119;
  assign n99421 = ~n99079 & n99099;
  assign n99422 = ~n99420 & ~n99421;
  assign n99423 = n99073 & ~n99422;
  assign n99424 = ~n99419 & ~n99423;
  assign n99425 = ~n99073 & n99108;
  assign n99426 = ~n99393 & ~n99425;
  assign n99427 = ~n99073 & n99098;
  assign n99428 = n99073 & n99131;
  assign n99429 = ~n99427 & ~n99428;
  assign n99430 = ~n99116 & n99429;
  assign n99431 = ~n99114 & n99430;
  assign n99432 = n99079 & ~n99431;
  assign n99433 = n99073 & n99132;
  assign n99434 = ~n99432 & ~n99433;
  assign n99435 = n99426 & n99434;
  assign n99436 = n99424 & n99435;
  assign n99437 = ~n99088 & ~n99436;
  assign n99438 = ~n99418 & ~n99437;
  assign n99439 = n99402 & n99438;
  assign n99440 = pi8793 & ~n99439;
  assign n99441 = ~pi8793 & n99439;
  assign po5816 = n99440 | n99441;
  assign n99443 = n99073 & ~n99079;
  assign n99444 = n99061 & n99443;
  assign n99445 = ~n99061 & n99139;
  assign n99446 = ~n99132 & ~n99445;
  assign n99447 = n99079 & ~n99446;
  assign n99448 = n99400 & ~n99447;
  assign n99449 = ~n99444 & n99448;
  assign n99450 = ~n99088 & ~n99449;
  assign n99451 = ~n99079 & n99425;
  assign n99452 = n99073 & n99079;
  assign n99453 = n99108 & n99452;
  assign n99454 = ~n99130 & ~n99453;
  assign n99455 = ~n99099 & ~n99132;
  assign n99456 = n99073 & n99098;
  assign n99457 = n99455 & ~n99456;
  assign n99458 = ~n99079 & ~n99457;
  assign n99459 = n99079 & n99137;
  assign n99460 = n99121 & ~n99459;
  assign n99461 = ~n99458 & n99460;
  assign n99462 = n99454 & n99461;
  assign n99463 = n99088 & ~n99462;
  assign n99464 = ~n99451 & ~n99463;
  assign n99465 = ~n99450 & n99464;
  assign n99466 = n99099 & n99452;
  assign n99467 = ~n99073 & n99096;
  assign n99468 = ~n99466 & ~n99467;
  assign n99469 = n99079 & n99399;
  assign n99470 = n99468 & ~n99469;
  assign n99471 = n99465 & n99470;
  assign n99472 = ~pi8744 & ~n99471;
  assign n99473 = pi8744 & n99470;
  assign n99474 = n99464 & n99473;
  assign n99475 = ~n99450 & n99474;
  assign po5817 = n99472 | n99475;
  assign n99477 = n99162 & n99181;
  assign n99478 = ~n99220 & ~n99477;
  assign n99479 = ~n99192 & n99478;
  assign n99480 = ~n99162 & n99277;
  assign n99481 = ~n99184 & ~n99204;
  assign n99482 = n99168 & ~n99481;
  assign n99483 = ~n99174 & n99193;
  assign n99484 = ~n99162 & n99184;
  assign n99485 = ~n99483 & ~n99484;
  assign n99486 = n99192 & n99485;
  assign n99487 = ~n99482 & n99486;
  assign n99488 = ~n99480 & n99487;
  assign n99489 = ~n99479 & ~n99488;
  assign n99490 = ~n99162 & n99482;
  assign n99491 = ~n99222 & ~n99490;
  assign n99492 = ~n99489 & n99491;
  assign n99493 = n99218 & ~n99492;
  assign n99494 = ~n99192 & ~n99481;
  assign n99495 = n99162 & n99494;
  assign n99496 = ~n99162 & n99201;
  assign n99497 = ~n99260 & ~n99496;
  assign n99498 = ~n99192 & ~n99497;
  assign n99499 = ~n99168 & n99494;
  assign n99500 = ~n99498 & ~n99499;
  assign n99501 = ~n99495 & n99500;
  assign n99502 = ~n99218 & ~n99501;
  assign n99503 = ~n99493 & ~n99502;
  assign n99504 = n99192 & ~n99478;
  assign n99505 = ~n99226 & ~n99504;
  assign n99506 = ~n99218 & ~n99505;
  assign n99507 = ~n99192 & n99226;
  assign n99508 = n99192 & ~n99491;
  assign n99509 = ~n99507 & ~n99508;
  assign n99510 = ~n99506 & n99509;
  assign n99511 = n99503 & n99510;
  assign n99512 = pi8718 & ~n99511;
  assign n99513 = ~pi8718 & n99510;
  assign n99514 = ~n99502 & n99513;
  assign n99515 = ~n99493 & n99514;
  assign po5828 = n99512 | n99515;
  assign n99517 = pi7971 & ~pi9040;
  assign n99518 = pi8000 & pi9040;
  assign n99519 = ~n99517 & ~n99518;
  assign n99520 = pi8726 & n99519;
  assign n99521 = ~pi8726 & ~n99519;
  assign n99522 = ~n99520 & ~n99521;
  assign n99523 = pi7986 & ~pi9040;
  assign n99524 = pi8022 & pi9040;
  assign n99525 = ~n99523 & ~n99524;
  assign n99526 = ~pi8776 & n99525;
  assign n99527 = pi8776 & ~n99525;
  assign n99528 = ~n99526 & ~n99527;
  assign n99529 = pi7975 & ~pi9040;
  assign n99530 = pi8030 & pi9040;
  assign n99531 = ~n99529 & ~n99530;
  assign n99532 = ~pi8750 & n99531;
  assign n99533 = pi8750 & ~n99531;
  assign n99534 = ~n99532 & ~n99533;
  assign n99535 = pi8010 & ~pi9040;
  assign n99536 = pi8005 & pi9040;
  assign n99537 = ~n99535 & ~n99536;
  assign n99538 = pi8743 & n99537;
  assign n99539 = ~pi8743 & ~n99537;
  assign n99540 = ~n99538 & ~n99539;
  assign n99541 = pi8016 & ~pi9040;
  assign n99542 = pi8023 & pi9040;
  assign n99543 = ~n99541 & ~n99542;
  assign n99544 = pi8761 & n99543;
  assign n99545 = ~pi8761 & ~n99543;
  assign n99546 = ~n99544 & ~n99545;
  assign n99547 = n99540 & n99546;
  assign n99548 = n99534 & n99547;
  assign n99549 = ~n99528 & n99548;
  assign n99550 = n99540 & ~n99546;
  assign n99551 = n99528 & n99550;
  assign n99552 = ~n99549 & ~n99551;
  assign n99553 = ~n99522 & ~n99552;
  assign n99554 = pi8036 & pi9040;
  assign n99555 = pi8007 & ~pi9040;
  assign n99556 = ~n99554 & ~n99555;
  assign n99557 = pi8713 & n99556;
  assign n99558 = ~pi8713 & ~n99556;
  assign n99559 = ~n99557 & ~n99558;
  assign n99560 = n99522 & ~n99540;
  assign n99561 = ~n99528 & n99560;
  assign n99562 = ~n99528 & n99534;
  assign n99563 = ~n99546 & n99562;
  assign n99564 = ~n99528 & ~n99534;
  assign n99565 = n99546 & n99564;
  assign n99566 = ~n99563 & ~n99565;
  assign n99567 = n99528 & n99534;
  assign n99568 = n99546 & n99567;
  assign n99569 = n99540 & n99568;
  assign n99570 = n99566 & ~n99569;
  assign n99571 = n99522 & ~n99570;
  assign n99572 = ~n99561 & ~n99571;
  assign n99573 = n99528 & ~n99534;
  assign n99574 = ~n99546 & n99573;
  assign n99575 = n99540 & n99574;
  assign n99576 = n99572 & ~n99575;
  assign n99577 = ~n99540 & n99567;
  assign n99578 = n99528 & n99546;
  assign n99579 = ~n99534 & n99578;
  assign n99580 = ~n99577 & ~n99579;
  assign n99581 = ~n99522 & ~n99580;
  assign n99582 = ~n99546 & n99564;
  assign n99583 = ~n99540 & n99582;
  assign n99584 = ~n99581 & ~n99583;
  assign n99585 = n99576 & n99584;
  assign n99586 = n99559 & ~n99585;
  assign n99587 = ~n99553 & ~n99586;
  assign n99588 = n99522 & ~n99559;
  assign n99589 = ~n99580 & n99588;
  assign n99590 = ~n99546 & n99567;
  assign n99591 = ~n99582 & ~n99590;
  assign n99592 = n99540 & ~n99591;
  assign n99593 = ~n99549 & ~n99592;
  assign n99594 = ~n99559 & ~n99593;
  assign n99595 = ~n99589 & ~n99594;
  assign n99596 = ~n99522 & ~n99559;
  assign n99597 = ~n99540 & n99562;
  assign n99598 = ~n99574 & ~n99597;
  assign n99599 = ~n99528 & n99546;
  assign n99600 = n99598 & ~n99599;
  assign n99601 = n99596 & ~n99600;
  assign n99602 = n99595 & ~n99601;
  assign n99603 = n99587 & n99602;
  assign n99604 = ~pi8771 & ~n99603;
  assign n99605 = pi8771 & n99595;
  assign n99606 = n99587 & n99605;
  assign n99607 = ~n99601 & n99606;
  assign po5837 = n99604 | n99607;
  assign n99609 = ~n99316 & n99322;
  assign n99610 = n99298 & n99609;
  assign n99611 = ~n99304 & n99610;
  assign n99612 = n99304 & n99310;
  assign n99613 = n99316 & n99612;
  assign n99614 = ~n99324 & ~n99613;
  assign n99615 = n99298 & ~n99614;
  assign n99616 = ~n99611 & ~n99615;
  assign n99617 = ~n99298 & n99352;
  assign n99618 = ~n99304 & n99617;
  assign n99619 = ~n99298 & n99327;
  assign n99620 = ~n99618 & ~n99619;
  assign n99621 = n99616 & n99620;
  assign n99622 = n99316 & n99331;
  assign n99623 = ~n99328 & ~n99622;
  assign n99624 = ~n99384 & n99623;
  assign n99625 = n99621 & n99624;
  assign n99626 = ~n99340 & ~n99625;
  assign n99627 = ~n99324 & ~n99333;
  assign n99628 = ~n99367 & n99627;
  assign n99629 = ~n99298 & ~n99628;
  assign n99630 = n99310 & n99609;
  assign n99631 = n99304 & n99630;
  assign n99632 = ~n99354 & ~n99631;
  assign n99633 = n99298 & n99377;
  assign n99634 = n99632 & ~n99633;
  assign n99635 = ~n99310 & n99326;
  assign n99636 = n99298 & n99635;
  assign n99637 = n99634 & ~n99636;
  assign n99638 = ~n99629 & n99637;
  assign n99639 = n99340 & ~n99638;
  assign n99640 = ~n99363 & ~n99373;
  assign n99641 = ~n99328 & n99632;
  assign n99642 = ~n99298 & ~n99641;
  assign n99643 = n99640 & ~n99642;
  assign n99644 = ~n99639 & n99643;
  assign n99645 = ~n99626 & n99644;
  assign n99646 = pi8722 & ~n99645;
  assign n99647 = ~pi8722 & n99645;
  assign po5880 = n99646 | n99647;
  assign n99649 = n99304 & n99341;
  assign n99650 = ~n99304 & n99635;
  assign n99651 = ~n99649 & ~n99650;
  assign n99652 = ~n99310 & n99609;
  assign n99653 = n99304 & n99652;
  assign n99654 = n99304 & n99352;
  assign n99655 = ~n99304 & n99630;
  assign n99656 = ~n99654 & ~n99655;
  assign n99657 = ~n99298 & ~n99656;
  assign n99658 = ~n99653 & ~n99657;
  assign n99659 = n99304 & n99610;
  assign n99660 = ~n99374 & ~n99659;
  assign n99661 = n99658 & n99660;
  assign n99662 = n99651 & n99661;
  assign n99663 = n99340 & ~n99662;
  assign n99664 = ~n99298 & ~n99340;
  assign n99665 = ~n99316 & n99612;
  assign n99666 = n99310 & ~n99322;
  assign n99667 = ~n99665 & ~n99666;
  assign n99668 = n99664 & ~n99667;
  assign n99669 = ~n99333 & ~n99345;
  assign n99670 = ~n99310 & ~n99609;
  assign n99671 = n99371 & n99670;
  assign n99672 = ~n99342 & ~n99671;
  assign n99673 = n99669 & n99672;
  assign n99674 = ~n99340 & ~n99673;
  assign n99675 = ~n99298 & n99324;
  assign n99676 = ~n99304 & n99675;
  assign n99677 = ~n99304 & n99353;
  assign n99678 = ~n99650 & ~n99677;
  assign n99679 = ~n99298 & ~n99678;
  assign n99680 = ~n99676 & ~n99679;
  assign n99681 = n99298 & n99333;
  assign n99682 = n99680 & ~n99681;
  assign n99683 = ~n99674 & n99682;
  assign n99684 = ~n99668 & n99683;
  assign n99685 = ~n99663 & n99684;
  assign n99686 = ~n99633 & n99685;
  assign n99687 = ~pi8701 & ~n99686;
  assign n99688 = pi8701 & ~n99633;
  assign n99689 = n99684 & n99688;
  assign n99690 = ~n99663 & n99689;
  assign po5888 = n99687 | n99690;
  assign n99692 = n98708 & ~n98720;
  assign n99693 = n98702 & n99692;
  assign n99694 = ~n98835 & ~n99693;
  assign n99695 = n98714 & n98745;
  assign n99696 = n98720 & n99695;
  assign n99697 = n98720 & ~n98729;
  assign n99698 = ~n98817 & ~n99697;
  assign n99699 = ~n98714 & ~n99698;
  assign n99700 = ~n99696 & ~n99699;
  assign n99701 = n99694 & n99700;
  assign n99702 = n98739 & ~n99701;
  assign n99703 = ~n98741 & ~n98783;
  assign n99704 = n98720 & n98760;
  assign n99705 = n99703 & ~n99704;
  assign n99706 = n98714 & ~n99705;
  assign n99707 = n98745 & n98776;
  assign n99708 = ~n98732 & ~n99707;
  assign n99709 = ~n99706 & n99708;
  assign n99710 = ~n98753 & ~n98762;
  assign n99711 = ~n98714 & ~n99710;
  assign n99712 = n99709 & ~n99711;
  assign n99713 = ~n98739 & ~n99712;
  assign n99714 = ~n99702 & ~n99713;
  assign n99715 = ~n98720 & n98757;
  assign n99716 = n98720 & ~n98752;
  assign n99717 = ~n99715 & ~n99716;
  assign n99718 = ~n98714 & n99717;
  assign n99719 = n98714 & ~n98720;
  assign n99720 = ~n98768 & ~n98771;
  assign n99721 = ~n98741 & n99720;
  assign n99722 = n99719 & ~n99721;
  assign n99723 = ~n99718 & ~n99722;
  assign n99724 = n99714 & n99723;
  assign n99725 = ~pi8790 & ~n99724;
  assign n99726 = pi8790 & n99723;
  assign n99727 = ~n99713 & n99726;
  assign n99728 = ~n99702 & n99727;
  assign po5904 = n99725 | n99728;
  assign n99730 = ~n98985 & ~n98992;
  assign n99731 = ~n98958 & ~n99730;
  assign n99732 = ~n99049 & ~n99731;
  assign n99733 = ~n98964 & ~n98970;
  assign n99734 = n98958 & n99733;
  assign n99735 = n98984 & n99734;
  assign n99736 = n98984 & n98999;
  assign n99737 = ~n99733 & ~n99736;
  assign n99738 = n98964 & ~n98984;
  assign n99739 = n98970 & n99738;
  assign n99740 = n99737 & ~n99739;
  assign n99741 = n98958 & ~n99740;
  assign n99742 = ~n98995 & ~n99741;
  assign n99743 = ~n99023 & ~n99742;
  assign n99744 = ~n98958 & n98977;
  assign n99745 = n98984 & n99744;
  assign n99746 = ~n98958 & n99035;
  assign n99747 = ~n99745 & ~n99746;
  assign n99748 = ~n99023 & ~n99747;
  assign n99749 = ~n99743 & ~n99748;
  assign n99750 = ~n99735 & n99749;
  assign n99751 = n98970 & n99029;
  assign n99752 = ~n99011 & ~n99030;
  assign n99753 = ~n99040 & n99752;
  assign n99754 = ~n98958 & ~n99753;
  assign n99755 = n98976 & n99738;
  assign n99756 = ~n98970 & n99755;
  assign n99757 = ~n99014 & ~n99756;
  assign n99758 = n98958 & ~n99757;
  assign n99759 = ~n99754 & ~n99758;
  assign n99760 = ~n99751 & n99759;
  assign n99761 = ~n99001 & ~n99041;
  assign n99762 = n99760 & n99761;
  assign n99763 = n99023 & ~n99762;
  assign n99764 = n99750 & ~n99763;
  assign n99765 = n99732 & n99764;
  assign n99766 = ~pi8755 & ~n99765;
  assign n99767 = pi8755 & n99750;
  assign n99768 = n99732 & n99767;
  assign n99769 = ~n99763 & n99768;
  assign po5914 = n99766 | n99769;
  assign n99771 = pi7939 & ~pi9040;
  assign n99772 = pi8025 & pi9040;
  assign n99773 = ~n99771 & ~n99772;
  assign n99774 = pi8773 & n99773;
  assign n99775 = ~pi8773 & ~n99773;
  assign n99776 = ~n99774 & ~n99775;
  assign n99777 = pi7963 & ~pi9040;
  assign n99778 = pi8034 & pi9040;
  assign n99779 = ~n99777 & ~n99778;
  assign n99780 = ~pi8782 & n99779;
  assign n99781 = pi8782 & ~n99779;
  assign n99782 = ~n99780 & ~n99781;
  assign n99783 = pi7949 & ~pi9040;
  assign n99784 = pi8031 & pi9040;
  assign n99785 = ~n99783 & ~n99784;
  assign n99786 = ~pi8750 & n99785;
  assign n99787 = pi8750 & ~n99785;
  assign n99788 = ~n99786 & ~n99787;
  assign n99789 = n99782 & ~n99788;
  assign n99790 = n99776 & n99789;
  assign n99791 = pi7929 & ~pi9040;
  assign n99792 = pi8020 & pi9040;
  assign n99793 = ~n99791 & ~n99792;
  assign n99794 = pi8713 & n99793;
  assign n99795 = ~pi8713 & ~n99793;
  assign n99796 = ~n99794 & ~n99795;
  assign n99797 = n99776 & n99796;
  assign n99798 = ~n99788 & n99797;
  assign n99799 = ~n99776 & n99796;
  assign n99800 = n99788 & n99799;
  assign n99801 = ~n99798 & ~n99800;
  assign n99802 = ~n99790 & n99801;
  assign n99803 = pi7931 & ~pi9040;
  assign n99804 = pi7986 & pi9040;
  assign n99805 = ~n99803 & ~n99804;
  assign n99806 = ~pi8795 & n99805;
  assign n99807 = pi8795 & ~n99805;
  assign n99808 = ~n99806 & ~n99807;
  assign n99809 = pi7977 & pi9040;
  assign n99810 = pi7959 & ~pi9040;
  assign n99811 = ~n99809 & ~n99810;
  assign n99812 = ~pi8775 & n99811;
  assign n99813 = pi8775 & ~n99811;
  assign n99814 = ~n99812 & ~n99813;
  assign n99815 = n99808 & ~n99814;
  assign n99816 = ~n99802 & n99815;
  assign n99817 = ~n99776 & ~n99796;
  assign n99818 = ~n99788 & n99817;
  assign n99819 = ~n99782 & ~n99814;
  assign n99820 = n99818 & n99819;
  assign n99821 = ~n99788 & n99799;
  assign n99822 = ~n99808 & n99821;
  assign n99823 = n99776 & ~n99796;
  assign n99824 = ~n99782 & n99823;
  assign n99825 = n99776 & n99788;
  assign n99826 = ~n99824 & ~n99825;
  assign n99827 = ~n99808 & ~n99826;
  assign n99828 = ~n99822 & ~n99827;
  assign n99829 = ~n99814 & ~n99828;
  assign n99830 = ~n99820 & ~n99829;
  assign n99831 = ~n99782 & n99788;
  assign n99832 = n99776 & n99831;
  assign n99833 = n99782 & n99817;
  assign n99834 = n99788 & n99833;
  assign n99835 = ~n99832 & ~n99834;
  assign n99836 = ~n99808 & ~n99835;
  assign n99837 = n99830 & ~n99836;
  assign n99838 = ~n99782 & n99808;
  assign n99839 = n99823 & n99838;
  assign n99840 = ~n99788 & n99839;
  assign n99841 = ~n99797 & ~n99817;
  assign n99842 = n99789 & ~n99841;
  assign n99843 = n99782 & n99788;
  assign n99844 = ~n99776 & n99843;
  assign n99845 = n99796 & n99844;
  assign n99846 = ~n99842 & ~n99845;
  assign n99847 = n99788 & n99823;
  assign n99848 = n99782 & n99808;
  assign n99849 = n99847 & n99848;
  assign n99850 = n99831 & ~n99841;
  assign n99851 = ~n99782 & n99821;
  assign n99852 = ~n99850 & ~n99851;
  assign n99853 = ~n99849 & n99852;
  assign n99854 = n99846 & n99853;
  assign n99855 = ~n99840 & n99854;
  assign n99856 = n99782 & ~n99808;
  assign n99857 = ~n99788 & n99856;
  assign n99858 = ~n99796 & n99857;
  assign n99859 = n99855 & ~n99858;
  assign n99860 = n99814 & ~n99859;
  assign n99861 = n99837 & ~n99860;
  assign n99862 = ~n99816 & n99861;
  assign n99863 = ~pi8721 & ~n99862;
  assign n99864 = pi8721 & n99837;
  assign n99865 = ~n99816 & n99864;
  assign n99866 = ~n99860 & n99865;
  assign po5920 = n99863 | n99866;
  assign n99868 = ~n98714 & n98801;
  assign n99869 = ~n98830 & ~n99868;
  assign n99870 = n98714 & n98813;
  assign n99871 = ~n98720 & n98771;
  assign n99872 = ~n98714 & n98781;
  assign n99873 = ~n99871 & ~n99872;
  assign n99874 = ~n98780 & n99873;
  assign n99875 = ~n99870 & n99874;
  assign n99876 = ~n98785 & ~n98817;
  assign n99877 = n99875 & n99876;
  assign n99878 = ~n98822 & n99877;
  assign n99879 = n98739 & ~n99878;
  assign n99880 = ~n98720 & n98756;
  assign n99881 = ~n98714 & ~n99720;
  assign n99882 = ~n99880 & ~n99881;
  assign n99883 = ~n98720 & n98729;
  assign n99884 = ~n98781 & ~n99883;
  assign n99885 = ~n98753 & n99884;
  assign n99886 = n98714 & ~n99885;
  assign n99887 = n99882 & ~n99886;
  assign n99888 = ~n98739 & ~n99887;
  assign n99889 = ~n99879 & ~n99888;
  assign n99890 = ~n98833 & n99889;
  assign n99891 = n99869 & n99890;
  assign n99892 = pi8714 & n99891;
  assign n99893 = ~pi8714 & ~n99891;
  assign po5922 = n99892 | n99893;
  assign n99895 = ~n99522 & n99540;
  assign n99896 = ~n99567 & ~n99582;
  assign n99897 = n99895 & ~n99896;
  assign n99898 = ~n99522 & ~n99546;
  assign n99899 = n99567 & n99898;
  assign n99900 = ~n99897 & ~n99899;
  assign n99901 = n99559 & ~n99900;
  assign n99902 = ~n99540 & n99546;
  assign n99903 = n99564 & n99902;
  assign n99904 = ~n99599 & ~n99902;
  assign n99905 = n99522 & ~n99904;
  assign n99906 = ~n99540 & n99563;
  assign n99907 = ~n99905 & ~n99906;
  assign n99908 = ~n99903 & n99907;
  assign n99909 = n99559 & ~n99908;
  assign n99910 = ~n99901 & ~n99909;
  assign n99911 = n99540 & n99579;
  assign n99912 = ~n99540 & n99574;
  assign n99913 = ~n99911 & ~n99912;
  assign n99914 = ~n99522 & ~n99913;
  assign n99915 = ~n99562 & ~n99599;
  assign n99916 = n99540 & ~n99915;
  assign n99917 = ~n99574 & ~n99916;
  assign n99918 = ~n99522 & ~n99917;
  assign n99919 = ~n99534 & ~n99540;
  assign n99920 = n99898 & n99919;
  assign n99921 = n99534 & n99546;
  assign n99922 = ~n99574 & ~n99921;
  assign n99923 = ~n99540 & ~n99922;
  assign n99924 = n99522 & n99540;
  assign n99925 = n99564 & n99924;
  assign n99926 = ~n99546 & n99925;
  assign n99927 = ~n99923 & ~n99926;
  assign n99928 = ~n99920 & n99927;
  assign n99929 = ~n99918 & n99928;
  assign n99930 = ~n99911 & n99929;
  assign n99931 = ~n99559 & ~n99930;
  assign n99932 = n99540 & n99590;
  assign n99933 = ~n99540 & n99599;
  assign n99934 = ~n99932 & ~n99933;
  assign n99935 = n99522 & ~n99934;
  assign n99936 = ~n99931 & ~n99935;
  assign n99937 = ~n99914 & n99936;
  assign n99938 = n99910 & n99937;
  assign n99939 = pi8765 & n99938;
  assign n99940 = ~pi8765 & ~n99938;
  assign po5923 = n99939 | n99940;
  assign n99942 = ~n99649 & ~n99665;
  assign n99943 = n99340 & ~n99942;
  assign n99944 = ~n99332 & ~n99346;
  assign n99945 = ~n99652 & n99944;
  assign n99946 = ~n99298 & ~n99945;
  assign n99947 = n99340 & n99946;
  assign n99948 = ~n99943 & ~n99947;
  assign n99949 = n99341 & n99349;
  assign n99950 = ~n99351 & ~n99949;
  assign n99951 = ~n99345 & ~n99368;
  assign n99952 = n99298 & ~n99951;
  assign n99953 = n99340 & n99952;
  assign n99954 = n99950 & ~n99953;
  assign n99955 = ~n99304 & n99341;
  assign n99956 = ~n99304 & n99326;
  assign n99957 = ~n99325 & ~n99956;
  assign n99958 = n99298 & ~n99957;
  assign n99959 = ~n99333 & ~n99354;
  assign n99960 = ~n99304 & n99323;
  assign n99961 = ~n99376 & ~n99960;
  assign n99962 = ~n99298 & ~n99961;
  assign n99963 = n99959 & ~n99962;
  assign n99964 = ~n99958 & n99963;
  assign n99965 = ~n99955 & n99964;
  assign n99966 = ~n99340 & ~n99965;
  assign n99967 = ~n99384 & n99632;
  assign n99968 = n99298 & ~n99967;
  assign n99969 = ~n99966 & ~n99968;
  assign n99970 = n99954 & n99969;
  assign n99971 = n99948 & n99970;
  assign n99972 = ~pi8779 & ~n99971;
  assign n99973 = pi8779 & n99954;
  assign n99974 = n99948 & n99973;
  assign n99975 = n99969 & n99974;
  assign po5924 = n99972 | n99975;
  assign n99977 = ~n99192 & n99208;
  assign n99978 = n99193 & ~n99481;
  assign n99979 = ~n99202 & ~n99978;
  assign n99980 = ~n99222 & n99979;
  assign n99981 = n99192 & ~n99980;
  assign n99982 = ~n99162 & n99248;
  assign n99983 = ~n99981 & ~n99982;
  assign n99984 = ~n99168 & n99201;
  assign n99985 = n99162 & n99230;
  assign n99986 = ~n99484 & ~n99985;
  assign n99987 = ~n99984 & n99986;
  assign n99988 = ~n99192 & ~n99987;
  assign n99989 = n99983 & ~n99988;
  assign n99990 = n99218 & ~n99989;
  assign n99991 = ~n99977 & ~n99990;
  assign n99992 = n99162 & n99184;
  assign n99993 = ~n99182 & ~n99992;
  assign n99994 = ~n99192 & ~n99993;
  assign n99995 = ~n99203 & ~n99994;
  assign n99996 = ~n99208 & ~n99260;
  assign n99997 = n99162 & n99248;
  assign n99998 = ~n99162 & n99233;
  assign n99999 = ~n99230 & ~n99998;
  assign n100000 = ~n99984 & n99999;
  assign n100001 = n99192 & ~n100000;
  assign n100002 = ~n99997 & ~n100001;
  assign n100003 = n99996 & n100002;
  assign n100004 = n99995 & n100003;
  assign n100005 = ~n99218 & ~n100004;
  assign n100006 = ~n99270 & ~n99480;
  assign n100007 = n99192 & ~n100006;
  assign n100008 = ~n100005 & ~n100007;
  assign n100009 = n99991 & n100008;
  assign n100010 = pi8787 & n100009;
  assign n100011 = ~pi8787 & ~n100009;
  assign po5933 = n100010 | n100011;
  assign n100013 = ~n98856 & n98868;
  assign n100014 = ~n98938 & ~n100013;
  assign n100015 = ~n98869 & n100014;
  assign n100016 = n98876 & ~n100015;
  assign n100017 = ~n98868 & n98906;
  assign n100018 = ~n98856 & ~n98862;
  assign n100019 = n98885 & n100018;
  assign n100020 = n98862 & n98931;
  assign n100021 = ~n100019 & ~n100020;
  assign n100022 = n98856 & n98868;
  assign n100023 = n98862 & ~n98876;
  assign n100024 = n100022 & n100023;
  assign n100025 = n100021 & ~n100024;
  assign n100026 = ~n100017 & n100025;
  assign n100027 = ~n100016 & n100026;
  assign n100028 = ~n98850 & ~n100027;
  assign n100029 = ~n98856 & n98886;
  assign n100030 = n98862 & n100029;
  assign n100031 = ~n98856 & n98890;
  assign n100032 = ~n98862 & n100031;
  assign n100033 = ~n100030 & ~n100032;
  assign n100034 = n98876 & ~n100033;
  assign n100035 = ~n100028 & ~n100034;
  assign n100036 = ~n98862 & n98931;
  assign n100037 = ~n98897 & ~n98917;
  assign n100038 = n98876 & ~n100037;
  assign n100039 = ~n100036 & ~n100038;
  assign n100040 = ~n98920 & n100039;
  assign n100041 = n98850 & ~n100040;
  assign n100042 = ~n98890 & ~n98926;
  assign n100043 = n98856 & ~n100042;
  assign n100044 = ~n98911 & ~n100043;
  assign n100045 = ~n98876 & ~n100044;
  assign n100046 = n98850 & n100045;
  assign n100047 = ~n100041 & ~n100046;
  assign n100048 = n100035 & n100047;
  assign n100049 = pi8751 & n100048;
  assign n100050 = ~pi8751 & ~n100048;
  assign po5978 = n100049 | n100050;
  assign n100052 = ~n99833 & ~n99847;
  assign n100053 = ~n99798 & n100052;
  assign n100054 = n99808 & ~n100053;
  assign n100055 = ~n99788 & n99823;
  assign n100056 = n99788 & n99797;
  assign n100057 = ~n100055 & ~n100056;
  assign n100058 = ~n99808 & ~n100057;
  assign n100059 = ~n100054 & ~n100058;
  assign n100060 = ~n99822 & ~n99834;
  assign n100061 = n100059 & n100060;
  assign n100062 = n99814 & ~n100061;
  assign n100063 = ~n99782 & n99817;
  assign n100064 = n99788 & n100063;
  assign n100065 = ~n99851 & ~n100064;
  assign n100066 = ~n99808 & ~n100065;
  assign n100067 = n99782 & n99799;
  assign n100068 = ~n100063 & ~n100067;
  assign n100069 = n99808 & ~n100068;
  assign n100070 = ~n99782 & n100055;
  assign n100071 = ~n100069 & ~n100070;
  assign n100072 = ~n99808 & n99818;
  assign n100073 = n99801 & ~n100072;
  assign n100074 = ~n99847 & n100073;
  assign n100075 = n99782 & ~n100074;
  assign n100076 = n100071 & ~n100075;
  assign n100077 = ~n99814 & ~n100076;
  assign n100078 = n99788 & n99796;
  assign n100079 = n99838 & n100078;
  assign n100080 = ~n100077 & ~n100079;
  assign n100081 = ~n100066 & n100080;
  assign n100082 = ~n100062 & n100081;
  assign n100083 = ~pi8753 & ~n100082;
  assign n100084 = pi8753 & n100082;
  assign po5979 = n100083 | n100084;
  assign n100086 = ~n98984 & n99014;
  assign n100087 = n98984 & n99025;
  assign n100088 = ~n99011 & ~n100087;
  assign n100089 = n98958 & ~n100088;
  assign n100090 = ~n100086 & ~n100089;
  assign n100091 = ~n98976 & n99047;
  assign n100092 = n98970 & n100091;
  assign n100093 = n98993 & n99026;
  assign n100094 = ~n100092 & ~n100093;
  assign n100095 = ~n99746 & n100094;
  assign n100096 = ~n98988 & ~n99001;
  assign n100097 = ~n98991 & n100096;
  assign n100098 = n100095 & n100097;
  assign n100099 = n100090 & n100098;
  assign n100100 = ~n99023 & ~n100099;
  assign n100101 = ~n98987 & ~n99011;
  assign n100102 = n98984 & ~n100101;
  assign n100103 = ~n98984 & n98999;
  assign n100104 = ~n98964 & n98984;
  assign n100105 = ~n98976 & n100104;
  assign n100106 = n98970 & n100105;
  assign n100107 = ~n100103 & ~n100106;
  assign n100108 = ~n98958 & ~n100107;
  assign n100109 = ~n99040 & ~n99751;
  assign n100110 = n98964 & ~n98976;
  assign n100111 = n98984 & n100110;
  assign n100112 = n100109 & ~n100111;
  assign n100113 = n98958 & ~n100112;
  assign n100114 = ~n98984 & n98994;
  assign n100115 = ~n100113 & ~n100114;
  assign n100116 = ~n100108 & n100115;
  assign n100117 = ~n100102 & n100116;
  assign n100118 = n99023 & ~n100117;
  assign n100119 = n98958 & n99030;
  assign n100120 = ~n100118 & ~n100119;
  assign n100121 = ~n98958 & n100086;
  assign n100122 = n100120 & ~n100121;
  assign n100123 = ~n100100 & n100122;
  assign n100124 = ~pi8725 & ~n100123;
  assign n100125 = pi8725 & n100120;
  assign n100126 = ~n100100 & n100125;
  assign n100127 = ~n100121 & n100126;
  assign po5980 = n100124 | n100127;
  assign n100129 = ~n98964 & n99026;
  assign n100130 = n98970 & n100129;
  assign n100131 = ~n98984 & n100110;
  assign n100132 = ~n98992 & ~n100131;
  assign n100133 = ~n100106 & n100132;
  assign n100134 = ~n100130 & n100133;
  assign n100135 = n98958 & n98987;
  assign n100136 = n100134 & ~n100135;
  assign n100137 = n99023 & ~n100136;
  assign n100138 = ~n99041 & ~n100114;
  assign n100139 = n98958 & ~n100138;
  assign n100140 = ~n99023 & n99025;
  assign n100141 = ~n98958 & n100140;
  assign n100142 = ~n98970 & n99738;
  assign n100143 = ~n100110 & ~n100142;
  assign n100144 = ~n98994 & n100143;
  assign n100145 = n98958 & ~n100144;
  assign n100146 = ~n98984 & n99000;
  assign n100147 = ~n100145 & ~n100146;
  assign n100148 = ~n99023 & ~n100147;
  assign n100149 = ~n100141 & ~n100148;
  assign n100150 = ~n100139 & n100149;
  assign n100151 = ~n98988 & ~n98992;
  assign n100152 = ~n98984 & n99040;
  assign n100153 = ~n100087 & ~n100152;
  assign n100154 = n100151 & n100153;
  assign n100155 = ~n98958 & ~n100154;
  assign n100156 = n100150 & ~n100155;
  assign n100157 = ~n100137 & n100156;
  assign n100158 = pi8768 & n100157;
  assign n100159 = ~pi8768 & ~n100157;
  assign po6025 = n100158 | n100159;
  assign n100161 = ~n98887 & ~n98897;
  assign n100162 = ~n98917 & ~n100031;
  assign n100163 = n100161 & n100162;
  assign n100164 = ~n98862 & ~n100163;
  assign n100165 = ~n100020 & ~n100164;
  assign n100166 = ~n98896 & ~n100029;
  assign n100167 = n98927 & ~n100166;
  assign n100168 = n100165 & ~n100167;
  assign n100169 = ~n98850 & ~n100168;
  assign n100170 = n98862 & n98917;
  assign n100171 = ~n98862 & n100029;
  assign n100172 = ~n100170 & ~n100171;
  assign n100173 = ~n98876 & ~n100172;
  assign n100174 = ~n98862 & n100043;
  assign n100175 = ~n98885 & n100018;
  assign n100176 = ~n98892 & ~n100175;
  assign n100177 = ~n100031 & n100176;
  assign n100178 = n98876 & ~n100177;
  assign n100179 = ~n98876 & ~n100166;
  assign n100180 = ~n100178 & ~n100179;
  assign n100181 = ~n100174 & n100180;
  assign n100182 = ~n100170 & n100181;
  assign n100183 = n98850 & ~n100182;
  assign n100184 = ~n100173 & ~n100183;
  assign n100185 = ~n100169 & n100184;
  assign n100186 = pi8797 & n100185;
  assign n100187 = ~pi8797 & ~n100185;
  assign po6028 = n100186 | n100187;
  assign n100189 = n99528 & n99540;
  assign n100190 = ~n99534 & n100189;
  assign n100191 = ~n99540 & ~n99546;
  assign n100192 = n99534 & n100191;
  assign n100193 = ~n100190 & ~n100192;
  assign n100194 = n99522 & ~n100193;
  assign n100195 = ~n99540 & n99568;
  assign n100196 = ~n99920 & ~n100195;
  assign n100197 = n99534 & n99550;
  assign n100198 = ~n99582 & ~n100197;
  assign n100199 = ~n99522 & ~n100198;
  assign n100200 = n100196 & ~n100199;
  assign n100201 = ~n100194 & n100200;
  assign n100202 = ~n99549 & n100201;
  assign n100203 = ~n99903 & ~n99911;
  assign n100204 = n100202 & n100203;
  assign n100205 = n99559 & ~n100204;
  assign n100206 = ~n99528 & n99550;
  assign n100207 = n99540 & n99564;
  assign n100208 = ~n100206 & ~n100207;
  assign n100209 = n99522 & ~n100208;
  assign n100210 = n99560 & n99573;
  assign n100211 = ~n100209 & ~n100210;
  assign n100212 = n99562 & n99902;
  assign n100213 = n99591 & ~n100212;
  assign n100214 = n99522 & ~n100213;
  assign n100215 = ~n99540 & n99579;
  assign n100216 = ~n100214 & ~n100215;
  assign n100217 = n100211 & n100216;
  assign n100218 = ~n99559 & ~n100217;
  assign n100219 = ~n99568 & ~n99906;
  assign n100220 = ~n99575 & n100219;
  assign n100221 = n99596 & ~n100220;
  assign n100222 = ~n100218 & ~n100221;
  assign n100223 = ~n99549 & ~n99903;
  assign n100224 = ~n99522 & ~n100223;
  assign n100225 = n100222 & ~n100224;
  assign n100226 = ~n100205 & n100225;
  assign n100227 = ~pi8729 & n100226;
  assign n100228 = pi8729 & ~n100226;
  assign po6035 = n100227 | n100228;
  assign n100230 = n98876 & n100031;
  assign n100231 = ~n98862 & n98888;
  assign n100232 = ~n100019 & ~n100231;
  assign n100233 = ~n100230 & n100232;
  assign n100234 = n98862 & n98896;
  assign n100235 = ~n98862 & n98926;
  assign n100236 = ~n98877 & ~n100235;
  assign n100237 = ~n98876 & ~n100236;
  assign n100238 = ~n100234 & ~n100237;
  assign n100239 = n100233 & n100238;
  assign n100240 = n98850 & ~n100239;
  assign n100241 = ~n98905 & ~n98938;
  assign n100242 = n98876 & n100029;
  assign n100243 = ~n98933 & ~n100242;
  assign n100244 = n100241 & n100243;
  assign n100245 = ~n98850 & ~n100244;
  assign n100246 = ~n98850 & ~n98876;
  assign n100247 = n98856 & n98930;
  assign n100248 = ~n98862 & n100247;
  assign n100249 = ~n100031 & ~n100248;
  assign n100250 = ~n98887 & n100249;
  assign n100251 = n100246 & ~n100250;
  assign n100252 = ~n100245 & ~n100251;
  assign n100253 = n98862 & n98887;
  assign n100254 = ~n100020 & ~n100253;
  assign n100255 = ~n98876 & ~n100254;
  assign n100256 = n98906 & n98917;
  assign n100257 = ~n100255 & ~n100256;
  assign n100258 = ~n98946 & n100257;
  assign n100259 = n98862 & n100230;
  assign n100260 = n100258 & ~n100259;
  assign n100261 = n100252 & n100260;
  assign n100262 = ~n100240 & n100261;
  assign n100263 = pi8767 & n100262;
  assign n100264 = ~pi8767 & ~n100262;
  assign po6043 = n100263 | n100264;
  assign n100266 = ~n99453 & ~n99469;
  assign n100267 = ~n99421 & ~n99425;
  assign n100268 = ~n99397 & ~n99428;
  assign n100269 = n99079 & ~n100268;
  assign n100270 = ~n99126 & ~n100269;
  assign n100271 = n100267 & n100270;
  assign n100272 = ~n99088 & ~n100271;
  assign n100273 = ~n99067 & n99094;
  assign n100274 = ~n99102 & ~n100273;
  assign n100275 = ~n99073 & ~n100274;
  assign n100276 = ~n99116 & ~n99456;
  assign n100277 = n99079 & ~n100276;
  assign n100278 = ~n99073 & n99094;
  assign n100279 = ~n99132 & ~n100278;
  assign n100280 = ~n99118 & n100279;
  assign n100281 = ~n99079 & ~n100280;
  assign n100282 = ~n100277 & ~n100281;
  assign n100283 = ~n100275 & n100282;
  assign n100284 = n99088 & ~n100283;
  assign n100285 = ~n99393 & ~n99445;
  assign n100286 = ~n99410 & n100285;
  assign n100287 = ~n99079 & ~n100286;
  assign n100288 = ~n100284 & ~n100287;
  assign n100289 = ~n100272 & n100288;
  assign n100290 = n100266 & n100289;
  assign n100291 = pi8720 & n100290;
  assign n100292 = ~pi8720 & ~n100290;
  assign po6071 = n100291 | n100292;
  assign n100294 = n99808 & n99814;
  assign n100295 = ~n99821 & ~n99824;
  assign n100296 = ~n99841 & n99843;
  assign n100297 = n100295 & ~n100296;
  assign n100298 = n100294 & ~n100297;
  assign n100299 = n99782 & n99823;
  assign n100300 = ~n99782 & n99796;
  assign n100301 = n99788 & n100300;
  assign n100302 = ~n100063 & ~n100301;
  assign n100303 = ~n99818 & n100302;
  assign n100304 = ~n100299 & n100303;
  assign n100305 = ~n99808 & ~n100304;
  assign n100306 = ~n99782 & n99800;
  assign n100307 = ~n100305 & ~n100306;
  assign n100308 = n99814 & ~n100307;
  assign n100309 = ~n100298 & ~n100308;
  assign n100310 = ~n99845 & ~n99849;
  assign n100311 = ~n99788 & n99796;
  assign n100312 = ~n99782 & n100311;
  assign n100313 = ~n99824 & ~n100312;
  assign n100314 = ~n99808 & ~n100313;
  assign n100315 = ~n99841 & ~n99843;
  assign n100316 = n99808 & n100315;
  assign n100317 = ~n99823 & n99856;
  assign n100318 = n99788 & n100317;
  assign n100319 = ~n100316 & ~n100318;
  assign n100320 = ~n100314 & n100319;
  assign n100321 = n100310 & n100320;
  assign n100322 = ~n99814 & ~n100321;
  assign n100323 = n100309 & ~n100322;
  assign n100324 = n99798 & n99808;
  assign n100325 = ~n99782 & n100324;
  assign n100326 = ~n99808 & n100055;
  assign n100327 = n99782 & n100326;
  assign n100328 = n99799 & n99856;
  assign n100329 = n99788 & n100328;
  assign n100330 = ~n100327 & ~n100329;
  assign n100331 = ~n100325 & n100330;
  assign n100332 = n100323 & n100331;
  assign n100333 = pi8747 & n100332;
  assign n100334 = ~pi8747 & ~n100332;
  assign po6086 = n100333 | n100334;
  assign n100336 = n99522 & n99565;
  assign n100337 = n99540 & n99582;
  assign n100338 = n99546 & n99895;
  assign n100339 = ~n100191 & ~n100338;
  assign n100340 = n99528 & ~n100339;
  assign n100341 = ~n100192 & ~n100340;
  assign n100342 = ~n99549 & n100341;
  assign n100343 = ~n100337 & n100342;
  assign n100344 = ~n100336 & n100343;
  assign n100345 = ~n99559 & ~n100344;
  assign n100346 = ~n99540 & n99564;
  assign n100347 = ~n99563 & ~n100346;
  assign n100348 = ~n99522 & ~n100347;
  assign n100349 = n99522 & ~n99922;
  assign n100350 = ~n99932 & ~n100349;
  assign n100351 = ~n100348 & n100350;
  assign n100352 = n99559 & ~n100351;
  assign n100353 = ~n100195 & ~n100207;
  assign n100354 = n99522 & ~n100353;
  assign n100355 = ~n99522 & n99579;
  assign n100356 = ~n100354 & ~n100355;
  assign n100357 = ~n100352 & n100356;
  assign n100358 = ~n100345 & n100357;
  assign n100359 = pi8693 & n100358;
  assign n100360 = ~pi8693 & ~n100358;
  assign po6118 = n100359 | n100360;
  assign n100362 = ~n100063 & ~n100299;
  assign n100363 = ~n99808 & ~n100362;
  assign n100364 = ~n100329 & ~n100363;
  assign n100365 = ~n99814 & ~n100364;
  assign n100366 = ~n99797 & ~n100078;
  assign n100367 = n99782 & ~n100366;
  assign n100368 = ~n100055 & ~n100367;
  assign n100369 = n99808 & ~n100368;
  assign n100370 = ~n100296 & ~n100369;
  assign n100371 = ~n99782 & n99847;
  assign n100372 = ~n99776 & n99789;
  assign n100373 = ~n99782 & ~n100366;
  assign n100374 = ~n100372 & ~n100373;
  assign n100375 = ~n99808 & ~n100374;
  assign n100376 = ~n100371 & ~n100375;
  assign n100377 = n100370 & n100376;
  assign n100378 = n99814 & ~n100377;
  assign n100379 = ~n99782 & ~n99788;
  assign n100380 = ~n99797 & n100379;
  assign n100381 = ~n99814 & n100380;
  assign n100382 = n99797 & n99831;
  assign n100383 = ~n99808 & n100382;
  assign n100384 = ~n99788 & n99838;
  assign n100385 = ~n99776 & n100384;
  assign n100386 = ~n100383 & ~n100385;
  assign n100387 = ~n100381 & n100386;
  assign n100388 = ~n99818 & ~n100300;
  assign n100389 = n99815 & ~n100388;
  assign n100390 = n100387 & ~n100389;
  assign n100391 = ~n100378 & n100390;
  assign n100392 = ~n100365 & n100391;
  assign n100393 = pi8784 & n100392;
  assign n100394 = ~pi8784 & ~n100392;
  assign po6125 = n100393 | n100394;
  assign n100396 = pi9007 & ~pi9040;
  assign n100397 = pi8895 & pi9040;
  assign po8158 = n100396 | n100397;
  assign n100399 = pi8925 & ~pi9040;
  assign n100400 = pi9037 & pi9040;
  assign po8159 = n100399 | n100400;
  assign n100402 = pi8993 & ~pi9040;
  assign n100403 = pi8881 & pi9040;
  assign po8160 = n100402 | n100403;
  assign n100405 = pi8906 & ~pi9040;
  assign n100406 = pi9018 & pi9040;
  assign po8161 = n100405 | n100406;
  assign n100408 = pi9024 & ~pi9040;
  assign n100409 = pi8912 & pi9040;
  assign po8162 = n100408 | n100409;
  assign n100411 = pi8992 & ~pi9040;
  assign n100412 = pi8880 & pi9040;
  assign po8163 = n100411 | n100412;
  assign n100414 = pi9009 & ~pi9040;
  assign n100415 = pi8897 & pi9040;
  assign po8164 = n100414 | n100415;
  assign n100417 = pi8875 & ~pi9040;
  assign n100418 = pi8987 & pi9040;
  assign po8165 = n100417 | n100418;
  assign n100420 = pi9029 & ~pi9040;
  assign n100421 = pi8917 & pi9040;
  assign po8166 = n100420 | n100421;
  assign n100423 = pi8914 & ~pi9040;
  assign n100424 = pi9026 & pi9040;
  assign po8167 = n100423 | n100424;
  assign n100426 = pi8994 & ~pi9040;
  assign n100427 = pi8882 & pi9040;
  assign po8168 = n100426 | n100427;
  assign n100429 = pi8877 & ~pi9040;
  assign n100430 = pi8989 & pi9040;
  assign po8169 = n100429 | n100430;
  assign n100432 = pi8916 & ~pi9040;
  assign n100433 = pi9028 & pi9040;
  assign po8170 = n100432 | n100433;
  assign n100435 = pi9010 & ~pi9040;
  assign n100436 = pi8898 & pi9040;
  assign po8171 = n100435 | n100436;
  assign n100438 = pi8902 & ~pi9040;
  assign n100439 = pi9014 & pi9040;
  assign po8172 = n100438 | n100439;
  assign n100441 = pi8924 & ~pi9040;
  assign n100442 = pi9036 & pi9040;
  assign po8173 = n100441 | n100442;
  assign n100444 = pi9039 & ~pi9040;
  assign n100445 = pi8927 & pi9040;
  assign po8174 = n100444 | n100445;
  assign n100447 = pi8988 & ~pi9040;
  assign n100448 = pi8876 & pi9040;
  assign po8175 = n100447 | n100448;
  assign n100450 = pi8909 & ~pi9040;
  assign n100451 = pi9021 & pi9040;
  assign po8176 = n100450 | n100451;
  assign n100453 = pi9004 & ~pi9040;
  assign n100454 = pi8892 & pi9040;
  assign po8177 = n100453 | n100454;
  assign n100456 = pi9002 & ~pi9040;
  assign n100457 = pi8890 & pi9040;
  assign po8178 = n100456 | n100457;
  assign n100459 = pi8897 & ~pi9040;
  assign n100460 = pi9009 & pi9040;
  assign po8179 = n100459 | n100460;
  assign n100462 = pi9018 & ~pi9040;
  assign n100463 = pi8906 & pi9040;
  assign po8180 = n100462 | n100463;
  assign n100465 = pi9017 & ~pi9040;
  assign n100466 = pi8905 & pi9040;
  assign po8181 = n100465 | n100466;
  assign n100468 = pi8912 & ~pi9040;
  assign n100469 = pi9024 & pi9040;
  assign po8182 = n100468 | n100469;
  assign n100471 = pi9037 & ~pi9040;
  assign n100472 = pi8925 & pi9040;
  assign po8183 = n100471 | n100472;
  assign n100474 = pi8881 & ~pi9040;
  assign n100475 = pi8993 & pi9040;
  assign po8184 = n100474 | n100475;
  assign n100477 = pi9032 & ~pi9040;
  assign n100478 = pi8920 & pi9040;
  assign po8185 = n100477 | n100478;
  assign n100480 = pi9035 & ~pi9040;
  assign n100481 = pi8923 & pi9040;
  assign po8186 = n100480 | n100481;
  assign n100483 = pi8917 & ~pi9040;
  assign n100484 = pi9029 & pi9040;
  assign po8187 = n100483 | n100484;
  assign n100486 = pi8907 & ~pi9040;
  assign n100487 = pi9019 & pi9040;
  assign po8188 = n100486 | n100487;
  assign n100489 = pi8889 & ~pi9040;
  assign n100490 = pi9001 & pi9040;
  assign po8189 = n100489 | n100490;
  assign n100492 = pi8985 & ~pi9040;
  assign n100493 = pi8873 & pi9040;
  assign po8190 = n100492 | n100493;
  assign n100495 = pi8880 & ~pi9040;
  assign n100496 = pi8992 & pi9040;
  assign po8191 = n100495 | n100496;
  assign n100498 = pi9026 & ~pi9040;
  assign n100499 = pi8914 & pi9040;
  assign po8192 = n100498 | n100499;
  assign n100501 = pi8905 & ~pi9040;
  assign n100502 = pi9017 & pi9040;
  assign po8193 = n100501 | n100502;
  assign n100504 = pi8991 & ~pi9040;
  assign n100505 = pi8879 & pi9040;
  assign po8194 = n100504 | n100505;
  assign n100507 = pi8915 & ~pi9040;
  assign n100508 = pi9027 & pi9040;
  assign po8195 = n100507 | n100508;
  assign n100510 = pi8903 & ~pi9040;
  assign n100511 = pi9015 & pi9040;
  assign po8196 = n100510 | n100511;
  assign n100513 = pi9016 & ~pi9040;
  assign n100514 = pi8904 & pi9040;
  assign po8197 = n100513 | n100514;
  assign n100516 = pi8888 & ~pi9040;
  assign n100517 = pi9000 & pi9040;
  assign po8198 = n100516 | n100517;
  assign n100519 = pi9028 & ~pi9040;
  assign n100520 = pi8916 & pi9040;
  assign po8199 = n100519 | n100520;
  assign n100522 = pi8999 & ~pi9040;
  assign n100523 = pi8887 & pi9040;
  assign po8200 = n100522 | n100523;
  assign n100525 = pi8920 & ~pi9040;
  assign n100526 = pi9032 & pi9040;
  assign po8201 = n100525 | n100526;
  assign n100528 = pi8876 & ~pi9040;
  assign n100529 = pi8988 & pi9040;
  assign po8202 = n100528 | n100529;
  assign n100531 = pi9015 & ~pi9040;
  assign n100532 = pi8903 & pi9040;
  assign po8203 = n100531 | n100532;
  assign n100534 = pi8883 & ~pi9040;
  assign n100535 = pi8995 & pi9040;
  assign po8204 = n100534 | n100535;
  assign n100537 = pi8891 & ~pi9040;
  assign n100538 = pi9003 & pi9040;
  assign po8205 = n100537 | n100538;
  assign n100540 = pi9019 & ~pi9040;
  assign n100541 = pi8907 & pi9040;
  assign po8206 = n100540 | n100541;
  assign n100543 = pi8882 & ~pi9040;
  assign n100544 = pi8994 & pi9040;
  assign po8207 = n100543 | n100544;
  assign n100546 = pi8895 & ~pi9040;
  assign n100547 = pi9007 & pi9040;
  assign po8208 = n100546 | n100547;
  assign n100549 = pi8894 & ~pi9040;
  assign n100550 = pi9006 & pi9040;
  assign po8209 = n100549 | n100550;
  assign n100552 = pi9038 & ~pi9040;
  assign n100553 = pi8926 & pi9040;
  assign po8210 = n100552 | n100553;
  assign n100555 = pi9021 & ~pi9040;
  assign n100556 = pi8909 & pi9040;
  assign po8211 = n100555 | n100556;
  assign n100558 = pi8987 & ~pi9040;
  assign n100559 = pi8875 & pi9040;
  assign po8212 = n100558 | n100559;
  assign n100561 = pi9003 & ~pi9040;
  assign n100562 = pi8891 & pi9040;
  assign po8213 = n100561 | n100562;
  assign n100564 = pi8996 & ~pi9040;
  assign n100565 = pi8884 & pi9040;
  assign po8214 = n100564 | n100565;
  assign n100567 = pi8997 & ~pi9040;
  assign n100568 = pi8885 & pi9040;
  assign po8215 = n100567 | n100568;
  assign n100570 = pi8899 & ~pi9040;
  assign n100571 = pi9011 & pi9040;
  assign po8216 = n100570 | n100571;
  assign n100573 = pi8995 & ~pi9040;
  assign n100574 = pi8883 & pi9040;
  assign po8217 = n100573 | n100574;
  assign n100576 = pi9013 & ~pi9040;
  assign n100577 = pi8901 & pi9040;
  assign po8218 = n100576 | n100577;
  assign n100579 = pi9014 & ~pi9040;
  assign n100580 = pi8902 & pi9040;
  assign po8219 = n100579 | n100580;
  assign n100582 = pi9025 & ~pi9040;
  assign n100583 = pi8913 & pi9040;
  assign po8220 = n100582 | n100583;
  assign n100585 = pi8900 & ~pi9040;
  assign n100586 = pi9012 & pi9040;
  assign po8221 = n100585 | n100586;
  assign n100588 = pi9005 & ~pi9040;
  assign n100589 = pi8893 & pi9040;
  assign po8222 = n100588 | n100589;
  assign n100591 = pi9011 & ~pi9040;
  assign n100592 = pi8899 & pi9040;
  assign po8223 = n100591 | n100592;
  assign n100594 = pi9012 & ~pi9040;
  assign n100595 = pi8900 & pi9040;
  assign po8224 = n100594 | n100595;
  assign n100597 = pi9022 & ~pi9040;
  assign n100598 = pi8910 & pi9040;
  assign po8225 = n100597 | n100598;
  assign n100600 = pi9006 & ~pi9040;
  assign n100601 = pi8894 & pi9040;
  assign po8226 = n100600 | n100601;
  assign n100603 = pi8923 & ~pi9040;
  assign n100604 = pi9035 & pi9040;
  assign po8227 = n100603 | n100604;
  assign n100606 = pi8885 & ~pi9040;
  assign n100607 = pi8997 & pi9040;
  assign po8228 = n100606 | n100607;
  assign n100609 = pi8901 & ~pi9040;
  assign n100610 = pi9013 & pi9040;
  assign po8229 = n100609 | n100610;
  assign n100612 = pi8913 & ~pi9040;
  assign n100613 = pi9025 & pi9040;
  assign po8230 = n100612 | n100613;
  assign n100615 = pi8908 & ~pi9040;
  assign n100616 = pi9020 & pi9040;
  assign po8231 = n100615 | n100616;
  assign n100618 = pi8990 & ~pi9040;
  assign n100619 = pi8878 & pi9040;
  assign po8232 = n100618 | n100619;
  assign n100621 = pi8893 & ~pi9040;
  assign n100622 = pi9005 & pi9040;
  assign po8233 = n100621 | n100622;
  assign n100624 = pi8886 & ~pi9040;
  assign n100625 = pi8998 & pi9040;
  assign po8234 = n100624 | n100625;
  assign n100627 = pi8919 & ~pi9040;
  assign n100628 = pi9031 & pi9040;
  assign po8235 = n100627 | n100628;
  assign n100630 = pi9020 & ~pi9040;
  assign n100631 = pi8908 & pi9040;
  assign po8236 = n100630 | n100631;
  assign n100633 = pi8911 & ~pi9040;
  assign n100634 = pi9023 & pi9040;
  assign po8237 = n100633 | n100634;
  assign n100636 = pi9008 & ~pi9040;
  assign n100637 = pi8896 & pi9040;
  assign po8238 = n100636 | n100637;
  assign n100639 = pi9000 & ~pi9040;
  assign n100640 = pi8888 & pi9040;
  assign po8239 = n100639 | n100640;
  assign n100642 = pi8926 & ~pi9040;
  assign n100643 = pi9038 & pi9040;
  assign po8240 = n100642 | n100643;
  assign n100645 = pi8910 & ~pi9040;
  assign n100646 = pi9022 & pi9040;
  assign po8241 = n100645 | n100646;
  assign n100648 = pi8989 & ~pi9040;
  assign n100649 = pi8877 & pi9040;
  assign po8242 = n100648 | n100649;
  assign n100651 = pi8873 & ~pi9040;
  assign n100652 = pi8985 & pi9040;
  assign po8243 = n100651 | n100652;
  assign n100654 = pi8998 & ~pi9040;
  assign n100655 = pi8886 & pi9040;
  assign po8244 = n100654 | n100655;
  assign n100657 = pi8921 & ~pi9040;
  assign n100658 = pi9033 & pi9040;
  assign po8245 = n100657 | n100658;
  assign n100660 = pi8878 & ~pi9040;
  assign n100661 = pi8990 & pi9040;
  assign po8246 = n100660 | n100661;
  assign n100663 = pi8887 & ~pi9040;
  assign n100664 = pi8999 & pi9040;
  assign po8247 = n100663 | n100664;
  assign n100666 = pi9030 & ~pi9040;
  assign n100667 = pi8918 & pi9040;
  assign po8248 = n100666 | n100667;
  assign n100669 = pi9034 & ~pi9040;
  assign n100670 = pi8922 & pi9040;
  assign po8249 = n100669 | n100670;
  assign n100672 = pi8918 & ~pi9040;
  assign n100673 = pi9030 & pi9040;
  assign po8250 = n100672 | n100673;
  assign n100675 = pi9023 & ~pi9040;
  assign n100676 = pi8911 & pi9040;
  assign po8251 = n100675 | n100676;
  assign n100678 = pi8892 & ~pi9040;
  assign n100679 = pi9004 & pi9040;
  assign po8252 = n100678 | n100679;
  assign n100681 = pi8896 & ~pi9040;
  assign n100682 = pi9008 & pi9040;
  assign po8253 = n100681 | n100682;
  assign n100684 = pi9033 & ~pi9040;
  assign n100685 = pi8921 & pi9040;
  assign po8254 = n100684 | n100685;
  assign n100687 = pi8927 & ~pi9040;
  assign n100688 = pi9039 & pi9040;
  assign po8255 = n100687 | n100688;
  assign n100690 = pi8986 & ~pi9040;
  assign n100691 = pi8874 & pi9040;
  assign po8256 = n100690 | n100691;
  assign n100693 = pi9031 & ~pi9040;
  assign n100694 = pi8919 & pi9040;
  assign po8257 = n100693 | n100694;
  assign n100696 = pi8879 & ~pi9040;
  assign n100697 = pi8991 & pi9040;
  assign po8258 = n100696 | n100697;
  assign n100699 = pi9036 & ~pi9040;
  assign n100700 = pi8924 & pi9040;
  assign po8259 = n100699 | n100700;
  assign n100702 = pi8884 & ~pi9040;
  assign n100703 = pi8996 & pi9040;
  assign po8260 = n100702 | n100703;
  assign n100705 = pi8890 & ~pi9040;
  assign n100706 = pi9002 & pi9040;
  assign po8261 = n100705 | n100706;
  assign n100708 = pi9001 & ~pi9040;
  assign n100709 = pi8889 & pi9040;
  assign po8262 = n100708 | n100709;
  assign n100711 = pi8874 & ~pi9040;
  assign n100712 = pi8986 & pi9040;
  assign po8263 = n100711 | n100712;
  assign n100714 = pi8898 & ~pi9040;
  assign n100715 = pi9010 & pi9040;
  assign po8264 = n100714 | n100715;
  assign n100717 = pi9027 & ~pi9040;
  assign n100718 = pi8915 & pi9040;
  assign po8265 = n100717 | n100718;
  assign n100720 = pi8904 & ~pi9040;
  assign n100721 = pi9016 & pi9040;
  assign po8266 = n100720 | n100721;
  assign n100723 = pi8984 & ~pi9040;
  assign n100724 = pi8872 & pi9040;
  assign po8267 = n100723 | n100724;
  assign n100726 = pi8922 & ~pi9040;
  assign n100727 = pi9034 & pi9040;
  assign po8268 = n100726 | n100727;
  assign n100729 = pi8872 & ~pi9040;
  assign n100730 = pi8984 & pi9040;
  assign po8269 = n100729 | n100730;
  assign po0064 = 1'b1;
  assign po0066 = ~po0068;
  assign po0071 = ~pi0105;
  assign po0074 = ~pi0110;
  assign po0077 = ~pi0108;
  assign po0080 = ~pi0104;
  assign po0083 = ~pi0103;
  assign po0086 = ~pi0125;
  assign po0089 = ~pi0100;
  assign po0092 = ~pi0099;
  assign po0095 = ~pi0139;
  assign po0098 = ~pi0096;
  assign po0101 = ~pi0102;
  assign po0104 = ~pi0111;
  assign po0107 = ~pi0115;
  assign po0110 = ~pi0117;
  assign po0113 = ~pi0098;
  assign po0116 = ~pi0097;
  assign po0119 = ~pi0121;
  assign po0122 = ~pi0116;
  assign po0125 = ~pi0101;
  assign po0128 = ~pi0126;
  assign po0131 = ~pi0123;
  assign po0134 = ~pi0158;
  assign po0137 = ~pi0137;
  assign po0140 = ~po0138;
  assign po0143 = ~pi0128;
  assign po0146 = ~pi0135;
  assign po0149 = ~pi0124;
  assign po0152 = ~pi0130;
  assign po0155 = ~pi0136;
  assign po0158 = ~pi0138;
  assign po0161 = ~pi0109;
  assign po0177 = ~pi0069;
  assign po1125 = ~po1127;
  assign po1133 = ~pi1203;
  assign po1139 = ~pi1189;
  assign po1147 = ~pi1195;
  assign po1155 = ~pi1197;
  assign po1158 = ~pi1204;
  assign po1166 = ~po1164;
  assign po1172 = ~pi1185;
  assign po1176 = ~pi1191;
  assign po1179 = ~pi1187;
  assign po1182 = ~pi1188;
  assign po1185 = ~pi1194;
  assign po1188 = ~pi1190;
  assign po1191 = ~pi1211;
  assign po1194 = ~pi1218;
  assign po1200 = ~pi1228;
  assign po1205 = ~pi1207;
  assign po1208 = ~pi1199;
  assign po1211 = ~pi1186;
  assign po1214 = ~pi1196;
  assign po1217 = ~pi1205;
  assign po1221 = ~pi1201;
  assign po1224 = ~pi1233;
  assign po1227 = ~pi1184;
  assign po1231 = ~pi1202;
  assign po1234 = ~pi1192;
  assign po1238 = ~pi1193;
  assign po1241 = ~pi1212;
  assign po1298 = ~pi1145;
  assign po1311 = ~pi1153;
  assign po1318 = ~pi1163;
  assign po1335 = ~pi1174;
  assign po1342 = ~pi1181;
  assign po2271 = ~pi2303;
  assign po2279 = ~pi2290;
  assign po2292 = ~pi2279;
  assign po2296 = ~pi2302;
  assign po2302 = ~pi2309;
  assign po2305 = ~pi2277;
  assign po2308 = ~pi2299;
  assign po2313 = ~pi2294;
  assign po2318 = ~pi2286;
  assign po2321 = ~pi2317;
  assign po2323 = ~po2325;
  assign po2328 = ~pi2278;
  assign po2332 = ~pi2293;
  assign po2336 = ~pi2287;
  assign po2339 = ~po2337;
  assign po2342 = ~pi2284;
  assign po2349 = ~pi2300;
  assign po2355 = ~pi2283;
  assign po2358 = ~pi2273;
  assign po2361 = ~pi2292;
  assign po2365 = ~pi2280;
  assign po2373 = ~pi2282;
  assign po2400 = ~pi2198;
  assign po2417 = ~pi2216;
  assign po2444 = ~pi2247;
  assign po2469 = ~pi2263;
  assign po2480 = ~pi2269;
  assign po2489 = ~pi2270;
  assign po2704 = ~pi2498;
  assign po3551 = ~pi3361;
  assign po3712 = ~pi3524;
  assign po3872 = ~pi3689;
  assign po5562 = ~pi5546;
  assign po5635 = ~pi5567;
  assign po5727 = ~pi5684;
  assign po5896 = ~pi5835;
  assign po6380 = ~pi6315;
  assign po6400 = ~pi6383;
  assign po6968 = ~pi6918;
  assign po6999 = ~pi6868;
  assign po0000 = pi0012;
  assign po0001 = pi0046;
  assign po0002 = pi0001;
  assign po0003 = pi0042;
  assign po0004 = pi0003;
  assign po0005 = pi0057;
  assign po0006 = pi0014;
  assign po0007 = pi0041;
  assign po0008 = pi0020;
  assign po0009 = pi0040;
  assign po0010 = pi0023;
  assign po0011 = pi0082;
  assign po0012 = pi0018;
  assign po0013 = pi0054;
  assign po0014 = pi0013;
  assign po0015 = pi0039;
  assign po0016 = pi0026;
  assign po0017 = pi0047;
  assign po0018 = pi0011;
  assign po0019 = pi0072;
  assign po0020 = pi0015;
  assign po0021 = pi0062;
  assign po0022 = pi0022;
  assign po0023 = pi0073;
  assign po0024 = pi0005;
  assign po0025 = pi0037;
  assign po0026 = pi0008;
  assign po0027 = pi0033;
  assign po0028 = pi0016;
  assign po0029 = pi0034;
  assign po0030 = pi0007;
  assign po0031 = pi0045;
  assign po0032 = pi0010;
  assign po0033 = pi0043;
  assign po0034 = pi0024;
  assign po0035 = pi0038;
  assign po0036 = pi0002;
  assign po0037 = pi0056;
  assign po0038 = pi0019;
  assign po0039 = pi0032;
  assign po0040 = pi0030;
  assign po0041 = pi0081;
  assign po0042 = pi0004;
  assign po0043 = pi0044;
  assign po0044 = pi0009;
  assign po0045 = pi0079;
  assign po0046 = pi0029;
  assign po0047 = pi0078;
  assign po0048 = pi0000;
  assign po0049 = pi0053;
  assign po0050 = pi0006;
  assign po0051 = pi0080;
  assign po0052 = pi0028;
  assign po0053 = pi0048;
  assign po0054 = pi0025;
  assign po0055 = pi0055;
  assign po0056 = pi0021;
  assign po0057 = pi0035;
  assign po0058 = pi0027;
  assign po0059 = pi0052;
  assign po0060 = pi0031;
  assign po0061 = pi0063;
  assign po0062 = pi0017;
  assign po0063 = pi0051;
  assign po0065 = pi9041;
  assign po0067 = pi0113;
  assign po0069 = pi0105;
  assign po0072 = pi0110;
  assign po0075 = pi0108;
  assign po0078 = pi0104;
  assign po0081 = pi0103;
  assign po0084 = pi0125;
  assign po0087 = pi0100;
  assign po0090 = pi0099;
  assign po0093 = pi0139;
  assign po0096 = pi0096;
  assign po0099 = pi0102;
  assign po0102 = pi0111;
  assign po0105 = pi0115;
  assign po0108 = pi0117;
  assign po0111 = pi0098;
  assign po0114 = pi0097;
  assign po0117 = pi0121;
  assign po0120 = pi0116;
  assign po0123 = pi0101;
  assign po0126 = pi0126;
  assign po0129 = pi0123;
  assign po0132 = pi0158;
  assign po0135 = pi0137;
  assign po0139 = pi0118;
  assign po0141 = pi0128;
  assign po0144 = pi0135;
  assign po0147 = pi0124;
  assign po0150 = pi0130;
  assign po0153 = pi0136;
  assign po0156 = pi0138;
  assign po0159 = pi0109;
  assign po0162 = pi0036;
  assign po0163 = pi0058;
  assign po0164 = pi0049;
  assign po0165 = pi0070;
  assign po0167 = pi0061;
  assign po0168 = pi0060;
  assign po0169 = pi0067;
  assign po0170 = pi0050;
  assign po0171 = pi0066;
  assign po0172 = pi0083;
  assign po0173 = pi0068;
  assign po0174 = pi0064;
  assign po0175 = pi0077;
  assign po0176 = pi0076;
  assign po0178 = pi0059;
  assign po0181 = pi0086;
  assign po0182 = pi0087;
  assign po0183 = pi0074;
  assign po0184 = pi0065;
  assign po0185 = pi0071;
  assign po0186 = pi0084;
  assign po0187 = pi0088;
  assign po0192 = pi0075;
  assign po0193 = pi0092;
  assign po0202 = pi0085;
  assign po0203 = pi0095;
  assign po0208 = pi0091;
  assign po0209 = pi0089;
  assign po0210 = pi0090;
  assign po0211 = pi0093;
  assign po0212 = pi0094;
  assign po0226 = pi0107;
  assign po0227 = pi0122;
  assign po0228 = pi0106;
  assign po0229 = pi0132;
  assign po0230 = pi0119;
  assign po0231 = pi0120;
  assign po0232 = pi0112;
  assign po0233 = pi0127;
  assign po0234 = pi0114;
  assign po0235 = pi0131;
  assign po0238 = pi0152;
  assign po0239 = pi0153;
  assign po0240 = pi0140;
  assign po0241 = pi0142;
  assign po0243 = pi0129;
  assign po0245 = pi0133;
  assign po0246 = pi0134;
  assign po0247 = pi0146;
  assign po0248 = pi0147;
  assign po0251 = pi0148;
  assign po0253 = pi0150;
  assign po0254 = pi0155;
  assign po0255 = pi0141;
  assign po0256 = pi0143;
  assign po0258 = pi0144;
  assign po0260 = pi0145;
  assign po0265 = pi0149;
  assign po0266 = pi0151;
  assign po0267 = pi0154;
  assign po0268 = pi0156;
  assign po0269 = pi0157;
  assign po0288 = pi0159;
  assign po0290 = pi0177;
  assign po0291 = pi0176;
  assign po0292 = pi0180;
  assign po0293 = pi0181;
  assign po0294 = pi0182;
  assign po0295 = pi0198;
  assign po0296 = pi0203;
  assign po0297 = pi0193;
  assign po0298 = pi0184;
  assign po0299 = pi0196;
  assign po0300 = pi0205;
  assign po0301 = pi0201;
  assign po0302 = pi0202;
  assign po0303 = pi0204;
  assign po0304 = pi0207;
  assign po0305 = pi0185;
  assign po0308 = pi0206;
  assign po0309 = pi0208;
  assign po0313 = pi0221;
  assign po0316 = pi0211;
  assign po0317 = pi0212;
  assign po0318 = pi0213;
  assign po0319 = pi0214;
  assign po0320 = pi0215;
  assign po0321 = pi0216;
  assign po0322 = pi0217;
  assign po0324 = pi0209;
  assign po0325 = pi0218;
  assign po0327 = pi0223;
  assign po0329 = pi0219;
  assign po0330 = pi0220;
  assign po0340 = pi0222;
  assign po0354 = pi0251;
  assign po0355 = pi0245;
  assign po0356 = pi0256;
  assign po0357 = pi0250;
  assign po0358 = pi0254;
  assign po0359 = pi0255;
  assign po0360 = pi0257;
  assign po0361 = pi0266;
  assign po0362 = pi0274;
  assign po0363 = pi0261;
  assign po0364 = pi0262;
  assign po0365 = pi0263;
  assign po0366 = pi0275;
  assign po0367 = pi0271;
  assign po0368 = pi0264;
  assign po0369 = pi0265;
  assign po0370 = pi0269;
  assign po0371 = pi0270;
  assign po0372 = pi0272;
  assign po0373 = pi0280;
  assign po0374 = pi0273;
  assign po0376 = pi0277;
  assign po0377 = pi0278;
  assign po0378 = pi0276;
  assign po0379 = pi0279;
  assign po0382 = pi0281;
  assign po0383 = pi0286;
  assign po0388 = pi0283;
  assign po0389 = pi0284;
  assign po0390 = pi0285;
  assign po0397 = pi0282;
  assign po0398 = pi0287;
  assign po0418 = pi0302;
  assign po0419 = pi0323;
  assign po0420 = pi0312;
  assign po0421 = pi0315;
  assign po0422 = pi0322;
  assign po0423 = pi0326;
  assign po0424 = pi0335;
  assign po0425 = pi0329;
  assign po0426 = pi0324;
  assign po0427 = pi0330;
  assign po0428 = pi0341;
  assign po0429 = pi0325;
  assign po0430 = pi0327;
  assign po0431 = pi0328;
  assign po0433 = pi0344;
  assign po0434 = pi0346;
  assign po0435 = pi0332;
  assign po0436 = pi0342;
  assign po0437 = pi0331;
  assign po0438 = pi0333;
  assign po0439 = pi0336;
  assign po0440 = pi0334;
  assign po0441 = pi0337;
  assign po0443 = pi0338;
  assign po0444 = pi0339;
  assign po0446 = pi0343;
  assign po0447 = pi0345;
  assign po0448 = pi0350;
  assign po0449 = pi0347;
  assign po0450 = pi0348;
  assign po0451 = pi0349;
  assign po0470 = pi0351;
  assign po0482 = pi0376;
  assign po0483 = pi0386;
  assign po0484 = pi0382;
  assign po0485 = pi0395;
  assign po0486 = pi0383;
  assign po0487 = pi0384;
  assign po0488 = pi0389;
  assign po0489 = pi0387;
  assign po0490 = pi0388;
  assign po0491 = pi0391;
  assign po0492 = pi0404;
  assign po0493 = pi0408;
  assign po0494 = pi0392;
  assign po0495 = pi0394;
  assign po0496 = pi0396;
  assign po0497 = pi0393;
  assign po0498 = pi0397;
  assign po0499 = pi0399;
  assign po0500 = pi0413;
  assign po0501 = pi0400;
  assign po0502 = pi0401;
  assign po0503 = pi0402;
  assign po0504 = pi0403;
  assign po0505 = pi0405;
  assign po0507 = pi0406;
  assign po0508 = pi0407;
  assign po0509 = pi0410;
  assign po0510 = pi0409;
  assign po0511 = pi0411;
  assign po0515 = pi0412;
  assign po0520 = pi0415;
  assign po0528 = pi0414;
  assign po0546 = pi0443;
  assign po0547 = pi0455;
  assign po0548 = pi0440;
  assign po0549 = pi0442;
  assign po0550 = pi0446;
  assign po0551 = pi0448;
  assign po0552 = pi0450;
  assign po0553 = pi0451;
  assign po0554 = pi0466;
  assign po0555 = pi0467;
  assign po0556 = pi0453;
  assign po0557 = pi0460;
  assign po0558 = pi0468;
  assign po0559 = pi0463;
  assign po0560 = pi0472;
  assign po0561 = pi0457;
  assign po0562 = pi0456;
  assign po0563 = pi0459;
  assign po0564 = pi0461;
  assign po0565 = pi0462;
  assign po0566 = pi0464;
  assign po0567 = pi0465;
  assign po0568 = pi0469;
  assign po0569 = pi0470;
  assign po0571 = pi0473;
  assign po0574 = pi0474;
  assign po0575 = pi0475;
  assign po0577 = pi0476;
  assign po0579 = pi0477;
  assign po0582 = pi0478;
  assign po0584 = pi0471;
  assign po0588 = pi0479;
  assign po0610 = pi0494;
  assign po0611 = pi0520;
  assign po0612 = pi0515;
  assign po0613 = pi0524;
  assign po0614 = pi0509;
  assign po0615 = pi0510;
  assign po0616 = pi0512;
  assign po0617 = pi0517;
  assign po0618 = pi0513;
  assign po0619 = pi0514;
  assign po0620 = pi0528;
  assign po0621 = pi0518;
  assign po0622 = pi0519;
  assign po0623 = pi0521;
  assign po0625 = pi0537;
  assign po0626 = pi0525;
  assign po0627 = pi0526;
  assign po0628 = pi0527;
  assign po0629 = pi0529;
  assign po0630 = pi0530;
  assign po0631 = pi0531;
  assign po0632 = pi0540;
  assign po0633 = pi0534;
  assign po0634 = pi0533;
  assign po0635 = pi0535;
  assign po0636 = pi0532;
  assign po0637 = pi0536;
  assign po0638 = pi0539;
  assign po0641 = pi0541;
  assign po0646 = pi0542;
  assign po0652 = pi0543;
  assign po0653 = pi0538;
  assign po0674 = pi0558;
  assign po0675 = pi0575;
  assign po0676 = pi0582;
  assign po0677 = pi0572;
  assign po0678 = pi0576;
  assign po0679 = pi0577;
  assign po0680 = pi0579;
  assign po0681 = pi0584;
  assign po0682 = pi0592;
  assign po0683 = pi0581;
  assign po0684 = pi0596;
  assign po0685 = pi0583;
  assign po0686 = pi0585;
  assign po0687 = pi0586;
  assign po0689 = pi0587;
  assign po0690 = pi0588;
  assign po0691 = pi0602;
  assign po0692 = pi0590;
  assign po0693 = pi0591;
  assign po0694 = pi0605;
  assign po0695 = pi0593;
  assign po0696 = pi0594;
  assign po0697 = pi0599;
  assign po0698 = pi0606;
  assign po0699 = pi0595;
  assign po0700 = pi0597;
  assign po0701 = pi0598;
  assign po0703 = pi0600;
  assign po0704 = pi0601;
  assign po0708 = pi0604;
  assign po0710 = pi0607;
  assign po0719 = pi0603;
  assign po0738 = pi0634;
  assign po0739 = pi0646;
  assign po0740 = pi0639;
  assign po0741 = pi0651;
  assign po0742 = pi0636;
  assign po0743 = pi0638;
  assign po0744 = pi0654;
  assign po0745 = pi0648;
  assign po0746 = pi0642;
  assign po0747 = pi0643;
  assign po0748 = pi0653;
  assign po0749 = pi0644;
  assign po0750 = pi0645;
  assign po0751 = pi0647;
  assign po0752 = pi0650;
  assign po0753 = pi0664;
  assign po0754 = pi0652;
  assign po0755 = pi0656;
  assign po0756 = pi0666;
  assign po0757 = pi0655;
  assign po0758 = pi0657;
  assign po0759 = pi0658;
  assign po0760 = pi0660;
  assign po0761 = pi0661;
  assign po0762 = pi0662;
  assign po0763 = pi0668;
  assign po0765 = pi0663;
  assign po0767 = pi0667;
  assign po0770 = pi0669;
  assign po0771 = pi0670;
  assign po0779 = pi0665;
  assign po0789 = pi0671;
  assign po0802 = pi0691;
  assign po0803 = pi0703;
  assign po0804 = pi0717;
  assign po0805 = pi0704;
  assign po0806 = pi0710;
  assign po0807 = pi0718;
  assign po0808 = pi0705;
  assign po0809 = pi0706;
  assign po0810 = pi0723;
  assign po0811 = pi0708;
  assign po0812 = pi0709;
  assign po0813 = pi0711;
  assign po0814 = pi0712;
  assign po0815 = pi0713;
  assign po0816 = pi0728;
  assign po0817 = pi0715;
  assign po0818 = pi0716;
  assign po0819 = pi0719;
  assign po0820 = pi0720;
  assign po0822 = pi0721;
  assign po0823 = pi0722;
  assign po0824 = pi0724;
  assign po0825 = pi0725;
  assign po0826 = pi0726;
  assign po0827 = pi0727;
  assign po0828 = pi0729;
  assign po0829 = pi0731;
  assign po0830 = pi0730;
  assign po0831 = pi0734;
  assign po0832 = pi0735;
  assign po0837 = pi0732;
  assign po0844 = pi0733;
  assign po0866 = pi0745;
  assign po0867 = pi0772;
  assign po0868 = pi0762;
  assign po0869 = pi0766;
  assign po0870 = pi0774;
  assign po0871 = pi0781;
  assign po0872 = pi0771;
  assign po0873 = pi0778;
  assign po0874 = pi0773;
  assign po0876 = pi0775;
  assign po0877 = pi0791;
  assign po0878 = pi0776;
  assign po0879 = pi0777;
  assign po0880 = pi0779;
  assign po0881 = pi0780;
  assign po0882 = pi0782;
  assign po0883 = pi0797;
  assign po0884 = pi0784;
  assign po0885 = pi0785;
  assign po0886 = pi0786;
  assign po0887 = pi0787;
  assign po0888 = pi0788;
  assign po0889 = pi0789;
  assign po0890 = pi0790;
  assign po0891 = pi0792;
  assign po0893 = pi0794;
  assign po0894 = pi0795;
  assign po0895 = pi0793;
  assign po0897 = pi0796;
  assign po0898 = pi0783;
  assign po0899 = pi0798;
  assign po0900 = pi0799;
  assign po0930 = pi0819;
  assign po0931 = pi0826;
  assign po0932 = pi0828;
  assign po0933 = pi0842;
  assign po0934 = pi0835;
  assign po0935 = pi0834;
  assign po0936 = pi0840;
  assign po0937 = pi0848;
  assign po0938 = pi0836;
  assign po0939 = pi0837;
  assign po0940 = pi0845;
  assign po0941 = pi0838;
  assign po0942 = pi0839;
  assign po0943 = pi0841;
  assign po0944 = pi0843;
  assign po0945 = pi0844;
  assign po0946 = pi0858;
  assign po0947 = pi0861;
  assign po0948 = pi0847;
  assign po0950 = pi0849;
  assign po0951 = pi0850;
  assign po0952 = pi0851;
  assign po0953 = pi0852;
  assign po0954 = pi0853;
  assign po0955 = pi0854;
  assign po0957 = pi0855;
  assign po0959 = pi0863;
  assign po0960 = pi0856;
  assign po0961 = pi0857;
  assign po0962 = pi0859;
  assign po0963 = pi0860;
  assign po0976 = pi0862;
  assign po0994 = pi0891;
  assign po0995 = pi0905;
  assign po0996 = pi0890;
  assign po0997 = pi0893;
  assign po0998 = pi0904;
  assign po0999 = pi0895;
  assign po1000 = pi0897;
  assign po1001 = pi0896;
  assign po1002 = pi0899;
  assign po1003 = pi0901;
  assign po1004 = pi0898;
  assign po1005 = pi0909;
  assign po1006 = pi0916;
  assign po1007 = pi0918;
  assign po1008 = pi0903;
  assign po1009 = pi0920;
  assign po1010 = pi0906;
  assign po1011 = pi0907;
  assign po1012 = pi0910;
  assign po1013 = pi0911;
  assign po1014 = pi0912;
  assign po1015 = pi0914;
  assign po1016 = pi0915;
  assign po1017 = pi0917;
  assign po1018 = pi0921;
  assign po1019 = pi0922;
  assign po1022 = pi0923;
  assign po1024 = pi0924;
  assign po1030 = pi0925;
  assign po1032 = pi0919;
  assign po1038 = pi0926;
  assign po1043 = pi0927;
  assign po1058 = pi0945;
  assign po1059 = pi0967;
  assign po1060 = pi0953;
  assign po1061 = pi0954;
  assign po1062 = pi0961;
  assign po1063 = pi0968;
  assign po1064 = pi0958;
  assign po1065 = pi0962;
  assign po1066 = pi0963;
  assign po1067 = pi0972;
  assign po1068 = pi0977;
  assign po1069 = pi0964;
  assign po1070 = pi0969;
  assign po1071 = pi0970;
  assign po1072 = pi0971;
  assign po1073 = pi0973;
  assign po1074 = pi0985;
  assign po1076 = pi0979;
  assign po1077 = pi0974;
  assign po1078 = pi0975;
  assign po1079 = pi0976;
  assign po1080 = pi0978;
  assign po1081 = pi0988;
  assign po1082 = pi0981;
  assign po1085 = pi0982;
  assign po1086 = pi0983;
  assign po1087 = pi0984;
  assign po1089 = pi0986;
  assign po1090 = pi0987;
  assign po1095 = pi0989;
  assign po1096 = pi0990;
  assign po1110 = pi0991;
  assign po1122 = pi0995;
  assign po1123 = pi0999;
  assign po1124 = pi1003;
  assign po1126 = pi1198;
  assign po1128 = pi1009;
  assign po1129 = pi1013;
  assign po1130 = pi1015;
  assign po1131 = pi1203;
  assign po1134 = pi1016;
  assign po1135 = pi1023;
  assign po1136 = pi1022;
  assign po1137 = pi1189;
  assign po1140 = pi1026;
  assign po1141 = pi1031;
  assign po1142 = pi1028;
  assign po1143 = pi1029;
  assign po1144 = pi1030;
  assign po1145 = pi1195;
  assign po1148 = pi1032;
  assign po1149 = pi1034;
  assign po1150 = pi1033;
  assign po1152 = pi1038;
  assign po1153 = pi1197;
  assign po1156 = pi1204;
  assign po1159 = pi1043;
  assign po1160 = pi1045;
  assign po1161 = pi1041;
  assign po1162 = pi1042;
  assign po1163 = pi1044;
  assign po1165 = pi1215;
  assign po1168 = pi1047;
  assign po1169 = pi1048;
  assign po1170 = pi1185;
  assign po1173 = pi1049;
  assign po1174 = pi1191;
  assign po1177 = pi1187;
  assign po1180 = pi1188;
  assign po1183 = pi1194;
  assign po1186 = pi1190;
  assign po1189 = pi1211;
  assign po1192 = pi1218;
  assign po1195 = pi1052;
  assign po1196 = pi1051;
  assign po1197 = pi1050;
  assign po1198 = pi1228;
  assign po1201 = pi1053;
  assign po1202 = pi1054;
  assign po1203 = pi1207;
  assign po1206 = pi1199;
  assign po1209 = pi1186;
  assign po1212 = pi1196;
  assign po1215 = pi1205;
  assign po1218 = pi1055;
  assign po1219 = pi1201;
  assign po1222 = pi1233;
  assign po1225 = pi1184;
  assign po1229 = pi1202;
  assign po1232 = pi1192;
  assign po1236 = pi1193;
  assign po1239 = pi1212;
  assign po1242 = pi1082;
  assign po1243 = pi1080;
  assign po1244 = pi1089;
  assign po1245 = pi1074;
  assign po1246 = pi1073;
  assign po1247 = pi1083;
  assign po1248 = pi1092;
  assign po1249 = pi1099;
  assign po1250 = pi1110;
  assign po1251 = pi1094;
  assign po1252 = pi1095;
  assign po1253 = pi1098;
  assign po1254 = pi1102;
  assign po1255 = pi1122;
  assign po1256 = pi1103;
  assign po1257 = pi1104;
  assign po1258 = pi1105;
  assign po1259 = pi1090;
  assign po1260 = pi1091;
  assign po1261 = pi1109;
  assign po1262 = pi1111;
  assign po1263 = pi1114;
  assign po1264 = pi1115;
  assign po1265 = pi1116;
  assign po1266 = pi1097;
  assign po1267 = pi1117;
  assign po1268 = pi1101;
  assign po1269 = pi1100;
  assign po1270 = pi1120;
  assign po1271 = pi1121;
  assign po1272 = pi1127;
  assign po1273 = pi1128;
  assign po1274 = pi1129;
  assign po1275 = pi1106;
  assign po1276 = pi1130;
  assign po1277 = pi1131;
  assign po1278 = pi1108;
  assign po1279 = pi1133;
  assign po1280 = pi1112;
  assign po1281 = pi1113;
  assign po1282 = pi1136;
  assign po1283 = pi1155;
  assign po1284 = pi1118;
  assign po1285 = pi1119;
  assign po1286 = pi1161;
  assign po1287 = pi1159;
  assign po1288 = pi1123;
  assign po1289 = pi1124;
  assign po1290 = pi1125;
  assign po1291 = pi1126;
  assign po1292 = pi1146;
  assign po1293 = pi1150;
  assign po1294 = pi1151;
  assign po1295 = pi1132;
  assign po1296 = pi1134;
  assign po1297 = pi1135;
  assign po1299 = pi1173;
  assign po1300 = pi1138;
  assign po1301 = pi1137;
  assign po1302 = pi1139;
  assign po1303 = pi1140;
  assign po1304 = pi1169;
  assign po1305 = pi1158;
  assign po1306 = pi1142;
  assign po1307 = pi1143;
  assign po1308 = pi1144;
  assign po1309 = pi1177;
  assign po1310 = pi1166;
  assign po1312 = pi1167;
  assign po1313 = pi1147;
  assign po1314 = pi1148;
  assign po1315 = pi1149;
  assign po1319 = pi1152;
  assign po1320 = pi1171;
  assign po1321 = pi1154;
  assign po1322 = pi1156;
  assign po1323 = pi1157;
  assign po1324 = pi1176;
  assign po1325 = pi1175;
  assign po1326 = pi1160;
  assign po1327 = pi1162;
  assign po1328 = pi1164;
  assign po1329 = pi1165;
  assign po1330 = pi1178;
  assign po1333 = pi1168;
  assign po1334 = pi1180;
  assign po1336 = pi1170;
  assign po1338 = pi1172;
  assign po1348 = pi1179;
  assign po1356 = pi1182;
  assign po1365 = pi1183;
  assign po1370 = pi1200;
  assign po1371 = pi1206;
  assign po1372 = pi1208;
  assign po1373 = pi1209;
  assign po1374 = pi1210;
  assign po1375 = pi1216;
  assign po1376 = pi1219;
  assign po1377 = pi1220;
  assign po1378 = pi1235;
  assign po1379 = pi1226;
  assign po1380 = pi1224;
  assign po1381 = pi1225;
  assign po1382 = pi1229;
  assign po1383 = pi1230;
  assign po1384 = pi1214;
  assign po1385 = pi1217;
  assign po1387 = pi1234;
  assign po1388 = pi1236;
  assign po1389 = pi1222;
  assign po1390 = pi1223;
  assign po1391 = pi1238;
  assign po1393 = pi1239;
  assign po1397 = pi1242;
  assign po1398 = pi1243;
  assign po1399 = pi1231;
  assign po1401 = pi1245;
  assign po1404 = pi1246;
  assign po1407 = pi1237;
  assign po1413 = pi1240;
  assign po1414 = pi1241;
  assign po1418 = pi1244;
  assign po1419 = pi1247;
  assign po1434 = pi1259;
  assign po1435 = pi1271;
  assign po1436 = pi1268;
  assign po1437 = pi1279;
  assign po1438 = pi1291;
  assign po1439 = pi1275;
  assign po1440 = pi1287;
  assign po1441 = pi1281;
  assign po1442 = pi1280;
  assign po1443 = pi1299;
  assign po1444 = pi1289;
  assign po1446 = pi1294;
  assign po1447 = pi1277;
  assign po1448 = pi1295;
  assign po1449 = pi1296;
  assign po1450 = pi1298;
  assign po1451 = pi1297;
  assign po1452 = pi1290;
  assign po1453 = pi1300;
  assign po1455 = pi1302;
  assign po1456 = pi1288;
  assign po1458 = pi1293;
  assign po1459 = pi1304;
  assign po1460 = pi1305;
  assign po1462 = pi1306;
  assign po1464 = pi1307;
  assign po1468 = pi1308;
  assign po1469 = pi1309;
  assign po1470 = pi1310;
  assign po1471 = pi1301;
  assign po1472 = pi1303;
  assign po1478 = pi1311;
  assign po1498 = pi1335;
  assign po1499 = pi1334;
  assign po1500 = pi1339;
  assign po1501 = pi1352;
  assign po1502 = pi1341;
  assign po1503 = pi1350;
  assign po1504 = pi1345;
  assign po1505 = pi1346;
  assign po1506 = pi1351;
  assign po1507 = pi1353;
  assign po1508 = pi1355;
  assign po1509 = pi1356;
  assign po1510 = pi1371;
  assign po1511 = pi1357;
  assign po1512 = pi1372;
  assign po1513 = pi1343;
  assign po1514 = pi1358;
  assign po1515 = pi1360;
  assign po1516 = pi1359;
  assign po1517 = pi1362;
  assign po1518 = pi1363;
  assign po1519 = pi1364;
  assign po1522 = pi1365;
  assign po1523 = pi1367;
  assign po1524 = pi1368;
  assign po1526 = pi1369;
  assign po1528 = pi1373;
  assign po1530 = pi1361;
  assign po1533 = pi1374;
  assign po1534 = pi1375;
  assign po1535 = pi1366;
  assign po1540 = pi1370;
  assign po1562 = pi1395;
  assign po1563 = pi1400;
  assign po1564 = pi1404;
  assign po1565 = pi1415;
  assign po1566 = pi1420;
  assign po1567 = pi1406;
  assign po1568 = pi1410;
  assign po1569 = pi1411;
  assign po1570 = pi1413;
  assign po1571 = pi1412;
  assign po1572 = pi1414;
  assign po1573 = pi1416;
  assign po1574 = pi1426;
  assign po1575 = pi1418;
  assign po1576 = pi1419;
  assign po1577 = pi1421;
  assign po1578 = pi1405;
  assign po1579 = pi1422;
  assign po1580 = pi1423;
  assign po1582 = pi1424;
  assign po1583 = pi1433;
  assign po1584 = pi1427;
  assign po1585 = pi1428;
  assign po1587 = pi1429;
  assign po1588 = pi1431;
  assign po1589 = pi1432;
  assign po1593 = pi1434;
  assign po1594 = pi1435;
  assign po1595 = pi1436;
  assign po1603 = pi1430;
  assign po1611 = pi1438;
  assign po1623 = pi1439;
  assign po1626 = pi1473;
  assign po1627 = pi1464;
  assign po1628 = pi1463;
  assign po1629 = pi1467;
  assign po1630 = pi1470;
  assign po1631 = pi1469;
  assign po1632 = pi1476;
  assign po1633 = pi1480;
  assign po1634 = pi1482;
  assign po1635 = pi1475;
  assign po1636 = pi1477;
  assign po1637 = pi1478;
  assign po1638 = pi1481;
  assign po1639 = pi1483;
  assign po1640 = pi1484;
  assign po1641 = pi1485;
  assign po1642 = pi1486;
  assign po1643 = pi1487;
  assign po1644 = pi1488;
  assign po1645 = pi1489;
  assign po1646 = pi1497;
  assign po1647 = pi1490;
  assign po1648 = pi1491;
  assign po1651 = pi1493;
  assign po1652 = pi1494;
  assign po1654 = pi1495;
  assign po1657 = pi1499;
  assign po1658 = pi1500;
  assign po1660 = pi1501;
  assign po1665 = pi1496;
  assign po1678 = pi1502;
  assign po1684 = pi1503;
  assign po1690 = pi1524;
  assign po1691 = pi1528;
  assign po1692 = pi1529;
  assign po1693 = pi1545;
  assign po1694 = pi1534;
  assign po1695 = pi1535;
  assign po1696 = pi1536;
  assign po1697 = pi1538;
  assign po1698 = pi1539;
  assign po1699 = pi1544;
  assign po1700 = pi1546;
  assign po1701 = pi1548;
  assign po1702 = pi1541;
  assign po1703 = pi1551;
  assign po1704 = pi1542;
  assign po1705 = pi1547;
  assign po1706 = pi1550;
  assign po1707 = pi1549;
  assign po1708 = pi1552;
  assign po1709 = pi1565;
  assign po1711 = pi1554;
  assign po1712 = pi1555;
  assign po1713 = pi1556;
  assign po1716 = pi1564;
  assign po1717 = pi1559;
  assign po1718 = pi1561;
  assign po1719 = pi1560;
  assign po1723 = pi1562;
  assign po1726 = pi1563;
  assign po1729 = pi1558;
  assign po1739 = pi1566;
  assign po1743 = pi1567;
  assign po1754 = pi1591;
  assign po1755 = pi1600;
  assign po1756 = pi1593;
  assign po1757 = pi1598;
  assign po1758 = pi1614;
  assign po1759 = pi1599;
  assign po1760 = pi1618;
  assign po1761 = pi1603;
  assign po1762 = pi1605;
  assign po1763 = pi1608;
  assign po1764 = pi1607;
  assign po1765 = pi1609;
  assign po1766 = pi1610;
  assign po1767 = pi1611;
  assign po1768 = pi1612;
  assign po1769 = pi1615;
  assign po1770 = pi1613;
  assign po1771 = pi1622;
  assign po1772 = pi1616;
  assign po1773 = pi1617;
  assign po1774 = pi1604;
  assign po1775 = pi1620;
  assign po1776 = pi1621;
  assign po1778 = pi1623;
  assign po1780 = pi1628;
  assign po1781 = pi1626;
  assign po1782 = pi1624;
  assign po1783 = pi1627;
  assign po1787 = pi1629;
  assign po1788 = pi1630;
  assign po1792 = pi1625;
  assign po1805 = pi1631;
  assign po1818 = pi1662;
  assign po1819 = pi1672;
  assign po1820 = pi1657;
  assign po1821 = pi1652;
  assign po1822 = pi1663;
  assign po1823 = pi1664;
  assign po1824 = pi1665;
  assign po1825 = pi1667;
  assign po1826 = pi1659;
  assign po1827 = pi1661;
  assign po1828 = pi1670;
  assign po1829 = pi1677;
  assign po1830 = pi1669;
  assign po1831 = pi1676;
  assign po1832 = pi1668;
  assign po1833 = pi1678;
  assign po1834 = pi1679;
  assign po1835 = pi1690;
  assign po1836 = pi1684;
  assign po1837 = pi1685;
  assign po1839 = pi1689;
  assign po1840 = pi1687;
  assign po1841 = pi1688;
  assign po1842 = pi1675;
  assign po1844 = pi1683;
  assign po1846 = pi1680;
  assign po1852 = pi1691;
  assign po1857 = pi1686;
  assign po1859 = pi1693;
  assign po1860 = pi1694;
  assign po1867 = pi1695;
  assign po1868 = pi1692;
  assign po1882 = pi1702;
  assign po1883 = pi1709;
  assign po1884 = pi1723;
  assign po1885 = pi1724;
  assign po1886 = pi1732;
  assign po1887 = pi1725;
  assign po1889 = pi1731;
  assign po1890 = pi1734;
  assign po1891 = pi1742;
  assign po1892 = pi1736;
  assign po1893 = pi1743;
  assign po1894 = pi1738;
  assign po1896 = pi1739;
  assign po1897 = pi1744;
  assign po1898 = pi1741;
  assign po1899 = pi1728;
  assign po1900 = pi1745;
  assign po1901 = pi1746;
  assign po1902 = pi1747;
  assign po1903 = pi1748;
  assign po1904 = pi1749;
  assign po1905 = pi1755;
  assign po1906 = pi1740;
  assign po1907 = pi1750;
  assign po1908 = pi1751;
  assign po1912 = pi1752;
  assign po1913 = pi1753;
  assign po1915 = pi1754;
  assign po1916 = pi1756;
  assign po1919 = pi1757;
  assign po1921 = pi1758;
  assign po1923 = pi1759;
  assign po1946 = pi1775;
  assign po1947 = pi1785;
  assign po1948 = pi1786;
  assign po1949 = pi1787;
  assign po1950 = pi1791;
  assign po1951 = pi1792;
  assign po1952 = pi1799;
  assign po1953 = pi1794;
  assign po1954 = pi1804;
  assign po1955 = pi1812;
  assign po1956 = pi1798;
  assign po1957 = pi1800;
  assign po1958 = pi1802;
  assign po1959 = pi1801;
  assign po1960 = pi1806;
  assign po1962 = pi1803;
  assign po1963 = pi1805;
  assign po1964 = pi1807;
  assign po1965 = pi1808;
  assign po1966 = pi1809;
  assign po1967 = pi1811;
  assign po1968 = pi1813;
  assign po1969 = pi1797;
  assign po1970 = pi1815;
  assign po1974 = pi1820;
  assign po1975 = pi1816;
  assign po1976 = pi1817;
  assign po1979 = pi1818;
  assign po1981 = pi1821;
  assign po1982 = pi1822;
  assign po1996 = pi1819;
  assign po2000 = pi1823;
  assign po2010 = pi1843;
  assign po2011 = pi1849;
  assign po2012 = pi1848;
  assign po2013 = pi1855;
  assign po2014 = pi1860;
  assign po2015 = pi1857;
  assign po2016 = pi1861;
  assign po2017 = pi1856;
  assign po2018 = pi1858;
  assign po2019 = pi1874;
  assign po2020 = pi1868;
  assign po2021 = pi1862;
  assign po2022 = pi1864;
  assign po2023 = pi1866;
  assign po2024 = pi1869;
  assign po2025 = pi1854;
  assign po2026 = pi1872;
  assign po2027 = pi1871;
  assign po2028 = pi1873;
  assign po2030 = pi1875;
  assign po2031 = pi1876;
  assign po2032 = pi1877;
  assign po2033 = pi1878;
  assign po2036 = pi1879;
  assign po2037 = pi1881;
  assign po2038 = pi1882;
  assign po2039 = pi1883;
  assign po2045 = pi1885;
  assign po2049 = pi1880;
  assign po2051 = pi1886;
  assign po2053 = pi1887;
  assign po2056 = pi1884;
  assign po2074 = pi1900;
  assign po2075 = pi1906;
  assign po2076 = pi1919;
  assign po2077 = pi1920;
  assign po2078 = pi1926;
  assign po2079 = pi1922;
  assign po2080 = pi1924;
  assign po2081 = pi1923;
  assign po2082 = pi1928;
  assign po2083 = pi1925;
  assign po2084 = pi1927;
  assign po2085 = pi1929;
  assign po2087 = pi1937;
  assign po2088 = pi1932;
  assign po2089 = pi1938;
  assign po2090 = pi1934;
  assign po2091 = pi1935;
  assign po2093 = pi1936;
  assign po2094 = pi1939;
  assign po2095 = pi1940;
  assign po2096 = pi1941;
  assign po2097 = pi1942;
  assign po2098 = pi1943;
  assign po2099 = pi1944;
  assign po2100 = pi1945;
  assign po2101 = pi1933;
  assign po2102 = pi1946;
  assign po2103 = pi1947;
  assign po2104 = pi1948;
  assign po2107 = pi1949;
  assign po2116 = pi1950;
  assign po2117 = pi1951;
  assign po2138 = pi1983;
  assign po2139 = pi1978;
  assign po2140 = pi1974;
  assign po2141 = pi1990;
  assign po2142 = pi1975;
  assign po2143 = pi1972;
  assign po2144 = pi1989;
  assign po2145 = pi1982;
  assign po2146 = pi1985;
  assign po2147 = pi1991;
  assign po2148 = pi1981;
  assign po2149 = pi1997;
  assign po2150 = pi1993;
  assign po2151 = pi1992;
  assign po2152 = pi2000;
  assign po2153 = pi1999;
  assign po2154 = pi2001;
  assign po2155 = pi1998;
  assign po2156 = pi2002;
  assign po2157 = pi2005;
  assign po2159 = pi2003;
  assign po2162 = pi2013;
  assign po2163 = pi2004;
  assign po2165 = pi2006;
  assign po2166 = pi2007;
  assign po2170 = pi2010;
  assign po2172 = pi2011;
  assign po2173 = pi2012;
  assign po2174 = pi2008;
  assign po2180 = pi2015;
  assign po2181 = pi2014;
  assign po2182 = pi2009;
  assign po2202 = pi2032;
  assign po2203 = pi2043;
  assign po2204 = pi2037;
  assign po2205 = pi2036;
  assign po2206 = pi2056;
  assign po2207 = pi2045;
  assign po2208 = pi2055;
  assign po2209 = pi2049;
  assign po2210 = pi2054;
  assign po2211 = pi2052;
  assign po2212 = pi2069;
  assign po2213 = pi2058;
  assign po2214 = pi2061;
  assign po2215 = pi2059;
  assign po2216 = pi2060;
  assign po2217 = pi2065;
  assign po2219 = pi2072;
  assign po2220 = pi2074;
  assign po2221 = pi2067;
  assign po2224 = pi2066;
  assign po2225 = pi2053;
  assign po2226 = pi2073;
  assign po2227 = pi2077;
  assign po2228 = pi2068;
  assign po2230 = pi2062;
  assign po2232 = pi2064;
  assign po2233 = pi2070;
  assign po2234 = pi2075;
  assign po2236 = pi2076;
  assign po2237 = pi2078;
  assign po2243 = pi2079;
  assign po2249 = pi2071;
  assign po2266 = pi2083;
  assign po2267 = pi2089;
  assign po2268 = pi2100;
  assign po2269 = pi2303;
  assign po2272 = pi2102;
  assign po2273 = pi2106;
  assign po2274 = pi2107;
  assign po2275 = pi2108;
  assign po2276 = pi2109;
  assign po2277 = pi2290;
  assign po2280 = pi2115;
  assign po2281 = pi2114;
  assign po2282 = pi2117;
  assign po2283 = pi2110;
  assign po2284 = pi2118;
  assign po2285 = pi2120;
  assign po2286 = pi2122;
  assign po2287 = pi2111;
  assign po2288 = pi2123;
  assign po2289 = pi2124;
  assign po2290 = pi2279;
  assign po2293 = pi2128;
  assign po2294 = pi2302;
  assign po2297 = pi2132;
  assign po2298 = pi2129;
  assign po2299 = pi2133;
  assign po2300 = pi2309;
  assign po2303 = pi2277;
  assign po2306 = pi2299;
  assign po2311 = pi2294;
  assign po2314 = pi2135;
  assign po2315 = pi2136;
  assign po2316 = pi2286;
  assign po2319 = pi2317;
  assign po2322 = pi2139;
  assign po2324 = pi2285;
  assign po2326 = pi2278;
  assign po2329 = pi2134;
  assign po2330 = pi2293;
  assign po2333 = pi2137;
  assign po2334 = pi2287;
  assign po2338 = pi2274;
  assign po2340 = pi2284;
  assign po2343 = pi2141;
  assign po2344 = pi2138;
  assign po2345 = pi2140;
  assign po2347 = pi2300;
  assign po2350 = pi2143;
  assign po2351 = pi2142;
  assign po2353 = pi2283;
  assign po2356 = pi2273;
  assign po2359 = pi2292;
  assign po2363 = pi2280;
  assign po2371 = pi2282;
  assign po2374 = pi2159;
  assign po2375 = pi2162;
  assign po2376 = pi2158;
  assign po2377 = pi2160;
  assign po2378 = pi2178;
  assign po2379 = pi2164;
  assign po2380 = pi2185;
  assign po2381 = pi2168;
  assign po2382 = pi2174;
  assign po2383 = pi2176;
  assign po2384 = pi2199;
  assign po2385 = pi2183;
  assign po2386 = pi2184;
  assign po2387 = pi2182;
  assign po2388 = pi2167;
  assign po2389 = pi2166;
  assign po2390 = pi2170;
  assign po2391 = pi2192;
  assign po2392 = pi2175;
  assign po2393 = pi2189;
  assign po2394 = pi2181;
  assign po2395 = pi2196;
  assign po2396 = pi2222;
  assign po2397 = pi2206;
  assign po2398 = pi2187;
  assign po2399 = pi2209;
  assign po2401 = pi2210;
  assign po2402 = pi2211;
  assign po2403 = pi2212;
  assign po2404 = pi2190;
  assign po2405 = pi2227;
  assign po2406 = pi2193;
  assign po2407 = pi2221;
  assign po2408 = pi2194;
  assign po2409 = pi2215;
  assign po2410 = pi2208;
  assign po2411 = pi2217;
  assign po2412 = pi2207;
  assign po2413 = pi2202;
  assign po2414 = pi2203;
  assign po2415 = pi2204;
  assign po2416 = pi2224;
  assign po2418 = pi2225;
  assign po2419 = pi2214;
  assign po2420 = pi2230;
  assign po2421 = pi2229;
  assign po2422 = pi2213;
  assign po2423 = pi2233;
  assign po2424 = pi2234;
  assign po2425 = pi2242;
  assign po2426 = pi2220;
  assign po2427 = pi2243;
  assign po2429 = pi2219;
  assign po2430 = pi2218;
  assign po2431 = pi2244;
  assign po2432 = pi2223;
  assign po2433 = pi2241;
  assign po2434 = pi2246;
  assign po2435 = pi2238;
  assign po2437 = pi2240;
  assign po2438 = pi2236;
  assign po2439 = pi2228;
  assign po2440 = pi2226;
  assign po2441 = pi2231;
  assign po2442 = pi2232;
  assign po2443 = pi2254;
  assign po2445 = pi2235;
  assign po2448 = pi2239;
  assign po2449 = pi2258;
  assign po2450 = pi2245;
  assign po2451 = pi2237;
  assign po2454 = pi2248;
  assign po2455 = pi2249;
  assign po2456 = pi2253;
  assign po2458 = pi2251;
  assign po2459 = pi2250;
  assign po2461 = pi2262;
  assign po2462 = pi2252;
  assign po2465 = pi2255;
  assign po2466 = pi2264;
  assign po2467 = pi2271;
  assign po2468 = pi2260;
  assign po2472 = pi2256;
  assign po2473 = pi2257;
  assign po2474 = pi2259;
  assign po2478 = pi2266;
  assign po2479 = pi2261;
  assign po2486 = pi2267;
  assign po2487 = pi2268;
  assign po2490 = pi2265;
  assign po2502 = pi2275;
  assign po2503 = pi2295;
  assign po2504 = pi2296;
  assign po2506 = pi2304;
  assign po2507 = pi2305;
  assign po2508 = pi2291;
  assign po2509 = pi2310;
  assign po2510 = pi2312;
  assign po2511 = pi2313;
  assign po2512 = pi2308;
  assign po2513 = pi2314;
  assign po2514 = pi2301;
  assign po2515 = pi2298;
  assign po2516 = pi2316;
  assign po2517 = pi2320;
  assign po2518 = pi2307;
  assign po2519 = pi2315;
  assign po2520 = pi2328;
  assign po2522 = pi2326;
  assign po2523 = pi2324;
  assign po2524 = pi2327;
  assign po2527 = pi2322;
  assign po2529 = pi2334;
  assign po2530 = pi2318;
  assign po2532 = pi2319;
  assign po2533 = pi2333;
  assign po2536 = pi2329;
  assign po2539 = pi2325;
  assign po2541 = pi2323;
  assign po2547 = pi2332;
  assign po2551 = pi2330;
  assign po2561 = pi2335;
  assign po2566 = pi2346;
  assign po2567 = pi2360;
  assign po2568 = pi2352;
  assign po2569 = pi2355;
  assign po2570 = pi2370;
  assign po2571 = pi2364;
  assign po2572 = pi2365;
  assign po2573 = pi2376;
  assign po2574 = pi2367;
  assign po2575 = pi2366;
  assign po2577 = pi2371;
  assign po2578 = pi2377;
  assign po2579 = pi2381;
  assign po2580 = pi2385;
  assign po2581 = pi2380;
  assign po2583 = pi2379;
  assign po2584 = pi2384;
  assign po2586 = pi2383;
  assign po2587 = pi2392;
  assign po2588 = pi2388;
  assign po2589 = pi2387;
  assign po2591 = pi2389;
  assign po2592 = pi2390;
  assign po2593 = pi2386;
  assign po2598 = pi2397;
  assign po2599 = pi2394;
  assign po2602 = pi2395;
  assign po2603 = pi2393;
  assign po2604 = pi2391;
  assign po2605 = pi2398;
  assign po2608 = pi2396;
  assign po2612 = pi2399;
  assign po2630 = pi2424;
  assign po2631 = pi2417;
  assign po2632 = pi2423;
  assign po2633 = pi2421;
  assign po2634 = pi2435;
  assign po2635 = pi2426;
  assign po2636 = pi2428;
  assign po2637 = pi2429;
  assign po2638 = pi2437;
  assign po2639 = pi2439;
  assign po2640 = pi2432;
  assign po2641 = pi2433;
  assign po2642 = pi2440;
  assign po2643 = pi2434;
  assign po2644 = pi2438;
  assign po2645 = pi2447;
  assign po2646 = pi2448;
  assign po2648 = pi2444;
  assign po2649 = pi2430;
  assign po2650 = pi2453;
  assign po2652 = pi2450;
  assign po2655 = pi2452;
  assign po2657 = pi2442;
  assign po2661 = pi2456;
  assign po2666 = pi2454;
  assign po2671 = pi2457;
  assign po2673 = pi2458;
  assign po2675 = pi2461;
  assign po2676 = pi2459;
  assign po2679 = pi2462;
  assign po2681 = pi2455;
  assign po2690 = pi2463;
  assign po2694 = pi2469;
  assign po2695 = pi2472;
  assign po2696 = pi2482;
  assign po2697 = pi2493;
  assign po2698 = pi2481;
  assign po2700 = pi2499;
  assign po2701 = pi2487;
  assign po2703 = pi2504;
  assign po2705 = pi2508;
  assign po2706 = pi2505;
  assign po2707 = pi2510;
  assign po2708 = pi2491;
  assign po2709 = pi2506;
  assign po2710 = pi2511;
  assign po2713 = pi2512;
  assign po2714 = pi2507;
  assign po2715 = pi2515;
  assign po2716 = pi2514;
  assign po2718 = pi2518;
  assign po2719 = pi2513;
  assign po2720 = pi2516;
  assign po2722 = pi2519;
  assign po2724 = pi2526;
  assign po2725 = pi2517;
  assign po2726 = pi2520;
  assign po2727 = pi2522;
  assign po2730 = pi2523;
  assign po2731 = pi2524;
  assign po2732 = pi2521;
  assign po2733 = pi2525;
  assign po2739 = pi2527;
  assign po2758 = pi2537;
  assign po2759 = pi2564;
  assign po2760 = pi2548;
  assign po2761 = pi2557;
  assign po2762 = pi2560;
  assign po2763 = pi2554;
  assign po2764 = pi2559;
  assign po2765 = pi2561;
  assign po2766 = pi2563;
  assign po2768 = pi2565;
  assign po2769 = pi2566;
  assign po2770 = pi2569;
  assign po2771 = pi2571;
  assign po2772 = pi2570;
  assign po2773 = pi2575;
  assign po2774 = pi2558;
  assign po2775 = pi2572;
  assign po2776 = pi2578;
  assign po2777 = pi2579;
  assign po2779 = pi2587;
  assign po2780 = pi2577;
  assign po2781 = pi2576;
  assign po2782 = pi2582;
  assign po2783 = pi2580;
  assign po2785 = pi2583;
  assign po2786 = pi2581;
  assign po2792 = pi2584;
  assign po2797 = pi2585;
  assign po2798 = pi2586;
  assign po2803 = pi2589;
  assign po2804 = pi2591;
  assign po2818 = pi2590;
  assign po2822 = pi2613;
  assign po2823 = pi2610;
  assign po2824 = pi2616;
  assign po2825 = pi2636;
  assign po2826 = pi2617;
  assign po2827 = pi2630;
  assign po2828 = pi2624;
  assign po2829 = pi2626;
  assign po2830 = pi2629;
  assign po2831 = pi2638;
  assign po2832 = pi2625;
  assign po2833 = pi2637;
  assign po2834 = pi2628;
  assign po2835 = pi2631;
  assign po2836 = pi2639;
  assign po2837 = pi2633;
  assign po2838 = pi2632;
  assign po2839 = pi2634;
  assign po2841 = pi2640;
  assign po2842 = pi2644;
  assign po2844 = pi2642;
  assign po2845 = pi2643;
  assign po2848 = pi2646;
  assign po2849 = pi2647;
  assign po2850 = pi2649;
  assign po2851 = pi2650;
  assign po2852 = pi2648;
  assign po2853 = pi2645;
  assign po2857 = pi2651;
  assign po2865 = pi2654;
  assign po2871 = pi2653;
  assign po2882 = pi2655;
  assign po2886 = pi2668;
  assign po2887 = pi2683;
  assign po2888 = pi2674;
  assign po2889 = pi2694;
  assign po2890 = pi2684;
  assign po2891 = pi2690;
  assign po2892 = pi2695;
  assign po2893 = pi2692;
  assign po2894 = pi2691;
  assign po2895 = pi2699;
  assign po2896 = pi2686;
  assign po2897 = pi2702;
  assign po2899 = pi2701;
  assign po2900 = pi2697;
  assign po2901 = pi2700;
  assign po2902 = pi2703;
  assign po2903 = pi2705;
  assign po2905 = pi2709;
  assign po2906 = pi2707;
  assign po2907 = pi2706;
  assign po2908 = pi2708;
  assign po2909 = pi2713;
  assign po2910 = pi2710;
  assign po2911 = pi2711;
  assign po2912 = pi2712;
  assign po2915 = pi2718;
  assign po2917 = pi2715;
  assign po2918 = pi2716;
  assign po2919 = pi2719;
  assign po2923 = pi2704;
  assign po2926 = pi2717;
  assign po2928 = pi2714;
  assign po2950 = pi2738;
  assign po2951 = pi2741;
  assign po2952 = pi2753;
  assign po2953 = pi2748;
  assign po2954 = pi2757;
  assign po2955 = pi2759;
  assign po2956 = pi2739;
  assign po2957 = pi2754;
  assign po2958 = pi2755;
  assign po2959 = pi2758;
  assign po2960 = pi2765;
  assign po2961 = pi2764;
  assign po2962 = pi2766;
  assign po2963 = pi2760;
  assign po2964 = pi2769;
  assign po2965 = pi2762;
  assign po2966 = pi2768;
  assign po2967 = pi2761;
  assign po2970 = pi2776;
  assign po2972 = pi2772;
  assign po2973 = pi2771;
  assign po2974 = pi2773;
  assign po2975 = pi2775;
  assign po2976 = pi2777;
  assign po2977 = pi2770;
  assign po2979 = pi2779;
  assign po2980 = pi2780;
  assign po2981 = pi2778;
  assign po2982 = pi2767;
  assign po2986 = pi2781;
  assign po2993 = pi2783;
  assign po3004 = pi2782;
  assign po3014 = pi2802;
  assign po3015 = pi2818;
  assign po3016 = pi2812;
  assign po3017 = pi2817;
  assign po3018 = pi2832;
  assign po3019 = pi2813;
  assign po3020 = pi2820;
  assign po3021 = pi2822;
  assign po3022 = pi2823;
  assign po3023 = pi2827;
  assign po3024 = pi2826;
  assign po3025 = pi2821;
  assign po3026 = pi2824;
  assign po3027 = pi2825;
  assign po3028 = pi2831;
  assign po3029 = pi2835;
  assign po3030 = pi2834;
  assign po3031 = pi2830;
  assign po3033 = pi2833;
  assign po3034 = pi2819;
  assign po3035 = pi2839;
  assign po3036 = pi2838;
  assign po3037 = pi2828;
  assign po3038 = pi2836;
  assign po3039 = pi2837;
  assign po3040 = pi2841;
  assign po3041 = pi2842;
  assign po3044 = pi2844;
  assign po3045 = pi2846;
  assign po3046 = pi2845;
  assign po3059 = pi2840;
  assign po3073 = pi2847;
  assign po3078 = pi2868;
  assign po3079 = pi2880;
  assign po3080 = pi2882;
  assign po3081 = pi2879;
  assign po3082 = pi2872;
  assign po3083 = pi2888;
  assign po3084 = pi2881;
  assign po3085 = pi2890;
  assign po3086 = pi2878;
  assign po3087 = pi2873;
  assign po3088 = pi2885;
  assign po3089 = pi2891;
  assign po3090 = pi2901;
  assign po3091 = pi2887;
  assign po3092 = pi2886;
  assign po3093 = pi2892;
  assign po3094 = pi2894;
  assign po3095 = pi2895;
  assign po3096 = pi2904;
  assign po3097 = pi2899;
  assign po3099 = pi2897;
  assign po3100 = pi2900;
  assign po3101 = pi2896;
  assign po3104 = pi2905;
  assign po3105 = pi2906;
  assign po3106 = pi2903;
  assign po3107 = pi2907;
  assign po3113 = pi2908;
  assign po3114 = pi2910;
  assign po3119 = pi2911;
  assign po3123 = pi2902;
  assign po3128 = pi2909;
  assign po3142 = pi2930;
  assign po3143 = pi2936;
  assign po3144 = pi2938;
  assign po3145 = pi2944;
  assign po3146 = pi2941;
  assign po3147 = pi2960;
  assign po3148 = pi2961;
  assign po3149 = pi2946;
  assign po3150 = pi2937;
  assign po3151 = pi2953;
  assign po3152 = pi2954;
  assign po3153 = pi2962;
  assign po3154 = pi2945;
  assign po3155 = pi2947;
  assign po3156 = pi2952;
  assign po3157 = pi2966;
  assign po3158 = pi2959;
  assign po3159 = pi2956;
  assign po3161 = pi2967;
  assign po3162 = pi2957;
  assign po3163 = pi2949;
  assign po3164 = pi2968;
  assign po3165 = pi2964;
  assign po3169 = pi2965;
  assign po3170 = pi2970;
  assign po3172 = pi2971;
  assign po3173 = pi2969;
  assign po3178 = pi2963;
  assign po3180 = pi2972;
  assign po3181 = pi2973;
  assign po3185 = pi2974;
  assign po3188 = pi2975;
  assign po3206 = pi3035;
  assign po3207 = pi3022;
  assign po3208 = pi3023;
  assign po3209 = pi3048;
  assign po3210 = pi3029;
  assign po3211 = pi3031;
  assign po3212 = pi3050;
  assign po3213 = pi3021;
  assign po3214 = pi3041;
  assign po3215 = pi3030;
  assign po3216 = pi3020;
  assign po3217 = pi3014;
  assign po3218 = pi3017;
  assign po3219 = pi3032;
  assign po3220 = pi3013;
  assign po3221 = pi3025;
  assign po3222 = pi3012;
  assign po3223 = pi3055;
  assign po3224 = pi3015;
  assign po3225 = pi3034;
  assign po3226 = pi3026;
  assign po3227 = pi3054;
  assign po3228 = pi3037;
  assign po3229 = pi3036;
  assign po3230 = pi3049;
  assign po3231 = pi3056;
  assign po3232 = pi3027;
  assign po3233 = pi3024;
  assign po3234 = pi3018;
  assign po3235 = pi3051;
  assign po3236 = pi3039;
  assign po3237 = pi3019;
  assign po3238 = pi3052;
  assign po3239 = pi3057;
  assign po3240 = pi3061;
  assign po3241 = pi3067;
  assign po3242 = pi3086;
  assign po3243 = pi3077;
  assign po3244 = pi3094;
  assign po3245 = pi3080;
  assign po3246 = pi3065;
  assign po3247 = pi3078;
  assign po3248 = pi3070;
  assign po3249 = pi3093;
  assign po3250 = pi3111;
  assign po3251 = pi3091;
  assign po3252 = pi3108;
  assign po3253 = pi3079;
  assign po3254 = pi3071;
  assign po3255 = pi3073;
  assign po3256 = pi3082;
  assign po3257 = pi3088;
  assign po3258 = pi3060;
  assign po3259 = pi3084;
  assign po3260 = pi3069;
  assign po3261 = pi3104;
  assign po3262 = pi3083;
  assign po3263 = pi3062;
  assign po3264 = pi3109;
  assign po3265 = pi3074;
  assign po3266 = pi3075;
  assign po3267 = pi3081;
  assign po3268 = pi3059;
  assign po3269 = pi3076;
  assign po3270 = pi3095;
  assign po3271 = pi3072;
  assign po3272 = pi3097;
  assign po3273 = pi3101;
  assign po3274 = pi3100;
  assign po3275 = pi3098;
  assign po3276 = pi3096;
  assign po3277 = pi3099;
  assign po3278 = pi3107;
  assign po3279 = pi3112;
  assign po3280 = pi3085;
  assign po3281 = pi3090;
  assign po3282 = pi3087;
  assign po3283 = pi3102;
  assign po3284 = pi3089;
  assign po3285 = pi3110;
  assign po3286 = pi3092;
  assign po3287 = pi3113;
  assign po3288 = pi3114;
  assign po3289 = pi3122;
  assign po3290 = pi3115;
  assign po3291 = pi3118;
  assign po3292 = pi3116;
  assign po3293 = pi3124;
  assign po3294 = pi3123;
  assign po3295 = pi3120;
  assign po3296 = pi3126;
  assign po3297 = pi3119;
  assign po3298 = pi3127;
  assign po3299 = pi3152;
  assign po3300 = pi3158;
  assign po3301 = pi3141;
  assign po3302 = pi3154;
  assign po3303 = pi3167;
  assign po3304 = pi3148;
  assign po3305 = pi3146;
  assign po3306 = pi3136;
  assign po3307 = pi3129;
  assign po3308 = pi3142;
  assign po3309 = pi3147;
  assign po3310 = pi3139;
  assign po3311 = pi3131;
  assign po3312 = pi3135;
  assign po3313 = pi3155;
  assign po3314 = pi3134;
  assign po3315 = pi3159;
  assign po3316 = pi3156;
  assign po3317 = pi3133;
  assign po3318 = pi3128;
  assign po3319 = pi3132;
  assign po3320 = pi3166;
  assign po3321 = pi3170;
  assign po3322 = pi3161;
  assign po3323 = pi3140;
  assign po3324 = pi3149;
  assign po3325 = pi3168;
  assign po3326 = pi3157;
  assign po3327 = pi3169;
  assign po3328 = pi3163;
  assign po3329 = pi3117;
  assign po3330 = pi3160;
  assign po3331 = pi3137;
  assign po3332 = pi3121;
  assign po3333 = pi3125;
  assign po3334 = pi3130;
  assign po3335 = pi3164;
  assign po3336 = pi3165;
  assign po3337 = pi3150;
  assign po3338 = pi3151;
  assign po3339 = pi3143;
  assign po3340 = pi3145;
  assign po3341 = pi3144;
  assign po3342 = pi3138;
  assign po3343 = pi3171;
  assign po3344 = pi3172;
  assign po3345 = pi3176;
  assign po3346 = pi3179;
  assign po3347 = pi3182;
  assign po3348 = pi3177;
  assign po3349 = pi3181;
  assign po3350 = pi3183;
  assign po3351 = pi3175;
  assign po3352 = pi3178;
  assign po3353 = pi3162;
  assign po3354 = pi3180;
  assign po3355 = pi3184;
  assign po3356 = pi3153;
  assign po3357 = pi3188;
  assign po3358 = pi3219;
  assign po3359 = pi3205;
  assign po3360 = pi3213;
  assign po3361 = pi3221;
  assign po3362 = pi3199;
  assign po3363 = pi3239;
  assign po3364 = pi3197;
  assign po3365 = pi3223;
  assign po3366 = pi3214;
  assign po3367 = pi3196;
  assign po3368 = pi3202;
  assign po3369 = pi3208;
  assign po3370 = pi3229;
  assign po3371 = pi3210;
  assign po3372 = pi3201;
  assign po3373 = pi3234;
  assign po3374 = pi3204;
  assign po3375 = pi3232;
  assign po3376 = pi3207;
  assign po3377 = pi3226;
  assign po3378 = pi3209;
  assign po3379 = pi3220;
  assign po3380 = pi3230;
  assign po3381 = pi3211;
  assign po3382 = pi3218;
  assign po3383 = pi3174;
  assign po3384 = pi3200;
  assign po3385 = pi3212;
  assign po3386 = pi3233;
  assign po3387 = pi3227;
  assign po3388 = pi3215;
  assign po3389 = pi3222;
  assign po3390 = pi3235;
  assign po3391 = pi3216;
  assign po3392 = pi3224;
  assign po3393 = pi3217;
  assign po3394 = pi3225;
  assign po3395 = pi3228;
  assign po3396 = pi3206;
  assign po3397 = pi3238;
  assign po3398 = pi3198;
  assign po3399 = pi3194;
  assign po3400 = pi3203;
  assign po3401 = pi3250;
  assign po3402 = pi3240;
  assign po3403 = pi3270;
  assign po3404 = pi3258;
  assign po3405 = pi3257;
  assign po3406 = pi3255;
  assign po3407 = pi3259;
  assign po3408 = pi3263;
  assign po3409 = pi3253;
  assign po3410 = pi3251;
  assign po3411 = pi3252;
  assign po3412 = pi3256;
  assign po3413 = pi3254;
  assign po3414 = pi3195;
  assign po3415 = pi3311;
  assign po3416 = pi3310;
  assign po3417 = pi3267;
  assign po3418 = pi3246;
  assign po3419 = pi3268;
  assign po3420 = pi3269;
  assign po3421 = pi3266;
  assign po3422 = pi3265;
  assign po3423 = pi3272;
  assign po3424 = pi3302;
  assign po3425 = pi3294;
  assign po3426 = pi3295;
  assign po3427 = pi3313;
  assign po3428 = pi3290;
  assign po3429 = pi3287;
  assign po3430 = pi3317;
  assign po3431 = pi3289;
  assign po3432 = pi3318;
  assign po3433 = pi3316;
  assign po3434 = pi3279;
  assign po3435 = pi3280;
  assign po3436 = pi3274;
  assign po3437 = pi3304;
  assign po3438 = pi3291;
  assign po3439 = pi3288;
  assign po3440 = pi3319;
  assign po3441 = pi3277;
  assign po3442 = pi3306;
  assign po3443 = pi3293;
  assign po3444 = pi3285;
  assign po3445 = pi3303;
  assign po3446 = pi3312;
  assign po3447 = pi3298;
  assign po3448 = pi3284;
  assign po3449 = pi3286;
  assign po3450 = pi3281;
  assign po3451 = pi3299;
  assign po3452 = pi3275;
  assign po3453 = pi3276;
  assign po3454 = pi3307;
  assign po3455 = pi3308;
  assign po3456 = pi3297;
  assign po3457 = pi3292;
  assign po3458 = pi3296;
  assign po3459 = pi3300;
  assign po3460 = pi3315;
  assign po3461 = pi3314;
  assign po3462 = pi3283;
  assign po3463 = pi3278;
  assign po3464 = pi3305;
  assign po3465 = pi3282;
  assign po3466 = pi3324;
  assign po3467 = pi3309;
  assign po3468 = pi3320;
  assign po3469 = pi3301;
  assign po3470 = pi3322;
  assign po3471 = pi3346;
  assign po3472 = pi3327;
  assign po3473 = pi3332;
  assign po3474 = pi3326;
  assign po3475 = pi3356;
  assign po3476 = pi3333;
  assign po3477 = pi3330;
  assign po3478 = pi3325;
  assign po3479 = pi3347;
  assign po3480 = pi3321;
  assign po3481 = pi3345;
  assign po3482 = pi3340;
  assign po3483 = pi3355;
  assign po3484 = pi3334;
  assign po3485 = pi3352;
  assign po3486 = pi3335;
  assign po3487 = pi3354;
  assign po3488 = pi3339;
  assign po3489 = pi3338;
  assign po3490 = pi3348;
  assign po3491 = pi3353;
  assign po3492 = pi3351;
  assign po3493 = pi3341;
  assign po3494 = pi3359;
  assign po3501 = pi3357;
  assign po3503 = pi3360;
  assign po3504 = pi3394;
  assign po3505 = pi3367;
  assign po3506 = pi3365;
  assign po3507 = pi3375;
  assign po3508 = pi3388;
  assign po3509 = pi3376;
  assign po3510 = pi3383;
  assign po3511 = pi3397;
  assign po3512 = pi3342;
  assign po3513 = pi3371;
  assign po3514 = pi3392;
  assign po3515 = pi3373;
  assign po3516 = pi3399;
  assign po3517 = pi3368;
  assign po3518 = pi3363;
  assign po3519 = pi3393;
  assign po3520 = pi3380;
  assign po3521 = pi3398;
  assign po3522 = pi3336;
  assign po3523 = pi3396;
  assign po3524 = pi3364;
  assign po3525 = pi3337;
  assign po3526 = pi3385;
  assign po3527 = pi3374;
  assign po3528 = pi3400;
  assign po3529 = pi3384;
  assign po3530 = pi3377;
  assign po3531 = pi3389;
  assign po3532 = pi3344;
  assign po3533 = pi3372;
  assign po3534 = pi3390;
  assign po3535 = pi3362;
  assign po3536 = pi3381;
  assign po3537 = pi3386;
  assign po3538 = pi3343;
  assign po3542 = pi3391;
  assign po3543 = pi3395;
  assign po3545 = pi3379;
  assign po3546 = pi3382;
  assign po3547 = pi3369;
  assign po3548 = pi3366;
  assign po3549 = pi3378;
  assign po3550 = pi3370;
  assign po3552 = pi3402;
  assign po3553 = pi3358;
  assign po3558 = pi3405;
  assign po3559 = pi3403;
  assign po3561 = pi3404;
  assign po3563 = pi3401;
  assign po3564 = pi3406;
  assign po3565 = pi3407;
  assign po3566 = pi3410;
  assign po3567 = pi3409;
  assign po3568 = pi3416;
  assign po3569 = pi3418;
  assign po3570 = pi3411;
  assign po3571 = pi3408;
  assign po3572 = pi3415;
  assign po3573 = pi3414;
  assign po3574 = pi3419;
  assign po3575 = pi3417;
  assign po3579 = pi3387;
  assign po3580 = pi3422;
  assign po3582 = pi3413;
  assign po3584 = pi3420;
  assign po3585 = pi3412;
  assign po3591 = pi3425;
  assign po3592 = pi3430;
  assign po3593 = pi3439;
  assign po3594 = pi3455;
  assign po3595 = pi3436;
  assign po3596 = pi3438;
  assign po3597 = pi3459;
  assign po3598 = pi3435;
  assign po3599 = pi3460;
  assign po3600 = pi3449;
  assign po3601 = pi3426;
  assign po3602 = pi3442;
  assign po3603 = pi3427;
  assign po3604 = pi3437;
  assign po3605 = pi3432;
  assign po3606 = pi3443;
  assign po3607 = pi3446;
  assign po3608 = pi3444;
  assign po3609 = pi3450;
  assign po3610 = pi3457;
  assign po3611 = pi3445;
  assign po3612 = pi3440;
  assign po3613 = pi3429;
  assign po3614 = pi3462;
  assign po3615 = pi3421;
  assign po3616 = pi3456;
  assign po3618 = pi3424;
  assign po3619 = pi3434;
  assign po3620 = pi3461;
  assign po3621 = pi3453;
  assign po3622 = pi3451;
  assign po3623 = pi3431;
  assign po3624 = pi3441;
  assign po3625 = pi3448;
  assign po3626 = pi3463;
  assign po3627 = pi3428;
  assign po3628 = pi3447;
  assign po3629 = pi3433;
  assign po3630 = pi3452;
  assign po3631 = pi3464;
  assign po3632 = pi3423;
  assign po3636 = pi3477;
  assign po3637 = pi3466;
  assign po3638 = pi3474;
  assign po3639 = pi3478;
  assign po3640 = pi3473;
  assign po3641 = pi3470;
  assign po3642 = pi3467;
  assign po3643 = pi3479;
  assign po3644 = pi3454;
  assign po3645 = pi3475;
  assign po3646 = pi3472;
  assign po3647 = pi3458;
  assign po3648 = pi3465;
  assign po3649 = pi3468;
  assign po3650 = pi3476;
  assign po3651 = pi3480;
  assign po3653 = pi3481;
  assign po3654 = pi3502;
  assign po3655 = pi3519;
  assign po3656 = pi3520;
  assign po3657 = pi3517;
  assign po3658 = pi3498;
  assign po3659 = pi3522;
  assign po3660 = pi3485;
  assign po3661 = pi3523;
  assign po3662 = pi3488;
  assign po3663 = pi3515;
  assign po3664 = pi3489;
  assign po3665 = pi3516;
  assign po3666 = pi3513;
  assign po3667 = pi3503;
  assign po3668 = pi3487;
  assign po3669 = pi3484;
  assign po3670 = pi3504;
  assign po3671 = pi3496;
  assign po3672 = pi3518;
  assign po3673 = pi3483;
  assign po3674 = pi3493;
  assign po3675 = pi3492;
  assign po3676 = pi3505;
  assign po3677 = pi3501;
  assign po3678 = pi3500;
  assign po3679 = pi3495;
  assign po3680 = pi3521;
  assign po3681 = pi3497;
  assign po3682 = pi3508;
  assign po3683 = pi3494;
  assign po3684 = pi3512;
  assign po3685 = pi3511;
  assign po3686 = pi3509;
  assign po3687 = pi3469;
  assign po3688 = pi3471;
  assign po3689 = pi3491;
  assign po3690 = pi3514;
  assign po3691 = pi3507;
  assign po3692 = pi3506;
  assign po3693 = pi3499;
  assign po3694 = pi3482;
  assign po3695 = pi3537;
  assign po3696 = pi3526;
  assign po3697 = pi3530;
  assign po3698 = pi3533;
  assign po3699 = pi3486;
  assign po3700 = pi3538;
  assign po3701 = pi3532;
  assign po3702 = pi3490;
  assign po3703 = pi3525;
  assign po3704 = pi3528;
  assign po3705 = pi3534;
  assign po3706 = pi3527;
  assign po3707 = pi3531;
  assign po3708 = pi3536;
  assign po3709 = pi3529;
  assign po3710 = pi3510;
  assign po3711 = pi3539;
  assign po3713 = pi3553;
  assign po3714 = pi3552;
  assign po3715 = pi3575;
  assign po3716 = pi3543;
  assign po3717 = pi3549;
  assign po3718 = pi3551;
  assign po3719 = pi3579;
  assign po3720 = pi3568;
  assign po3721 = pi3545;
  assign po3722 = pi3560;
  assign po3723 = pi3576;
  assign po3724 = pi3540;
  assign po3725 = pi3565;
  assign po3726 = pi3556;
  assign po3727 = pi3555;
  assign po3728 = pi3564;
  assign po3729 = pi3566;
  assign po3730 = pi3546;
  assign po3731 = pi3544;
  assign po3732 = pi3548;
  assign po3733 = pi3571;
  assign po3734 = pi3541;
  assign po3735 = pi3577;
  assign po3736 = pi3570;
  assign po3737 = pi3550;
  assign po3738 = pi3562;
  assign po3739 = pi3559;
  assign po3740 = pi3535;
  assign po3741 = pi3580;
  assign po3742 = pi3567;
  assign po3743 = pi3542;
  assign po3744 = pi3569;
  assign po3745 = pi3547;
  assign po3746 = pi3573;
  assign po3747 = pi3563;
  assign po3748 = pi3572;
  assign po3749 = pi3554;
  assign po3750 = pi3578;
  assign po3751 = pi3558;
  assign po3752 = pi3574;
  assign po3753 = pi3561;
  assign po3754 = pi3595;
  assign po3755 = pi3590;
  assign po3756 = pi3586;
  assign po3757 = pi3587;
  assign po3758 = pi3583;
  assign po3759 = pi3585;
  assign po3760 = pi3584;
  assign po3761 = pi3593;
  assign po3762 = pi3557;
  assign po3763 = pi3591;
  assign po3764 = pi3582;
  assign po3765 = pi3594;
  assign po3766 = pi3589;
  assign po3767 = pi3592;
  assign po3768 = pi3596;
  assign po3769 = pi3581;
  assign po3770 = pi3621;
  assign po3771 = pi3609;
  assign po3772 = pi3620;
  assign po3773 = pi3627;
  assign po3774 = pi3610;
  assign po3775 = pi3622;
  assign po3776 = pi3631;
  assign po3777 = pi3600;
  assign po3778 = pi3625;
  assign po3779 = pi3604;
  assign po3780 = pi3635;
  assign po3781 = pi3617;
  assign po3782 = pi3636;
  assign po3783 = pi3634;
  assign po3784 = pi3601;
  assign po3785 = pi3599;
  assign po3786 = pi3618;
  assign po3787 = pi3608;
  assign po3788 = pi3614;
  assign po3789 = pi3613;
  assign po3790 = pi3629;
  assign po3791 = pi3624;
  assign po3792 = pi3616;
  assign po3793 = pi3619;
  assign po3794 = pi3597;
  assign po3795 = pi3602;
  assign po3796 = pi3598;
  assign po3797 = pi3588;
  assign po3798 = pi3630;
  assign po3799 = pi3612;
  assign po3800 = pi3637;
  assign po3801 = pi3628;
  assign po3802 = pi3638;
  assign po3803 = pi3603;
  assign po3804 = pi3605;
  assign po3805 = pi3632;
  assign po3806 = pi3626;
  assign po3807 = pi3623;
  assign po3808 = pi3607;
  assign po3809 = pi3633;
  assign po3810 = pi3615;
  assign po3811 = pi3642;
  assign po3812 = pi3641;
  assign po3813 = pi3649;
  assign po3814 = pi3651;
  assign po3815 = pi3648;
  assign po3816 = pi3647;
  assign po3817 = pi3650;
  assign po3818 = pi3653;
  assign po3819 = pi3606;
  assign po3820 = pi3639;
  assign po3821 = pi3611;
  assign po3822 = pi3646;
  assign po3823 = pi3652;
  assign po3824 = pi3640;
  assign po3825 = pi3643;
  assign po3826 = pi3645;
  assign po3827 = pi3693;
  assign po3828 = pi3682;
  assign po3829 = pi3658;
  assign po3830 = pi3672;
  assign po3831 = pi3670;
  assign po3832 = pi3692;
  assign po3833 = pi3664;
  assign po3834 = pi3673;
  assign po3835 = pi3685;
  assign po3836 = pi3677;
  assign po3837 = pi3675;
  assign po3838 = pi3668;
  assign po3839 = pi3696;
  assign po3840 = pi3671;
  assign po3841 = pi3667;
  assign po3842 = pi3694;
  assign po3843 = pi3654;
  assign po3844 = pi3663;
  assign po3845 = pi3698;
  assign po3846 = pi3644;
  assign po3847 = pi3681;
  assign po3848 = pi3669;
  assign po3849 = pi3690;
  assign po3850 = pi3660;
  assign po3851 = pi3661;
  assign po3852 = pi3665;
  assign po3853 = pi3662;
  assign po3854 = pi3695;
  assign po3855 = pi3666;
  assign po3856 = pi3659;
  assign po3857 = pi3678;
  assign po3858 = pi3683;
  assign po3859 = pi3679;
  assign po3860 = pi3691;
  assign po3861 = pi3676;
  assign po3862 = pi3697;
  assign po3863 = pi3699;
  assign po3864 = pi3656;
  assign po3865 = pi3680;
  assign po3866 = pi3674;
  assign po3867 = pi3686;
  assign po3868 = pi3684;
  assign po3869 = pi3687;
  assign po3870 = pi3655;
  assign po3871 = pi3657;
  assign po3873 = pi3706;
  assign po3874 = pi3708;
  assign po3875 = pi3701;
  assign po3876 = pi3702;
  assign po3877 = pi3704;
  assign po3878 = pi3705;
  assign po3879 = pi3700;
  assign po3880 = pi3703;
  assign po3881 = pi3709;
  assign po3882 = pi3707;
  assign po3883 = pi3688;
  assign po3884 = pi3755;
  assign po3885 = pi3722;
  assign po3886 = pi3720;
  assign po3887 = pi3733;
  assign po3888 = pi3758;
  assign po3889 = pi3711;
  assign po3890 = pi3730;
  assign po3891 = pi3732;
  assign po3892 = pi3721;
  assign po3893 = pi3753;
  assign po3894 = pi3750;
  assign po3895 = pi3745;
  assign po3896 = pi3756;
  assign po3897 = pi3716;
  assign po3898 = pi3743;
  assign po3899 = pi3723;
  assign po3900 = pi3747;
  assign po3901 = pi3742;
  assign po3902 = pi3715;
  assign po3903 = pi3734;
  assign po3904 = pi3712;
  assign po3905 = pi3735;
  assign po3906 = pi3725;
  assign po3907 = pi3726;
  assign po3908 = pi3751;
  assign po3909 = pi3740;
  assign po3910 = pi3739;
  assign po3911 = pi3714;
  assign po3912 = pi3749;
  assign po3913 = pi3731;
  assign po3914 = pi3746;
  assign po3915 = pi3717;
  assign po3916 = pi3724;
  assign po3917 = pi3728;
  assign po3918 = pi3737;
  assign po3919 = pi3738;
  assign po3920 = pi3754;
  assign po3921 = pi3741;
  assign po3922 = pi3729;
  assign po3923 = pi3713;
  assign po3924 = pi3757;
  assign po3925 = pi3748;
  assign po3926 = pi3719;
  assign po3927 = pi3718;
  assign po3928 = pi3752;
  assign po3929 = pi3736;
  assign po3930 = pi3772;
  assign po3931 = pi3769;
  assign po3932 = pi3765;
  assign po3933 = pi3777;
  assign po3934 = pi3766;
  assign po3935 = pi3768;
  assign po3936 = pi3727;
  assign po3937 = pi3774;
  assign po3938 = pi3744;
  assign po3939 = pi3773;
  assign po3940 = pi3782;
  assign po3941 = pi3785;
  assign po3942 = pi3838;
  assign po3943 = pi3820;
  assign po3944 = pi3794;
  assign po3945 = pi3830;
  assign po3946 = pi3831;
  assign po3947 = pi3799;
  assign po3948 = pi3826;
  assign po3949 = pi3792;
  assign po3950 = pi3833;
  assign po3951 = pi3811;
  assign po3952 = pi3827;
  assign po3953 = pi3807;
  assign po3954 = pi3818;
  assign po3955 = pi3822;
  assign po3956 = pi3806;
  assign po3957 = pi3796;
  assign po3958 = pi3825;
  assign po3959 = pi3788;
  assign po3960 = pi3813;
  assign po3961 = pi3814;
  assign po3962 = pi3828;
  assign po3963 = pi3804;
  assign po3964 = pi3819;
  assign po3965 = pi3795;
  assign po3966 = pi3823;
  assign po3967 = pi3791;
  assign po3968 = pi3805;
  assign po3969 = pi3836;
  assign po3970 = pi3834;
  assign po3971 = pi3784;
  assign po3972 = pi3787;
  assign po3973 = pi3835;
  assign po3974 = pi3837;
  assign po3975 = pi3829;
  assign po3976 = pi3790;
  assign po3977 = pi3803;
  assign po3978 = pi3817;
  assign po3979 = pi3832;
  assign po3980 = pi3812;
  assign po3981 = pi3786;
  assign po3982 = pi3775;
  assign po3983 = pi3802;
  assign po3984 = pi3801;
  assign po3985 = pi3816;
  assign po3986 = pi3821;
  assign po3987 = pi3808;
  assign po3988 = pi3815;
  assign po3989 = pi3839;
  assign po3990 = pi3866;
  assign po3991 = pi3840;
  assign po3992 = pi3842;
  assign po3993 = pi3845;
  assign po3994 = pi3853;
  assign po3995 = pi3797;
  assign po3996 = pi3798;
  assign po3997 = pi3852;
  assign po3998 = pi3859;
  assign po3999 = pi3858;
  assign po4000 = pi3863;
  assign po4001 = pi3851;
  assign po4002 = pi3855;
  assign po4003 = pi3854;
  assign po4004 = pi3848;
  assign po4005 = pi3850;
  assign po4006 = pi3915;
  assign po4007 = pi3793;
  assign po4008 = pi3865;
  assign po4009 = pi3892;
  assign po4010 = pi3862;
  assign po4011 = pi3861;
  assign po4013 = pi3846;
  assign po4014 = pi3906;
  assign po4015 = pi3923;
  assign po4016 = pi3888;
  assign po4017 = pi3897;
  assign po4018 = pi3886;
  assign po4019 = pi3870;
  assign po4020 = pi3879;
  assign po4021 = pi3913;
  assign po4022 = pi3894;
  assign po4023 = pi3893;
  assign po4024 = pi3890;
  assign po4025 = pi3919;
  assign po4026 = pi3910;
  assign po4027 = pi3904;
  assign po4028 = pi3905;
  assign po4029 = pi3927;
  assign po4030 = pi3940;
  assign po4031 = pi3918;
  assign po4032 = pi3887;
  assign po4033 = pi3873;
  assign po4034 = pi3871;
  assign po4035 = pi3903;
  assign po4036 = pi3911;
  assign po4037 = pi3924;
  assign po4038 = pi3881;
  assign po4039 = pi3912;
  assign po4040 = pi3930;
  assign po4041 = pi3877;
  assign po4042 = pi3916;
  assign po4043 = pi3909;
  assign po4044 = pi3900;
  assign po4045 = pi3868;
  assign po4046 = pi3860;
  assign po4047 = pi3889;
  assign po4048 = pi3901;
  assign po4049 = pi3876;
  assign po4050 = pi3922;
  assign po4051 = pi3908;
  assign po4052 = pi3882;
  assign po4053 = pi3872;
  assign po4054 = pi3895;
  assign po4055 = pi3920;
  assign po4056 = pi3874;
  assign po4057 = pi3896;
  assign po4058 = pi3869;
  assign po4059 = pi3925;
  assign po4060 = pi3880;
  assign po4061 = pi3883;
  assign po4062 = pi3884;
  assign po4063 = pi3878;
  assign po4064 = pi3907;
  assign po4065 = pi3926;
  assign po4066 = pi3899;
  assign po4067 = pi3928;
  assign po4068 = pi3891;
  assign po4071 = pi3931;
  assign po4073 = pi3929;
  assign po4074 = pi3936;
  assign po4077 = pi3935;
  assign po4078 = pi3885;
  assign po4079 = pi3875;
  assign po4080 = pi3902;
  assign po4084 = pi3944;
  assign po4085 = pi3898;
  assign po4086 = pi3943;
  assign po4087 = pi3958;
  assign po4088 = pi3942;
  assign po4089 = pi3914;
  assign po4090 = pi3941;
  assign po4094 = pi3960;
  assign po4097 = pi3939;
  assign po4098 = pi3984;
  assign po4099 = pi3998;
  assign po4101 = pi3982;
  assign po4102 = pi4007;
  assign po4103 = pi4006;
  assign po4104 = pi4004;
  assign po4106 = pi4010;
  assign po4107 = pi4018;
  assign po4108 = pi4027;
  assign po4109 = pi3981;
  assign po4110 = pi3992;
  assign po4111 = pi3983;
  assign po4112 = pi4031;
  assign po4113 = pi3993;
  assign po4114 = pi3994;
  assign po4115 = pi4019;
  assign po4116 = pi4017;
  assign po4117 = pi3991;
  assign po4118 = pi4035;
  assign po4119 = pi4009;
  assign po4120 = pi3974;
  assign po4121 = pi4001;
  assign po4123 = pi4016;
  assign po4124 = pi4026;
  assign po4126 = pi3990;
  assign po4127 = pi3999;
  assign po4128 = pi3979;
  assign po4129 = pi3976;
  assign po4130 = pi3975;
  assign po4131 = pi4013;
  assign po4132 = pi4014;
  assign po4133 = pi4003;
  assign po4134 = pi3988;
  assign po4135 = pi4012;
  assign po4136 = pi3985;
  assign po4137 = pi3987;
  assign po4138 = pi4008;
  assign po4139 = pi4015;
  assign po4140 = pi4034;
  assign po4141 = pi3973;
  assign po4143 = pi4030;
  assign po4144 = pi4005;
  assign po4146 = pi4002;
  assign po4147 = pi3972;
  assign po4148 = pi4033;
  assign po4149 = pi3977;
  assign po4150 = pi3997;
  assign po4151 = pi3989;
  assign po4152 = pi3986;
  assign po4153 = pi4028;
  assign po4154 = pi3980;
  assign po4155 = pi3995;
  assign po4156 = pi3996;
  assign po4157 = pi4032;
  assign po4158 = pi4000;
  assign po4162 = pi4037;
  assign po4163 = pi4044;
  assign po4164 = pi4042;
  assign po4167 = pi4045;
  assign po4168 = pi4036;
  assign po4171 = pi4011;
  assign po4172 = pi3978;
  assign po4174 = pi4020;
  assign po4175 = pi4106;
  assign po4176 = pi4038;
  assign po4177 = pi4097;
  assign po4178 = pi4111;
  assign po4179 = pi4075;
  assign po4180 = pi4114;
  assign po4181 = pi4100;
  assign po4182 = pi4099;
  assign po4183 = pi4120;
  assign po4184 = pi4101;
  assign po4185 = pi4110;
  assign po4186 = pi4105;
  assign po4187 = pi4088;
  assign po4189 = pi4121;
  assign po4191 = pi4122;
  assign po4192 = pi4124;
  assign po4193 = pi4125;
  assign po4194 = pi4137;
  assign po4195 = pi4123;
  assign po4196 = pi4127;
  assign po4197 = pi4135;
  assign po4198 = pi4069;
  assign po4199 = pi4104;
  assign po4200 = pi4098;
  assign po4201 = pi4129;
  assign po4203 = pi4046;
  assign po4204 = pi4094;
  assign po4205 = pi4096;
  assign po4206 = pi4066;
  assign po4207 = pi4081;
  assign po4208 = pi4112;
  assign po4209 = pi4076;
  assign po4210 = pi4062;
  assign po4211 = pi4058;
  assign po4212 = pi4074;
  assign po4213 = pi4061;
  assign po4214 = pi4092;
  assign po4215 = pi4060;
  assign po4216 = pi4103;
  assign po4217 = pi4109;
  assign po4218 = pi4115;
  assign po4220 = pi4091;
  assign po4221 = pi4072;
  assign po4222 = pi4087;
  assign po4223 = pi4116;
  assign po4224 = pi4086;
  assign po4225 = pi4064;
  assign po4226 = pi4051;
  assign po4227 = pi4070;
  assign po4228 = pi4102;
  assign po4229 = pi4057;
  assign po4230 = pi4084;
  assign po4231 = pi4052;
  assign po4232 = pi4049;
  assign po4233 = pi4068;
  assign po4234 = pi4108;
  assign po4235 = pi4113;
  assign po4236 = pi4090;
  assign po4237 = pi4047;
  assign po4238 = pi4083;
  assign po4239 = pi4050;
  assign po4240 = pi4080;
  assign po4241 = pi4085;
  assign po4242 = pi4089;
  assign po4243 = pi4053;
  assign po4244 = pi4065;
  assign po4245 = pi4067;
  assign po4246 = pi4055;
  assign po4247 = pi4056;
  assign po4248 = pi4054;
  assign po4249 = pi4078;
  assign po4250 = pi4071;
  assign po4251 = pi4190;
  assign po4252 = pi4203;
  assign po4253 = pi4136;
  assign po4254 = pi4200;
  assign po4255 = pi4159;
  assign po4256 = pi4048;
  assign po4257 = pi4095;
  assign po4258 = pi4059;
  assign po4259 = pi4169;
  assign po4260 = pi4079;
  assign po4261 = pi4073;
  assign po4262 = pi4082;
  assign po4263 = pi4077;
  assign po4264 = pi4093;
  assign po4265 = pi4063;
  assign po4266 = pi4213;
  assign po4267 = pi4215;
  assign po4268 = pi4208;
  assign po4269 = pi4209;
  assign po4270 = pi4128;
  assign po4271 = pi4207;
  assign po4272 = pi4205;
  assign po4273 = pi4212;
  assign po4274 = pi4214;
  assign po4275 = pi4206;
  assign po4276 = pi4161;
  assign po4277 = pi4154;
  assign po4278 = pi4153;
  assign po4279 = pi4142;
  assign po4280 = pi4150;
  assign po4281 = pi4189;
  assign po4282 = pi4177;
  assign po4283 = pi4155;
  assign po4284 = pi4187;
  assign po4285 = pi4201;
  assign po4286 = pi4165;
  assign po4287 = pi4174;
  assign po4288 = pi4197;
  assign po4289 = pi4149;
  assign po4290 = pi4144;
  assign po4291 = pi4172;
  assign po4292 = pi4158;
  assign po4293 = pi4182;
  assign po4294 = pi4170;
  assign po4295 = pi4185;
  assign po4296 = pi4199;
  assign po4297 = pi4146;
  assign po4298 = pi4178;
  assign po4299 = pi4220;
  assign po4300 = pi4171;
  assign po4301 = pi4176;
  assign po4302 = pi4145;
  assign po4303 = pi4167;
  assign po4304 = pi4148;
  assign po4305 = pi4285;
  assign po4306 = pi4198;
  assign po4307 = pi4162;
  assign po4308 = pi4160;
  assign po4309 = pi4147;
  assign po4310 = pi4164;
  assign po4311 = pi4166;
  assign po4312 = pi4183;
  assign po4313 = pi4194;
  assign po4314 = pi4181;
  assign po4315 = pi4152;
  assign po4316 = pi4151;
  assign po4317 = pi4175;
  assign po4318 = pi4293;
  assign po4319 = pi4140;
  assign po4320 = pi4163;
  assign po4321 = pi4139;
  assign po4322 = pi4157;
  assign po4323 = pi4195;
  assign po4324 = pi4180;
  assign po4325 = pi4141;
  assign po4326 = pi4188;
  assign po4327 = pi4246;
  assign po4328 = pi4280;
  assign po4329 = pi4292;
  assign po4330 = pi4247;
  assign po4331 = pi4211;
  assign po4332 = pi4156;
  assign po4333 = pi4196;
  assign po4334 = pi4204;
  assign po4335 = pi4249;
  assign po4336 = pi4287;
  assign po4337 = pi4184;
  assign po4338 = pi4168;
  assign po4339 = pi4143;
  assign po4340 = pi4284;
  assign po4341 = pi4288;
  assign po4342 = pi4202;
  assign po4343 = pi4173;
  assign po4344 = pi4254;
  assign po4345 = pi4179;
  assign po4346 = pi4186;
  assign po4347 = pi4279;
  assign po4348 = pi4191;
  assign po4349 = pi4252;
  assign po4350 = pi4286;
  assign po4351 = pi4228;
  assign po4352 = pi4297;
  assign po4353 = pi4221;
  assign po4354 = pi4303;
  assign po4355 = pi4294;
  assign po4356 = pi4301;
  assign po4357 = pi4296;
  assign po4358 = pi4309;
  assign po4359 = pi4308;
  assign po4360 = pi4298;
  assign po4361 = pi4299;
  assign po4362 = pi4216;
  assign po4363 = pi4300;
  assign po4364 = pi4295;
  assign po4365 = pi4281;
  assign po4366 = pi4282;
  assign po4367 = pi4302;
  assign po4368 = pi4307;
  assign po4369 = pi4226;
  assign po4370 = pi4283;
  assign po4371 = pi4225;
  assign po4372 = pi4251;
  assign po4373 = pi4245;
  assign po4374 = pi4256;
  assign po4375 = pi4255;
  assign po4376 = pi4275;
  assign po4377 = pi4239;
  assign po4378 = pi4250;
  assign po4379 = pi4274;
  assign po4380 = pi4248;
  assign po4381 = pi4233;
  assign po4382 = pi4217;
  assign po4383 = pi4231;
  assign po4384 = pi4235;
  assign po4385 = pi4278;
  assign po4386 = pi4242;
  assign po4387 = pi4229;
  assign po4388 = pi4272;
  assign po4389 = pi4306;
  assign po4390 = pi4223;
  assign po4391 = pi4289;
  assign po4392 = pi4270;
  assign po4393 = pi4222;
  assign po4394 = pi4258;
  assign po4395 = pi4224;
  assign po4396 = pi4264;
  assign po4397 = pi4236;
  assign po4398 = pi4291;
  assign po4399 = pi4379;
  assign po4400 = pi4268;
  assign po4401 = pi4257;
  assign po4402 = pi4237;
  assign po4403 = pi4262;
  assign po4404 = pi4241;
  assign po4405 = pi4261;
  assign po4406 = pi4232;
  assign po4407 = pi4263;
  assign po4408 = pi4227;
  assign po4409 = pi4243;
  assign po4410 = pi4259;
  assign po4411 = pi4219;
  assign po4412 = pi4238;
  assign po4413 = pi4273;
  assign po4414 = pi4316;
  assign po4415 = pi4230;
  assign po4416 = pi4253;
  assign po4417 = pi4244;
  assign po4418 = pi4276;
  assign po4419 = pi4218;
  assign po4420 = pi4373;
  assign po4421 = pi4311;
  assign po4422 = pi4317;
  assign po4423 = pi4375;
  assign po4424 = pi4265;
  assign po4425 = pi4240;
  assign po4426 = pi4234;
  assign po4427 = pi4290;
  assign po4428 = pi4260;
  assign po4429 = pi4267;
  assign po4430 = pi4310;
  assign po4431 = pi4269;
  assign po4432 = pi4271;
  assign po4433 = pi4374;
  assign po4434 = pi4381;
  assign po4435 = pi4397;
  assign po4436 = pi4385;
  assign po4437 = pi4304;
  assign po4438 = pi4400;
  assign po4439 = pi4380;
  assign po4440 = pi4305;
  assign po4441 = pi4399;
  assign po4442 = pi4382;
  assign po4443 = pi4393;
  assign po4444 = pi4394;
  assign po4445 = pi4392;
  assign po4446 = pi4384;
  assign po4447 = pi4338;
  assign po4448 = pi4357;
  assign po4449 = pi4333;
  assign po4450 = pi4408;
  assign po4451 = pi4490;
  assign po4452 = pi4361;
  assign po4453 = pi4362;
  assign po4454 = pi4354;
  assign po4455 = pi4345;
  assign po4456 = pi4325;
  assign po4457 = pi4319;
  assign po4458 = pi4403;
  assign po4459 = pi4363;
  assign po4460 = pi4364;
  assign po4461 = pi4334;
  assign po4462 = pi4368;
  assign po4463 = pi4340;
  assign po4464 = pi4360;
  assign po4465 = pi4322;
  assign po4466 = pi4342;
  assign po4467 = pi4366;
  assign po4468 = pi4318;
  assign po4469 = pi4371;
  assign po4470 = pi4353;
  assign po4471 = pi4356;
  assign po4472 = pi4359;
  assign po4473 = pi4344;
  assign po4474 = pi4336;
  assign po4475 = pi4335;
  assign po4476 = pi4481;
  assign po4477 = pi4401;
  assign po4478 = pi4332;
  assign po4479 = pi4396;
  assign po4480 = pi4369;
  assign po4481 = pi4372;
  assign po4482 = pi4404;
  assign po4483 = pi4330;
  assign po4484 = pi4473;
  assign po4485 = pi4331;
  assign po4486 = pi4326;
  assign po4487 = pi4337;
  assign po4488 = pi4350;
  assign po4489 = pi4365;
  assign po4490 = pi4347;
  assign po4491 = pi4358;
  assign po4492 = pi4349;
  assign po4493 = pi4370;
  assign po4494 = pi4376;
  assign po4495 = pi4355;
  assign po4496 = pi4383;
  assign po4497 = pi4377;
  assign po4498 = pi4343;
  assign po4499 = pi4315;
  assign po4500 = pi4346;
  assign po4501 = pi4339;
  assign po4502 = pi4351;
  assign po4503 = pi4367;
  assign po4504 = pi4314;
  assign po4505 = pi4327;
  assign po4506 = pi4378;
  assign po4507 = pi4446;
  assign po4508 = pi4329;
  assign po4509 = pi4484;
  assign po4510 = pi4475;
  assign po4511 = pi4413;
  assign po4512 = pi4409;
  assign po4513 = pi4341;
  assign po4514 = pi4483;
  assign po4515 = pi4402;
  assign po4516 = pi4480;
  assign po4517 = pi4425;
  assign po4518 = pi4477;
  assign po4519 = pi4328;
  assign po4520 = pi4348;
  assign po4521 = pi4352;
  assign po4522 = pi4419;
  assign po4523 = pi4482;
  assign po4524 = pi4506;
  assign po4525 = pi4398;
  assign po4526 = pi4479;
  assign po4527 = pi4485;
  assign po4528 = pi4391;
  assign po4529 = pi4497;
  assign po4530 = pi4493;
  assign po4531 = pi4505;
  assign po4532 = pi4494;
  assign po4533 = pi4511;
  assign po4534 = pi4507;
  assign po4535 = pi4491;
  assign po4536 = pi4510;
  assign po4537 = pi4495;
  assign po4538 = pi4492;
  assign po4539 = pi4509;
  assign po4540 = pi4579;
  assign po4541 = pi4521;
  assign po4542 = pi4543;
  assign po4543 = pi4542;
  assign po4544 = pi4436;
  assign po4545 = pi4428;
  assign po4546 = pi4561;
  assign po4547 = pi4489;
  assign po4548 = pi4467;
  assign po4549 = pi4435;
  assign po4550 = pi4538;
  assign po4551 = pi4544;
  assign po4552 = pi4463;
  assign po4553 = pi4541;
  assign po4554 = pi4540;
  assign po4555 = pi4486;
  assign po4556 = pi4447;
  assign po4557 = pi4456;
  assign po4558 = pi4426;
  assign po4559 = pi4437;
  assign po4560 = pi4429;
  assign po4561 = pi4416;
  assign po4562 = pi4454;
  assign po4563 = pi4452;
  assign po4564 = pi4462;
  assign po4565 = pi4455;
  assign po4566 = pi4406;
  assign po4567 = pi4469;
  assign po4568 = pi4427;
  assign po4569 = pi4422;
  assign po4570 = pi4405;
  assign po4571 = pi4464;
  assign po4572 = pi4415;
  assign po4573 = pi4410;
  assign po4574 = pi4432;
  assign po4575 = pi4430;
  assign po4576 = pi4414;
  assign po4577 = pi4411;
  assign po4578 = pi4421;
  assign po4579 = pi4448;
  assign po4580 = pi4470;
  assign po4581 = pi4471;
  assign po4582 = pi4451;
  assign po4583 = pi4444;
  assign po4584 = pi4466;
  assign po4585 = pi4438;
  assign po4586 = pi4442;
  assign po4587 = pi4412;
  assign po4588 = pi4468;
  assign po4589 = pi4417;
  assign po4590 = pi4433;
  assign po4591 = pi4418;
  assign po4592 = pi4431;
  assign po4593 = pi4449;
  assign po4594 = pi4461;
  assign po4595 = pi4420;
  assign po4596 = pi4450;
  assign po4597 = pi4453;
  assign po4598 = pi4459;
  assign po4599 = pi4465;
  assign po4600 = pi4424;
  assign po4601 = pi4472;
  assign po4602 = pi4457;
  assign po4603 = pi4508;
  assign po4604 = pi4578;
  assign po4605 = pi4588;
  assign po4606 = pi4460;
  assign po4607 = pi4441;
  assign po4608 = pi4458;
  assign po4609 = pi4583;
  assign po4610 = pi4603;
  assign po4611 = pi4590;
  assign po4612 = pi4615;
  assign po4613 = pi4593;
  assign po4614 = pi4553;
  assign po4615 = pi4607;
  assign po4616 = pi4599;
  assign po4617 = pi4614;
  assign po4618 = pi4598;
  assign po4619 = pi4592;
  assign po4620 = pi4514;
  assign po4621 = pi4512;
  assign po4622 = pi4613;
  assign po4623 = pi4619;
  assign po4624 = pi4605;
  assign po4625 = pi4600;
  assign po4626 = pi4617;
  assign po4627 = pi4611;
  assign po4628 = pi4602;
  assign po4629 = pi4620;
  assign po4630 = pi4616;
  assign po4631 = pi4692;
  assign po4632 = pi4604;
  assign po4633 = pi4690;
  assign po4634 = pi4650;
  assign po4635 = pi4527;
  assign po4636 = pi4513;
  assign po4637 = pi4663;
  assign po4638 = pi4695;
  assign po4639 = pi4691;
  assign po4640 = pi4587;
  assign po4641 = pi4576;
  assign po4642 = pi4556;
  assign po4643 = pi4612;
  assign po4644 = pi4554;
  assign po4645 = pi4515;
  assign po4646 = pi4552;
  assign po4647 = pi4571;
  assign po4648 = pi4566;
  assign po4649 = pi4699;
  assign po4650 = pi4549;
  assign po4651 = pi4545;
  assign po4652 = pi4562;
  assign po4653 = pi4664;
  assign po4654 = pi4589;
  assign po4655 = pi4685;
  assign po4656 = pi4520;
  assign po4657 = pi4557;
  assign po4658 = pi4572;
  assign po4659 = pi4581;
  assign po4660 = pi4559;
  assign po4661 = pi4516;
  assign po4662 = pi4575;
  assign po4663 = pi4582;
  assign po4664 = pi4595;
  assign po4665 = pi4569;
  assign po4666 = pi4570;
  assign po4667 = pi4535;
  assign po4668 = pi4539;
  assign po4669 = pi4658;
  assign po4670 = pi4594;
  assign po4671 = pi4550;
  assign po4672 = pi4574;
  assign po4673 = pi4672;
  assign po4674 = pi4564;
  assign po4675 = pi4669;
  assign po4676 = pi4698;
  assign po4677 = pi4524;
  assign po4678 = pi4577;
  assign po4679 = pi4565;
  assign po4680 = pi4563;
  assign po4681 = pi4551;
  assign po4682 = pi4568;
  assign po4683 = pi4525;
  assign po4684 = pi4526;
  assign po4685 = pi4518;
  assign po4686 = pi4580;
  assign po4687 = pi4519;
  assign po4688 = pi4547;
  assign po4689 = pi4529;
  assign po4690 = pi4558;
  assign po4691 = pi4586;
  assign po4692 = pi4528;
  assign po4693 = pi4531;
  assign po4694 = pi4523;
  assign po4695 = pi4567;
  assign po4696 = pi4548;
  assign po4697 = pi4555;
  assign po4698 = pi4533;
  assign po4699 = pi4517;
  assign po4700 = pi4530;
  assign po4701 = pi4522;
  assign po4702 = pi4573;
  assign po4703 = pi4654;
  assign po4704 = pi4668;
  assign po4705 = pi4689;
  assign po4706 = pi4661;
  assign po4707 = pi4606;
  assign po4708 = pi4667;
  assign po4709 = pi4608;
  assign po4710 = pi4652;
  assign po4711 = pi4623;
  assign po4712 = pi4710;
  assign po4713 = pi4709;
  assign po4714 = pi4678;
  assign po4715 = pi4618;
  assign po4716 = pi4560;
  assign po4717 = pi4659;
  assign po4718 = pi4660;
  assign po4719 = pi4711;
  assign po4720 = pi4675;
  assign po4721 = pi4591;
  assign po4722 = pi4610;
  assign po4723 = pi4718;
  assign po4724 = pi4716;
  assign po4725 = pi4730;
  assign po4726 = pi4724;
  assign po4727 = pi4735;
  assign po4728 = pi4674;
  assign po4729 = pi4728;
  assign po4730 = pi4726;
  assign po4731 = pi4719;
  assign po4732 = pi4732;
  assign po4733 = pi4722;
  assign po4734 = pi4721;
  assign po4735 = pi4609;
  assign po4736 = pi4715;
  assign po4737 = pi4733;
  assign po4738 = pi4707;
  assign po4739 = pi4734;
  assign po4740 = pi4738;
  assign po4741 = pi4737;
  assign po4742 = pi4736;
  assign po4743 = pi4697;
  assign po4744 = pi4800;
  assign po4745 = pi4641;
  assign po4746 = pi4625;
  assign po4747 = pi4643;
  assign po4748 = pi4631;
  assign po4749 = pi4680;
  assign po4750 = pi4628;
  assign po4751 = pi4754;
  assign po4752 = pi4696;
  assign po4753 = pi4624;
  assign po4754 = pi4673;
  assign po4755 = pi4653;
  assign po4756 = pi4632;
  assign po4757 = pi4621;
  assign po4758 = pi4687;
  assign po4759 = pi4636;
  assign po4760 = pi4679;
  assign po4761 = pi4714;
  assign po4762 = pi4727;
  assign po4763 = pi4644;
  assign po4764 = pi4666;
  assign po4765 = pi4648;
  assign po4766 = pi4756;
  assign po4767 = pi4665;
  assign po4768 = pi4752;
  assign po4769 = pi4712;
  assign po4770 = pi4761;
  assign po4771 = pi4759;
  assign po4772 = pi4758;
  assign po4773 = pi4751;
  assign po4774 = pi4750;
  assign po4775 = pi4703;
  assign po4776 = pi4763;
  assign po4777 = pi4683;
  assign po4778 = pi4708;
  assign po4779 = pi4713;
  assign po4780 = pi4701;
  assign po4781 = pi4639;
  assign po4782 = pi4627;
  assign po4783 = pi4780;
  assign po4784 = pi4681;
  assign po4785 = pi4629;
  assign po4786 = pi4635;
  assign po4787 = pi4676;
  assign po4788 = pi4694;
  assign po4789 = pi4630;
  assign po4790 = pi4677;
  assign po4791 = pi4781;
  assign po4792 = pi4651;
  assign po4793 = pi4622;
  assign po4794 = pi4702;
  assign po4795 = pi4626;
  assign po4796 = pi4704;
  assign po4797 = pi4655;
  assign po4798 = pi4637;
  assign po4799 = pi4640;
  assign po4800 = pi4688;
  assign po4801 = pi4700;
  assign po4802 = pi4693;
  assign po4803 = pi4671;
  assign po4804 = pi4633;
  assign po4805 = pi4638;
  assign po4806 = pi4634;
  assign po4807 = pi4649;
  assign po4808 = pi4774;
  assign po4809 = pi4794;
  assign po4810 = pi4642;
  assign po4811 = pi4684;
  assign po4812 = pi4682;
  assign po4813 = pi4772;
  assign po4814 = pi4725;
  assign po4815 = pi4670;
  assign po4816 = pi4686;
  assign po4817 = pi4647;
  assign po4818 = pi4805;
  assign po4819 = pi4705;
  assign po4820 = pi4821;
  assign po4821 = pi4839;
  assign po4822 = pi4824;
  assign po4823 = pi4731;
  assign po4824 = pi4826;
  assign po4825 = pi4825;
  assign po4826 = pi4830;
  assign po4827 = pi4723;
  assign po4828 = pi4828;
  assign po4829 = pi4819;
  assign po4830 = pi4820;
  assign po4831 = pi4823;
  assign po4832 = pi4815;
  assign po4833 = pi4816;
  assign po4834 = pi4841;
  assign po4835 = pi4844;
  assign po4836 = pi4818;
  assign po4837 = pi4846;
  assign po4838 = pi4843;
  assign po4839 = pi4817;
  assign po4840 = pi4840;
  assign po4841 = pi4833;
  assign po4842 = pi4842;
  assign po4843 = pi4834;
  assign po4844 = pi4829;
  assign po4845 = pi4831;
  assign po4846 = pi4845;
  assign po4847 = pi4849;
  assign po4848 = pi4838;
  assign po4849 = pi4847;
  assign po4850 = pi4835;
  assign po4851 = pi4770;
  assign po4852 = pi4790;
  assign po4853 = pi4923;
  assign po4854 = pi4786;
  assign po4855 = pi4788;
  assign po4856 = pi4766;
  assign po4857 = pi4783;
  assign po4858 = pi4744;
  assign po4859 = pi4777;
  assign po4860 = pi4806;
  assign po4861 = pi4741;
  assign po4862 = pi4768;
  assign po4863 = pi4739;
  assign po4864 = pi4814;
  assign po4865 = pi4762;
  assign po4866 = pi4808;
  assign po4867 = pi4775;
  assign po4868 = pi4779;
  assign po4869 = pi4795;
  assign po4870 = pi4798;
  assign po4871 = pi4753;
  assign po4872 = pi4789;
  assign po4873 = pi4765;
  assign po4874 = pi4740;
  assign po4875 = pi4873;
  assign po4876 = pi4860;
  assign po4877 = pi4776;
  assign po4878 = pi4799;
  assign po4879 = pi4797;
  assign po4880 = pi4891;
  assign po4881 = pi4792;
  assign po4882 = pi4854;
  assign po4883 = pi4745;
  assign po4884 = pi4836;
  assign po4885 = pi4785;
  assign po4886 = pi4867;
  assign po4887 = pi4858;
  assign po4888 = pi4938;
  assign po4889 = pi4827;
  assign po4890 = pi4941;
  assign po4891 = pi4862;
  assign po4892 = pi4864;
  assign po4893 = pi4863;
  assign po4894 = pi4868;
  assign po4895 = pi4859;
  assign po4896 = pi4866;
  assign po4897 = pi4856;
  assign po4898 = pi4939;
  assign po4899 = pi4942;
  assign po4900 = pi4855;
  assign po4901 = pi4746;
  assign po4902 = pi4848;
  assign po4903 = pi4769;
  assign po4904 = pi4869;
  assign po4905 = pi4890;
  assign po4906 = pi4791;
  assign po4907 = pi4793;
  assign po4908 = pi4883;
  assign po4909 = pi4767;
  assign po4910 = pi4809;
  assign po4911 = pi4812;
  assign po4912 = pi4755;
  assign po4913 = pi4811;
  assign po4914 = pi4784;
  assign po4915 = pi4943;
  assign po4916 = pi4771;
  assign po4917 = pi4747;
  assign po4918 = pi4810;
  assign po4919 = pi4881;
  assign po4920 = pi4837;
  assign po4921 = pi4874;
  assign po4922 = pi4906;
  assign po4923 = pi4796;
  assign po4924 = pi4743;
  assign po4925 = pi4911;
  assign po4926 = pi4787;
  assign po4927 = pi4801;
  assign po4928 = pi4852;
  assign po4929 = pi4882;
  assign po4930 = pi4749;
  assign po4931 = pi4742;
  assign po4932 = pi4802;
  assign po4933 = pi4778;
  assign po4934 = pi4748;
  assign po4935 = pi4807;
  assign po4936 = pi4872;
  assign po4937 = pi4898;
  assign po4938 = pi4773;
  assign po4939 = pi4876;
  assign po4940 = pi4832;
  assign po4941 = pi4850;
  assign po4942 = pi4760;
  assign po4943 = pi4813;
  assign po4944 = pi4782;
  assign po4945 = pi4964;
  assign po4946 = pi4961;
  assign po4947 = pi4950;
  assign po4948 = pi4947;
  assign po4949 = pi4870;
  assign po4950 = pi4955;
  assign po4951 = pi4865;
  assign po4952 = pi4956;
  assign po4953 = pi4952;
  assign po4954 = pi4953;
  assign po4955 = pi4954;
  assign po4956 = pi4951;
  assign po4957 = pi4857;
  assign po4958 = pi4968;
  assign po4959 = pi4871;
  assign po4960 = pi4959;
  assign po4961 = pi4958;
  assign po4962 = pi4948;
  assign po4963 = pi4957;
  assign po4964 = pi4962;
  assign po4965 = pi4949;
  assign po4966 = pi4967;
  assign po4967 = pi4963;
  assign po4968 = pi4909;
  assign po4969 = pi4936;
  assign po4970 = pi4932;
  assign po4971 = pi4908;
  assign po4972 = pi4880;
  assign po4973 = pi4895;
  assign po4974 = pi4946;
  assign po4975 = pi4878;
  assign po4976 = pi4901;
  assign po4977 = pi4907;
  assign po4978 = pi4879;
  assign po4979 = pi4851;
  assign po4980 = pi4971;
  assign po4981 = pi5036;
  assign po4982 = pi4989;
  assign po4983 = pi4886;
  assign po4984 = pi5038;
  assign po4985 = pi4917;
  assign po4986 = pi4977;
  assign po4987 = pi4975;
  assign po4988 = pi4976;
  assign po4989 = pi4974;
  assign po4990 = pi4912;
  assign po4991 = pi5042;
  assign po4992 = pi4929;
  assign po4993 = pi4893;
  assign po4994 = pi4980;
  assign po4995 = pi4920;
  assign po4996 = pi4944;
  assign po4997 = pi4913;
  assign po4998 = pi4927;
  assign po4999 = pi4925;
  assign po5000 = pi4914;
  assign po5001 = pi4853;
  assign po5002 = pi4984;
  assign po5003 = pi4889;
  assign po5004 = pi4987;
  assign po5005 = pi4894;
  assign po5006 = pi4928;
  assign po5007 = pi4904;
  assign po5008 = pi4924;
  assign po5009 = pi4919;
  assign po5010 = pi4990;
  assign po5011 = pi4988;
  assign po5012 = pi4902;
  assign po5013 = pi4877;
  assign po5014 = pi4888;
  assign po5015 = pi4900;
  assign po5016 = pi4935;
  assign po5017 = pi4892;
  assign po5018 = pi4930;
  assign po5019 = pi4915;
  assign po5020 = pi4934;
  assign po5021 = pi4875;
  assign po5022 = pi4933;
  assign po5023 = pi4905;
  assign po5024 = pi5039;
  assign po5025 = pi4903;
  assign po5026 = pi4931;
  assign po5027 = pi4921;
  assign po5028 = pi4896;
  assign po5029 = pi4884;
  assign po5030 = pi4979;
  assign po5031 = pi4916;
  assign po5032 = pi4945;
  assign po5033 = pi4969;
  assign po5034 = pi4861;
  assign po5035 = pi4937;
  assign po5036 = pi4922;
  assign po5037 = pi4918;
  assign po5038 = pi4910;
  assign po5039 = pi4885;
  assign po5040 = pi4897;
  assign po5041 = pi4887;
  assign po5042 = pi4940;
  assign po5043 = pi4899;
  assign po5044 = pi4926;
  assign po5045 = pi5060;
  assign po5046 = pi4960;
  assign po5047 = pi4966;
  assign po5048 = pi5058;
  assign po5049 = pi5080;
  assign po5050 = pi5057;
  assign po5051 = pi5065;
  assign po5052 = pi5054;
  assign po5053 = pi5052;
  assign po5054 = pi5051;
  assign po5055 = pi5055;
  assign po5056 = pi5049;
  assign po5057 = pi5047;
  assign po5058 = pi5046;
  assign po5059 = pi5082;
  assign po5060 = pi5081;
  assign po5061 = pi4965;
  assign po5062 = pi5079;
  assign po5063 = pi5068;
  assign po5064 = pi5062;
  assign po5065 = pi5066;
  assign po5066 = pi5072;
  assign po5067 = pi5078;
  assign po5068 = pi5061;
  assign po5069 = pi5063;
  assign po5070 = pi5064;
  assign po5071 = pi5075;
  assign po5072 = pi5076;
  assign po5073 = pi5067;
  assign po5074 = pi5074;
  assign po5075 = pi5083;
  assign po5076 = pi5069;
  assign po5077 = pi5070;
  assign po5078 = pi5056;
  assign po5079 = pi5071;
  assign po5080 = pi5059;
  assign po5081 = pi5014;
  assign po5082 = pi5037;
  assign po5083 = pi5040;
  assign po5084 = pi5154;
  assign po5085 = pi5053;
  assign po5086 = pi5094;
  assign po5087 = pi5093;
  assign po5088 = pi5090;
  assign po5089 = pi5106;
  assign po5090 = pi5111;
  assign po5091 = pi5114;
  assign po5092 = pi5096;
  assign po5093 = pi5099;
  assign po5094 = pi4970;
  assign po5095 = pi5108;
  assign po5096 = pi5109;
  assign po5097 = pi5095;
  assign po5098 = pi5101;
  assign po5099 = pi5091;
  assign po5100 = pi5105;
  assign po5101 = pi5092;
  assign po5102 = pi5087;
  assign po5103 = pi4978;
  assign po5104 = pi5156;
  assign po5105 = pi5032;
  assign po5106 = pi5164;
  assign po5107 = pi5017;
  assign po5108 = pi4997;
  assign po5109 = pi5001;
  assign po5110 = pi5030;
  assign po5111 = pi5112;
  assign po5112 = pi5144;
  assign po5113 = pi5043;
  assign po5114 = pi4983;
  assign po5115 = pi5031;
  assign po5116 = pi5029;
  assign po5117 = pi4985;
  assign po5118 = pi4972;
  assign po5119 = pi5022;
  assign po5120 = pi5151;
  assign po5121 = pi5116;
  assign po5122 = pi5007;
  assign po5123 = pi5104;
  assign po5124 = pi4986;
  assign po5125 = pi5006;
  assign po5126 = pi5021;
  assign po5127 = pi5008;
  assign po5128 = pi5152;
  assign po5129 = pi5016;
  assign po5130 = pi5020;
  assign po5131 = pi5010;
  assign po5132 = pi4999;
  assign po5133 = pi5005;
  assign po5134 = pi4982;
  assign po5135 = pi5041;
  assign po5136 = pi5155;
  assign po5137 = pi5024;
  assign po5138 = pi5015;
  assign po5139 = pi5117;
  assign po5140 = pi5023;
  assign po5141 = pi5143;
  assign po5142 = pi4992;
  assign po5143 = pi5044;
  assign po5144 = pi4993;
  assign po5145 = pi4991;
  assign po5146 = pi4995;
  assign po5147 = pi4981;
  assign po5148 = pi5002;
  assign po5149 = pi5012;
  assign po5150 = pi5019;
  assign po5151 = pi5004;
  assign po5152 = pi4994;
  assign po5153 = pi5073;
  assign po5154 = pi5013;
  assign po5155 = pi5018;
  assign po5156 = pi5027;
  assign po5157 = pi5025;
  assign po5158 = pi4998;
  assign po5159 = pi5009;
  assign po5160 = pi5035;
  assign po5161 = pi5033;
  assign po5162 = pi5045;
  assign po5163 = pi5028;
  assign po5164 = pi4996;
  assign po5165 = pi4973;
  assign po5166 = pi5000;
  assign po5167 = pi5150;
  assign po5168 = pi5048;
  assign po5169 = pi5097;
  assign po5170 = pi5026;
  assign po5171 = pi5107;
  assign po5172 = pi5103;
  assign po5173 = pi5089;
  assign po5174 = pi5034;
  assign po5175 = pi5011;
  assign po5176 = pi5003;
  assign po5177 = pi5077;
  assign po5178 = pi5088;
  assign po5179 = pi5185;
  assign po5180 = pi5050;
  assign po5181 = pi5180;
  assign po5182 = pi5181;
  assign po5183 = pi5179;
  assign po5184 = pi5178;
  assign po5185 = pi5186;
  assign po5186 = pi5110;
  assign po5187 = pi5194;
  assign po5188 = pi5187;
  assign po5189 = pi5184;
  assign po5190 = pi5189;
  assign po5191 = pi5190;
  assign po5192 = pi5196;
  assign po5193 = pi5193;
  assign po5194 = pi5188;
  assign po5195 = pi5182;
  assign po5196 = pi5195;
  assign po5197 = pi5192;
  assign po5198 = pi5102;
  assign po5199 = pi5211;
  assign po5200 = pi5100;
  assign po5201 = pi5214;
  assign po5202 = pi5129;
  assign po5203 = pi5175;
  assign po5204 = pi5213;
  assign po5205 = pi5210;
  assign po5206 = pi5215;
  assign po5207 = pi5208;
  assign po5208 = pi5206;
  assign po5209 = pi5207;
  assign po5210 = pi5277;
  assign po5211 = pi5177;
  assign po5212 = pi5120;
  assign po5213 = pi5086;
  assign po5214 = pi5252;
  assign po5215 = pi5165;
  assign po5216 = pi5137;
  assign po5217 = pi5253;
  assign po5218 = pi5250;
  assign po5219 = pi5204;
  assign po5220 = pi5262;
  assign po5221 = pi5141;
  assign po5222 = pi5134;
  assign po5223 = pi5124;
  assign po5224 = pi5149;
  assign po5225 = pi5169;
  assign po5226 = pi5145;
  assign po5227 = pi5133;
  assign po5228 = pi5121;
  assign po5229 = pi5123;
  assign po5230 = pi5142;
  assign po5231 = pi5172;
  assign po5232 = pi5127;
  assign po5233 = pi5132;
  assign po5234 = pi5085;
  assign po5235 = pi5167;
  assign po5236 = pi5148;
  assign po5237 = pi5139;
  assign po5238 = pi5131;
  assign po5239 = pi5115;
  assign po5240 = pi5140;
  assign po5241 = pi5126;
  assign po5242 = pi5157;
  assign po5243 = pi5138;
  assign po5244 = pi5163;
  assign po5245 = pi5170;
  assign po5246 = pi5168;
  assign po5247 = pi5176;
  assign po5248 = pi5166;
  assign po5249 = pi5158;
  assign po5250 = pi5162;
  assign po5251 = pi5147;
  assign po5252 = pi5118;
  assign po5253 = pi5119;
  assign po5254 = pi5128;
  assign po5255 = pi5084;
  assign po5256 = pi5125;
  assign po5257 = pi5153;
  assign po5258 = pi5171;
  assign po5259 = pi5159;
  assign po5260 = pi5130;
  assign po5261 = pi5160;
  assign po5262 = pi5146;
  assign po5263 = pi5136;
  assign po5264 = pi5122;
  assign po5265 = pi5173;
  assign po5266 = pi5203;
  assign po5267 = pi5278;
  assign po5268 = pi5245;
  assign po5269 = pi5267;
  assign po5270 = pi5174;
  assign po5271 = pi5135;
  assign po5272 = pi5212;
  assign po5273 = pi5255;
  assign po5274 = pi5161;
  assign po5275 = pi5113;
  assign po5276 = pi5288;
  assign po5277 = pi5287;
  assign po5278 = pi5289;
  assign po5279 = pi5297;
  assign po5280 = pi5291;
  assign po5281 = pi5296;
  assign po5282 = pi5290;
  assign po5283 = pi5283;
  assign po5284 = pi5295;
  assign po5285 = pi5286;
  assign po5286 = pi5284;
  assign po5287 = pi5285;
  assign po5288 = pi5318;
  assign po5289 = pi5314;
  assign po5290 = pi5302;
  assign po5291 = pi5303;
  assign po5292 = pi5306;
  assign po5293 = pi5315;
  assign po5294 = pi5313;
  assign po5295 = pi5316;
  assign po5296 = pi5321;
  assign po5297 = pi5309;
  assign po5298 = pi5319;
  assign po5299 = pi5325;
  assign po5300 = pi5324;
  assign po5301 = pi5305;
  assign po5302 = pi5308;
  assign po5303 = pi5299;
  assign po5304 = pi5322;
  assign po5305 = pi5323;
  assign po5306 = pi5317;
  assign po5307 = pi5312;
  assign po5308 = pi5293;
  assign po5309 = pi5311;
  assign po5310 = pi5298;
  assign po5311 = pi5281;
  assign po5312 = pi5205;
  assign po5313 = pi5320;
  assign po5314 = pi5266;
  assign po5315 = pi5220;
  assign po5316 = pi5246;
  assign po5317 = pi5418;
  assign po5318 = pi5333;
  assign po5319 = pi5310;
  assign po5320 = pi5332;
  assign po5321 = pi5346;
  assign po5322 = pi5343;
  assign po5323 = pi5378;
  assign po5324 = pi5336;
  assign po5325 = pi5327;
  assign po5326 = pi5338;
  assign po5327 = pi5337;
  assign po5328 = pi5512;
  assign po5329 = pi5421;
  assign po5330 = pi5345;
  assign po5331 = pi5344;
  assign po5332 = pi5335;
  assign po5333 = pi5341;
  assign po5334 = pi5330;
  assign po5335 = pi5422;
  assign po5336 = pi5334;
  assign po5337 = pi5358;
  assign po5338 = pi5348;
  assign po5339 = pi5340;
  assign po5340 = pi5292;
  assign po5341 = pi5342;
  assign po5342 = pi5392;
  assign po5343 = pi5224;
  assign po5344 = pi5209;
  assign po5345 = pi5269;
  assign po5346 = pi5416;
  assign po5347 = pi5403;
  assign po5348 = pi5197;
  assign po5349 = pi5235;
  assign po5350 = pi5243;
  assign po5351 = pi5272;
  assign po5352 = pi5264;
  assign po5353 = pi5270;
  assign po5354 = pi5260;
  assign po5355 = pi5247;
  assign po5356 = pi5271;
  assign po5357 = pi5276;
  assign po5358 = pi5261;
  assign po5359 = pi5241;
  assign po5360 = pi5236;
  assign po5361 = pi5227;
  assign po5362 = pi5237;
  assign po5363 = pi5225;
  assign po5364 = pi5263;
  assign po5365 = pi5279;
  assign po5366 = pi5198;
  assign po5367 = pi5244;
  assign po5368 = pi5228;
  assign po5369 = pi5199;
  assign po5370 = pi5258;
  assign po5371 = pi5239;
  assign po5372 = pi5218;
  assign po5373 = pi5400;
  assign po5374 = pi5408;
  assign po5375 = pi5221;
  assign po5376 = pi5200;
  assign po5377 = pi5256;
  assign po5378 = pi5222;
  assign po5379 = pi5232;
  assign po5380 = pi5251;
  assign po5381 = pi5396;
  assign po5382 = pi5398;
  assign po5383 = pi5273;
  assign po5384 = pi5304;
  assign po5385 = pi5415;
  assign po5386 = pi5401;
  assign po5387 = pi5275;
  assign po5388 = pi5248;
  assign po5389 = pi5257;
  assign po5390 = pi5240;
  assign po5391 = pi5249;
  assign po5392 = pi5274;
  assign po5393 = pi5226;
  assign po5394 = pi5407;
  assign po5395 = pi5259;
  assign po5396 = pi5219;
  assign po5397 = pi5242;
  assign po5398 = pi5231;
  assign po5399 = pi5268;
  assign po5400 = pi5254;
  assign po5401 = pi5201;
  assign po5402 = pi5265;
  assign po5403 = pi5234;
  assign po5404 = pi5233;
  assign po5405 = pi5230;
  assign po5406 = pi5223;
  assign po5407 = pi5229;
  assign po5408 = pi5430;
  assign po5409 = pi5347;
  assign po5410 = pi5294;
  assign po5411 = pi5429;
  assign po5412 = pi5434;
  assign po5413 = pi5534;
  assign po5414 = pi5326;
  assign po5415 = pi5439;
  assign po5416 = pi5282;
  assign po5417 = pi5440;
  assign po5418 = pi5402;
  assign po5419 = pi5438;
  assign po5420 = pi5399;
  assign po5421 = pi5431;
  assign po5422 = pi5442;
  assign po5423 = pi5328;
  assign po5424 = pi5441;
  assign po5425 = pi5437;
  assign po5426 = pi5436;
  assign po5427 = pi5371;
  assign po5428 = pi5373;
  assign po5429 = pi5353;
  assign po5430 = pi5423;
  assign po5431 = pi5381;
  assign po5432 = pi5446;
  assign po5433 = pi5459;
  assign po5434 = pi5450;
  assign po5435 = pi5455;
  assign po5436 = pi5461;
  assign po5437 = pi5460;
  assign po5438 = pi5456;
  assign po5439 = pi5506;
  assign po5440 = pi5458;
  assign po5441 = pi5447;
  assign po5442 = pi5454;
  assign po5443 = pi5464;
  assign po5444 = pi5453;
  assign po5445 = pi5452;
  assign po5446 = pi5585;
  assign po5447 = pi5475;
  assign po5448 = pi5372;
  assign po5449 = pi5382;
  assign po5450 = pi5406;
  assign po5451 = pi5388;
  assign po5452 = pi5374;
  assign po5453 = pi5391;
  assign po5454 = pi5424;
  assign po5455 = pi5375;
  assign po5456 = pi5331;
  assign po5457 = pi5393;
  assign po5458 = pi5413;
  assign po5459 = pi5370;
  assign po5460 = pi5412;
  assign po5461 = pi5384;
  assign po5462 = pi5425;
  assign po5463 = pi5410;
  assign po5464 = pi5329;
  assign po5465 = pi5395;
  assign po5466 = pi5411;
  assign po5467 = pi5380;
  assign po5468 = pi5465;
  assign po5469 = pi5420;
  assign po5470 = pi5361;
  assign po5471 = pi5419;
  assign po5472 = pi5417;
  assign po5473 = pi5390;
  assign po5474 = pi5394;
  assign po5475 = pi5510;
  assign po5476 = pi5351;
  assign po5477 = pi5369;
  assign po5478 = pi5404;
  assign po5479 = pi5354;
  assign po5480 = pi5443;
  assign po5481 = pi5514;
  assign po5482 = pi5502;
  assign po5483 = pi5509;
  assign po5484 = pi5377;
  assign po5485 = pi5513;
  assign po5486 = pi5409;
  assign po5487 = pi5389;
  assign po5488 = pi5367;
  assign po5489 = pi5397;
  assign po5490 = pi5366;
  assign po5491 = pi5386;
  assign po5492 = pi5511;
  assign po5493 = pi5368;
  assign po5494 = pi5357;
  assign po5495 = pi5364;
  assign po5496 = pi5385;
  assign po5497 = pi5405;
  assign po5498 = pi5365;
  assign po5499 = pi5387;
  assign po5500 = pi5360;
  assign po5501 = pi5359;
  assign po5502 = pi5379;
  assign po5503 = pi5383;
  assign po5504 = pi5362;
  assign po5505 = pi5376;
  assign po5506 = pi5414;
  assign po5507 = pi5339;
  assign po5508 = pi5355;
  assign po5509 = pi5363;
  assign po5510 = pi5607;
  assign po5511 = pi5584;
  assign po5512 = pi5543;
  assign po5513 = pi5562;
  assign po5514 = pi5538;
  assign po5515 = pi5537;
  assign po5516 = pi5539;
  assign po5517 = pi5535;
  assign po5518 = pi5547;
  assign po5519 = pi5548;
  assign po5520 = pi5583;
  assign po5521 = pi5545;
  assign po5522 = pi5533;
  assign po5523 = pi5560;
  assign po5524 = pi5536;
  assign po5525 = pi5542;
  assign po5526 = pi5449;
  assign po5527 = pi5552;
  assign po5528 = pi5530;
  assign po5529 = pi5569;
  assign po5530 = pi5586;
  assign po5531 = pi5587;
  assign po5532 = pi5566;
  assign po5533 = pi5581;
  assign po5534 = pi5563;
  assign po5535 = pi5564;
  assign po5536 = pi5578;
  assign po5537 = pi5550;
  assign po5538 = pi5555;
  assign po5539 = pi5574;
  assign po5540 = pi5575;
  assign po5541 = pi5582;
  assign po5542 = pi5505;
  assign po5543 = pi5553;
  assign po5544 = pi5576;
  assign po5545 = pi5573;
  assign po5546 = pi5579;
  assign po5547 = pi5554;
  assign po5548 = pi5571;
  assign po5549 = pi5580;
  assign po5550 = pi5577;
  assign po5551 = pi5559;
  assign po5552 = pi5558;
  assign po5553 = pi5557;
  assign po5554 = pi5556;
  assign po5555 = pi5568;
  assign po5556 = pi5435;
  assign po5557 = pi5544;
  assign po5558 = pi5663;
  assign po5559 = pi5527;
  assign po5560 = pi5619;
  assign po5561 = pi5526;
  assign po5563 = pi5606;
  assign po5564 = pi5626;
  assign po5565 = pi5608;
  assign po5566 = pi5541;
  assign po5567 = pi5532;
  assign po5568 = pi5624;
  assign po5569 = pi5630;
  assign po5570 = pi5631;
  assign po5571 = pi5616;
  assign po5572 = pi5641;
  assign po5573 = pi5662;
  assign po5574 = pi5625;
  assign po5575 = pi5636;
  assign po5576 = pi5549;
  assign po5577 = pi5668;
  assign po5578 = pi5609;
  assign po5579 = pi5598;
  assign po5580 = pi5658;
  assign po5581 = pi5504;
  assign po5582 = pi5650;
  assign po5583 = pi5472;
  assign po5584 = pi5468;
  assign po5585 = pi5665;
  assign po5586 = pi5703;
  assign po5587 = pi5503;
  assign po5588 = pi5634;
  assign po5589 = pi5491;
  assign po5590 = pi5500;
  assign po5591 = pi5496;
  assign po5592 = pi5477;
  assign po5593 = pi5525;
  assign po5594 = pi5470;
  assign po5595 = pi5501;
  assign po5596 = pi5490;
  assign po5597 = pi5489;
  assign po5598 = pi5469;
  assign po5599 = pi5462;
  assign po5600 = pi5507;
  assign po5601 = pi5520;
  assign po5602 = pi5494;
  assign po5603 = pi5515;
  assign po5604 = pi5482;
  assign po5605 = pi5480;
  assign po5606 = pi5445;
  assign po5607 = pi5483;
  assign po5608 = pi5618;
  assign po5609 = pi5516;
  assign po5610 = pi5484;
  assign po5611 = pi5474;
  assign po5612 = pi5519;
  assign po5613 = pi5528;
  assign po5614 = pi5448;
  assign po5615 = pi5488;
  assign po5616 = pi5522;
  assign po5617 = pi5485;
  assign po5618 = pi5466;
  assign po5619 = pi5521;
  assign po5620 = pi5498;
  assign po5621 = pi5495;
  assign po5622 = pi5666;
  assign po5623 = pi5451;
  assign po5624 = pi5518;
  assign po5625 = pi5486;
  assign po5626 = pi5664;
  assign po5627 = pi5479;
  assign po5628 = pi5671;
  assign po5629 = pi5561;
  assign po5630 = pi5669;
  assign po5631 = pi5661;
  assign po5632 = pi5572;
  assign po5633 = pi5677;
  assign po5634 = pi5463;
  assign po5636 = pi5529;
  assign po5637 = pi5672;
  assign po5638 = pi5667;
  assign po5639 = pi5492;
  assign po5640 = pi5471;
  assign po5641 = pi5524;
  assign po5642 = pi5473;
  assign po5643 = pi5481;
  assign po5644 = pi5493;
  assign po5645 = pi5588;
  assign po5646 = pi5508;
  assign po5647 = pi5478;
  assign po5648 = pi5628;
  assign po5649 = pi5444;
  assign po5650 = pi5517;
  assign po5651 = pi5633;
  assign po5652 = pi5540;
  assign po5653 = pi5457;
  assign po5654 = pi5487;
  assign po5655 = pi5476;
  assign po5656 = pi5674;
  assign po5657 = pi5694;
  assign po5658 = pi5692;
  assign po5659 = pi5687;
  assign po5660 = pi5670;
  assign po5662 = pi5693;
  assign po5663 = pi5690;
  assign po5664 = pi5699;
  assign po5665 = pi5704;
  assign po5666 = pi5698;
  assign po5667 = pi5706;
  assign po5668 = pi5695;
  assign po5669 = pi5570;
  assign po5670 = pi5565;
  assign po5671 = pi5697;
  assign po5672 = pi5701;
  assign po5673 = pi5696;
  assign po5674 = pi5591;
  assign po5675 = pi5610;
  assign po5677 = pi5738;
  assign po5678 = pi5644;
  assign po5679 = pi5747;
  assign po5680 = pi5781;
  assign po5681 = pi5604;
  assign po5682 = pi5746;
  assign po5683 = pi5741;
  assign po5684 = pi5723;
  assign po5685 = pi5735;
  assign po5686 = pi5740;
  assign po5687 = pi5680;
  assign po5688 = pi5736;
  assign po5689 = pi5737;
  assign po5690 = pi5727;
  assign po5691 = pi5734;
  assign po5692 = pi5635;
  assign po5693 = pi5649;
  assign po5694 = pi5732;
  assign po5696 = pi5657;
  assign po5697 = pi5750;
  assign po5698 = pi5640;
  assign po5699 = pi5659;
  assign po5700 = pi5652;
  assign po5701 = pi5648;
  assign po5702 = pi5600;
  assign po5703 = pi5601;
  assign po5704 = pi5681;
  assign po5706 = pi5622;
  assign po5707 = pi5639;
  assign po5708 = pi5612;
  assign po5709 = pi5593;
  assign po5710 = pi5673;
  assign po5711 = pi5642;
  assign po5712 = pi5654;
  assign po5713 = pi5637;
  assign po5714 = pi5653;
  assign po5715 = pi5595;
  assign po5716 = pi5632;
  assign po5717 = pi5660;
  assign po5718 = pi5638;
  assign po5719 = pi5602;
  assign po5720 = pi5617;
  assign po5721 = pi5597;
  assign po5722 = pi5605;
  assign po5723 = pi5678;
  assign po5724 = pi5589;
  assign po5725 = pi5623;
  assign po5726 = pi5590;
  assign po5728 = pi5655;
  assign po5729 = pi5748;
  assign po5730 = pi5643;
  assign po5731 = pi5682;
  assign po5732 = pi5779;
  assign po5733 = pi5676;
  assign po5734 = pi5683;
  assign po5735 = pi5700;
  assign po5736 = pi5722;
  assign po5737 = pi5679;
  assign po5738 = pi5675;
  assign po5739 = pi5784;
  assign po5740 = pi5782;
  assign po5741 = pi5783;
  assign po5743 = pi5780;
  assign po5744 = pi5785;
  assign po5745 = pi5627;
  assign po5746 = pi5594;
  assign po5747 = pi5621;
  assign po5748 = pi5645;
  assign po5749 = pi5614;
  assign po5750 = pi5596;
  assign po5751 = pi5592;
  assign po5752 = pi5651;
  assign po5753 = pi5749;
  assign po5754 = pi5611;
  assign po5755 = pi5620;
  assign po5756 = pi5615;
  assign po5757 = pi5656;
  assign po5758 = pi5629;
  assign po5759 = pi5613;
  assign po5760 = pi5814;
  assign po5761 = pi5841;
  assign po5762 = pi5810;
  assign po5763 = pi5800;
  assign po5765 = pi5743;
  assign po5766 = pi5807;
  assign po5767 = pi5811;
  assign po5768 = pi5801;
  assign po5769 = pi5806;
  assign po5770 = pi5839;
  assign po5771 = pi5812;
  assign po5772 = pi5688;
  assign po5773 = pi5802;
  assign po5774 = pi5808;
  assign po5775 = pi5794;
  assign po5776 = pi5793;
  assign po5777 = pi5791;
  assign po5778 = pi5803;
  assign po5779 = pi5797;
  assign po5781 = pi5805;
  assign po5782 = pi5745;
  assign po5783 = pi5840;
  assign po5784 = pi5824;
  assign po5785 = pi5837;
  assign po5786 = pi5820;
  assign po5787 = pi5792;
  assign po5788 = pi5829;
  assign po5789 = pi5832;
  assign po5790 = pi5823;
  assign po5791 = pi5818;
  assign po5792 = pi5804;
  assign po5793 = pi5836;
  assign po5794 = pi5828;
  assign po5795 = pi5705;
  assign po5796 = pi5830;
  assign po5797 = pi5833;
  assign po5798 = pi5827;
  assign po5799 = pi5822;
  assign po5800 = pi5702;
  assign po5801 = pi5843;
  assign po5802 = pi5831;
  assign po5803 = pi5826;
  assign po5804 = pi5825;
  assign po5805 = pi5838;
  assign po5806 = pi5834;
  assign po5807 = pi5842;
  assign po5808 = pi5817;
  assign po5809 = pi5796;
  assign po5810 = pi5819;
  assign po5811 = pi5815;
  assign po5812 = pi5821;
  assign po5813 = pi5685;
  assign po5814 = pi5686;
  assign po5818 = pi5909;
  assign po5819 = pi5708;
  assign po5820 = pi5773;
  assign po5821 = pi5728;
  assign po5822 = pi5719;
  assign po5823 = pi5761;
  assign po5824 = pi5718;
  assign po5825 = pi5726;
  assign po5826 = pi5790;
  assign po5827 = pi5721;
  assign po5829 = pi5856;
  assign po5830 = pi5709;
  assign po5831 = pi5716;
  assign po5832 = pi5768;
  assign po5833 = pi5888;
  assign po5834 = pi5769;
  assign po5835 = pi5766;
  assign po5836 = pi5884;
  assign po5838 = pi5879;
  assign po5839 = pi5799;
  assign po5840 = pi5730;
  assign po5841 = pi5714;
  assign po5842 = pi5786;
  assign po5843 = pi5752;
  assign po5844 = pi5758;
  assign po5845 = pi5755;
  assign po5846 = pi5874;
  assign po5847 = pi5753;
  assign po5848 = pi5862;
  assign po5849 = pi5871;
  assign po5850 = pi5754;
  assign po5851 = pi5772;
  assign po5852 = pi5789;
  assign po5853 = pi5707;
  assign po5854 = pi5877;
  assign po5855 = pi5849;
  assign po5856 = pi5873;
  assign po5857 = pi5765;
  assign po5858 = pi5742;
  assign po5859 = pi5763;
  assign po5860 = pi5733;
  assign po5861 = pi5844;
  assign po5862 = pi5762;
  assign po5863 = pi5910;
  assign po5864 = pi5725;
  assign po5865 = pi5757;
  assign po5866 = pi5891;
  assign po5867 = pi5776;
  assign po5868 = pi5744;
  assign po5869 = pi5777;
  assign po5870 = pi5731;
  assign po5871 = pi5878;
  assign po5872 = pi5770;
  assign po5873 = pi5712;
  assign po5874 = pi5774;
  assign po5875 = pi5739;
  assign po5876 = pi5895;
  assign po5877 = pi5798;
  assign po5878 = pi5713;
  assign po5879 = pi5767;
  assign po5881 = pi5764;
  assign po5882 = pi5720;
  assign po5883 = pi5788;
  assign po5884 = pi5724;
  assign po5885 = pi5751;
  assign po5886 = pi5759;
  assign po5887 = pi5787;
  assign po5889 = pi5717;
  assign po5890 = pi5778;
  assign po5891 = pi5929;
  assign po5892 = pi5809;
  assign po5893 = pi5921;
  assign po5894 = pi5916;
  assign po5895 = pi5919;
  assign po5897 = pi5918;
  assign po5898 = pi5881;
  assign po5899 = pi5920;
  assign po5900 = pi5883;
  assign po5901 = pi5922;
  assign po5902 = pi5913;
  assign po5903 = pi5710;
  assign po5905 = pi5911;
  assign po5906 = pi5715;
  assign po5907 = pi5923;
  assign po5908 = pi5771;
  assign po5909 = pi5760;
  assign po5910 = pi5729;
  assign po5911 = pi5711;
  assign po5912 = pi5775;
  assign po5913 = pi5756;
  assign po5915 = pi5944;
  assign po5916 = pi5934;
  assign po5917 = pi5932;
  assign po5918 = pi5936;
  assign po5919 = pi5813;
  assign po5921 = pi5795;
  assign po5925 = pi5947;
  assign po5926 = pi5940;
  assign po5927 = pi5942;
  assign po5928 = pi5946;
  assign po5929 = pi5938;
  assign po5930 = pi5937;
  assign po5931 = pi5943;
  assign po5932 = pi5941;
  assign po5934 = pi5816;
  assign po5935 = pi5945;
  assign po5936 = pi5948;
  assign po5937 = pi5887;
  assign po5938 = pi5861;
  assign po5939 = pi5925;
  assign po5940 = pi5889;
  assign po5941 = pi5885;
  assign po5942 = pi5864;
  assign po5943 = pi5872;
  assign po5944 = pi5869;
  assign po5945 = pi5880;
  assign po5946 = pi5852;
  assign po5947 = pi5894;
  assign po5948 = pi5846;
  assign po5949 = pi5853;
  assign po5950 = pi5892;
  assign po5951 = pi5890;
  assign po5952 = pi5951;
  assign po5953 = pi5956;
  assign po5954 = pi5851;
  assign po5955 = pi6010;
  assign po5956 = pi5845;
  assign po5957 = pi6007;
  assign po5958 = pi5901;
  assign po5959 = pi5903;
  assign po5960 = pi5899;
  assign po5961 = pi5866;
  assign po5962 = pi5963;
  assign po5963 = pi6002;
  assign po5964 = pi6016;
  assign po5965 = pi5952;
  assign po5966 = pi5882;
  assign po5967 = pi6017;
  assign po5968 = pi5931;
  assign po5969 = pi5886;
  assign po5970 = pi5933;
  assign po5971 = pi5965;
  assign po5972 = pi6011;
  assign po5973 = pi5991;
  assign po5974 = pi5867;
  assign po5975 = pi5964;
  assign po5976 = pi5960;
  assign po5977 = pi6025;
  assign po5981 = pi5865;
  assign po5982 = pi5847;
  assign po5983 = pi5855;
  assign po5984 = pi5860;
  assign po5985 = pi5904;
  assign po5986 = pi5870;
  assign po5987 = pi5930;
  assign po5988 = pi5905;
  assign po5989 = pi5854;
  assign po5990 = pi5908;
  assign po5991 = pi5897;
  assign po5992 = pi5926;
  assign po5993 = pi5896;
  assign po5994 = pi5928;
  assign po5995 = pi5848;
  assign po5996 = pi5858;
  assign po5997 = pi5898;
  assign po5998 = pi5893;
  assign po5999 = pi5914;
  assign po6000 = pi5907;
  assign po6001 = pi5863;
  assign po6002 = pi5924;
  assign po6003 = pi5900;
  assign po6004 = pi5927;
  assign po6005 = pi5859;
  assign po6006 = pi5876;
  assign po6007 = pi5850;
  assign po6008 = pi5906;
  assign po6009 = pi5917;
  assign po6010 = pi5939;
  assign po6011 = pi5950;
  assign po6012 = pi6013;
  assign po6013 = pi6015;
  assign po6014 = pi6012;
  assign po6015 = pi5915;
  assign po6016 = pi5868;
  assign po6017 = pi5912;
  assign po6018 = pi5875;
  assign po6019 = pi5857;
  assign po6020 = pi5902;
  assign po6021 = pi6043;
  assign po6022 = pi6058;
  assign po6023 = pi5935;
  assign po6024 = pi6036;
  assign po6026 = pi6050;
  assign po6027 = pi6029;
  assign po6029 = pi6042;
  assign po6030 = pi6044;
  assign po6031 = pi6032;
  assign po6032 = pi6037;
  assign po6033 = pi6068;
  assign po6034 = pi6073;
  assign po6036 = pi6047;
  assign po6037 = pi6074;
  assign po6038 = pi6045;
  assign po6039 = pi6033;
  assign po6040 = pi6030;
  assign po6041 = pi6075;
  assign po6042 = pi6048;
  assign po6044 = pi6034;
  assign po6045 = pi6038;
  assign po6046 = pi6057;
  assign po6047 = pi6035;
  assign po6048 = pi6084;
  assign po6049 = pi6041;
  assign po6050 = pi6060;
  assign po6051 = pi6031;
  assign po6052 = pi6082;
  assign po6053 = pi6071;
  assign po6054 = pi6026;
  assign po6055 = pi6056;
  assign po6056 = pi6076;
  assign po6057 = pi6078;
  assign po6058 = pi6053;
  assign po6059 = pi6062;
  assign po6060 = pi6080;
  assign po6061 = pi6066;
  assign po6062 = pi6059;
  assign po6063 = pi6051;
  assign po6064 = pi6069;
  assign po6065 = pi6063;
  assign po6066 = pi6070;
  assign po6067 = pi6081;
  assign po6068 = pi6052;
  assign po6069 = pi6046;
  assign po6070 = pi6064;
  assign po6072 = pi6067;
  assign po6073 = pi6027;
  assign po6074 = pi6139;
  assign po6075 = pi6005;
  assign po6076 = pi5992;
  assign po6077 = pi6001;
  assign po6078 = pi5969;
  assign po6079 = pi6089;
  assign po6080 = pi5961;
  assign po6081 = pi5997;
  assign po6082 = pi5987;
  assign po6083 = pi6019;
  assign po6084 = pi5959;
  assign po6085 = pi5989;
  assign po6087 = pi5966;
  assign po6088 = pi6022;
  assign po6089 = pi6021;
  assign po6090 = pi5995;
  assign po6091 = pi6024;
  assign po6092 = pi6040;
  assign po6093 = pi5974;
  assign po6094 = pi5990;
  assign po6095 = pi5970;
  assign po6096 = pi5980;
  assign po6097 = pi5982;
  assign po6098 = pi5993;
  assign po6099 = pi5958;
  assign po6100 = pi5967;
  assign po6101 = pi6093;
  assign po6102 = pi6023;
  assign po6103 = pi6094;
  assign po6104 = pi6142;
  assign po6105 = pi5978;
  assign po6106 = pi6009;
  assign po6107 = pi6079;
  assign po6108 = pi6018;
  assign po6109 = pi6124;
  assign po6110 = pi5979;
  assign po6111 = pi6121;
  assign po6112 = pi6158;
  assign po6113 = pi6144;
  assign po6114 = pi6072;
  assign po6115 = pi5976;
  assign po6116 = pi5957;
  assign po6117 = pi6008;
  assign po6119 = pi6014;
  assign po6120 = pi5994;
  assign po6121 = pi6088;
  assign po6122 = pi5968;
  assign po6123 = pi5962;
  assign po6124 = pi6003;
  assign po6126 = pi5973;
  assign po6127 = pi5985;
  assign po6128 = pi6020;
  assign po6129 = pi5984;
  assign po6130 = pi5954;
  assign po6131 = pi5972;
  assign po6132 = pi5975;
  assign po6133 = pi5971;
  assign po6134 = pi5981;
  assign po6135 = pi6006;
  assign po6136 = pi5988;
  assign po6137 = pi5999;
  assign po6138 = pi5986;
  assign po6139 = pi6148;
  assign po6140 = pi6039;
  assign po6141 = pi6159;
  assign po6142 = pi5983;
  assign po6143 = pi6061;
  assign po6144 = pi6004;
  assign po6145 = pi6150;
  assign po6146 = pi6133;
  assign po6147 = pi6154;
  assign po6148 = pi6147;
  assign po6149 = pi5949;
  assign po6150 = pi6152;
  assign po6151 = pi6143;
  assign po6152 = pi6149;
  assign po6153 = pi6151;
  assign po6154 = pi5955;
  assign po6155 = pi5977;
  assign po6156 = pi5998;
  assign po6157 = pi6000;
  assign po6158 = pi5996;
  assign po6159 = pi6153;
  assign po6160 = pi5953;
  assign po6161 = pi6146;
  assign po6162 = pi6165;
  assign po6163 = pi6086;
  assign po6164 = pi6167;
  assign po6165 = pi6166;
  assign po6166 = pi6028;
  assign po6167 = pi6077;
  assign po6168 = pi6049;
  assign po6169 = pi6055;
  assign po6170 = pi6169;
  assign po6171 = pi6083;
  assign po6172 = pi6168;
  assign po6173 = pi6174;
  assign po6174 = pi6173;
  assign po6175 = pi6175;
  assign po6176 = pi6176;
  assign po6177 = pi6065;
  assign po6178 = pi6054;
  assign po6179 = pi6259;
  assign po6180 = pi6258;
  assign po6181 = pi6256;
  assign po6182 = pi6227;
  assign po6183 = pi6107;
  assign po6184 = pi6162;
  assign po6185 = pi6120;
  assign po6186 = pi6245;
  assign po6187 = pi6131;
  assign po6188 = pi6100;
  assign po6189 = pi6110;
  assign po6190 = pi6232;
  assign po6191 = pi6119;
  assign po6192 = pi6116;
  assign po6193 = pi6234;
  assign po6194 = pi6228;
  assign po6195 = pi6255;
  assign po6196 = pi6097;
  assign po6197 = pi6108;
  assign po6198 = pi6122;
  assign po6199 = pi6087;
  assign po6200 = pi6134;
  assign po6201 = pi6125;
  assign po6202 = pi6099;
  assign po6203 = pi6114;
  assign po6204 = pi6090;
  assign po6205 = pi6104;
  assign po6206 = pi6155;
  assign po6207 = pi6128;
  assign po6208 = pi6117;
  assign po6209 = pi6130;
  assign po6210 = pi6160;
  assign po6211 = pi6106;
  assign po6212 = pi6157;
  assign po6213 = pi6109;
  assign po6214 = pi6096;
  assign po6215 = pi6115;
  assign po6216 = pi6129;
  assign po6217 = pi6127;
  assign po6218 = pi6091;
  assign po6219 = pi6101;
  assign po6220 = pi6113;
  assign po6221 = pi6244;
  assign po6222 = pi6095;
  assign po6223 = pi6135;
  assign po6224 = pi6140;
  assign po6225 = pi6103;
  assign po6226 = pi6141;
  assign po6227 = pi6112;
  assign po6228 = pi6156;
  assign po6229 = pi6098;
  assign po6230 = pi6085;
  assign po6231 = pi6132;
  assign po6232 = pi6183;
  assign po6233 = pi6138;
  assign po6234 = pi6137;
  assign po6235 = pi6163;
  assign po6236 = pi6102;
  assign po6237 = pi6242;
  assign po6238 = pi6111;
  assign po6239 = pi6123;
  assign po6240 = pi6231;
  assign po6241 = pi6179;
  assign po6242 = pi6225;
  assign po6243 = pi6233;
  assign po6244 = pi6105;
  assign po6245 = pi6257;
  assign po6246 = pi6241;
  assign po6247 = pi6188;
  assign po6248 = pi6145;
  assign po6249 = pi6092;
  assign po6250 = pi6136;
  assign po6251 = pi6161;
  assign po6252 = pi6164;
  assign po6253 = pi6118;
  assign po6254 = pi6126;
  assign po6255 = pi6243;
  assign po6256 = pi6296;
  assign po6257 = pi6311;
  assign po6258 = pi6266;
  assign po6259 = pi6262;
  assign po6260 = pi6264;
  assign po6261 = pi6260;
  assign po6262 = pi6310;
  assign po6263 = pi6172;
  assign po6264 = pi6273;
  assign po6265 = pi6281;
  assign po6266 = pi6275;
  assign po6267 = pi6170;
  assign po6268 = pi6287;
  assign po6269 = pi6240;
  assign po6270 = pi6181;
  assign po6271 = pi6280;
  assign po6272 = pi6305;
  assign po6273 = pi6279;
  assign po6274 = pi6269;
  assign po6275 = pi6171;
  assign po6276 = pi6283;
  assign po6277 = pi6246;
  assign po6278 = pi6248;
  assign po6279 = pi6286;
  assign po6280 = pi6261;
  assign po6281 = pi6289;
  assign po6282 = pi6313;
  assign po6283 = pi6282;
  assign po6284 = pi6306;
  assign po6285 = pi6277;
  assign po6286 = pi6314;
  assign po6287 = pi6300;
  assign po6288 = pi6270;
  assign po6289 = pi6285;
  assign po6290 = pi6263;
  assign po6291 = pi6304;
  assign po6292 = pi6268;
  assign po6293 = pi6288;
  assign po6294 = pi6284;
  assign po6295 = pi6278;
  assign po6296 = pi6271;
  assign po6297 = pi6290;
  assign po6298 = pi6276;
  assign po6299 = pi6294;
  assign po6300 = pi6308;
  assign po6301 = pi6292;
  assign po6302 = pi6177;
  assign po6303 = pi6302;
  assign po6304 = pi6303;
  assign po6305 = pi6301;
  assign po6306 = pi6298;
  assign po6307 = pi6309;
  assign po6308 = pi6272;
  assign po6309 = pi6247;
  assign po6310 = pi6297;
  assign po6311 = pi6291;
  assign po6312 = pi6295;
  assign po6313 = pi6293;
  assign po6314 = pi6307;
  assign po6315 = pi6194;
  assign po6316 = pi6274;
  assign po6317 = pi6199;
  assign po6318 = pi6393;
  assign po6319 = pi6384;
  assign po6320 = pi6216;
  assign po6321 = pi6250;
  assign po6322 = pi6222;
  assign po6323 = pi6366;
  assign po6324 = pi6385;
  assign po6325 = pi6226;
  assign po6326 = pi6219;
  assign po6327 = pi6211;
  assign po6328 = pi6223;
  assign po6329 = pi6193;
  assign po6330 = pi6251;
  assign po6331 = pi6195;
  assign po6332 = pi6235;
  assign po6333 = pi6205;
  assign po6334 = pi6184;
  assign po6335 = pi6230;
  assign po6336 = pi6229;
  assign po6337 = pi6237;
  assign po6338 = pi6212;
  assign po6339 = pi6238;
  assign po6340 = pi6218;
  assign po6341 = pi6224;
  assign po6342 = pi6203;
  assign po6343 = pi6221;
  assign po6344 = pi6190;
  assign po6345 = pi6239;
  assign po6346 = pi6191;
  assign po6347 = pi6249;
  assign po6348 = pi6208;
  assign po6349 = pi6186;
  assign po6350 = pi6214;
  assign po6351 = pi6320;
  assign po6352 = pi6187;
  assign po6353 = pi6196;
  assign po6354 = pi6379;
  assign po6355 = pi6189;
  assign po6356 = pi6252;
  assign po6357 = pi6207;
  assign po6358 = pi6198;
  assign po6359 = pi6206;
  assign po6360 = pi6185;
  assign po6361 = pi6180;
  assign po6362 = pi6253;
  assign po6363 = pi6372;
  assign po6364 = pi6220;
  assign po6365 = pi6200;
  assign po6366 = pi6217;
  assign po6367 = pi6178;
  assign po6368 = pi6213;
  assign po6369 = pi6392;
  assign po6370 = pi6192;
  assign po6371 = pi6202;
  assign po6372 = pi6373;
  assign po6373 = pi6367;
  assign po6374 = pi6377;
  assign po6375 = pi6365;
  assign po6376 = pi6265;
  assign po6377 = pi6374;
  assign po6378 = pi6322;
  assign po6379 = pi6312;
  assign po6381 = pi6319;
  assign po6382 = pi6375;
  assign po6383 = pi6369;
  assign po6384 = pi6382;
  assign po6385 = pi6210;
  assign po6386 = pi6201;
  assign po6387 = pi6182;
  assign po6388 = pi6204;
  assign po6389 = pi6368;
  assign po6390 = pi6209;
  assign po6391 = pi6197;
  assign po6392 = pi6236;
  assign po6393 = pi6215;
  assign po6394 = pi6254;
  assign po6395 = pi6381;
  assign po6396 = pi6398;
  assign po6397 = pi6400;
  assign po6398 = pi6397;
  assign po6399 = pi6402;
  assign po6401 = pi6267;
  assign po6402 = pi6299;
  assign po6403 = pi6399;
  assign po6404 = pi6396;
  assign po6405 = pi6395;
  assign po6406 = pi6401;
  assign po6407 = pi6464;
  assign po6408 = pi6333;
  assign po6409 = pi6407;
  assign po6410 = pi6371;
  assign po6411 = pi6480;
  assign po6412 = pi6335;
  assign po6413 = pi6469;
  assign po6414 = pi6356;
  assign po6415 = pi6344;
  assign po6416 = pi6358;
  assign po6417 = pi6359;
  assign po6418 = pi6485;
  assign po6419 = pi6345;
  assign po6420 = pi6342;
  assign po6421 = pi6350;
  assign po6422 = pi6378;
  assign po6423 = pi6394;
  assign po6424 = pi6380;
  assign po6425 = pi6326;
  assign po6426 = pi6391;
  assign po6427 = pi6390;
  assign po6428 = pi6346;
  assign po6429 = pi6351;
  assign po6430 = pi6318;
  assign po6431 = pi6325;
  assign po6432 = pi6338;
  assign po6433 = pi6364;
  assign po6434 = pi6387;
  assign po6435 = pi6330;
  assign po6436 = pi6334;
  assign po6437 = pi6389;
  assign po6438 = pi6388;
  assign po6439 = pi6340;
  assign po6440 = pi6339;
  assign po6441 = pi6341;
  assign po6442 = pi6357;
  assign po6443 = pi6316;
  assign po6444 = pi6332;
  assign po6445 = pi6353;
  assign po6446 = pi6361;
  assign po6447 = pi6355;
  assign po6448 = pi6348;
  assign po6449 = pi6354;
  assign po6450 = pi6323;
  assign po6451 = pi6328;
  assign po6452 = pi6331;
  assign po6453 = pi6349;
  assign po6454 = pi6343;
  assign po6455 = pi6467;
  assign po6456 = pi6386;
  assign po6457 = pi6483;
  assign po6458 = pi6481;
  assign po6459 = pi6362;
  assign po6460 = pi6327;
  assign po6461 = pi6419;
  assign po6462 = pi6409;
  assign po6463 = pi6466;
  assign po6464 = pi6408;
  assign po6465 = pi6317;
  assign po6466 = pi6337;
  assign po6467 = pi6324;
  assign po6468 = pi6321;
  assign po6469 = pi6363;
  assign po6470 = pi6404;
  assign po6471 = pi6472;
  assign po6472 = pi6465;
  assign po6473 = pi6468;
  assign po6474 = pi6405;
  assign po6475 = pi6460;
  assign po6476 = pi6461;
  assign po6477 = pi6421;
  assign po6478 = pi6484;
  assign po6479 = pi6360;
  assign po6480 = pi6347;
  assign po6481 = pi6336;
  assign po6482 = pi6329;
  assign po6483 = pi6370;
  assign po6484 = pi6352;
  assign po6485 = pi6463;
  assign po6486 = pi6474;
  assign po6487 = pi6403;
  assign po6488 = pi6416;
  assign po6489 = pi6376;
  assign po6490 = pi6525;
  assign po6491 = pi6521;
  assign po6492 = pi6499;
  assign po6493 = pi6517;
  assign po6494 = pi6491;
  assign po6495 = pi6470;
  assign po6496 = pi6538;
  assign po6497 = pi6495;
  assign po6498 = pi6539;
  assign po6499 = pi6501;
  assign po6500 = pi6526;
  assign po6501 = pi6536;
  assign po6502 = pi6516;
  assign po6503 = pi6542;
  assign po6504 = pi6503;
  assign po6505 = pi6537;
  assign po6506 = pi6498;
  assign po6507 = pi6530;
  assign po6508 = pi6497;
  assign po6509 = pi6500;
  assign po6510 = pi6490;
  assign po6511 = pi6519;
  assign po6512 = pi6512;
  assign po6513 = pi6507;
  assign po6514 = pi6524;
  assign po6515 = pi6487;
  assign po6516 = pi6518;
  assign po6517 = pi6520;
  assign po6518 = pi6488;
  assign po6519 = pi6509;
  assign po6520 = pi6486;
  assign po6521 = pi6515;
  assign po6522 = pi6489;
  assign po6523 = pi6527;
  assign po6524 = pi6533;
  assign po6525 = pi6529;
  assign po6526 = pi6493;
  assign po6527 = pi6531;
  assign po6528 = pi6535;
  assign po6529 = pi6508;
  assign po6530 = pi6543;
  assign po6531 = pi6494;
  assign po6532 = pi6541;
  assign po6533 = pi6514;
  assign po6534 = pi6532;
  assign po6535 = pi6504;
  assign po6536 = pi6510;
  assign po6537 = pi6496;
  assign po6538 = pi6522;
  assign po6539 = pi6513;
  assign po6540 = pi6502;
  assign po6541 = pi6540;
  assign po6542 = pi6511;
  assign po6543 = pi6534;
  assign po6544 = pi6523;
  assign po6545 = pi6528;
  assign po6546 = pi6415;
  assign po6547 = pi6452;
  assign po6548 = pi6438;
  assign po6549 = pi6546;
  assign po6550 = pi6551;
  assign po6551 = pi6445;
  assign po6552 = pi6492;
  assign po6553 = pi6475;
  assign po6554 = pi6476;
  assign po6555 = pi6430;
  assign po6556 = pi6447;
  assign po6557 = pi6434;
  assign po6558 = pi6448;
  assign po6559 = pi6477;
  assign po6560 = pi6429;
  assign po6561 = pi6424;
  assign po6562 = pi6453;
  assign po6563 = pi6455;
  assign po6564 = pi6446;
  assign po6565 = pi6482;
  assign po6566 = pi6444;
  assign po6567 = pi6454;
  assign po6568 = pi6436;
  assign po6569 = pi6457;
  assign po6570 = pi6478;
  assign po6571 = pi6442;
  assign po6572 = pi6410;
  assign po6573 = pi6450;
  assign po6574 = pi6417;
  assign po6575 = pi6420;
  assign po6576 = pi6462;
  assign po6577 = pi6458;
  assign po6578 = pi6471;
  assign po6579 = pi6433;
  assign po6580 = pi6432;
  assign po6581 = pi6473;
  assign po6582 = pi6437;
  assign po6583 = pi6428;
  assign po6584 = pi6426;
  assign po6585 = pi6479;
  assign po6586 = pi6435;
  assign po6587 = pi6441;
  assign po6588 = pi6443;
  assign po6589 = pi6413;
  assign po6590 = pi6431;
  assign po6591 = pi6412;
  assign po6592 = pi6411;
  assign po6593 = pi6406;
  assign po6594 = pi6423;
  assign po6595 = pi6459;
  assign po6596 = pi6613;
  assign po6597 = pi6606;
  assign po6598 = pi6621;
  assign po6599 = pi6609;
  assign po6600 = pi6439;
  assign po6601 = pi6414;
  assign po6602 = pi6600;
  assign po6603 = pi6506;
  assign po6604 = pi6605;
  assign po6605 = pi6607;
  assign po6606 = pi6608;
  assign po6607 = pi6603;
  assign po6608 = pi6427;
  assign po6609 = pi6577;
  assign po6610 = pi6456;
  assign po6611 = pi6598;
  assign po6612 = pi6620;
  assign po6613 = pi6555;
  assign po6614 = pi6610;
  assign po6615 = pi6599;
  assign po6616 = pi6425;
  assign po6617 = pi6619;
  assign po6618 = pi6449;
  assign po6619 = pi6418;
  assign po6620 = pi6422;
  assign po6621 = pi6451;
  assign po6622 = pi6602;
  assign po6623 = pi6604;
  assign po6624 = pi6440;
  assign po6625 = pi6544;
  assign po6626 = pi6628;
  assign po6627 = pi6626;
  assign po6628 = pi6505;
  assign po6629 = pi6627;
  assign po6630 = pi6614;
  assign po6631 = pi6623;
  assign po6632 = pi6625;
  assign po6633 = pi6629;
  assign po6634 = pi6655;
  assign po6635 = pi6634;
  assign po6636 = pi6596;
  assign po6637 = pi6637;
  assign po6638 = pi6663;
  assign po6639 = pi6661;
  assign po6640 = pi6574;
  assign po6641 = pi6553;
  assign po6642 = pi6554;
  assign po6643 = pi6581;
  assign po6644 = pi6587;
  assign po6645 = pi6569;
  assign po6646 = pi6699;
  assign po6647 = pi6617;
  assign po6648 = pi6547;
  assign po6649 = pi6676;
  assign po6650 = pi6575;
  assign po6651 = pi6664;
  assign po6652 = pi6572;
  assign po6653 = pi6582;
  assign po6654 = pi6563;
  assign po6655 = pi6585;
  assign po6656 = pi6568;
  assign po6657 = pi6584;
  assign po6658 = pi6612;
  assign po6659 = pi6616;
  assign po6660 = pi6601;
  assign po6661 = pi6590;
  assign po6662 = pi6618;
  assign po6663 = pi6565;
  assign po6664 = pi6545;
  assign po6665 = pi6611;
  assign po6666 = pi6579;
  assign po6667 = pi6567;
  assign po6668 = pi6583;
  assign po6669 = pi6566;
  assign po6670 = pi6556;
  assign po6671 = pi6578;
  assign po6672 = pi6558;
  assign po6673 = pi6562;
  assign po6674 = pi6580;
  assign po6675 = pi6549;
  assign po6676 = pi6589;
  assign po6677 = pi6595;
  assign po6678 = pi6548;
  assign po6679 = pi6571;
  assign po6680 = pi6592;
  assign po6681 = pi6560;
  assign po6682 = pi6573;
  assign po6683 = pi6576;
  assign po6684 = pi6557;
  assign po6685 = pi6597;
  assign po6686 = pi6550;
  assign po6687 = pi6586;
  assign po6688 = pi6564;
  assign po6689 = pi6671;
  assign po6690 = pi6667;
  assign po6691 = pi6673;
  assign po6692 = pi6559;
  assign po6693 = pi6658;
  assign po6694 = pi6674;
  assign po6695 = pi6660;
  assign po6696 = pi6695;
  assign po6697 = pi6693;
  assign po6698 = pi6669;
  assign po6699 = pi6680;
  assign po6700 = pi6681;
  assign po6701 = pi6552;
  assign po6702 = pi6698;
  assign po6703 = pi6615;
  assign po6704 = pi6707;
  assign po6705 = pi6591;
  assign po6706 = pi6594;
  assign po6707 = pi6593;
  assign po6708 = pi6588;
  assign po6709 = pi6570;
  assign po6710 = pi6670;
  assign po6711 = pi6662;
  assign po6712 = pi6561;
  assign po6713 = pi6632;
  assign po6714 = pi6668;
  assign po6715 = pi6684;
  assign po6716 = pi6758;
  assign po6717 = pi6749;
  assign po6718 = pi6724;
  assign po6719 = pi6755;
  assign po6720 = pi6771;
  assign po6721 = pi6672;
  assign po6722 = pi6779;
  assign po6723 = pi6742;
  assign po6724 = pi6726;
  assign po6725 = pi6763;
  assign po6726 = pi6747;
  assign po6727 = pi6725;
  assign po6728 = pi6774;
  assign po6729 = pi6766;
  assign po6730 = pi6734;
  assign po6731 = pi6727;
  assign po6732 = pi6722;
  assign po6733 = pi6736;
  assign po6734 = pi6731;
  assign po6735 = pi6769;
  assign po6736 = pi6765;
  assign po6737 = pi6730;
  assign po6738 = pi6735;
  assign po6739 = pi6772;
  assign po6740 = pi6760;
  assign po6741 = pi6741;
  assign po6742 = pi6768;
  assign po6743 = pi6750;
  assign po6744 = pi6738;
  assign po6745 = pi6761;
  assign po6746 = pi6723;
  assign po6747 = pi6751;
  assign po6748 = pi6757;
  assign po6749 = pi6743;
  assign po6750 = pi6777;
  assign po6751 = pi6759;
  assign po6752 = pi6717;
  assign po6753 = pi6720;
  assign po6754 = pi6715;
  assign po6755 = pi6764;
  assign po6756 = pi6753;
  assign po6757 = pi6773;
  assign po6758 = pi6754;
  assign po6759 = pi6728;
  assign po6760 = pi6744;
  assign po6761 = pi6718;
  assign po6762 = pi6733;
  assign po6763 = pi6729;
  assign po6764 = pi6748;
  assign po6765 = pi6622;
  assign po6766 = pi6775;
  assign po6767 = pi6745;
  assign po6768 = pi6624;
  assign po6769 = pi6752;
  assign po6770 = pi6762;
  assign po6771 = pi6737;
  assign po6772 = pi6732;
  assign po6773 = pi6767;
  assign po6774 = pi6719;
  assign po6775 = pi6712;
  assign po6776 = pi6746;
  assign po6777 = pi6665;
  assign po6778 = pi6646;
  assign po6779 = pi6701;
  assign po6780 = pi6630;
  assign po6781 = pi6799;
  assign po6782 = pi6644;
  assign po6783 = pi6645;
  assign po6784 = pi6685;
  assign po6785 = pi6828;
  assign po6786 = pi6642;
  assign po6787 = pi6683;
  assign po6788 = pi6703;
  assign po6789 = pi6638;
  assign po6790 = pi6709;
  assign po6791 = pi6631;
  assign po6792 = pi6639;
  assign po6793 = pi6678;
  assign po6794 = pi6710;
  assign po6795 = pi6682;
  assign po6796 = pi6649;
  assign po6797 = pi6675;
  assign po6798 = pi6653;
  assign po6799 = pi6689;
  assign po6800 = pi6635;
  assign po6801 = pi6659;
  assign po6802 = pi6711;
  assign po6803 = pi6657;
  assign po6804 = pi6686;
  assign po6805 = pi6690;
  assign po6806 = pi6666;
  assign po6807 = pi6739;
  assign po6808 = pi6677;
  assign po6809 = pi6643;
  assign po6810 = pi6704;
  assign po6811 = pi6688;
  assign po6812 = pi6652;
  assign po6813 = pi6708;
  assign po6814 = pi6696;
  assign po6815 = pi6636;
  assign po6816 = pi6700;
  assign po6817 = pi6647;
  assign po6818 = pi6692;
  assign po6819 = pi6650;
  assign po6820 = pi6633;
  assign po6821 = pi6640;
  assign po6822 = pi6654;
  assign po6823 = pi6641;
  assign po6824 = pi6656;
  assign po6825 = pi6651;
  assign po6826 = pi6714;
  assign po6827 = pi6648;
  assign po6828 = pi6794;
  assign po6829 = pi6839;
  assign po6830 = pi6778;
  assign po6831 = pi6694;
  assign po6832 = pi6809;
  assign po6833 = pi6721;
  assign po6834 = pi6801;
  assign po6835 = pi6782;
  assign po6836 = pi6780;
  assign po6837 = pi6827;
  assign po6838 = pi6756;
  assign po6839 = pi6821;
  assign po6840 = pi6800;
  assign po6841 = pi6691;
  assign po6842 = pi6702;
  assign po6843 = pi6806;
  assign po6844 = pi6697;
  assign po6845 = pi6679;
  assign po6846 = pi6705;
  assign po6847 = pi6713;
  assign po6848 = pi6687;
  assign po6849 = pi6706;
  assign po6850 = pi6716;
  assign po6851 = pi6849;
  assign po6852 = pi6857;
  assign po6853 = pi6859;
  assign po6854 = pi6853;
  assign po6855 = pi6855;
  assign po6856 = pi6770;
  assign po6857 = pi6740;
  assign po6858 = pi6776;
  assign po6859 = pi6858;
  assign po6860 = pi6796;
  assign po6861 = pi6824;
  assign po6862 = pi6885;
  assign po6863 = pi6825;
  assign po6864 = pi6897;
  assign po6865 = pi6836;
  assign po6866 = pi6803;
  assign po6867 = pi6811;
  assign po6868 = pi6851;
  assign po6869 = pi6843;
  assign po6870 = pi6787;
  assign po6871 = pi6841;
  assign po6872 = pi6840;
  assign po6873 = pi6845;
  assign po6874 = pi6837;
  assign po6875 = pi6805;
  assign po6876 = pi6829;
  assign po6877 = pi6790;
  assign po6878 = pi6833;
  assign po6879 = pi6784;
  assign po6880 = pi6808;
  assign po6881 = pi6817;
  assign po6882 = pi6842;
  assign po6883 = pi6831;
  assign po6884 = pi6783;
  assign po6885 = pi6864;
  assign po6886 = pi6846;
  assign po6887 = pi6810;
  assign po6888 = pi6937;
  assign po6889 = pi6834;
  assign po6890 = pi6884;
  assign po6891 = pi6861;
  assign po6892 = pi6922;
  assign po6893 = pi6870;
  assign po6894 = pi6917;
  assign po6895 = pi6785;
  assign po6896 = pi6802;
  assign po6897 = pi6905;
  assign po6898 = pi6874;
  assign po6899 = pi6895;
  assign po6900 = pi6913;
  assign po6901 = pi6860;
  assign po6902 = pi6879;
  assign po6903 = pi6911;
  assign po6904 = pi6867;
  assign po6905 = pi6820;
  assign po6906 = pi6936;
  assign po6907 = pi6812;
  assign po6908 = pi6789;
  assign po6909 = pi6832;
  assign po6910 = pi6807;
  assign po6911 = pi6844;
  assign po6912 = pi6822;
  assign po6913 = pi6835;
  assign po6914 = pi6909;
  assign po6915 = pi6848;
  assign po6916 = pi6826;
  assign po6917 = pi6823;
  assign po6918 = pi6795;
  assign po6919 = pi6793;
  assign po6920 = pi6797;
  assign po6921 = pi6818;
  assign po6922 = pi6838;
  assign po6923 = pi6941;
  assign po6924 = pi6781;
  assign po6925 = pi6854;
  assign po6926 = pi6788;
  assign po6927 = pi6878;
  assign po6928 = pi6896;
  assign po6929 = pi6889;
  assign po6930 = pi6816;
  assign po6931 = pi6791;
  assign po6932 = pi6847;
  assign po6933 = pi6792;
  assign po6934 = pi6804;
  assign po6935 = pi6815;
  assign po6936 = pi6915;
  assign po6937 = pi6866;
  assign po6938 = pi6798;
  assign po6939 = pi6830;
  assign po6940 = pi6850;
  assign po6941 = pi6786;
  assign po6942 = pi6814;
  assign po6943 = pi6813;
  assign po6944 = pi6819;
  assign po6945 = pi6947;
  assign po6946 = pi6972;
  assign po6947 = pi6962;
  assign po6948 = pi6852;
  assign po6949 = pi6993;
  assign po6950 = pi6961;
  assign po6951 = pi7010;
  assign po6952 = pi6977;
  assign po6953 = pi6945;
  assign po6954 = pi6992;
  assign po6955 = pi6975;
  assign po6956 = pi6999;
  assign po6957 = pi6963;
  assign po6958 = pi6965;
  assign po6959 = pi6856;
  assign po6960 = pi7000;
  assign po6961 = pi6998;
  assign po6962 = pi6927;
  assign po6963 = pi6980;
  assign po6964 = pi6872;
  assign po6965 = pi6971;
  assign po6966 = pi6964;
  assign po6967 = pi7013;
  assign po6969 = pi6989;
  assign po6970 = pi7011;
  assign po6971 = pi6957;
  assign po6972 = pi6955;
  assign po6973 = pi6969;
  assign po6974 = pi6973;
  assign po6975 = pi6987;
  assign po6976 = pi6994;
  assign po6977 = pi6950;
  assign po6978 = pi6948;
  assign po6979 = pi6968;
  assign po6980 = pi6986;
  assign po6981 = pi7012;
  assign po6982 = pi6981;
  assign po6983 = pi6956;
  assign po6984 = pi6983;
  assign po6985 = pi6952;
  assign po6986 = pi6967;
  assign po6987 = pi6979;
  assign po6988 = pi6959;
  assign po6989 = pi7003;
  assign po6990 = pi7008;
  assign po6991 = pi6988;
  assign po6992 = pi7009;
  assign po6993 = pi6991;
  assign po6994 = pi7004;
  assign po6995 = pi6997;
  assign po6996 = pi6970;
  assign po6997 = pi6958;
  assign po6998 = pi6974;
  assign po7000 = pi6966;
  assign po7001 = pi6985;
  assign po7002 = pi6951;
  assign po7003 = pi7005;
  assign po7004 = pi6995;
  assign po7005 = pi7002;
  assign po7006 = pi6953;
  assign po7007 = pi7006;
  assign po7008 = pi6984;
  assign po7009 = pi6946;
  assign po7010 = pi7068;
  assign po7011 = pi6890;
  assign po7012 = pi6954;
  assign po7013 = pi6914;
  assign po7014 = pi6907;
  assign po7015 = pi6934;
  assign po7016 = pi6883;
  assign po7017 = pi6899;
  assign po7018 = pi6880;
  assign po7019 = pi6865;
  assign po7020 = pi6876;
  assign po7021 = pi6904;
  assign po7022 = pi6881;
  assign po7023 = pi6877;
  assign po7024 = pi7048;
  assign po7025 = pi6921;
  assign po7026 = pi6929;
  assign po7027 = pi6933;
  assign po7028 = pi6925;
  assign po7029 = pi7001;
  assign po7030 = pi7020;
  assign po7031 = pi7063;
  assign po7032 = pi6930;
  assign po7033 = pi6894;
  assign po7034 = pi6875;
  assign po7035 = pi6892;
  assign po7036 = pi7016;
  assign po7037 = pi7073;
  assign po7038 = pi6887;
  assign po7039 = pi7022;
  assign po7040 = pi6943;
  assign po7041 = pi7028;
  assign po7042 = pi6903;
  assign po7043 = pi6900;
  assign po7044 = pi6901;
  assign po7045 = pi6908;
  assign po7046 = pi6873;
  assign po7047 = pi6863;
  assign po7048 = pi6902;
  assign po7049 = pi6926;
  assign po7050 = pi6923;
  assign po7051 = pi6982;
  assign po7052 = pi6871;
  assign po7053 = pi6893;
  assign po7054 = pi6935;
  assign po7055 = pi6916;
  assign po7056 = pi6924;
  assign po7057 = pi6960;
  assign po7058 = pi7080;
  assign po7059 = pi6862;
  assign po7060 = pi6939;
  assign po7061 = pi6919;
  assign po7062 = pi6940;
  assign po7063 = pi6932;
  assign po7064 = pi6931;
  assign po7065 = pi6891;
  assign po7066 = pi6886;
  assign po7067 = pi6928;
  assign po7068 = pi6898;
  assign po7069 = pi7018;
  assign po7070 = pi6869;
  assign po7071 = pi6944;
  assign po7072 = pi6938;
  assign po7073 = pi6912;
  assign po7074 = pi7025;
  assign po7075 = pi6942;
  assign po7076 = pi6910;
  assign po7077 = pi6906;
  assign po7078 = pi6888;
  assign po7079 = pi6990;
  assign po7080 = pi6920;
  assign po7081 = pi6882;
  assign po7082 = pi7081;
  assign po7083 = pi6976;
  assign po7084 = pi7007;
  assign po7085 = pi7083;
  assign po7086 = pi7082;
  assign po7087 = pi6949;
  assign po7088 = pi6978;
  assign po7089 = pi6996;
  assign po7090 = pi7159;
  assign po7091 = pi7169;
  assign po7092 = pi7036;
  assign po7093 = pi7069;
  assign po7094 = pi7154;
  assign po7095 = pi7053;
  assign po7096 = pi7134;
  assign po7097 = pi7151;
  assign po7098 = pi7177;
  assign po7099 = pi7064;
  assign po7100 = pi7143;
  assign po7101 = pi7062;
  assign po7102 = pi7142;
  assign po7103 = pi7021;
  assign po7104 = pi7146;
  assign po7105 = pi7035;
  assign po7106 = pi7029;
  assign po7107 = pi7051;
  assign po7108 = pi7153;
  assign po7109 = pi7117;
  assign po7110 = pi7067;
  assign po7111 = pi7078;
  assign po7112 = pi7077;
  assign po7113 = pi7060;
  assign po7114 = pi7161;
  assign po7115 = pi7166;
  assign po7116 = pi7027;
  assign po7117 = pi7026;
  assign po7118 = pi7047;
  assign po7119 = pi7101;
  assign po7120 = pi7043;
  assign po7121 = pi7033;
  assign po7122 = pi7076;
  assign po7123 = pi7071;
  assign po7124 = pi7059;
  assign po7125 = pi7158;
  assign po7126 = pi7167;
  assign po7127 = pi7162;
  assign po7128 = pi7037;
  assign po7129 = pi7057;
  assign po7130 = pi7058;
  assign po7131 = pi7045;
  assign po7132 = pi7039;
  assign po7133 = pi7044;
  assign po7134 = pi7038;
  assign po7135 = pi7140;
  assign po7136 = pi7015;
  assign po7137 = pi7041;
  assign po7138 = pi7055;
  assign po7139 = pi7144;
  assign po7140 = pi7074;
  assign po7141 = pi7145;
  assign po7142 = pi7024;
  assign po7143 = pi7165;
  assign po7144 = pi7040;
  assign po7145 = pi7148;
  assign po7146 = pi7046;
  assign po7147 = pi7160;
  assign po7148 = pi7157;
  assign po7149 = pi7052;
  assign po7150 = pi7017;
  assign po7151 = pi7023;
  assign po7152 = pi7141;
  assign po7153 = pi7049;
  assign po7154 = pi7070;
  assign po7155 = pi7056;
  assign po7156 = pi7075;
  assign po7157 = pi7135;
  assign po7158 = pi7032;
  assign po7159 = pi7019;
  assign po7160 = pi7066;
  assign po7161 = pi7050;
  assign po7162 = pi7034;
  assign po7163 = pi7014;
  assign po7164 = pi7031;
  assign po7165 = pi7079;
  assign po7166 = pi7137;
  assign po7167 = pi7147;
  assign po7168 = pi7065;
  assign po7169 = pi7054;
  assign po7170 = pi7072;
  assign po7171 = pi7084;
  assign po7172 = pi7030;
  assign po7173 = pi7042;
  assign po7174 = pi7061;
  assign po7175 = pi7191;
  assign po7176 = pi7220;
  assign po7177 = pi7183;
  assign po7178 = pi7219;
  assign po7179 = pi7181;
  assign po7180 = pi7217;
  assign po7181 = pi7199;
  assign po7182 = pi7245;
  assign po7183 = pi7195;
  assign po7184 = pi7187;
  assign po7185 = pi7182;
  assign po7186 = pi7241;
  assign po7187 = pi7188;
  assign po7188 = pi7223;
  assign po7189 = pi7197;
  assign po7190 = pi7202;
  assign po7191 = pi7192;
  assign po7192 = pi7226;
  assign po7193 = pi7118;
  assign po7194 = pi7230;
  assign po7195 = pi7205;
  assign po7196 = pi7216;
  assign po7197 = pi7208;
  assign po7198 = pi7238;
  assign po7199 = pi7221;
  assign po7200 = pi7231;
  assign po7201 = pi7218;
  assign po7202 = pi7198;
  assign po7203 = pi7184;
  assign po7204 = pi7215;
  assign po7205 = pi7225;
  assign po7206 = pi7235;
  assign po7207 = pi7228;
  assign po7208 = pi7190;
  assign po7209 = pi7196;
  assign po7210 = pi7201;
  assign po7211 = pi7180;
  assign po7212 = pi7185;
  assign po7213 = pi7200;
  assign po7214 = pi7239;
  assign po7215 = pi7207;
  assign po7216 = pi7242;
  assign po7217 = pi7098;
  assign po7218 = pi7186;
  assign po7219 = pi7164;
  assign po7220 = pi7212;
  assign po7221 = pi7138;
  assign po7222 = pi7189;
  assign po7223 = pi7206;
  assign po7224 = pi7243;
  assign po7225 = pi7155;
  assign po7226 = pi7203;
  assign po7227 = pi7229;
  assign po7228 = pi7234;
  assign po7229 = pi7150;
  assign po7230 = pi7233;
  assign po7231 = pi7236;
  assign po7232 = pi7209;
  assign po7233 = pi7213;
  assign po7234 = pi7204;
  assign po7235 = pi7244;
  assign po7236 = pi7214;
  assign po7237 = pi7237;
  assign po7238 = pi7193;
  assign po7239 = pi7240;
  assign po7240 = pi7224;
  assign po7241 = pi7136;
  assign po7242 = pi7227;
  assign po7243 = pi7156;
  assign po7244 = pi7114;
  assign po7245 = pi7102;
  assign po7246 = pi7285;
  assign po7247 = pi7172;
  assign po7248 = pi7248;
  assign po7249 = pi7116;
  assign po7250 = pi7294;
  assign po7251 = pi7092;
  assign po7252 = pi7292;
  assign po7253 = pi7091;
  assign po7254 = pi7100;
  assign po7255 = pi7272;
  assign po7256 = pi7123;
  assign po7257 = pi7128;
  assign po7258 = pi7232;
  assign po7259 = pi7108;
  assign po7260 = pi7111;
  assign po7261 = pi7095;
  assign po7262 = pi7124;
  assign po7263 = pi7103;
  assign po7264 = pi7132;
  assign po7265 = pi7130;
  assign po7266 = pi7133;
  assign po7267 = pi7119;
  assign po7268 = pi7149;
  assign po7269 = pi7121;
  assign po7270 = pi7086;
  assign po7271 = pi7131;
  assign po7272 = pi7173;
  assign po7273 = pi7104;
  assign po7274 = pi7112;
  assign po7275 = pi7109;
  assign po7276 = pi7129;
  assign po7277 = pi7097;
  assign po7278 = pi7250;
  assign po7279 = pi7093;
  assign po7280 = pi7125;
  assign po7281 = pi7105;
  assign po7282 = pi7115;
  assign po7283 = pi7176;
  assign po7284 = pi7122;
  assign po7285 = pi7152;
  assign po7286 = pi7087;
  assign po7287 = pi7106;
  assign po7288 = pi7168;
  assign po7289 = pi7178;
  assign po7290 = pi7096;
  assign po7291 = pi7171;
  assign po7292 = pi7120;
  assign po7293 = pi7246;
  assign po7294 = pi7175;
  assign po7295 = pi7099;
  assign po7296 = pi7126;
  assign po7297 = pi7110;
  assign po7298 = pi7210;
  assign po7299 = pi7127;
  assign po7300 = pi7113;
  assign po7301 = pi7089;
  assign po7302 = pi7090;
  assign po7303 = pi7085;
  assign po7304 = pi7094;
  assign po7305 = pi7139;
  assign po7306 = pi7170;
  assign po7307 = pi7088;
  assign po7308 = pi7107;
  assign po7309 = pi7174;
  assign po7310 = pi7163;
  assign po7311 = pi7194;
  assign po7312 = pi7211;
  assign po7313 = pi7222;
  assign po7314 = pi7179;
  assign po7315 = pi7446;
  assign po7316 = pi7302;
  assign po7317 = pi7282;
  assign po7318 = pi7257;
  assign po7319 = pi7270;
  assign po7320 = pi7264;
  assign po7321 = pi7283;
  assign po7322 = pi7273;
  assign po7323 = pi7253;
  assign po7324 = pi7309;
  assign po7325 = pi7254;
  assign po7326 = pi7296;
  assign po7327 = pi7306;
  assign po7328 = pi7423;
  assign po7329 = pi7262;
  assign po7330 = pi7256;
  assign po7331 = pi7369;
  assign po7332 = pi7276;
  assign po7333 = pi7281;
  assign po7334 = pi7298;
  assign po7335 = pi7265;
  assign po7336 = pi7288;
  assign po7337 = pi7252;
  assign po7338 = pi7304;
  assign po7339 = pi7301;
  assign po7340 = pi7263;
  assign po7341 = pi7277;
  assign po7342 = pi7279;
  assign po7343 = pi7287;
  assign po7344 = pi7286;
  assign po7345 = pi7259;
  assign po7346 = pi7261;
  assign po7347 = pi7461;
  assign po7348 = pi7422;
  assign po7349 = pi7268;
  assign po7350 = pi7271;
  assign po7351 = pi7305;
  assign po7352 = pi7249;
  assign po7353 = pi7295;
  assign po7354 = pi7308;
  assign po7355 = pi7300;
  assign po7356 = pi7266;
  assign po7357 = pi7255;
  assign po7358 = pi7307;
  assign po7359 = pi7303;
  assign po7360 = pi7290;
  assign po7361 = pi7274;
  assign po7362 = pi7297;
  assign po7363 = pi7251;
  assign po7364 = pi7293;
  assign po7365 = pi7462;
  assign po7366 = pi7409;
  assign po7367 = pi7444;
  assign po7368 = pi7436;
  assign po7369 = pi7278;
  assign po7370 = pi7366;
  assign po7371 = pi7429;
  assign po7372 = pi7383;
  assign po7373 = pi7411;
  assign po7374 = pi7433;
  assign po7375 = pi7414;
  assign po7376 = pi7424;
  assign po7377 = pi7415;
  assign po7378 = pi7386;
  assign po7379 = pi7299;
  assign po7380 = pi7454;
  assign po7381 = pi7428;
  assign po7382 = pi7280;
  assign po7383 = pi7453;
  assign po7384 = pi7413;
  assign po7385 = pi7421;
  assign po7386 = pi7376;
  assign po7387 = pi7456;
  assign po7388 = pi7385;
  assign po7389 = pi7410;
  assign po7390 = pi7460;
  assign po7391 = pi7450;
  assign po7392 = pi7434;
  assign po7393 = pi7425;
  assign po7394 = pi7417;
  assign po7395 = pi7412;
  assign po7396 = pi7440;
  assign po7397 = pi7426;
  assign po7398 = pi7275;
  assign po7399 = pi7379;
  assign po7400 = pi7284;
  assign po7401 = pi7269;
  assign po7402 = pi7291;
  assign po7403 = pi7258;
  assign po7404 = pi7267;
  assign po7405 = pi7247;
  assign po7406 = pi7289;
  assign po7407 = pi7431;
  assign po7408 = pi7260;
  assign po7409 = pi7335;
  assign po7410 = pi7314;
  assign po7411 = pi7315;
  assign po7412 = pi7359;
  assign po7413 = pi7320;
  assign po7414 = pi7348;
  assign po7415 = pi7322;
  assign po7416 = pi7352;
  assign po7417 = pi7344;
  assign po7418 = pi7331;
  assign po7419 = pi7360;
  assign po7420 = pi7321;
  assign po7421 = pi7333;
  assign po7422 = pi7327;
  assign po7423 = pi7310;
  assign po7424 = pi7356;
  assign po7425 = pi7345;
  assign po7426 = pi7353;
  assign po7427 = pi7343;
  assign po7428 = pi7355;
  assign po7429 = pi7324;
  assign po7430 = pi7357;
  assign po7431 = pi7358;
  assign po7432 = pi7346;
  assign po7433 = pi7329;
  assign po7434 = pi7364;
  assign po7435 = pi7330;
  assign po7436 = pi7350;
  assign po7437 = pi7319;
  assign po7438 = pi7365;
  assign po7439 = pi7341;
  assign po7440 = pi7334;
  assign po7441 = pi7323;
  assign po7442 = pi7311;
  assign po7443 = pi7318;
  assign po7444 = pi7325;
  assign po7445 = pi7354;
  assign po7446 = pi7338;
  assign po7447 = pi7332;
  assign po7448 = pi7466;
  assign po7449 = pi7351;
  assign po7450 = pi7361;
  assign po7451 = pi7339;
  assign po7452 = pi7313;
  assign po7453 = pi7347;
  assign po7454 = pi7401;
  assign po7455 = pi7312;
  assign po7456 = pi7340;
  assign po7457 = pi7349;
  assign po7458 = pi7439;
  assign po7459 = pi7511;
  assign po7460 = pi7519;
  assign po7461 = pi7522;
  assign po7462 = pi7518;
  assign po7463 = pi7397;
  assign po7464 = pi7430;
  assign po7465 = pi7396;
  assign po7466 = pi7521;
  assign po7467 = pi7362;
  assign po7468 = pi7328;
  assign po7469 = pi7317;
  assign po7470 = pi7336;
  assign po7471 = pi7337;
  assign po7472 = pi7363;
  assign po7473 = pi7342;
  assign po7474 = pi7316;
  assign po7475 = pi7326;
  assign po7476 = pi7449;
  assign po7477 = pi7464;
  assign po7478 = pi7534;
  assign po7479 = pi7458;
  assign po7480 = pi7568;
  assign po7481 = pi7371;
  assign po7482 = pi7420;
  assign po7483 = pi7442;
  assign po7484 = pi7387;
  assign po7485 = pi7378;
  assign po7486 = pi7402;
  assign po7487 = pi7381;
  assign po7488 = pi7432;
  assign po7489 = pi7373;
  assign po7490 = pi7405;
  assign po7491 = pi7380;
  assign po7492 = pi7451;
  assign po7493 = pi7445;
  assign po7494 = pi7400;
  assign po7495 = pi7367;
  assign po7496 = pi7465;
  assign po7497 = pi7416;
  assign po7498 = pi7399;
  assign po7499 = pi7394;
  assign po7500 = pi7403;
  assign po7501 = pi7408;
  assign po7502 = pi7591;
  assign po7503 = pi7435;
  assign po7504 = pi7459;
  assign po7505 = pi7447;
  assign po7506 = pi7384;
  assign po7507 = pi7407;
  assign po7508 = pi7418;
  assign po7509 = pi7463;
  assign po7510 = pi7452;
  assign po7511 = pi7437;
  assign po7512 = pi7375;
  assign po7513 = pi7393;
  assign po7514 = pi7374;
  assign po7515 = pi7427;
  assign po7516 = pi7448;
  assign po7517 = pi7398;
  assign po7518 = pi7392;
  assign po7519 = pi7370;
  assign po7520 = pi7406;
  assign po7521 = pi7441;
  assign po7522 = pi7528;
  assign po7523 = pi7537;
  assign po7524 = pi7589;
  assign po7525 = pi7438;
  assign po7526 = pi7368;
  assign po7527 = pi7391;
  assign po7528 = pi7455;
  assign po7529 = pi7377;
  assign po7530 = pi7389;
  assign po7531 = pi7457;
  assign po7532 = pi7372;
  assign po7533 = pi7404;
  assign po7534 = pi7419;
  assign po7535 = pi7443;
  assign po7536 = pi7390;
  assign po7537 = pi7395;
  assign po7538 = pi7382;
  assign po7539 = pi7388;
  assign po7540 = pi7483;
  assign po7541 = pi7474;
  assign po7542 = pi7494;
  assign po7543 = pi7503;
  assign po7544 = pi7477;
  assign po7545 = pi7491;
  assign po7546 = pi7497;
  assign po7547 = pi7488;
  assign po7548 = pi7485;
  assign po7549 = pi7484;
  assign po7550 = pi7499;
  assign po7551 = pi7512;
  assign po7552 = pi7473;
  assign po7553 = pi7505;
  assign po7554 = pi7510;
  assign po7555 = pi7527;
  assign po7556 = pi7487;
  assign po7557 = pi7472;
  assign po7558 = pi7516;
  assign po7559 = pi7482;
  assign po7560 = pi7506;
  assign po7561 = pi7523;
  assign po7562 = pi7524;
  assign po7563 = pi7480;
  assign po7564 = pi7514;
  assign po7565 = pi7504;
  assign po7566 = pi7515;
  assign po7567 = pi7517;
  assign po7568 = pi7508;
  assign po7569 = pi7509;
  assign po7570 = pi7513;
  assign po7571 = pi7493;
  assign po7572 = pi7489;
  assign po7573 = pi7475;
  assign po7574 = pi7476;
  assign po7575 = pi7486;
  assign po7576 = pi7525;
  assign po7577 = pi7496;
  assign po7578 = pi7469;
  assign po7579 = pi7490;
  assign po7580 = pi7471;
  assign po7581 = pi7502;
  assign po7582 = pi7526;
  assign po7583 = pi7467;
  assign po7584 = pi7479;
  assign po7585 = pi7495;
  assign po7586 = pi7520;
  assign po7587 = pi7498;
  assign po7588 = pi7492;
  assign po7589 = pi7468;
  assign po7590 = pi7478;
  assign po7591 = pi7501;
  assign po7592 = pi7507;
  assign po7593 = pi7470;
  assign po7594 = pi7500;
  assign po7595 = pi7481;
  assign po7596 = pi7703;
  assign po7597 = pi7555;
  assign po7598 = pi7587;
  assign po7599 = pi7726;
  assign po7600 = pi7570;
  assign po7601 = pi7564;
  assign po7602 = pi7531;
  assign po7603 = pi7574;
  assign po7604 = pi7580;
  assign po7605 = pi7538;
  assign po7606 = pi7744;
  assign po7607 = pi7560;
  assign po7608 = pi7562;
  assign po7609 = pi7674;
  assign po7610 = pi7541;
  assign po7611 = pi7585;
  assign po7612 = pi7563;
  assign po7613 = pi7711;
  assign po7614 = pi7586;
  assign po7615 = pi7660;
  assign po7616 = pi7745;
  assign po7617 = pi7567;
  assign po7618 = pi7552;
  assign po7619 = pi7532;
  assign po7620 = pi7583;
  assign po7621 = pi7565;
  assign po7622 = pi7536;
  assign po7623 = pi7543;
  assign po7624 = pi7561;
  assign po7625 = pi7571;
  assign po7626 = pi7649;
  assign po7627 = pi7684;
  assign po7628 = pi7550;
  assign po7629 = pi7549;
  assign po7630 = pi7533;
  assign po7631 = pi7661;
  assign po7632 = pi7529;
  assign po7633 = pi7539;
  assign po7634 = pi7548;
  assign po7635 = pi7578;
  assign po7636 = pi7559;
  assign po7637 = pi7545;
  assign po7638 = pi7572;
  assign po7639 = pi7736;
  assign po7640 = pi7727;
  assign po7641 = pi7648;
  assign po7642 = pi7659;
  assign po7643 = pi7693;
  assign po7644 = pi7651;
  assign po7645 = pi7668;
  assign po7646 = pi7557;
  assign po7647 = pi7663;
  assign po7648 = pi7546;
  assign po7649 = pi7576;
  assign po7650 = pi7553;
  assign po7651 = pi7683;
  assign po7652 = pi7741;
  assign po7653 = pi7590;
  assign po7654 = pi7725;
  assign po7655 = pi7670;
  assign po7656 = pi7575;
  assign po7657 = pi7653;
  assign po7658 = pi7742;
  assign po7659 = pi7658;
  assign po7660 = pi7708;
  assign po7661 = pi7739;
  assign po7662 = pi7573;
  assign po7663 = pi7664;
  assign po7664 = pi7733;
  assign po7665 = pi7558;
  assign po7666 = pi7705;
  assign po7667 = pi7584;
  assign po7668 = pi7566;
  assign po7669 = pi7689;
  assign po7670 = pi7677;
  assign po7671 = pi7588;
  assign po7672 = pi7542;
  assign po7673 = pi7530;
  assign po7674 = pi7662;
  assign po7675 = pi7581;
  assign po7676 = pi7752;
  assign po7677 = pi7544;
  assign po7678 = pi7554;
  assign po7679 = pi7749;
  assign po7680 = pi7666;
  assign po7681 = pi7577;
  assign po7682 = pi7569;
  assign po7683 = pi7679;
  assign po7684 = pi7655;
  assign po7685 = pi7582;
  assign po7686 = pi7721;
  assign po7687 = pi7551;
  assign po7688 = pi7556;
  assign po7689 = pi7547;
  assign po7690 = pi7698;
  assign po7691 = pi7720;
  assign po7692 = pi7675;
  assign po7693 = pi7540;
  assign po7694 = pi7579;
  assign po7695 = pi7535;
  assign po7696 = pi7723;
  assign po7697 = pi7634;
  assign po7698 = pi7641;
  assign po7699 = pi7621;
  assign po7700 = pi7626;
  assign po7701 = pi7645;
  assign po7702 = pi7612;
  assign po7703 = pi7624;
  assign po7704 = pi7604;
  assign po7705 = pi7628;
  assign po7706 = pi7616;
  assign po7707 = pi7630;
  assign po7708 = pi7618;
  assign po7709 = pi7633;
  assign po7710 = pi7622;
  assign po7711 = pi7640;
  assign po7712 = pi7639;
  assign po7713 = pi7593;
  assign po7714 = pi7637;
  assign po7715 = pi7625;
  assign po7716 = pi7614;
  assign po7717 = pi7608;
  assign po7718 = pi7603;
  assign po7719 = pi7598;
  assign po7720 = pi7623;
  assign po7721 = pi7611;
  assign po7722 = pi7596;
  assign po7723 = pi7642;
  assign po7724 = pi7617;
  assign po7725 = pi7632;
  assign po7726 = pi7595;
  assign po7727 = pi7619;
  assign po7728 = pi7631;
  assign po7729 = pi7635;
  assign po7730 = pi7610;
  assign po7731 = pi7600;
  assign po7732 = pi7605;
  assign po7733 = pi7644;
  assign po7734 = pi7606;
  assign po7735 = pi7599;
  assign po7736 = pi7602;
  assign po7737 = pi7646;
  assign po7738 = pi7620;
  assign po7739 = pi7592;
  assign po7740 = pi7597;
  assign po7741 = pi7686;
  assign po7742 = pi7615;
  assign po7743 = pi7607;
  assign po7744 = pi7601;
  assign po7745 = pi7594;
  assign po7746 = pi7627;
  assign po7747 = pi7647;
  assign po7748 = pi7795;
  assign po7749 = pi7811;
  assign po7750 = pi7643;
  assign po7751 = pi7803;
  assign po7752 = pi7700;
  assign po7753 = pi7609;
  assign po7754 = pi7629;
  assign po7755 = pi7636;
  assign po7756 = pi7613;
  assign po7757 = pi7638;
  assign po7758 = pi7746;
  assign po7759 = pi7738;
  assign po7760 = pi7713;
  assign po7761 = pi7716;
  assign po7762 = pi7718;
  assign po7763 = pi7737;
  assign po7764 = pi7750;
  assign po7765 = pi7728;
  assign po7766 = pi7687;
  assign po7767 = pi7652;
  assign po7768 = pi7696;
  assign po7769 = pi7680;
  assign po7770 = pi7730;
  assign po7771 = pi7732;
  assign po7772 = pi7747;
  assign po7773 = pi7734;
  assign po7774 = pi7702;
  assign po7775 = pi7715;
  assign po7776 = pi7722;
  assign po7777 = pi7740;
  assign po7778 = pi7719;
  assign po7779 = pi7731;
  assign po7780 = pi7673;
  assign po7781 = pi7690;
  assign po7782 = pi7717;
  assign po7783 = pi7714;
  assign po7784 = pi7712;
  assign po7785 = pi7697;
  assign po7786 = pi7706;
  assign po7787 = pi7704;
  assign po7788 = pi7656;
  assign po7789 = pi7709;
  assign po7790 = pi7751;
  assign po7791 = pi7665;
  assign po7792 = pi7724;
  assign po7793 = pi7688;
  assign po7794 = pi7748;
  assign po7795 = pi7654;
  assign po7796 = pi7710;
  assign po7797 = pi7676;
  assign po7798 = pi7821;
  assign po7799 = pi7692;
  assign po7800 = pi7671;
  assign po7801 = pi7743;
  assign po7802 = pi7699;
  assign po7803 = pi7694;
  assign po7804 = pi7707;
  assign po7805 = pi7817;
  assign po7806 = pi7735;
  assign po7807 = pi7685;
  assign po7808 = pi7667;
  assign po7809 = pi7657;
  assign po7810 = pi7695;
  assign po7811 = pi7701;
  assign po7812 = pi7678;
  assign po7813 = pi7682;
  assign po7814 = pi7691;
  assign po7815 = pi7672;
  assign po7816 = pi7669;
  assign po7817 = pi7729;
  assign po7818 = pi7681;
  assign po7819 = pi7813;
  assign po7820 = pi7846;
  assign po7821 = pi7650;
  assign po7822 = pi7754;
  assign po7823 = pi7809;
  assign po7824 = pi7789;
  assign po7825 = pi7775;
  assign po7826 = pi7800;
  assign po7827 = pi7797;
  assign po7828 = pi7801;
  assign po7829 = pi7804;
  assign po7830 = pi7762;
  assign po7831 = pi7776;
  assign po7832 = pi7759;
  assign po7833 = pi7771;
  assign po7834 = pi7757;
  assign po7835 = pi7792;
  assign po7836 = pi7779;
  assign po7837 = pi7778;
  assign po7838 = pi7772;
  assign po7839 = pi7769;
  assign po7840 = pi7791;
  assign po7841 = pi7785;
  assign po7842 = pi7798;
  assign po7843 = pi7794;
  assign po7844 = pi7773;
  assign po7845 = pi7787;
  assign po7846 = pi7783;
  assign po7847 = pi7755;
  assign po7848 = pi7766;
  assign po7849 = pi7781;
  assign po7850 = pi7796;
  assign po7851 = pi7782;
  assign po7852 = pi7780;
  assign po7853 = pi7802;
  assign po7854 = pi7799;
  assign po7855 = pi7761;
  assign po7856 = pi7786;
  assign po7857 = pi7764;
  assign po7858 = pi7784;
  assign po7859 = pi7777;
  assign po7860 = pi7760;
  assign po7861 = pi7810;
  assign po7862 = pi7808;
  assign po7863 = pi7758;
  assign po7864 = pi7793;
  assign po7865 = pi7770;
  assign po7866 = pi7805;
  assign po7867 = pi7774;
  assign po7868 = pi7768;
  assign po7869 = pi7788;
  assign po7870 = pi7753;
  assign po7871 = pi7756;
  assign po7872 = pi7806;
  assign po7873 = pi7807;
  assign po7874 = pi7790;
  assign po7875 = pi7767;
  assign po7876 = pi7763;
  assign po7877 = pi7765;
  assign po7878 = pi7961;
  assign po7879 = pi7998;
  assign po7880 = pi8023;
  assign po7881 = pi8005;
  assign po7882 = pi7929;
  assign po7883 = pi7940;
  assign po7884 = pi7826;
  assign po7885 = pi8001;
  assign po7886 = pi7851;
  assign po7887 = pi7868;
  assign po7888 = pi8004;
  assign po7889 = pi7991;
  assign po7890 = pi8038;
  assign po7891 = pi8020;
  assign po7892 = pi7954;
  assign po7893 = pi8017;
  assign po7894 = pi8003;
  assign po7895 = pi7869;
  assign po7896 = pi8015;
  assign po7897 = pi7838;
  assign po7898 = pi7975;
  assign po7899 = pi7849;
  assign po7900 = pi7942;
  assign po7901 = pi7866;
  assign po7902 = pi7862;
  assign po7903 = pi7854;
  assign po7904 = pi7939;
  assign po7905 = pi7999;
  assign po7906 = pi7819;
  assign po7907 = pi8036;
  assign po7908 = pi7844;
  assign po7909 = pi8033;
  assign po7910 = pi7816;
  assign po7911 = pi7864;
  assign po7912 = pi7833;
  assign po7913 = pi7971;
  assign po7914 = pi7972;
  assign po7915 = pi7814;
  assign po7916 = pi7935;
  assign po7917 = pi7870;
  assign po7918 = pi7839;
  assign po7919 = pi8030;
  assign po7920 = pi7832;
  assign po7921 = pi7858;
  assign po7922 = pi7824;
  assign po7923 = pi7968;
  assign po7924 = pi7853;
  assign po7925 = pi7836;
  assign po7926 = pi7850;
  assign po7927 = pi7848;
  assign po7928 = pi7959;
  assign po7929 = pi7837;
  assign po7930 = pi8022;
  assign po7931 = pi7820;
  assign po7932 = pi7861;
  assign po7933 = pi8016;
  assign po7934 = pi7831;
  assign po7935 = pi8025;
  assign po7936 = pi7818;
  assign po7937 = pi7842;
  assign po7938 = pi7931;
  assign po7939 = pi7815;
  assign po7940 = pi7845;
  assign po7941 = pi8011;
  assign po7942 = pi7860;
  assign po7943 = pi7863;
  assign po7944 = pi7843;
  assign po7945 = pi7827;
  assign po7946 = pi7828;
  assign po7947 = pi7867;
  assign po7948 = pi7822;
  assign po7949 = pi7865;
  assign po7950 = pi7997;
  assign po7951 = pi8000;
  assign po7952 = pi7829;
  assign po7953 = pi8034;
  assign po7954 = pi7857;
  assign po7955 = pi7965;
  assign po7956 = pi7979;
  assign po7957 = pi7946;
  assign po7958 = pi7840;
  assign po7959 = pi7841;
  assign po7960 = pi7825;
  assign po7961 = pi7852;
  assign po7962 = pi7830;
  assign po7963 = pi7974;
  assign po7964 = pi7847;
  assign po7965 = pi7855;
  assign po7966 = pi7966;
  assign po7967 = pi7856;
  assign po7968 = pi7823;
  assign po7969 = pi7957;
  assign po7970 = pi7871;
  assign po7971 = pi8031;
  assign po7972 = pi8010;
  assign po7973 = pi7812;
  assign po7974 = pi7943;
  assign po7975 = pi7978;
  assign po7976 = pi7949;
  assign po7977 = pi7834;
  assign po7978 = pi7859;
  assign po7979 = pi8028;
  assign po7980 = pi8013;
  assign po7981 = pi7835;
  assign po7982 = pi7986;
  assign po7983 = pi7894;
  assign po7984 = pi7876;
  assign po7985 = pi7874;
  assign po7986 = pi7892;
  assign po7987 = pi7882;
  assign po7988 = pi7917;
  assign po7989 = pi7907;
  assign po7990 = pi7890;
  assign po7991 = pi7872;
  assign po7992 = pi7923;
  assign po7993 = pi7902;
  assign po7994 = pi7877;
  assign po7995 = pi7916;
  assign po7996 = pi7880;
  assign po7997 = pi7881;
  assign po7998 = pi7915;
  assign po7999 = pi7900;
  assign po8000 = pi7886;
  assign po8001 = pi7908;
  assign po8002 = pi7914;
  assign po8003 = pi7899;
  assign po8004 = pi7896;
  assign po8005 = pi7924;
  assign po8006 = pi7926;
  assign po8007 = pi7879;
  assign po8008 = pi7878;
  assign po8009 = pi7912;
  assign po8010 = pi7895;
  assign po8011 = pi7904;
  assign po8012 = pi7910;
  assign po8013 = pi7898;
  assign po8014 = pi7922;
  assign po8015 = pi7887;
  assign po8016 = pi7875;
  assign po8017 = pi7903;
  assign po8018 = pi7897;
  assign po8019 = pi7893;
  assign po8020 = pi7911;
  assign po8021 = pi7883;
  assign po8022 = pi7918;
  assign po8023 = pi7906;
  assign po8024 = pi7909;
  assign po8025 = pi8039;
  assign po8026 = pi7884;
  assign po8027 = pi7901;
  assign po8028 = pi7919;
  assign po8029 = pi7873;
  assign po8030 = pi7891;
  assign po8031 = pi7905;
  assign po8032 = pi7913;
  assign po8033 = pi7952;
  assign po8034 = pi7885;
  assign po8035 = pi7888;
  assign po8036 = pi7925;
  assign po8037 = pi7921;
  assign po8038 = pi7889;
  assign po8039 = pi7927;
  assign po8040 = pi7920;
  assign po8041 = pi7963;
  assign po8042 = pi8008;
  assign po8043 = pi7937;
  assign po8044 = pi8006;
  assign po8045 = pi7984;
  assign po8046 = pi7985;
  assign po8047 = pi7977;
  assign po8048 = pi7948;
  assign po8049 = pi7969;
  assign po8050 = pi7989;
  assign po8051 = pi7958;
  assign po8052 = pi7953;
  assign po8053 = pi7973;
  assign po8054 = pi7928;
  assign po8055 = pi7987;
  assign po8056 = pi7990;
  assign po8057 = pi7947;
  assign po8058 = pi7994;
  assign po8059 = pi7951;
  assign po8060 = pi8024;
  assign po8061 = pi7992;
  assign po8062 = pi7988;
  assign po8063 = pi7933;
  assign po8064 = pi7936;
  assign po8065 = pi8027;
  assign po8066 = pi8002;
  assign po8067 = pi7995;
  assign po8068 = pi7982;
  assign po8069 = pi8029;
  assign po8070 = pi8032;
  assign po8071 = pi8012;
  assign po8072 = pi7964;
  assign po8073 = pi7932;
  assign po8074 = pi7976;
  assign po8075 = pi7980;
  assign po8076 = pi8007;
  assign po8077 = pi7930;
  assign po8078 = pi7950;
  assign po8079 = pi7981;
  assign po8080 = pi7955;
  assign po8081 = pi7962;
  assign po8082 = pi7967;
  assign po8083 = pi7941;
  assign po8084 = pi7934;
  assign po8085 = pi7993;
  assign po8086 = pi7938;
  assign po8087 = pi8019;
  assign po8088 = pi7956;
  assign po8089 = pi7945;
  assign po8090 = pi8021;
  assign po8091 = pi7996;
  assign po8092 = pi8018;
  assign po8093 = pi7983;
  assign po8094 = pi8035;
  assign po8095 = pi8037;
  assign po8096 = pi8014;
  assign po8097 = pi7970;
  assign po8098 = pi8026;
  assign po8099 = pi8009;
  assign po8100 = pi7944;
  assign po8101 = pi7960;
  assign po8102 = pi8059;
  assign po8103 = pi8091;
  assign po8104 = pi8043;
  assign po8105 = pi8071;
  assign po8106 = pi8040;
  assign po8107 = pi8082;
  assign po8108 = pi8046;
  assign po8109 = pi8053;
  assign po8110 = pi8086;
  assign po8111 = pi8088;
  assign po8112 = pi8056;
  assign po8113 = pi8070;
  assign po8114 = pi8061;
  assign po8115 = pi8047;
  assign po8116 = pi8084;
  assign po8117 = pi8054;
  assign po8118 = pi8078;
  assign po8119 = pi8081;
  assign po8120 = pi8057;
  assign po8121 = pi8063;
  assign po8122 = pi8087;
  assign po8123 = pi8092;
  assign po8124 = pi8072;
  assign po8125 = pi8068;
  assign po8126 = pi8049;
  assign po8127 = pi8073;
  assign po8128 = pi8064;
  assign po8129 = pi8058;
  assign po8130 = pi8069;
  assign po8131 = pi8074;
  assign po8132 = pi8066;
  assign po8133 = pi8055;
  assign po8134 = pi8051;
  assign po8135 = pi8050;
  assign po8136 = pi8065;
  assign po8137 = pi8042;
  assign po8138 = pi8060;
  assign po8139 = pi8094;
  assign po8140 = pi8083;
  assign po8141 = pi8044;
  assign po8142 = pi8045;
  assign po8143 = pi8095;
  assign po8144 = pi8090;
  assign po8145 = pi8089;
  assign po8146 = pi8085;
  assign po8147 = pi8067;
  assign po8148 = pi8079;
  assign po8149 = pi8052;
  assign po8150 = pi8076;
  assign po8151 = pi8041;
  assign po8152 = pi8077;
  assign po8153 = pi8048;
  assign po8154 = pi8080;
  assign po8155 = pi8093;
  assign po8156 = pi8062;
  assign po8157 = pi8075;
  assign po8270 = pi8125;
  assign po8271 = pi8099;
  assign po8272 = pi8131;
  assign po8273 = pi8096;
  assign po8274 = pi8134;
  assign po8275 = pi8097;
  assign po8276 = pi8123;
  assign po8277 = pi8145;
  assign po8278 = pi8142;
  assign po8279 = pi8135;
  assign po8280 = pi8098;
  assign po8281 = pi8103;
  assign po8282 = pi8129;
  assign po8283 = pi8122;
  assign po8284 = pi8109;
  assign po8285 = pi8149;
  assign po8286 = pi8128;
  assign po8287 = pi8138;
  assign po8288 = pi8108;
  assign po8289 = pi8100;
  assign po8290 = pi8111;
  assign po8291 = pi8124;
  assign po8292 = pi8139;
  assign po8293 = pi8116;
  assign po8294 = pi8140;
  assign po8295 = pi8137;
  assign po8296 = pi8148;
  assign po8297 = pi8120;
  assign po8298 = pi8107;
  assign po8299 = pi8114;
  assign po8300 = pi8126;
  assign po8301 = pi8102;
  assign po8302 = pi8130;
  assign po8303 = pi8150;
  assign po8304 = pi8115;
  assign po8305 = pi8112;
  assign po8306 = pi8133;
  assign po8307 = pi8117;
  assign po8308 = pi8104;
  assign po8309 = pi8143;
  assign po8310 = pi8144;
  assign po8311 = pi8106;
  assign po8312 = pi8147;
  assign po8313 = pi8118;
  assign po8314 = pi8113;
  assign po8315 = pi8110;
  assign po8316 = pi8119;
  assign po8317 = pi8151;
  assign po8318 = pi8121;
  assign po8319 = pi8101;
  assign po8320 = pi8132;
  assign po8321 = pi8141;
  assign po8322 = pi8105;
  assign po8323 = pi8136;
  assign po8324 = pi8146;
  assign po8325 = pi8127;
  assign po8326 = pi8184;
  assign po8327 = pi8203;
  assign po8328 = pi8163;
  assign po8329 = pi8205;
  assign po8330 = pi8158;
  assign po8331 = pi8202;
  assign po8332 = pi8178;
  assign po8333 = pi8177;
  assign po8334 = pi8193;
  assign po8335 = pi8195;
  assign po8336 = pi8155;
  assign po8337 = pi8179;
  assign po8338 = pi8198;
  assign po8339 = pi8187;
  assign po8340 = pi8191;
  assign po8341 = pi8156;
  assign po8342 = pi8173;
  assign po8343 = pi8160;
  assign po8344 = pi8189;
  assign po8345 = pi8152;
  assign po8346 = pi8186;
  assign po8347 = pi8188;
  assign po8348 = pi8197;
  assign po8349 = pi8196;
  assign po8350 = pi8181;
  assign po8351 = pi8182;
  assign po8352 = pi8185;
  assign po8353 = pi8183;
  assign po8354 = pi8207;
  assign po8355 = pi8171;
  assign po8356 = pi8157;
  assign po8357 = pi8167;
  assign po8358 = pi8199;
  assign po8359 = pi8153;
  assign po8360 = pi8175;
  assign po8361 = pi8154;
  assign po8362 = pi8170;
  assign po8363 = pi8161;
  assign po8364 = pi8194;
  assign po8365 = pi8166;
  assign po8366 = pi8201;
  assign po8367 = pi8200;
  assign po8368 = pi8190;
  assign po8369 = pi8164;
  assign po8370 = pi8169;
  assign po8371 = pi8176;
  assign po8372 = pi8159;
  assign po8373 = pi8165;
  assign po8374 = pi8174;
  assign po8375 = pi8206;
  assign po8376 = pi8162;
  assign po8377 = pi8204;
  assign po8378 = pi8172;
  assign po8379 = pi8168;
  assign po8380 = pi8180;
  assign po8381 = pi8192;
  assign po8382 = pi8226;
  assign po8383 = pi8258;
  assign po8384 = pi8262;
  assign po8385 = pi8221;
  assign po8386 = pi8242;
  assign po8387 = pi8215;
  assign po8388 = pi8249;
  assign po8389 = pi8240;
  assign po8390 = pi8260;
  assign po8391 = pi8227;
  assign po8392 = pi8235;
  assign po8393 = pi8231;
  assign po8394 = pi8212;
  assign po8395 = pi8225;
  assign po8396 = pi8234;
  assign po8397 = pi8255;
  assign po8398 = pi8253;
  assign po8399 = pi8230;
  assign po8400 = pi8229;
  assign po8401 = pi8236;
  assign po8402 = pi8219;
  assign po8403 = pi8228;
  assign po8404 = pi8250;
  assign po8405 = pi8224;
  assign po8406 = pi8256;
  assign po8407 = pi8252;
  assign po8408 = pi8263;
  assign po8409 = pi8237;
  assign po8410 = pi8246;
  assign po8411 = pi8245;
  assign po8412 = pi8243;
  assign po8413 = pi8217;
  assign po8414 = pi8241;
  assign po8415 = pi8248;
  assign po8416 = pi8213;
  assign po8417 = pi8216;
  assign po8418 = pi8218;
  assign po8419 = pi8222;
  assign po8420 = pi8209;
  assign po8421 = pi8211;
  assign po8422 = pi8223;
  assign po8423 = pi8254;
  assign po8424 = pi8247;
  assign po8425 = pi8208;
  assign po8426 = pi8214;
  assign po8427 = pi8244;
  assign po8428 = pi8220;
  assign po8429 = pi8257;
  assign po8430 = pi8232;
  assign po8431 = pi8251;
  assign po8432 = pi8259;
  assign po8433 = pi8239;
  assign po8434 = pi8210;
  assign po8435 = pi8233;
  assign po8436 = pi8261;
  assign po8437 = pi8238;
  assign po8438 = pi8273;
  assign po8439 = pi8306;
  assign po8440 = pi8315;
  assign po8441 = pi8311;
  assign po8442 = pi8299;
  assign po8443 = pi8296;
  assign po8444 = pi8301;
  assign po8445 = pi8295;
  assign po8446 = pi8274;
  assign po8447 = pi8280;
  assign po8448 = pi8271;
  assign po8449 = pi8310;
  assign po8450 = pi8272;
  assign po8451 = pi8304;
  assign po8452 = pi8302;
  assign po8453 = pi8282;
  assign po8454 = pi8270;
  assign po8455 = pi8285;
  assign po8456 = pi8314;
  assign po8457 = pi8313;
  assign po8458 = pi8279;
  assign po8459 = pi8278;
  assign po8460 = pi8281;
  assign po8461 = pi8275;
  assign po8462 = pi8266;
  assign po8463 = pi8298;
  assign po8464 = pi8297;
  assign po8465 = pi8303;
  assign po8466 = pi8265;
  assign po8467 = pi8312;
  assign po8468 = pi8289;
  assign po8469 = pi8309;
  assign po8470 = pi8288;
  assign po8471 = pi8269;
  assign po8472 = pi8300;
  assign po8473 = pi8284;
  assign po8474 = pi8268;
  assign po8475 = pi8318;
  assign po8476 = pi8277;
  assign po8477 = pi8292;
  assign po8478 = pi8316;
  assign po8479 = pi8317;
  assign po8480 = pi8290;
  assign po8481 = pi8286;
  assign po8482 = pi8319;
  assign po8483 = pi8307;
  assign po8484 = pi8294;
  assign po8485 = pi8293;
  assign po8486 = pi8276;
  assign po8487 = pi8283;
  assign po8488 = pi8291;
  assign po8489 = pi8308;
  assign po8490 = pi8287;
  assign po8491 = pi8264;
  assign po8492 = pi8267;
  assign po8493 = pi8305;
  assign po8494 = pi8365;
  assign po8495 = pi8348;
  assign po8496 = pi8354;
  assign po8497 = pi8341;
  assign po8498 = pi8327;
  assign po8499 = pi8339;
  assign po8500 = pi8340;
  assign po8501 = pi8331;
  assign po8502 = pi8328;
  assign po8503 = pi8325;
  assign po8504 = pi8369;
  assign po8505 = pi8371;
  assign po8506 = pi8364;
  assign po8507 = pi8336;
  assign po8508 = pi8329;
  assign po8509 = pi8338;
  assign po8510 = pi8363;
  assign po8511 = pi8346;
  assign po8512 = pi8333;
  assign po8513 = pi8361;
  assign po8514 = pi8349;
  assign po8515 = pi8326;
  assign po8516 = pi8332;
  assign po8517 = pi8356;
  assign po8518 = pi8362;
  assign po8519 = pi8347;
  assign po8520 = pi8367;
  assign po8521 = pi8352;
  assign po8522 = pi8324;
  assign po8523 = pi8330;
  assign po8524 = pi8360;
  assign po8525 = pi8322;
  assign po8526 = pi8374;
  assign po8527 = pi8343;
  assign po8528 = pi8370;
  assign po8529 = pi8337;
  assign po8530 = pi8372;
  assign po8531 = pi8355;
  assign po8532 = pi8353;
  assign po8533 = pi8345;
  assign po8534 = pi8334;
  assign po8535 = pi8335;
  assign po8536 = pi8350;
  assign po8537 = pi8359;
  assign po8538 = pi8321;
  assign po8539 = pi8375;
  assign po8540 = pi8358;
  assign po8541 = pi8351;
  assign po8542 = pi8366;
  assign po8543 = pi8323;
  assign po8544 = pi8368;
  assign po8545 = pi8342;
  assign po8546 = pi8373;
  assign po8547 = pi8344;
  assign po8548 = pi8320;
  assign po8549 = pi8357;
  assign po8550 = pi8407;
  assign po8551 = pi8383;
  assign po8552 = pi8398;
  assign po8553 = pi8418;
  assign po8554 = pi8394;
  assign po8555 = pi8382;
  assign po8556 = pi8430;
  assign po8557 = pi8409;
  assign po8558 = pi8390;
  assign po8559 = pi8389;
  assign po8560 = pi8401;
  assign po8561 = pi8406;
  assign po8562 = pi8376;
  assign po8563 = pi8427;
  assign po8564 = pi8413;
  assign po8565 = pi8379;
  assign po8566 = pi8412;
  assign po8567 = pi8403;
  assign po8568 = pi8419;
  assign po8569 = pi8391;
  assign po8570 = pi8426;
  assign po8571 = pi8425;
  assign po8572 = pi8402;
  assign po8573 = pi8414;
  assign po8574 = pi8411;
  assign po8575 = pi8385;
  assign po8576 = pi8377;
  assign po8577 = pi8395;
  assign po8578 = pi8424;
  assign po8579 = pi8423;
  assign po8580 = pi8422;
  assign po8581 = pi8408;
  assign po8582 = pi8388;
  assign po8583 = pi8393;
  assign po8584 = pi8387;
  assign po8585 = pi8392;
  assign po8586 = pi8410;
  assign po8587 = pi8380;
  assign po8588 = pi8396;
  assign po8589 = pi8421;
  assign po8590 = pi8386;
  assign po8591 = pi8420;
  assign po8592 = pi8381;
  assign po8593 = pi8384;
  assign po8594 = pi8429;
  assign po8595 = pi8431;
  assign po8596 = pi8416;
  assign po8597 = pi8397;
  assign po8598 = pi8378;
  assign po8599 = pi8400;
  assign po8600 = pi8417;
  assign po8601 = pi8399;
  assign po8602 = pi8405;
  assign po8603 = pi8404;
  assign po8604 = pi8428;
  assign po8605 = pi8415;
  assign po8606 = pi8463;
  assign po8607 = pi8480;
  assign po8608 = pi8481;
  assign po8609 = pi8456;
  assign po8610 = pi8439;
  assign po8611 = pi8455;
  assign po8612 = pi8447;
  assign po8613 = pi8451;
  assign po8614 = pi8448;
  assign po8615 = pi8437;
  assign po8616 = pi8436;
  assign po8617 = pi8457;
  assign po8618 = pi8468;
  assign po8619 = pi8452;
  assign po8620 = pi8446;
  assign po8621 = pi8469;
  assign po8622 = pi8434;
  assign po8623 = pi8484;
  assign po8624 = pi8474;
  assign po8625 = pi8473;
  assign po8626 = pi8466;
  assign po8627 = pi8470;
  assign po8628 = pi8485;
  assign po8629 = pi8433;
  assign po8630 = pi8479;
  assign po8631 = pi8432;
  assign po8632 = pi8454;
  assign po8633 = pi8453;
  assign po8634 = pi8444;
  assign po8635 = pi8461;
  assign po8636 = pi8460;
  assign po8637 = pi8482;
  assign po8638 = pi8443;
  assign po8639 = pi8458;
  assign po8640 = pi8449;
  assign po8641 = pi8467;
  assign po8642 = pi8487;
  assign po8643 = pi8486;
  assign po8644 = pi8464;
  assign po8645 = pi8478;
  assign po8646 = pi8440;
  assign po8647 = pi8472;
  assign po8648 = pi8477;
  assign po8649 = pi8476;
  assign po8650 = pi8459;
  assign po8651 = pi8475;
  assign po8652 = pi8438;
  assign po8653 = pi8462;
  assign po8654 = pi8441;
  assign po8655 = pi8471;
  assign po8656 = pi8435;
  assign po8657 = pi8483;
  assign po8658 = pi8445;
  assign po8659 = pi8442;
  assign po8660 = pi8465;
  assign po8661 = pi8450;
  assign po8662 = pi8493;
  assign po8663 = pi8542;
  assign po8664 = pi8510;
  assign po8665 = pi8512;
  assign po8666 = pi8515;
  assign po8667 = pi8508;
  assign po8668 = pi8495;
  assign po8669 = pi8524;
  assign po8670 = pi8527;
  assign po8671 = pi8513;
  assign po8672 = pi8505;
  assign po8673 = pi8517;
  assign po8674 = pi8529;
  assign po8675 = pi8500;
  assign po8676 = pi8534;
  assign po8677 = pi8525;
  assign po8678 = pi8546;
  assign po8679 = pi8492;
  assign po8680 = pi8543;
  assign po8681 = pi8537;
  assign po8682 = pi8504;
  assign po8683 = pi8496;
  assign po8684 = pi8516;
  assign po8685 = pi8545;
  assign po8686 = pi8535;
  assign po8687 = pi8541;
  assign po8688 = pi8540;
  assign po8689 = pi8532;
  assign po8690 = pi8533;
  assign po8691 = pi8523;
  assign po8692 = pi8536;
  assign po8693 = pi8498;
  assign po8694 = pi8531;
  assign po8695 = pi8522;
  assign po8696 = pi8490;
  assign po8697 = pi8502;
  assign po8698 = pi8518;
  assign po8699 = pi8530;
  assign po8700 = pi8544;
  assign po8701 = pi8521;
  assign po8702 = pi8488;
  assign po8703 = pi8489;
  assign po8704 = pi8526;
  assign po8705 = pi8501;
  assign po8706 = pi8519;
  assign po8707 = pi8514;
  assign po8708 = pi8538;
  assign po8709 = pi8497;
  assign po8710 = pi8509;
  assign po8711 = pi8506;
  assign po8712 = pi8511;
  assign po8713 = pi8499;
  assign po8714 = pi8491;
  assign po8715 = pi8494;
  assign po8716 = pi8539;
  assign po8717 = pi8507;
  assign po8718 = pi8617;
  assign po8719 = pi8596;
  assign po8720 = pi8562;
  assign po8721 = pi8604;
  assign po8722 = pi8608;
  assign po8723 = pi8588;
  assign po8724 = pi8586;
  assign po8725 = pi8618;
  assign po8726 = pi8577;
  assign po8727 = pi8595;
  assign po8728 = pi8593;
  assign po8729 = pi8574;
  assign po8730 = pi8551;
  assign po8731 = pi8581;
  assign po8732 = pi8567;
  assign po8733 = pi8742;
  assign po8734 = pi8578;
  assign po8735 = pi8623;
  assign po8736 = pi8614;
  assign po8737 = pi8611;
  assign po8738 = pi8612;
  assign po8739 = pi8563;
  assign po8740 = pi8566;
  assign po8741 = pi8589;
  assign po8742 = pi8571;
  assign po8743 = pi8626;
  assign po8744 = pi8587;
  assign po8745 = pi8552;
  assign po8746 = pi8564;
  assign po8747 = pi8616;
  assign po8748 = pi8573;
  assign po8749 = pi8610;
  assign po8750 = pi8752;
  assign po8751 = pi8591;
  assign po8752 = pi8607;
  assign po8753 = pi8620;
  assign po8754 = pi8572;
  assign po8755 = pi8576;
  assign po8756 = pi8560;
  assign po8757 = pi8584;
  assign po8758 = pi8802;
  assign po8759 = pi8553;
  assign po8760 = pi8619;
  assign po8761 = pi8598;
  assign po8762 = pi8627;
  assign po8763 = pi8606;
  assign po8764 = pi8603;
  assign po8765 = pi8555;
  assign po8766 = pi8621;
  assign po8767 = pi8569;
  assign po8768 = pi8625;
  assign po8769 = pi8558;
  assign po8770 = pi8613;
  assign po8771 = pi8599;
  assign po8772 = pi8580;
  assign po8773 = pi8565;
  assign po8774 = pi8609;
  assign po8775 = pi8597;
  assign po8776 = pi8590;
  assign po8777 = pi8748;
  assign po8778 = pi8713;
  assign po8779 = pi8712;
  assign po8780 = pi8726;
  assign po8781 = pi8687;
  assign po8782 = pi8653;
  assign po8783 = pi8631;
  assign po8784 = pi8782;
  assign po8785 = pi8661;
  assign po8786 = pi8766;
  assign po8787 = pi8761;
  assign po8788 = pi8657;
  assign po8789 = pi8803;
  assign po8790 = pi8658;
  assign po8791 = pi8796;
  assign po8792 = pi8632;
  assign po8793 = pi8683;
  assign po8794 = pi8676;
  assign po8795 = pi8636;
  assign po8796 = pi8679;
  assign po8797 = pi8643;
  assign po8798 = pi8727;
  assign po8799 = pi8674;
  assign po8800 = pi8776;
  assign po8801 = pi8656;
  assign po8802 = pi8677;
  assign po8803 = pi8647;
  assign po8804 = pi8655;
  assign po8805 = pi8781;
  assign po8806 = pi8639;
  assign po8807 = pi8659;
  assign po8808 = pi8663;
  assign po8809 = pi8717;
  assign po8810 = pi8654;
  assign po8811 = pi8641;
  assign po8812 = pi8743;
  assign po8813 = pi8719;
  assign po8814 = pi8640;
  assign po8815 = pi8773;
  assign po8816 = pi8644;
  assign po8817 = pi8637;
  assign po8818 = pi8686;
  assign po8819 = pi8634;
  assign po8820 = pi8638;
  assign po8821 = pi8672;
  assign po8822 = pi8795;
  assign po8823 = pi8667;
  assign po8824 = pi8738;
  assign po8825 = pi8645;
  assign po8826 = pi8662;
  assign po8827 = pi8642;
  assign po8828 = pi8673;
  assign po8829 = pi8664;
  assign po8830 = pi8715;
  assign po8831 = pi8778;
  assign po8832 = pi8775;
  assign po8833 = pi8652;
  assign po8834 = pi8660;
  assign po8835 = pi8705;
  assign po8836 = pi8650;
  assign po8837 = pi8630;
  assign po8838 = pi8648;
  assign po8839 = pi8681;
  assign po8840 = pi8668;
  assign po8841 = pi8670;
  assign po8842 = pi8675;
  assign po8843 = pi8635;
  assign po8844 = pi8628;
  assign po8845 = pi8750;
  assign po8846 = pi8684;
  assign po8847 = pi8680;
  assign po8848 = pi8669;
  assign po8849 = pi8646;
  assign po8850 = pi8671;
  assign po8851 = pi8651;
  assign po8852 = pi8798;
  assign po8853 = pi8682;
  assign po8854 = pi8799;
  assign po8855 = pi8665;
  assign po8856 = pi8649;
  assign po8857 = pi8666;
  assign po8858 = pi8794;
  assign po8859 = pi8807;
  assign po8860 = pi8737;
  assign po8861 = pi8732;
  assign po8862 = pi8792;
  assign po8863 = pi8702;
  assign po8864 = pi8774;
  assign po8865 = pi8791;
  assign po8866 = pi8731;
  assign po8867 = pi8733;
  assign po8868 = pi8694;
  assign po8869 = pi8756;
  assign po8870 = pi8758;
  assign po8871 = pi8801;
  assign po8872 = pi8706;
  assign po8873 = pi8711;
  assign po8874 = pi8703;
  assign po8875 = pi8730;
  assign po8876 = pi8740;
  assign po8877 = pi8800;
  assign po8878 = pi8757;
  assign po8879 = pi8739;
  assign po8880 = pi8741;
  assign po8881 = pi8699;
  assign po8882 = pi8759;
  assign po8883 = pi8764;
  assign po8884 = pi8692;
  assign po8885 = pi8690;
  assign po8886 = pi8691;
  assign po8887 = pi8760;
  assign po8888 = pi8698;
  assign po8889 = pi8700;
  assign po8890 = pi8786;
  assign po8891 = pi8704;
  assign po8892 = pi8708;
  assign po8893 = pi8785;
  assign po8894 = pi8736;
  assign po8895 = pi8724;
  assign po8896 = pi8789;
  assign po8897 = pi8805;
  assign po8898 = pi8762;
  assign po8899 = pi8689;
  assign po8900 = pi8777;
  assign po8901 = pi8745;
  assign po8902 = pi8804;
  assign po8903 = pi8770;
  assign po8904 = pi8746;
  assign po8905 = pi8707;
  assign po8906 = pi8723;
  assign po8907 = pi8688;
  assign po8908 = pi8772;
  assign po8909 = pi8735;
  assign po8910 = pi8728;
  assign po8911 = pi8734;
  assign po8912 = pi8783;
  assign po8913 = pi8769;
  assign po8914 = pi8780;
  assign po8915 = pi8710;
  assign po8916 = pi8763;
  assign po8917 = pi8806;
  assign po8918 = pi8951;
  assign po8919 = pi8947;
  assign po8920 = pi8966;
  assign po8921 = pi8941;
  assign po8922 = pi8932;
  assign po8923 = pi8818;
  assign po8924 = pi8975;
  assign po8925 = pi8834;
  assign po8926 = pi8840;
  assign po8927 = pi8808;
  assign po8928 = pi8963;
  assign po8929 = pi8958;
  assign po8930 = pi8961;
  assign po8931 = pi8816;
  assign po8932 = pi8827;
  assign po8933 = pi8979;
  assign po8934 = pi8952;
  assign po8935 = pi8841;
  assign po8936 = pi8943;
  assign po8937 = pi8971;
  assign po8938 = pi8972;
  assign po8939 = pi8850;
  assign po8940 = pi8825;
  assign po8941 = pi8956;
  assign po8942 = pi8833;
  assign po8943 = pi8871;
  assign po8944 = pi8826;
  assign po8945 = pi8823;
  assign po8946 = pi8828;
  assign po8947 = pi8817;
  assign po8948 = pi8862;
  assign po8949 = pi8815;
  assign po8950 = pi8830;
  assign po8951 = pi8854;
  assign po8952 = pi8820;
  assign po8953 = pi8939;
  assign po8954 = pi8970;
  assign po8955 = pi8842;
  assign po8956 = pi8863;
  assign po8957 = pi8851;
  assign po8958 = pi8938;
  assign po8959 = pi8844;
  assign po8960 = pi8981;
  assign po8961 = pi8967;
  assign po8962 = pi8945;
  assign po8963 = pi8973;
  assign po8964 = pi8965;
  assign po8965 = pi8937;
  assign po8966 = pi8959;
  assign po8967 = pi8982;
  assign po8968 = pi8859;
  assign po8969 = pi8968;
  assign po8970 = pi8928;
  assign po8971 = pi8977;
  assign po8972 = pi8835;
  assign po8973 = pi8855;
  assign po8974 = pi8870;
  assign po8975 = pi8936;
  assign po8976 = pi8946;
  assign po8977 = pi8866;
  assign po8978 = pi8809;
  assign po8979 = pi8846;
  assign po8980 = pi8813;
  assign po8981 = pi8810;
  assign po8982 = pi8869;
  assign po8983 = pi8868;
  assign po8984 = pi8856;
  assign po8985 = pi8824;
  assign po8986 = pi8957;
  assign po8987 = pi8969;
  assign po8988 = pi8934;
  assign po8989 = pi8935;
  assign po8990 = pi8940;
  assign po8991 = pi8847;
  assign po8992 = pi8955;
  assign po8993 = pi8933;
  assign po8994 = pi8949;
  assign po8995 = pi8822;
  assign po8996 = pi8857;
  assign po8997 = pi8858;
  assign po8998 = pi8860;
  assign po8999 = pi8948;
  assign po9000 = pi8962;
  assign po9001 = pi8832;
  assign po9002 = pi8861;
  assign po9003 = pi8845;
  assign po9004 = pi8976;
  assign po9005 = pi8837;
  assign po9006 = pi8839;
  assign po9007 = pi8953;
  assign po9008 = pi8853;
  assign po9009 = pi8814;
  assign po9010 = pi8964;
  assign po9011 = pi8811;
  assign po9012 = pi8821;
  assign po9013 = pi8942;
  assign po9014 = pi8848;
  assign po9015 = pi8974;
  assign po9016 = pi8960;
  assign po9017 = pi8864;
  assign po9018 = pi8836;
  assign po9019 = pi8954;
  assign po9020 = pi8838;
  assign po9021 = pi8930;
  assign po9022 = pi8929;
  assign po9023 = pi8852;
  assign po9024 = pi8983;
  assign po9025 = pi8829;
  assign po9026 = pi8865;
  assign po9027 = pi8812;
  assign po9028 = pi8831;
  assign po9029 = pi8819;
  assign po9030 = pi8950;
  assign po9031 = pi8980;
  assign po9032 = pi8867;
  assign po9033 = pi8843;
  assign po9034 = pi8931;
  assign po9035 = pi8944;
  assign po9036 = pi8978;
  assign po9037 = pi8849;
endmodule


