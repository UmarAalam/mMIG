//Written by the Majority Logic Package Thu Apr 30 22:51:15 2015
module top (
            pi00, pi01, pi02, pi03, pi04, pi05, pi06, pi07, pi08, pi09, pi10, pi11, pi12, pi13, pi14, pi15, pi16, pi17, pi18, pi19, pi20, pi21, pi22, pi23, pi24, pi25, pi26, pi27, pi28, pi29, pi30, pi31, 
            po00, po01, po02, po03, po04, po05, po06, po07, po08, po09, po10, po11, po12, po13, po14, po15, po16, po17, po18, po19, po20, po21, po22, po23, po24, po25, po26, po27, po28, po29, po30, po31);
input pi00, pi01, pi02, pi03, pi04, pi05, pi06, pi07, pi08, pi09, pi10, pi11, pi12, pi13, pi14, pi15, pi16, pi17, pi18, pi19, pi20, pi21, pi22, pi23, pi24, pi25, pi26, pi27, pi28, pi29, pi30, pi31;
output po00, po01, po02, po03, po04, po05, po06, po07, po08, po09, po10, po11, po12, po13, po14, po15, po16, po17, po18, po19, po20, po21, po22, po23, po24, po25, po26, po27, po28, po29, po30, po31;
wire one, v0, v1, v2, v3, v4, v5, v6, v7, v8, v9, v10, v11, v12, v13, v14, v15, v16, v17, v18, v19, v20, v21, v22, v23, v24, v25, v26, v27, v28, v29, v30, v31, v32, v33, v34, v35, v36, v37, v38, v39, v40, v41, v42, v43, v44, v45, v46, v47, v48, v49, v50, v51, v52, v53, v54, v55, v56, v57, v58, v59, v60, v61, v62, v63, v64, v65, v66, v67, v68, v69, v70, v71, v72, v73, v74, v75, v76, v77, v78, v79, v80, v81, v82, v83, v84, v85, v86, v87, v88, v89, v90, v91, v92, v93, v94, v95, v96, v97, v98, v99, v100, v101, v102, v103, v104, v105, v106, v107, v108, v109, v110, v111, v112, v113, v114, v115, v116, v117, v118, v119, v120, v121, v122, v123, v124, v125, v126, v127, v128, v129, v130, v131, v132, v133, v134, v135, v136, v137, v138, v139, v140, v141, v142, v143, v144, v145, v146, v147, v148, v149, v150, v151, v152, v153, v154, v155, v156, v157, v158, v159, v160, v161, v162, v163, v164, v165, v166, v167, v168, v169, v170, v171, v172, v173, v174, v175, v176, v177, v178, v179, v180, v181, v182, v183, v184, v185, v186, v187, v188, v189, v190, v191, v192, v193, v194, v195, v196, v197, v198, v199, v200, v201, v202, v203, v204, v205, v206, v207, v208, v209, v210, v211, v212, v213, v214, v215, v216, v217, v218, v219, v220, v221, v222, v223, v224, v225, v226, v227, v228, v229, v230, v231, v232, v233, v234, v235, v236, v237, v238, v239, v240, v241, v242, v243, v244, v245, v246, v247, v248, v249, v250, v251, v252, v253, v254, v255, v256, v257, v258, v259, v260, v261, v262, v263, v264, v265, v266, v267, v268, v269, v270, v271, v272, v273, v274, v275, v276, v277, v278, v279, v280, v281, v282, v283, v284, v285, v286, v287, v288, v289, v290, v291, v292, v293, v294, v295, v296, v297, v298, v299, v300, v301, v302, v303, v304, v305, v306, v307, v308, v309, v310, v311, v312, v313, v314, v315, v316, v317, v318, v319, v320, v321, v322, v323, v324, v325, v326, v327, v328, v329, v330, v331, v332, v333, v334, v335, v336, v337, v338, v339, v340, v341, v342, v343, v344, v345, v346, v347, v348, v349, v350, v351, v352, v353, v354, v355, v356, v357, v358, v359, v360, v361, v362, v363, v364, v365, v366, v367, v368, v369, v370, v371, v372, v373, v374, v375, v376, v377, v378, v379, v380, v381, v382, v383, v384, v385, v386, v387, v388, v389, v390, v391, v392, v393, v394, v395, v396, v397, v398, v399, v400, v401, v402, v403, v404, v405, v406, v407, v408, v409, v410, v411, v412, v413, v414, v415, v416, v417, v418, v419, v420, v421, v422, v423, v424, v425, v426, v427, v428, v429, v430, v431, v432, v433, v434, v435, v436, v437, v438, v439, v440, v441, v442, v443, v444, v445, v446, v447, v448, v449, v450, v451, v452, v453, v454, v455, v456, v457, v458, v459, v460, v461, v462, v463, v464, v465, v466, v467, v468, v469, v470, v471, v472, v473, v474, v475, v476, v477, v478, v479, v480, v481, v482, v483, v484, v485, v486, v487, v488, v489, v490, v491, v492, v493, v494, v495, v496, v497, v498, v499, v500, v501, v502, v503, v504, v505, v506, v507, v508, v509, v510, v511, v512, v513, v514, v515, v516, v517, v518, v519, v520, v521, v522, v523, v524, v525, v526, v527, v528, v529, v530, v531, v532, v533, v534, v535, v536, v537, v538, v539, v540, v541, v542, v543, v544, v545, v546, v547, v548, v549, v550, v551, v552, v553, v554, v555, v556, v557, v558, v559, v560, v561, v562, v563, v564, v565, v566, v567, v568, v569, v570, v571, v572, v573, v574, v575, v576, v577, v578, v579, v580, v581, v582, v583, v584, v585, v586, v587, v588, v589, v590, v591, v592, v593, v594, v595, v596, v597, v598, v599, v600, v601, v602, v603, v604, v605, v606, v607, v608, v609, v610, v611, v612, v613, v614, v615, v616, v617, v618, v619, v620, v621, v622, v623, v624, v625, v626, v627, v628, v629, v630, v631, v632, v633, v634, v635, v636, v637, v638, v639, v640, v641, v642, v643, v644, v645, v646, v647, v648, v649, v650, v651, v652, v653, v654, v655, v656, v657, v658, v659, v660, v661, v662, v663, v664, v665, v666, v667, v668, v669, v670, v671, v672, v673, v674, v675, v676, v677, v678, v679, v680, v681, v682, v683, v684, v685, v686, v687, v688, v689, v690, v691, v692, v693, v694, v695, v696, v697, v698, v699, v700, v701, v702, v703, v704, v705, v706, v707, v708, v709, v710, v711, v712, v713, v714, v715, v716, v717, v718, v719, v720, v721, v722, v723, v724, v725, v726, v727, v728, v729, v730, v731, v732, v733, v734, v735, v736, v737, v738, v739, v740, v741, v742, v743, v744, v745, v746, v747, v748, v749, v750, v751, v752, v753, v754, v755, v756, v757, v758, v759, v760, v761, v762, v763, v764, v765, v766, v767, v768, v769, v770, v771, v772, v773, v774, v775, v776, v777, v778, v779, v780, v781, v782, v783, v784, v785, v786, v787, v788, v789, v790, v791, v792, v793, v794, v795, v796, v797, v798, v799, v800, v801, 
w0, w1, w2, w3, w4, w5, w6, w7, w8, w9, w10, w11, w12, w13, w14, w15, w16, w17, w18, w19, w20, w21, w22, w23, w24, w25, w26, w27, w28, w29, w30, w31, w32, w33, w34, w35, w36, w37, w38, w39, w40, w41, w42, w43, w44, w45, w46, w47, w48, w49, w50, w51, w52, w53, w54, w55, w56, w57, w58, w59, w60, w61, w62, w63, w64, w65, w66, w67, w68, w69, w70, w71, w72, w73, w74, w75, w76, w77, w78, w79, w80, w81, w82, w83, w84, w85, w86, w87, w88, w89, w90, w91, w92, w93, w94, w95, w96, w97, w98, w99, w100, w101, w102, w103, w104, w105, w106, w107, w108, w109, w110, w111, w112, w113, w114, w115, w116, w117, w118, w119, w120, w121, w122, w123, w124, w125, w126, w127, w128, w129, w130, w131, w132, w133, w134, w135, w136, w137, w138, w139, w140, w141, w142, w143, w144, w145, w146, w147, w148, w149, w150, w151, w152, w153, w154, w155, w156, w157, w158, w159, w160, w161, w162, w163, w164, w165, w166, w167, w168, w169, w170, w171, w172, w173, w174, w175, w176, w177, w178, w179, w180, w181, w182, w183, w184, w185, w186, w187, w188, w189, w190, w191, w192, w193, w194, w195, w196, w197, w198, w199, w200, w201, w202, w203, w204, w205, w206, w207, w208, w209, w210, w211, w212, w213, w214, w215, w216, w217, w218, w219, w220, w221, w222, w223, w224, w225, w226, w227, w228, w229, w230, w231, w232, w233, w234, w235, w236, w237, w238, w239, w240, w241, w242, w243, w244, w245, w246, w247, w248, w249, w250, w251, w252, w253, w254, w255, w256, w257, w258, w259, w260, w261, w262, w263, w264, w265, w266, w267, w268, w269, w270, w271, w272, w273, w274, w275, w276, w277, w278, w279, w280, w281, w282, w283, w284, w285, w286, w287, w288, w289, w290, w291, w292, w293, w294, w295, w296, w297, w298, w299, w300, w301, w302, w303, w304, w305, w306, w307, w308, w309, w310, w311, w312, w313, w314, w315, w316, w317, w318, w319, w320, w321, w322, w323, w324, w325, w326, w327, w328, w329, w330, w331, w332, w333, w334, w335, w336, w337, w338, w339, w340, w341, w342, w343, w344, w345, w346, w347, w348, w349, w350, w351, w352, w353, w354, w355, w356, w357, w358, w359, w360, w361, w362, w363, w364, w365, w366, w367, w368, w369, w370, w371, w372, w373, w374, w375, w376, w377, w378, w379, w380, w381, w382, w383, w384, w385, w386, w387, w388, w389, w390, w391, w392, w393, w394, w395, w396, w397, w398, w399, w400, w401, w402, w403, w404, w405, w406, w407, w408, w409, w410, w411, w412, w413, w414, w415, w416, w417, w418, w419, w420, w421, w422, w423, w424, w425, w426, w427, w428, w429, w430, w431, w432, w433, w434, w435, w436, w437, w438, w439, w440, w441, w442, w443, w444, w445, w446, w447, w448, w449, w450, w451, w452, w453, w454, w455, w456, w457, w458, w459, w460, w461, w462, w463, w464, w465, w466, w467, w468, w469, w470, w471, w472, w473, w474, w475, w476, w477, w478, w479, w480, w481, w482, w483, w484, w485, w486, w487, w488, w489, w490, w491, w492, w493, w494, w495, w496, w497, w498, w499, w500, w501, w502, w503, w504, w505, w506, w507, w508, w509, w510, w511, w512, w513, w514, w515, w516, w517, w518, w519, w520, w521, w522, w523, w524, w525, w526, w527, w528, w529, w530, w531, w532, w533, w534, w535, w536, w537, w538, w539, w540, w541, w542, w543, w544, w545, w546, w547, w548, w549, w550, w551, w552, w553, w554, w555, w556, w557, w558, w559, w560, w561, w562, w563, w564, w565, w566, w567, w568, w569, w570, w571, w572, w573, w574, w575, w576, w577, w578, w579, w580, w581, w582, w583, w584, w585, w586, w587, w588, w589, w590, w591, w592, w593, w594, w595, w596, w597, w598, w599, w600, w601, w602, w603, w604, w605, w606, w607, w608, w609, w610, w611, w612, w613, w614, w615, w616, w617, w618, w619, w620, w621, w622, w623, w624, w625, w626, w627, w628, w629, w630, w631, w632, w633, w634, w635, w636, w637, w638, w639, w640, w641, w642, w643, w644, w645, w646, w647, w648, w649, w650, w651, w652, w653, w654, w655, w656, w657, w658, w659, w660, w661, w662, w663, w664, w665, w666, w667, w668, w669, w670, w671, w672, w673, w674, w675, w676, w677, w678, w679, w680, w681, w682, w683, w684, w685, w686, w687, w688, w689, w690, w691, w692, w693, w694, w695, w696, w697, w698, w699, w700, w701, w702, w703, w704, w705, w706, w707, w708, w709, w710, w711, w712, w713, w714, w715, w716, w717, w718, w719, w720, w721, w722, w723, w724, w725, w726, w727, w728, w729, w730, w731, w732, w733, w734, w735, w736, w737, w738, w739, w740, w741, w742, w743, w744, w745, w746, w747, w748, w749, w750, w751, w752, w753, w754, w755, w756, w757, w758, w759, w760, w761, w762, w763, w764, w765, w766, w767, w768, w769, w770, w771, w772, w773, w774, w775, w776, w777, w778, w779, w780, w781, w782, w783, w784, w785, w786, w787, w788, w789, w790, w791, w792, w793, w794, w795, w796, w797, w798, w799, w800, w801, w802, w803, w804, w805, w806, w807, w808, w809, w810, w811, w812, w813, w814, w815, w816, w817, w818, w819, w820, w821, w822, w823, w824, w825, w826, w827, w828, w829, w830, w831, w832, w833, w834, w835, w836, w837, w838, w839, w840, w841, w842, w843, w844, w845, w846, w847, w848, w849, w850, w851, w852, w853, w854, w855, w856, w857, w858, w859, w860, w861, w862, w863, w864, w865, w866, w867, w868, w869, w870, w871, w872, w873, w874, w875, w876, w877, w878, w879, w880, w881, w882, w883, w884, w885, w886, w887, w888, w889, w890, w891, w892, w893, w894, w895, w896, w897, w898, w899, w900, w901, w902, w903, w904, w905, w906, w907, w908, w909, w910, w911, w912, w913, w914, w915, w916, w917, w918, w919, w920, w921, w922, w923, w924, w925, w926, w927, w928, w929, w930, w931, w932, w933, w934, w935, w936, w937, w938, w939, w940, w941, w942, w943, w944, w945, w946, w947, w948, w949, w950, w951, w952, w953, w954, w955, w956, w957, w958, w959, w960, w961, w962, w963, w964, w965, w966, w967, w968, w969, w970, w971, w972, w973, w974, w975, w976, w977, w978, w979, w980, w981, w982, w983, w984, w985, w986, w987, w988, w989, w990, w991, w992, w993, w994, w995, w996, w997, w998, w999, w1000, w1001, w1002, w1003, w1004, w1005, w1006, w1007, w1008, w1009, w1010, w1011, w1012, w1013, w1014, w1015, w1016, w1017, w1018, w1019, w1020, w1021, w1022, w1023, w1024, w1025, w1026, w1027, w1028, w1029, w1030, w1031, w1032, w1033, w1034, w1035, w1036, w1037, w1038, w1039, w1040, w1041, w1042, w1043, w1044, w1045, w1046, w1047, w1048, w1049, w1050, w1051, w1052, w1053, w1054, w1055, w1056, w1057, w1058, w1059, w1060, w1061, w1062, w1063, w1064, w1065, w1066, w1067, w1068, w1069, w1070, w1071, w1072, w1073, w1074, w1075, w1076, w1077, w1078, w1079, w1080, w1081, w1082, w1083, w1084, w1085, w1086, w1087, w1088, w1089, w1090, w1091, w1092, w1093, w1094, w1095, w1096, w1097, w1098, w1099, w1100, w1101, w1102, w1103, w1104, w1105, w1106, w1107, w1108, w1109, w1110, w1111, w1112, w1113, w1114, w1115, w1116, w1117, w1118, w1119, w1120, w1121, w1122, w1123, w1124, w1125, w1126, w1127, w1128, w1129, w1130, w1131, w1132, w1133, w1134, w1135, w1136, w1137, w1138, w1139, w1140, w1141, w1142, w1143, w1144, w1145, w1146, w1147, w1148, w1149, w1150, w1151, w1152, w1153, w1154, w1155, w1156, w1157, w1158, w1159, w1160, w1161, w1162, w1163, w1164, w1165, w1166, w1167, w1168, w1169, w1170, w1171, w1172, w1173, w1174, w1175, w1176, w1177, w1178, w1179, w1180, w1181, w1182, w1183, w1184, w1185, w1186, w1187, w1188, w1189, w1190, w1191, w1192, w1193, w1194, w1195, w1196, w1197, w1198, w1199, w1200, w1201, w1202, w1203, w1204, w1205, w1206, w1207, w1208, w1209, w1210, w1211, w1212, w1213, w1214, w1215, w1216, w1217, w1218, w1219, w1220, w1221, w1222, w1223, w1224, w1225, w1226, w1227, w1228, w1229, w1230, w1231, w1232, w1233, w1234, w1235, w1236, w1237, w1238, w1239, w1240, w1241, w1242, w1243, w1244, w1245, w1246, w1247, w1248, w1249, w1250, w1251, w1252, w1253, w1254, w1255, w1256, w1257, w1258, w1259, w1260, w1261, w1262, w1263, w1264, w1265, w1266, w1267, w1268, w1269, w1270, w1271, w1272, w1273, w1274, w1275, w1276, w1277, w1278, w1279, w1280, w1281, w1282, w1283, w1284, w1285, w1286, w1287, w1288, w1289, w1290, w1291, w1292, w1293, w1294, w1295, w1296, w1297, w1298, w1299, w1300, w1301, w1302, w1303, w1304, w1305, w1306, w1307, w1308, w1309, w1310, w1311, w1312, w1313, w1314, w1315, w1316, w1317, w1318, w1319, w1320, w1321, w1322, w1323, w1324, w1325, w1326, w1327, w1328, w1329, w1330, w1331, w1332, w1333, w1334, w1335, w1336, w1337, w1338, w1339, w1340, w1341, w1342, w1343, w1344, w1345, w1346, w1347, w1348, w1349, w1350, w1351, w1352, w1353, w1354, w1355, w1356, w1357, w1358, w1359, w1360, w1361, w1362, w1363, w1364, w1365, w1366, w1367, w1368, w1369, w1370, w1371, w1372, w1373, w1374, w1375, w1376, w1377, w1378, w1379, w1380, w1381, w1382, w1383, w1384, w1385, w1386, w1387, w1388, w1389, w1390, w1391, w1392, w1393, w1394, w1395, w1396, w1397, w1398, w1399, w1400, w1401, w1402, w1403, w1404, w1405, w1406, w1407, w1408, w1409, w1410, w1411, w1412, w1413, w1414, w1415, w1416, w1417, w1418, w1419, w1420, w1421, w1422, w1423, w1424, w1425, w1426, w1427, w1428, w1429, w1430, w1431, w1432, w1433, w1434, w1435, w1436, w1437, w1438, w1439, w1440, w1441, w1442, w1443, w1444, w1445, w1446, w1447, w1448, w1449, w1450, w1451, w1452, w1453, w1454, w1455, w1456, w1457, w1458, w1459, w1460, w1461, w1462, w1463, w1464, w1465, w1466, w1467, w1468, w1469, w1470, w1471, w1472, w1473, w1474, w1475, w1476, w1477, w1478, w1479, w1480, w1481, w1482, w1483, w1484, w1485, w1486, w1487, w1488, w1489, w1490, w1491, w1492, w1493, w1494, w1495, w1496, w1497, w1498, w1499, w1500, w1501, w1502, w1503, w1504, w1505, w1506, w1507, w1508, w1509, w1510, w1511, w1512, w1513, w1514, w1515, w1516, w1517, w1518, w1519, w1520, w1521, w1522, w1523, w1524, w1525, w1526, w1527, w1528, w1529, w1530, w1531, w1532, w1533, w1534, w1535, w1536, w1537, w1538, w1539, w1540, w1541, w1542, w1543, w1544, w1545, w1546, w1547, w1548, w1549, w1550, w1551, w1552, w1553, w1554, w1555, w1556, w1557, w1558, w1559, w1560, w1561, w1562, w1563, w1564, w1565, w1566, w1567, w1568, w1569, w1570, w1571, w1572, w1573, w1574, w1575, w1576, w1577, w1578, w1579, w1580, w1581, w1582, w1583, w1584, w1585, w1586, w1587, w1588, w1589, w1590, w1591, w1592, w1593, w1594, w1595, w1596, w1597, w1598, w1599, w1600, w1601, w1602, w1603, w1604, w1605, w1606, w1607, w1608, w1609, w1610, w1611, w1612, w1613, w1614, w1615, w1616, w1617, w1618, w1619, w1620, w1621, w1622, w1623, w1624, w1625, w1626, w1627, w1628, w1629, w1630, w1631, w1632, w1633, w1634, w1635, w1636, w1637, w1638, w1639, w1640, w1641, w1642, w1643, w1644, w1645, w1646, w1647, w1648, w1649, w1650, w1651, w1652, w1653, w1654, w1655, w1656, w1657, w1658, w1659, w1660, w1661, w1662, w1663, w1664, w1665, w1666, w1667, w1668, w1669, w1670, w1671, w1672, w1673, w1674, w1675, w1676, w1677, w1678, w1679, w1680, w1681, w1682, w1683, w1684, w1685, w1686, w1687, w1688, w1689, w1690, w1691, w1692, w1693, w1694, w1695, w1696, w1697, w1698, w1699, w1700, w1701, w1702, w1703, w1704, w1705, w1706, w1707, w1708, w1709, w1710, w1711, w1712, w1713, w1714, w1715, w1716, w1717, w1718, w1719, w1720, w1721, w1722, w1723, w1724, w1725, w1726, w1727, w1728, w1729, w1730, w1731, w1732, w1733, w1734, w1735, w1736, w1737, w1738, w1739, w1740, w1741, w1742, w1743, w1744, w1745, w1746, w1747, w1748, w1749, w1750, w1751, w1752, w1753, w1754, w1755, w1756, w1757, w1758, w1759, w1760, w1761, w1762, w1763, w1764, w1765, w1766, w1767, w1768, w1769, w1770, w1771, w1772, w1773, w1774, w1775, w1776, w1777, w1778, w1779, w1780, w1781, w1782, w1783, w1784, w1785, w1786, w1787, w1788, w1789, w1790, w1791, w1792, w1793, w1794, w1795, w1796, w1797, w1798, w1799, w1800, w1801, w1802, w1803, w1804, w1805, w1806, w1807, w1808, w1809, w1810, w1811, w1812, w1813, w1814, w1815, w1816, w1817, w1818, w1819, w1820, w1821, w1822, w1823, w1824, w1825, w1826, w1827, w1828, w1829, w1830, w1831, w1832, w1833, w1834, w1835, w1836, w1837, w1838, w1839, w1840, w1841, w1842, w1843, w1844, w1845, w1846, w1847, w1848, w1849, w1850, w1851, w1852, w1853, w1854, w1855, w1856, w1857, w1858, w1859, w1860, w1861, w1862, w1863, w1864, w1865, w1866, w1867, w1868, w1869, w1870, w1871, w1872, w1873, w1874, w1875, w1876, w1877, w1878, w1879, w1880, w1881, w1882, w1883, w1884, w1885, w1886, w1887, w1888, w1889, w1890, w1891, w1892, w1893, w1894, w1895, w1896, w1897, w1898, w1899, w1900, w1901, w1902, w1903, w1904, w1905, w1906, w1907, w1908, w1909, w1910, w1911, w1912, w1913, w1914, w1915, w1916, w1917, w1918, w1919, w1920, w1921, w1922, w1923, w1924, w1925, w1926, w1927, w1928, w1929, w1930, w1931, w1932, w1933, w1934, w1935, w1936, w1937, w1938, w1939, w1940, w1941, w1942, w1943, w1944, w1945, w1946, w1947, w1948, w1949, w1950, w1951, w1952, w1953, w1954, w1955, w1956, w1957, w1958, w1959, w1960, w1961, w1962, w1963, w1964, w1965, w1966, w1967, w1968, w1969, w1970, w1971, w1972, w1973, w1974, w1975, w1976, w1977, w1978, w1979, w1980, w1981, w1982, w1983, w1984, w1985, w1986, w1987, w1988, w1989, w1990, w1991, w1992, w1993, w1994, w1995, w1996, w1997, w1998, w1999, w2000, w2001, w2002, w2003, w2004, w2005, w2006, w2007, w2008, w2009, w2010, w2011, w2012, w2013, w2014, w2015, w2016, w2017, w2018, w2019, w2020, w2021, w2022, w2023, w2024, w2025, w2026, w2027, w2028, w2029, w2030, w2031, w2032, w2033, w2034, w2035, w2036, w2037, w2038, w2039, w2040, w2041, w2042, w2043, w2044, w2045, w2046, w2047, w2048, w2049, w2050, w2051, w2052, w2053, w2054, w2055, w2056, w2057, w2058, w2059, w2060, w2061, w2062, w2063, w2064, w2065, w2066, w2067, w2068, w2069, w2070, w2071, w2072, w2073, w2074, w2075, w2076, w2077, w2078, w2079, w2080, w2081, w2082, w2083, w2084, w2085, w2086, w2087, w2088, w2089, w2090, w2091, w2092, w2093, w2094, w2095, w2096, w2097, w2098, w2099, w2100, w2101, w2102, w2103, w2104, w2105, w2106, w2107, w2108, w2109, w2110, w2111, w2112, w2113, w2114, w2115, w2116, w2117, w2118, w2119, w2120, w2121, w2122, w2123, w2124, w2125, w2126, w2127, w2128, w2129, w2130, w2131, w2132, w2133, w2134, w2135, w2136, w2137, w2138, w2139, w2140, w2141, w2142, w2143, w2144, w2145, w2146, w2147, w2148, w2149, w2150, w2151, w2152, w2153, w2154, w2155, w2156, w2157, w2158, w2159, w2160, w2161, w2162, w2163, w2164, w2165, w2166, w2167, w2168, w2169, w2170, w2171, w2172, w2173, w2174, w2175, w2176, w2177, w2178, w2179, w2180, w2181, w2182, w2183, w2184, w2185, w2186, w2187, w2188, w2189, w2190, w2191, w2192, w2193, w2194, w2195, w2196, w2197, w2198, w2199, w2200, w2201, w2202, w2203, w2204, w2205, w2206, w2207, w2208, w2209, w2210, w2211, w2212, w2213, w2214, w2215, w2216, w2217, w2218, w2219, w2220, w2221, w2222, w2223, w2224, w2225, w2226, w2227, w2228, w2229, w2230, w2231, w2232, w2233, w2234, w2235, w2236, w2237, w2238, w2239, w2240, w2241, w2242, w2243, w2244, w2245, w2246, w2247, w2248, w2249, w2250, w2251, w2252, w2253, w2254, w2255, w2256, w2257, w2258, w2259, w2260, w2261, w2262, w2263, w2264, w2265, w2266, w2267, w2268, w2269, w2270, w2271, w2272, w2273, w2274, w2275, w2276, w2277, w2278, w2279, w2280, w2281, w2282, w2283, w2284, w2285, w2286, w2287, w2288, w2289, w2290, w2291, w2292, w2293, w2294, w2295, w2296, w2297, w2298, w2299, w2300, w2301, w2302, w2303, w2304, w2305, w2306, w2307, w2308, w2309, w2310, w2311, w2312, w2313, w2314, w2315, w2316, w2317, w2318, w2319, w2320, w2321, w2322, w2323, w2324, w2325, w2326, w2327, w2328, w2329, w2330, w2331, w2332, w2333, w2334, w2335, w2336, w2337, w2338, w2339, w2340, w2341, w2342, w2343, w2344, w2345, w2346, w2347, w2348, w2349, w2350, w2351, w2352, w2353, w2354, w2355, w2356, w2357, w2358, w2359, w2360, w2361, w2362, w2363, w2364, w2365, w2366, w2367, w2368, w2369, w2370, w2371, w2372, w2373, w2374, w2375, w2376, w2377, w2378, w2379, w2380, w2381, w2382, w2383, w2384, w2385, w2386, w2387, w2388, w2389, w2390, w2391, w2392, w2393, w2394, w2395, w2396, w2397, w2398, w2399, w2400, w2401, w2402, w2403, w2404, w2405, w2406, w2407, w2408, w2409, w2410, w2411, w2412, w2413, w2414, w2415, w2416, w2417, w2418, w2419, w2420, w2421, w2422, w2423, w2424, w2425, w2426, w2427, w2428, w2429, w2430, w2431, w2432, w2433, w2434, w2435, w2436, w2437, w2438, w2439, w2440, w2441, w2442, w2443, w2444, w2445, w2446, w2447, w2448, w2449, w2450, w2451, w2452, w2453, w2454, w2455, w2456, w2457, w2458, w2459, w2460, w2461, w2462, w2463, w2464, w2465, w2466, w2467, w2468, w2469, w2470, w2471, w2472, w2473, w2474, w2475, w2476, w2477, w2478, w2479, w2480, w2481, w2482, w2483, w2484, w2485, w2486, w2487, w2488, w2489, w2490, w2491, w2492, w2493, w2494, w2495, w2496, w2497, w2498, w2499, w2500, w2501, w2502, w2503, w2504, w2505, w2506, w2507, w2508, w2509, w2510, w2511, w2512, w2513, w2514, w2515, w2516, w2517, w2518, w2519, w2520, w2521, w2522, w2523, w2524, w2525, w2526, w2527, w2528, w2529, w2530, w2531, w2532, w2533, w2534, w2535, w2536, w2537, w2538, w2539, w2540, w2541, w2542, w2543, w2544, w2545, w2546, w2547, w2548, w2549, w2550, w2551, w2552, w2553, w2554, w2555, w2556, w2557, w2558, w2559, w2560, w2561, w2562, w2563, w2564, w2565, w2566, w2567, w2568, w2569, w2570, w2571, w2572, w2573, w2574, w2575, w2576, w2577, w2578, w2579, w2580, w2581, w2582, w2583, w2584, w2585, w2586, w2587, w2588, w2589, w2590, w2591, w2592, w2593, w2594, w2595, w2596, w2597, w2598, w2599, w2600, w2601, w2602, w2603, w2604, w2605, w2606, w2607, w2608, w2609, w2610, w2611, w2612, w2613, w2614, w2615, w2616, w2617, w2618, w2619, w2620, w2621, w2622, w2623, w2624, w2625, w2626, w2627, w2628, w2629, w2630, w2631, w2632, w2633, w2634, w2635, w2636, w2637, w2638, w2639, w2640, w2641, w2642, w2643, w2644, w2645, w2646, w2647, w2648, w2649, w2650, w2651, w2652, w2653, w2654, w2655, w2656, w2657, w2658, w2659, w2660, w2661, w2662, w2663, w2664, w2665, w2666, w2667, w2668, w2669, w2670, w2671, w2672, w2673, w2674, w2675, w2676, w2677, w2678, w2679, w2680, w2681, w2682, w2683, w2684, w2685, w2686, w2687, w2688, w2689, w2690, w2691, w2692, w2693, w2694, w2695, w2696, w2697, w2698, w2699, w2700, w2701, w2702, w2703, w2704, w2705, w2706, w2707, w2708, w2709, w2710, w2711, w2712, w2713, w2714, w2715, w2716, w2717, w2718, w2719, w2720, w2721, w2722, w2723, w2724, w2725, w2726, w2727, w2728, w2729, w2730, w2731, w2732, w2733, w2734, w2735, w2736, w2737, w2738, w2739, w2740, w2741, w2742, w2743, w2744, w2745, w2746, w2747, w2748, w2749, w2750, w2751, w2752, w2753, w2754, w2755, w2756, w2757, w2758, w2759, w2760, w2761, w2762, w2763, w2764, w2765, w2766, w2767, w2768, w2769, w2770, w2771, w2772, w2773, w2774, w2775, w2776, w2777, w2778, w2779, w2780, w2781, w2782, w2783, w2784, w2785, w2786, w2787, w2788, w2789, w2790, w2791, w2792, w2793, w2794, w2795, w2796, w2797, w2798, w2799, w2800, w2801, w2802, w2803, w2804, w2805, w2806, w2807, w2808, w2809, w2810, w2811, w2812, w2813, w2814, w2815, w2816, w2817, w2818, w2819, w2820, w2821, w2822, w2823, w2824, w2825, w2826, w2827, w2828, w2829, w2830, w2831, w2832, w2833, w2834, w2835, w2836, w2837, w2838, w2839, w2840, w2841, w2842, w2843, w2844, w2845, w2846, w2847, w2848, w2849, w2850, w2851, w2852, w2853, w2854, w2855, w2856, w2857, w2858, w2859, w2860, w2861, w2862, w2863, w2864, w2865, w2866, w2867, w2868, w2869, w2870, w2871, w2872, w2873, w2874, w2875, w2876, w2877, w2878, w2879, w2880, w2881, w2882, w2883, w2884, w2885, w2886, w2887, w2888, w2889, w2890, w2891, w2892, w2893, w2894, w2895, w2896, w2897, w2898, w2899, w2900, w2901, w2902, w2903, w2904, w2905, w2906, w2907, w2908, w2909, w2910, w2911, w2912, w2913, w2914, w2915, w2916, w2917, w2918, w2919, w2920, w2921, w2922, w2923, w2924, w2925, w2926, w2927, w2928, w2929, w2930, w2931, w2932, w2933, w2934, w2935, w2936, w2937, w2938, w2939, w2940, w2941, w2942, w2943, w2944, w2945, w2946, w2947, w2948, w2949, w2950, w2951, w2952, w2953, w2954, w2955, w2956, w2957, w2958, w2959, w2960, w2961, w2962, w2963, w2964, w2965, w2966, w2967, w2968, w2969, w2970, w2971, w2972, w2973, w2974, w2975, w2976, w2977, w2978, w2979, w2980, w2981, w2982, w2983, w2984, w2985, w2986, w2987, w2988, w2989, w2990, w2991, w2992, w2993, w2994, w2995, w2996, w2997, w2998, w2999, w3000, w3001, w3002, w3003, w3004, w3005, w3006, w3007, w3008, w3009, w3010, w3011, w3012, w3013, w3014, w3015, w3016, w3017, w3018, w3019, w3020, w3021, w3022, w3023, w3024, w3025, w3026, w3027, w3028, w3029, w3030, w3031, w3032, w3033, w3034, w3035, w3036, w3037, w3038, w3039, w3040, w3041, w3042, w3043, w3044, w3045, w3046, w3047, w3048, w3049, w3050, w3051, w3052, w3053, w3054, w3055, w3056, w3057, w3058, w3059, w3060, w3061, w3062, w3063, w3064, w3065, w3066, w3067, w3068, w3069, w3070, w3071, w3072, w3073, w3074, w3075, w3076, w3077, w3078, w3079, w3080, w3081, w3082, w3083, w3084, w3085, w3086, w3087, w3088, w3089, w3090, w3091, w3092, w3093, w3094, w3095, w3096, w3097, w3098, w3099, w3100, w3101, w3102, w3103, w3104, w3105, w3106, w3107, w3108, w3109, w3110, w3111, w3112, w3113, w3114, w3115, w3116, w3117, w3118, w3119, w3120, w3121, w3122, w3123, w3124, w3125, w3126, w3127, w3128, w3129, w3130, w3131, w3132, w3133, w3134, w3135, w3136, w3137, w3138, w3139, w3140, w3141, w3142, w3143, w3144, w3145, w3146, w3147, w3148, w3149, w3150, w3151, w3152, w3153, w3154, w3155, w3156, w3157, w3158, w3159, w3160, w3161, w3162, w3163, w3164, w3165, w3166, w3167, w3168, w3169, w3170, w3171, w3172, w3173, w3174, w3175, w3176, w3177, w3178, w3179, w3180, w3181, w3182, w3183, w3184, w3185, w3186, w3187, w3188, w3189, w3190, w3191, w3192, w3193, w3194, w3195, w3196, w3197, w3198, w3199, w3200, w3201, w3202, w3203, w3204, w3205, w3206, w3207, w3208, w3209, w3210, w3211, w3212, w3213, w3214, w3215, w3216, w3217, w3218, w3219, w3220, w3221, w3222, w3223, w3224, w3225, w3226, w3227, w3228, w3229, w3230, w3231, w3232, w3233, w3234, w3235, w3236, w3237, w3238, w3239, w3240, w3241, w3242, w3243, w3244, w3245, w3246, w3247, w3248, w3249, w3250, w3251, w3252, w3253, w3254, w3255, w3256, w3257, w3258, w3259, w3260, w3261, w3262, w3263, w3264, w3265, w3266, w3267, w3268, w3269, w3270, w3271, w3272, w3273, w3274, w3275, w3276, w3277, w3278, w3279, w3280, w3281, w3282, w3283, w3284, w3285, w3286, w3287, w3288, w3289, w3290, w3291, w3292, w3293, w3294, w3295, w3296, w3297, w3298, w3299, w3300, w3301, w3302, w3303, w3304, w3305, w3306, w3307, w3308, w3309, w3310, w3311, w3312, w3313, w3314, w3315, w3316, w3317, w3318, w3319, w3320, w3321, w3322, w3323, w3324, w3325, w3326, w3327, w3328, w3329, w3330, w3331, w3332, w3333, w3334, w3335, w3336, w3337, w3338, w3339, w3340, w3341, w3342, w3343, w3344, w3345, w3346, w3347, w3348, w3349, w3350, w3351, w3352, w3353, w3354, w3355, w3356, w3357, w3358, w3359, w3360, w3361, w3362, w3363, w3364, w3365, w3366, w3367, w3368, w3369, w3370, w3371, w3372, w3373, w3374, w3375, w3376, w3377, w3378, w3379, w3380, w3381, w3382, w3383, w3384, w3385, w3386, w3387, w3388, w3389, w3390, w3391, w3392, w3393, w3394, w3395, w3396, w3397, w3398, w3399, w3400, w3401, w3402, w3403, w3404, w3405, w3406, w3407, w3408, w3409, w3410, w3411, w3412, w3413, w3414, w3415, w3416, w3417, w3418, w3419, w3420, w3421, w3422, w3423, w3424, w3425, w3426, w3427, w3428, w3429, w3430, w3431, w3432, w3433, w3434, w3435, w3436, w3437, w3438, w3439, w3440, w3441, w3442, w3443, w3444, w3445, w3446, w3447, w3448, w3449, w3450, w3451, w3452, w3453, w3454, w3455, w3456, w3457, w3458, w3459, w3460, w3461, w3462, w3463, w3464, w3465, w3466, w3467, w3468, w3469, w3470, w3471, w3472, w3473, w3474, w3475, w3476, w3477, w3478, w3479, w3480, w3481, w3482, w3483, w3484, w3485, w3486, w3487, w3488, w3489, w3490, w3491, w3492, w3493, w3494, w3495, w3496, w3497, w3498, w3499, w3500, w3501, w3502, w3503, w3504, w3505, w3506, w3507, w3508, w3509, w3510, w3511, w3512, w3513, w3514, w3515, w3516, w3517, w3518, w3519, w3520, w3521, w3522, w3523, w3524, w3525, w3526, w3527, w3528, w3529, w3530, w3531, w3532, w3533, w3534, w3535, w3536, w3537, w3538, w3539, w3540, w3541, w3542, w3543, w3544, w3545, w3546, w3547, w3548, w3549, w3550, w3551, w3552, w3553, w3554, w3555, w3556, w3557, w3558, w3559, w3560, w3561, w3562, w3563, w3564, w3565, w3566, w3567, w3568, w3569, w3570, w3571, w3572, w3573, w3574, w3575, w3576, w3577, w3578, w3579, w3580, w3581, w3582, w3583, w3584, w3585, w3586, w3587, w3588, w3589, w3590, w3591, w3592, w3593, w3594, w3595, w3596, w3597, w3598, w3599, w3600, w3601, w3602, w3603, w3604, w3605, w3606, w3607, w3608, w3609, w3610, w3611, w3612, w3613, w3614, w3615, w3616, w3617, w3618, w3619, w3620, w3621, w3622, w3623, w3624, w3625, w3626, w3627, w3628, w3629, w3630, w3631, w3632, w3633, w3634, w3635, w3636, w3637, w3638, w3639, w3640, w3641, w3642, w3643, w3644, w3645, w3646, w3647, w3648, w3649, w3650, w3651, w3652, w3653, w3654, w3655, w3656, w3657, w3658, w3659, w3660, w3661, w3662, w3663, w3664, w3665, w3666, w3667, w3668, w3669, w3670, w3671, w3672, w3673, w3674, w3675, w3676, w3677, w3678, w3679, w3680, w3681, w3682, w3683, w3684, w3685, w3686, w3687, w3688, w3689, w3690, w3691, w3692, w3693, w3694, w3695, w3696, w3697, w3698, w3699, w3700, w3701, w3702, w3703, w3704, w3705, w3706, w3707, w3708, w3709, w3710, w3711, w3712, w3713, w3714, w3715, w3716, w3717, w3718, w3719, w3720, w3721, w3722, w3723, w3724, w3725, w3726, w3727, w3728, w3729, w3730, w3731, w3732, w3733, w3734, w3735, w3736, w3737, w3738, w3739, w3740, w3741, w3742, w3743, w3744, w3745, w3746, w3747, w3748, w3749, w3750, w3751, w3752, w3753, w3754, w3755, w3756, w3757, w3758, w3759, w3760, w3761, w3762, w3763, w3764, w3765, w3766, w3767, w3768, w3769, w3770, w3771, w3772, w3773, w3774, w3775, w3776, w3777, w3778, w3779, w3780, w3781, w3782, w3783, w3784, w3785, w3786, w3787, w3788, w3789, w3790, w3791, w3792, w3793, w3794, w3795, w3796, w3797, w3798, w3799, w3800, w3801, w3802, w3803, w3804, w3805, w3806, w3807, w3808, w3809, w3810, w3811, w3812, w3813, w3814, w3815, w3816, w3817, w3818, w3819, w3820, w3821, w3822, w3823, w3824, w3825, w3826, w3827, w3828, w3829, w3830, w3831, w3832, w3833, w3834, w3835, w3836, w3837, w3838, w3839, w3840, w3841, w3842, w3843, w3844, w3845, w3846, w3847, w3848, w3849, w3850, w3851, w3852, w3853, w3854, w3855, w3856, w3857, w3858, w3859, w3860, w3861, w3862, w3863, w3864, w3865, w3866, w3867, w3868, w3869, w3870, w3871, w3872, w3873, w3874, w3875, w3876, w3877, w3878, w3879, w3880, w3881, w3882, w3883, w3884, w3885, w3886, w3887, w3888, w3889, w3890, w3891, w3892, w3893, w3894, w3895, w3896, w3897, w3898, w3899, w3900, w3901, w3902, w3903, w3904, w3905, w3906, w3907, w3908, w3909, w3910, w3911, w3912, w3913, w3914, w3915, w3916, w3917, w3918, w3919, w3920, w3921, w3922, w3923, w3924, w3925, w3926, w3927, w3928, w3929, w3930, w3931, w3932, w3933, w3934, w3935, w3936, w3937, w3938, w3939, w3940, w3941, w3942, w3943, w3944, w3945, w3946, w3947, w3948, w3949, w3950, w3951, w3952, w3953, w3954, w3955, w3956, w3957, w3958, w3959, w3960, w3961, w3962, w3963, w3964, w3965, w3966, w3967, w3968, w3969, w3970, w3971, w3972, w3973, w3974, w3975, w3976, w3977, w3978, w3979, w3980, w3981, w3982, w3983, w3984, w3985, w3986, w3987, w3988, w3989, w3990, w3991, w3992, w3993, w3994, w3995, w3996, w3997, w3998, w3999, w4000, w4001, w4002, w4003, w4004, w4005, w4006, w4007, w4008, w4009, w4010, w4011, w4012, w4013, w4014, w4015, w4016, w4017, w4018, w4019, w4020, w4021, w4022, w4023, w4024, w4025, w4026, w4027, w4028, w4029, w4030, w4031, w4032, w4033, w4034, w4035, w4036, w4037, w4038, w4039, w4040, w4041, w4042, w4043, w4044, w4045, w4046, w4047, w4048, w4049, w4050, w4051, w4052, w4053, w4054, w4055, w4056, w4057, w4058, w4059, w4060, w4061, w4062, w4063, w4064, w4065, w4066, w4067, w4068, w4069, w4070, w4071, w4072, w4073, w4074, w4075, w4076, w4077, w4078, w4079, w4080, w4081, w4082, w4083, w4084, w4085, w4086, w4087, w4088, w4089, w4090, w4091, w4092, w4093, w4094, w4095, w4096, w4097, w4098, w4099, w4100, w4101, w4102, w4103, w4104, w4105, w4106, w4107, w4108, w4109, w4110, w4111, w4112, w4113, w4114, w4115, w4116, w4117, w4118, w4119, w4120, w4121, w4122, w4123, w4124, w4125, w4126, w4127, w4128, w4129, w4130, w4131, w4132, w4133, w4134, w4135, w4136, w4137, w4138, w4139, w4140, w4141, w4142, w4143, w4144, w4145, w4146, w4147, w4148, w4149, w4150, w4151, w4152, w4153, w4154, w4155, w4156, w4157, w4158, w4159, w4160, w4161, w4162, w4163, w4164, w4165, w4166, w4167, w4168, w4169, w4170, w4171, w4172, w4173, w4174, w4175, w4176, w4177, w4178, w4179, w4180, w4181, w4182, w4183, w4184, w4185, w4186, w4187, w4188, w4189, w4190, w4191, w4192, w4193, w4194, w4195, w4196, w4197, w4198, w4199, w4200, w4201, w4202, w4203, w4204, w4205, w4206, w4207, w4208, w4209, w4210, w4211, w4212, w4213, w4214, w4215, w4216, w4217, w4218, w4219, w4220, w4221, w4222, w4223, w4224, w4225, w4226, w4227, w4228, w4229, w4230, w4231, w4232, w4233, w4234, w4235, w4236, w4237, w4238, w4239, w4240, w4241, w4242, w4243, w4244, w4245, w4246, w4247, w4248, w4249, w4250, w4251, w4252, w4253, w4254, w4255, w4256, w4257, w4258, w4259, w4260, w4261, w4262, w4263, w4264, w4265, w4266, w4267, w4268, w4269, w4270, w4271, w4272, w4273, w4274, w4275, w4276, w4277, w4278, w4279, w4280, w4281, w4282, w4283, w4284, w4285, w4286, w4287, w4288, w4289, w4290, w4291, w4292, w4293, w4294, w4295, w4296, w4297, w4298, w4299, w4300, w4301, w4302, w4303, w4304, w4305, w4306, w4307, w4308, w4309, w4310, w4311, w4312, w4313, w4314, w4315, w4316, w4317, w4318, w4319, w4320, w4321, w4322, w4323, w4324, w4325, w4326, w4327, w4328, w4329, w4330, w4331, w4332, w4333, w4334, w4335, w4336, w4337, w4338, w4339, w4340, w4341, w4342, w4343, w4344, w4345, w4346, w4347, w4348, w4349, w4350, w4351, w4352, w4353, w4354, w4355, w4356, w4357, w4358, w4359, w4360, w4361, w4362, w4363, w4364, w4365, w4366, w4367, w4368, w4369, w4370, w4371, w4372, w4373;
assign w0 = pi01 & ~pi02;
assign v0 = ~(pi03 | w0);
assign w1 = v0;
assign w2 = pi01 & pi03;
assign w3 = ~pi14 & w2;
assign w4 = pi01 & ~pi26;
assign v1 = ~(pi03 | w4);
assign w5 = v1;
assign w6 = pi01 & ~pi11;
assign w7 = pi03 & ~pi30;
assign w8 = ~pi13 & w6;
assign w9 = (pi28 & ~w8) | (pi28 & w2106) | (~w8 & w2106);
assign v2 = ~(w5 | w9);
assign w10 = v2;
assign w11 = pi03 & w4;
assign v3 = ~(pi07 | pi09);
assign w12 = v3;
assign w13 = w6 & w12;
assign v4 = ~(pi29 | pi31);
assign w14 = v4;
assign v5 = ~(pi25 | pi27);
assign w15 = v5;
assign v6 = ~(pi21 | pi23);
assign w16 = v6;
assign v7 = ~(pi13 | pi15);
assign w17 = v7;
assign v8 = ~(pi17 | pi19);
assign w18 = v8;
assign w19 = w17 & w18;
assign w20 = ~pi05 & w19;
assign w21 = w3796 & w20;
assign w22 = ~w11 & w13;
assign w23 = w21 & w22;
assign w24 = ~w10 & w23;
assign v9 = ~(pi05 | pi07);
assign w25 = v9;
assign v10 = ~(pi01 | pi03);
assign w26 = v10;
assign w27 = ~pi28 & w2;
assign v11 = ~(pi09 | pi11);
assign w28 = v11;
assign w29 = w25 & ~w26;
assign w30 = w28 & w29;
assign w31 = ~w27 & w30;
assign w32 = w3796 & w19;
assign w33 = w31 & w32;
assign w34 = (pi28 & ~w4) | (pi28 & w2107) | (~w4 & w2107);
assign w35 = (pi05 & w4) | (pi05 & w2108) | (w4 & w2108);
assign w36 = ~w34 & w35;
assign w37 = w3062 & w19;
assign w38 = pi30 & w16;
assign w39 = w13 & w38;
assign w40 = w37 & w39;
assign w41 = ~w36 & w40;
assign w42 = ~w33 & w41;
assign w43 = pi26 & ~w42;
assign w44 = ~pi26 & w42;
assign v12 = ~(w43 | w44);
assign w45 = v12;
assign v13 = ~(w24 | w45);
assign w46 = v13;
assign w47 = ~pi24 & w2;
assign w48 = pi01 & ~pi24;
assign v14 = ~(pi03 | w48);
assign w49 = v14;
assign v15 = ~(w47 | w49);
assign w50 = v15;
assign w51 = ~pi11 & w19;
assign w52 = w12 & w2721;
assign w53 = (pi28 & ~w2) | (pi28 & w2920) | (~w2 & w2920);
assign w54 = pi05 & ~w53;
assign w55 = pi03 & ~pi07;
assign w56 = ~w4 & w55;
assign w57 = w28 & w56;
assign v16 = ~(w13 | w57);
assign w58 = v16;
assign w59 = w3796 & w2757;
assign w60 = (pi30 & w4) | (pi30 & w2758) | (w4 & w2758);
assign w61 = w34 & w60;
assign w62 = ~w58 & w61;
assign w63 = w59 & w62;
assign w64 = (~w54 & ~w62) | (~w54 & w2852) | (~w62 & w2852);
assign w65 = w52 & w64;
assign w66 = (~pi05 & ~w4) | (~pi05 & w2101) | (~w4 & w2101);
assign w67 = (w66 & w9) | (w66 & w2921) | (w9 & w2921);
assign w68 = w2721 & w2109;
assign w69 = ~w67 & w68;
assign w70 = w37 & w38;
assign w71 = ~w31 & w70;
assign w72 = ~w69 & w2359;
assign w73 = ~w48 & w2107;
assign w74 = pi05 & pi07;
assign w75 = ~w73 & w74;
assign w76 = (w75 & w42) | (w75 & w2360) | (w42 & w2360);
assign w77 = w72 & ~w76;
assign w78 = (w50 & w77) | (w50 & w2922) | (w77 & w2922);
assign w79 = w46 & ~w78;
assign w80 = (~w47 & ~w23) | (~w47 & w2111) | (~w23 & w2111);
assign w81 = w43 & w80;
assign w82 = (~pi26 & ~w2) | (~pi26 & w2923) | (~w2 & w2923);
assign w83 = (~w49 & ~w42) | (~w49 & w2112) | (~w42 & w2112);
assign w84 = ~w81 & w83;
assign w85 = (pi28 & ~w21) | (pi28 & w2113) | (~w21 & w2113);
assign w86 = ~w36 & w57;
assign w87 = w71 & w86;
assign v17 = ~(w85 | w87);
assign w88 = v17;
assign v18 = ~(w63 | w88);
assign w89 = v18;
assign w90 = w9 & w57;
assign w91 = w21 & w90;
assign w92 = ~w88 & w2114;
assign w93 = w84 & ~w92;
assign w94 = pi05 & ~w73;
assign w95 = (~w94 & ~w62) | (~w94 & w2924) | (~w62 & w2924);
assign w96 = (w65 & ~w45) | (w65 & w2853) | (~w45 & w2853);
assign w97 = ~w93 & w96;
assign w98 = pi07 & ~pi28;
assign w99 = ~w49 & w98;
assign w100 = (w99 & ~w43) | (w99 & w2115) | (~w43 & w2115);
assign w101 = w77 & ~w100;
assign w102 = (~w101 & w93) | (~w101 & w2854) | (w93 & w2854);
assign w103 = (w50 & w45) | (w50 & w2361) | (w45 & w2361);
assign w104 = (~w97 & w4098) | (~w97 & w4099) | (w4098 & w4099);
assign w105 = w3796 & w3773;
assign w106 = w64 & w105;
assign w107 = (w106 & ~w45) | (w106 & w2855) | (~w45 & w2855);
assign w108 = ~w93 & w107;
assign w109 = w3062 & w2925;
assign w110 = ~pi17 & w109;
assign w111 = pi01 & ~pi13;
assign w112 = pi30 & w28;
assign w113 = (w112 & ~w30) | (w112 & w2927) | (~w30 & w2927);
assign w114 = (w113 & ~w68) | (w113 & w2928) | (~w68 & w2928);
assign w115 = w3701 & w114;
assign w116 = ~w100 & w115;
assign w117 = ~w100 & w2929;
assign w118 = (~w117 & w93) | (~w117 & w2930) | (w93 & w2930);
assign w119 = ~pi22 & w2;
assign w120 = pi01 & ~pi22;
assign v19 = ~(pi03 | w120);
assign w121 = v19;
assign w122 = (~pi24 & w120) | (~pi24 & w2931) | (w120 & w2931);
assign v20 = ~(w119 | w122);
assign w123 = v20;
assign w124 = ~pi05 & w123;
assign w125 = (w2117 & w93) | (w2117 & w4039) | (w93 & w4039);
assign w126 = (pi24 & w120) | (pi24 & w2932) | (w120 & w2932);
assign v21 = ~(w119 | w126);
assign w127 = v21;
assign w128 = ~pi05 & w127;
assign w129 = (~w93 & w4100) | (~w93 & w4101) | (w4100 & w4101);
assign v22 = ~(w125 | w129);
assign w130 = v22;
assign w131 = w104 & w130;
assign w132 = (~pi05 & w81) | (~pi05 & w2119) | (w81 & w2119);
assign w133 = w92 & w132;
assign w134 = w101 & ~w133;
assign w135 = ~pi07 & w92;
assign w136 = (w135 & ~w96) | (w135 & w2120) | (~w96 & w2120);
assign w137 = ~w134 & w136;
assign w138 = (w94 & w42) | (w94 & w2759) | (w42 & w2759);
assign w139 = (~pi07 & w138) | (~pi07 & w2933) | (w138 & w2933);
assign w140 = (w139 & ~w84) | (w139 & w2934) | (~w84 & w2934);
assign w141 = ~w102 & w140;
assign v23 = ~(w137 | w141);
assign w142 = v23;
assign w143 = pi07 & pi30;
assign w144 = (w132 & w3774) | (w132 & w3775) | (w3774 & w3775);
assign w145 = pi30 & ~w33;
assign w146 = ~w69 & w145;
assign w147 = (w2721 & w146) | (w2721 & w3751) | (w146 & w3751);
assign w148 = (w133 & w2856) | (w133 & w2857) | (w2856 & w2857);
assign w149 = ~w141 & w2761;
assign w150 = ~w131 & w149;
assign w151 = ~w138 & w2858;
assign v24 = ~(w76 | w100);
assign w152 = v24;
assign w153 = (w152 & w93) | (w152 & w2762) | (w93 & w2762);
assign w154 = w72 & ~w153;
assign w155 = ~w141 & w2763;
assign w156 = (w141 & w2764) | (w141 & w2765) | (w2764 & w2765);
assign w157 = (w127 & w108) | (w127 & w2362) | (w108 & w2362);
assign w158 = (pi05 & w2363) | (pi05 & w108) | (w2363 & w108);
assign w159 = ~w157 & w158;
assign w160 = w130 & ~w159;
assign w161 = (w160 & w150) | (w160 & w2122) | (w150 & w2122);
assign v25 = ~(w104 | w161);
assign w162 = v25;
assign w163 = w131 & ~w159;
assign w164 = (pi07 & ~w163) | (pi07 & w2859) | (~w163 & w2859);
assign w165 = (w164 & w161) | (w164 & w4040) | (w161 & w4040);
assign w166 = (~w156 & ~w173) | (~w156 & w2766) | (~w173 & w2766);
assign w167 = w131 & w2936;
assign w168 = ~w166 & w167;
assign v26 = ~(pi07 | w104);
assign w169 = v26;
assign w170 = ~w161 & w169;
assign v27 = ~(w168 | w170);
assign w171 = v27;
assign w172 = ~w165 & w171;
assign v28 = ~(w131 | w159);
assign w173 = v28;
assign v29 = ~(w119 | w121);
assign w174 = v29;
assign w175 = (w146 & w2937) | (w146 & w2938) | (w2937 & w2938);
assign w176 = (w133 & w2939) | (w133 & w2940) | (w2939 & w2940);
assign w177 = ~w141 & w2767;
assign w178 = w173 & w177;
assign w179 = (w175 & ~w142) | (w175 & w2123) | (~w142 & w2123);
assign w180 = pi05 & ~pi24;
assign w181 = ~pi05 & pi24;
assign v30 = ~(w180 | w181);
assign w182 = v30;
assign w183 = ~w108 & w2860;
assign w184 = (~w182 & w108) | (~w182 & w2861) | (w108 & w2861);
assign v31 = ~(w183 | w184);
assign w185 = v31;
assign v32 = ~(w179 | w185);
assign w186 = v32;
assign w187 = ~w178 & w186;
assign w188 = w177 & w185;
assign w189 = w173 & w188;
assign w190 = w179 & w185;
assign v33 = ~(w189 | w190);
assign w191 = v33;
assign w192 = ~w187 & w191;
assign w193 = ~pi20 & w2;
assign w194 = (w146 & w2941) | (w146 & w2942) | (w2941 & w2942);
assign w195 = w2124 & w2862;
assign w196 = pi01 & ~pi20;
assign v34 = ~(pi03 | w196);
assign w197 = v34;
assign w198 = (~pi22 & w196) | (~pi22 & w2943) | (w196 & w2943);
assign v35 = ~(w193 | w198);
assign w199 = v35;
assign w200 = (w142 & w2768) | (w142 & w2769) | (w2768 & w2769);
assign w201 = (w200 & ~w173) | (w200 & w2944) | (~w173 & w2944);
assign w202 = (w146 & w2945) | (w146 & w2946) | (w2945 & w2946);
assign w203 = (w202 & ~w2763) | (w202 & w2947) | (~w2763 & w2947);
assign w204 = w2124 & w2863;
assign w205 = (~w203 & ~w173) | (~w203 & w2948) | (~w173 & w2948);
assign w206 = ~w201 & w205;
assign w207 = ~w192 & w206;
assign v36 = ~(pi24 | w118);
assign w208 = v36;
assign w209 = pi24 & w118;
assign v37 = ~(w208 | w209);
assign w210 = v37;
assign w211 = ~pi05 & w210;
assign w212 = (~w2864 & w4102) | (~w2864 & w4103) | (w4102 & w4103);
assign v38 = ~(pi05 | w210);
assign w213 = v38;
assign w214 = ~w178 & w2364;
assign v39 = ~(w212 | w214);
assign w215 = v39;
assign w216 = (w215 & w192) | (w215 & w4104) | (w192 & w4104);
assign w217 = w172 & w216;
assign w218 = ~w153 & w3776;
assign w219 = (~w2365 & w4105) | (~w2365 & w4106) | (w4105 & w4106);
assign v40 = ~(w173 | w219);
assign w220 = v40;
assign w221 = (w92 & w102) | (w92 & w133) | (w102 & w133);
assign w222 = w2763 & w3777;
assign w223 = (~w222 & ~w173) | (~w222 & w3778) | (~w173 & w3778);
assign w224 = (pi09 & ~w223) | (pi09 & w2366) | (~w223 & w2366);
assign v41 = ~(w165 | w224);
assign w225 = v41;
assign w226 = ~pi11 & w225;
assign w227 = (w226 & ~w216) | (w226 & w4041) | (~w216 & w4041);
assign w228 = (w173 & w2770) | (w173 & w2771) | (w2770 & w2771);
assign v42 = ~(w166 | w228);
assign w229 = v42;
assign w230 = (w2865 & w166) | (w2865 & w4328) | (w166 & w4328);
assign w231 = w223 & w2866;
assign v43 = ~(w230 | w231);
assign w232 = v43;
assign w233 = (w232 & w217) | (w232 & w2368) | (w217 & w2368);
assign w234 = w223 & w2369;
assign w235 = (pi11 & ~w2369) | (pi11 & w3779) | (~w2369 & w3779);
assign w236 = ~w225 & w235;
assign w237 = (w32 & w225) | (w32 & w2370) | (w225 & w2370);
assign w238 = (pi11 & w178) | (pi11 & w2949) | (w178 & w2949);
assign w239 = w171 & w238;
assign w240 = (~w234 & w192) | (~w234 & w2371) | (w192 & w2371);
assign w241 = w239 & w240;
assign w242 = w237 & ~w241;
assign w243 = ~w233 & w242;
assign w244 = (w2950 & w161) | (w2950 & w4107) | (w161 & w4107);
assign w245 = (~w244 & w233) | (~w244 & w2125) | (w233 & w2125);
assign w246 = (~pi09 & w2951) | (~pi09 & w162) | (w2951 & w162);
assign w247 = w245 & ~w246;
assign v44 = ~(w172 | w216);
assign w248 = v44;
assign v45 = ~(w217 | w248);
assign w249 = v45;
assign w250 = pi09 & w249;
assign w251 = w243 & ~w250;
assign v46 = ~(pi09 | w249);
assign w252 = v46;
assign w253 = w243 & w2126;
assign v47 = ~(w247 | w253);
assign w254 = v47;
assign w255 = ~w210 & w4341;
assign w256 = ~w179 & w4342;
assign v48 = ~(w255 | w256);
assign w257 = v48;
assign w258 = ~w243 & w257;
assign w259 = w192 & ~w206;
assign v49 = ~(w207 | w259);
assign w260 = v49;
assign w261 = w243 & w260;
assign v50 = ~(w258 | w261);
assign w262 = v50;
assign v51 = ~(w193 | w197);
assign w263 = v51;
assign w264 = (w263 & ~w240) | (w263 & w2127) | (~w240 & w2127);
assign w265 = (~w2766 & w4042) | (~w2766 & w4043) | (w4042 & w4043);
assign w266 = (w2772 & w4044) | (w2772 & w4045) | (w4044 & w4045);
assign v52 = ~(w265 | w266);
assign w267 = v52;
assign w268 = pi05 & w267;
assign v53 = ~(pi05 | w267);
assign w269 = v53;
assign v54 = ~(w268 | w269);
assign w270 = v54;
assign w271 = (w270 & w233) | (w270 & w2128) | (w233 & w2128);
assign w272 = ~w233 & w2129;
assign v55 = ~(w271 | w272);
assign w273 = v55;
assign w274 = (w3701 & ~w240) | (w3701 & w2130) | (~w240 & w2130);
assign w275 = ~pi03 & pi18;
assign w276 = ~pi18 & w2;
assign v56 = ~(w26 | w275);
assign w277 = v56;
assign w278 = ~pi20 & w277;
assign v57 = ~(w276 | w278);
assign w279 = v57;
assign w280 = (w279 & w233) | (w279 & w2131) | (w233 & w2131);
assign w281 = (~pi20 & ~w2) | (~pi20 & w2952) | (~w2 & w2952);
assign w282 = w109 & w2953;
assign w283 = (w282 & w225) | (w282 & w2372) | (w225 & w2372);
assign w284 = ~w241 & w283;
assign w285 = ~w233 & w284;
assign v58 = ~(w280 | w285);
assign w286 = v58;
assign w287 = ~w273 & w286;
assign w288 = ~w236 & w264;
assign w289 = ~w233 & w288;
assign w290 = w59 & ~w267;
assign w291 = w289 & w290;
assign w292 = (~w2132 & w2373) | (~w2132 & w2374) | (w2373 & w2374);
assign w293 = ~w291 & w292;
assign w294 = ~w287 & w293;
assign w295 = ~w254 & w262;
assign w296 = ~w294 & w295;
assign w297 = w21 & w267;
assign w298 = ~w233 & w2133;
assign w299 = (w269 & w233) | (w269 & w2134) | (w233 & w2134);
assign w300 = (pi07 & w233) | (pi07 & w2135) | (w233 & w2135);
assign w301 = ~w280 & w300;
assign v59 = ~(w298 | w299);
assign w302 = v59;
assign w303 = w301 & w302;
assign w304 = (~w267 & w233) | (~w267 & w2136) | (w233 & w2136);
assign w305 = ~w233 & w2137;
assign v60 = ~(w304 | w305);
assign w306 = v60;
assign w307 = w74 & w306;
assign v61 = ~(w303 | w307);
assign w308 = v61;
assign v62 = ~(w254 | w308);
assign w309 = v62;
assign v63 = ~(w296 | w309);
assign w310 = v63;
assign v64 = ~(w224 | w234);
assign w311 = v64;
assign w312 = w216 & w2375;
assign w313 = w165 & ~w311;
assign w314 = ~w165 & w311;
assign w315 = ~w217 & w2138;
assign v65 = ~(w312 | w315);
assign w316 = v65;
assign w317 = (w4041 & w4109) | (w4041 & w4110) | (w4109 & w4110);
assign w318 = ~w316 & w317;
assign w319 = w223 & w2954;
assign w320 = (w319 & w233) | (w319 & w2140) | (w233 & w2140);
assign v66 = ~(w318 | w320);
assign w321 = v66;
assign v67 = ~(w245 | w251);
assign w322 = v67;
assign w323 = w321 & w322;
assign w324 = (~w229 & w3605) | (~w229 & w2955) | (w3605 & w2955);
assign w325 = (pi11 & ~w223) | (pi11 & w4111) | (~w223 & w4111);
assign w326 = (w325 & w233) | (w325 & w2141) | (w233 & w2141);
assign w327 = (w2956 & w166) | (w2956 & w4329) | (w166 & w4329);
assign w328 = ~w241 & w2868;
assign w329 = ~w315 & w328;
assign v68 = ~(w326 | w329);
assign w330 = v68;
assign w331 = w324 & w330;
assign w332 = ~w323 & w331;
assign w333 = (~w231 & w225) | (~w231 & w3780) | (w225 & w3780);
assign w334 = ~w241 & w333;
assign w335 = ~w227 & w334;
assign w336 = ~w229 & w2957;
assign w337 = ~w335 & w336;
assign w338 = (~w337 & w323) | (~w337 & w2142) | (w323 & w2142);
assign w339 = ~w296 & w2619;
assign w340 = (~w2376 & w2773) | (~w2376 & w2774) | (w2773 & w2774);
assign w341 = (w340 & ~w310) | (w340 & w2143) | (~w310 & w2143);
assign w342 = pi01 & ~pi16;
assign v69 = ~(w2 | w342);
assign w343 = v69;
assign w344 = pi18 & ~w343;
assign w345 = (w310 & w2377) | (w310 & w2378) | (w2377 & w2378);
assign v70 = ~(pi03 | w342);
assign w346 = v70;
assign w347 = (~pi18 & w342) | (~pi18 & w2958) | (w342 & w2958);
assign w348 = ~pi16 & w2;
assign w349 = ~pi01 & w347;
assign v71 = ~(w348 | w349);
assign w350 = v71;
assign w351 = (w310 & w2379) | (w310 & w2380) | (w2379 & w2380);
assign w352 = ~w345 & w351;
assign w353 = ~w276 & w277;
assign w354 = (~w2774 & w2871) | (~w2774 & w2872) | (w2871 & w2872);
assign w355 = (~w323 & w2873) | (~w323 & w2874) | (w2873 & w2874);
assign w356 = ~w296 & w2959;
assign w357 = ~w236 & w274;
assign w358 = (pi20 & w233) | (pi20 & w4046) | (w233 & w4046);
assign w359 = ~w233 & w4047;
assign v72 = ~(w358 | w359);
assign w360 = v72;
assign w361 = (pi05 & w358) | (pi05 & w4330) | (w358 & w4330);
assign w362 = ~w358 & w4331;
assign v73 = ~(w361 | w362);
assign w363 = v73;
assign w364 = (w2144 & ~w310) | (w2144 & w2381) | (~w310 & w2381);
assign w365 = (w310 & w2382) | (w310 & w2383) | (w2382 & w2383);
assign v74 = ~(w364 | w365);
assign w366 = v74;
assign w367 = ~w352 & w366;
assign w368 = pi05 & w360;
assign w369 = (w2146 & ~w310) | (w2146 & w2384) | (~w310 & w2384);
assign w370 = (w310 & w2385) | (w310 & w2386) | (w2385 & w2386);
assign v75 = ~(w369 | w370);
assign w371 = v75;
assign w372 = w273 & ~w286;
assign v76 = ~(w287 | w372);
assign w373 = v76;
assign v77 = ~(pi07 | w373);
assign w374 = v77;
assign w375 = pi07 & w373;
assign v78 = ~(w374 | w375);
assign w376 = v78;
assign w377 = (w310 & w2620) | (w310 & w2621) | (w2620 & w2621);
assign v79 = ~(pi07 | w306);
assign w378 = v79;
assign w379 = pi07 & w306;
assign v80 = ~(w378 | w379);
assign w380 = v80;
assign w381 = (~w310 & w2387) | (~w310 & w2388) | (w2387 & w2388);
assign v81 = ~(w377 | w381);
assign w382 = v81;
assign w383 = w371 & ~w382;
assign w384 = ~w367 & w383;
assign w385 = ~w296 & w332;
assign w386 = ~w294 & w308;
assign w387 = pi09 & ~w262;
assign w388 = ~pi09 & w262;
assign v82 = ~(w387 | w388);
assign w389 = v82;
assign w390 = (w385 & w2622) | (w385 & w2623) | (w2622 & w2623);
assign w391 = (~w385 & w2624) | (~w385 & w2625) | (w2624 & w2625);
assign v83 = ~(w390 | w391);
assign w392 = v83;
assign w393 = (w310 & w2389) | (w310 & w2390) | (w2389 & w2390);
assign w394 = (~w310 & w2391) | (~w310 & w2392) | (w2391 & w2392);
assign v84 = ~(w393 | w394);
assign w395 = v84;
assign w396 = ~w392 & w395;
assign w397 = (w396 & ~w383) | (w396 & w2798) | (~w383 & w2798);
assign w398 = (~w385 & w2626) | (~w385 & w2627) | (w2626 & w2627);
assign w399 = (w385 & w2628) | (w385 & w2629) | (w2628 & w2629);
assign v85 = ~(w398 | w399);
assign w400 = v85;
assign w401 = pi09 & ~w400;
assign w402 = (w262 & w287) | (w262 & w2875) | (w287 & w2875);
assign w403 = w254 & w308;
assign w404 = ~w402 & w403;
assign w405 = w339 & ~w404;
assign w406 = (~pi09 & w253) | (~pi09 & w2876) | (w253 & w2876);
assign v86 = ~(w322 | w406);
assign w407 = v86;
assign w408 = w340 & ~w407;
assign w409 = ~w339 & w408;
assign v87 = ~(w405 | w409);
assign w410 = v87;
assign w411 = ~pi11 & w410;
assign w412 = pi11 & ~w410;
assign v88 = ~(w411 | w412);
assign w413 = v88;
assign w414 = ~w401 & w413;
assign w415 = (w110 & w146) | (w110 & w2960) | (w146 & w2960);
assign w416 = w321 & w330;
assign w417 = ~w296 & w2630;
assign w418 = (w296 & w2631) | (w296 & w2632) | (w2631 & w2632);
assign v89 = ~(w417 | w418);
assign w419 = v89;
assign v90 = ~(w341 | w419);
assign w420 = v90;
assign w421 = pi11 & w330;
assign w422 = w321 & ~w421;
assign w423 = (~w310 & w2393) | (~w310 & w2394) | (w2393 & w2394);
assign w424 = (w310 & w2877) | (w310 & w2878) | (w2877 & w2878);
assign w425 = ~w420 & w424;
assign w426 = (w415 & w420) | (w415 & w2961) | (w420 & w2961);
assign w427 = w413 & w2962;
assign w428 = ~w397 & w427;
assign w429 = ~w341 & w419;
assign w430 = (w310 & w2879) | (w310 & w2880) | (w2879 & w2880);
assign w431 = ~w429 & w430;
assign w432 = (~w310 & w2397) | (~w310 & w2398) | (w2397 & w2398);
assign w433 = ~w323 & w2633;
assign w434 = (w2399 & w433) | (w2399 & w310) | (w433 & w310);
assign v91 = ~(w432 | w434);
assign w435 = v91;
assign w436 = (w2960 & w432) | (w2960 & w4048) | (w432 & w4048);
assign v92 = ~(w431 | w436);
assign w437 = v92;
assign w438 = w411 & ~w425;
assign w439 = w437 & ~w438;
assign w440 = w415 & ~w439;
assign v93 = ~(w428 | w440);
assign w441 = v93;
assign w442 = ~w428 & w2150;
assign w443 = w427 & w2151;
assign w444 = ~pi01 & pi16;
assign w445 = pi01 & ~pi14;
assign v94 = ~(pi03 | w445);
assign w446 = v94;
assign v95 = ~(w444 | w446);
assign w447 = v95;
assign w448 = (w447 & w439) | (w447 & w2400) | (w439 & w2400);
assign w449 = ~w443 & w448;
assign w450 = ~w442 & w449;
assign v96 = ~(w3 | w450);
assign w451 = v96;
assign v97 = ~(w346 | w348);
assign w452 = v97;
assign w453 = (w452 & w428) | (w452 & w2152) | (w428 & w2152);
assign w454 = (w310 & w3781) | (w310 & w3782) | (w3781 & w3782);
assign w455 = (~w310 & w4112) | (~w310 & w4113) | (w4112 & w4113);
assign v98 = ~(w454 | w455);
assign w456 = v98;
assign w457 = pi05 & ~w456;
assign w458 = ~pi05 & w456;
assign v99 = ~(w457 | w458);
assign w459 = v99;
assign w460 = (w428 & w2401) | (w428 & w2402) | (w2401 & w2402);
assign w461 = (~w428 & w2403) | (~w428 & w2404) | (w2403 & w2404);
assign v100 = ~(w460 | w461);
assign w462 = v100;
assign v101 = ~(w451 | w462);
assign w463 = v101;
assign w464 = (~w360 & w356) | (~w360 & w2634) | (w356 & w2634);
assign w465 = ~w356 & w2635;
assign v102 = ~(w464 | w465);
assign w466 = v102;
assign w467 = ~pi07 & w466;
assign w468 = ~w428 & w2153;
assign w469 = pi07 & ~w466;
assign w470 = ~w428 & w2405;
assign w471 = w352 & ~w366;
assign v103 = ~(w367 | w471);
assign w472 = v103;
assign v104 = ~(pi07 | w472);
assign w473 = v104;
assign w474 = (~w473 & w428) | (~w473 & w2154) | (w428 & w2154);
assign w475 = pi07 & w472;
assign w476 = (w428 & w2775) | (w428 & w2776) | (w2775 & w2776);
assign v105 = ~(w470 | w476);
assign w477 = v105;
assign w478 = (w428 & w2406) | (w428 & w2407) | (w2406 & w2407);
assign w479 = pi05 & w456;
assign w480 = (~w428 & w2408) | (~w428 & w2409) | (w2408 & w2409);
assign v106 = ~(w478 | w480);
assign w481 = v106;
assign w482 = ~w477 & w481;
assign w483 = ~w463 & w482;
assign v107 = ~(w468 | w474);
assign w484 = v107;
assign w485 = w392 & ~w395;
assign v108 = ~(w396 | w485);
assign w486 = v108;
assign w487 = w384 & w486;
assign v109 = ~(w384 | w486);
assign w488 = v109;
assign v110 = ~(w487 | w488);
assign w489 = v110;
assign v111 = ~(pi11 | w489);
assign w490 = v111;
assign w491 = ~w441 & w490;
assign w492 = ~pi11 & w400;
assign w493 = ~w428 & w2155;
assign v112 = ~(w491 | w493);
assign w494 = v112;
assign w495 = (w382 & w367) | (w382 & w2636) | (w367 & w2636);
assign v113 = ~(w384 | w495);
assign w496 = v113;
assign w497 = pi09 & ~w496;
assign w498 = (w497 & w428) | (w497 & w2410) | (w428 & w2410);
assign w499 = (w310 & w2966) | (w310 & w2967) | (w2966 & w2967);
assign w500 = (~w310 & w3439) | (~w310 & w2968) | (w3439 & w2968);
assign v114 = ~(w499 | w500);
assign w501 = v114;
assign w502 = pi09 & w501;
assign w503 = ~w428 & w2156;
assign v115 = ~(w498 | w503);
assign w504 = v115;
assign v116 = ~(pi09 | w501);
assign w505 = v116;
assign w506 = ~w428 & w2157;
assign w507 = ~pi09 & w496;
assign w508 = (w507 & w428) | (w507 & w2411) | (w428 & w2411);
assign v117 = ~(w506 | w508);
assign w509 = v117;
assign w510 = w504 & w509;
assign w511 = ~w484 & w494;
assign w512 = w510 & w511;
assign w513 = ~w483 & w512;
assign w514 = w396 & ~w411;
assign w515 = ~w384 & w514;
assign w516 = (~w411 & ~w413) | (~w411 & w2158) | (~w413 & w2158);
assign v118 = ~(w425 | w431);
assign w517 = v118;
assign w518 = w436 & w517;
assign w519 = (~w518 & w515) | (~w518 & w2799) | (w515 & w2799);
assign v119 = ~(w437 | w517);
assign w520 = v119;
assign w521 = ~w515 & w2800;
assign v120 = ~(w519 | w521);
assign w522 = v120;
assign v121 = ~(w420 | w423);
assign w523 = v121;
assign w524 = ~w428 & w2159;
assign v122 = ~(w522 | w524);
assign w525 = v122;
assign w526 = ~w522 & w2969;
assign w527 = ~w429 & w2970;
assign w528 = (~pi15 & w420) | (~pi15 & w2971) | (w420 & w2971);
assign w529 = (~w527 & w428) | (~w527 & w2160) | (w428 & w2160);
assign w530 = (~pi17 & w432) | (~pi17 & w4114) | (w432 & w4114);
assign w531 = (w530 & ~w529) | (w530 & w2412) | (~w529 & w2412);
assign w532 = (w432 & w4115) | (w432 & w4116) | (w4115 & w4116);
assign w533 = (w532 & ~w526) | (w532 & w2413) | (~w526 & w2413);
assign w534 = pi11 & ~w400;
assign w535 = ~w428 & w2161;
assign w536 = pi11 & w489;
assign w537 = ~w441 & w536;
assign v123 = ~(w535 | w537);
assign w538 = v123;
assign w539 = w504 & w538;
assign w540 = w494 & ~w539;
assign w541 = ~w428 & w2162;
assign w542 = ~w413 & w3757;
assign w543 = ~w397 & w414;
assign w544 = w440 & ~w543;
assign w545 = ~w542 & w544;
assign v124 = ~(w541 | w545);
assign w546 = v124;
assign w547 = (~pi13 & w545) | (~pi13 & w2972) | (w545 & w2972);
assign w548 = ~w545 & w2973;
assign v125 = ~(w547 | w548);
assign w549 = v125;
assign w550 = ~w540 & w549;
assign w551 = ~w540 & w2415;
assign w552 = ~w513 & w551;
assign w553 = (~pi15 & w522) | (~pi15 & w2974) | (w522 & w2974);
assign v126 = ~(w526 | w553);
assign w554 = v126;
assign w555 = ~w547 & w554;
assign w556 = w533 & ~w555;
assign w557 = (~w556 & ~w551) | (~w556 & w2163) | (~w551 & w2163);
assign w558 = w511 & w2416;
assign w559 = ~w483 & w558;
assign w560 = (~w547 & w540) | (~w547 & w2164) | (w540 & w2164);
assign w561 = ~w559 & w2165;
assign v127 = ~(w557 | w561);
assign w562 = v127;
assign w563 = (w110 & w432) | (w110 & w4117) | (w432 & w4117);
assign w564 = (w563 & ~w529) | (w563 & w2417) | (~w529 & w2417);
assign v128 = ~(w547 | w564);
assign w565 = v128;
assign w566 = w554 & w565;
assign w567 = w525 & w566;
assign w568 = (w567 & w559) | (w567 & w2166) | (w559 & w2166);
assign w569 = w525 & ~w533;
assign w570 = (~pi17 & w533) | (~pi17 & w2975) | (w533 & w2975);
assign w571 = (~w2166 & w2418) | (~w2166 & w2419) | (w2418 & w2419);
assign w572 = ~w562 & w571;
assign w573 = ~w559 & w2167;
assign w574 = (~w435 & ~w529) | (~w435 & w2420) | (~w529 & w2420);
assign w575 = (w2977 & w3783) | (w2977 & w3784) | (w3783 & w3784);
assign w576 = pi17 & ~w553;
assign w577 = w575 & w576;
assign w578 = (~w2421 & w2802) | (~w2421 & w2803) | (w2802 & w2803);
assign w579 = (w578 & w562) | (w578 & w4049) | (w562 & w4049);
assign w580 = ~w109 & w4343;
assign w581 = (~w580 & w572) | (~w580 & w2422) | (w572 & w2422);
assign w582 = ~w533 & w2978;
assign w583 = w576 & w3785;
assign w584 = w553 & w575;
assign w585 = (~w584 & ~w566) | (~w584 & w3786) | (~w566 & w3786);
assign w586 = (w559 & w3787) | (w559 & w3788) | (w3787 & w3788);
assign w587 = (w559 & w4050) | (w559 & w4051) | (w4050 & w4051);
assign w588 = ~w586 & w587;
assign w589 = ~w572 & w588;
assign w590 = ~w513 & w550;
assign w591 = w513 & ~w549;
assign v129 = ~(w590 | w591);
assign w592 = v129;
assign w593 = w533 & ~w566;
assign w594 = w540 & ~w549;
assign w595 = w593 & ~w594;
assign w596 = w592 & w595;
assign w597 = (~w546 & w566) | (~w546 & w2979) | (w566 & w2979);
assign w598 = ~w552 & w597;
assign w599 = (pi15 & w552) | (pi15 & w2170) | (w552 & w2170);
assign w600 = ~w596 & w599;
assign w601 = (~w580 & w596) | (~w580 & w2423) | (w596 & w2423);
assign w602 = w589 & w601;
assign v130 = ~(w581 | w602);
assign w603 = v130;
assign w604 = (~w444 & w439) | (~w444 & w2980) | (w439 & w2980);
assign w605 = ~w443 & w604;
assign w606 = ~w442 & w605;
assign w607 = pi05 & w606;
assign w608 = w566 & w607;
assign v131 = ~(w3 | w446);
assign w609 = v131;
assign w610 = w609 & w532;
assign w611 = (w610 & ~w526) | (w610 & w2424) | (~w526 & w2424);
assign w612 = w607 & ~w611;
assign w613 = (~w593 & ~w551) | (~w593 & w2171) | (~w551 & w2171);
assign w614 = pi05 & w609;
assign w615 = ~w606 & w614;
assign w616 = (~w2171 & w2425) | (~w2171 & w2426) | (w2425 & w2426);
assign w617 = (~pi09 & w611) | (~pi09 & w2981) | (w611 & w2981);
assign w618 = (w617 & w590) | (w617 & w2427) | (w590 & w2427);
assign w619 = ~w616 & w618;
assign w620 = (w477 & w463) | (w477 & w2982) | (w463 & w2982);
assign v132 = ~(w483 | w620);
assign w621 = v132;
assign w622 = (~w2171 & w4118) | (~w2171 & w4119) | (w4118 & w4119);
assign w623 = w441 & ~w466;
assign w624 = ~w441 & w472;
assign v133 = ~(w623 | w624);
assign w625 = v133;
assign w626 = (w2171 & w2428) | (w2171 & w2429) | (w2428 & w2429);
assign v134 = ~(w622 | w626);
assign w627 = v134;
assign w628 = ~w619 & w627;
assign w629 = ~pi12 & w2;
assign w630 = w445 & ~w629;
assign w631 = ~pi05 & w609;
assign w632 = (~w630 & ~w606) | (~w630 & w2983) | (~w606 & w2983);
assign w633 = (~w2171 & w2430) | (~w2171 & w2431) | (w2430 & w2431);
assign w634 = (pi14 & ~w2) | (pi14 & w2984) | (~w2 & w2984);
assign w635 = (~w634 & w606) | (~w634 & w2985) | (w606 & w2985);
assign w636 = w566 & ~w635;
assign w637 = pi01 & w533;
assign w638 = (w526 & w3789) | (w526 & w3790) | (w3789 & w3790);
assign w639 = pi01 & ~pi12;
assign v135 = ~(pi03 | w639);
assign w640 = v135;
assign w641 = (~w640 & w611) | (~w640 & w2987) | (w611 & w2987);
assign w642 = ~w638 & w641;
assign w643 = (w642 & w590) | (w642 & w2988) | (w590 & w2988);
assign w644 = ~w633 & w643;
assign w645 = (~w612 & w590) | (~w612 & w2432) | (w590 & w2432);
assign w646 = ~w616 & w645;
assign w647 = ~w644 & w646;
assign w648 = w451 & w462;
assign v136 = ~(w463 | w648);
assign w649 = v136;
assign w650 = (~w2171 & w2433) | (~w2171 & w2434) | (w2433 & w2434);
assign v137 = ~(w453 | w456);
assign w651 = v137;
assign w652 = w453 & w456;
assign v138 = ~(w651 | w652);
assign w653 = v138;
assign w654 = (~w653 & w566) | (~w653 & w2637) | (w566 & w2637);
assign w655 = ~w552 & w654;
assign v139 = ~(w650 | w655);
assign w656 = v139;
assign w657 = pi07 & w656;
assign w658 = w647 & ~w657;
assign w659 = ~w628 & w658;
assign w660 = w12 & ~w656;
assign w661 = pi09 & w566;
assign w662 = (~w526 & w4120) | (~w526 & w4121) | (w4120 & w4121);
assign w663 = (pi09 & w649) | (pi09 & w3791) | (w649 & w3791);
assign w664 = (~w663 & w590) | (~w663 & w4122) | (w590 & w4122);
assign w665 = ~w552 & w2172;
assign v140 = ~(w664 | w665);
assign w666 = v140;
assign v141 = ~(w627 | w666);
assign w667 = v141;
assign w668 = ~w667 & w2435;
assign w669 = ~w659 & w668;
assign w670 = ~w483 & w2436;
assign w671 = w504 & ~w670;
assign w672 = ~w498 & w3792;
assign w673 = (w672 & w483) | (w672 & w2638) | (w483 & w2638);
assign w674 = (~w2171 & w4123) | (~w2171 & w4124) | (w4123 & w4124);
assign v142 = ~(w441 | w489);
assign w675 = v142;
assign w676 = w400 & w441;
assign v143 = ~(w675 | w676);
assign w677 = v143;
assign w678 = pi13 & w677;
assign v144 = ~(pi13 | w677);
assign w679 = v144;
assign v145 = ~(w678 | w679);
assign w680 = v145;
assign w681 = (~w680 & ~w674) | (~w680 & w2437) | (~w674 & w2437);
assign w682 = w674 & w2438;
assign v146 = ~(w681 | w682);
assign w683 = v146;
assign w684 = ~w441 & w496;
assign w685 = w441 & ~w501;
assign v147 = ~(w684 | w685);
assign w686 = v147;
assign w687 = (w2171 & w2989) | (w2171 & w2990) | (w2989 & w2990);
assign w688 = (~w510 & w483) | (~w510 & w2991) | (w483 & w2991);
assign v148 = ~(w670 | w688);
assign w689 = v148;
assign w690 = ~w613 & w689;
assign v149 = ~(w687 | w690);
assign w691 = v149;
assign w692 = w683 & w691;
assign w693 = (w692 & w659) | (w692 & w2439) | (w659 & w2439);
assign v150 = ~(pi11 | w680);
assign w694 = v150;
assign w695 = ~w613 & w2440;
assign w696 = ~pi11 & w680;
assign w697 = (w696 & w613) | (w696 & w2441) | (w613 & w2441);
assign v151 = ~(w695 | w697);
assign w698 = v151;
assign v152 = ~(w628 | w698);
assign w699 = v152;
assign w700 = w658 & w699;
assign w701 = (~w698 & w667) | (~w698 & w2442) | (w667 & w2442);
assign v153 = ~(w700 | w701);
assign w702 = v153;
assign w703 = (w677 & ~w674) | (w677 & w2443) | (~w674 & w2443);
assign v154 = ~(w513 | w540);
assign w704 = v154;
assign w705 = ~w613 & w2444;
assign v155 = ~(pi13 | w705);
assign w706 = v155;
assign w707 = ~w703 & w706;
assign w708 = ~w552 & w2173;
assign w709 = w109 & w4344;
assign w710 = ~w566 & w709;
assign w711 = ~w594 & w710;
assign w712 = w592 & w711;
assign v156 = ~(w708 | w712);
assign w713 = v156;
assign w714 = ~w600 & w713;
assign w715 = ~w707 & w714;
assign w716 = ~w700 & w2445;
assign w717 = ~w693 & w716;
assign w718 = (~w603 & ~w716) | (~w603 & w4125) | (~w716 & w4125);
assign w719 = ~w700 & w2446;
assign w720 = (~w714 & ~w719) | (~w714 & w4126) | (~w719 & w4126);
assign w721 = w718 & ~w720;
assign w722 = w579 & w714;
assign w723 = ~w707 & w722;
assign w724 = w702 & w723;
assign w725 = (~w603 & ~w702) | (~w603 & w742) | (~w702 & w742);
assign w726 = (w692 & w602) | (w692 & w2639) | (w602 & w2639);
assign v157 = ~(w596 | w598);
assign w727 = v157;
assign w728 = (w727 & ~w726) | (w727 & w2993) | (~w726 & w2993);
assign w729 = ~w725 & w728;
assign v158 = ~(w721 | w729);
assign w730 = v158;
assign w731 = (pi17 & w721) | (pi17 & w2174) | (w721 & w2174);
assign w732 = (~pi17 & ~w728) | (~pi17 & w2175) | (~w728 & w2175);
assign w733 = ~w721 & w732;
assign w734 = (~pi11 & w667) | (~pi11 & w2447) | (w667 & w2447);
assign w735 = (w4032 & w691) | (w4032 & w4052) | (w691 & w4052);
assign w736 = ~w669 & w735;
assign w737 = (~pi11 & ~w627) | (~pi11 & w2448) | (~w627 & w2448);
assign w738 = w658 & w737;
assign v159 = ~(w734 | w738);
assign w739 = v159;
assign w740 = ~w738 & w2449;
assign w741 = ~w736 & w740;
assign v160 = ~(w603 | w723);
assign w742 = v160;
assign w743 = w742 & w4127;
assign w744 = ~w741 & w743;
assign v161 = ~(w703 | w705);
assign w745 = v161;
assign w746 = (w745 & w669) | (w745 & w2640) | (w669 & w2640);
assign w747 = ~w725 & w746;
assign v162 = ~(w744 | w747);
assign w748 = v162;
assign w749 = ~w744 & w2641;
assign v163 = ~(w733 | w749);
assign w750 = v163;
assign w751 = ~w731 & w750;
assign w752 = ~w693 & w724;
assign v164 = ~(w603 | w738);
assign w753 = v164;
assign w754 = w736 & w753;
assign w755 = ~w752 & w754;
assign w756 = ~w669 & w739;
assign w757 = (~w691 & ~w756) | (~w691 & w2176) | (~w756 & w2176);
assign v165 = ~(w755 | w757);
assign w758 = v165;
assign w759 = ~w755 & w2177;
assign w760 = (~pi15 & w744) | (~pi15 & w2642) | (w744 & w2642);
assign v166 = ~(w759 | w760);
assign w761 = v166;
assign w762 = w751 & ~w761;
assign w763 = (w742 & w2994) | (w742 & w2995) | (w2994 & w2995);
assign v167 = ~(w718 | w763);
assign w764 = v167;
assign w765 = w589 & ~w600;
assign w766 = ~w589 & w600;
assign w767 = (w716 & w4128) | (w716 & w4129) | (w4128 & w4129);
assign w768 = ~w764 & w767;
assign v168 = ~(w568 | w569);
assign w769 = v168;
assign w770 = ~w562 & w769;
assign w771 = (w770 & w669) | (w770 & w2643) | (w669 & w2643);
assign w772 = ~w725 & w771;
assign w773 = (pi19 & ~w771) | (pi19 & w2179) | (~w771 & w2179);
assign w774 = w771 & w2180;
assign v169 = ~(w773 | w774);
assign w775 = v169;
assign w776 = w768 & w775;
assign v170 = ~(w768 | w775);
assign w777 = v170;
assign v171 = ~(w776 | w777);
assign w778 = v171;
assign w779 = (w2977 & w3793) | (w2977 & w3794) | (w3793 & w3794);
assign w780 = (w2997 & w2998) | (w2997 & ~w717) | (w2998 & ~w717);
assign w781 = (w780 & w721) | (w780 & w3795) | (w721 & w3795);
assign w782 = w778 & w781;
assign w783 = ~pi23 & w3062;
assign w784 = pi21 & ~w574;
assign w785 = (w783 & w574) | (w783 & w3796) | (w574 & w3796);
assign w786 = (~w2179 & w2644) | (~w2179 & w2645) | (w2644 & w2645);
assign w787 = ~w768 & w3000;
assign w788 = ~pi10 & w2;
assign w789 = pi01 & ~pi10;
assign v172 = ~(pi03 | w789);
assign w790 = v172;
assign v173 = ~(w788 | w790);
assign w791 = v173;
assign w792 = (w768 & w3001) | (w768 & w3002) | (w3001 & w3002);
assign w793 = (w792 & w762) | (w792 & w2450) | (w762 & w2450);
assign w794 = (~w590 & w3003) | (~w590 & w3004) | (w3003 & w3004);
assign w795 = (~w2171 & w4130) | (~w2171 & w4131) | (w4130 & w4131);
assign v174 = ~(w794 | w795);
assign w796 = v174;
assign v175 = ~(w629 | w640);
assign w797 = v175;
assign w798 = (w797 & w602) | (w797 & w3005) | (w602 & w3005);
assign w799 = (~w796 & w752) | (~w796 & w2183) | (w752 & w2183);
assign w800 = ~w752 & w2184;
assign v176 = ~(w799 | w800);
assign w801 = v176;
assign v177 = ~(pi05 | w801);
assign w802 = v177;
assign w803 = w724 & w2451;
assign w804 = (w579 & ~w589) | (w579 & w4132) | (~w589 & w4132);
assign w805 = (w2977 & w3798) | (w2977 & w3799) | (w3798 & w3799);
assign w806 = (w805 & w765) | (w805 & w3007) | (w765 & w3007);
assign w807 = ~w724 & w806;
assign v178 = ~(w2 | w789);
assign w808 = v178;
assign w809 = (w2977 & w3800) | (w2977 & w3801) | (w3800 & w3801);
assign w810 = (~pi12 & w789) | (~pi12 & w3009) | (w789 & w3009);
assign v179 = ~(w788 | w810);
assign w811 = v179;
assign w812 = (~w765 & w4133) | (~w765 & w4134) | (w4133 & w4134);
assign w813 = ~w690 & w3010;
assign w814 = w683 & w813;
assign w815 = ~w804 & w814;
assign w816 = ~w669 & w815;
assign w817 = (~w812 & ~w815) | (~w812 & w3802) | (~w815 & w3802);
assign w818 = ~w807 & w817;
assign w819 = (~w788 & ~w818) | (~w788 & w2452) | (~w818 & w2452);
assign w820 = (pi05 & w795) | (pi05 & w3011) | (w795 & w3011);
assign w821 = ~w795 & w3012;
assign v180 = ~(w820 | w821);
assign w822 = v180;
assign w823 = ~w752 & w2186;
assign w824 = (~w822 & w752) | (~w822 & w2187) | (w752 & w2187);
assign v181 = ~(w823 | w824);
assign w825 = v181;
assign w826 = w819 & ~w825;
assign v182 = ~(w802 | w826);
assign w827 = v182;
assign w828 = (w656 & w669) | (w656 & w2646) | (w669 & w2646);
assign w829 = ~w725 & w828;
assign v183 = ~(pi07 | w656);
assign w830 = v183;
assign v184 = ~(w657 | w830);
assign w831 = v184;
assign w832 = ~w647 & w831;
assign w833 = w647 & ~w831;
assign w834 = ~w603 & w3013;
assign w835 = ~w752 & w834;
assign v185 = ~(w829 | w835);
assign w836 = v185;
assign w837 = (pi09 & w835) | (pi09 & w2647) | (w835 & w2647);
assign w838 = w647 & w2909;
assign w839 = (w666 & ~w647) | (w666 & w2910) | (~w647 & w2910);
assign w840 = (~w660 & w602) | (~w660 & w2911) | (w602 & w2911);
assign v186 = ~(w838 | w839);
assign w841 = v186;
assign w842 = w840 & w841;
assign w843 = ~pi11 & w627;
assign w844 = pi11 & ~w627;
assign v187 = ~(w843 | w844);
assign w845 = v187;
assign w846 = ~w752 & w2188;
assign w847 = (~w845 & w752) | (~w845 & w2189) | (w752 & w2189);
assign v188 = ~(w846 | w847);
assign w848 = v188;
assign v189 = ~(w837 | w848);
assign w849 = v189;
assign w850 = w3015 & w4345;
assign w851 = (w3014 & w3803) | (w3014 & w3804) | (w3803 & w3804);
assign w852 = (w590 & w3805) | (w590 & w3806) | (w3805 & w3806);
assign w853 = (~w590 & w3018) | (~w590 & w3019) | (w3018 & w3019);
assign v190 = ~(w852 | w853);
assign w854 = v190;
assign w855 = ~w852 & w3020;
assign w856 = (pi07 & w852) | (pi07 & w3021) | (w852 & w3021);
assign v191 = ~(w855 | w856);
assign w857 = v191;
assign w858 = ~w752 & w2912;
assign w859 = (~w857 & w752) | (~w857 & w2913) | (w752 & w2913);
assign v192 = ~(w858 | w859);
assign w860 = v192;
assign w861 = ~w837 & w3022;
assign w862 = ~w827 & w861;
assign w863 = ~w835 & w2648;
assign w864 = (~pi07 & w852) | (~pi07 & w3023) | (w852 & w3023);
assign w865 = ~w752 & w2190;
assign w866 = (w855 & w752) | (w855 & w2191) | (w752 & w2191);
assign v193 = ~(w865 | w866);
assign w867 = v193;
assign w868 = ~w863 & w867;
assign w869 = w849 & ~w868;
assign w870 = ~pi11 & w848;
assign v194 = ~(w869 | w870);
assign w871 = v194;
assign w872 = ~w862 & w871;
assign w873 = (pi13 & w755) | (pi13 & w2192) | (w755 & w2192);
assign v195 = ~(w759 | w873);
assign w874 = v195;
assign w875 = w874 & w751;
assign w876 = w2193 & w3024;
assign w877 = ~w872 & w876;
assign w878 = pi12 & w4370;
assign v196 = ~(w816 | w878);
assign w879 = v196;
assign w880 = ~w807 & w879;
assign w881 = w879 & w3807;
assign w882 = (~pi05 & ~w880) | (~pi05 & w3025) | (~w880 & w3025);
assign w883 = ~w877 & w2453;
assign w884 = w880 & w3026;
assign w885 = (w884 & w877) | (w884 & w2454) | (w877 & w2454);
assign v197 = ~(w883 | w885);
assign w886 = v197;
assign w887 = w2193 & w3027;
assign w888 = ~w872 & w887;
assign w889 = (~w787 & w762) | (~w787 & w2455) | (w762 & w2455);
assign v198 = ~(w888 | w889);
assign w890 = v198;
assign w891 = pi07 & ~w801;
assign w892 = ~pi07 & w801;
assign v199 = ~(w891 | w892);
assign w893 = v199;
assign w894 = ~w888 & w2456;
assign w895 = ~w819 & w825;
assign v200 = ~(w826 | w895);
assign w896 = v200;
assign v201 = ~(pi07 | w896);
assign w897 = v201;
assign w898 = pi07 & w896;
assign v202 = ~(w897 | w898);
assign w899 = v202;
assign w900 = (w899 & w888) | (w899 & w2457) | (w888 & w2457);
assign v203 = ~(w894 | w900);
assign w901 = v203;
assign w902 = ~w872 & w875;
assign w903 = ~pi08 & w2;
assign w904 = pi01 & ~pi08;
assign v204 = ~(pi03 | w904);
assign w905 = v204;
assign w906 = (~pi10 & w904) | (~pi10 & w3028) | (w904 & w3028);
assign v205 = ~(w903 | w906);
assign w907 = v205;
assign v206 = ~(w2 | w904);
assign w908 = v206;
assign w909 = (w3797 & w4135) | (w3797 & w4136) | (w4135 & w4136);
assign w910 = w789 & ~w903;
assign w911 = (w910 & w768) | (w910 & w3808) | (w768 & w3808);
assign v207 = ~(w909 | w911);
assign w912 = v207;
assign w913 = (~w912 & w902) | (~w912 & w2459) | (w902 & w2459);
assign w914 = ~w762 & w2804;
assign w915 = ~w902 & w914;
assign v208 = ~(w913 | w915);
assign w916 = v208;
assign w917 = w880 & w3029;
assign w918 = ~w877 & w2460;
assign w919 = (pi05 & ~w880) | (pi05 & w3030) | (~w880 & w3030);
assign w920 = (w919 & w877) | (w919 & w2461) | (w877 & w2461);
assign v209 = ~(w918 | w920);
assign w921 = v209;
assign w922 = ~w916 & w921;
assign w923 = w886 & w901;
assign w924 = ~w922 & w923;
assign w925 = (~w896 & w888) | (~w896 & w2462) | (w888 & w2462);
assign w926 = ~w888 & w2463;
assign v210 = ~(w925 | w926);
assign w927 = v210;
assign w928 = pi07 & ~w927;
assign w929 = ~w752 & w3031;
assign w930 = (~w854 & w752) | (~w854 & w3032) | (w752 & w3032);
assign v211 = ~(w929 | w930);
assign w931 = v211;
assign w932 = pi09 & ~w931;
assign w933 = ~pi09 & w931;
assign v212 = ~(w932 | w933);
assign w934 = v212;
assign w935 = ~w888 & w2805;
assign w936 = (w860 & w826) | (w860 & w2194) | (w826 & w2194);
assign w937 = ~w826 & w3033;
assign v213 = ~(w936 | w937);
assign w938 = v213;
assign v214 = ~(pi09 | w938);
assign w939 = v214;
assign w940 = pi09 & w938;
assign v215 = ~(w939 | w940);
assign w941 = v215;
assign w942 = ~w890 & w941;
assign v216 = ~(w935 | w942);
assign w943 = v216;
assign w944 = ~w928 & w943;
assign w945 = ~w924 & w944;
assign w946 = (~w938 & w888) | (~w938 & w2464) | (w888 & w2464);
assign w947 = ~w888 & w2465;
assign v217 = ~(w946 | w947);
assign w948 = v217;
assign w949 = ~w946 & w2777;
assign w950 = ~w888 & w2466;
assign v218 = ~(w837 | w863);
assign w951 = v218;
assign w952 = w867 & w951;
assign w953 = ~w936 & w952;
assign v219 = ~(w867 | w951);
assign w954 = v219;
assign w955 = w860 & ~w951;
assign w956 = ~w827 & w955;
assign v220 = ~(w954 | w956);
assign w957 = v220;
assign w958 = ~w953 & w957;
assign w959 = ~w890 & w958;
assign v221 = ~(w950 | w959);
assign w960 = v221;
assign w961 = ~w959 & w2467;
assign v222 = ~(w949 | w961);
assign w962 = v222;
assign w963 = (w962 & w924) | (w962 & w2914) | (w924 & w2914);
assign w964 = (~w733 & ~w751) | (~w733 & w2195) | (~w751 & w2195);
assign w965 = (~w2196 & w4053) | (~w2196 & w4054) | (w4053 & w4054);
assign w966 = (~w772 & w764) | (~w772 & w2197) | (w764 & w2197);
assign w967 = (w3034 & w780) | (w3034 & w4033) | (w780 & w4033);
assign w968 = (w2196 & w4055) | (w2196 & w4056) | (w4055 & w4056);
assign w969 = w778 & w964;
assign w970 = ~w902 & w969;
assign w971 = (w2915 & w3809) | (w2915 & w3810) | (w3809 & w3810);
assign w972 = (w2915 & w3811) | (w2915 & w3812) | (w3811 & w3812);
assign v223 = ~(w778 | w972);
assign w973 = v223;
assign w974 = (~w2196 & w4057) | (~w2196 & w4058) | (w4057 & w4058);
assign v224 = ~(w970 | w974);
assign w975 = v224;
assign w976 = (w2197 & w4137) | (w2197 & w4138) | (w4137 & w4138);
assign v225 = ~(w3410 | w976);
assign w977 = v225;
assign w978 = ~w888 & w3813;
assign w979 = (~w978 & ~w975) | (~w978 & w3814) | (~w975 & w3814);
assign w980 = ~w888 & w2470;
assign v226 = ~(w731 | w733);
assign w981 = v226;
assign w982 = (~w749 & ~w873) | (~w749 & w4139) | (~w873 & w4139);
assign v227 = ~(w981 | w982);
assign w983 = v227;
assign w984 = w761 & ~w981;
assign w985 = w871 & w3815;
assign w986 = (~w787 & ~w751) | (~w787 & w2471) | (~w751 & w2471);
assign v228 = ~(w782 | w983);
assign w987 = v228;
assign w988 = w986 & w987;
assign w989 = w988 & w4059;
assign w990 = ~w989 & w2472;
assign v229 = ~(w979 | w990);
assign w991 = v229;
assign w992 = ~w870 & w874;
assign w993 = ~w869 & w992;
assign w994 = ~w862 & w993;
assign w995 = (~w874 & ~w871) | (~w874 & w3816) | (~w871 & w3816);
assign v230 = ~(w994 | w995);
assign w996 = v230;
assign v231 = ~(w890 | w996);
assign w997 = v231;
assign w998 = ~w888 & w2473;
assign w999 = ~w997 & w2474;
assign w1000 = pi11 & ~w848;
assign v232 = ~(w870 | w1000);
assign w1001 = v232;
assign w1002 = pi13 & w1001;
assign w1003 = ~w888 & w2475;
assign w1004 = w951 & w2198;
assign w1005 = ~w936 & w1004;
assign w1006 = w837 & w848;
assign v233 = ~(w869 | w1006);
assign w1007 = v233;
assign w1008 = ~w862 & w1007;
assign w1009 = ~w1005 & w1008;
assign w1010 = (pi13 & ~w1008) | (pi13 & w2199) | (~w1008 & w2199);
assign v234 = ~(w890 | w1010);
assign w1011 = v234;
assign v235 = ~(w1003 | w1011);
assign w1012 = v235;
assign w1013 = pi11 & ~w836;
assign w1014 = ~w888 & w2476;
assign w1015 = w957 & w2200;
assign v236 = ~(w890 | w1015);
assign w1016 = v236;
assign v237 = ~(w1014 | w1016);
assign w1017 = v237;
assign v238 = ~(w1012 | w1017);
assign w1018 = v238;
assign w1019 = ~w888 & w2477;
assign v239 = ~(w749 | w760);
assign w1020 = v239;
assign w1021 = w993 & w3817;
assign v240 = ~(w873 | w1020);
assign w1022 = v240;
assign w1023 = w873 & w1020;
assign v241 = ~(w1022 | w1023);
assign w1024 = v241;
assign w1025 = (w1024 & ~w993) | (w1024 & w4140) | (~w993 & w4140);
assign v242 = ~(w1021 | w1025);
assign w1026 = v242;
assign v243 = ~(w890 | w1026);
assign w1027 = v243;
assign v244 = ~(w1019 | w1027);
assign w1028 = v244;
assign w1029 = ~w1027 & w2478;
assign w1030 = (pi17 & w1027) | (pi17 & w2479) | (w1027 & w2479);
assign v245 = ~(w1029 | w1030);
assign w1031 = v245;
assign w1032 = ~w999 & w1018;
assign w1033 = w1031 & w1032;
assign w1034 = w1032 & w3818;
assign w1035 = ~w963 & w1034;
assign w1036 = ~w888 & w2480;
assign w1037 = ~w890 & w1009;
assign v246 = ~(w1036 | w1037);
assign w1038 = v246;
assign w1039 = (~pi13 & w1037) | (~pi13 & w2481) | (w1037 & w2481);
assign w1040 = (~pi15 & w997) | (~pi15 & w2482) | (w997 & w2482);
assign v247 = ~(w1039 | w1040);
assign w1041 = v247;
assign v248 = ~(w999 | w1030);
assign w1042 = v248;
assign w1043 = ~w1041 & w1042;
assign w1044 = (~pi19 & w989) | (~pi19 & w2483) | (w989 & w2483);
assign v249 = ~(w1029 | w1044);
assign w1045 = v249;
assign w1046 = (w991 & w1043) | (w991 & w2201) | (w1043 & w2201);
assign w1047 = (~w2806 & w3036) | (~w2806 & w3037) | (w3036 & w3037);
assign w1048 = (w789 & w888) | (w789 & w3819) | (w888 & w3819);
assign v250 = ~(w1047 | w1048);
assign w1049 = v250;
assign w1050 = pi23 & w3062;
assign w1051 = (w2420 & w3038) | (w2420 & w3039) | (w3038 & w3039);
assign v251 = ~(w903 | w905);
assign w1052 = v251;
assign w1053 = (w3039 & w3820) | (w3039 & w3821) | (w3820 & w3821);
assign v252 = ~(pi05 | w1053);
assign w1054 = v252;
assign w1055 = (w3039 & w3822) | (w3039 & w3823) | (w3822 & w3823);
assign v253 = ~(w1054 | w1055);
assign w1056 = v253;
assign w1057 = (~w1056 & w1047) | (~w1056 & w4141) | (w1047 & w4141);
assign w1058 = ~w1047 & w4142;
assign v254 = ~(w1057 | w1058);
assign w1059 = v254;
assign w1060 = (~w787 & w902) | (~w787 & w2202) | (w902 & w2202);
assign w1061 = ~w965 & w1060;
assign w1062 = ~w888 & w3824;
assign w1063 = (w888 & ~pi21) | (w888 & w2807) | (~pi21 & w2807);
assign w1064 = ~w1061 & w1063;
assign w1065 = (w971 & w902) | (w971 & w2203) | (w902 & w2203);
assign w1066 = w3796 & w778;
assign w1067 = w964 & w1066;
assign w1068 = (pi17 & w573) | (pi17 & w3041) | (w573 & w3041);
assign w1069 = (~pi19 & w573) | (~pi19 & w3825) | (w573 & w3825);
assign w1070 = ~w1068 & w1069;
assign w1071 = (w716 & w4143) | (w716 & w4144) | (w4143 & w4144);
assign w1072 = (w574 & w2919) | (w574 & w4371) | (w2919 & w4371);
assign w1073 = (~w966 & w4145) | (~w966 & w4146) | (w4145 & w4146);
assign w1074 = (w1073 & w902) | (w1073 & w2204) | (w902 & w2204);
assign w1075 = ~w1065 & w1074;
assign w1076 = (w1053 & ~w1074) | (w1053 & w4060) | (~w1074 & w4060);
assign w1077 = ~w1064 & w1076;
assign w1078 = ~w1059 & w1077;
assign w1079 = ~w1035 & w2205;
assign w1080 = (w2808 & w2201) | (w2808 & w3826) | (w2201 & w3826);
assign w1081 = (w1077 & ~w1033) | (w1077 & w2206) | (~w1033 & w2206);
assign w1082 = w962 & w1077;
assign w1083 = (w1059 & w945) | (w1059 & w3043) | (w945 & w3043);
assign w1084 = ~w1081 & w1083;
assign v255 = ~(w1080 | w1084);
assign w1085 = v255;
assign w1086 = ~w1079 & w1085;
assign w1087 = ~pi06 & w2;
assign w1088 = (pi08 & ~w2) | (pi08 & w3044) | (~w2 & w3044);
assign w1089 = (w3039 & w3827) | (w3039 & w3828) | (w3827 & w3828);
assign w1090 = w1088 & ~w1089;
assign w1091 = (w2201 & w2809) | (w2201 & w2810) | (w2809 & w2810);
assign w1092 = ~w1075 & w1088;
assign w1093 = ~w1064 & w1092;
assign w1094 = (w1093 & ~w1033) | (w1093 & w2207) | (~w1033 & w2207);
assign w1095 = (~w1090 & w945) | (~w1090 & w2778) | (w945 & w2778);
assign w1096 = ~w1094 & w1095;
assign v256 = ~(w1091 | w1096);
assign w1097 = v256;
assign w1098 = pi01 & ~pi06;
assign v257 = ~(pi03 | w1098);
assign w1099 = v257;
assign w1100 = w904 & ~w1087;
assign w1101 = ~w1099 & w4346;
assign w1102 = (w2201 & w2811) | (w2201 & w2812) | (w2811 & w2812);
assign w1103 = (~w1099 & ~w1074) | (~w1099 & w4061) | (~w1074 & w4061);
assign w1104 = ~w1064 & w1103;
assign w1105 = (w1104 & ~w1033) | (w1104 & w2208) | (~w1033 & w2208);
assign w1106 = w962 & w1104;
assign w1107 = (~w1101 & w945) | (~w1101 & w2779) | (w945 & w2779);
assign w1108 = ~w1105 & w1107;
assign v258 = ~(w1102 | w1108);
assign w1109 = v258;
assign w1110 = ~w1097 & w1109;
assign w1111 = ~w1086 & w1110;
assign v259 = ~(w1064 | w1075);
assign w1112 = v259;
assign w1113 = ~w991 & w1112;
assign w1114 = w1045 & w1112;
assign w1115 = ~w1043 & w1114;
assign v260 = ~(w1113 | w1115);
assign w1116 = v260;
assign v261 = ~(w1035 | w1116);
assign w1117 = v261;
assign w1118 = (w2209 & w1035) | (w2209 & w2813) | (w1035 & w2813);
assign w1119 = (~w1035 & w2814) | (~w1035 & w2815) | (w2814 & w2815);
assign v262 = ~(w1118 | w1119);
assign w1120 = v262;
assign w1121 = (w1120 & w1086) | (w1120 & w2881) | (w1086 & w2881);
assign w1122 = (~w881 & w877) | (~w881 & w3829) | (w877 & w3829);
assign w1123 = ~w877 & w3830;
assign v263 = ~(w1122 | w1123);
assign w1124 = v263;
assign w1125 = pi07 & ~w1124;
assign w1126 = ~pi07 & w1124;
assign v264 = ~(w1125 | w1126);
assign w1127 = v264;
assign w1128 = ~w913 & w3048;
assign w1129 = (~pi05 & w913) | (~pi05 & w3049) | (w913 & w3049);
assign v265 = ~(w4147 | w1128);
assign w1130 = v265;
assign w1131 = ~w1129 & w1130;
assign w1132 = (w2816 & w3831) | (w2816 & w3832) | (w3831 & w3832);
assign w1133 = (~w2816 & w3833) | (~w2816 & w3834) | (w3833 & w3834);
assign v266 = ~(w1132 | w1133);
assign w1134 = v266;
assign w1135 = (w2881 & w3835) | (w2881 & w3836) | (w3835 & w3836);
assign w1136 = (~w4147 & w1035) | (~w4147 & w2484) | (w1035 & w2484);
assign w1137 = (w886 & w916) | (w886 & w2882) | (w916 & w2882);
assign v267 = ~(w901 | w1137);
assign w1138 = v267;
assign v268 = ~(w924 | w1138);
assign w1139 = v268;
assign w1140 = (w2210 & w1035) | (w2210 & w3765) | (w1035 & w3765);
assign w1141 = ~pi09 & w927;
assign w1142 = ~w1051 & w4373;
assign w1143 = (~w1142 & w1035) | (~w1142 & w2817) | (w1035 & w2817);
assign w1144 = ~w1140 & w1143;
assign w1145 = (~w1035 & w2818) | (~w1035 & w2819) | (w2818 & w2819);
assign w1146 = w1127 & w1137;
assign w1147 = (w2211 & w1035) | (w2211 & w2820) | (w1035 & w2820);
assign v269 = ~(w1145 | w1147);
assign w1148 = v269;
assign w1149 = ~w1144 & w1148;
assign w1150 = (~w943 & w924) | (~w943 & w2883) | (w924 & w2883);
assign v270 = ~(w945 | w1150);
assign w1151 = v270;
assign w1152 = ~pi11 & w1151;
assign w1153 = (w2484 & w3837) | (w2484 & w3838) | (w3837 & w3838);
assign w1154 = ~w946 & w3050;
assign w1155 = w4147 & ~w1154;
assign w1156 = ~w1064 & w3839;
assign w1157 = (~w1155 & w1035) | (~w1155 & w2821) | (w1035 & w2821);
assign w1158 = ~w1153 & w1157;
assign w1159 = pi11 & ~w1151;
assign w1160 = (w2484 & w3840) | (w2484 & w3841) | (w3840 & w3841);
assign w1161 = (pi11 & w946) | (pi11 & w3051) | (w946 & w3051);
assign w1162 = (~w1035 & w4084) | (~w1035 & w4085) | (w4084 & w4085);
assign v271 = ~(w1160 | w1162);
assign w1163 = v271;
assign v272 = ~(w1158 | w1163);
assign w1164 = v272;
assign w1165 = w1149 & w1164;
assign w1166 = ~w1135 & w1165;
assign w1167 = (~w1038 & w2213) | (~w1038 & w1117) | (w2213 & w1117);
assign v273 = ~(w1012 | w1039);
assign w1168 = v273;
assign w1169 = ~w1168 & w3758;
assign w1170 = (w945 & w2884) | (w945 & w2885) | (w2884 & w2885);
assign v274 = ~(w1169 | w1170);
assign w1171 = v274;
assign w1172 = w1136 & w1171;
assign v275 = ~(w1167 | w1172);
assign w1173 = v275;
assign w1174 = (~pi15 & w1172) | (~pi15 & w2215) | (w1172 & w2215);
assign w1175 = ~w1037 & w3052;
assign w1176 = (w3039 & w3842) | (w3039 & w3843) | (w3842 & w3843);
assign w1177 = (~w1175 & w2216) | (~w1175 & w1117) | (w2216 & w1117);
assign v276 = ~(w1172 | w1177);
assign w1178 = v276;
assign v277 = ~(w1174 | w1178);
assign w1179 = v277;
assign w1180 = (w2217 & w1035) | (w2217 & w3766) | (w1035 & w3766);
assign w1181 = pi09 & ~w927;
assign w1182 = (w4147 & w927) | (w4147 & w3054) | (w927 & w3054);
assign w1183 = (~w1182 & w1035) | (~w1182 & w2822) | (w1035 & w2822);
assign w1184 = ~w1180 & w1183;
assign w1185 = ~w1158 & w1184;
assign w1186 = (~pi13 & w1160) | (~pi13 & w2218) | (w1160 & w2218);
assign w1187 = ~w1185 & w1186;
assign w1188 = w1179 & w1187;
assign w1189 = ~w1166 & w1188;
assign w1190 = (pi13 & w1153) | (pi13 & w2219) | (w1153 & w2219);
assign w1191 = w1149 & w1190;
assign w1192 = ~w1135 & w1191;
assign v278 = ~(w1163 | w1184);
assign w1193 = v278;
assign w1194 = w1190 & ~w1193;
assign w1195 = (~w949 & w924) | (~w949 & w2886) | (w924 & w2886);
assign w1196 = w1034 & ~w1195;
assign w1197 = (~w960 & w2220) | (~w960 & w3772) | (w2220 & w3772);
assign v279 = ~(w961 | w1017);
assign w1198 = v279;
assign v280 = ~(w1198 | w1195);
assign w1199 = v280;
assign w1200 = (w3844 & w2886) | (w3844 & w4062) | (w2886 & w4062);
assign v281 = ~(w1199 | w1200);
assign w1201 = v281;
assign w1202 = (w2484 & w3845) | (w2484 & w3846) | (w3845 & w3846);
assign v282 = ~(w1197 | w1202);
assign w1203 = v282;
assign w1204 = ~w1178 & w1203;
assign w1205 = ~w1174 & w1204;
assign w1206 = ~w1194 & w1205;
assign w1207 = ~w1192 & w1206;
assign v283 = ~(w1189 | w1207);
assign w1208 = v283;
assign v284 = ~(w1018 | w1039);
assign w1209 = v284;
assign w1210 = w962 & ~w1039;
assign w1211 = ~w945 & w1210;
assign v285 = ~(w999 | w1040);
assign w1212 = v285;
assign w1213 = (w1212 & w1211) | (w1212 & w2221) | (w1211 & w2221);
assign w1214 = ~w1211 & w2222;
assign v286 = ~(w1213 | w1214);
assign w1215 = v286;
assign w1216 = w1136 & w1215;
assign w1217 = (w1117 & w3767) | (w1117 & w2223) | (w3767 & w2223);
assign v287 = ~(w1216 | w1217);
assign w1218 = v287;
assign w1219 = ~w1216 & w2224;
assign v288 = ~(w1174 | w1219);
assign w1220 = v288;
assign w1221 = ~w990 & w1018;
assign w1222 = w1221 & w2485;
assign w1223 = ~w963 & w1222;
assign v289 = ~(w990 | w1044);
assign w1224 = v289;
assign w1225 = (w1224 & w1043) | (w1224 & w2225) | (w1043 & w2225);
assign w1226 = (~w1225 & w963) | (~w1225 & w2887) | (w963 & w2887);
assign w1227 = ~w963 & w1033;
assign w1228 = ~w1043 & w2226;
assign w1229 = (w1228 & w963) | (w1228 & w2888) | (w963 & w2888);
assign w1230 = w1226 & ~w1229;
assign w1231 = w1136 & ~w1230;
assign w1232 = (w1117 & w3847) | (w1117 & w2227) | (w3847 & w2227);
assign v290 = ~(w1231 | w1232);
assign w1233 = v290;
assign w1234 = (pi21 & w1231) | (pi21 & w2228) | (w1231 & w2228);
assign w1235 = (w1211 & w2651) | (w1211 & w2652) | (w2651 & w2652);
assign w1236 = ~w1029 & w1043;
assign w1237 = w999 & ~w1031;
assign w1238 = (w3039 & w3848) | (w3039 & w3849) | (w3848 & w3849);
assign w1239 = (w1238 & w1031) | (w1238 & w2229) | (w1031 & w2229);
assign w1240 = ~w1236 & w1239;
assign w1241 = w1116 & w1240;
assign w1242 = w1241 & w2653;
assign w1243 = (w1117 & w4063) | (w1117 & w4064) | (w4063 & w4064);
assign v291 = ~(w1242 | w1243);
assign w1244 = v291;
assign w1245 = (~pi21 & w989) | (~pi21 & w3057) | (w989 & w3057);
assign w1246 = (w3039 & w3850) | (w3039 & w3851) | (w3850 & w3851);
assign w1247 = (~w1245 & w2230) | (~w1245 & w1117) | (w2230 & w1117);
assign v292 = ~(w1231 | w1247);
assign w1248 = v292;
assign w1249 = w1244 & ~w1248;
assign v293 = ~(w1234 | w1249);
assign w1250 = v293;
assign w1251 = w1220 & ~w1250;
assign w1252 = (~w2484 & w2654) | (~w2484 & w2655) | (w2654 & w2655);
assign v294 = ~(w1236 | w1237);
assign w1253 = v294;
assign w1254 = ~w1227 & w1253;
assign w1255 = w1136 & w2231;
assign v295 = ~(w1252 | w1255);
assign w1256 = v295;
assign w1257 = ~w1255 & w2656;
assign w1258 = (pi17 & w1216) | (pi17 & w2232) | (w1216 & w2232);
assign w1259 = (w1244 & w1257) | (w1244 & w2823) | (w1257 & w2823);
assign v296 = ~(w1234 | w1248);
assign w1260 = v296;
assign w1261 = ~w1259 & w1260;
assign v297 = ~(w1250 | w1261);
assign w1262 = v297;
assign w1263 = (~w1262 & ~w1208) | (~w1262 & w2657) | (~w1208 & w2657);
assign v298 = ~(w1061 | w1062);
assign w1264 = v298;
assign w1265 = (pi23 & w1061) | (pi23 & w3852) | (w1061 & w3852);
assign w1266 = (~w1265 & w2233) | (~w1265 & w1117) | (w2233 & w1117);
assign w1267 = w979 & w1224;
assign w1268 = ~w1223 & w2234;
assign w1269 = w979 & w990;
assign w1270 = ~w1269 & w2486;
assign w1271 = ~w1035 & w2235;
assign w1272 = ~w1268 & w1271;
assign v299 = ~(w1266 | w1272);
assign w1273 = v299;
assign w1274 = ~w1249 & w2236;
assign w1275 = (w2237 & w1035) | (w2237 & w2487) | (w1035 & w2487);
assign w1276 = (w1072 & w902) | (w1072 & w3058) | (w902 & w3058);
assign w1277 = ~w1065 & w1276;
assign w1278 = (~w902 & w3059) | (~w902 & w3060) | (w3059 & w3060);
assign w1279 = ~w1035 & w2238;
assign w1280 = ~w1061 & w3853;
assign w1281 = (w1280 & w1279) | (w1280 & w2824) | (w1279 & w2824);
assign w1282 = ~w1269 & w3061;
assign w1283 = ~w1035 & w2825;
assign w1284 = ~w1268 & w1283;
assign v300 = ~(w1281 | w1284);
assign w1285 = v300;
assign w1286 = ~w2488 & w1285;
assign w1287 = w1220 & w1286;
assign w1288 = ~w1274 & w1287;
assign w1289 = ~w1207 & w3854;
assign w1290 = ~pi27 & w14;
assign w1291 = (w1290 & w1277) | (w1290 & w3062) | (w1277 & w3062);
assign w1292 = (w1291 & ~w1273) | (w1291 & w2488) | (~w1273 & w2488);
assign w1293 = ~w1249 & w2658;
assign w1294 = (w1291 & ~w1285) | (w1291 & w2488) | (~w1285 & w2488);
assign w1295 = (~w1294 & ~w2658) | (~w1294 & w2826) | (~w2658 & w2826);
assign w1296 = w1244 & ~w1257;
assign v301 = ~(w1234 | w1258);
assign w1297 = v301;
assign w1298 = w1292 & w1297;
assign w1299 = w1296 & w1298;
assign w1300 = w1295 & ~w1299;
assign w1301 = ~w1273 & w1285;
assign w1302 = (w1301 & ~w1295) | (w1301 & w2239) | (~w1295 & w2239);
assign w1303 = ~w1289 & w1302;
assign w1304 = w1263 & w1303;
assign w1305 = (~w1300 & ~w1208) | (~w1300 & w2663) | (~w1208 & w2663);
assign w1306 = w1264 & ~w1136;
assign v302 = ~(w1272 | w1306);
assign w1307 = v302;
assign w1308 = (w1307 & w1289) | (w1307 & w2240) | (w1289 & w2240);
assign v303 = ~(w1300 | w1301);
assign w1309 = v303;
assign w1310 = ~w1263 & w1309;
assign w1311 = (~pi25 & w1263) | (~pi25 & w2241) | (w1263 & w2241);
assign w1312 = ~w1304 & w2659;
assign w1313 = (~w1289 & w3478) | (~w1289 & w3063) | (w3478 & w3063);
assign w1314 = w14 & ~w1313;
assign w1315 = (w1314 & ~w2659) | (w1314 & w3855) | (~w2659 & w3855);
assign w1316 = (~w1233 & w1289) | (~w1233 & w2242) | (w1289 & w2242);
assign w1317 = ~w1219 & w4148;
assign w1318 = ~w1207 & w3856;
assign w1319 = w1261 & ~w1300;
assign w1320 = ~w1318 & w1319;
assign w1321 = (w1207 & w3857) | (w1207 & w3858) | (w3857 & w3858);
assign v304 = ~(w1260 | w1295);
assign w1322 = v304;
assign w1323 = (w1208 & w3064) | (w1208 & w3065) | (w3064 & w3065);
assign v305 = ~(w1316 | w1320);
assign w1324 = v305;
assign w1325 = ~w1323 & w1324;
assign w1326 = (pi23 & ~w1324) | (pi23 & w2489) | (~w1324 & w2489);
assign w1327 = ~w1304 & w3066;
assign w1328 = (w1304 & pi25) | (w1304 & w2660) | (pi25 & w2660);
assign v306 = ~(w1326 | w1328);
assign w1329 = v306;
assign w1330 = w1315 & w1329;
assign w1331 = (~w1289 & w3481) | (~w1289 & w3067) | (w3481 & w3067);
assign w1332 = (w1289 & w4086) | (w1289 & w4087) | (w4086 & w4087);
assign w1333 = (~w1332 & ~w2659) | (~w1332 & w3859) | (~w2659 & w3859);
assign w1334 = (w1314 & w1312) | (w1314 & w2245) | (w1312 & w2245);
assign v307 = ~(w1330 | w1334);
assign w1335 = v307;
assign w1336 = pi01 & ~pi04;
assign w1337 = ~pi02 & w2;
assign w1338 = w1336 & ~w1337;
assign w1339 = ~w1 & w4097;
assign w1340 = ~pi04 & w2;
assign w1341 = (pi06 & w1289) | (pi06 & w2247) | (w1289 & w2247);
assign v308 = ~(pi03 | w1336);
assign w1342 = v308;
assign w1343 = (w1098 & ~w1295) | (w1098 & w2248) | (~w1295 & w2248);
assign w1344 = ~w1289 & w1343;
assign w1345 = (~w1342 & w1289) | (~w1342 & w2249) | (w1289 & w2249);
assign w1346 = ~w1341 & w1345;
assign v309 = ~(w1340 | w1346);
assign w1347 = v309;
assign v310 = ~(w1087 | w1099);
assign w1348 = v310;
assign w1349 = (w1348 & ~w1295) | (w1348 & w2250) | (~w1295 & w2250);
assign w1350 = pi08 & w4034;
assign w1351 = w904 & w1136;
assign v311 = ~(w1350 | w1351);
assign w1352 = v311;
assign w1353 = (pi05 & w1351) | (pi05 & w3860) | (w1351 & w3860);
assign w1354 = ~w1351 & w3861;
assign v312 = ~(w1353 | w1354);
assign w1355 = v312;
assign w1356 = ~w1289 & w2490;
assign w1357 = (~w1355 & w1289) | (~w1355 & w2491) | (w1289 & w2491);
assign v313 = ~(w1356 | w1357);
assign w1358 = v313;
assign v314 = ~(w1347 | w1358);
assign w1359 = v314;
assign w1360 = ~w1289 & w2251;
assign w1361 = ~w1351 & w3862;
assign w1362 = (w1361 & w1289) | (w1361 & w2252) | (w1289 & w2252);
assign v315 = ~(w1360 | w1362);
assign w1363 = v315;
assign w1364 = w1086 & ~w1110;
assign v316 = ~(w1111 | w1364);
assign w1365 = v316;
assign w1366 = pi07 & ~w1365;
assign w1367 = ~pi07 & w1365;
assign v317 = ~(w1366 | w1367);
assign w1368 = v317;
assign w1369 = ~w1289 & w2253;
assign w1370 = w1049 & w4035;
assign w1371 = (w3047 & w3863) | (w3047 & w3864) | (w3863 & w3864);
assign v318 = ~(w1370 | w1371);
assign w1372 = v318;
assign v319 = ~(pi07 | w1372);
assign w1373 = v319;
assign w1374 = pi07 & w1372;
assign v320 = ~(w1373 | w1374);
assign w1375 = v320;
assign w1376 = (w1375 & w1289) | (w1375 & w2254) | (w1289 & w2254);
assign v321 = ~(w1369 | w1376);
assign w1377 = v321;
assign w1378 = w1363 & w1377;
assign w1379 = w1134 & ~w1121;
assign v322 = ~(w1135 | w1379);
assign w1380 = v322;
assign w1381 = pi09 & ~w1380;
assign w1382 = ~w1289 & w2255;
assign w1383 = ~w1124 & w4036;
assign w1384 = (w2816 & w3865) | (w2816 & w3866) | (w3865 & w3866);
assign v323 = ~(w1383 | w1384);
assign w1385 = v323;
assign w1386 = pi09 & ~w1385;
assign w1387 = (~w1386 & w1289) | (~w1386 & w2256) | (w1289 & w2256);
assign v324 = ~(w1382 | w1387);
assign w1388 = v324;
assign w1389 = w1378 & ~w1388;
assign w1390 = ~w1359 & w1389;
assign w1391 = (~w1365 & ~w1295) | (~w1365 & w2257) | (~w1295 & w2257);
assign w1392 = ~w1289 & w1391;
assign w1393 = w1295 & w2258;
assign w1394 = w1287 & w2492;
assign w1395 = w1208 & w1394;
assign v325 = ~(w1393 | w1395);
assign w1396 = v325;
assign w1397 = ~w1392 & w1396;
assign w1398 = (~pi07 & ~w1396) | (~pi07 & w3867) | (~w1396 & w3867);
assign w1399 = ~pi09 & w1380;
assign v326 = ~(w1381 | w1399);
assign w1400 = v326;
assign w1401 = ~w1289 & w2259;
assign w1402 = ~pi09 & w1385;
assign v327 = ~(w1386 | w1402);
assign w1403 = v327;
assign w1404 = (w1403 & w1289) | (w1403 & w2260) | (w1289 & w2260);
assign v328 = ~(w1401 | w1404);
assign w1405 = v328;
assign v329 = ~(w1398 | w1405);
assign w1406 = v329;
assign w1407 = (~w2261 & w4088) | (~w2261 & w4089) | (w4088 & w4089);
assign w1408 = ~w1390 & w1407;
assign v330 = ~(pi11 | w1388);
assign w1409 = v330;
assign w1410 = w1378 & w1409;
assign w1411 = ~w1359 & w1410;
assign w1412 = ~w1406 & w1409;
assign w1413 = w927 & ~w1136;
assign w1414 = (w2484 & w3868) | (w2484 & w3869) | (w3868 & w3869);
assign v331 = ~(w1413 | w1414);
assign w1415 = v331;
assign w1416 = (w1415 & w1289) | (w1415 & w2493) | (w1289 & w2493);
assign v332 = ~(w1144 | w1184);
assign w1417 = v332;
assign w1418 = (w1121 & w3870) | (w1121 & w3871) | (w3870 & w3871);
assign w1419 = w1148 & w1417;
assign w1420 = ~w1135 & w1419;
assign v333 = ~(w1418 | w1420);
assign w1421 = v333;
assign w1422 = ~w1289 & w2494;
assign v334 = ~(w1416 | w1422);
assign w1423 = v334;
assign w1424 = (~w1423 & w1406) | (~w1423 & w2262) | (w1406 & w2262);
assign w1425 = ~w1411 & w1424;
assign v335 = ~(w1408 | w1425);
assign w1426 = v335;
assign w1427 = w1296 & ~w1295;
assign w1428 = (w1208 & w3070) | (w1208 & w3071) | (w3070 & w3071);
assign w1429 = ~w1207 & w3872;
assign w1430 = (w1293 & w2827) | (w1293 & w2828) | (w2827 & w2828);
assign w1431 = (w1430 & ~w1208) | (w1430 & w2661) | (~w1208 & w2661);
assign w1432 = ~w1274 & w4332;
assign w1433 = (~w1256 & ~w1297) | (~w1256 & w3873) | (~w1297 & w3873);
assign w1434 = w1295 & w1433;
assign w1435 = (~w1434 & ~w1208) | (~w1434 & w2662) | (~w1208 & w2662);
assign w1436 = ~w1431 & w1435;
assign w1437 = w1435 & w4149;
assign w1438 = w1435 & w4333;
assign w1439 = (~pi21 & ~w1436) | (~pi21 & w2265) | (~w1436 & w2265);
assign v336 = ~(w1438 | w1439);
assign w1440 = v336;
assign w1441 = (~w1293 & w3072) | (~w1293 & w3073) | (w3072 & w3073);
assign w1442 = w1218 & w1300;
assign v337 = ~(w1219 | w1258);
assign w1443 = v337;
assign w1444 = ~w1207 & w3874;
assign v338 = ~(w1300 | w1443);
assign w1445 = v338;
assign w1446 = ~w1444 & w1445;
assign w1447 = (~w1442 & ~w1429) | (~w1442 & w3074) | (~w1429 & w3074);
assign w1448 = ~w1446 & w1447;
assign w1449 = w1447 & w2266;
assign w1450 = ~w1439 & w4334;
assign w1451 = w1164 & ~w1184;
assign w1452 = ~w1164 & w1184;
assign v339 = ~(w1451 | w1452);
assign w1453 = v339;
assign w1454 = ~w1420 & w1453;
assign v340 = ~(w1166 | w1454);
assign w1455 = v340;
assign w1456 = ~w1300 & w1455;
assign w1457 = ~w1289 & w1456;
assign w1458 = (w2484 & w3875) | (w2484 & w3876) | (w3875 & w3876);
assign v341 = ~(w948 | w1136);
assign w1459 = v341;
assign v342 = ~(w1458 | w1459);
assign w1460 = v342;
assign w1461 = w1295 & w2267;
assign w1462 = w1287 & w2495;
assign w1463 = w1208 & w1462;
assign v343 = ~(w1461 | w1463);
assign w1464 = v343;
assign w1465 = ~w1457 & w1464;
assign w1466 = (pi13 & ~w1464) | (pi13 & w3877) | (~w1464 & w3877);
assign w1467 = w1464 & w3878;
assign v344 = ~(w1466 | w1467);
assign w1468 = v344;
assign w1469 = ~w1172 & w3075;
assign w1470 = (~w1469 & w1289) | (~w1469 & w2269) | (w1289 & w2269);
assign w1471 = (w1187 & w1135) | (w1187 & w2780) | (w1135 & w2780);
assign w1472 = (~w1194 & w1135) | (~w1194 & w2781) | (w1135 & w2781);
assign w1473 = (w2781 & w3076) | (w2781 & w3077) | (w3076 & w3077);
assign v345 = ~(w1179 | w1471);
assign w1474 = v345;
assign w1475 = ~w1473 & w1474;
assign w1476 = w2663 & w4150;
assign v346 = ~(w1470 | w1476);
assign w1477 = v346;
assign w1478 = ~w1471 & w1472;
assign w1479 = ~w1300 & w1478;
assign w1480 = ~w1289 & w1479;
assign w1481 = ~w1202 & w3078;
assign w1482 = ~w1289 & w2782;
assign w1483 = (pi15 & w1202) | (pi15 & w3079) | (w1202 & w3079);
assign w1484 = (w1483 & w1289) | (w1483 & w2783) | (w1289 & w2783);
assign v347 = ~(w1482 | w1484);
assign w1485 = v347;
assign w1486 = ~w1477 & w1485;
assign w1487 = w1468 & w1486;
assign w1488 = w1450 & w1487;
assign w1489 = w1426 & w1488;
assign w1490 = ~w1202 & w3080;
assign v348 = ~(w1483 | w1490);
assign w1491 = v348;
assign w1492 = w1480 & w1491;
assign v349 = ~(w1480 | w1491);
assign w1493 = v349;
assign v350 = ~(w1492 | w1493);
assign w1494 = v350;
assign w1495 = ~w1467 & w1494;
assign w1496 = w1486 & ~w1495;
assign w1497 = (~pi19 & ~w1447) | (~pi19 & w2270) | (~w1447 & w2270);
assign w1498 = (~w1173 & w1289) | (~w1173 & w2271) | (w1289 & w2271);
assign v351 = ~(w1476 | w1498);
assign w1499 = v351;
assign w1500 = (~pi17 & w1476) | (~pi17 & w2272) | (w1476 & w2272);
assign v352 = ~(w1497 | w1500);
assign w1501 = v352;
assign w1502 = ~w1496 & w1501;
assign w1503 = (w1450 & w1496) | (w1450 & w2664) | (w1496 & w2664);
assign w1504 = w1324 & w2496;
assign v353 = ~(w1439 | w1504);
assign w1505 = v353;
assign w1506 = (w1312 & w3879) | (w1312 & w3880) | (w3879 & w3880);
assign w1507 = (~w1 & w3081) | (~w1 & ~w1334) | (w3081 & ~w1334);
assign w1508 = (w1502 & w3082) | (w1502 & w3083) | (w3082 & w3083);
assign w1509 = (~w1339 & w1489) | (~w1339 & w3084) | (w1489 & w3084);
assign w1510 = (pi04 & ~w2) | (pi04 & w3881) | (~w2 & w3881);
assign w1511 = (pi01 & w1330) | (pi01 & w3085) | (w1330 & w3085);
assign w1512 = w1510 & ~w1511;
assign w1513 = ~pi01 & pi04;
assign w1514 = (w1312 & w3882) | (w1312 & w3883) | (w3882 & w3883);
assign w1515 = (w1502 & w4090) | (w1502 & w4091) | (w4090 & w4091);
assign w1516 = (~w1512 & w1489) | (~w1512 & w4092) | (w1489 & w4092);
assign w1517 = ~w1509 & w1516;
assign v354 = ~(w1340 | w1342);
assign w1518 = v354;
assign w1519 = ~w1313 & w3087;
assign w1520 = ~w1312 & w3088;
assign w1521 = w1329 & w1520;
assign w1522 = (~w1502 & w4093) | (~w1502 & w4094) | (w4093 & w4094);
assign w1523 = w1488 & w1521;
assign w1524 = w1426 & w1523;
assign v355 = ~(w1341 | w1344);
assign w1525 = v355;
assign w1526 = (~w3859 & w4151) | (~w3859 & w4152) | (w4151 & w4152);
assign w1527 = (w3859 & w4153) | (w3859 & w4154) | (w4153 & w4154);
assign v356 = ~(w1526 | w1527);
assign w1528 = v356;
assign w1529 = ~w1525 & w1528;
assign w1530 = w1525 & ~w1528;
assign v357 = ~(w1529 | w1530);
assign w1531 = v357;
assign w1532 = ~w1524 & w4335;
assign w1533 = (~w1531 & w1524) | (~w1531 & w4336) | (w1524 & w4336);
assign v358 = ~(w1532 | w1533);
assign w1534 = v358;
assign v359 = ~(w1517 | w1534);
assign w1535 = v359;
assign w1536 = w1333 & w1505;
assign w1537 = (~w2664 & w3884) | (~w2664 & w3885) | (w3884 & w3885);
assign v360 = ~(w1335 | w1537);
assign w1538 = v360;
assign w1539 = w1330 & w1488;
assign w1540 = w1426 & w1539;
assign v361 = ~(w1538 | w1540);
assign w1541 = v361;
assign w1542 = w1518 & w1525;
assign w1543 = (w1542 & w1538) | (w1542 & w2276) | (w1538 & w2276);
assign w1544 = (~pi05 & w1543) | (~pi05 & w3089) | (w1543 & w3089);
assign v362 = ~(w1535 | w1544);
assign w1545 = v362;
assign w1546 = w1347 & w1358;
assign v363 = ~(w1359 | w1546);
assign w1547 = v363;
assign w1548 = (~w1547 & w1538) | (~w1547 & w2278) | (w1538 & w2278);
assign w1549 = (~w1352 & w1289) | (~w1352 & w3090) | (w1289 & w3090);
assign w1550 = ~w1289 & w3091;
assign v364 = ~(w1549 | w1550);
assign w1551 = v364;
assign w1552 = ~w1538 & w2279;
assign v365 = ~(w1548 | w1552);
assign w1553 = v365;
assign w1554 = pi07 & w1553;
assign v366 = ~(pi07 | w1553);
assign w1555 = v366;
assign v367 = ~(w1554 | w1555);
assign w1556 = v367;
assign w1557 = w1545 & w1556;
assign w1558 = (w1363 & w1347) | (w1363 & w3092) | (w1347 & w3092);
assign v368 = ~(w1377 | w1558);
assign w1559 = v368;
assign w1560 = ~w1359 & w1378;
assign v369 = ~(w1559 | w1560);
assign w1561 = v369;
assign w1562 = (w1561 & w1538) | (w1561 & w2280) | (w1538 & w2280);
assign w1563 = ~w1538 & w2281;
assign v370 = ~(w1562 | w1563);
assign w1564 = v370;
assign v371 = ~(pi09 | w1564);
assign w1565 = v371;
assign w1566 = pi09 & w1564;
assign v372 = ~(w1565 | w1566);
assign w1567 = v372;
assign w1568 = ~w1554 & w1567;
assign w1569 = ~w1557 & w1568;
assign v373 = ~(w1411 | w1412);
assign w1570 = v373;
assign w1571 = ~w1408 & w1570;
assign w1572 = (~w2282 & w2665) | (~w2282 & w2666) | (w2665 & w2666);
assign w1573 = w1423 & w1571;
assign w1574 = (w1573 & w1538) | (w1573 & w2283) | (w1538 & w2283);
assign w1575 = (~w2283 & w2667) | (~w2283 & w2668) | (w2667 & w2668);
assign w1576 = ~w1572 & w1575;
assign w1577 = pi13 & ~w1426;
assign w1578 = ~pi13 & w1426;
assign v374 = ~(w1577 | w1578);
assign w1579 = v374;
assign w1580 = (pi15 & ~w1464) | (pi15 & w3886) | (~w1464 & w3886);
assign w1581 = w1464 & w3887;
assign v375 = ~(w1580 | w1581);
assign w1582 = v375;
assign w1583 = ~w1541 & w2284;
assign w1584 = (~w1582 & w1541) | (~w1582 & w2285) | (w1541 & w2285);
assign v376 = ~(w1583 | w1584);
assign w1585 = v376;
assign w1586 = ~w1576 & w1585;
assign w1587 = w1385 & ~w1305;
assign w1588 = ~w1300 & w4347;
assign v377 = ~(w1587 | w1588);
assign w1589 = v377;
assign v378 = ~(pi11 | w1589);
assign w1590 = v378;
assign w1591 = pi11 & w1589;
assign v379 = ~(w1590 | w1591);
assign w1592 = v379;
assign w1593 = ~w1538 & w2497;
assign w1594 = (~w1398 & w1359) | (~w1398 & w2498) | (w1359 & w2498);
assign w1595 = ~w1405 & w1594;
assign w1596 = w1405 & ~w1594;
assign v380 = ~(w1595 | w1596);
assign w1597 = v380;
assign v381 = ~(pi11 | w1597);
assign w1598 = v381;
assign w1599 = pi11 & w1597;
assign w1600 = ~w1541 & w2286;
assign v382 = ~(w1593 | w1600);
assign w1601 = v382;
assign v383 = ~(w1565 | w1601);
assign w1602 = v383;
assign w1603 = w1586 & w1602;
assign w1604 = (w1603 & w1557) | (w1603 & w2287) | (w1557 & w2287);
assign w1605 = ~w1499 & w1541;
assign v384 = ~(w1477 | w1500);
assign w1606 = v384;
assign w1607 = w1495 & w1606;
assign w1608 = w1495 & w2669;
assign w1609 = w1426 & w1608;
assign w1610 = w1426 & w1468;
assign w1611 = ~w1495 & w3093;
assign w1612 = (w1606 & w1495) | (w1606 & w3094) | (w1495 & w3094);
assign v385 = ~(w1611 | w1612);
assign w1613 = v385;
assign w1614 = (w1613 & ~w1426) | (w1613 & w3095) | (~w1426 & w3095);
assign w1615 = (w3096 & w3888) | (w3096 & w3889) | (w3888 & w3889);
assign v386 = ~(w1605 | w1615);
assign w1616 = v386;
assign w1617 = ~w1615 & w3890;
assign w1618 = (~w1500 & ~w1485) | (~w1500 & w2671) | (~w1485 & w2671);
assign v387 = ~(w1449 | w1497);
assign w1619 = v387;
assign w1620 = ~w1618 & w1619;
assign w1621 = w1618 & ~w1619;
assign v388 = ~(w1620 | w1621);
assign w1622 = v388;
assign w1623 = w1426 & w3097;
assign w1624 = ~w1607 & w1622;
assign w1625 = w1607 & ~w1622;
assign v389 = ~(w1624 | w1625);
assign w1626 = v389;
assign v390 = ~(w1609 | w1626);
assign w1627 = v390;
assign w1628 = ~w1627 & w3891;
assign w1629 = (~pi21 & ~w2288) | (~pi21 & w3098) | (~w2288 & w3098);
assign w1630 = ~w1628 & w1629;
assign w1631 = (~w1541 & w1627) | (~w1541 & w3892) | (w1627 & w3892);
assign w1632 = ~w1538 & w2289;
assign w1633 = (pi21 & ~w2289) | (pi21 & w3099) | (~w2289 & w3099);
assign w1634 = ~w1631 & w1633;
assign v391 = ~(w1630 | w1634);
assign w1635 = v391;
assign w1636 = ~w1617 & w1635;
assign w1637 = ~w1538 & w2290;
assign w1638 = (~w1597 & w1538) | (~w1597 & w2291) | (w1538 & w2291);
assign v392 = ~(w1637 | w1638);
assign w1639 = v392;
assign w1640 = pi11 & w1639;
assign w1641 = (w2283 & w2672) | (w2283 & w2673) | (w2672 & w2673);
assign w1642 = pi13 & ~w1423;
assign w1643 = (~w2282 & w2674) | (~w2282 & w2675) | (w2674 & w2675);
assign v393 = ~(w1641 | w1643);
assign w1644 = v393;
assign w1645 = ~w1640 & w1644;
assign w1646 = w1586 & ~w1645;
assign w1647 = (w1495 & ~w1426) | (w1495 & w2499) | (~w1426 & w2499);
assign v394 = ~(w1466 | w1494);
assign w1648 = v394;
assign w1649 = (w1648 & w1426) | (w1648 & w2500) | (w1426 & w2500);
assign w1650 = ~w1541 & w2292;
assign w1651 = w1203 & ~w1480;
assign w1652 = ~w1203 & w1480;
assign v395 = ~(w1651 | w1652);
assign w1653 = v395;
assign w1654 = ~w1538 & w2293;
assign v396 = ~(w1650 | w1654);
assign w1655 = v396;
assign w1656 = (pi17 & w1650) | (pi17 & w2501) | (w1650 & w2501);
assign w1657 = (~pi17 & ~w2293) | (~pi17 & w2676) | (~w2293 & w2676);
assign w1658 = ~w1650 & w1657;
assign v397 = ~(w1426 | w1468);
assign w1659 = v397;
assign v398 = ~(w1610 | w1659);
assign w1660 = v398;
assign w1661 = ~w1541 & w1660;
assign w1662 = ~w1538 & w2294;
assign v399 = ~(w1661 | w1662);
assign w1663 = v399;
assign w1664 = ~w1661 & w2295;
assign v400 = ~(w1658 | w1664);
assign w1665 = v400;
assign w1666 = ~w1656 & w1665;
assign w1667 = ~w1646 & w1666;
assign w1668 = w1636 & w1667;
assign w1669 = ~w1604 & w1668;
assign w1670 = (~pi19 & w1615) | (~pi19 & w2677) | (w1615 & w2677);
assign v401 = ~(w1658 | w1670);
assign w1671 = v401;
assign w1672 = w1635 & w4156;
assign w1673 = ~w1437 & w1541;
assign v402 = ~(w1440 | w1497);
assign w1674 = v402;
assign w1675 = (~w1626 & w2502) | (~w1626 & w2503) | (w2502 & w2503);
assign w1676 = (~w1503 & ~w1426) | (~w1503 & w2678) | (~w1426 & w2678);
assign w1677 = w1538 & w1676;
assign w1678 = ~w1675 & w1677;
assign v403 = ~(w1673 | w1678);
assign w1679 = v403;
assign w1680 = (~pi23 & w1678) | (~pi23 & w2679) | (w1678 & w2679);
assign v404 = ~(w1630 | w1680);
assign w1681 = v404;
assign w1682 = (w1681 & ~w1636) | (w1681 & w2504) | (~w1636 & w2504);
assign v405 = ~(w1312 | w1328);
assign w1683 = v405;
assign w1684 = ~w1326 & w1683;
assign w1685 = (w1684 & w1489) | (w1684 & w2505) | (w1489 & w2505);
assign w1686 = (w1489 & w4095) | (w1489 & w4096) | (w4095 & w4096);
assign w1687 = (w1502 & w2680) | (w1502 & w2681) | (w2680 & w2681);
assign w1688 = w1326 & ~w1683;
assign w1689 = w1334 & ~w1688;
assign w1690 = (w1689 & w1489) | (w1689 & w2682) | (w1489 & w2682);
assign w1691 = ~w1685 & w1690;
assign w1692 = ~w1538 & w2296;
assign w1693 = (pi27 & ~w2296) | (pi27 & w2683) | (~w2296 & w2683);
assign w1694 = ~w1691 & w1693;
assign w1695 = (~w1691 & w3893) | (~w1691 & w3894) | (w3893 & w3894);
assign v406 = ~(w1691 | w1692);
assign w1696 = v406;
assign w1697 = (~pi27 & w1691) | (~pi27 & w3895) | (w1691 & w3895);
assign w1698 = ~w1489 & w2684;
assign v407 = ~(w1326 | w1504);
assign w1699 = v407;
assign w1700 = w1487 & w3102;
assign w1701 = w1426 & w1700;
assign w1702 = ~w1699 & w4348;
assign v408 = ~(w1701 | w1702);
assign w1703 = v408;
assign w1704 = ~w1541 & w1703;
assign w1705 = ~w1698 & w1704;
assign w1706 = ~w1538 & w2298;
assign w1707 = (~pi25 & ~w2298) | (~pi25 & w3103) | (~w2298 & w3103);
assign w1708 = ~w1705 & w1707;
assign w1709 = (w1686 & w1705) | (w1686 & w2507) | (w1705 & w2507);
assign w1710 = ~w1697 & w1709;
assign v409 = ~(w1695 | w1710);
assign w1711 = v409;
assign v410 = ~(w1 | w1337);
assign w1712 = v410;
assign w1713 = ~w1710 & w2299;
assign w1714 = w1682 & ~w1713;
assign w1715 = ~w1678 & w2685;
assign w1716 = (~w1706 & ~w1704) | (~w1706 & w2508) | (~w1704 & w2508);
assign w1717 = (~w2508 & w2686) | (~w2508 & w2687) | (w2686 & w2687);
assign v411 = ~(w1708 | w1717);
assign w1718 = v411;
assign v412 = ~(w1695 | w1715);
assign w1719 = v412;
assign w1720 = w1718 & w1719;
assign v413 = ~(w1711 | w1720);
assign w1721 = v413;
assign w1722 = ~pi04 & w1541;
assign v414 = ~(w1336 | w1513);
assign w1723 = v414;
assign w1724 = ~w1541 & w1723;
assign v415 = ~(w1722 | w1724);
assign w1725 = v415;
assign w1726 = w1712 & ~w1725;
assign w1727 = ~w1721 & w1726;
assign w1728 = (w1727 & w1669) | (w1727 & w3104) | (w1669 & w3104);
assign w1729 = (w2300 & w1669) | (w2300 & w3105) | (w1669 & w3105);
assign w1730 = ~pi05 & w1725;
assign w1731 = w1725 & w3106;
assign w1732 = w1720 & ~w1731;
assign w1733 = ~w1713 & w1730;
assign w1734 = (~w1669 & w3896) | (~w1669 & w3897) | (w3896 & w3897);
assign v416 = ~(w1729 | w1734);
assign w1735 = v416;
assign w1736 = w1682 & ~w1711;
assign w1737 = ~w1669 & w1736;
assign w1738 = (~w1721 & w1669) | (~w1721 & w2688) | (w1669 & w2688);
assign w1739 = ~pi00 & pi01;
assign w1740 = pi03 & w1739;
assign v417 = ~(pi03 | w1739);
assign w1741 = v417;
assign w1742 = (~pi02 & w1739) | (~pi02 & w3107) | (w1739 & w3107);
assign v418 = ~(w1740 | w1742);
assign w1743 = v418;
assign w1744 = (~w1669 & w3898) | (~w1669 & w3899) | (w3898 & w3899);
assign w1745 = ~pi01 & w1742;
assign v419 = ~(w2 | w1739);
assign w1746 = v419;
assign w1747 = (~pi02 & ~w1739) | (~pi02 & w3108) | (~w1739 & w3108);
assign v420 = ~(w1746 | w1747);
assign w1748 = v420;
assign v421 = ~(w1745 | w1748);
assign w1749 = v421;
assign w1750 = (w1669 & w3109) | (w1669 & w3110) | (w3109 & w3110);
assign v422 = ~(w1744 | w1750);
assign w1751 = v422;
assign w1752 = w1735 & w1751;
assign w1753 = (~w1669 & w3111) | (~w1669 & w3112) | (w3111 & w3112);
assign w1754 = (~w1669 & w4157) | (~w1669 & w4158) | (w4157 & w4158);
assign w1755 = ~w1753 & w1754;
assign w1756 = (~w1525 & w1541) | (~w1525 & w3113) | (w1541 & w3113);
assign v423 = ~(w1543 | w1756);
assign w1757 = v423;
assign w1758 = pi07 & w1757;
assign w1759 = pi09 & w1553;
assign w1760 = pi13 & w1639;
assign w1761 = pi11 & w1564;
assign v424 = ~(w1759 | w1760);
assign w1762 = v424;
assign w1763 = ~w1761 & w1762;
assign w1764 = w1762 & w3114;
assign w1765 = (~w1669 & w3900) | (~w1669 & w3901) | (w3900 & w3901);
assign w1766 = (w1765 & ~w1754) | (w1765 & w2303) | (~w1754 & w2303);
assign w1767 = ~w1752 & w1766;
assign w1768 = (w2517 & w2516) | (w2517 & ~w2301) | (w2516 & ~w2301);
assign w1769 = (~pi11 & ~w1639) | (~pi11 & w3115) | (~w1639 & w3115);
assign w1770 = (w2691 & w2690) | (w2691 & ~w2301) | (w2690 & ~w2301);
assign v425 = ~(pi07 | w1757);
assign w1771 = v425;
assign v426 = ~(pi09 | w1553);
assign w1772 = v426;
assign v427 = ~(w1771 | w1772);
assign w1773 = v427;
assign w1774 = w1763 & ~w1773;
assign w1775 = ~w1738 & w1774;
assign v428 = ~(w1770 | w1775);
assign w1776 = v428;
assign w1777 = ~w1767 & w1776;
assign v429 = ~(w1572 | w1574);
assign w1778 = v429;
assign w1779 = (w2519 & w2518) | (w2519 & ~w2301) | (w2518 & ~w2301);
assign w1780 = ~w1576 & w1644;
assign w1781 = (w1602 & w1557) | (w1602 & w2304) | (w1557 & w2304);
assign w1782 = (w2304 & w3116) | (w2304 & w3117) | (w3116 & w3117);
assign w1783 = ~w1640 & w1780;
assign w1784 = (~w2304 & w3902) | (~w2304 & w3903) | (w3902 & w3903);
assign v430 = ~(w1782 | w1784);
assign w1785 = v430;
assign w1786 = w1738 & w1785;
assign v431 = ~(w1779 | w1786);
assign w1787 = v431;
assign w1788 = ~w1786 & w2521;
assign w1789 = (~w1585 & w1784) | (~w1585 & w3118) | (w1784 & w3118);
assign w1790 = (~w2287 & w3904) | (~w2287 & w3905) | (w3904 & w3905);
assign w1791 = ~w1721 & w1790;
assign w1792 = ~w1737 & w3119;
assign w1793 = (w2523 & w2522) | (w2523 & ~w2301) | (w2522 & ~w2301);
assign v432 = ~(w1792 | w1793);
assign w1794 = v432;
assign w1795 = (pi17 & w1792) | (pi17 & w2305) | (w1792 & w2305);
assign v433 = ~(w1788 | w1795);
assign w1796 = v433;
assign w1797 = ~w1777 & w1796;
assign v434 = ~(w1752 | w1755);
assign w1798 = v434;
assign w1799 = w1517 & w1534;
assign v435 = ~(w1535 | w1799);
assign w1800 = v435;
assign w1801 = (w1669 & w3120) | (w1669 & w3121) | (w3120 & w3121);
assign w1802 = (~w1669 & w3906) | (~w1669 & w3907) | (w3906 & w3907);
assign v436 = ~(w1801 | w1802);
assign w1803 = v436;
assign w1804 = ~pi07 & w1803;
assign v437 = ~(w1545 | w1556);
assign w1805 = v437;
assign v438 = ~(w1557 | w1805);
assign w1806 = v438;
assign v439 = ~(pi09 | w1806);
assign w1807 = v439;
assign w1808 = (~w2528 & w3908) | (~w2528 & w3909) | (w3908 & w3909);
assign v440 = ~(w1569 | w1808);
assign w1809 = v440;
assign w1810 = ~pi11 & w1809;
assign v441 = ~(w1807 | w1810);
assign w1811 = v441;
assign w1812 = (~w1557 & w2529) | (~w1557 & w2530) | (w2529 & w2530);
assign v442 = ~(w1781 | w1812);
assign w1813 = v442;
assign v443 = ~(pi13 | w1813);
assign w1814 = v443;
assign w1815 = w1738 & ~w1814;
assign v444 = ~(pi13 | w1639);
assign w1816 = v444;
assign w1817 = (~w1669 & w3910) | (~w1669 & w3911) | (w3910 & w3911);
assign v445 = ~(w1815 | w1817);
assign w1818 = v445;
assign w1819 = (w1811 & w1815) | (w1811 & w2533) | (w1815 & w2533);
assign w1820 = ~w1804 & w1819;
assign w1821 = ~w1798 & w1820;
assign w1822 = pi11 & ~w1809;
assign w1823 = pi07 & ~w1800;
assign w1824 = (~w1823 & ~w1806) | (~w1823 & w3122) | (~w1806 & w3122);
assign w1825 = ~w1810 & w3912;
assign w1826 = pi13 & w1813;
assign w1827 = w2534 & w3913;
assign v446 = ~(w1818 | w1827);
assign w1828 = v446;
assign w1829 = w1796 & ~w1828;
assign w1830 = ~w1821 & w1829;
assign v447 = ~(w1797 | w1830);
assign w1831 = v447;
assign v448 = ~(w1669 | w1672);
assign w1832 = v448;
assign w1833 = w1738 & ~w1832;
assign v449 = ~(w1617 | w1670);
assign w1834 = v449;
assign w1835 = w1603 & ~w1658;
assign w1836 = ~w1569 & w1835;
assign w1837 = ~w1836 & w2307;
assign v450 = ~(w1680 | w1715);
assign w1838 = v450;
assign w1839 = ~w1711 & w3123;
assign v451 = ~(w1635 | w1670);
assign w1840 = v451;
assign w1841 = ~w1721 & w1840;
assign w1842 = ~w1839 & w1841;
assign w1843 = ~w1837 & w1842;
assign v452 = ~(w1833 | w1843);
assign w1844 = v452;
assign v453 = ~(w1631 | w1632);
assign w1845 = v453;
assign w1846 = (w2536 & w2535) | (w2536 & ~w2301) | (w2535 & ~w2301);
assign w1847 = (w2301 & w3124) | (w2301 & w3125) | (w3124 & w3125);
assign w1848 = w1844 & w1847;
assign w1849 = (w2538 & w2537) | (w2538 & ~w2301) | (w2537 & ~w2301);
assign w1850 = (~w1630 & ~w1636) | (~w1630 & w2539) | (~w1636 & w2539);
assign w1851 = w1711 & w1838;
assign w1852 = ~w1669 & w2540;
assign v454 = ~(w1721 | w1838);
assign w1853 = v454;
assign w1854 = (~w1853 & w1669) | (~w1853 & w3126) | (w1669 & w3126);
assign v455 = ~(w1852 | w1854);
assign w1855 = v455;
assign v456 = ~(w1849 | w1855);
assign w1856 = v456;
assign w1857 = (~pi25 & w1855) | (~pi25 & w2541) | (w1855 & w2541);
assign w1858 = ~w1855 & w2542;
assign v457 = ~(w1857 | w1858);
assign w1859 = v457;
assign w1860 = w1848 & w1859;
assign w1861 = (w2544 & w2543) | (w2544 & ~w2301) | (w2543 & ~w2301);
assign w1862 = ~w1672 & w2308;
assign w1863 = w1715 & w1718;
assign w1864 = (~w1863 & w1669) | (~w1863 & w2692) | (w1669 & w2692);
assign v458 = ~(w1694 | w1697);
assign w1865 = v458;
assign v459 = ~(w1717 | w1865);
assign w1866 = v459;
assign w1867 = w1711 & w1866;
assign w1868 = (w2545 & w1669) | (w2545 & w3127) | (w1669 & w3127);
assign w1869 = (w2546 & w1669) | (w2546 & w2693) | (w1669 & w2693);
assign w1870 = (w1865 & w1711) | (w1865 & w3128) | (w1711 & w3128);
assign w1871 = ~w1721 & w1870;
assign w1872 = w1871 & ~w1869;
assign v460 = ~(w1861 | w1868);
assign w1873 = v460;
assign w1874 = ~w1872 & w1873;
assign w1875 = (~pi29 & ~w1873) | (~pi29 & w2694) | (~w1873 & w2694);
assign w1876 = (w2548 & w2547) | (w2548 & ~w2301) | (w2547 & ~w2301);
assign w1877 = (w2696 & w2695) | (w2696 & ~w2301) | (w2695 & ~w2301);
assign v461 = ~(w1715 | w1718);
assign w1878 = v461;
assign w1879 = (w1878 & w1669) | (w1878 & w2549) | (w1669 & w2549);
assign w1880 = w1864 & ~w1879;
assign w1881 = ~w1710 & w3129;
assign w1882 = (w1881 & ~w1864) | (w1881 & w2550) | (~w1864 & w2550);
assign v462 = ~(w1877 | w1882);
assign w1883 = v462;
assign w1884 = ~w1857 & w1883;
assign w1885 = ~w1875 & w1884;
assign w1886 = ~w1860 & w1885;
assign w1887 = (w2552 & w2551) | (w2552 & ~w2301) | (w2551 & ~w2301);
assign w1888 = (~w1834 & w1836) | (~w1834 & w2309) | (w1836 & w2309);
assign v463 = ~(w1837 | w1888);
assign w1889 = v463;
assign w1890 = w1738 & ~w1889;
assign v464 = ~(w1887 | w1890);
assign w1891 = v464;
assign w1892 = ~w1890 & w2553;
assign w1893 = (~w1664 & ~w1665) | (~w1664 & w3914) | (~w1665 & w3914);
assign w1894 = ~w1604 & w2554;
assign w1895 = (~w1656 & w1836) | (~w1656 & w2310) | (w1836 & w2310);
assign v465 = ~(w1894 | w1895);
assign w1896 = v465;
assign w1897 = w1738 & ~w1896;
assign w1898 = (w2556 & w2555) | (w2556 & ~w2301) | (w2555 & ~w2301);
assign v466 = ~(w1897 | w1898);
assign w1899 = v466;
assign w1900 = (~pi19 & w1897) | (~pi19 & w2557) | (w1897 & w2557);
assign v467 = ~(w1892 | w1900);
assign w1901 = v467;
assign w1902 = ~w1792 & w2311;
assign w1903 = (~pi15 & w1786) | (~pi15 & w2558) | (w1786 & w2558);
assign v468 = ~(w1902 | w1903);
assign w1904 = v468;
assign v469 = ~(w1795 | w1904);
assign w1905 = v469;
assign w1906 = (w1901 & w1904) | (w1901 & w2697) | (w1904 & w2697);
assign w1907 = w1886 & w1906;
assign w1908 = w1831 & w1907;
assign w1909 = (pi21 & w1890) | (pi21 & w2559) | (w1890 & w2559);
assign w1910 = ~w1897 & w2560;
assign v470 = ~(w1909 | w1910);
assign w1911 = v470;
assign v471 = ~(w1848 | w1892);
assign w1912 = v471;
assign w1913 = ~w1911 & w1912;
assign w1914 = ~w1833 & w3915;
assign w1915 = (pi23 & ~w1844) | (pi23 & w2312) | (~w1844 & w2312);
assign w1916 = w1859 & ~w1915;
assign w1917 = ~w1913 & w1916;
assign w1918 = w1711 & ~w1880;
assign w1919 = (~w1876 & w1880) | (~w1876 & w3130) | (w1880 & w3130);
assign w1920 = ~w1918 & w2313;
assign w1921 = ~w1875 & w1920;
assign w1922 = w1873 & w2698;
assign w1923 = (~pi31 & ~w2698) | (~pi31 & w3131) | (~w2698 & w3131);
assign w1924 = ~w1921 & w1923;
assign w1925 = (w1924 & w1917) | (w1924 & w2561) | (w1917 & w2561);
assign w1926 = ~w1908 & w1925;
assign w1927 = ~w1857 & w2784;
assign w1928 = ~w1875 & w1901;
assign w1929 = ~w1860 & w1928;
assign w1930 = ~w1905 & w1927;
assign w1931 = w1929 & w1930;
assign w1932 = w1831 & w1931;
assign v472 = ~(w1920 | w1922);
assign w1933 = v472;
assign w1934 = (w1873 & w2699) | (w1873 & w2700) | (w2699 & w2700);
assign w1935 = (w1934 & w1920) | (w1934 & w3916) | (w1920 & w3916);
assign w1936 = (~w434 & w1738) | (~w434 & w3135) | (w1738 & w3135);
assign w1937 = w1884 & w2701;
assign w1938 = (~w1936 & w1933) | (~w1936 & w2315) | (w1933 & w2315);
assign w1939 = (w1938 & w1917) | (w1938 & w2562) | (w1917 & w2562);
assign w1940 = ~w1932 & w1939;
assign v473 = ~(w1926 | w1940);
assign w1941 = v473;
assign w1942 = (pi00 & w1941) | (pi00 & w2316) | (w1941 & w2316);
assign w1943 = w1739 & ~w1941;
assign v474 = ~(w1942 | w1943);
assign w1944 = v474;
assign v475 = ~(w1740 | w1741);
assign w1945 = v475;
assign w1946 = (pi02 & ~w1738) | (pi02 & w3136) | (~w1738 & w3136);
assign w1947 = w1738 & w0;
assign v476 = ~(w1946 | w1947);
assign w1948 = v476;
assign w1949 = ~w1941 & w2317;
assign w1950 = (~w1948 & w1941) | (~w1948 & w2318) | (w1941 & w2318);
assign v477 = ~(w1949 | w1950);
assign w1951 = v477;
assign w1952 = (~w1751 & w1755) | (~w1751 & w3137) | (w1755 & w3137);
assign w1953 = ~w1755 & w1752;
assign v478 = ~(w1952 | w1953);
assign w1954 = v478;
assign w1955 = ~w1941 & w1954;
assign v479 = ~(w1728 | w1753);
assign w1956 = v479;
assign w1957 = w1941 & w1956;
assign v480 = ~(w1955 | w1957);
assign w1958 = v480;
assign w1959 = pi07 & ~w1803;
assign v481 = ~(w1804 | w1959);
assign w1960 = v481;
assign w1961 = w1798 & ~w1960;
assign w1962 = ~w1798 & w1960;
assign v482 = ~(w1961 | w1962);
assign w1963 = v482;
assign v483 = ~(w1941 | w1963);
assign w1964 = v483;
assign w1965 = w1803 & w1941;
assign v484 = ~(w1964 | w1965);
assign w1966 = v484;
assign w1967 = ~w1721 & w3759;
assign w1968 = (~w1669 & w3917) | (~w1669 & w3918) | (w3917 & w3918);
assign v485 = ~(w1967 | w1968);
assign w1969 = v485;
assign w1970 = w1941 & ~w1969;
assign w1971 = w1798 & ~w1959;
assign w1972 = (pi09 & w1967) | (pi09 & w3138) | (w1967 & w3138);
assign w1973 = ~w1967 & w3139;
assign v486 = ~(w1972 | w1973);
assign w1974 = v486;
assign w1975 = ~w1804 & w1974;
assign w1976 = ~w1971 & w1975;
assign w1977 = (~w1804 & ~w1798) | (~w1804 & w3140) | (~w1798 & w3140);
assign v487 = ~(w1974 | w1977);
assign w1978 = v487;
assign v488 = ~(w1976 | w1978);
assign w1979 = v488;
assign w1980 = ~w1941 & w1979;
assign v489 = ~(w1970 | w1980);
assign w1981 = v489;
assign w1982 = w1738 & w1809;
assign v490 = ~(w1768 | w1982);
assign w1983 = v490;
assign w1984 = (~w1935 & w1917) | (~w1935 & w2566) | (w1917 & w2566);
assign w1985 = ~w1932 & w1984;
assign w1986 = (~w1738 & w3141) | (~w1738 & w3142) | (w3141 & w3142);
assign w1987 = ~w1976 & w2319;
assign w1988 = (~w1738 & w3143) | (~w1738 & w3144) | (w3143 & w3144);
assign w1989 = (w1988 & w1976) | (w1988 & w2320) | (w1976 & w2320);
assign v491 = ~(w1987 | w1989);
assign w1990 = v491;
assign w1991 = ~w1932 & w3145;
assign w1992 = (~w1921 & w1917) | (~w1921 & w2567) | (w1917 & w2567);
assign w1993 = ~w1908 & w1992;
assign w1994 = ~w1976 & w2702;
assign w1995 = (w3131 & w3919) | (w3131 & w3920) | (w3919 & w3920);
assign w1996 = (w1995 & w1976) | (w1995 & w2703) | (w1976 & w2703);
assign v492 = ~(w1994 | w1996);
assign w1997 = v492;
assign w1998 = ~w1908 & w3146;
assign v493 = ~(w1991 | w1998);
assign w1999 = v493;
assign w2000 = ~w1983 & w1999;
assign w2001 = w1983 & ~w1999;
assign v494 = ~(w2000 | w2001);
assign w2002 = v494;
assign v495 = ~(w603 | w752);
assign w2003 = v495;
assign w2004 = w1738 & ~w1813;
assign v496 = ~(w1639 | w1738);
assign w2005 = v496;
assign v497 = ~(w2004 | w2005);
assign w2006 = v497;
assign w2007 = w1941 & ~w2006;
assign w2008 = pi13 & w2006;
assign v498 = ~(w1818 | w2008);
assign w2009 = v498;
assign w2010 = (~pi11 & w1982) | (~pi11 & w3147) | (w1982 & w3147);
assign w2011 = ~w1982 & w3148;
assign w2012 = (~w2010 & w1976) | (~w2010 & w3149) | (w1976 & w3149);
assign w2013 = (~w1976 & w4159) | (~w1976 & w4160) | (w4159 & w4160);
assign w2014 = (w1976 & w3150) | (w1976 & w3151) | (w3150 & w3151);
assign w2015 = ~w1941 & w2322;
assign v499 = ~(w2007 | w2015);
assign w2016 = v499;
assign w2017 = w1787 & w1941;
assign v500 = ~(w1788 | w1903);
assign w2018 = v500;
assign w2019 = ~w2012 & w3152;
assign w2020 = w1818 & ~w2018;
assign w2021 = w1776 & ~w1903;
assign w2022 = (~w1788 & w1767) | (~w1788 & w2704) | (w1767 & w2704);
assign w2023 = (~w1788 & w1827) | (~w1788 & w3153) | (w1827 & w3153);
assign w2024 = ~w1821 & w2023;
assign v501 = ~(w2022 | w2024);
assign w2025 = v501;
assign w2026 = (~w2020 & ~w2025) | (~w2020 & w3154) | (~w2025 & w3154);
assign w2027 = ~w1941 & w3155;
assign v502 = ~(w2017 | w2027);
assign w2028 = v502;
assign w2029 = (w3131 & w3921) | (w3131 & w3922) | (w3921 & w3922);
assign w2030 = ~w2024 & w2705;
assign w2031 = (w3131 & w3923) | (w3131 & w3924) | (w3923 & w3924);
assign w2032 = (w2031 & w2024) | (w2031 & w2706) | (w2024 & w2706);
assign v503 = ~(w2030 | w2032);
assign w2033 = v503;
assign w2034 = w1993 & ~w2033;
assign w2035 = (~w1738 & w3156) | (~w1738 & w3157) | (w3156 & w3157);
assign w2036 = ~w2024 & w2707;
assign w2037 = (~w1738 & w3158) | (~w1738 & w3159) | (w3158 & w3159);
assign w2038 = (w2037 & w2024) | (w2037 & w2708) | (w2024 & w2708);
assign v504 = ~(w2036 | w2038);
assign w2039 = v504;
assign w2040 = w1985 & ~w2039;
assign v505 = ~(w2034 | w2040);
assign w2041 = v505;
assign w2042 = ~w1794 & w2041;
assign w2043 = w1794 & ~w2041;
assign v506 = ~(w2042 | w2043);
assign w2044 = v506;
assign w2045 = w1899 & w1941;
assign v507 = ~(w1900 | w1910);
assign w2046 = v507;
assign w2047 = ~w1830 & w3161;
assign w2048 = (~w2046 & ~w3160) | (~w2046 & w3925) | (~w3160 & w3925);
assign v508 = ~(w2047 | w2048);
assign w2049 = v508;
assign w2050 = ~w1941 & w2049;
assign v509 = ~(w2045 | w2050);
assign w2051 = v509;
assign v510 = ~(w1892 | w1911);
assign w2052 = v510;
assign w2053 = (w1831 & w3510) | (w1831 & w3162) | (w3510 & w3162);
assign v511 = ~(w1892 | w1909);
assign w2054 = v511;
assign v512 = ~(w1910 | w2054);
assign w2055 = v512;
assign w2056 = (w2055 & ~w3161) | (w2055 & w3926) | (~w3161 & w3926);
assign v513 = ~(w2053 | w2056);
assign w2057 = v513;
assign v514 = ~(w1941 | w2057);
assign w2058 = v514;
assign w2059 = w1891 & w1941;
assign v515 = ~(w2058 | w2059);
assign w2060 = v515;
assign w2061 = w1914 & w1941;
assign v516 = ~(w1848 | w1915);
assign w2062 = v516;
assign w2063 = (w1831 & w3163) | (w1831 & w3164) | (w3163 & w3164);
assign w2064 = (~w1831 & w3165) | (~w1831 & w3166) | (w3165 & w3166);
assign w2065 = ~w1941 & w2324;
assign v517 = ~(w2061 | w2065);
assign w2066 = v517;
assign w2067 = ~w1856 & w1941;
assign v518 = ~(w1848 | w1859);
assign w2068 = v518;
assign w2069 = ~w2064 & w2068;
assign w2070 = (w1917 & ~w1831) | (w1917 & w3167) | (~w1831 & w3167);
assign w2071 = ~w1941 & w3168;
assign v519 = ~(w2067 | w2071);
assign w2072 = v519;
assign w2073 = (~w67 & w33) | (~w67 & w3169) | (w33 & w3169);
assign w2074 = w68 & ~w2073;
assign w2075 = w1919 & w1941;
assign w2076 = (~w1857 & ~w1859) | (~w1857 & w2326) | (~w1859 & w2326);
assign w2077 = w1906 & w2076;
assign w2078 = w1831 & w2077;
assign w2079 = (~w1857 & w1913) | (~w1857 & w2568) | (w1913 & w2568);
assign w2080 = w1883 & ~w1920;
assign w2081 = (w2080 & w2078) | (w2080 & w2327) | (w2078 & w2327);
assign w2082 = (w4065 & w4161) | (w4065 & w4162) | (w4161 & w4162);
assign w2083 = ~w1941 & w3170;
assign v520 = ~(w2075 | w2083);
assign w2084 = v520;
assign w2085 = pi01 & ~pi28;
assign w2086 = ~w7 & w25;
assign w2087 = ~w2085 & w2086;
assign w2088 = w3751 & w2087;
assign w2089 = w1874 & w1941;
assign v521 = ~(w1875 | w1922);
assign w2090 = v521;
assign w2091 = (w2078 & w3171) | (w2078 & w3172) | (w3171 & w3172);
assign w2092 = w1920 & ~w2090;
assign w2093 = ~w1920 & w2090;
assign v522 = ~(w2092 | w2093);
assign w2094 = v522;
assign w2095 = ~w2080 & w2094;
assign w2096 = ~w2079 & w2094;
assign w2097 = (~w2095 & w2078) | (~w2095 & w2785) | (w2078 & w2785);
assign w2098 = ~w1941 & w3173;
assign v523 = ~(w2089 | w2098);
assign w2099 = v523;
assign w2100 = pi01 & ~pi30;
assign v524 = ~(pi03 | pi05);
assign w2101 = v524;
assign w2102 = ~w2100 & w2101;
assign w2103 = w52 & w2102;
assign w2104 = ~w1932 & w3174;
assign v525 = ~(w1936 | w2104);
assign w2105 = v525;
assign w2106 = w7 & pi28;
assign w2107 = ~pi03 & pi28;
assign w2108 = pi03 & pi05;
assign w2109 = w12 & ~w36;
assign w2110 = pi26 & w53;
assign w2111 = ~w9 & w2328;
assign v526 = ~(w82 | w49);
assign w2112 = v526;
assign w2113 = (pi28 & ~w13) | (pi28 & w2106) | (~w13 & w2106);
assign v527 = ~(w63 | w91);
assign w2114 = v527;
assign w2115 = (w23 & w2329) | (w23 & w2330) | (w2329 & w2330);
assign w2116 = w101 & w103;
assign w2117 = (w100 & w3927) | (w100 & w3928) | (w3927 & w3928);
assign w2118 = ~w100 & w3175;
assign w2119 = (w42 & w2709) | (w42 & w2710) | (w2709 & w2710);
assign w2120 = w132 & w135;
assign w2121 = ~w153 & w2332;
assign w2122 = w156 & w160;
assign w2123 = ~w153 & w2711;
assign w2124 = ~w137 & w144;
assign w2125 = (~w244 & w241) | (~w244 & w2829) | (w241 & w2829);
assign v528 = ~(w250 | w252);
assign w2126 = v528;
assign w2127 = (w263 & ~w171) | (w263 & w2569) | (~w171 & w2569);
assign w2128 = (w270 & ~w264) | (w270 & w2889) | (~w264 & w2889);
assign w2129 = w264 & w2890;
assign w2130 = (w3701 & ~w171) | (w3701 & w2570) | (~w171 & w2570);
assign w2131 = (w279 & ~w274) | (w279 & w2786) | (~w274 & w2786);
assign w2132 = (w268 & ~w264) | (w268 & w3176) | (~w264 & w3176);
assign w2133 = w264 & w2787;
assign w2134 = (w269 & ~w264) | (w269 & w2788) | (~w264 & w2788);
assign w2135 = (pi07 & w241) | (pi07 & w2789) | (w241 & w2789);
assign w2136 = (~w267 & ~w264) | (~w267 & w2790) | (~w264 & w2790);
assign w2137 = w264 & w2791;
assign v529 = ~(w313 | w314);
assign w2138 = v529;
assign w2139 = (w2721 & w230) | (w2721 & w2333) | (w230 & w2333);
assign w2140 = (w319 & w241) | (w319 & w2830) | (w241 & w2830);
assign w2141 = (w325 & w241) | (w325 & w2831) | (w241 & w2831);
assign w2142 = (~w337 & ~w330) | (~w337 & w2773) | (~w330 & w2773);
assign w2143 = w338 & w340;
assign w2144 = ~w354 & w363;
assign w2145 = w354 & ~w363;
assign w2146 = ~w354 & w368;
assign w2147 = ~w294 & w2792;
assign v530 = ~(w322 | w416);
assign w2148 = v530;
assign w2149 = w322 & w416;
assign w2150 = (pi16 & w439) | (pi16 & w2571) | (w439 & w2571);
assign w2151 = (w342 & w384) | (w342 & w2334) | (w384 & w2334);
assign w2152 = ~w439 & w2335;
assign w2153 = (~w467 & w439) | (~w467 & w2336) | (w439 & w2336);
assign w2154 = ~w439 & w2572;
assign w2155 = (w492 & w439) | (w492 & w3177) | (w439 & w3177);
assign w2156 = (w502 & w439) | (w502 & w3178) | (w439 & w3178);
assign w2157 = (w505 & w439) | (w505 & w3179) | (w439 & w3179);
assign w2158 = w401 & ~w411;
assign w2159 = (~w523 & w439) | (~w523 & w2337) | (w439 & w2337);
assign w2160 = ~w439 & w2338;
assign w2161 = (w534 & w439) | (w534 & w3180) | (w439 & w3180);
assign w2162 = (w410 & w439) | (w410 & w2339) | (w439 & w2339);
assign w2163 = w513 & ~w556;
assign v531 = ~(w549 | w547);
assign w2164 = v531;
assign w2165 = (~w2164 & w2793) | (~w2164 & w2794) | (w2793 & w2794);
assign w2166 = w560 & w567;
assign v532 = ~(w560 | w526);
assign w2167 = v532;
assign w2168 = (w2795 & w3768) | (w2795 & w2164) | (w3768 & w2164);
assign v533 = ~(w583 | w582);
assign w2169 = v533;
assign w2170 = (pi15 & w2340) | (pi15 & w593) | (w2340 & w593);
assign w2171 = w513 & ~w593;
assign w2172 = (w2341 & w566) | (w2341 & w3181) | (w566 & w3181);
assign w2173 = (w2342 & w566) | (w2342 & w3182) | (w566 & w3182);
assign w2174 = w728 & w2891;
assign w2175 = (w742 & w3183) | (w742 & w3184) | (w3183 & w3184);
assign v534 = ~(w742 | w691);
assign w2176 = v534;
assign w2177 = (~w2176 & w3186) | (~w2176 & w3187) | (w3186 & w3187);
assign v535 = ~(w765 | w766);
assign w2178 = v535;
assign w2179 = (w742 & w3188) | (w742 & w3189) | (w3188 & w3189);
assign w2180 = (~w742 & w3190) | (~w742 & w3191) | (w3190 & w3191);
assign w2181 = (~w572 & ~w589) | (~w572 & w3192) | (~w589 & w3192);
assign w2182 = (w716 & w4163) | (w716 & w4164) | (w4163 & w4164);
assign v536 = ~(w798 | w796);
assign w2183 = v536;
assign w2184 = w798 & w796;
assign w2185 = (w809 & w3195) | (w809 & w572) | (w3195 & w572);
assign w2186 = w798 & w822;
assign v537 = ~(w798 | w822);
assign w2187 = v537;
assign w2188 = w842 & w845;
assign v538 = ~(w842 | w845);
assign w2189 = v538;
assign w2190 = ~w603 & w3196;
assign w2191 = (w603 & w855) | (w603 & w3197) | (w855 & w3197);
assign w2192 = pi13 & w757;
assign w2193 = ~w731 & w874;
assign w2194 = w802 & w860;
assign w2195 = ~w760 & w2573;
assign w2196 = ~w875 & w964;
assign v539 = ~(w767 | w772);
assign w2197 = v539;
assign w2198 = w867 & w848;
assign w2199 = ~w936 & w2894;
assign w2200 = (pi11 & w936) | (pi11 & w2895) | (w936 & w2895);
assign w2201 = ~w1045 & w991;
assign w2202 = (~w787 & ~w964) | (~w787 & w2574) | (~w964 & w2574);
assign w2203 = (w971 & ~w964) | (w971 & w2575) | (~w964 & w2575);
assign w2204 = ~w1067 & w1073;
assign w2205 = ~w1046 & w1078;
assign w2206 = ~w991 & w1077;
assign w2207 = ~w991 & w1093;
assign w2208 = ~w991 & w1104;
assign w2209 = ~w1049 & w3198;
assign w2210 = (~w4147 & w1139) | (~w4147 & w3200) | (w1139 & w3200);
assign w2211 = w1131 & w1146;
assign w2212 = w4147 & ~w1161;
assign w2213 = (w4147 & w1037) | (w4147 & w3201) | (w1037 & w3201);
assign v540 = ~(w962 | w1017);
assign w2214 = v540;
assign w2215 = (w2577 & w2576) | (w2577 & w1117) | (w2576 & w1117);
assign w2216 = (~w1176 & w1037) | (~w1176 & w3929) | (w1037 & w3929);
assign w2217 = (~w4147 & ~w1139) | (~w4147 & w3202) | (~w1139 & w3202);
assign w2218 = (w1117 & w3769) | (w1117 & w3770) | (w3769 & w3770);
assign w2219 = (~w1035 & w3203) | (~w1035 & w3204) | (w3203 & w3204);
assign w2220 = (w4147 & w959) | (w4147 & w3930) | (w959 & w3930);
assign w2221 = w1209 & w1212;
assign v541 = ~(w1209 | w1212);
assign w2222 = v541;
assign w2223 = ~w997 & w3205;
assign v542 = ~(pi17 | w1217);
assign w2224 = v542;
assign w2225 = w1029 & w1224;
assign v543 = ~(w1029 | w1224);
assign w2226 = v543;
assign w2227 = ~w989 & w3206;
assign w2228 = (w1117 & w4066) | (w1117 & w4067) | (w4066 & w4067);
assign w2229 = (w1238 & w997) | (w1238 & w3931) | (w997 & w3931);
assign v544 = ~(w1246 | w1245);
assign w2230 = v544;
assign w2231 = w1254 & ~w1235;
assign w2232 = (w1117 & w4068) | (w1117 & w4069) | (w4068 & w4069);
assign w2233 = (w3207 & ~w1051) | (w3207 & w1264) | (~w1051 & w1264);
assign w2234 = ~w1225 & w1267;
assign w2235 = ~w1046 & w1270;
assign v545 = ~(w1234 | w1273);
assign w2236 = v545;
assign w2237 = (w3039 & w3933) | (w3039 & w3934) | (w3933 & w3934);
assign w2238 = (~w2201 & w3209) | (~w2201 & w3210) | (w3209 & w3210);
assign w2239 = w1298 & w3935;
assign w2240 = w1300 & w1307;
assign w2241 = (~pi25 & w1300) | (~pi25 & w3211) | (w1300 & w3211);
assign w2242 = w1295 & w2343;
assign v546 = ~(w1317 | w1259);
assign w2243 = v546;
assign w2244 = ~w1263 & w2344;
assign w2245 = w1332 & w1314;
assign w2246 = w1298 & w2713;
assign w2247 = pi06 & w3760;
assign w2248 = w1298 & w2714;
assign v547 = ~(w1342 | w1343);
assign w2249 = v547;
assign w2250 = w1298 & w2715;
assign w2251 = (w2250 & w2832) | (w2250 & w2833) | (w2832 & w2833);
assign w2252 = (w4037 & w4070) | (w4037 & w4071) | (w4070 & w4071);
assign w2253 = (w1368 & ~w1295) | (w1368 & w2345) | (~w1295 & w2345);
assign w2254 = w1295 & w2346;
assign v548 = ~(w1300 | w1381);
assign w2255 = v548;
assign w2256 = w1295 & w2347;
assign w2257 = w1298 & w3936;
assign w2258 = (w1372 & ~w1298) | (w1372 & w3937) | (~w1298 & w3937);
assign w2259 = ~w1300 & w1400;
assign w2260 = w1295 & w2348;
assign w2261 = w1405 & ~w1388;
assign v549 = ~(w1409 | w1423);
assign w2262 = v549;
assign w2263 = w1294 & ~w1258;
assign w2264 = (w3858 & w4165) | (w3858 & w4166) | (w4165 & w4166);
assign w2265 = ~w1321 & w2350;
assign w2266 = (pi19 & w1444) | (pi19 & w3212) | (w1444 & w3212);
assign w2267 = (~w1460 & ~w1298) | (~w1460 & w3938) | (~w1298 & w3938);
assign w2268 = w1298 & w3939;
assign w2269 = ~w1469 & w3761;
assign w2270 = w1446 & ~pi19;
assign w2271 = w1295 & w2579;
assign w2272 = (w1289 & w2580) | (w1289 & w2581) | (w2580 & w2581);
assign w2273 = ~w1450 & w1505;
assign w2274 = ~w1313 & w3213;
assign w2275 = (pi05 & w1313) | (pi05 & w3214) | (w1313 & w3214);
assign w2276 = w1540 & w1542;
assign w2277 = w1529 & ~w1522;
assign w2278 = w1540 & ~w1547;
assign v550 = ~(w1540 | w1551);
assign w2279 = v550;
assign w2280 = w1540 & w1561;
assign v551 = ~(w1540 | w1397);
assign w2281 = v551;
assign w2282 = w1540 & w1571;
assign w2283 = w1540 & w1573;
assign w2284 = w1579 & w1582;
assign v552 = ~(w1579 | w1582);
assign w2285 = v552;
assign v553 = ~(w1598 | w1599);
assign w2286 = v553;
assign w2287 = ~w1568 & w1603;
assign w2288 = ~w1540 & w1448;
assign v554 = ~(w1540 | w1448);
assign w2289 = v554;
assign v555 = ~(w1540 | w1589);
assign w2290 = v555;
assign w2291 = w1540 & ~w1597;
assign v556 = ~(w1647 | w1649);
assign w2292 = v556;
assign w2293 = ~w1540 & w1653;
assign w2294 = ~w1540 & w1465;
assign w2295 = (pi15 & ~w2294) | (pi15 & w2716) | (~w2294 & w2716);
assign w2296 = ~w1540 & w1327;
assign w2297 = (~w1439 & ~w1440) | (~w1439 & w3215) | (~w1440 & w3215);
assign v557 = ~(w1540 | w1325);
assign w2298 = v557;
assign w2299 = ~w1695 & w1712;
assign w2300 = ~w1721 & w2352;
assign w2301 = w1669 & ~w1721;
assign w2302 = (w1725 & w1721) | (w1725 & w2353) | (w1721 & w2353);
assign w2303 = w1753 & w1765;
assign w2304 = ~w1568 & w1602;
assign w2305 = (w2583 & w2582) | (w2583 & ~w2301) | (w2582 & ~w2301);
assign w2306 = (~w1565 & ~w1567) | (~w1565 & w2355) | (~w1567 & w2355);
assign w2307 = (~w1646 & w4337) | (~w1646 & w4338) | (w4337 & w4338);
assign w2308 = w1681 & w1718;
assign w2309 = (w2357 & w1646) | (w2357 & w4339) | (w1646 & w4339);
assign w2310 = (w2358 & w1646) | (w2358 & w3216) | (w1646 & w3216);
assign w2311 = (w1669 & w3940) | (w1669 & w3941) | (w3940 & w3941);
assign w2312 = (~w2301 & w3217) | (~w2301 & w3218) | (w3217 & w3218);
assign w2313 = ~w1876 & pi27;
assign w2314 = pi29 & pi31;
assign w2315 = (~w2700 & w3219) | (~w2700 & w3220) | (w3219 & w3220);
assign w2316 = ~pi01 & pi00;
assign w2317 = w1945 & w1948;
assign v558 = ~(w1945 | w1948);
assign w2318 = v558;
assign w2319 = ~w1972 & w1986;
assign w2320 = w1972 & w1988;
assign v559 = ~(w1972 | w2011);
assign w2321 = v559;
assign v560 = ~(w2013 | w2014);
assign w2322 = v560;
assign w2323 = ~w1905 & w2046;
assign v561 = ~(w2063 | w2064);
assign w2324 = v561;
assign w2325 = w1906 & ~w1860;
assign v562 = ~(w1848 | w1857);
assign w2326 = v562;
assign w2327 = w2079 & w2080;
assign v563 = ~(w5 | w47);
assign w2328 = v563;
assign w2329 = w99 & w47;
assign w2330 = w99 & ~w2111;
assign w2331 = (w42 & w3221) | (w42 & w3222) | (w3221 & w3222);
assign w2332 = w72 & w147;
assign w2333 = w223 & w3224;
assign w2334 = ~w396 & w342;
assign w2335 = (w146 & w3226) | (w146 & w3227) | (w3226 & w3227);
assign w2336 = (~w415 & ~w466) | (~w415 & w3228) | (~w466 & w3228);
assign w2337 = (~w415 & w420) | (~w415 & w3229) | (w420 & w3229);
assign w2338 = w415 & ~w527;
assign w2339 = ~w415 & w410;
assign w2340 = ~w545 & w3230;
assign v564 = ~(w653 | pi07);
assign w2341 = v564;
assign w2342 = (~pi15 & w545) | (~pi15 & w3231) | (w545 & w3231);
assign w2343 = (~w1233 & ~w1298) | (~w1233 & w3944) | (~w1298 & w3944);
assign w2344 = ~w1300 & w3234;
assign w2345 = w1299 & w1368;
assign w2346 = (w1375 & ~w1298) | (w1375 & w3945) | (~w1298 & w3945);
assign w2347 = (~w1386 & ~w1298) | (~w1386 & w3946) | (~w1298 & w3946);
assign w2348 = (w1403 & ~w1298) | (w1403 & w3947) | (~w1298 & w3947);
assign w2349 = (w2826 & w3948) | (w2826 & w3949) | (w3948 & w3949);
assign w2350 = w3236 & ~w1295;
assign w2351 = w1608 & w1620;
assign w2352 = ~w1725 & w3237;
assign w2353 = ~w1712 & w1725;
assign w2354 = w1663 & pi17;
assign w2355 = w1554 & ~w1565;
assign w2356 = ~w1617 & w4167;
assign w2357 = (~w1658 & w1617) | (~w1658 & w4168) | (w1617 & w4168);
assign v565 = ~(w1658 | w1656);
assign w2358 = v565;
assign w2359 = w71 & w28;
assign w2360 = ~w2110 & w75;
assign w2361 = w23 & w3238;
assign w2362 = w116 & w2836;
assign w2363 = (w2837 & w2838) | (w2837 & w116) | (w2838 & w116);
assign w2364 = ~w179 & w213;
assign w2365 = w137 & w147;
assign w2366 = ~w173 & w3950;
assign w2367 = (w144 & w141) | (w144 & w2720) | (w141 & w2720);
assign w2368 = ~w226 & w232;
assign w2369 = (~pi09 & w173) | (~pi09 & w3951) | (w173 & w3951);
assign w2370 = (w32 & w234) | (w32 & w2721) | (w234 & w2721);
assign v566 = ~(w206 | w234);
assign w2371 = v566;
assign w2372 = (w282 & w234) | (w282 & w2723) | (w234 & w2723);
assign w2373 = (~pi07 & ~w267) | (~pi07 & w25) | (~w267 & w25);
assign v567 = ~(pi07 | w233);
assign w2374 = v567;
assign w2375 = w172 & w311;
assign w2376 = w320 & w324;
assign w2377 = (~w2774 & w3239) | (~w2774 & w3240) | (w3239 & w3240);
assign w2378 = (w344 & ~w338) | (w344 & w2377) | (~w338 & w2377);
assign w2379 = w350 & w4349;
assign w2380 = (w350 & ~w338) | (w350 & w2379) | (~w338 & w2379);
assign w2381 = ~w355 & w2144;
assign w2382 = w2145 & ~w363;
assign w2383 = (~w363 & w2145) | (~w363 & w355) | (w2145 & w355);
assign w2384 = ~w355 & w2146;
assign w2385 = w354 & w361;
assign w2386 = (w361 & w2385) | (w361 & w355) | (w2385 & w355);
assign w2387 = w380 & w340;
assign w2388 = w338 & w2387;
assign w2389 = ~w373 & w2839;
assign w2390 = w374 & ~w2143;
assign w2391 = w378 & w340;
assign w2392 = w338 & w2391;
assign w2393 = ~w422 & w340;
assign w2394 = w338 & w2393;
assign w2395 = w422 & w340;
assign w2396 = w338 & w2395;
assign w2397 = (w323 & w3241) | (w323 & w3242) | (w3241 & w3242);
assign w2398 = (w323 & w3243) | (w323 & w3244) | (w3243 & w3244);
assign w2399 = ~w323 & w3952;
assign w2400 = w447 & w4350;
assign w2401 = w459 & w452;
assign w2402 = ~w439 & w3953;
assign v568 = ~(w459 | w452);
assign w2403 = v568;
assign w2404 = (~w459 & w439) | (~w459 & w3954) | (w439 & w3954);
assign w2405 = (w439 & w3245) | (w439 & w3246) | (w3245 & w3246);
assign w2406 = ~w456 & w3247;
assign w2407 = ~w439 & w3248;
assign w2408 = w456 & w3249;
assign w2409 = (w479 & w439) | (w479 & w3250) | (w439 & w3250);
assign w2410 = w440 & w497;
assign w2411 = w440 & w507;
assign w2412 = ~w515 & w2840;
assign w2413 = (~w529 & w2585) | (~w529 & w2586) | (w2585 & w2586);
assign v569 = ~(w396 | w401);
assign w2414 = v569;
assign w2415 = w549 & w533;
assign w2416 = w510 & ~w547;
assign w2417 = w2801 & w3251;
assign w2418 = w570 & ~w567;
assign w2419 = (w570 & ~w558) | (w570 & w3252) | (~w558 & w3252);
assign w2420 = w2801 & w3253;
assign w2421 = w558 & w3955;
assign v570 = ~(w578 | w580);
assign w2422 = v570;
assign w2423 = (~w552 & w3254) | (~w552 & w3255) | (w3254 & w3255);
assign w2424 = w531 & w610;
assign w2425 = ~w566 & w3256;
assign w2426 = w615 & w551;
assign w2427 = ~w608 & w617;
assign w2428 = (w625 & w566) | (w625 & w3257) | (w566 & w3257);
assign w2429 = w625 & ~w551;
assign w2430 = ~w566 & w3258;
assign w2431 = ~w632 & w551;
assign v571 = ~(w608 | w612);
assign w2432 = v571;
assign w2433 = ~w566 & w2796;
assign w2434 = w2415 & w2797;
assign w2435 = (pi11 & w656) | (pi11 & w2587) | (w656 & w2587);
assign w2436 = ~w484 & w510;
assign w2437 = ~w671 & w2588;
assign w2438 = (w680 & w671) | (w680 & w696) | (w671 & w696);
assign w2439 = ~w668 & w692;
assign w2440 = ~w673 & w694;
assign w2441 = w673 & w696;
assign w2442 = w660 & ~w698;
assign w2443 = (w2589 & w670) | (w2589 & w3259) | (w670 & w3259);
assign w2444 = ~w673 & w704;
assign w2445 = ~w701 & w715;
assign v572 = ~(w701 | w707);
assign w2446 = v572;
assign w2447 = ~w656 & w3260;
assign w2448 = w619 & ~pi11;
assign v573 = ~(w734 | w683);
assign w2449 = v573;
assign w2450 = (w792 & ~w778) | (w792 & w3261) | (~w778 & w3261);
assign w2451 = (~w2439 & w3262) | (~w2439 & w3263) | (w3262 & w3263);
assign w2452 = w724 & w4169;
assign w2453 = (~w2450 & w2724) | (~w2450 & w2725) | (w2724 & w2725);
assign w2454 = (w2450 & w2726) | (w2450 & w2727) | (w2726 & w2727);
assign w2455 = (~w787 & ~w778) | (~w787 & w3264) | (~w778 & w3264);
assign w2456 = (~w2455 & w2728) | (~w2455 & w2729) | (w2728 & w2729);
assign w2457 = w889 & w899;
assign w2458 = w778 & w3956;
assign w2459 = (~w912 & ~w2458) | (~w912 & w3265) | (~w2458 & w3265);
assign w2460 = (~w2450 & w2730) | (~w2450 & w2731) | (w2730 & w2731);
assign w2461 = (w2450 & w2732) | (w2450 & w2733) | (w2732 & w2733);
assign w2462 = (w2455 & w2734) | (w2455 & w2735) | (w2734 & w2735);
assign w2463 = (~w2455 & w2736) | (~w2455 & w2737) | (w2736 & w2737);
assign w2464 = w889 & ~w938;
assign w2465 = (~w2455 & w2738) | (~w2455 & w2739) | (w2738 & w2739);
assign w2466 = (~w2455 & w2740) | (~w2455 & w2741) | (w2740 & w2741);
assign w2467 = (~pi11 & w888) | (~pi11 & w3266) | (w888 & w3266);
assign w2468 = ~w718 & w3267;
assign w2469 = w778 & w967;
assign w2470 = (~w2455 & w2742) | (~w2455 & w2743) | (w2742 & w2743);
assign w2471 = w761 & ~w787;
assign w2472 = (pi19 & w888) | (pi19 & w3268) | (w888 & w3268);
assign w2473 = (~w2455 & w2744) | (~w2455 & w2745) | (w2744 & w2745);
assign w2474 = (pi15 & w888) | (pi15 & w3269) | (w888 & w3269);
assign v574 = ~(w1002 | w889);
assign w2475 = v574;
assign w2476 = (~w2455 & w2896) | (~w2455 & w2897) | (w2896 & w2897);
assign w2477 = (~w2455 & w2746) | (~w2455 & w2747) | (w2746 & w2747);
assign w2478 = (~pi17 & w888) | (~pi17 & w3270) | (w888 & w3270);
assign w2479 = ~w888 & w3271;
assign w2480 = (~w2455 & w2748) | (~w2455 & w2749) | (w2748 & w2749);
assign w2481 = ~w888 & w3771;
assign w2482 = ~w888 & w3272;
assign w2483 = ~w888 & w3273;
assign w2484 = ~w1115 & w3957;
assign w2485 = w1042 & w1045;
assign w2486 = (~w4147 & w1064) | (~w4147 & w3274) | (w1064 & w3274);
assign w2487 = ~w1115 & w3958;
assign w2488 = ~w1275 & w2590;
assign w2489 = w1323 & pi23;
assign w2490 = (w2250 & w3275) | (w2250 & w3276) | (w3275 & w3276);
assign v575 = ~(w1355 | w1349);
assign w2491 = v575;
assign w2492 = ~w1274 & w1372;
assign w2493 = w1300 & w1415;
assign w2494 = ~w1300 & w1421;
assign v576 = ~(w1274 | w1460);
assign w2495 = v576;
assign v577 = ~(w1323 | pi23);
assign w2496 = v577;
assign w2497 = ~w1540 & w1592;
assign v578 = ~(w1378 | w1398);
assign w2498 = v578;
assign w2499 = ~w1468 & w1495;
assign w2500 = w1467 & w1648;
assign w2501 = w2293 & w3277;
assign w2502 = w1674 & ~w1620;
assign w2503 = (w1674 & ~w1426) | (w1674 & w3278) | (~w1426 & w3278);
assign w2504 = w1671 & w1681;
assign w2505 = w1684 & w4351;
assign w2506 = (w1489 & w4074) | (w1489 & w4075) | (w4074 & w4075);
assign w2507 = ~w1707 & w1686;
assign w2508 = w1698 & ~w1706;
assign w2509 = ~w1682 & w1732;
assign w2510 = w1743 & w1721;
assign w2511 = w1682 & w2592;
assign w2512 = w1749 & ~w1721;
assign w2513 = (w1749 & ~w1682) | (w1749 & w2593) | (~w1682 & w2593);
assign w2514 = w1764 & w1721;
assign w2515 = w1682 & w2594;
assign w2516 = ~w1564 & w1721;
assign w2517 = w1682 & w2595;
assign w2518 = w1778 & w1721;
assign w2519 = w1682 & w2596;
assign w2520 = w1640 & ~w1780;
assign w2521 = (w1669 & w3959) | (w1669 & w3960) | (w3959 & w3960);
assign w2522 = w1663 & w1721;
assign w2523 = w1682 & w2599;
assign v579 = ~(w1800 | w1721);
assign w2524 = v579;
assign w2525 = (~w1800 & ~w1682) | (~w1800 & w2600) | (~w1682 & w2600);
assign w2526 = w1757 & w1721;
assign w2527 = w1682 & w2601;
assign v580 = ~(w1556 | w1554);
assign w2528 = v580;
assign w2529 = w1601 & w1565;
assign w2530 = w1601 & ~w2306;
assign w2531 = ~w1816 & w1721;
assign w2532 = w1682 & w2602;
assign w2533 = w1817 & w1811;
assign v581 = ~(w1822 | w1826);
assign w2534 = v581;
assign w2535 = w1845 & w1721;
assign w2536 = w1682 & w3280;
assign w2537 = ~w1679 & w1721;
assign w2538 = w1682 & w2603;
assign w2539 = w1671 & ~w1630;
assign w2540 = w1850 & ~w1851;
assign w2541 = (w2605 & w2604) | (w2605 & ~w2301) | (w2604 & ~w2301);
assign w2542 = (w1669 & w3961) | (w1669 & w3962) | (w3961 & w3962);
assign w2543 = ~w1696 & w1721;
assign w2544 = w1682 & w2608;
assign w2545 = ~w1863 & w1867;
assign w2546 = (~w1717 & ~w1718) | (~w1717 & w3281) | (~w1718 & w3281);
assign w2547 = w1716 & w1721;
assign w2548 = w1682 & w2609;
assign w2549 = ~w1682 & w1878;
assign w2550 = (w1669 & w2750) | (w1669 & w2751) | (w2750 & w2751);
assign w2551 = w1616 & w1721;
assign w2552 = w1682 & w2610;
assign w2553 = (w1669 & w3963) | (w1669 & w3964) | (w3963 & w3964);
assign w2554 = ~w1646 & w1893;
assign w2555 = w1655 & w1721;
assign w2556 = w1682 & w2613;
assign w2557 = (w2615 & w2614) | (w2615 & ~w2301) | (w2614 & ~w2301);
assign w2558 = (w2617 & w2616) | (w2617 & ~w2301) | (w2616 & ~w2301);
assign w2559 = w1887 & pi21;
assign w2560 = ~w1898 & pi19;
assign w2561 = ~w1886 & w1924;
assign w2562 = ~w1937 & w1938;
assign w2563 = w1806 & ~w1736;
assign w2564 = w1553 & w1721;
assign w2565 = w1682 & w2618;
assign v582 = ~(w1937 | w1935);
assign w2566 = v582;
assign v583 = ~(w1886 | w1921);
assign w2567 = v583;
assign w2568 = (~w1857 & ~w1859) | (~w1857 & w2752) | (~w1859 & w2752);
assign w2569 = (w263 & w2753) | (w263 & w214) | (w2753 & w214);
assign w2570 = (w214 & w3701) | (w214 & w4170) | (w3701 & w4170);
assign w2571 = (pi16 & w3965) | (pi16 & w3764) | (w3965 & w3764);
assign w2572 = (w415 & w472) | (w415 & w2754) | (w472 & w2754);
assign v584 = ~(w759 | w733);
assign w2573 = v584;
assign v585 = ~(w778 | w787);
assign w2574 = v585;
assign w2575 = ~w778 & w971;
assign w2576 = (~pi15 & w1037) | (~pi15 & w3284) | (w1037 & w3284);
assign w2577 = (w1037 & w3966) | (w1037 & w3967) | (w3966 & w3967);
assign w2578 = ~w1154 & w3286;
assign w2579 = (~w1173 & ~w1298) | (~w1173 & w3968) | (~w1298 & w3968);
assign w2580 = (~pi17 & w1172) | (~pi17 & w3287) | (w1172 & w3287);
assign w2581 = w2579 & w3288;
assign w2582 = w2354 & w1721;
assign w2583 = w1682 & w3289;
assign w2584 = w528 & w530;
assign w2585 = w532 & w530;
assign w2586 = w2840 & w3290;
assign w2587 = ~w12 & pi11;
assign w2588 = pi11 & ~w680;
assign w2589 = pi11 & w677;
assign w2590 = w3062 & w1277;
assign w2591 = (w1331 & w3291) | (w1331 & w3292) | (w3291 & w3292);
assign w2592 = (w1743 & w1710) | (w1743 & w3969) | (w1710 & w3969);
assign w2593 = ~w1710 & w3293;
assign w2594 = ~w1711 & w1764;
assign w2595 = (~w1564 & w1710) | (~w1564 & w3294) | (w1710 & w3294);
assign w2596 = (w1778 & w1710) | (w1778 & w3295) | (w1710 & w3295);
assign w2597 = (pi15 & ~w1682) | (pi15 & w3296) | (~w1682 & w3296);
assign w2598 = (pi15 & ~w1721) | (pi15 & w3297) | (~w1721 & w3297);
assign w2599 = (w1663 & w1710) | (w1663 & w3298) | (w1710 & w3298);
assign w2600 = ~w1710 & w4340;
assign w2601 = (w1757 & w1710) | (w1757 & w3299) | (w1710 & w3299);
assign w2602 = (~w1816 & w1710) | (~w1816 & w3300) | (w1710 & w3300);
assign w2603 = (~w1679 & w1710) | (~w1679 & w3301) | (w1710 & w3301);
assign w2604 = w1682 & w3302;
assign w2605 = w1721 & w3303;
assign w2606 = (pi25 & ~w1682) | (pi25 & w3304) | (~w1682 & w3304);
assign w2607 = (pi25 & ~w1721) | (pi25 & w3305) | (~w1721 & w3305);
assign w2608 = (~w1696 & w1710) | (~w1696 & w3306) | (w1710 & w3306);
assign w2609 = (w1716 & w1710) | (w1716 & w3307) | (w1710 & w3307);
assign w2610 = (w1616 & w1710) | (w1616 & w3308) | (w1710 & w3308);
assign w2611 = (~pi21 & ~w1682) | (~pi21 & w3309) | (~w1682 & w3309);
assign w2612 = (~pi21 & ~w1721) | (~pi21 & w3310) | (~w1721 & w3310);
assign w2613 = (w1655 & w1710) | (w1655 & w3311) | (w1710 & w3311);
assign w2614 = w1682 & w3312;
assign w2615 = w1721 & w3313;
assign w2616 = w1682 & w3314;
assign w2617 = w1721 & w3315;
assign w2618 = (w1553 & w1710) | (w1553 & w3316) | (w1710 & w3316);
assign v586 = ~(w309 | w338);
assign w2619 = v586;
assign w2620 = w376 & ~w340;
assign w2621 = w376 & ~w2143;
assign w2622 = w389 & w386;
assign w2623 = w389 & w2147;
assign v587 = ~(w389 | w386);
assign w2624 = v587;
assign v588 = ~(w389 | w2147);
assign w2625 = v588;
assign w2626 = (w262 & w294) | (w262 & w2841) | (w294 & w2841);
assign w2627 = (w262 & ~w386) | (w262 & w2755) | (~w386 & w2755);
assign w2628 = ~w294 & w2842;
assign w2629 = w386 & w2756;
assign w2630 = ~w309 & w2148;
assign w2631 = w2149 | w416;
assign w2632 = (w416 & w2149) | (w416 & w309) | (w2149 & w309);
assign w2633 = w330 & w337;
assign w2634 = w354 & ~w360;
assign w2635 = ~w354 & w360;
assign w2636 = ~w371 & w382;
assign v589 = ~(w533 | w653);
assign w2637 = v589;
assign w2638 = (w672 & ~w510) | (w672 & w3970) | (~w510 & w3970);
assign w2639 = w581 & w692;
assign w2640 = (~w2639 & w2843) | (~w2639 & w2844) | (w2843 & w2844);
assign w2641 = (pi15 & w725) | (pi15 & w3971) | (w725 & w3971);
assign w2642 = ~w725 & w3972;
assign w2643 = (~w2639 & w2845) | (~w2639 & w2846) | (w2845 & w2846);
assign w2644 = (w3055 & w574) | (w3055 & w3973) | (w574 & w3973);
assign w2645 = (w2643 & w3317) | (w2643 & w3318) | (w3317 & w3318);
assign w2646 = (~w2639 & w2847) | (~w2639 & w2848) | (w2847 & w2848);
assign w2647 = ~w725 & w3974;
assign w2648 = (~pi09 & w725) | (~pi09 & w3975) | (w725 & w3975);
assign w2649 = w907 & w908;
assign w2650 = (~w717 & w3319) | (~w717 & w3320) | (w3319 & w3320);
assign w2651 = ~w1031 & w1212;
assign w2652 = w1209 & w2651;
assign v590 = ~(w1227 | w1235);
assign w2653 = v590;
assign w2654 = ~w1027 & w3321;
assign w2655 = (w1028 & ~w1034) | (w1028 & w3322) | (~w1034 & w3322);
assign w2656 = pi19 & ~w1252;
assign v591 = ~(w1251 | w1262);
assign w2657 = v591;
assign w2658 = ~w1234 & w1292;
assign w2659 = ~w1308 & w1311;
assign w2660 = (pi25 & w2244) | (pi25 & w1308) | (w2244 & w1308);
assign w2661 = ~w1220 & w1430;
assign v592 = ~(w1432 | w1434);
assign w2662 = v592;
assign v593 = ~(w1288 | w1300);
assign w2663 = v593;
assign w2664 = ~w1501 & w1450;
assign v594 = ~(w1423 | w1571);
assign w2665 = v594;
assign w2666 = (~w1423 & w1537) | (~w1423 & w3323) | (w1537 & w3323);
assign w2667 = (~pi13 & ~w1571) | (~pi13 & w3324) | (~w1571 & w3324);
assign w2668 = (~pi13 & w1537) | (~pi13 & w3325) | (w1537 & w3325);
assign w2669 = w1606 & ~w1466;
assign w2670 = w1468 & w1494;
assign w2671 = w1477 & ~w1500;
assign w2672 = w1571 & w3326;
assign w2673 = ~w1537 & w3327;
assign w2674 = w1642 & ~w1571;
assign w2675 = (w1642 & w1537) | (w1642 & w3328) | (w1537 & w3328);
assign w2676 = ~w1537 & w3329;
assign w2677 = w1541 & w3330;
assign v595 = ~(w1488 | w1503);
assign w2678 = v595;
assign w2679 = w1541 & w3331;
assign w2680 = ~w1683 & w1505;
assign w2681 = ~w1450 & w2680;
assign w2682 = ~w1687 & w1689;
assign w2683 = ~w1537 & w3332;
assign w2684 = (w1502 & w3333) | (w1502 & w3334) | (w3333 & w3334);
assign w2685 = (pi23 & ~w1541) | (pi23 & w3335) | (~w1541 & w3335);
assign w2686 = w2298 & w3336;
assign w2687 = pi25 & w1704;
assign v596 = ~(w1721 | w1736);
assign w2688 = v596;
assign w2689 = (pi05 & w1721) | (pi05 & w3337) | (w1721 & w3337);
assign w2690 = w1682 & w3338;
assign w2691 = w1721 & w3339;
assign w2692 = (~w1863 & w1672) | (~w1863 & w3340) | (w1672 & w3340);
assign w2693 = (w2546 & w1672) | (w2546 & w3341) | (w1672 & w3341);
assign w2694 = ~w1869 & w3342;
assign w2695 = w1682 & w3343;
assign w2696 = w1721 & w3344;
assign w2697 = w1795 & w1901;
assign w2698 = (pi29 & w1869) | (pi29 & w3345) | (w1869 & w3345);
assign w2699 = w2314 & pi31;
assign w2700 = (w1869 & w3346) | (w1869 & w3347) | (w3346 & w3347);
assign w2701 = pi31 & ~w1875;
assign w2702 = w1923 & w3348;
assign w2703 = w1972 & w1995;
assign v597 = ~(w2021 | w1788);
assign w2704 = v597;
assign w2705 = (~w2704 & w3976) | (~w2704 & w3977) | (w3976 & w3977);
assign w2706 = (w2704 & w3978) | (w2704 & w3979) | (w3978 & w3979);
assign w2707 = w2035 & ~w2022;
assign w2708 = w2037 & w2022;
assign w2709 = ~w48 & w2101;
assign v598 = ~(pi05 | w2112);
assign w2710 = v598;
assign w2711 = w72 & w175;
assign w2712 = w146 & w4352;
assign w2713 = ~w1257 & w3349;
assign w2714 = ~w1257 & w3350;
assign w2715 = ~w1257 & w3351;
assign w2716 = ~w1537 & w3352;
assign w2717 = (~pi17 & ~w1682) | (~pi17 & w3353) | (~w1682 & w3353);
assign w2718 = (~pi17 & ~w1721) | (~pi17 & w3354) | (~w1721 & w3354);
assign v599 = ~(w336 | w324);
assign w2719 = v599;
assign w2720 = w137 & w144;
assign w2721 = w3796 & w51;
assign v600 = ~(pi11 | w275);
assign w2722 = v600;
assign w2723 = ~pi11 & w282;
assign w2724 = w882 & ~w792;
assign w2725 = (w882 & ~w751) | (w882 & w3355) | (~w751 & w3355);
assign w2726 = w884 & w792;
assign w2727 = w751 & w3356;
assign w2728 = w893 & w787;
assign w2729 = (w893 & ~w751) | (w893 & w3357) | (~w751 & w3357);
assign w2730 = w917 & ~w792;
assign w2731 = (w917 & ~w751) | (w917 & w3358) | (~w751 & w3358);
assign w2732 = w919 & w792;
assign w2733 = w751 & w3359;
assign v601 = ~(w896 | w787);
assign w2734 = v601;
assign w2735 = w751 & w3980;
assign w2736 = ~w768 & w3360;
assign w2737 = (w801 & ~w751) | (w801 & w3361) | (~w751 & w3361);
assign w2738 = ~w768 & w3362;
assign w2739 = (~w931 & ~w751) | (~w931 & w2898) | (~w751 & w2898);
assign w2740 = ~w768 & w3363;
assign w2741 = (~w836 & ~w751) | (~w836 & w2899) | (~w751 & w2899);
assign w2742 = w730 & w787;
assign w2743 = (w730 & ~w751) | (w730 & w2900) | (~w751 & w2900);
assign w2744 = ~w768 & w3364;
assign w2745 = (w758 & ~w751) | (w758 & w2901) | (~w751 & w2901);
assign w2746 = w748 & w787;
assign w2747 = (w748 & ~w751) | (w748 & w2902) | (~w751 & w2902);
assign w2748 = ~w1001 & w787;
assign w2749 = (~w1001 & ~w751) | (~w1001 & w3365) | (~w751 & w3365);
assign w2750 = w1881 & w1878;
assign w2751 = ~w1682 & w2750;
assign w2752 = w1915 & ~w1857;
assign w2753 = ~pi11 & w263;
assign w2754 = (w146 & w3367) | (w146 & w3368) | (w3367 & w3368);
assign w2755 = w340 & w262;
assign v602 = ~(w340 | w262);
assign w2756 = v602;
assign w2757 = w19 & pi05;
assign w2758 = pi03 & pi30;
assign w2759 = ~w73 & w3369;
assign w2760 = (w138 & ~w98) | (w138 & w3370) | (~w98 & w3370);
assign w2761 = ~w137 & w148;
assign w2762 = ~w151 & w152;
assign v603 = ~(w137 | w154);
assign w2763 = v603;
assign w2764 = (w147 & ~w153) | (w147 & w2850) | (~w153 & w2850);
assign w2765 = (w147 & w2121) | (w147 & w137) | (w2121 & w137);
assign v604 = ~(w149 | w156);
assign w2766 = v604;
assign w2767 = ~w137 & w176;
assign v605 = ~(w199 | w194);
assign w2768 = v605;
assign w2769 = (~w199 & w153) | (~w199 & w3371) | (w153 & w3371);
assign w2770 = ~pi09 & w144;
assign w2771 = w144 & w4353;
assign w2772 = w155 & ~w2367;
assign w2773 = (~w324 & w2719) | (~w324 & w335) | (w2719 & w335);
assign v606 = ~(w337 | w318);
assign w2774 = v606;
assign v607 = ~(w475 | w473);
assign w2775 = v607;
assign w2776 = ~w475 & w2154;
assign w2777 = (~pi09 & w888) | (~pi09 & w3374) | (w888 & w3374);
assign w2778 = (~w1090 & ~w1093) | (~w1090 & w3981) | (~w1093 & w3981);
assign v608 = ~(w1106 | w1101);
assign w2779 = v608;
assign w2780 = ~w1165 & w1187;
assign v609 = ~(w1191 | w1194);
assign w2781 = v609;
assign w2782 = w1478 & w2903;
assign w2783 = (w1483 & ~w1478) | (w1483 & w2904) | (~w1478 & w2904);
assign w2784 = ~w1882 & w3982;
assign v610 = ~(w2096 | w2095);
assign w2785 = v610;
assign w2786 = (~w225 & w3983) | (~w225 & w3984) | (w3983 & w3984);
assign w2787 = ~w236 & w297;
assign w2788 = ~w237 & w269;
assign w2789 = (~w225 & w3985) | (~w225 & w3986) | (w3985 & w3986);
assign w2790 = (~w225 & w3987) | (~w225 & w3988) | (w3987 & w3988);
assign w2791 = (w225 & w3989) | (w225 & w3990) | (w3989 & w3990);
assign w2792 = w308 & ~w340;
assign w2793 = ~w554 & w547;
assign v611 = ~(w554 | w540);
assign w2794 = v611;
assign w2795 = ~w539 & w2851;
assign w2796 = w533 & ~w649;
assign v612 = ~(w540 | w649);
assign w2797 = v612;
assign w2798 = w367 & w396;
assign w2799 = w516 & ~w518;
assign v613 = ~(w516 | w520);
assign w2800 = v613;
assign w2801 = ~w516 & w528;
assign w2802 = (~w434 & ~w576) | (~w434 & w3991) | (~w576 & w3991);
assign w2803 = ~w560 & w3375;
assign w2804 = w778 & w3376;
assign v614 = ~(w889 | w934);
assign w2805 = v614;
assign w2806 = w889 & pi01;
assign w2807 = (w2455 & w2905) | (w2455 & w2906) | (w2905 & w2906);
assign w2808 = w1059 & w1043;
assign w2809 = ~w979 & w3377;
assign w2810 = ~w1090 & w1043;
assign w2811 = ~w979 & w3378;
assign w2812 = ~w1101 & w1043;
assign w2813 = ~w1115 & w3992;
assign w2814 = w1049 & w3199;
assign w2815 = (w4038 & w4076) | (w4038 & w4077) | (w4076 & w4077);
assign w2816 = ~w1115 & w3994;
assign w2817 = (~w1142 & w1046) | (~w1142 & w3995) | (w1046 & w3995);
assign w2818 = ~w1131 & w1126;
assign w2819 = (w1115 & w3996) | (w1115 & w3997) | (w3996 & w3997);
assign w2820 = w1116 & w2211;
assign w2821 = (~w1155 & w1046) | (~w1155 & w3998) | (w1046 & w3998);
assign w2822 = (~w1182 & w1046) | (~w1182 & w3999) | (w1046 & w3999);
assign w2823 = w1258 & w1244;
assign w2824 = ~w1061 & w4000;
assign w2825 = ~w1046 & w1282;
assign w2826 = w1249 & ~w1294;
assign w2827 = (~w1258 & w1257) | (~w1258 & w4171) | (w1257 & w4171);
assign w2828 = ~w1296 & w2263;
assign v615 = ~(w244 | w237);
assign w2829 = v615;
assign w2830 = w319 & ~w237;
assign w2831 = (~w225 & w4001) | (~w225 & w4002) | (w4001 & w4002);
assign w2832 = ~w1352 & w3380;
assign w2833 = w1353 & ~w1295;
assign w2834 = w1352 & w3381;
assign w2835 = w28 & w2721;
assign w2836 = w127 & ~w76;
assign w2837 = pi05 & ~w123;
assign w2838 = (~w42 & w3382) | (~w42 & w3383) | (w3382 & w3383);
assign v616 = ~(pi07 | w340);
assign w2839 = v616;
assign w2840 = ~w516 & w2584;
assign w2841 = ~w308 & w262;
assign w2842 = w308 & ~w262;
assign w2843 = w745 & ~w692;
assign w2844 = (w745 & ~w589) | (w745 & w2907) | (~w589 & w2907);
assign w2845 = (w770 & ~w683) | (w770 & w3384) | (~w683 & w3384);
assign w2846 = (w770 & ~w589) | (w770 & w3385) | (~w589 & w3385);
assign w2847 = (w656 & ~w683) | (w656 & w3386) | (~w683 & w3386);
assign w2848 = (w656 & ~w589) | (w656 & w2908) | (~w589 & w2908);
assign w2849 = (~w98 & ~w2721) | (~w98 & w3387) | (~w2721 & w3387);
assign w2850 = w2332 | w147;
assign w2851 = ~w491 & w3388;
assign v617 = ~(w59 | w54);
assign w2852 = v617;
assign w2853 = w95 & w65;
assign v618 = ~(w96 | w101);
assign w2854 = v618;
assign w2855 = w95 & w106;
assign w2856 = (w146 & w3389) | (w146 & w3390) | (w3389 & w3390);
assign w2857 = w147 & w2760;
assign w2858 = w64 & ~pi07;
assign w2859 = (~w2765 & w3391) | (~w2765 & w3392) | (w3391 & w3392);
assign w2860 = ~w117 & w182;
assign w2861 = w117 & ~w182;
assign w2862 = (w194 & w102) | (w194 & w3393) | (w102 & w3393);
assign w2863 = (w202 & w102) | (w202 & w3394) | (w102 & w3394);
assign v619 = ~(w177 | w179);
assign w2864 = v619;
assign w2865 = (w146 & ~w153) | (w146 & w3395) | (~w153 & w3395);
assign w2866 = (w28 & w173) | (w28 & w4004) | (w173 & w4004);
assign w2867 = (pi22 & ~w2721) | (pi22 & w4354) | (~w2721 & w4354);
assign w2868 = (w225 & w4005) | (w225 & w4006) | (w4005 & w4006);
assign w2869 = (w347 & w3396) | (w347 & ~w320) | (w3396 & ~w320);
assign w2870 = (w3396 & w3397) | (w3396 & w335) | (w3397 & w335);
assign w2871 = (w233 & w4007) | (w233 & w4008) | (w4007 & w4008);
assign w2872 = (w227 & w4009) | (w227 & w4010) | (w4009 & w4010);
assign w2873 = (w3400 & w227) | (w3400 & w4011) | (w227 & w4011);
assign w2874 = w353 & ~w2142;
assign w2875 = ~w293 & w262;
assign w2876 = (w233 & w4012) | (w233 & w4013) | (w4012 & w4013);
assign w2877 = pi13 & ~w2393;
assign w2878 = pi13 & ~w2394;
assign v620 = ~(pi13 | w2395);
assign w2879 = v620;
assign v621 = ~(pi13 | w2396);
assign w2880 = v621;
assign w2881 = ~w1110 & w1120;
assign w2882 = ~w921 & w886;
assign w2883 = w928 & ~w943;
assign w2884 = w1168 & ~w1017;
assign w2885 = w1168 & w2214;
assign v622 = ~(w944 | w949);
assign w2886 = v622;
assign v623 = ~(w1222 | w1225);
assign w2887 = v623;
assign w2888 = ~w1033 & w1228;
assign w2889 = ~w237 & w270;
assign w2890 = w237 & ~w270;
assign w2891 = (~w742 & w3402) | (~w742 & w3403) | (w3402 & w3403);
assign w2892 = ~w851 & w864;
assign w2893 = w851 & w855;
assign w2894 = w951 & w3404;
assign w2895 = (pi11 & ~w951) | (pi11 & w3405) | (~w951 & w3405);
assign w2896 = ~w1013 & w787;
assign w2897 = (~w1013 & ~w751) | (~w1013 & w3406) | (~w751 & w3406);
assign w2898 = ~w760 & w3407;
assign w2899 = ~w760 & w3408;
assign w2900 = w761 & w730;
assign w2901 = ~w760 & w3409;
assign w2902 = w761 & w748;
assign w2903 = ~w1300 & w1481;
assign w2904 = w1300 & w1483;
assign w2905 = (~pi21 & w3410) | (~pi21 & ~w787) | (w3410 & ~w787);
assign w2906 = (w751 & w3410) | (w751 & w3411) | (w3410 & w3411);
assign w2907 = ~w601 & w745;
assign w2908 = ~w601 & w656;
assign w2909 = (~pi09 & ~w656) | (~pi09 & w12) | (~w656 & w12);
assign w2910 = w657 & w666;
assign w2911 = w581 & ~w660;
assign w2912 = ~w603 & w3412;
assign w2913 = (~w857 & w603) | (~w857 & w3413) | (w603 & w3413);
assign w2914 = ~w944 & w962;
assign w2915 = (w783 & w772) | (w783 & w4172) | (w772 & w4172);
assign w2916 = (w772 & w783) | (w772 & w3055) | (w783 & w3055);
assign w2917 = (pi19 & w562) | (pi19 & w4014) | (w562 & w4014);
assign w2918 = pi19 & w2181;
assign w2919 = (~w717 & w3414) | (~w717 & w3415) | (w3414 & w3415);
assign w2920 = pi24 & pi28;
assign w2921 = w5 & w66;
assign w2922 = w64 & w3416;
assign w2923 = pi24 & ~pi26;
assign v624 = ~(w59 | w94);
assign w2924 = v624;
assign w2925 = w16 & ~pi19;
assign v625 = ~(pi17 | pi15);
assign w2926 = v625;
assign w2927 = w27 & w112;
assign w2928 = w67 & w113;
assign w2929 = w115 & ~w76;
assign v626 = ~(w107 | w117);
assign w2930 = v626;
assign w2931 = pi03 & ~pi24;
assign w2932 = pi03 & pi24;
assign v627 = ~(w64 | pi07);
assign w2933 = v627;
assign w2934 = w89 & w139;
assign w2935 = ~pi09 & w143;
assign v628 = ~(w159 | pi07);
assign w2936 = v628;
assign w2937 = w174 & w2721;
assign w2938 = w2721 & w3417;
assign w2939 = (w146 & w3418) | (w146 & w3419) | (w3418 & w3419);
assign w2940 = w175 & w2760;
assign w2941 = w2721 & w3421;
assign w2942 = w2721 & w3422;
assign w2943 = pi03 & ~pi22;
assign w2944 = ~w195 & w200;
assign w2945 = w2721 & w3423;
assign w2946 = w2721 & w3424;
assign w2947 = ~w102 & w3425;
assign v629 = ~(w204 | w203);
assign w2948 = v629;
assign w2949 = ~w2364 & pi11;
assign w2950 = (pi09 & ~w163) | (pi09 & w3426) | (~w163 & w3426);
assign w2951 = w163 & w3427;
assign w2952 = pi18 & ~pi20;
assign w2953 = w3752 & w281;
assign w2954 = (~pi11 & w173) | (~pi11 & w4015) | (w173 & w4015);
assign w2955 = (~w153 & w3429) | (~w153 & w3430) | (w3429 & w3430);
assign w2956 = pi11 & w2865;
assign w2957 = ~w69 & w4355;
assign w2958 = pi03 & ~pi18;
assign w2959 = ~w309 & w355;
assign w2960 = w109 & w2926;
assign w2961 = ~w424 & w415;
assign w2962 = ~w401 & w426;
assign w2963 = w109 & w3432;
assign w2964 = w109 & w3433;
assign w2965 = (pi01 & ~w338) | (pi01 & w3436) | (~w338 & w3436);
assign v630 = ~(w373 | w340);
assign w2966 = v630;
assign w2967 = (~w373 & ~w338) | (~w373 & w2966) | (~w338 & w2966);
assign w2968 = w338 & w3439;
assign w2969 = ~w524 & pi15;
assign w2970 = w430 & ~pi15;
assign v631 = ~(w424 | pi15);
assign w2971 = v631;
assign w2972 = w541 & ~pi13;
assign w2973 = ~w541 & pi13;
assign w2974 = w524 & ~pi15;
assign w2975 = (~pi17 & w522) | (~pi17 & w3440) | (w522 & w3440);
assign w2976 = (w3796 & w432) | (w3796 & w4173) | (w432 & w4173);
assign w2977 = w3796 & ~w529;
assign w2978 = ~w522 & w3441;
assign v632 = ~(w533 | w546);
assign w2979 = v632;
assign w2980 = (~w444 & w4016) | (~w444 & w4356) | (w4016 & w4356);
assign w2981 = (~pi09 & ~w606) | (~pi09 & w3442) | (~w606 & w3442);
assign w2982 = ~w481 & w477;
assign v633 = ~(w631 | w630);
assign w2983 = v633;
assign w2984 = pi12 & pi14;
assign w2985 = pi05 & ~w634;
assign w2986 = ~pi01 & w634;
assign w2987 = (~w640 & w606) | (~w640 & w3015) | (w606 & w3015);
assign w2988 = ~w636 & w642;
assign w2989 = (w686 & w566) | (w686 & w3443) | (w566 & w3443);
assign w2990 = w686 & ~w551;
assign w2991 = w484 & ~w510;
assign w2992 = ~pi15 & w109;
assign w2993 = ~w659 & w4174;
assign w2994 = (w589 & w602) | (w589 & w3444) | (w602 & w3444);
assign w2995 = w589 & ~w702;
assign w2996 = (w779 & w562) | (w779 & w3445) | (w562 & w3445);
assign v634 = ~(w434 | w2996);
assign w2997 = v634;
assign w2998 = (~w434 & ~w2181) | (~w434 & w3446) | (~w2181 & w3446);
assign w2999 = pi21 & w529;
assign w3000 = ~w786 & w780;
assign w3001 = (w716 & w4175) | (w716 & w4176) | (w4175 & w4176);
assign w3002 = (w791 & w2182) | (w791 & w786) | (w2182 & w786);
assign w3003 = (w526 & w4017) | (w526 & w4018) | (w4017 & w4018);
assign w3004 = (pi14 & w566) | (pi14 & w4019) | (w566 & w4019);
assign w3005 = (w572 & w4177) | (w572 & w4178) | (w4177 & w4178);
assign w3006 = w109 & w639;
assign w3007 = (w805 & w3450) | (w805 & w572) | (w3450 & w572);
assign w3008 = w109 & ~w808;
assign w3009 = pi03 & ~pi12;
assign w3010 = ~w687 & w805;
assign w3011 = pi05 & w794;
assign w3012 = (w590 & w4020) | (w590 & w4021) | (w4020 & w4021);
assign v635 = ~(w832 | w833);
assign w3013 = v635;
assign w3014 = ~w629 & w794;
assign w3015 = (pi05 & w639) | (pi05 & w2108) | (w639 & w2108);
assign w3016 = ~w639 & w2101;
assign v636 = ~(w850 | w851);
assign w3017 = v636;
assign w3018 = w606 & ~w611;
assign w3019 = (w606 & w566) | (w606 & w3018) | (w566 & w3018);
assign w3020 = (w590 & w3451) | (w590 & w3452) | (w3451 & w3452);
assign w3021 = (~w590 & w3453) | (~w590 & w3454) | (w3453 & w3454);
assign w3022 = ~w848 & w860;
assign w3023 = (~w590 & w3455) | (~w590 & w3456) | (w3455 & w3456);
assign w3024 = w750 & w792;
assign w3025 = w724 & w4179;
assign w3026 = (~pi05 & ~w724) | (~pi05 & w4180) | (~w724 & w4180);
assign w3027 = w750 & ~w787;
assign w3028 = pi03 & ~pi10;
assign w3029 = (pi05 & ~w724) | (pi05 & w4181) | (~w724 & w4181);
assign w3030 = w724 & w4182;
assign w3031 = ~w603 & w3457;
assign w3032 = (~w854 & w603) | (~w854 & w3458) | (w603 & w3458);
assign v637 = ~(w802 | w860);
assign w3033 = v637;
assign w3034 = (w3459 & w3460) | (w3459 & ~w717) | (w3460 & ~w717);
assign w3035 = pi21 & w574;
assign w3036 = pi10 & ~pi01;
assign w3037 = (pi10 & w872) | (pi10 & w3461) | (w872 & w3461);
assign w3038 = (w1050 & w432) | (w1050 & w4183) | (w432 & w4183);
assign w3039 = w1050 & ~w529;
assign w3040 = w783 & w1052;
assign w3041 = w553 & pi17;
assign w3042 = (w3796 & ~w1070) | (w3796 & w3462) | (~w1070 & w3462);
assign w3043 = ~w1082 & w1059;
assign w3044 = pi06 & pi08;
assign w3045 = w3062 & w3463;
assign w3046 = w783 & w1100;
assign w3047 = ~w1115 & w4024;
assign w3048 = (pi05 & w902) | (pi05 & w3464) | (w902 & w3464);
assign w3049 = ~w902 & w3465;
assign w3050 = (~pi11 & w888) | (~pi11 & w3467) | (w888 & w3467);
assign w3051 = ~w888 & w3468;
assign w3052 = (pi15 & w888) | (pi15 & w3469) | (w888 & w3469);
assign w3053 = w3062 & w3470;
assign w3054 = w3471 & ~w1051;
assign w3055 = w3062 & w3472;
assign w3056 = (~pi19 & w888) | (~pi19 & w3473) | (w888 & w3473);
assign w3057 = ~w888 & w3474;
assign w3058 = ~w1067 & w1072;
assign w3059 = (w3475 & ~w784) | (w3475 & w4033) | (~w784 & w4033);
assign v638 = ~(w784 | w2203);
assign w3060 = v638;
assign w3061 = (w783 & w1064) | (w783 & w3476) | (w1064 & w3476);
assign w3062 = w14 & w15;
assign w3063 = (pi27 & ~w1300) | (pi27 & w3478) | (~w1300 & w3478);
assign w3064 = ~w1295 & w3479;
assign w3065 = w1322 & ~w2243;
assign v639 = ~(w1308 | w1310);
assign w3066 = v639;
assign w3067 = (~w434 & ~w1300) | (~w434 & w3481) | (~w1300 & w3481);
assign w3068 = ~w1115 & w4025;
assign w3069 = w1134 & w1148;
assign w3070 = ~w1295 & w3482;
assign w3071 = w1427 & ~w2243;
assign w3072 = ~w1218 & w1258;
assign w3073 = (~w1218 & ~w1294) | (~w1218 & w3072) | (~w1294 & w3072);
assign w3074 = (w1441 & ~w1300) | (w1441 & w4026) | (~w1300 & w4026);
assign w3075 = pi17 & ~w1167;
assign w3076 = (w1203 & w1193) | (w1203 & w3483) | (w1193 & w3483);
assign w3077 = w1121 & w3484;
assign w3078 = pi15 & ~w1197;
assign w3079 = (w3772 & w4027) | (w3772 & w4028) | (w4027 & w4028);
assign v640 = ~(pi15 | w1197);
assign w3080 = v640;
assign v641 = ~(w1338 | w1);
assign w3081 = v641;
assign w3082 = w1507 & w1505;
assign w3083 = w1507 & w2273;
assign v642 = ~(w1508 | w1339);
assign w3084 = v642;
assign w3085 = w1334 & pi01;
assign w3086 = (~w1513 & w1337) | (~w1513 & w3485) | (w1337 & w3485);
assign w3087 = w14 & w1518;
assign w3088 = ~w1332 & w1519;
assign w3089 = w2277 & w4029;
assign v643 = ~(w1349 | w1352);
assign w3090 = v643;
assign w3091 = w1349 & w1352;
assign w3092 = w1358 & w1363;
assign w3093 = w1485 & ~w1606;
assign w3094 = ~w1485 & w1606;
assign w3095 = ~w2670 & w1613;
assign w3096 = ~w1614 & w1538;
assign w3097 = w1608 & w1622;
assign w3098 = ~w1537 & w3486;
assign w3099 = ~w1537 & w3487;
assign w3100 = ~w1313 & w3488;
assign w3101 = (~w434 & w1312) | (~w434 & w3489) | (w1312 & w3489);
assign w3102 = w1450 & ~w1699;
assign w3103 = ~w1537 & w3490;
assign w3104 = ~w1714 & w1727;
assign w3105 = ~w1714 & w2300;
assign v644 = ~(pi05 | w1712);
assign w3106 = v644;
assign w3107 = pi03 & ~pi02;
assign v645 = ~(pi03 | pi02);
assign w3108 = v645;
assign w3109 = w2512 & w2513;
assign w3110 = (w2513 & w2512) | (w2513 & ~w1721) | (w2512 & ~w1721);
assign w3111 = (w1725 & w1721) | (w1725 & w3491) | (w1721 & w3491);
assign w3112 = (w1725 & w2302) | (w1725 & w1736) | (w2302 & w1736);
assign v646 = ~(w1518 | w1525);
assign w3113 = v646;
assign v647 = ~(w1761 | w1758);
assign w3114 = v647;
assign v648 = ~(pi13 | pi11);
assign w3115 = v648;
assign w3116 = (~w1780 & w2520) | (~w1780 & w1602) | (w2520 & w1602);
assign w3117 = (~w1780 & w2520) | (~w1780 & w1557) | (w2520 & w1557);
assign w3118 = w1576 & ~w1585;
assign w3119 = w1791 & ~w1789;
assign w3120 = w2524 & w2525;
assign w3121 = (w2525 & w2524) | (w2525 & ~w1721) | (w2524 & ~w1721);
assign w3122 = (~pi09 & w1800) | (~pi09 & w12) | (w1800 & w12);
assign w3123 = w1838 & pi21;
assign w3124 = (~pi23 & ~w1721) | (~pi23 & w3492) | (~w1721 & w3492);
assign v649 = ~(pi23 | w2536);
assign w3125 = v649;
assign v650 = ~(w1850 | w1853);
assign w3126 = v650;
assign w3127 = ~w1862 & w2545;
assign w3128 = ~w1838 & w1865;
assign w3129 = (~w1694 & w3493) | (~w1694 & w3494) | (w3493 & w3494);
assign v651 = ~(w1711 | w1876);
assign w3130 = v651;
assign v652 = ~(w1873 | pi31);
assign w3131 = v652;
assign w3132 = (~w310 & w3495) | (~w310 & w3496) | (w3495 & w3496);
assign w3133 = (w1289 & w3497) | (w1289 & w3498) | (w3497 & w3498);
assign w3134 = (w3499 & ~w1331) | (w3499 & ~w3101) | (~w1331 & ~w3101);
assign w3135 = (w1685 & w4030) | (w1685 & w4031) | (w4030 & w4031);
assign w3136 = ~pi01 & pi02;
assign v653 = ~(w1735 | w1751);
assign w3137 = v653;
assign w3138 = w1968 & pi09;
assign v654 = ~(w1968 | pi09);
assign w3139 = v654;
assign w3140 = w1959 & ~w1804;
assign w3141 = (w310 & w3640) | (w310 & w3500) | (w3640 & w3500);
assign w3142 = (pi11 & w3501) | (pi11 & w4357) | (w3501 & w4357);
assign w3143 = (w310 & w3643) | (w310 & w3502) | (w3643 & w3502);
assign w3144 = (~pi11 & w3503) | (~pi11 & w4357) | (w3503 & w4357);
assign w3145 = w1984 & ~w1990;
assign w3146 = w1992 & ~w1997;
assign w3147 = w1768 & ~pi11;
assign w3148 = ~w1768 & pi11;
assign v655 = ~(w2321 | w2010);
assign w3149 = v655;
assign w3150 = (~w2010 & w2008) | (~w2010 & w3504) | (w2008 & w3504);
assign w3151 = ~w2009 & w3149;
assign w3152 = w2009 & ~w2018;
assign w3153 = w1818 & ~w1788;
assign w3154 = (w1788 & w2018) | (w1788 & w3505) | (w2018 & w3505);
assign w3155 = w2026 & ~w2019;
assign w3156 = (w310 & w3646) | (w310 & w3506) | (w3646 & w3506);
assign w3157 = (~pi17 & w3507) | (~pi17 & w4357) | (w3507 & w4357);
assign w3158 = (w310 & w3649) | (w310 & w3508) | (w3649 & w3508);
assign w3159 = (pi17 & w3509) | (pi17 & w4357) | (w3509 & w4357);
assign v656 = ~(w1797 | w1905);
assign w3160 = v656;
assign w3161 = ~w1797 & w2323;
assign w3162 = (~w1909 & w1906) | (~w1909 & w3510) | (w1906 & w3510);
assign w3163 = ~w2062 & w2052;
assign w3164 = (~w2062 & w1906) | (~w2062 & w3163) | (w1906 & w3163);
assign w3165 = w2062 & ~w2052;
assign w3166 = ~w1906 & w3165;
assign w3167 = ~w2325 & w1917;
assign v657 = ~(w2070 | w2069);
assign w3168 = v657;
assign v658 = ~(pi30 | w67);
assign w3169 = v658;
assign v659 = ~(w2081 | w2082);
assign w3170 = v659;
assign w3171 = w2090 & w2080;
assign w3172 = w2079 & w3171;
assign w3173 = w2097 & ~w2091;
assign w3174 = (w1917 & w4184) | (w1917 & w4185) | (w4184 & w4185);
assign w3175 = w114 & w3511;
assign w3176 = ~w237 & w268;
assign w3177 = w400 & w3512;
assign w3178 = w501 & w3513;
assign w3179 = ~w501 & w3514;
assign w3180 = ~w400 & w3515;
assign w3181 = ~w533 & w2341;
assign w3182 = ~w533 & w2342;
assign w3183 = (~pi17 & w602) | (~pi17 & w3516) | (w602 & w3516);
assign v660 = ~(pi17 | w702);
assign w3184 = v660;
assign w3185 = ~w687 & pi11;
assign w3186 = ~w690 & w3517;
assign w3187 = ~pi13 & w756;
assign w3188 = (pi19 & w602) | (pi19 & w3518) | (w602 & w3518);
assign w3189 = pi19 & ~w702;
assign w3190 = ~w602 & w3519;
assign w3191 = ~pi19 & w702;
assign w3192 = w600 & ~w572;
assign w3193 = (w791 & w2996) | (w791 & w3520) | (w2996 & w3520);
assign w3194 = (w2181 & w3520) | (w2181 & w3521) | (w3520 & w3521);
assign w3195 = (w2421 & w3522) | (w2421 & w3523) | (w3522 & w3523);
assign w3196 = ~w850 & w2892;
assign w3197 = (w855 & w2893) | (w855 & w850) | (w2893 & w850);
assign w3198 = ~w1056 & w1053;
assign w3199 = pi05 & ~w1053;
assign w3200 = (w3039 & w4186) | (w3039 & w4187) | (w4186 & w4187);
assign w3201 = ~w888 & w3527;
assign w3202 = (w3039 & w4188) | (w3039 & w4189) | (w4188 & w4189);
assign w3203 = ~w1154 & w3529;
assign w3204 = (pi13 & w2578) | (pi13 & w4358) | (w2578 & w4358);
assign w3205 = (w4147 & w888) | (w4147 & w3530) | (w888 & w3530);
assign w3206 = (w4147 & w888) | (w4147 & w3531) | (w888 & w3531);
assign w3207 = (~w3039 & ~pi23) | (~w3039 & w3532) | (~pi23 & w3532);
assign w3208 = (~w310 & w3533) | (~w310 & w3534) | (w3533 & w3534);
assign w3209 = (~w1278 & w979) | (~w1278 & w3535) | (w979 & w3535);
assign v661 = ~(w1278 | w1043);
assign w3210 = v661;
assign w3211 = w1301 & ~pi25;
assign w3212 = (pi19 & w1300) | (pi19 & w3536) | (w1300 & w3536);
assign w3213 = w1518 & w3537;
assign w3214 = (pi05 & ~w1518) | (pi05 & w3538) | (~w1518 & w3538);
assign w3215 = w1449 & ~w1439;
assign w3216 = ~w1666 & w2358;
assign w3217 = w1721 & w3539;
assign w3218 = pi23 & w2536;
assign w3219 = (~w1738 & w3540) | (~w1738 & w3541) | (w3540 & w3541);
assign v662 = ~(w1936 | w1873);
assign w3220 = v662;
assign w3221 = w124 & w75;
assign w3222 = w124 & w2360;
assign w3223 = w123 & w75;
assign w3224 = ~w220 & w2835;
assign v663 = ~(w32 | w2960);
assign w3225 = v663;
assign w3226 = w452 & w110;
assign w3227 = w452 & w2960;
assign w3228 = (pi07 & w3764) | (pi07 & w4190) | (w3764 & w4190);
assign w3229 = ~w415 & w423;
assign w3230 = ~w541 & pi15;
assign w3231 = w541 & ~pi15;
assign w3232 = (pi21 & w888) | (pi21 & w3542) | (w888 & w3542);
assign w3233 = (pi17 & w888) | (pi17 & w3543) | (w888 & w3543);
assign w3234 = ~w1301 & pi25;
assign w3235 = (pi21 & w1257) | (pi21 & w3544) | (w1257 & w3544);
assign w3236 = ~w1257 & w3545;
assign w3237 = w1712 & ~pi05;
assign w3238 = ~w10 & w50;
assign w3239 = w320 & w3546;
assign w3240 = w344 & ~w2773;
assign w3241 = w146 & ~w32;
assign w3242 = w146 & w4372;
assign w3243 = (w321 & w3241) | (w321 & w4191) | (w3241 & w4191);
assign w3244 = (w3241 & w321) | (w3241 & w2712) | (w321 & w2712);
assign w3245 = ~w469 & w2336;
assign v664 = ~(w469 | w467);
assign w3246 = v664;
assign w3247 = pi05 & w452;
assign w3248 = ~w456 & w3547;
assign w3249 = pi05 & ~w452;
assign w3250 = w456 & w3548;
assign w3251 = ~w515 & w563;
assign w3252 = w483 & w570;
assign v665 = ~(w515 | w435);
assign w3253 = v665;
assign w3254 = (w2977 & w4192) | (w2977 & w4193) | (w4192 & w4193);
assign v666 = ~(w580 | w2170);
assign w3255 = v666;
assign w3256 = w533 & w615;
assign w3257 = ~w533 & w625;
assign w3258 = w533 & ~w632;
assign w3259 = ~w504 & w2589;
assign w3260 = w12 & ~pi11;
assign w3261 = ~w781 & w792;
assign w3262 = (pi12 & ~w683) | (pi12 & w3549) | (~w683 & w3549);
assign w3263 = (pi12 & ~w658) | (pi12 & w3550) | (~w658 & w3550);
assign v667 = ~(w781 | w787);
assign w3264 = v667;
assign w3265 = w762 & ~w912;
assign v668 = ~(w2466 | pi11);
assign w3266 = v668;
assign w3267 = ~w763 & pi19;
assign w3268 = ~w2470 & pi19;
assign w3269 = ~w2473 & pi15;
assign v669 = ~(w2477 | pi17);
assign w3270 = v669;
assign w3271 = w2477 & pi17;
assign w3272 = w2473 & ~pi15;
assign w3273 = w2470 & ~pi19;
assign w3274 = w1075 & ~w4147;
assign w3275 = w1355 & w1348;
assign w3276 = w1355 & ~w1295;
assign w3277 = (pi17 & w1537) | (pi17 & w3551) | (w1537 & w3551);
assign w3278 = ~w2351 & w1674;
assign w3279 = (w2591 & w1312) | (w2591 & w3552) | (w1312 & w3552);
assign w3280 = (w1845 & w1710) | (w1845 & w4194) | (w1710 & w4194);
assign v670 = ~(w1715 | w1717);
assign w3281 = v670;
assign w3282 = ~w323 & w3553;
assign w3283 = ~w323 & w4195;
assign w3284 = ~w888 & w3555;
assign w3285 = w3556 & ~w1051;
assign w3286 = w3557 & ~w1051;
assign w3287 = (w1117 & w4196) | (w1117 & w4197) | (w4196 & w4197);
assign w3288 = ~w1294 & w4359;
assign w3289 = (w2354 & w1710) | (w2354 & w3558) | (w1710 & w3558);
assign w3290 = ~w515 & w532;
assign w3291 = (~w310 & w3559) | (~w310 & w3560) | (w3559 & w3560);
assign w3292 = (~w310 & w3561) | (~w310 & w3562) | (w3561 & w3562);
assign w3293 = (~w1694 & w3563) | (~w1694 & w3564) | (w3563 & w3564);
assign w3294 = w1695 & ~w1564;
assign w3295 = w1695 & w1778;
assign w3296 = ~w2596 & pi15;
assign w3297 = ~w1778 & pi15;
assign w3298 = w1695 & w1663;
assign w3299 = w1695 & w1757;
assign w3300 = w1695 & ~w1816;
assign w3301 = w1695 & ~w1679;
assign w3302 = w2603 & ~pi25;
assign w3303 = (~pi25 & w1678) | (~pi25 & w4199) | (w1678 & w4199);
assign w3304 = ~w2603 & pi25;
assign w3305 = ~w1678 & w4200;
assign w3306 = w1695 & ~w1696;
assign w3307 = w1695 & w1716;
assign w3308 = w1695 & w1616;
assign v671 = ~(w2610 | pi21);
assign w3309 = v671;
assign v672 = ~(w1616 | pi21);
assign w3310 = v672;
assign w3311 = w1695 & w1655;
assign w3312 = w2613 & ~pi19;
assign w3313 = w1655 & ~pi19;
assign w3314 = w2596 & ~pi15;
assign w3315 = w1778 & ~pi15;
assign w3316 = w1695 & w1553;
assign w3317 = w785 & w770;
assign w3318 = ~w659 & w4201;
assign w3319 = (~w2996 & w2649) | (~w2996 & w3565) | (w2649 & w3565);
assign w3320 = w907 & w4360;
assign w3321 = (w4147 & w888) | (w4147 & w3566) | (w888 & w3566);
assign w3322 = w1028 & w963;
assign w3323 = ~w1330 & w3567;
assign v673 = ~(w1423 | pi13);
assign w3324 = v673;
assign w3325 = ~w1330 & w3568;
assign w3326 = w1423 & pi13;
assign w3327 = (pi13 & w1330) | (pi13 & w3569) | (w1330 & w3569);
assign w3328 = ~w1330 & w3570;
assign w3329 = (~pi17 & w1330) | (~pi17 & w3571) | (w1330 & w3571);
assign v674 = ~(w1499 | pi19);
assign w3330 = v674;
assign w3331 = (~pi23 & ~w1436) | (~pi23 & w3572) | (~w1436 & w3572);
assign w3332 = (pi27 & w1330) | (pi27 & w3573) | (w1330 & w3573);
assign w3333 = ~w1326 & w1505;
assign w3334 = ~w1450 & w3333;
assign w3335 = w1436 & w3574;
assign w3336 = (pi25 & w1537) | (pi25 & w3575) | (w1537 & w3575);
assign w3337 = (pi05 & w1725) | (pi05 & w3576) | (w1725 & w3576);
assign w3338 = w2595 & w1769;
assign w3339 = ~w1564 & w1769;
assign v675 = ~(w2308 | w1863);
assign w3340 = v675;
assign w3341 = ~w2308 & w2546;
assign w3342 = w1871 & ~pi29;
assign w3343 = w2609 & ~pi27;
assign w3344 = (w2508 & w3577) | (w2508 & w3578) | (w3577 & w3578);
assign w3345 = ~w1871 & pi29;
assign w3346 = w2314 | pi31;
assign w3347 = (pi31 & w2314) | (pi31 & ~w1871) | (w2314 & ~w1871);
assign w3348 = pi11 & ~w1972;
assign w3349 = w1244 & pi01;
assign w3350 = w1244 & w1098;
assign w3351 = w1244 & w1348;
assign w3352 = (pi15 & w1330) | (pi15 & w3579) | (w1330 & w3579);
assign v676 = ~(w2599 | pi17);
assign w3353 = v676;
assign v677 = ~(w1663 | pi17);
assign w3354 = v677;
assign w3355 = w761 & w882;
assign w3356 = ~w761 & w884;
assign w3357 = w761 & w893;
assign w3358 = w761 & w917;
assign w3359 = ~w761 & w919;
assign w3360 = w3000 & w801;
assign w3361 = ~w760 & w3580;
assign w3362 = w3000 & ~w931;
assign w3363 = w3000 & ~w836;
assign w3364 = w3000 & w758;
assign w3365 = w761 & ~w1001;
assign w3366 = w3752 & ~pi11;
assign w3367 = w109 & w3581;
assign w3368 = w109 & w3582;
assign w3369 = pi05 & ~pi26;
assign w3370 = (~w98 & w2849) | (~w98 & ~w64) | (w2849 & ~w64);
assign w3371 = (~w199 & ~w194) | (~w199 & w3583) | (~w194 & w3583);
assign w3372 = ~w102 & w4202;
assign w3373 = (~w144 & w102) | (~w144 & w4203) | (w102 & w4203);
assign v678 = ~(w2465 | pi09);
assign w3374 = v678;
assign v679 = ~(w526 | w434);
assign w3375 = v679;
assign w3376 = ~w733 & w3584;
assign w3377 = (~w1090 & w989) | (~w1090 & w3585) | (w989 & w3585);
assign w3378 = (~w1101 & w989) | (~w1101 & w3586) | (w989 & w3586);
assign v680 = ~(pi23 | w3062);
assign w3379 = v680;
assign w3380 = pi05 & w1348;
assign w3381 = pi05 & ~w1348;
assign w3382 = pi05 & ~w3223;
assign w3383 = (pi05 & ~w2360) | (pi05 & w2837) | (~w2360 & w2837);
assign w3384 = ~w691 & w770;
assign w3385 = ~w601 & w770;
assign w3386 = ~w691 & w656;
assign v681 = ~(w2935 | w98);
assign w3387 = v681;
assign w3388 = ~w493 & pi17;
assign w3389 = ~w98 & w2721;
assign w3390 = w2721 & w3587;
assign w3391 = (pi07 & w102) | (pi07 & w3588) | (w102 & w3588);
assign w3392 = (w153 & w3589) | (w153 & w3590) | (w3589 & w3590);
assign w3393 = ~w140 & w194;
assign w3394 = ~w140 & w202;
assign w3395 = ~w3751 & w146;
assign w3396 = (w229 & w3591) | (w229 & w3592) | (w3591 & w3592);
assign w3397 = w347 & w2719;
assign w3398 = (w166 & w4204) | (w166 & w4205) | (w4204 & w4205);
assign w3399 = w353 & ~w2719;
assign w3400 = (w3594 & w166) | (w3594 & w4206) | (w166 & w4206);
assign w3401 = ~w162 & w3595;
assign w3402 = ~w602 & w3596;
assign w3403 = pi17 & w702;
assign w3404 = w2198 & pi13;
assign w3405 = ~w867 & pi11;
assign w3406 = w761 & ~w1013;
assign v682 = ~(w759 | w931);
assign w3407 = v682;
assign v683 = ~(w759 | w836);
assign w3408 = v683;
assign w3409 = ~w759 & w758;
assign v684 = ~(pi21 | w966);
assign w3410 = v684;
assign w3411 = (~pi21 & w3410) | (~pi21 & ~w761) | (w3410 & ~w761);
assign w3412 = w3017 & w857;
assign v685 = ~(w3017 | w857);
assign w3413 = v685;
assign w3414 = w574 & ~w3042;
assign w3415 = (w574 & w3597) | (w574 & w4361) | (w3597 & w4361);
assign w3416 = w52 & w50;
assign w3417 = ~pi09 & w174;
assign w3418 = ~w98 & w2938;
assign w3419 = w2721 & w3598;
assign w3420 = ~pi09 & pi01;
assign w3421 = (pi01 & ~w2) | (pi01 & w3599) | (~w2 & w3599);
assign w3422 = w3420 & ~w193;
assign w3423 = ~w197 & w3600;
assign w3424 = ~w197 & w3601;
assign w3425 = w140 & w202;
assign w3426 = (~w2765 & w3602) | (~w2765 & w3603) | (w3602 & w3603);
assign w3427 = (w2765 & w3372) | (w2765 & w3751) | (w3372 & w3751);
assign w3428 = w2926 & ~pi13;
assign w3429 = (w2960 & w146) | (w2960 & w3605) | (w146 & w3605);
assign w3430 = (w146 & w4207) | (w146 & w4208) | (w4207 & w4208);
assign w3431 = ~w69 & w3606;
assign w3432 = ~pi17 & w342;
assign w3433 = w2926 & w342;
assign w3434 = w320 & w3607;
assign w3435 = (~w335 & w3607) | (~w335 & w3608) | (w3607 & w3608);
assign w3436 = (~w2774 & w3609) | (~w2774 & w3610) | (w3609 & w3610);
assign v686 = ~(w306 | w2376);
assign w3437 = v686;
assign w3438 = ~w306 & w2773;
assign w3439 = (w2774 & w3437) | (w2774 & w3438) | (w3437 & w3438);
assign w3440 = w524 & ~pi17;
assign w3441 = ~w524 & pi17;
assign v687 = ~(pi05 | pi09);
assign w3442 = v687;
assign w3443 = ~w533 & w686;
assign w3444 = w581 & w589;
assign w3445 = ~w571 & w779;
assign w3446 = (~w434 & w3611) | (~w434 & w4343) | (w3611 & w4343);
assign w3447 = (w791 & w2996) | (w791 & w3612) | (w2996 & w3612);
assign w3448 = (w2181 & w3612) | (w2181 & w3613) | (w3612 & w3613);
assign w3449 = ~pi01 & pi14;
assign w3450 = (w2421 & w3614) | (w2421 & w3615) | (w3614 & w3615);
assign w3451 = (~pi07 & w611) | (~pi07 & w3616) | (w611 & w3616);
assign v688 = ~(pi07 | w3019);
assign w3452 = v688;
assign w3453 = ~w611 & w3617;
assign w3454 = pi07 & w3019;
assign w3455 = ~w611 & w3618;
assign w3456 = ~pi07 & w3019;
assign w3457 = w3017 & w854;
assign v689 = ~(w3017 | w854);
assign w3458 = v689;
assign w3459 = ~w2996 & w3619;
assign w3460 = (~w2181 & w3619) | (~w2181 & w3620) | (w3619 & w3620);
assign w3461 = ~w887 & pi10;
assign w3462 = (w3796 & w562) | (w3796 & w3621) | (w562 & w3621);
assign w3463 = ~pi23 & pi01;
assign w3464 = ~w914 & pi05;
assign w3465 = w914 & ~pi05;
assign w3466 = (pi09 & ~w3062) | (pi09 & w3622) | (~w3062 & w3622);
assign v690 = ~(w2465 | pi11);
assign w3467 = v690;
assign w3468 = w2465 & pi11;
assign w3469 = pi15 & ~w2480;
assign w3470 = ~pi23 & pi15;
assign w3471 = (~pi09 & ~w3062) | (~pi09 & w3623) | (~w3062 & w3623);
assign v691 = ~(pi23 | pi19);
assign w3472 = v691;
assign v692 = ~(w2477 | pi19);
assign w3473 = v692;
assign w3474 = w2470 & ~pi21;
assign w3475 = (~w2999 & ~pi21) | (~w2999 & w3624) | (~pi21 & w3624);
assign w3476 = w1075 & w783;
assign w3477 = ~w1277 & pi27;
assign w3478 = (pi27 & w1136) | (pi27 & w3477) | (w1136 & w3477);
assign w3479 = ~w1260 & w1259;
assign v693 = ~(w1277 | w434);
assign w3480 = v693;
assign w3481 = (~w434 & w1136) | (~w434 & w3480) | (w1136 & w3480);
assign w3482 = w1296 & w1259;
assign w3483 = ~w1190 & w1203;
assign w3484 = ~w1134 & w1203;
assign v694 = ~(pi04 | w1513);
assign w3485 = v694;
assign w3486 = (~pi21 & w1330) | (~pi21 & w3625) | (w1330 & w3625);
assign w3487 = (pi21 & w1330) | (pi21 & w3626) | (w1330 & w3626);
assign w3488 = w14 & pi27;
assign w3489 = (~w434 & w1313) | (~w434 & w3627) | (w1313 & w3627);
assign w3490 = (~pi25 & w1330) | (~pi25 & w3628) | (w1330 & w3628);
assign w3491 = w2353 & w1725;
assign w3492 = (~pi23 & w1631) | (~pi23 & w3629) | (w1631 & w3629);
assign v695 = ~(pi27 | w2506);
assign w3493 = v695;
assign w3494 = (~w1685 & w3630) | (~w1685 & w3631) | (w3630 & w3631);
assign w3495 = (w14 & w323) | (w14 & w3632) | (w323 & w3632);
assign w3496 = (w323 & w4209) | (w323 & w4210) | (w4209 & w4210);
assign w3497 = (~w1136 & w3634) | (~w1136 & w3635) | (w3634 & w3635);
assign w3498 = (w1300 & w3634) | (w1300 & w3636) | (w3634 & w3636);
assign w3499 = (w1289 & w3637) | (w1289 & w3638) | (w3637 & w3638);
assign w3500 = ~w323 & w4211;
assign w3501 = (w310 & w3640) | (w310 & w3641) | (w3640 & w3641);
assign w3502 = ~w323 & w4212;
assign w3503 = (w310 & w3643) | (w310 & w3644) | (w3643 & w3644);
assign w3504 = w1818 & ~w2010;
assign w3505 = ~w1818 & w1788;
assign w3506 = ~w323 & w4213;
assign w3507 = (w310 & w3646) | (w310 & w3647) | (w3646 & w3647);
assign w3508 = ~w323 & w4214;
assign w3509 = (w310 & w3649) | (w310 & w3650) | (w3649 & w3650);
assign w3510 = ~w1911 & w2054;
assign w3511 = w3701 & w128;
assign w3512 = (~pi11 & w3764) | (~pi11 & w4215) | (w3764 & w4215);
assign w3513 = (pi09 & w3764) | (pi09 & w4216) | (w3764 & w4216);
assign w3514 = (~pi09 & w3764) | (~pi09 & w4217) | (w3764 & w4217);
assign w3515 = (pi11 & w3764) | (pi11 & w4218) | (w3764 & w4218);
assign w3516 = (w572 & w4219) | (w572 & w4220) | (w4219 & w4220);
assign v696 = ~(w687 | pi13);
assign w3517 = v696;
assign w3518 = (w572 & w4221) | (w572 & w4222) | (w4221 & w4222);
assign v697 = ~(pi19 | w581);
assign w3519 = v697;
assign w3520 = (w310 & w3726) | (w310 & w3651) | (w3726 & w3651);
assign w3521 = (w2977 & w4223) | (w2977 & w4224) | (w4223 & w4224);
assign w3522 = (w809 & w577) | (w809 & w3654) | (w577 & w3654);
assign w3523 = (w809 & w560) | (w809 & w3655) | (w560 & w3655);
assign w3524 = (w310 & w3656) | (w310 & w3657) | (w3656 & w3657);
assign w3525 = (w2977 & w4225) | (w2977 & w4226) | (w4225 & w4226);
assign w3526 = w3062 & w3660;
assign w3527 = (w2749 & w4227) | (w2749 & w4228) | (w4227 & w4228);
assign w3528 = w3062 & w3661;
assign w3529 = w3662 & ~w1051;
assign w3530 = ~w2473 & w4147;
assign w3531 = ~w2470 & w4147;
assign v698 = ~(pi23 | w2420);
assign w3532 = v698;
assign w3533 = (w783 & w323) | (w783 & w3663) | (w323 & w3663);
assign w3534 = (w323 & w4229) | (w323 & w4230) | (w4229 & w4230);
assign w3535 = ~w989 & w3665;
assign w3536 = w1443 & pi19;
assign w3537 = w14 & ~pi05;
assign w3538 = ~w14 & pi05;
assign w3539 = ~w1631 & w3666;
assign w3540 = (w310 & w3737) | (w310 & w3667) | (w3737 & w3667);
assign w3541 = (~w2699 & w3668) | (~w2699 & w4357) | (w3668 & w4357);
assign w3542 = ~w2470 & pi21;
assign w3543 = ~w2473 & pi17;
assign w3544 = ~w1244 & pi21;
assign w3545 = w1244 & ~pi21;
assign w3546 = w344 & w324;
assign w3547 = (w146 & w3669) | (w146 & w3670) | (w3669 & w3670);
assign w3548 = (pi05 & w3249) | (pi05 & ~w415) | (w3249 & ~w415);
assign w3549 = (pi12 & w690) | (pi12 & w3671) | (w690 & w3671);
assign w3550 = w628 & pi12;
assign w3551 = ~w1330 & w3672;
assign w3552 = ~w3100 & w2591;
assign w3553 = w2633 & ~w908;
assign w3554 = (~w908 & w318) | (~w908 & w3673) | (w318 & w3673);
assign w3555 = (w2749 & w4231) | (w2749 & w4232) | (w4231 & w4232);
assign w3556 = (~pi13 & ~w3062) | (~pi13 & w3674) | (~w3062 & w3674);
assign w3557 = (pi13 & ~w3062) | (pi13 & w3675) | (~w3062 & w3675);
assign w3558 = w1695 & w2354;
assign w3559 = (pi31 & w323) | (pi31 & w3676) | (w323 & w3676);
assign w3560 = (w323 & w4233) | (w323 & w4234) | (w4233 & w4234);
assign w3561 = (~w14 & w323) | (~w14 & w3678) | (w323 & w3678);
assign w3562 = (w323 & w4235) | (w323 & w4236) | (w4235 & w4236);
assign w3563 = w1749 & ~w2506;
assign w3564 = (~w1685 & w3680) | (~w1685 & w3681) | (w3680 & w3681);
assign w3565 = (~w310 & w3682) | (~w310 & w3683) | (w3682 & w3683);
assign w3566 = ~w2477 & w4147;
assign v699 = ~(w1334 | w1423);
assign w3567 = v699;
assign v700 = ~(w1334 | pi13);
assign w3568 = v700;
assign w3569 = w1334 & pi13;
assign w3570 = ~w1334 & w1642;
assign w3571 = w1334 & ~pi17;
assign w3572 = w1428 & ~pi23;
assign w3573 = w1334 & pi27;
assign w3574 = ~w1428 & pi23;
assign w3575 = ~w1330 & w3684;
assign w3576 = ~w1712 & pi05;
assign w3577 = (~pi27 & ~w2298) | (~pi27 & w3685) | (~w2298 & w3685);
assign v701 = ~(pi27 | w1704);
assign w3578 = v701;
assign w3579 = w1334 & pi15;
assign w3580 = ~w759 & w801;
assign w3581 = ~pi17 & pi07;
assign w3582 = w2926 & pi07;
assign v702 = ~(w72 | w199);
assign w3583 = v702;
assign w3584 = (~w717 & w3686) | (~w717 & w3687) | (w3686 & w3687);
assign v703 = ~(w2472 | w1090);
assign w3585 = v703;
assign v704 = ~(w2472 | w1101);
assign w3586 = v704;
assign v705 = ~(pi09 | w98);
assign w3587 = v705;
assign w3588 = ~w140 & pi07;
assign w3589 = (pi07 & ~w2721) | (pi07 & w4362) | (~w2721 & w4362);
assign w3590 = ~w2332 & w3688;
assign w3591 = (w347 & ~w109) | (w347 & w3689) | (~w109 & w3689);
assign w3592 = (w153 & w3690) | (w153 & w3691) | (w3690 & w3691);
assign w3593 = (~w153 & w3692) | (~w153 & w3693) | (w3692 & w3693);
assign w3594 = (~w153 & w3694) | (~w153 & w3695) | (w3694 & w3695);
assign w3595 = (~pi09 & ~w163) | (~pi09 & w3696) | (~w163 & w3696);
assign w3596 = pi17 & ~w581;
assign w3597 = ~w3796 & w574;
assign w3598 = w174 & ~w98;
assign w3599 = pi20 & pi01;
assign w3600 = pi22 & pi01;
assign w3601 = pi22 & w3420;
assign w3602 = (pi09 & w102) | (pi09 & w3697) | (w102 & w3697);
assign w3603 = (w153 & w3698) | (w153 & w3699) | (w3698 & w3699);
assign w3604 = w2721 & w3700;
assign w3605 = w109 & w3428;
assign w3606 = w71 & ~w3751;
assign w3607 = (w166 & w4237) | (w166 & w4238) | (w4237 & w4238);
assign w3608 = pi01 & ~w2719;
assign w3609 = w320 & w3703;
assign w3610 = pi01 & ~w2773;
assign w3611 = (~w310 & w3704) | (~w310 & w3705) | (w3704 & w3705);
assign w3612 = (w310 & w4250) | (w310 & w4239) | (w4250 & w4239);
assign w3613 = (w2977 & w4240) | (w2977 & w4241) | (w4240 & w4241);
assign w3614 = (w805 & w577) | (w805 & w3707) | (w577 & w3707);
assign w3615 = (w805 & w560) | (w805 & w3708) | (w560 & w3708);
assign v706 = ~(w606 | pi07);
assign w3616 = v706;
assign w3617 = w606 & pi07;
assign w3618 = w606 & ~pi07;
assign w3619 = (~w310 & w3709) | (~w310 & w3710) | (w3709 & w3710);
assign w3620 = pi21 & w3446;
assign w3621 = ~w571 & w3796;
assign w3622 = pi23 & pi09;
assign w3623 = pi23 & ~pi09;
assign w3624 = ~pi21 & w2420;
assign w3625 = w1334 & ~pi21;
assign w3626 = w1334 & pi21;
assign v707 = ~(w3488 | w434);
assign w3627 = v707;
assign w3628 = w1334 & ~pi25;
assign w3629 = w2289 & w3711;
assign w3630 = (w310 & w3712) | (w310 & w3713) | (w3712 & w3713);
assign v708 = ~(pi27 | w3101);
assign w3631 = v708;
assign w3632 = ~w2633 & w14;
assign w3633 = ~w318 & w3714;
assign w3634 = ~w3132 & w434;
assign w3635 = (~w3132 & w1277) | (~w3132 & w3634) | (w1277 & w3634);
assign v709 = ~(w3132 | w3481);
assign w3636 = v709;
assign v710 = ~(w14 | w3481);
assign w3637 = v710;
assign w3638 = (w1300 & w3715) | (w1300 & w3637) | (w3715 & w3637);
assign w3639 = w2633 & pi11;
assign w3640 = ~w323 & w3639;
assign w3641 = w433 & w3717;
assign w3642 = w2633 & ~pi11;
assign w3643 = ~w323 & w3642;
assign w3644 = w433 & w3719;
assign w3645 = w2633 & ~pi17;
assign w3646 = ~w323 & w3645;
assign w3647 = w433 & w3721;
assign w3648 = w2633 & pi17;
assign w3649 = ~w323 & w3648;
assign w3650 = w433 & w3723;
assign w3651 = w433 & w3725;
assign w3652 = (w310 & w3726) | (w310 & w3727) | (w3726 & w3727);
assign w3653 = (w310 & w4242) | (w310 & w4243) | (w4242 & w4243);
assign w3654 = (w2977 & w4244) | (w2977 & w4245) | (w4244 & w4245);
assign w3655 = ~w3375 & w809;
assign w3656 = ~w908 & w3282;
assign w3657 = w433 & w3728;
assign w3658 = (w310 & w3656) | (w310 & w3729) | (w3656 & w3729);
assign w3659 = (w310 & w3730) | (w310 & w3731) | (w3730 & w3731);
assign w3660 = ~pi23 & pi09;
assign v711 = ~(pi23 | pi09);
assign w3661 = v711;
assign w3662 = (pi13 & ~w3062) | (pi13 & w3732) | (~w3062 & w3732);
assign w3663 = ~w2633 & w783;
assign w3664 = ~w318 & w3733;
assign w3665 = w2472 & ~w1278;
assign w3666 = (pi23 & ~w2289) | (pi23 & w3734) | (~w2289 & w3734);
assign w3667 = w433 & w3736;
assign w3668 = (w310 & w3737) | (w310 & w3738) | (w3737 & w3738);
assign w3669 = w2960 & w3247;
assign w3670 = w110 & w3247;
assign w3671 = w687 & pi12;
assign w3672 = ~w1334 & pi17;
assign w3673 = w320 & ~w908;
assign w3674 = pi23 & ~pi13;
assign w3675 = pi23 & pi13;
assign w3676 = ~w2633 & pi31;
assign w3677 = ~w318 & w3739;
assign v712 = ~(w2633 | w14);
assign w3678 = v712;
assign w3679 = ~w318 & w3740;
assign w3680 = (w310 & w3741) | (w310 & w3742) | (w3741 & w3742);
assign w3681 = w1749 & ~w3101;
assign w3682 = w907 & ~w3282;
assign w3683 = (w907 & ~w433) | (w907 & w3743) | (~w433 & w3743);
assign w3684 = ~w1334 & pi25;
assign w3685 = ~w1537 & w3744;
assign w3686 = ~w2996 & w3745;
assign w3687 = w907 & w2998;
assign w3688 = pi07 & ~w147;
assign w3689 = ~w3428 & w347;
assign w3690 = (~w146 & w4246) | (~w146 & w3747) | (w4246 & w3747);
assign w3691 = (w347 & w3747) | (w347 & w4363) | (w3747 & w4363);
assign w3692 = (w146 & w3748) | (w146 & w3749) | (w3748 & w3749);
assign w3693 = (w146 & w4247) | (w146 & w4248) | (w4247 & w4248);
assign w3694 = w353 & w3431;
assign w3695 = ~w69 & w3750;
assign v713 = ~(pi09 | w3427);
assign w3696 = v713;
assign w3697 = ~w140 & pi09;
assign w3698 = pi09 & ~w147;
assign w3699 = ~w2332 & w3698;
assign w3700 = ~pi09 & pi13;
assign w3701 = w109 & w3752;
assign w3702 = pi01 & w2955;
assign w3703 = pi01 & w324;
assign w3704 = (~pi19 & w323) | (~pi19 & w3753) | (w323 & w3753);
assign w3705 = (~pi19 & ~w433) | (~pi19 & w3754) | (~w433 & w3754);
assign w3706 = (w310 & w4249) | (w310 & w4250) | (w4249 & w4250);
assign w3707 = (w2977 & w4251) | (w2977 & w4252) | (w4251 & w4252);
assign w3708 = ~w3375 & w805;
assign w3709 = (pi21 & w323) | (pi21 & w3755) | (w323 & w3755);
assign w3710 = (pi21 & ~w433) | (pi21 & w3756) | (~w433 & w3756);
assign w3711 = (~pi23 & w1537) | (~pi23 & w4253) | (w1537 & w4253);
assign w3712 = ~w323 & w4254;
assign w3713 = ~pi27 & w2399;
assign w3714 = ~w320 & w14;
assign w3715 = ~w14 & w434;
assign w3716 = w320 & pi11;
assign w3717 = (pi11 & w318) | (pi11 & w3716) | (w318 & w3716);
assign w3718 = w320 & ~pi11;
assign w3719 = (~pi11 & w318) | (~pi11 & w3718) | (w318 & w3718);
assign w3720 = w320 & ~pi17;
assign w3721 = (~pi17 & w318) | (~pi17 & w3720) | (w318 & w3720);
assign w3722 = w320 & pi17;
assign w3723 = (pi17 & w318) | (pi17 & w3722) | (w318 & w3722);
assign w3724 = w2633 & w791;
assign w3725 = (w791 & w318) | (w791 & w4255) | (w318 & w4255);
assign w3726 = ~w323 & w3724;
assign w3727 = w791 & w2399;
assign w3728 = w3554 & ~w908;
assign w3729 = ~w908 & w3283;
assign w3730 = (pi19 & ~w908) | (pi19 & w3282) | (~w908 & w3282);
assign w3731 = (pi19 & ~w908) | (pi19 & w3283) | (~w908 & w3283);
assign w3732 = w3675 & pi13;
assign w3733 = ~w320 & w783;
assign w3734 = ~w1537 & w4256;
assign w3735 = w2633 & ~w2699;
assign w3736 = (~w2699 & w318) | (~w2699 & w4257) | (w318 & w4257);
assign w3737 = ~w323 & w3735;
assign w3738 = ~w2699 & w2399;
assign w3739 = ~w320 & pi31;
assign v714 = ~(w320 | w14);
assign w3740 = v714;
assign w3741 = ~w323 & w4258;
assign w3742 = w1749 & w2399;
assign w3743 = ~w3554 & w907;
assign w3744 = (~pi27 & w1330) | (~pi27 & w4259) | (w1330 & w4259);
assign w3745 = ~w434 & w907;
assign w3746 = pi09 & pi07;
assign w3747 = (w347 & ~w109) | (w347 & w4260) | (~w109 & w4260);
assign w3748 = w353 & w3605;
assign w3749 = w353 & w2960;
assign w3750 = w71 & w353;
assign w3751 = w2721 & ~pi09;
assign w3752 = w2926 & w111;
assign v715 = ~(w2633 | pi19);
assign w3753 = v715;
assign w3754 = ~w318 & w4261;
assign w3755 = ~w2633 & pi21;
assign w3756 = ~w318 & w4262;
assign w3757 = (w401 & ~w2414) | (w401 & ~w384) | (~w2414 & ~w384);
assign w3758 = (w1017 & ~w2214) | (w1017 & ~w945) | (~w2214 & ~w945);
assign w3759 = (w1669 & w1806) | (w1669 & w2563) | (w1806 & w2563);
assign w3760 = (~pi01 & w1295) | (~pi01 & ~w2246) | (w1295 & ~w2246);
assign w3761 = (~pi17 & w1295) | (~pi17 & ~w2268) | (w1295 & ~w2268);
assign w3762 = w3225 | ~w32;
assign w3763 = w3225 & ~w32;
assign w3764 = (pi17 & ~w2926) | (pi17 & ~w146) | (~w2926 & ~w146);
assign w3765 = w1116 & w2210;
assign w3766 = w1116 & w2217;
assign v716 = ~(w997 | w998);
assign w3767 = v716;
assign w3768 = ~w547 & pi17;
assign v717 = ~(w1161 | pi13);
assign w3769 = v717;
assign w3770 = ~w1161 & w3285;
assign w3771 = (w2749 & w4263) | (w2749 & w4264) | (w4263 & w4264);
assign v718 = ~(w1116 | w1196);
assign w3772 = v718;
assign w3773 = w19 & w13;
assign w3774 = w2760 & ~w98;
assign w3775 = (~w98 & w2760) | (~w98 & w92) | (w2760 & w92);
assign w3776 = w72 & ~w144;
assign v719 = ~(w141 | w221);
assign w3777 = v719;
assign v720 = ~(w149 | w222);
assign w3778 = v720;
assign w3779 = pi11 & ~w223;
assign v721 = ~(w235 | w231);
assign w3780 = v721;
assign w3781 = ~pi18 & w4364;
assign w3782 = ~pi18 & w2965;
assign w3783 = ~pi19 & w2976;
assign w3784 = ~pi19 & w2420;
assign w3785 = w575 & ~w526;
assign v722 = ~(w525 | w584);
assign w3786 = v722;
assign w3787 = ~w585 & pi17;
assign w3788 = ~w585 & w2168;
assign w3789 = (w634 & w2986) | (w634 & ~w532) | (w2986 & ~w532);
assign w3790 = (w634 & w2986) | (w634 & ~w2413) | (w2986 & ~w2413);
assign w3791 = ~w662 & pi09;
assign v723 = ~(w503 | pi11);
assign w3792 = v723;
assign w3793 = pi19 & w2976;
assign w3794 = pi19 & w2420;
assign w3795 = ~w732 & w780;
assign w3796 = w3062 & w16;
assign v724 = ~(w767 | w786);
assign w3797 = v724;
assign w3798 = (w639 & w3006) | (w639 & w2976) | (w3006 & w2976);
assign w3799 = (w639 & w3006) | (w639 & w2420) | (w3006 & w2420);
assign w3800 = (~w808 & w3008) | (~w808 & w2976) | (w3008 & w2976);
assign w3801 = (~w808 & w3008) | (~w808 & w2420) | (w3008 & w2420);
assign w3802 = w669 & ~w812;
assign w3803 = (~pi05 & w3016) | (~pi05 & ~w629) | (w3016 & ~w629);
assign w3804 = (~pi05 & w3016) | (~pi05 & w795) | (w3016 & w795);
assign w3805 = ~w606 & w611;
assign w3806 = ~w566 & w3805;
assign v725 = ~(w807 | w803);
assign w3807 = v725;
assign w3808 = (w910 & w786) | (w910 & w4265) | (w786 & w4265);
assign w3809 = (w772 & w4266) | (w772 & w4267) | (w4266 & w4267);
assign w3810 = (pi21 & ~w3267) | (pi21 & w4268) | (~w3267 & w4268);
assign w3811 = (w772 & w4269) | (w772 & w4270) | (w4269 & w4270);
assign w3812 = (w3035 & ~w3267) | (w3035 & w4271) | (~w3267 & w4271);
assign w3813 = ~w889 & w977;
assign w3814 = w968 & ~w978;
assign w3815 = ~w862 & w984;
assign w3816 = w862 & ~w874;
assign v726 = ~(w862 | w1020);
assign w3817 = v726;
assign w3818 = w1031 & w991;
assign w3819 = w889 & w789;
assign w3820 = (w1052 & w3040) | (w1052 & w3038) | (w3040 & w3038);
assign w3821 = (w1052 & w3040) | (w1052 & w2420) | (w3040 & w2420);
assign w3822 = (w3038 & w4272) | (w3038 & w4273) | (w4272 & w4273);
assign w3823 = (w2420 & w4272) | (w2420 & w4273) | (w4272 & w4273);
assign w3824 = ~w889 & w966;
assign w3825 = (~pi19 & w553) | (~pi19 & w4274) | (w553 & w4274);
assign w3826 = w991 & w1059;
assign w3827 = (pi01 & w3045) | (pi01 & w3038) | (w3045 & w3038);
assign w3828 = (pi01 & w3045) | (pi01 & w2420) | (w3045 & w2420);
assign w3829 = w793 & ~w881;
assign w3830 = ~w793 & w881;
assign w3831 = ~w1127 & w1131;
assign w3832 = w1034 & w4078;
assign w3833 = w1127 & ~w1131;
assign w3834 = (w1127 & ~w1034) | (w1127 & w4079) | (~w1034 & w4079);
assign w3835 = ~w1134 & w1120;
assign w3836 = ~w1134 & w1086;
assign w3837 = (~w4147 & ~w1151) | (~w4147 & w4080) | (~w1151 & w4080);
assign w3838 = ~w1152 & w1035;
assign v727 = ~(w1075 | w1154);
assign w3839 = v727;
assign w3840 = (~w4147 & w1151) | (~w4147 & w4081) | (w1151 & w4081);
assign w3841 = ~w1159 & w1035;
assign w3842 = (pi15 & w3053) | (pi15 & w3038) | (w3053 & w3038);
assign w3843 = (pi15 & w3053) | (pi15 & w2420) | (w3053 & w2420);
assign w3844 = w1198 & w924;
assign w3845 = w1201 & ~w4147;
assign w3846 = w1201 & w1035;
assign v728 = ~(w989 | w980);
assign w3847 = v728;
assign w3848 = (~pi19 & w3055) | (~pi19 & w3038) | (w3055 & w3038);
assign w3849 = (~pi19 & w3055) | (~pi19 & w2420) | (w3055 & w2420);
assign w3850 = (~pi21 & w3796) | (~pi21 & w3038) | (w3796 & w3038);
assign w3851 = (~pi21 & w3796) | (~pi21 & w2420) | (w3796 & w2420);
assign w3852 = w1062 & pi23;
assign v729 = ~(w1062 | pi23);
assign w3853 = v729;
assign w3854 = ~w1189 & w1288;
assign w3855 = w1304 & w1314;
assign w3856 = ~w1189 & w1317;
assign w3857 = w2243 | ~w1259;
assign w3858 = (~w1259 & w2243) | (~w1259 & w1189) | (w2243 & w1189);
assign w3859 = w1304 & ~w1332;
assign w3860 = w4034 & w4275;
assign w3861 = (~pi05 & ~w4034) | (~pi05 & w4276) | (~w4034 & w4276);
assign w3862 = (pi05 & ~w4034) | (pi05 & w4277) | (~w4034 & w4277);
assign w3863 = ~w1049 & w1053;
assign w3864 = ~w1049 & w1035;
assign w3865 = w1130 & w4278;
assign w3866 = w1124 & w1035;
assign w3867 = ~w1289 & w4082;
assign v730 = ~(w1139 | w4147);
assign w3868 = v730;
assign w3869 = ~w1139 & w1035;
assign v731 = ~(w1417 | w1148);
assign w3870 = v731;
assign v732 = ~(w1417 | w3069);
assign w3871 = v732;
assign w3872 = ~w1189 & w1220;
assign v733 = ~(w1292 | w1256);
assign w3873 = v733;
assign v734 = ~(w1189 | w1174);
assign w3874 = v734;
assign v735 = ~(w1151 | w4147);
assign w3875 = v735;
assign w3876 = ~w1151 & w1035;
assign w3877 = w1457 & pi13;
assign v736 = ~(w1457 | pi13);
assign w3878 = v736;
assign w3879 = ~w1313 & w4279;
assign w3880 = w1338 & w2245;
assign w3881 = pi02 & pi04;
assign w3882 = (~w1513 & w3086) | (~w1513 & w1314) | (w3086 & w1314);
assign w3883 = (~w1513 & w3086) | (~w1513 & w2245) | (w3086 & w2245);
assign w3884 = w1536 & ~w1450;
assign w3885 = w1536 & ~w1496;
assign w3886 = w1457 & pi15;
assign v737 = ~(w1457 | pi15);
assign w3887 = v737;
assign w3888 = ~w1609 & w1540;
assign v738 = ~(w1609 | w1614);
assign w3889 = v738;
assign w3890 = (pi19 & ~w1541) | (pi19 & w4280) | (~w1541 & w4280);
assign v739 = ~(w1623 | w1541);
assign w3891 = v739;
assign w3892 = w1623 & ~w1541;
assign w3893 = w1686 & w2506;
assign w3894 = (w2506 & w1686) | (w2506 & w1693) | (w1686 & w1693);
assign w3895 = w2296 & w4083;
assign w3896 = w1733 & ~w1732;
assign w3897 = w1733 & ~w2509;
assign w3898 = w2510 | w2511;
assign w3899 = (w2511 & w2510) | (w2511 & w1721) | (w2510 & w1721);
assign w3900 = w2514 | w2515;
assign w3901 = (w2515 & w2514) | (w2515 & w1721) | (w2514 & w1721);
assign w3902 = w1783 & ~w1602;
assign w3903 = w1783 & ~w1557;
assign v740 = ~(w1646 | w1603);
assign w3904 = v740;
assign v741 = ~(w1646 | w1557);
assign w3905 = v741;
assign w3906 = w2526 | w2527;
assign w3907 = (w2527 & w2526) | (w2527 & w1721) | (w2526 & w1721);
assign w3908 = ~w1567 & w1554;
assign w3909 = ~w1567 & w1545;
assign w3910 = w2531 | w2532;
assign w3911 = (w2532 & w2531) | (w2532 & w1721) | (w2531 & w1721);
assign v742 = ~(w1807 | w1824);
assign w3912 = v742;
assign w3913 = w1738 & ~w1825;
assign w3914 = w1656 & ~w1664;
assign v743 = ~(w1843 | w1846);
assign w3915 = v743;
assign w3916 = w1922 & w1934;
assign w3917 = w2564 | w2565;
assign w3918 = (w2565 & w2564) | (w2565 & w1721) | (w2564 & w1721);
assign v744 = ~(pi11 | pi31);
assign w3919 = v744;
assign v745 = ~(pi11 | w2698);
assign w3920 = v745;
assign v746 = ~(pi17 | pi31);
assign w3921 = v746;
assign v747 = ~(pi17 | w2698);
assign w3922 = v747;
assign w3923 = pi17 & ~pi31;
assign w3924 = pi17 & ~w2698;
assign w3925 = w1830 & ~w2046;
assign w3926 = w1830 & w2055;
assign w3927 = (w42 & w4281) | (w42 & w4282) | (w4281 & w4282);
assign w3928 = (w124 & w2331) | (w124 & ~w115) | (w2331 & ~w115);
assign v748 = ~(w3052 | w1176);
assign w3929 = v748;
assign w3930 = ~w888 & w4283;
assign w3931 = ~w2474 & w1238;
assign w3932 = w3056 & w4147;
assign w3933 = (w3208 & ~w434) | (w3208 & w3038) | (~w434 & w3038);
assign w3934 = (w3208 & ~w434) | (w3208 & w2420) | (~w434 & w2420);
assign w3935 = w1296 & w1301;
assign w3936 = w1296 & ~w1365;
assign w3937 = (w1372 & w1257) | (w1372 & w4284) | (w1257 & w4284);
assign w3938 = (~w1460 & w1257) | (~w1460 & w4285) | (w1257 & w4285);
assign w3939 = ~w1257 & w4286;
assign w3940 = w2717 & w2718;
assign w3941 = (w2718 & w2717) | (w2718 & ~w1721) | (w2717 & ~w1721);
assign w3942 = w3206 & pi21;
assign w3943 = w3205 & pi17;
assign v749 = ~(w1296 | w1233);
assign w3944 = v749;
assign w3945 = ~w1296 & w1375;
assign v750 = ~(w1296 | w1386);
assign w3946 = v750;
assign w3947 = ~w1296 & w1403;
assign w3948 = (pi21 & w3235) | (pi21 & ~w1294) | (w3235 & ~w1294);
assign w3949 = (pi21 & w3235) | (pi21 & ~w2658) | (w3235 & ~w2658);
assign w3950 = ~w219 & pi09;
assign w3951 = w219 & ~pi09;
assign w3952 = w2633 & ~w321;
assign w3953 = w2335 & w459;
assign v751 = ~(w2335 | w459);
assign w3954 = v751;
assign w3955 = ~w483 & w577;
assign w3956 = w781 & ~w909;
assign v752 = ~(w1113 | w4147);
assign w3957 = v752;
assign w3958 = ~w1113 & w2237;
assign w3959 = w2597 & w2598;
assign w3960 = (w2598 & w2597) | (w2598 & ~w1721) | (w2597 & ~w1721);
assign w3961 = w2606 & w2607;
assign w3962 = (w2607 & w2606) | (w2607 & ~w1721) | (w2606 & ~w1721);
assign w3963 = w2611 & w2612;
assign w3964 = (w2612 & w2611) | (w2612 & ~w1721) | (w2611 & ~w1721);
assign w3965 = pi16 & ~w109;
assign w3966 = ~pi15 & w4147;
assign w3967 = ~pi15 & w3201;
assign w3968 = (~w1173 & w1257) | (~w1173 & w4287) | (w1257 & w4287);
assign w3969 = w1695 & w1743;
assign w3970 = w484 & w672;
assign w3971 = ~w746 & pi15;
assign w3972 = w746 & ~pi15;
assign w3973 = w3062 & w4288;
assign w3974 = w828 & pi09;
assign v753 = ~(w828 | pi09);
assign w3975 = v753;
assign w3976 = w2029 & w1788;
assign w3977 = w2029 & ~w1767;
assign w3978 = w2031 & ~w1788;
assign w3979 = w2031 & w1767;
assign v754 = ~(w761 | w896);
assign w3980 = v754;
assign w3981 = (~w1090 & w961) | (~w1090 & w4289) | (w961 & w4289);
assign w3982 = ~w1877 & pi31;
assign w3983 = ~w278 & w4290;
assign w3984 = w279 & w4365;
assign w3985 = pi07 & ~w282;
assign w3986 = pi07 & ~w2372;
assign v755 = ~(w267 | w32);
assign w3987 = v755;
assign v756 = ~(w267 | w2370);
assign w3988 = v756;
assign w3989 = w267 & w32;
assign w3990 = w267 & w2370;
assign v757 = ~(w575 | w434);
assign w3991 = v757;
assign w3992 = ~w1113 & w2209;
assign w3993 = w1049 & pi05;
assign w3994 = ~w1113 & w1131;
assign w3995 = (~w1142 & ~w1112) | (~w1142 & w4291) | (~w1112 & w4291);
assign w3996 = w2818 | w1126;
assign w3997 = (w1126 & w2818) | (w1126 & w1113) | (w2818 & w1113);
assign v758 = ~(w1156 | w1155);
assign w3998 = v758;
assign w3999 = (~w1182 & ~w1112) | (~w1182 & w4292) | (~w1112 & w4292);
assign w4000 = ~w1062 & w3379;
assign w4001 = w325 & ~w32;
assign w4002 = w325 & ~w2370;
assign w4003 = w1361 & ~w2658;
assign w4004 = w219 & w28;
assign w4005 = ~w229 & w4293;
assign w4006 = w327 & w2370;
assign w4007 = w3398 & w319;
assign w4008 = w3398 & w2140;
assign w4009 = (w3398 & ~w2719) | (w3398 & w4294) | (~w2719 & w4294);
assign w4010 = (w3398 & w3399) | (w3398 & ~w334) | (w3399 & ~w334);
assign w4011 = (w3400 & w241) | (w3400 & w4295) | (w241 & w4295);
assign w4012 = w3401 & ~w244;
assign w4013 = w3401 & w2125;
assign w4014 = ~w571 & pi19;
assign w4015 = w219 & ~pi11;
assign v759 = ~(w444 | w109);
assign w4016 = v759;
assign w4017 = (pi14 & w3449) | (pi14 & ~w532) | (w3449 & ~w532);
assign w4018 = (pi14 & w3449) | (pi14 & ~w2413) | (w3449 & ~w2413);
assign w4019 = ~w637 & pi14;
assign v760 = ~(pi05 | w3003);
assign w4020 = v760;
assign v761 = ~(pi05 | w3004);
assign w4021 = v761;
assign w4022 = pi01 & ~w580;
assign w4023 = ~w578 & w4022;
assign w4024 = ~w1113 & w1053;
assign w4025 = ~w1113 & w1089;
assign w4026 = ~w1218 & w1441;
assign w4027 = (pi15 & w959) | (pi15 & w4296) | (w959 & w4296);
assign w4028 = (w959 & w4297) | (w959 & w4298) | (w4297 & w4298);
assign v762 = ~(w1524 | pi05);
assign w4029 = v762;
assign v763 = ~(w434 | w3133);
assign w4030 = v763;
assign v764 = ~(w434 | w3134);
assign w4031 = v764;
assign v765 = ~(w660 | w667);
assign w4032 = v765;
assign w4033 = (~w2916 & w2468) | (~w2916 & ~w2915) | (w2468 & ~w2915);
assign w4034 = (~w1089 & ~w1035) | (~w1089 & ~w3068) | (~w1035 & ~w3068);
assign w4035 = (~w1053 & ~w1035) | (~w1053 & ~w3047) | (~w1035 & ~w3047);
assign w4036 = (~w1131 & ~w1035) | (~w1131 & ~w2816) | (~w1035 & ~w2816);
assign w4037 = (w1249 & w1361) | (w1249 & w4003) | (w1361 & w4003);
assign w4038 = (pi05 & w3199) | (pi05 & w1113) | (w3199 & w1113);
assign w4039 = ~w107 & w2117;
assign w4040 = w104 & w164;
assign w4041 = ~w172 & w226;
assign w4042 = (w2765 & w4299) | (w2765 & w4300) | (w4299 & w4300);
assign w4043 = w120 & w173;
assign w4044 = (pi22 & w2867) | (pi22 & ~w173) | (w2867 & ~w173);
assign w4045 = (w2763 & w4301) | (w2763 & w4302) | (w4301 & w4302);
assign w4046 = ~w357 & pi20;
assign w4047 = w274 & w4303;
assign w4048 = w434 & w2960;
assign w4049 = ~w571 & w578;
assign w4050 = w2169 | ~w582;
assign w4051 = (~w582 & w2169) | (~w582 & w560) | (w2169 & w560);
assign w4052 = ~w690 & w3185;
assign v766 = ~(w778 | w964);
assign w4053 = v766;
assign v767 = ~(w778 | w872);
assign w4054 = v767;
assign w4055 = (w967 & w2469) | (w967 & w964) | (w2469 & w964);
assign w4056 = (w967 & w2469) | (w967 & w872) | (w2469 & w872);
assign w4057 = w973 & ~w964;
assign w4058 = w973 & ~w872;
assign v768 = ~(w902 | w985);
assign w4059 = v768;
assign w4060 = (w902 & w4304) | (w902 & w4305) | (w4304 & w4305);
assign w4061 = (w902 & w4306) | (w902 & w4307) | (w4306 & w4307);
assign w4062 = ~w949 & w1198;
assign w4063 = ~w1027 & w3056;
assign w4064 = ~w1027 & w3932;
assign v769 = ~(w2079 | w2077);
assign w4065 = v769;
assign w4066 = ~w989 & w3232;
assign w4067 = ~w989 & w3942;
assign w4068 = ~w997 & w3233;
assign w4069 = ~w997 & w3943;
assign w4070 = (w2834 & ~w1298) | (w2834 & w4308) | (~w1298 & w4308);
assign w4071 = (~w1294 & w2834) | (~w1294 & ~w2250) | (w2834 & ~w2250);
assign w4072 = w1684 & ~w1505;
assign w4073 = w1684 & ~w2273;
assign w4074 = (w2591 & w3279) | (w2591 & w1684) | (w3279 & w1684);
assign w4075 = (w4073 & w4309) | (w4073 & w4310) | (w4309 & w4310);
assign w4076 = w1115 & w3993;
assign w4077 = (w3993 & w1115) | (w3993 & w1049) | (w1115 & w1049);
assign v770 = ~(w1127 | w963);
assign w4078 = v770;
assign w4079 = w962 & w4366;
assign w4080 = pi11 & ~w4147;
assign v771 = ~(pi11 | w4147);
assign w4081 = v771;
assign w4082 = w1391 & ~pi07;
assign w4083 = (~pi27 & w1537) | (~pi27 & w4312) | (w1537 & w4312);
assign w4084 = w2212 & ~w1161;
assign w4085 = (w1115 & w4313) | (w1115 & w4314) | (w4313 & w4314);
assign w4086 = w1290 & ~w3481;
assign w4087 = (w1300 & w4315) | (w1300 & w4086) | (w4315 & w4086);
assign w4088 = pi11 & w1388;
assign w4089 = pi11 & ~w1398;
assign w4090 = ~w1514 & w1505;
assign w4091 = ~w1514 & w2273;
assign v772 = ~(w1515 | w1512);
assign w4092 = v772;
assign w4093 = w1521 & ~w1505;
assign w4094 = w1521 & ~w2273;
assign w4095 = (~w434 & w3101) | (~w434 & w1684) | (w3101 & w1684);
assign w4096 = (w4073 & w4316) | (w4073 & w4317) | (w4316 & w4317);
assign w4097 = (~w1338 & ~w1506) | (~w1338 & ~w1330) | (~w1506 & ~w1330);
assign v773 = ~(w79 | w103);
assign w4098 = v773;
assign v774 = ~(w79 | w2116);
assign w4099 = v774;
assign w4100 = ~w100 & w4318;
assign w4101 = (w128 & w2118) | (w128 & w107) | (w2118 & w107);
assign w4102 = w211 & w179;
assign w4103 = w211 & w173;
assign w4104 = ~w206 & w215;
assign v775 = ~(w218 | w147);
assign w4105 = v775;
assign v776 = ~(w218 | w141);
assign w4106 = v776;
assign w4107 = w104 & w2950;
assign w4108 = w210 & ~w173;
assign w4109 = (w2721 & w2139) | (w2721 & w226) | (w2139 & w226);
assign w4110 = (w2721 & w2139) | (w2721 & ~w216) | (w2139 & ~w216);
assign w4111 = w220 & pi11;
assign w4112 = (w2774 & w4319) | (w2774 & w4320) | (w4319 & w4320);
assign w4113 = pi18 & ~w2965;
assign w4114 = w434 & ~pi17;
assign w4115 = w110 | w109;
assign w4116 = (w109 & w110) | (w109 & w434) | (w110 & w434);
assign w4117 = w434 & w110;
assign w4118 = w621 & w593;
assign w4119 = w621 & w551;
assign w4120 = ~pi07 & w532;
assign w4121 = ~pi07 & w2413;
assign v777 = ~(w661 | w663);
assign w4122 = v777;
assign w4123 = ~w673 & w593;
assign w4124 = ~w673 & w551;
assign w4125 = w693 & ~w603;
assign w4126 = w693 & ~w714;
assign w4127 = w702 & ~w693;
assign w4128 = w2178 & ~w766;
assign w4129 = (~w766 & w2178) | (~w766 & ~w693) | (w2178 & ~w693);
assign w4130 = ~w566 & w4321;
assign w4131 = w445 & w551;
assign w4132 = w600 & w579;
assign w4133 = w811 & ~w809;
assign w4134 = w811 & ~w2185;
assign w4135 = (w2649 & w2650) | (w2649 & ~w786) | (w2650 & ~w786);
assign w4136 = (w2649 & w2650) | (w2649 & w764) | (w2650 & w764);
assign w4137 = (pi21 & w725) | (pi21 & w4322) | (w725 & w4322);
assign w4138 = pi21 & w764;
assign w4139 = w760 & ~w749;
assign w4140 = w862 & w1024;
assign w4141 = w1048 & ~w1056;
assign w4142 = ~w1048 & w1056;
assign w4143 = w2181 & w4323;
assign w4144 = (w2917 & w2918) | (w2917 & ~w693) | (w2918 & ~w693);
assign w4145 = (w2919 & w4324) | (w2919 & w4325) | (w4324 & w4325);
assign w4146 = ~pi23 & w4368;
assign v778 = ~(w783 | w1051);
assign w4147 = v778;
assign w4148 = ~w1174 & w1244;
assign v779 = ~(w1431 | w1428);
assign w4149 = v779;
assign w4150 = w1208 & ~w1475;
assign w4151 = w2274 & w1332;
assign w4152 = w2274 & w2659;
assign w4153 = (pi05 & w2275) | (pi05 & ~w1332) | (w2275 & ~w1332);
assign w4154 = (pi05 & w2275) | (pi05 & ~w2659) | (w2275 & ~w2659);
assign w4155 = w1380 & ~w1208;
assign v780 = ~(w1617 | w1671);
assign w4156 = v780;
assign w4157 = (pi05 & w1721) | (pi05 & w4326) | (w1721 & w4326);
assign w4158 = (pi05 & w2689) | (pi05 & w1714) | (w2689 & w1714);
assign w4159 = ~w2008 & w4327;
assign w4160 = w2009 & ~w3149;
assign v781 = ~(w2080 | w1831);
assign w4161 = v781;
assign v782 = ~(w2080 | w2079);
assign w4162 = v782;
assign w4163 = w3194 & w3193;
assign w4164 = (w3193 & w3194) | (w3193 & ~w693) | (w3194 & ~w693);
assign w4165 = (pi21 & w2349) | (pi21 & w1207) | (w2349 & w1207);
assign w4166 = (pi21 & w2349) | (pi21 & w3857) | (w2349 & w3857);
assign w4167 = ~w1670 & w1658;
assign w4168 = w1670 & ~w1658;
assign w4169 = w2451 & ~w788;
assign w4170 = w109 & w3366;
assign v783 = ~(w1244 | w1258);
assign w4171 = v783;
assign w4172 = w767 & w783;
assign w4173 = w434 & w3796;
assign w4174 = w668 & w727;
assign w4175 = w3448 & w3447;
assign w4176 = (w3447 & w3448) | (w3447 & ~w693) | (w3448 & ~w693);
assign w4177 = w797 & ~w580;
assign w4178 = w797 & w2422;
assign w4179 = w2451 & ~pi05;
assign v784 = ~(w2451 | pi05);
assign w4180 = v784;
assign w4181 = ~w2451 & pi05;
assign w4182 = w2451 & pi05;
assign w4183 = w434 & w1050;
assign v785 = ~(w434 | w1935);
assign w4184 = v785;
assign w4185 = ~w434 & w2566;
assign w4186 = (pi09 & w3526) | (pi09 & w3038) | (w3526 & w3038);
assign w4187 = (pi09 & w3526) | (pi09 & w2420) | (w3526 & w2420);
assign w4188 = (~pi09 & w3528) | (~pi09 & w3038) | (w3528 & w3038);
assign w4189 = (~pi09 & w3528) | (~pi09 & w2420) | (w3528 & w2420);
assign w4190 = pi07 & ~w109;
assign w4191 = w146 & w3762;
assign w4192 = (~pi15 & w2992) | (~pi15 & w2976) | (w2992 & w2976);
assign w4193 = (~pi15 & w2992) | (~pi15 & w2420) | (w2992 & w2420);
assign w4194 = w1695 & w1845;
assign w4195 = w2633 & w3554;
assign v786 = ~(pi17 | w1038);
assign w4196 = v786;
assign w4197 = ~pi17 & w2213;
assign v787 = ~(pi17 | w2658);
assign w4198 = v787;
assign w4199 = w1673 & ~pi25;
assign w4200 = ~w1673 & pi25;
assign w4201 = w668 & w785;
assign w4202 = w140 & ~pi09;
assign v788 = ~(w140 | w144);
assign w4203 = v788;
assign w4204 = w3593 | w3748;
assign w4205 = (w3748 & w3593) | (w3748 & w228) | (w3593 & w228);
assign w4206 = w228 & w3594;
assign w4207 = w2960 & ~pi13;
assign w4208 = w2960 & ~w3604;
assign w4209 = w3633 | w14;
assign w4210 = (w14 & w3633) | (w14 & ~w2633) | (w3633 & ~w2633);
assign w4211 = w2633 & w3717;
assign w4212 = w2633 & w3719;
assign w4213 = w2633 & w3721;
assign w4214 = w2633 & w3723;
assign v789 = ~(pi11 | w109);
assign w4215 = v789;
assign w4216 = pi09 & ~w109;
assign v790 = ~(pi09 | w109);
assign w4217 = v790;
assign w4218 = pi11 & ~w109;
assign v791 = ~(pi17 | w580);
assign w4219 = v791;
assign w4220 = ~pi17 & w2422;
assign w4221 = pi19 & ~w580;
assign w4222 = pi19 & w2422;
assign w4223 = (w3652 & w3653) | (w3652 & w2976) | (w3653 & w2976);
assign w4224 = (w3652 & w3653) | (w3652 & w2420) | (w3653 & w2420);
assign w4225 = (w3659 & w3658) | (w3659 & w2976) | (w3658 & w2976);
assign w4226 = (w3659 & w3658) | (w3659 & w2420) | (w3658 & w2420);
assign w4227 = w4147 & ~w2455;
assign w4228 = w4147 & w2748;
assign w4229 = w3664 | w783;
assign w4230 = (w783 & w3664) | (w783 & ~w2633) | (w3664 & ~w2633);
assign v792 = ~(pi15 | w2455);
assign w4231 = v792;
assign w4232 = ~pi15 & w2748;
assign w4233 = w3677 | pi31;
assign w4234 = (pi31 & w3677) | (pi31 & ~w2633) | (w3677 & ~w2633);
assign w4235 = w3679 | ~w14;
assign w4236 = (~w14 & w3679) | (~w14 & ~w2633) | (w3679 & ~w2633);
assign w4237 = w3702 | w3701;
assign w4238 = (w3701 & w3702) | (w3701 & w228) | (w3702 & w228);
assign w4239 = w791 | w3651;
assign w4240 = (w791 & w3706) | (w791 & w2976) | (w3706 & w2976);
assign w4241 = (w791 & w3706) | (w791 & w2420) | (w3706 & w2420);
assign w4242 = w791 & ~w3704;
assign w4243 = w791 & ~w3705;
assign w4244 = w434 & w3800;
assign w4245 = w434 & w3801;
assign w4246 = w347 & ~w3605;
assign w4247 = w3749 & ~pi13;
assign w4248 = w3749 & ~w3604;
assign w4249 = w791 | w3727;
assign w4250 = w791 | w3726;
assign w4251 = w434 & w3798;
assign w4252 = w434 & w3799;
assign w4253 = w1335 & ~pi23;
assign w4254 = w2633 & ~pi27;
assign w4255 = w320 & w791;
assign w4256 = ~w1335 & pi23;
assign w4257 = w320 & ~w2699;
assign w4258 = w2633 & w1749;
assign w4259 = w1334 & ~pi27;
assign w4260 = ~w2926 & w347;
assign v793 = ~(w320 | pi19);
assign w4261 = v793;
assign w4262 = ~w320 & pi21;
assign v794 = ~(pi13 | w2455);
assign w4263 = v794;
assign w4264 = ~pi13 & w2748;
assign w4265 = ~w780 & w910;
assign w4266 = pi21 & w3055;
assign w4267 = pi21 & w783;
assign w4268 = w718 & pi21;
assign w4269 = w3035 & w3055;
assign w4270 = w3035 & w783;
assign w4271 = w718 & w3035;
assign w4272 = pi05 & w1052;
assign w4273 = pi05 & w3040;
assign w4274 = pi17 & ~pi19;
assign w4275 = pi08 & pi05;
assign v795 = ~(pi08 | pi05);
assign w4276 = v795;
assign w4277 = ~pi08 & pi05;
assign w4278 = ~w1129 & w1124;
assign w4279 = w14 & w1338;
assign w4280 = w1499 & pi19;
assign w4281 = w124 | w3222;
assign w4282 = w124 | w3221;
assign w4283 = w2466 & w4147;
assign w4284 = ~w1244 & w1372;
assign v796 = ~(w1244 | w1460);
assign w4285 = v796;
assign w4286 = w1244 & pi17;
assign v797 = ~(w1244 | w1173);
assign w4287 = v797;
assign w4288 = w3472 & ~pi21;
assign w4289 = w949 & ~w1090;
assign w4290 = ~w276 & w275;
assign w4291 = w1141 & ~w1142;
assign w4292 = w1181 & ~w1182;
assign w4293 = w2956 & w32;
assign w4294 = w353 | w3398;
assign w4295 = ~w333 & w3400;
assign w4296 = w950 & pi15;
assign w4297 = pi15 & w4147;
assign w4298 = pi15 & w3930;
assign w4299 = w120 & w141;
assign w4300 = w120 & w2764;
assign w4301 = w2867 & pi22;
assign w4302 = (pi22 & w2867) | (pi22 & w3373) | (w2867 & w3373);
assign v798 = ~(w236 | pi20);
assign w4303 = v798;
assign w4304 = w1053 & w971;
assign w4305 = w1053 & w2203;
assign w4306 = ~w1099 & w971;
assign w4307 = ~w1099 & w2203;
assign w4308 = ~w2715 & w2834;
assign w4309 = (w2591 & w3279) | (w2591 & ~w1502) | (w3279 & ~w1502);
assign w4310 = (w2591 & w3279) | (w2591 & w4072) | (w3279 & w4072);
assign w4311 = w1127 & w924;
assign w4312 = w1335 & ~pi27;
assign w4313 = w2212 | ~w1161;
assign w4314 = (~w1161 & w2212) | (~w1161 & w1113) | (w2212 & w1113);
assign w4315 = w1290 & w434;
assign w4316 = (~w434 & w3101) | (~w434 & ~w1502) | (w3101 & ~w1502);
assign w4317 = (~w434 & w3101) | (~w434 & w4072) | (w3101 & w4072);
assign w4318 = w3175 & w128;
assign w4319 = pi18 & ~w3435;
assign w4320 = pi18 & ~w3434;
assign w4321 = w533 & w445;
assign w4322 = ~w771 & pi21;
assign w4323 = pi19 & w2917;
assign w4324 = ~pi23 & w574;
assign w4325 = ~pi23 & w1071;
assign w4326 = w3337 & pi05;
assign w4327 = ~w1818 & w2010;
assign w4328 = w228 & w2865;
assign w4329 = w228 & w2956;
assign w4330 = w359 & pi05;
assign v799 = ~(w359 | pi05);
assign w4331 = v799;
assign w4332 = ~w1256 & w1287;
assign w4333 = ~w1431 & w2264;
assign v800 = ~(w1438 | w1449);
assign w4334 = v800;
assign w4335 = ~w1522 & w1531;
assign w4336 = w1522 & ~w1531;
assign w4337 = w2356 & w1834;
assign w4338 = (w1834 & w2356) | (w1834 & w1666) | (w2356 & w1666);
assign w4339 = ~w1666 & w2357;
assign v801 = ~(w1695 | w1800);
assign w4340 = v801;
assign w4341 = (w179 & w173) | (w179 & ~w2864) | (w173 & ~w2864);
assign w4342 = (~w177 & w210) | (~w177 & w4108) | (w210 & w4108);
assign w4343 = (~w2976 & ~w2420) | (~w2976 & ~w2977) | (~w2420 & ~w2977);
assign w4344 = (~pi15 & w2926) | (~pi15 & ~w435) | (w2926 & ~w435);
assign w4345 = (w629 & ~w795) | (w629 & ~w3014) | (~w795 & ~w3014);
assign w4346 = (~w1100 & ~w3046) | (~w1100 & ~w1051) | (~w3046 & ~w1051);
assign w4347 = (~w1288 & w1380) | (~w1288 & w4155) | (w1380 & w4155);
assign w4348 = (w1439 & ~w2297) | (w1439 & ~w1502) | (~w2297 & ~w1502);
assign w4349 = (~w2870 & ~w2869) | (~w2870 & ~w2774) | (~w2869 & ~w2774);
assign w4350 = (~w2963 & ~w2964) | (~w2963 & ~w146) | (~w2964 & ~w146);
assign w4351 = (~w1505 & ~w2273) | (~w1505 & ~w1502) | (~w2273 & ~w1502);
assign w4352 = (~w32 & w3225) | (~w32 & ~w330) | (w3225 & ~w330);
assign w4353 = (w137 & ~pi09) | (w137 & w3372) | (~pi09 & w3372);
assign w4354 = pi22 & w4369;
assign w4355 = (w71 & w3606) | (w71 & ~w153) | (w3606 & ~w153);
assign w4356 = (~w3433 & ~w3432) | (~w3433 & ~w146) | (~w3432 & ~w146);
assign w4357 = (w3133 & w3134) | (w3133 & ~w1685) | (w3134 & ~w1685);
assign w4358 = w1156 & ~w1046;
assign w4359 = (w1249 & ~pi17) | (w1249 & w4198) | (~pi17 & w4198);
assign w4360 = (~w3524 & ~w3525) | (~w3524 & ~w2181) | (~w3525 & ~w2181);
assign w4361 = w1070 & ~w2181;
assign w4362 = w3746 & ~w146;
assign w4363 = (pi13 & w3604) | (pi13 & ~w146) | (w3604 & ~w146);
assign w4364 = (w3435 & w3434) | (w3435 & ~w2774) | (w3434 & ~w2774);
assign w4365 = (w275 & ~w2722) | (w275 & ~w234) | (~w2722 & ~w234);
assign w4366 = (~w944 & w1127) | (~w944 & w4311) | (w1127 & w4311);
assign w4367 = (~w4022 & ~w4023) | (~w4022 & ~w572) | (~w4023 & ~w572);
assign w4368 = w574 & w2919;
assign w4369 = (~pi01 & ~w3420) | (~pi01 & ~w146) | (~w3420 & ~w146);
assign w4370 = (~pi01 & w4367) | (~pi01 & ~w602) | (w4367 & ~w602);
assign w4371 = w1071 & ~w966;
assign w4372 = (~w32 & w3763) | (~w32 & ~w330) | (w3763 & ~w330);
assign w4373 = (~w783 & w3466) | (~w783 & ~w927) | (w3466 & ~w927);
assign one = 1;
assign po00 = ~w1941;// level 99
assign po01 = ~w1944;// level 101
assign po02 = w1738;// level 90
assign po03 = ~w1951;// level 101
assign po04 = ~w1541;// level 81
assign po05 = w1958;// level 101
assign po06 = w1305;// level 73
assign po07 = ~w1966;// level 101
assign po08 = w1136;// level 64
assign po09 = w1981;// level 101
assign po10 = ~w890;// level 57
assign po11 = ~w2002;// level 102
assign po12 = w2003;// level 50
assign po13 = ~w2016;// level 101
assign po14 = ~w613;// level 42
assign po15 = w2028;// level 101
assign po16 = ~w441;// level 35
assign po17 = w2044;// level 102
assign po18 = ~w341;// level 29
assign po19 = w2051;// level 101
assign po20 = w243;// level 22
assign po21 = ~w2060;// level 101
assign po22 = ~w166;// level 16
assign po23 = ~w2066;// level 101
assign po24 = ~w102;// level 11
assign po25 = ~w2072;// level 102
assign po26 = w2074;// level 7
assign po27 = w2084;// level 101
assign po28 = w2088;// level 6
assign po29 = w2099;// level 102
assign po30 = w2103;// level 6
assign po31 = w2105;// level 100
endmodule
