// Benchmark "aes_core" written by ABC on Wed Apr 29 13:45:51 2015

module aes_core ( 
    pi000, pi001, pi002, pi003, pi004, pi005, pi006, pi007, pi008, pi009,
    pi010, pi011, pi012, pi013, pi014, pi015, pi016, pi017, pi018, pi019,
    pi020, pi021, pi022, pi023, pi024, pi025, pi026, pi027, pi028, pi029,
    pi030, pi031, pi032, pi033, pi034, pi035, pi036, pi037, pi038, pi039,
    pi040, pi041, pi042, pi043, pi044, pi045, pi046, pi047, pi048, pi049,
    pi050, pi051, pi052, pi053, pi054, pi055, pi056, pi057, pi058, pi059,
    pi060, pi061, pi062, pi063, pi064, pi065, pi066, pi067, pi068, pi069,
    pi070, pi071, pi072, pi073, pi074, pi075, pi076, pi077, pi078, pi079,
    pi080, pi081, pi082, pi083, pi084, pi085, pi086, pi087, pi088, pi089,
    pi090, pi091, pi092, pi093, pi094, pi095, pi096, pi097, pi098, pi099,
    pi100, pi101, pi102, pi103, pi104, pi105, pi106, pi107, pi108, pi109,
    pi110, pi111, pi112, pi113, pi114, pi115, pi116, pi117, pi118, pi119,
    pi120, pi121, pi122, pi123, pi124, pi125, pi126, pi127, pi128, pi129,
    pi130, pi131, pi132, pi133, pi134, pi135, pi136, pi137, pi138, pi139,
    pi140, pi141, pi142, pi143, pi144, pi145, pi146, pi147, pi148, pi149,
    pi150, pi151, pi152, pi153, pi154, pi155, pi156, pi157, pi158, pi159,
    pi160, pi161, pi162, pi163, pi164, pi165, pi166, pi167, pi168, pi169,
    pi170, pi171, pi172, pi173, pi174, pi175, pi176, pi177, pi178, pi179,
    pi180, pi181, pi182, pi183, pi184, pi185, pi186, pi187, pi188, pi189,
    pi190, pi191, pi192, pi193, pi194, pi195, pi196, pi197, pi198, pi199,
    pi200, pi201, pi202, pi203, pi204, pi205, pi206, pi207, pi208, pi209,
    pi210, pi211, pi212, pi213, pi214, pi215, pi216, pi217, pi218, pi219,
    pi220, pi221, pi222, pi223, pi224, pi225, pi226, pi227, pi228, pi229,
    pi230, pi231, pi232, pi233, pi234, pi235, pi236, pi237, pi238, pi239,
    pi240, pi241, pi242, pi243, pi244, pi245, pi246, pi247, pi248, pi249,
    pi250, pi251, pi252, pi253, pi254, pi255, pi256, pi257, pi258, pi259,
    pi260, pi261, pi262, pi263, pi264, pi265, pi266, pi267, pi268, pi269,
    pi270, pi271, pi272, pi273, pi274, pi275, pi276, pi277, pi278, pi279,
    pi280, pi281, pi282, pi283, pi284, pi285, pi286, pi287, pi288, pi289,
    pi290, pi291, pi292, pi293, pi294, pi295, pi296, pi297, pi298, pi299,
    pi300, pi301, pi302, pi303, pi304, pi305, pi306, pi307, pi308, pi309,
    pi310, pi311, pi312, pi313, pi314, pi315, pi316, pi317, pi318, pi319,
    pi320, pi321, pi322, pi323, pi324, pi325, pi326, pi327, pi328, pi329,
    pi330, pi331, pi332, pi333, pi334, pi335, pi336, pi337, pi338, pi339,
    pi340, pi341, pi342, pi343, pi344, pi345, pi346, pi347, pi348, pi349,
    pi350, pi351, pi352, pi353, pi354, pi355, pi356, pi357, pi358, pi359,
    pi360, pi361, pi362, pi363, pi364, pi365, pi366, pi367, pi368, pi369,
    pi370, pi371, pi372, pi373, pi374, pi375, pi376, pi377, pi378, pi379,
    pi380, pi381, pi382, pi383, pi384, pi385, pi386, pi387, pi388, pi389,
    pi390, pi391, pi392, pi393, pi394, pi395, pi396, pi397, pi398, pi399,
    pi400, pi401, pi402, pi403, pi404, pi405, pi406, pi407, pi408, pi409,
    pi410, pi411, pi412, pi413, pi414, pi415, pi416, pi417, pi418, pi419,
    pi420, pi421, pi422, pi423, pi424, pi425, pi426, pi427, pi428, pi429,
    pi430, pi431, pi432, pi433, pi434, pi435, pi436, pi437, pi438, pi439,
    pi440, pi441, pi442, pi443, pi444, pi445, pi446, pi447, pi448, pi449,
    pi450, pi451, pi452, pi453, pi454, pi455, pi456, pi457, pi458, pi459,
    pi460, pi461, pi462, pi463, pi464, pi465, pi466, pi467, pi468, pi469,
    pi470, pi471, pi472, pi473, pi474, pi475, pi476, pi477, pi478, pi479,
    pi480, pi481, pi482, pi483, pi484, pi485, pi486, pi487, pi488, pi489,
    pi490, pi491, pi492, pi493, pi494, pi495, pi496, pi497, pi498, pi499,
    pi500, pi501, pi502, pi503, pi504, pi505, pi506, pi507, pi508, pi509,
    pi510, pi511, pi512, pi513, pi514, pi515, pi516, pi517, pi518, pi519,
    pi520, pi521, pi522, pi523, pi524, pi525, pi526, pi527, pi528, pi529,
    pi530, pi531, pi532, pi533, pi534, pi535, pi536, pi537, pi538, pi539,
    pi540, pi541, pi542, pi543, pi544, pi545, pi546, pi547, pi548, pi549,
    pi550, pi551, pi552, pi553, pi554, pi555, pi556, pi557, pi558, pi559,
    pi560, pi561, pi562, pi563, pi564, pi565, pi566, pi567, pi568, pi569,
    pi570, pi571, pi572, pi573, pi574, pi575, pi576, pi577, pi578, pi579,
    pi580, pi581, pi582, pi583, pi584, pi585, pi586, pi587, pi588, pi589,
    pi590, pi591, pi592, pi593, pi594, pi595, pi596, pi597, pi598, pi599,
    pi600, pi601, pi602, pi603, pi604, pi605, pi606, pi607, pi608, pi609,
    pi610, pi611, pi612, pi613, pi614, pi615, pi616, pi617, pi618, pi619,
    pi620, pi621, pi622, pi623, pi624, pi625, pi626, pi627, pi628, pi629,
    pi630, pi631, pi632, pi633, pi634, pi635, pi636, pi637, pi638, pi639,
    pi640, pi641, pi642, pi643, pi644, pi645, pi646, pi647, pi648, pi649,
    pi650, pi651, pi652, pi653, pi654, pi655, pi656, pi657, pi658, pi659,
    pi660, pi661, pi662, pi663, pi664, pi665, pi666, pi667, pi668, pi669,
    pi670, pi671, pi672, pi673, pi674, pi675, pi676, pi677, pi678, pi679,
    pi680, pi681, pi682, pi683, pi684, pi685, pi686, pi687, pi688, pi689,
    pi690, pi691, pi692, pi693, pi694, pi695, pi696, pi697, pi698, pi699,
    pi700, pi701, pi702, pi703, pi704, pi705, pi706, pi707, pi708, pi709,
    pi710, pi711, pi712, pi713, pi714, pi715, pi716, pi717, pi718, pi719,
    pi720, pi721, pi722, pi723, pi724, pi725, pi726, pi727, pi728, pi729,
    pi730, pi731, pi732, pi733, pi734, pi735, pi736, pi737, pi738, pi739,
    pi740, pi741, pi742, pi743, pi744, pi745, pi746, pi747, pi748, pi749,
    pi750, pi751, pi752, pi753, pi754, pi755, pi756, pi757, pi758, pi759,
    pi760, pi761, pi762, pi763, pi764, pi765, pi766, pi767, pi768, pi769,
    pi770, pi771, pi772, pi773, pi774, pi775, pi776, pi777, pi778, pi779,
    pi780, pi781, pi782, pi783, pi784, pi785, pi786, pi787, pi788,
    po000, po001, po002, po003, po004, po005, po006, po007, po008, po009,
    po010, po011, po012, po013, po014, po015, po016, po017, po018, po019,
    po020, po021, po022, po023, po024, po025, po026, po027, po028, po029,
    po030, po031, po032, po033, po034, po035, po036, po037, po038, po039,
    po040, po041, po042, po043, po044, po045, po046, po047, po048, po049,
    po050, po051, po052, po053, po054, po055, po056, po057, po058, po059,
    po060, po061, po062, po063, po064, po065, po066, po067, po068, po069,
    po070, po071, po072, po073, po074, po075, po076, po077, po078, po079,
    po080, po081, po082, po083, po084, po085, po086, po087, po088, po089,
    po090, po091, po092, po093, po094, po095, po096, po097, po098, po099,
    po100, po101, po102, po103, po104, po105, po106, po107, po108, po109,
    po110, po111, po112, po113, po114, po115, po116, po117, po118, po119,
    po120, po121, po122, po123, po124, po125, po126, po127, po128, po129,
    po130, po131, po132, po133, po134, po135, po136, po137, po138, po139,
    po140, po141, po142, po143, po144, po145, po146, po147, po148, po149,
    po150, po151, po152, po153, po154, po155, po156, po157, po158, po159,
    po160, po161, po162, po163, po164, po165, po166, po167, po168, po169,
    po170, po171, po172, po173, po174, po175, po176, po177, po178, po179,
    po180, po181, po182, po183, po184, po185, po186, po187, po188, po189,
    po190, po191, po192, po193, po194, po195, po196, po197, po198, po199,
    po200, po201, po202, po203, po204, po205, po206, po207, po208, po209,
    po210, po211, po212, po213, po214, po215, po216, po217, po218, po219,
    po220, po221, po222, po223, po224, po225, po226, po227, po228, po229,
    po230, po231, po232, po233, po234, po235, po236, po237, po238, po239,
    po240, po241, po242, po243, po244, po245, po246, po247, po248, po249,
    po250, po251, po252, po253, po254, po255, po256, po257, po258, po259,
    po260, po261, po262, po263, po264, po265, po266, po267, po268, po269,
    po270, po271, po272, po273, po274, po275, po276, po277, po278, po279,
    po280, po281, po282, po283, po284, po285, po286, po287, po288, po289,
    po290, po291, po292, po293, po294, po295, po296, po297, po298, po299,
    po300, po301, po302, po303, po304, po305, po306, po307, po308, po309,
    po310, po311, po312, po313, po314, po315, po316, po317, po318, po319,
    po320, po321, po322, po323, po324, po325, po326, po327, po328, po329,
    po330, po331, po332, po333, po334, po335, po336, po337, po338, po339,
    po340, po341, po342, po343, po344, po345, po346, po347, po348, po349,
    po350, po351, po352, po353, po354, po355, po356, po357, po358, po359,
    po360, po361, po362, po363, po364, po365, po366, po367, po368, po369,
    po370, po371, po372, po373, po374, po375, po376, po377, po378, po379,
    po380, po381, po382, po383, po384, po385, po386, po387, po388, po389,
    po390, po391, po392, po393, po394, po395, po396, po397, po398, po399,
    po400, po401, po402, po403, po404, po405, po406, po407, po408, po409,
    po410, po411, po412, po413, po414, po415, po416, po417, po418, po419,
    po420, po421, po422, po423, po424, po425, po426, po427, po428, po429,
    po430, po431, po432, po433, po434, po435, po436, po437, po438, po439,
    po440, po441, po442, po443, po444, po445, po446, po447, po448, po449,
    po450, po451, po452, po453, po454, po455, po456, po457, po458, po459,
    po460, po461, po462, po463, po464, po465, po466, po467, po468, po469,
    po470, po471, po472, po473, po474, po475, po476, po477, po478, po479,
    po480, po481, po482, po483, po484, po485, po486, po487, po488, po489,
    po490, po491, po492, po493, po494, po495, po496, po497, po498, po499,
    po500, po501, po502, po503, po504, po505, po506, po507, po508, po509,
    po510, po511, po512, po513, po514, po515, po516, po517, po518, po519,
    po520, po521, po522, po523, po524, po525, po526, po527, po528, po529,
    po530, po531, po532, po533, po534, po535, po536, po537, po538, po539,
    po540, po541, po542, po543, po544, po545, po546, po547, po548, po549,
    po550, po551, po552, po553, po554, po555, po556, po557, po558, po559,
    po560, po561, po562, po563, po564, po565, po566, po567, po568, po569,
    po570, po571, po572, po573, po574, po575, po576, po577, po578, po579,
    po580, po581, po582, po583, po584, po585, po586, po587, po588, po589,
    po590, po591, po592, po593, po594, po595, po596, po597, po598, po599,
    po600, po601, po602, po603, po604, po605, po606, po607, po608, po609,
    po610, po611, po612, po613, po614, po615, po616, po617, po618, po619,
    po620, po621, po622, po623, po624, po625, po626, po627, po628, po629,
    po630, po631, po632, po633, po634, po635, po636, po637, po638, po639,
    po640, po641, po642, po643, po644, po645, po646, po647, po648, po649,
    po650, po651, po652, po653, po654, po655, po656, po657, po658, po659,
    po660, po661, po662, po663, po664, po665, po666, po667  );
  input  pi000, pi001, pi002, pi003, pi004, pi005, pi006, pi007, pi008,
    pi009, pi010, pi011, pi012, pi013, pi014, pi015, pi016, pi017, pi018,
    pi019, pi020, pi021, pi022, pi023, pi024, pi025, pi026, pi027, pi028,
    pi029, pi030, pi031, pi032, pi033, pi034, pi035, pi036, pi037, pi038,
    pi039, pi040, pi041, pi042, pi043, pi044, pi045, pi046, pi047, pi048,
    pi049, pi050, pi051, pi052, pi053, pi054, pi055, pi056, pi057, pi058,
    pi059, pi060, pi061, pi062, pi063, pi064, pi065, pi066, pi067, pi068,
    pi069, pi070, pi071, pi072, pi073, pi074, pi075, pi076, pi077, pi078,
    pi079, pi080, pi081, pi082, pi083, pi084, pi085, pi086, pi087, pi088,
    pi089, pi090, pi091, pi092, pi093, pi094, pi095, pi096, pi097, pi098,
    pi099, pi100, pi101, pi102, pi103, pi104, pi105, pi106, pi107, pi108,
    pi109, pi110, pi111, pi112, pi113, pi114, pi115, pi116, pi117, pi118,
    pi119, pi120, pi121, pi122, pi123, pi124, pi125, pi126, pi127, pi128,
    pi129, pi130, pi131, pi132, pi133, pi134, pi135, pi136, pi137, pi138,
    pi139, pi140, pi141, pi142, pi143, pi144, pi145, pi146, pi147, pi148,
    pi149, pi150, pi151, pi152, pi153, pi154, pi155, pi156, pi157, pi158,
    pi159, pi160, pi161, pi162, pi163, pi164, pi165, pi166, pi167, pi168,
    pi169, pi170, pi171, pi172, pi173, pi174, pi175, pi176, pi177, pi178,
    pi179, pi180, pi181, pi182, pi183, pi184, pi185, pi186, pi187, pi188,
    pi189, pi190, pi191, pi192, pi193, pi194, pi195, pi196, pi197, pi198,
    pi199, pi200, pi201, pi202, pi203, pi204, pi205, pi206, pi207, pi208,
    pi209, pi210, pi211, pi212, pi213, pi214, pi215, pi216, pi217, pi218,
    pi219, pi220, pi221, pi222, pi223, pi224, pi225, pi226, pi227, pi228,
    pi229, pi230, pi231, pi232, pi233, pi234, pi235, pi236, pi237, pi238,
    pi239, pi240, pi241, pi242, pi243, pi244, pi245, pi246, pi247, pi248,
    pi249, pi250, pi251, pi252, pi253, pi254, pi255, pi256, pi257, pi258,
    pi259, pi260, pi261, pi262, pi263, pi264, pi265, pi266, pi267, pi268,
    pi269, pi270, pi271, pi272, pi273, pi274, pi275, pi276, pi277, pi278,
    pi279, pi280, pi281, pi282, pi283, pi284, pi285, pi286, pi287, pi288,
    pi289, pi290, pi291, pi292, pi293, pi294, pi295, pi296, pi297, pi298,
    pi299, pi300, pi301, pi302, pi303, pi304, pi305, pi306, pi307, pi308,
    pi309, pi310, pi311, pi312, pi313, pi314, pi315, pi316, pi317, pi318,
    pi319, pi320, pi321, pi322, pi323, pi324, pi325, pi326, pi327, pi328,
    pi329, pi330, pi331, pi332, pi333, pi334, pi335, pi336, pi337, pi338,
    pi339, pi340, pi341, pi342, pi343, pi344, pi345, pi346, pi347, pi348,
    pi349, pi350, pi351, pi352, pi353, pi354, pi355, pi356, pi357, pi358,
    pi359, pi360, pi361, pi362, pi363, pi364, pi365, pi366, pi367, pi368,
    pi369, pi370, pi371, pi372, pi373, pi374, pi375, pi376, pi377, pi378,
    pi379, pi380, pi381, pi382, pi383, pi384, pi385, pi386, pi387, pi388,
    pi389, pi390, pi391, pi392, pi393, pi394, pi395, pi396, pi397, pi398,
    pi399, pi400, pi401, pi402, pi403, pi404, pi405, pi406, pi407, pi408,
    pi409, pi410, pi411, pi412, pi413, pi414, pi415, pi416, pi417, pi418,
    pi419, pi420, pi421, pi422, pi423, pi424, pi425, pi426, pi427, pi428,
    pi429, pi430, pi431, pi432, pi433, pi434, pi435, pi436, pi437, pi438,
    pi439, pi440, pi441, pi442, pi443, pi444, pi445, pi446, pi447, pi448,
    pi449, pi450, pi451, pi452, pi453, pi454, pi455, pi456, pi457, pi458,
    pi459, pi460, pi461, pi462, pi463, pi464, pi465, pi466, pi467, pi468,
    pi469, pi470, pi471, pi472, pi473, pi474, pi475, pi476, pi477, pi478,
    pi479, pi480, pi481, pi482, pi483, pi484, pi485, pi486, pi487, pi488,
    pi489, pi490, pi491, pi492, pi493, pi494, pi495, pi496, pi497, pi498,
    pi499, pi500, pi501, pi502, pi503, pi504, pi505, pi506, pi507, pi508,
    pi509, pi510, pi511, pi512, pi513, pi514, pi515, pi516, pi517, pi518,
    pi519, pi520, pi521, pi522, pi523, pi524, pi525, pi526, pi527, pi528,
    pi529, pi530, pi531, pi532, pi533, pi534, pi535, pi536, pi537, pi538,
    pi539, pi540, pi541, pi542, pi543, pi544, pi545, pi546, pi547, pi548,
    pi549, pi550, pi551, pi552, pi553, pi554, pi555, pi556, pi557, pi558,
    pi559, pi560, pi561, pi562, pi563, pi564, pi565, pi566, pi567, pi568,
    pi569, pi570, pi571, pi572, pi573, pi574, pi575, pi576, pi577, pi578,
    pi579, pi580, pi581, pi582, pi583, pi584, pi585, pi586, pi587, pi588,
    pi589, pi590, pi591, pi592, pi593, pi594, pi595, pi596, pi597, pi598,
    pi599, pi600, pi601, pi602, pi603, pi604, pi605, pi606, pi607, pi608,
    pi609, pi610, pi611, pi612, pi613, pi614, pi615, pi616, pi617, pi618,
    pi619, pi620, pi621, pi622, pi623, pi624, pi625, pi626, pi627, pi628,
    pi629, pi630, pi631, pi632, pi633, pi634, pi635, pi636, pi637, pi638,
    pi639, pi640, pi641, pi642, pi643, pi644, pi645, pi646, pi647, pi648,
    pi649, pi650, pi651, pi652, pi653, pi654, pi655, pi656, pi657, pi658,
    pi659, pi660, pi661, pi662, pi663, pi664, pi665, pi666, pi667, pi668,
    pi669, pi670, pi671, pi672, pi673, pi674, pi675, pi676, pi677, pi678,
    pi679, pi680, pi681, pi682, pi683, pi684, pi685, pi686, pi687, pi688,
    pi689, pi690, pi691, pi692, pi693, pi694, pi695, pi696, pi697, pi698,
    pi699, pi700, pi701, pi702, pi703, pi704, pi705, pi706, pi707, pi708,
    pi709, pi710, pi711, pi712, pi713, pi714, pi715, pi716, pi717, pi718,
    pi719, pi720, pi721, pi722, pi723, pi724, pi725, pi726, pi727, pi728,
    pi729, pi730, pi731, pi732, pi733, pi734, pi735, pi736, pi737, pi738,
    pi739, pi740, pi741, pi742, pi743, pi744, pi745, pi746, pi747, pi748,
    pi749, pi750, pi751, pi752, pi753, pi754, pi755, pi756, pi757, pi758,
    pi759, pi760, pi761, pi762, pi763, pi764, pi765, pi766, pi767, pi768,
    pi769, pi770, pi771, pi772, pi773, pi774, pi775, pi776, pi777, pi778,
    pi779, pi780, pi781, pi782, pi783, pi784, pi785, pi786, pi787, pi788;
  output po000, po001, po002, po003, po004, po005, po006, po007, po008, po009,
    po010, po011, po012, po013, po014, po015, po016, po017, po018, po019,
    po020, po021, po022, po023, po024, po025, po026, po027, po028, po029,
    po030, po031, po032, po033, po034, po035, po036, po037, po038, po039,
    po040, po041, po042, po043, po044, po045, po046, po047, po048, po049,
    po050, po051, po052, po053, po054, po055, po056, po057, po058, po059,
    po060, po061, po062, po063, po064, po065, po066, po067, po068, po069,
    po070, po071, po072, po073, po074, po075, po076, po077, po078, po079,
    po080, po081, po082, po083, po084, po085, po086, po087, po088, po089,
    po090, po091, po092, po093, po094, po095, po096, po097, po098, po099,
    po100, po101, po102, po103, po104, po105, po106, po107, po108, po109,
    po110, po111, po112, po113, po114, po115, po116, po117, po118, po119,
    po120, po121, po122, po123, po124, po125, po126, po127, po128, po129,
    po130, po131, po132, po133, po134, po135, po136, po137, po138, po139,
    po140, po141, po142, po143, po144, po145, po146, po147, po148, po149,
    po150, po151, po152, po153, po154, po155, po156, po157, po158, po159,
    po160, po161, po162, po163, po164, po165, po166, po167, po168, po169,
    po170, po171, po172, po173, po174, po175, po176, po177, po178, po179,
    po180, po181, po182, po183, po184, po185, po186, po187, po188, po189,
    po190, po191, po192, po193, po194, po195, po196, po197, po198, po199,
    po200, po201, po202, po203, po204, po205, po206, po207, po208, po209,
    po210, po211, po212, po213, po214, po215, po216, po217, po218, po219,
    po220, po221, po222, po223, po224, po225, po226, po227, po228, po229,
    po230, po231, po232, po233, po234, po235, po236, po237, po238, po239,
    po240, po241, po242, po243, po244, po245, po246, po247, po248, po249,
    po250, po251, po252, po253, po254, po255, po256, po257, po258, po259,
    po260, po261, po262, po263, po264, po265, po266, po267, po268, po269,
    po270, po271, po272, po273, po274, po275, po276, po277, po278, po279,
    po280, po281, po282, po283, po284, po285, po286, po287, po288, po289,
    po290, po291, po292, po293, po294, po295, po296, po297, po298, po299,
    po300, po301, po302, po303, po304, po305, po306, po307, po308, po309,
    po310, po311, po312, po313, po314, po315, po316, po317, po318, po319,
    po320, po321, po322, po323, po324, po325, po326, po327, po328, po329,
    po330, po331, po332, po333, po334, po335, po336, po337, po338, po339,
    po340, po341, po342, po343, po344, po345, po346, po347, po348, po349,
    po350, po351, po352, po353, po354, po355, po356, po357, po358, po359,
    po360, po361, po362, po363, po364, po365, po366, po367, po368, po369,
    po370, po371, po372, po373, po374, po375, po376, po377, po378, po379,
    po380, po381, po382, po383, po384, po385, po386, po387, po388, po389,
    po390, po391, po392, po393, po394, po395, po396, po397, po398, po399,
    po400, po401, po402, po403, po404, po405, po406, po407, po408, po409,
    po410, po411, po412, po413, po414, po415, po416, po417, po418, po419,
    po420, po421, po422, po423, po424, po425, po426, po427, po428, po429,
    po430, po431, po432, po433, po434, po435, po436, po437, po438, po439,
    po440, po441, po442, po443, po444, po445, po446, po447, po448, po449,
    po450, po451, po452, po453, po454, po455, po456, po457, po458, po459,
    po460, po461, po462, po463, po464, po465, po466, po467, po468, po469,
    po470, po471, po472, po473, po474, po475, po476, po477, po478, po479,
    po480, po481, po482, po483, po484, po485, po486, po487, po488, po489,
    po490, po491, po492, po493, po494, po495, po496, po497, po498, po499,
    po500, po501, po502, po503, po504, po505, po506, po507, po508, po509,
    po510, po511, po512, po513, po514, po515, po516, po517, po518, po519,
    po520, po521, po522, po523, po524, po525, po526, po527, po528, po529,
    po530, po531, po532, po533, po534, po535, po536, po537, po538, po539,
    po540, po541, po542, po543, po544, po545, po546, po547, po548, po549,
    po550, po551, po552, po553, po554, po555, po556, po557, po558, po559,
    po560, po561, po562, po563, po564, po565, po566, po567, po568, po569,
    po570, po571, po572, po573, po574, po575, po576, po577, po578, po579,
    po580, po581, po582, po583, po584, po585, po586, po587, po588, po589,
    po590, po591, po592, po593, po594, po595, po596, po597, po598, po599,
    po600, po601, po602, po603, po604, po605, po606, po607, po608, po609,
    po610, po611, po612, po613, po614, po615, po616, po617, po618, po619,
    po620, po621, po622, po623, po624, po625, po626, po627, po628, po629,
    po630, po631, po632, po633, po634, po635, po636, po637, po638, po639,
    po640, po641, po642, po643, po644, po645, po646, po647, po648, po649,
    po650, po651, po652, po653, po654, po655, po656, po657, po658, po659,
    po660, po661, po662, po663, po664, po665, po666, po667;
  wire n1459, n1460, n1461, n1462, n1463, n1464, n1465, n1466, n1467, n1468,
    n1469, n1470, n1471, n1472, n1473, n1474, n1475, n1476, n1477, n1478,
    n1479, n1480, n1481, n1482, n1483, n1484, n1485, n1486, n1487, n1488,
    n1489, n1490, n1491, n1492, n1493, n1494, n1495, n1496, n1497, n1498,
    n1499, n1500, n1501, n1502, n1503, n1504, n1505, n1506, n1507, n1508,
    n1509, n1510, n1511, n1512, n1513, n1514, n1515, n1516, n1517, n1518,
    n1519, n1520, n1521, n1522, n1523, n1524, n1525, n1526, n1527, n1528,
    n1529, n1530, n1531, n1532, n1533, n1534, n1535, n1536, n1537, n1538,
    n1539, n1540, n1541, n1542, n1543, n1544, n1545, n1546, n1547, n1548,
    n1549, n1550, n1551, n1552, n1553, n1554, n1555, n1556, n1557, n1558,
    n1559, n1560, n1561, n1562, n1563, n1564, n1565, n1566, n1567, n1568,
    n1569, n1570, n1571, n1572, n1573, n1574, n1575, n1576, n1577, n1578,
    n1579, n1580, n1581, n1582, n1583, n1584, n1585, n1586, n1587, n1588,
    n1589, n1590, n1591, n1592, n1593, n1594, n1595, n1596, n1597, n1598,
    n1599, n1600, n1601, n1602, n1603, n1604, n1605, n1606, n1607, n1608,
    n1609, n1610, n1611, n1612, n1613, n1614, n1615, n1616, n1617, n1618,
    n1619, n1620, n1621, n1622, n1623, n1624, n1625, n1626, n1627, n1628,
    n1629, n1630, n1631, n1632, n1633, n1634, n1635, n1636, n1637, n1638,
    n1639, n1640, n1641, n1642, n1643, n1644, n1645, n1646, n1647, n1648,
    n1649, n1650, n1651, n1652, n1653, n1654, n1655, n1656, n1657, n1658,
    n1659, n1660, n1661, n1662, n1663, n1664, n1665, n1666, n1667, n1668,
    n1669, n1670, n1671, n1672, n1673, n1674, n1675, n1676, n1677, n1678,
    n1679, n1680, n1681, n1682, n1683, n1684, n1685, n1686, n1687, n1688,
    n1689, n1690, n1691, n1692, n1693, n1694, n1695, n1696, n1697, n1698,
    n1699, n1700, n1701, n1702, n1703, n1704, n1705, n1706, n1707, n1708,
    n1709, n1710, n1711, n1712, n1713, n1714, n1715, n1716, n1717, n1718,
    n1719, n1720, n1721, n1722, n1723, n1724, n1725, n1726, n1727, n1728,
    n1729, n1730, n1731, n1732, n1733, n1734, n1735, n1736, n1737, n1738,
    n1739, n1740, n1741, n1742, n1743, n1744, n1745, n1746, n1747, n1748,
    n1749, n1750, n1751, n1752, n1753, n1754, n1755, n1756, n1757, n1758,
    n1759, n1760, n1761, n1762, n1763, n1764, n1765, n1766, n1767, n1768,
    n1769, n1770, n1771, n1772, n1773, n1774, n1775, n1776, n1777, n1778,
    n1779, n1780, n1781, n1782, n1783, n1784, n1785, n1786, n1787, n1788,
    n1789, n1790, n1791, n1792, n1793, n1794, n1795, n1796, n1797, n1798,
    n1799, n1800, n1801, n1802, n1803, n1804, n1805, n1806, n1807, n1808,
    n1809, n1810, n1811, n1812, n1813, n1814, n1815, n1816, n1817, n1818,
    n1819, n1820, n1821, n1822, n1823, n1824, n1825, n1826, n1827, n1828,
    n1829, n1830, n1831, n1832, n1833, n1834, n1835, n1836, n1837, n1838,
    n1839, n1840, n1841, n1842, n1843, n1844, n1845, n1846, n1847, n1848,
    n1849, n1850, n1851, n1852, n1853, n1854, n1855, n1856, n1857, n1858,
    n1859, n1860, n1861, n1862, n1863, n1864, n1865, n1866, n1867, n1868,
    n1869, n1870, n1871, n1872, n1873, n1874, n1875, n1876, n1877, n1878,
    n1879, n1880, n1881, n1882, n1883, n1884, n1885, n1886, n1887, n1888,
    n1889, n1890, n1891, n1892, n1893, n1894, n1895, n1896, n1897, n1898,
    n1899, n1900, n1901, n1902, n1903, n1904, n1905, n1906, n1907, n1908,
    n1909, n1910, n1911, n1912, n1913, n1914, n1915, n1916, n1917, n1918,
    n1919, n1920, n1921, n1922, n1923, n1924, n1925, n1926, n1927, n1928,
    n1929, n1930, n1931, n1932, n1933, n1934, n1935, n1936, n1937, n1938,
    n1939, n1940, n1941, n1942, n1943, n1944, n1945, n1946, n1947, n1948,
    n1949, n1950, n1951, n1952, n1953, n1954, n1955, n1956, n1957, n1958,
    n1959, n1960, n1961, n1962, n1963, n1964, n1965, n1966, n1967, n1968,
    n1969, n1970, n1971, n1972, n1973, n1974, n1975, n1976, n1977, n1978,
    n1979, n1980, n1981, n1982, n1983, n1984, n1985, n1986, n1987, n1988,
    n1989, n1990, n1991, n1992, n1993, n1994, n1995, n1996, n1997, n1998,
    n1999, n2000, n2001, n2002, n2003, n2004, n2005, n2006, n2007, n2008,
    n2009, n2010, n2011, n2012, n2013, n2014, n2015, n2016, n2017, n2018,
    n2019, n2020, n2021, n2022, n2023, n2024, n2025, n2026, n2027, n2028,
    n2029, n2030, n2031, n2032, n2033, n2034, n2035, n2036, n2037, n2038,
    n2039, n2040, n2041, n2042, n2043, n2044, n2045, n2046, n2047, n2048,
    n2049, n2050, n2051, n2052, n2053, n2054, n2055, n2056, n2057, n2058,
    n2059, n2060, n2061, n2062, n2063, n2064, n2065, n2066, n2067, n2068,
    n2069, n2070, n2071, n2072, n2073, n2074, n2075, n2076, n2077, n2078,
    n2079, n2080, n2081, n2082, n2083, n2084, n2085, n2086, n2087, n2088,
    n2089, n2090, n2091, n2092, n2093, n2094, n2095, n2096, n2097, n2098,
    n2099, n2100, n2101, n2102, n2103, n2104, n2105, n2106, n2107, n2108,
    n2109, n2110, n2111, n2112, n2113, n2114, n2115, n2116, n2117, n2118,
    n2119, n2120, n2121, n2122, n2123, n2124, n2125, n2126, n2127, n2128,
    n2129, n2130, n2131, n2132, n2133, n2134, n2135, n2136, n2137, n2138,
    n2139, n2140, n2141, n2142, n2143, n2144, n2145, n2146, n2147, n2148,
    n2149, n2150, n2151, n2152, n2153, n2154, n2155, n2156, n2157, n2158,
    n2159, n2160, n2161, n2162, n2163, n2164, n2165, n2166, n2167, n2168,
    n2169, n2170, n2171, n2172, n2173, n2174, n2175, n2176, n2177, n2178,
    n2179, n2180, n2181, n2182, n2183, n2184, n2185, n2186, n2187, n2188,
    n2189, n2190, n2191, n2192, n2193, n2194, n2195, n2196, n2197, n2198,
    n2199, n2200, n2201, n2202, n2203, n2204, n2205, n2206, n2207, n2208,
    n2209, n2210, n2211, n2212, n2213, n2214, n2215, n2216, n2217, n2218,
    n2219, n2220, n2221, n2222, n2223, n2224, n2225, n2226, n2227, n2228,
    n2229, n2230, n2231, n2232, n2233, n2234, n2235, n2236, n2237, n2238,
    n2239, n2240, n2241, n2242, n2243, n2244, n2245, n2246, n2247, n2248,
    n2249, n2250, n2251, n2252, n2253, n2254, n2255, n2256, n2257, n2258,
    n2259, n2260, n2261, n2262, n2263, n2264, n2265, n2266, n2267, n2268,
    n2269, n2270, n2271, n2272, n2273, n2274, n2275, n2276, n2277, n2278,
    n2279, n2280, n2281, n2282, n2283, n2284, n2285, n2286, n2287, n2288,
    n2289, n2290, n2291, n2292, n2293, n2294, n2295, n2296, n2297, n2298,
    n2299, n2300, n2301, n2302, n2303, n2304, n2305, n2306, n2307, n2308,
    n2309, n2310, n2311, n2312, n2313, n2314, n2315, n2316, n2317, n2318,
    n2319, n2320, n2321, n2322, n2323, n2324, n2325, n2326, n2327, n2328,
    n2329, n2330, n2331, n2332, n2333, n2334, n2335, n2336, n2337, n2338,
    n2339, n2340, n2341, n2342, n2343, n2344, n2345, n2346, n2347, n2348,
    n2349, n2350, n2351, n2352, n2353, n2354, n2355, n2356, n2357, n2358,
    n2359, n2360, n2361, n2362, n2363, n2364, n2365, n2366, n2367, n2368,
    n2369, n2370, n2371, n2372, n2373, n2374, n2375, n2376, n2377, n2378,
    n2379, n2380, n2381, n2382, n2383, n2384, n2385, n2386, n2387, n2388,
    n2389, n2390, n2391, n2392, n2393, n2394, n2395, n2396, n2397, n2398,
    n2399, n2400, n2401, n2402, n2403, n2404, n2405, n2406, n2407, n2408,
    n2409, n2410, n2411, n2412, n2413, n2414, n2415, n2416, n2417, n2418,
    n2419, n2420, n2421, n2422, n2423, n2424, n2425, n2426, n2427, n2428,
    n2429, n2430, n2431, n2432, n2433, n2434, n2435, n2436, n2437, n2438,
    n2439, n2440, n2441, n2442, n2443, n2444, n2445, n2446, n2447, n2448,
    n2449, n2450, n2451, n2452, n2453, n2454, n2455, n2456, n2457, n2458,
    n2459, n2460, n2461, n2462, n2463, n2464, n2465, n2466, n2467, n2468,
    n2469, n2470, n2471, n2472, n2473, n2474, n2475, n2476, n2477, n2478,
    n2479, n2480, n2481, n2482, n2483, n2484, n2486, n2487, n2488, n2489,
    n2490, n2491, n2492, n2493, n2494, n2495, n2496, n2497, n2498, n2499,
    n2500, n2501, n2502, n2503, n2504, n2505, n2506, n2507, n2508, n2509,
    n2510, n2511, n2512, n2513, n2514, n2515, n2516, n2517, n2518, n2519,
    n2520, n2521, n2522, n2523, n2524, n2525, n2526, n2527, n2528, n2529,
    n2530, n2531, n2532, n2533, n2534, n2535, n2536, n2537, n2538, n2539,
    n2540, n2541, n2542, n2543, n2544, n2545, n2546, n2547, n2548, n2549,
    n2550, n2551, n2552, n2553, n2554, n2555, n2556, n2557, n2558, n2559,
    n2560, n2561, n2562, n2563, n2564, n2565, n2566, n2567, n2568, n2569,
    n2570, n2571, n2572, n2573, n2574, n2575, n2576, n2577, n2578, n2579,
    n2580, n2581, n2582, n2583, n2584, n2585, n2586, n2587, n2588, n2589,
    n2590, n2591, n2592, n2593, n2594, n2595, n2596, n2597, n2598, n2599,
    n2600, n2601, n2602, n2603, n2604, n2605, n2606, n2607, n2608, n2609,
    n2610, n2611, n2612, n2613, n2614, n2615, n2616, n2617, n2618, n2619,
    n2620, n2621, n2622, n2623, n2624, n2625, n2626, n2627, n2628, n2629,
    n2630, n2631, n2632, n2633, n2634, n2635, n2636, n2637, n2638, n2639,
    n2640, n2641, n2642, n2643, n2644, n2645, n2646, n2647, n2648, n2649,
    n2650, n2651, n2652, n2653, n2654, n2655, n2656, n2657, n2658, n2659,
    n2660, n2661, n2662, n2663, n2664, n2665, n2666, n2667, n2668, n2669,
    n2670, n2671, n2672, n2673, n2674, n2675, n2676, n2677, n2678, n2679,
    n2680, n2681, n2682, n2683, n2684, n2685, n2686, n2687, n2688, n2689,
    n2690, n2691, n2692, n2693, n2694, n2695, n2696, n2697, n2698, n2699,
    n2700, n2701, n2702, n2703, n2704, n2705, n2706, n2707, n2708, n2709,
    n2710, n2711, n2712, n2713, n2714, n2715, n2716, n2717, n2718, n2719,
    n2720, n2721, n2722, n2723, n2724, n2725, n2726, n2727, n2728, n2729,
    n2730, n2731, n2732, n2733, n2734, n2735, n2736, n2737, n2738, n2739,
    n2740, n2741, n2742, n2743, n2744, n2745, n2746, n2747, n2748, n2749,
    n2750, n2751, n2752, n2753, n2754, n2755, n2756, n2757, n2758, n2759,
    n2760, n2761, n2762, n2763, n2764, n2765, n2766, n2767, n2768, n2769,
    n2770, n2771, n2772, n2773, n2774, n2775, n2776, n2777, n2778, n2779,
    n2780, n2781, n2782, n2783, n2784, n2785, n2786, n2787, n2788, n2789,
    n2790, n2791, n2792, n2793, n2794, n2795, n2796, n2797, n2798, n2799,
    n2800, n2801, n2802, n2803, n2804, n2805, n2806, n2807, n2808, n2809,
    n2810, n2811, n2812, n2813, n2814, n2815, n2816, n2817, n2818, n2819,
    n2820, n2821, n2822, n2823, n2824, n2825, n2826, n2827, n2828, n2829,
    n2830, n2831, n2832, n2833, n2834, n2835, n2836, n2837, n2838, n2839,
    n2840, n2841, n2842, n2843, n2844, n2845, n2846, n2847, n2848, n2849,
    n2850, n2851, n2852, n2853, n2854, n2855, n2856, n2857, n2858, n2859,
    n2860, n2861, n2862, n2863, n2864, n2865, n2866, n2867, n2868, n2869,
    n2870, n2871, n2872, n2873, n2874, n2875, n2876, n2877, n2878, n2879,
    n2880, n2881, n2882, n2883, n2884, n2885, n2886, n2887, n2888, n2889,
    n2890, n2891, n2892, n2893, n2894, n2895, n2896, n2897, n2898, n2899,
    n2900, n2901, n2902, n2903, n2904, n2905, n2906, n2907, n2908, n2909,
    n2910, n2911, n2912, n2913, n2914, n2915, n2916, n2917, n2918, n2919,
    n2920, n2921, n2922, n2923, n2924, n2925, n2926, n2927, n2928, n2929,
    n2930, n2931, n2932, n2933, n2934, n2935, n2936, n2937, n2938, n2939,
    n2940, n2941, n2942, n2943, n2944, n2945, n2946, n2947, n2948, n2949,
    n2950, n2951, n2952, n2953, n2954, n2955, n2956, n2957, n2958, n2959,
    n2960, n2961, n2962, n2963, n2964, n2965, n2966, n2967, n2968, n2969,
    n2970, n2971, n2972, n2973, n2974, n2975, n2976, n2977, n2978, n2979,
    n2980, n2981, n2982, n2983, n2984, n2985, n2986, n2987, n2988, n2989,
    n2990, n2991, n2992, n2993, n2994, n2995, n2996, n2997, n2998, n2999,
    n3000, n3001, n3002, n3003, n3004, n3005, n3006, n3007, n3008, n3009,
    n3010, n3011, n3012, n3013, n3014, n3015, n3016, n3017, n3018, n3019,
    n3020, n3021, n3022, n3023, n3024, n3025, n3026, n3027, n3028, n3029,
    n3030, n3031, n3032, n3033, n3034, n3035, n3036, n3037, n3038, n3039,
    n3040, n3041, n3042, n3043, n3044, n3045, n3046, n3047, n3048, n3049,
    n3050, n3051, n3052, n3053, n3054, n3055, n3056, n3057, n3058, n3059,
    n3060, n3061, n3062, n3063, n3064, n3065, n3066, n3067, n3068, n3069,
    n3070, n3071, n3072, n3073, n3074, n3075, n3076, n3077, n3078, n3079,
    n3080, n3081, n3082, n3083, n3084, n3085, n3086, n3087, n3088, n3089,
    n3090, n3091, n3092, n3093, n3094, n3095, n3096, n3097, n3098, n3099,
    n3100, n3101, n3102, n3103, n3104, n3105, n3106, n3107, n3108, n3109,
    n3110, n3111, n3112, n3113, n3114, n3115, n3116, n3117, n3118, n3119,
    n3120, n3121, n3122, n3123, n3124, n3125, n3126, n3127, n3128, n3129,
    n3130, n3131, n3132, n3133, n3134, n3135, n3136, n3137, n3138, n3139,
    n3140, n3141, n3142, n3143, n3144, n3145, n3146, n3147, n3148, n3149,
    n3150, n3151, n3152, n3153, n3154, n3155, n3156, n3157, n3158, n3159,
    n3160, n3161, n3162, n3163, n3164, n3165, n3166, n3167, n3168, n3169,
    n3170, n3171, n3172, n3173, n3174, n3175, n3176, n3177, n3178, n3179,
    n3180, n3181, n3182, n3183, n3184, n3185, n3186, n3187, n3188, n3189,
    n3190, n3191, n3192, n3193, n3194, n3195, n3196, n3197, n3198, n3199,
    n3200, n3201, n3202, n3203, n3204, n3205, n3206, n3207, n3208, n3209,
    n3210, n3211, n3212, n3213, n3214, n3215, n3216, n3217, n3218, n3219,
    n3220, n3221, n3222, n3223, n3224, n3225, n3226, n3227, n3228, n3229,
    n3230, n3231, n3232, n3233, n3234, n3235, n3236, n3237, n3238, n3239,
    n3240, n3241, n3242, n3243, n3244, n3245, n3246, n3247, n3248, n3249,
    n3250, n3251, n3253, n3254, n3255, n3256, n3257, n3258, n3259, n3260,
    n3261, n3262, n3263, n3264, n3265, n3266, n3267, n3268, n3269, n3270,
    n3271, n3272, n3273, n3274, n3275, n3276, n3277, n3278, n3279, n3280,
    n3281, n3282, n3283, n3284, n3285, n3286, n3287, n3288, n3289, n3290,
    n3291, n3292, n3293, n3294, n3295, n3296, n3297, n3298, n3299, n3300,
    n3301, n3302, n3303, n3304, n3305, n3306, n3307, n3308, n3309, n3310,
    n3311, n3312, n3313, n3314, n3315, n3316, n3317, n3318, n3319, n3320,
    n3321, n3322, n3323, n3324, n3325, n3326, n3327, n3328, n3329, n3330,
    n3331, n3332, n3333, n3334, n3335, n3336, n3337, n3338, n3339, n3340,
    n3341, n3342, n3343, n3344, n3345, n3346, n3347, n3348, n3349, n3350,
    n3351, n3352, n3353, n3354, n3355, n3356, n3357, n3358, n3359, n3360,
    n3361, n3362, n3363, n3364, n3365, n3366, n3367, n3368, n3369, n3370,
    n3371, n3372, n3373, n3374, n3375, n3376, n3377, n3378, n3379, n3380,
    n3381, n3382, n3383, n3384, n3385, n3386, n3387, n3388, n3389, n3390,
    n3391, n3392, n3393, n3394, n3395, n3396, n3397, n3398, n3399, n3400,
    n3401, n3402, n3403, n3404, n3405, n3406, n3407, n3408, n3409, n3410,
    n3411, n3412, n3413, n3414, n3415, n3416, n3417, n3418, n3419, n3420,
    n3421, n3422, n3423, n3424, n3425, n3426, n3427, n3428, n3429, n3430,
    n3431, n3432, n3433, n3434, n3435, n3436, n3437, n3438, n3439, n3440,
    n3441, n3442, n3443, n3444, n3445, n3446, n3447, n3448, n3449, n3450,
    n3451, n3452, n3453, n3454, n3455, n3456, n3457, n3458, n3459, n3460,
    n3461, n3462, n3463, n3464, n3465, n3466, n3467, n3468, n3469, n3470,
    n3471, n3472, n3473, n3474, n3475, n3476, n3477, n3478, n3479, n3480,
    n3481, n3482, n3483, n3484, n3485, n3486, n3487, n3488, n3489, n3490,
    n3491, n3492, n3493, n3494, n3495, n3496, n3497, n3498, n3499, n3500,
    n3501, n3502, n3503, n3504, n3505, n3506, n3507, n3508, n3509, n3510,
    n3511, n3512, n3513, n3514, n3515, n3516, n3517, n3518, n3519, n3520,
    n3521, n3522, n3523, n3524, n3525, n3526, n3527, n3528, n3529, n3530,
    n3531, n3532, n3533, n3534, n3535, n3536, n3537, n3538, n3539, n3540,
    n3541, n3542, n3543, n3544, n3545, n3546, n3547, n3548, n3549, n3550,
    n3551, n3552, n3553, n3554, n3555, n3556, n3557, n3558, n3559, n3560,
    n3561, n3562, n3563, n3564, n3565, n3566, n3567, n3568, n3569, n3570,
    n3571, n3572, n3573, n3574, n3575, n3576, n3577, n3578, n3579, n3580,
    n3581, n3582, n3583, n3584, n3585, n3586, n3587, n3588, n3589, n3590,
    n3591, n3592, n3593, n3594, n3595, n3596, n3597, n3598, n3599, n3600,
    n3601, n3602, n3603, n3604, n3605, n3606, n3607, n3608, n3609, n3610,
    n3611, n3612, n3613, n3614, n3615, n3616, n3617, n3618, n3619, n3620,
    n3621, n3622, n3623, n3624, n3625, n3626, n3627, n3628, n3629, n3630,
    n3631, n3632, n3633, n3634, n3635, n3636, n3637, n3638, n3639, n3640,
    n3641, n3642, n3643, n3644, n3645, n3646, n3647, n3648, n3649, n3650,
    n3651, n3652, n3653, n3654, n3655, n3656, n3657, n3658, n3659, n3660,
    n3661, n3662, n3663, n3664, n3665, n3666, n3667, n3668, n3669, n3670,
    n3671, n3672, n3673, n3674, n3675, n3676, n3677, n3678, n3679, n3680,
    n3681, n3682, n3683, n3684, n3685, n3686, n3687, n3688, n3689, n3690,
    n3691, n3692, n3693, n3694, n3695, n3696, n3697, n3698, n3699, n3700,
    n3701, n3702, n3703, n3704, n3705, n3706, n3707, n3708, n3709, n3710,
    n3711, n3712, n3713, n3714, n3715, n3716, n3717, n3718, n3719, n3720,
    n3721, n3722, n3723, n3724, n3725, n3726, n3727, n3728, n3729, n3730,
    n3731, n3732, n3733, n3734, n3735, n3736, n3737, n3738, n3739, n3740,
    n3741, n3742, n3743, n3744, n3745, n3746, n3747, n3748, n3749, n3750,
    n3751, n3752, n3753, n3754, n3755, n3756, n3757, n3758, n3759, n3760,
    n3761, n3762, n3763, n3764, n3765, n3766, n3767, n3768, n3769, n3770,
    n3771, n3772, n3773, n3774, n3775, n3776, n3777, n3778, n3779, n3780,
    n3781, n3782, n3783, n3784, n3785, n3786, n3787, n3788, n3789, n3790,
    n3791, n3792, n3793, n3794, n3795, n3796, n3797, n3798, n3799, n3800,
    n3801, n3802, n3803, n3804, n3805, n3806, n3807, n3808, n3809, n3810,
    n3811, n3812, n3813, n3814, n3815, n3816, n3817, n3818, n3819, n3820,
    n3821, n3822, n3823, n3824, n3825, n3826, n3827, n3828, n3829, n3830,
    n3831, n3832, n3833, n3834, n3835, n3836, n3837, n3838, n3839, n3840,
    n3841, n3842, n3843, n3844, n3845, n3846, n3847, n3848, n3849, n3850,
    n3851, n3852, n3853, n3854, n3855, n3856, n3857, n3858, n3859, n3860,
    n3861, n3862, n3863, n3864, n3865, n3866, n3867, n3868, n3869, n3870,
    n3871, n3872, n3873, n3874, n3875, n3876, n3877, n3878, n3879, n3880,
    n3881, n3882, n3883, n3884, n3885, n3886, n3887, n3888, n3889, n3890,
    n3891, n3892, n3893, n3894, n3895, n3896, n3897, n3898, n3899, n3900,
    n3901, n3902, n3903, n3904, n3905, n3906, n3907, n3908, n3909, n3910,
    n3911, n3912, n3913, n3914, n3915, n3916, n3917, n3918, n3919, n3920,
    n3921, n3922, n3923, n3924, n3925, n3926, n3927, n3928, n3929, n3930,
    n3931, n3932, n3933, n3934, n3935, n3936, n3937, n3938, n3939, n3940,
    n3941, n3942, n3943, n3944, n3945, n3946, n3947, n3948, n3949, n3950,
    n3951, n3952, n3953, n3954, n3955, n3956, n3957, n3958, n3959, n3960,
    n3961, n3962, n3963, n3964, n3965, n3966, n3967, n3968, n3969, n3970,
    n3971, n3972, n3973, n3974, n3975, n3976, n3977, n3978, n3979, n3980,
    n3981, n3982, n3983, n3984, n3985, n3986, n3987, n3988, n3989, n3990,
    n3991, n3992, n3993, n3994, n3995, n3996, n3997, n3998, n3999, n4000,
    n4001, n4002, n4003, n4004, n4005, n4006, n4007, n4008, n4009, n4010,
    n4011, n4012, n4013, n4014, n4015, n4016, n4017, n4018, n4019, n4020,
    n4021, n4022, n4023, n4024, n4025, n4026, n4027, n4028, n4029, n4030,
    n4031, n4032, n4033, n4034, n4035, n4036, n4037, n4038, n4039, n4040,
    n4041, n4042, n4043, n4044, n4045, n4046, n4047, n4048, n4049, n4050,
    n4051, n4052, n4053, n4054, n4055, n4056, n4057, n4058, n4059, n4060,
    n4061, n4062, n4063, n4064, n4065, n4066, n4067, n4068, n4069, n4070,
    n4071, n4072, n4073, n4074, n4075, n4076, n4077, n4078, n4079, n4080,
    n4081, n4082, n4083, n4084, n4085, n4086, n4087, n4088, n4089, n4090,
    n4091, n4092, n4093, n4094, n4095, n4096, n4097, n4098, n4099, n4100,
    n4101, n4102, n4103, n4104, n4105, n4106, n4107, n4108, n4109, n4110,
    n4111, n4112, n4113, n4114, n4115, n4116, n4117, n4118, n4119, n4120,
    n4121, n4122, n4123, n4124, n4125, n4126, n4127, n4128, n4129, n4130,
    n4131, n4132, n4133, n4134, n4135, n4136, n4137, n4138, n4139, n4140,
    n4141, n4142, n4143, n4144, n4145, n4146, n4147, n4148, n4149, n4150,
    n4151, n4152, n4153, n4154, n4155, n4156, n4157, n4158, n4159, n4160,
    n4161, n4162, n4163, n4164, n4165, n4166, n4167, n4168, n4169, n4170,
    n4171, n4172, n4173, n4174, n4175, n4176, n4177, n4178, n4179, n4180,
    n4181, n4182, n4183, n4184, n4185, n4186, n4187, n4188, n4189, n4190,
    n4191, n4192, n4193, n4194, n4195, n4196, n4197, n4198, n4199, n4200,
    n4201, n4202, n4203, n4204, n4205, n4206, n4207, n4208, n4209, n4210,
    n4211, n4212, n4213, n4214, n4215, n4216, n4217, n4218, n4219, n4220,
    n4221, n4222, n4223, n4224, n4225, n4226, n4227, n4228, n4229, n4230,
    n4231, n4232, n4233, n4234, n4235, n4236, n4237, n4238, n4239, n4240,
    n4241, n4242, n4243, n4244, n4245, n4246, n4247, n4248, n4249, n4250,
    n4251, n4252, n4253, n4254, n4255, n4256, n4257, n4258, n4259, n4260,
    n4261, n4262, n4263, n4264, n4265, n4266, n4267, n4268, n4269, n4270,
    n4271, n4272, n4273, n4274, n4275, n4276, n4277, n4278, n4279, n4280,
    n4282, n4283, n4284, n4285, n4286, n4287, n4288, n4289, n4290, n4291,
    n4292, n4293, n4294, n4295, n4296, n4297, n4298, n4299, n4300, n4301,
    n4302, n4303, n4304, n4305, n4306, n4307, n4308, n4309, n4310, n4311,
    n4312, n4313, n4314, n4315, n4316, n4317, n4318, n4319, n4320, n4321,
    n4322, n4323, n4324, n4325, n4326, n4327, n4328, n4329, n4330, n4331,
    n4332, n4333, n4334, n4335, n4336, n4337, n4338, n4339, n4340, n4341,
    n4342, n4343, n4344, n4345, n4346, n4347, n4348, n4349, n4350, n4351,
    n4352, n4353, n4354, n4355, n4356, n4357, n4358, n4359, n4360, n4361,
    n4362, n4363, n4364, n4365, n4366, n4367, n4368, n4369, n4370, n4371,
    n4372, n4373, n4374, n4375, n4376, n4377, n4378, n4379, n4380, n4381,
    n4382, n4383, n4384, n4385, n4386, n4387, n4388, n4389, n4390, n4391,
    n4392, n4393, n4394, n4395, n4396, n4397, n4398, n4399, n4400, n4401,
    n4402, n4403, n4404, n4405, n4406, n4407, n4408, n4409, n4410, n4411,
    n4412, n4413, n4414, n4415, n4416, n4417, n4418, n4419, n4420, n4421,
    n4422, n4423, n4424, n4425, n4426, n4427, n4428, n4429, n4430, n4431,
    n4432, n4433, n4434, n4435, n4436, n4437, n4438, n4439, n4440, n4441,
    n4442, n4443, n4444, n4445, n4446, n4447, n4448, n4449, n4450, n4451,
    n4452, n4453, n4454, n4455, n4456, n4457, n4458, n4459, n4460, n4461,
    n4462, n4463, n4464, n4465, n4466, n4467, n4468, n4469, n4470, n4471,
    n4472, n4473, n4474, n4475, n4476, n4477, n4478, n4479, n4480, n4481,
    n4482, n4483, n4484, n4485, n4486, n4487, n4488, n4489, n4490, n4491,
    n4492, n4493, n4494, n4495, n4496, n4497, n4498, n4499, n4500, n4501,
    n4502, n4503, n4504, n4505, n4506, n4507, n4508, n4509, n4510, n4511,
    n4512, n4513, n4514, n4515, n4516, n4517, n4518, n4519, n4520, n4521,
    n4522, n4523, n4524, n4525, n4526, n4527, n4528, n4529, n4530, n4531,
    n4532, n4533, n4534, n4535, n4536, n4537, n4538, n4539, n4540, n4541,
    n4542, n4543, n4544, n4545, n4546, n4547, n4548, n4549, n4550, n4551,
    n4552, n4553, n4554, n4555, n4556, n4557, n4558, n4559, n4560, n4561,
    n4562, n4563, n4564, n4565, n4566, n4567, n4568, n4569, n4570, n4571,
    n4572, n4573, n4574, n4575, n4576, n4577, n4578, n4579, n4580, n4581,
    n4582, n4583, n4584, n4585, n4586, n4587, n4588, n4589, n4590, n4591,
    n4592, n4593, n4594, n4595, n4596, n4597, n4598, n4599, n4600, n4601,
    n4602, n4603, n4604, n4605, n4606, n4607, n4608, n4609, n4610, n4611,
    n4612, n4613, n4614, n4615, n4616, n4617, n4618, n4619, n4620, n4621,
    n4622, n4623, n4624, n4625, n4626, n4627, n4628, n4629, n4630, n4631,
    n4632, n4633, n4634, n4635, n4636, n4637, n4638, n4639, n4640, n4641,
    n4642, n4643, n4644, n4645, n4646, n4647, n4648, n4649, n4650, n4651,
    n4652, n4653, n4654, n4655, n4656, n4657, n4658, n4659, n4660, n4661,
    n4662, n4663, n4664, n4665, n4666, n4667, n4668, n4669, n4670, n4671,
    n4672, n4673, n4674, n4675, n4676, n4677, n4678, n4679, n4680, n4681,
    n4682, n4683, n4684, n4685, n4686, n4687, n4688, n4689, n4690, n4691,
    n4692, n4693, n4694, n4695, n4696, n4697, n4698, n4699, n4700, n4701,
    n4702, n4703, n4704, n4705, n4706, n4707, n4708, n4709, n4710, n4711,
    n4712, n4713, n4714, n4715, n4716, n4717, n4718, n4719, n4720, n4721,
    n4722, n4723, n4724, n4725, n4726, n4727, n4728, n4729, n4730, n4731,
    n4732, n4733, n4734, n4735, n4736, n4737, n4738, n4739, n4740, n4741,
    n4742, n4743, n4744, n4745, n4746, n4747, n4748, n4749, n4750, n4751,
    n4752, n4753, n4754, n4755, n4756, n4757, n4758, n4759, n4760, n4761,
    n4762, n4763, n4764, n4765, n4766, n4767, n4768, n4769, n4770, n4771,
    n4772, n4773, n4774, n4775, n4776, n4777, n4778, n4779, n4780, n4781,
    n4782, n4783, n4784, n4785, n4786, n4787, n4788, n4789, n4790, n4791,
    n4792, n4793, n4794, n4795, n4796, n4797, n4798, n4799, n4800, n4801,
    n4802, n4803, n4804, n4805, n4806, n4807, n4808, n4809, n4810, n4811,
    n4812, n4813, n4814, n4815, n4816, n4817, n4818, n4819, n4820, n4821,
    n4822, n4823, n4824, n4825, n4826, n4827, n4828, n4829, n4830, n4831,
    n4832, n4833, n4834, n4835, n4836, n4837, n4838, n4839, n4840, n4841,
    n4842, n4843, n4844, n4845, n4846, n4847, n4848, n4849, n4850, n4851,
    n4852, n4853, n4854, n4855, n4856, n4857, n4858, n4859, n4860, n4861,
    n4862, n4863, n4864, n4865, n4866, n4867, n4868, n4869, n4870, n4871,
    n4872, n4873, n4874, n4875, n4876, n4877, n4878, n4879, n4880, n4881,
    n4882, n4883, n4884, n4885, n4886, n4887, n4888, n4889, n4890, n4891,
    n4892, n4893, n4894, n4895, n4896, n4897, n4898, n4899, n4900, n4901,
    n4902, n4903, n4904, n4905, n4906, n4907, n4908, n4909, n4910, n4911,
    n4912, n4913, n4914, n4915, n4916, n4917, n4918, n4919, n4920, n4921,
    n4922, n4923, n4924, n4925, n4926, n4927, n4928, n4929, n4930, n4931,
    n4932, n4933, n4934, n4935, n4936, n4937, n4938, n4939, n4940, n4941,
    n4942, n4943, n4944, n4945, n4946, n4947, n4948, n4949, n4950, n4951,
    n4952, n4953, n4954, n4955, n4956, n4957, n4958, n4959, n4960, n4961,
    n4962, n4963, n4964, n4965, n4966, n4967, n4968, n4969, n4970, n4971,
    n4972, n4973, n4974, n4975, n4976, n4977, n4978, n4979, n4980, n4981,
    n4982, n4983, n4984, n4985, n4986, n4987, n4988, n4989, n4990, n4991,
    n4992, n4993, n4994, n4995, n4996, n4997, n4998, n4999, n5000, n5001,
    n5002, n5003, n5004, n5005, n5006, n5007, n5008, n5009, n5010, n5011,
    n5012, n5013, n5014, n5015, n5016, n5017, n5018, n5019, n5020, n5021,
    n5022, n5023, n5024, n5025, n5026, n5027, n5028, n5029, n5030, n5031,
    n5032, n5033, n5034, n5035, n5036, n5037, n5038, n5039, n5040, n5041,
    n5042, n5043, n5044, n5045, n5046, n5047, n5048, n5049, n5050, n5051,
    n5052, n5053, n5054, n5055, n5056, n5057, n5058, n5059, n5060, n5061,
    n5062, n5063, n5064, n5065, n5066, n5067, n5068, n5069, n5070, n5071,
    n5072, n5073, n5074, n5075, n5076, n5077, n5078, n5079, n5080, n5081,
    n5082, n5083, n5084, n5085, n5086, n5087, n5088, n5089, n5090, n5091,
    n5092, n5093, n5094, n5095, n5096, n5097, n5098, n5099, n5100, n5101,
    n5102, n5103, n5104, n5105, n5106, n5107, n5108, n5109, n5110, n5111,
    n5112, n5113, n5114, n5115, n5116, n5117, n5118, n5119, n5120, n5121,
    n5122, n5123, n5124, n5125, n5126, n5127, n5128, n5129, n5130, n5131,
    n5132, n5133, n5134, n5135, n5136, n5137, n5138, n5139, n5140, n5141,
    n5142, n5143, n5144, n5145, n5146, n5147, n5148, n5149, n5150, n5151,
    n5152, n5153, n5154, n5155, n5156, n5157, n5158, n5159, n5160, n5161,
    n5162, n5163, n5164, n5165, n5166, n5167, n5168, n5169, n5170, n5171,
    n5172, n5173, n5174, n5175, n5176, n5177, n5178, n5179, n5180, n5181,
    n5182, n5183, n5184, n5185, n5186, n5187, n5188, n5189, n5190, n5191,
    n5192, n5193, n5194, n5195, n5196, n5197, n5198, n5199, n5200, n5201,
    n5202, n5203, n5204, n5205, n5206, n5207, n5208, n5209, n5210, n5211,
    n5212, n5213, n5214, n5215, n5216, n5217, n5218, n5219, n5220, n5221,
    n5222, n5223, n5224, n5225, n5226, n5227, n5228, n5229, n5230, n5231,
    n5232, n5233, n5234, n5235, n5236, n5237, n5238, n5239, n5240, n5241,
    n5242, n5243, n5244, n5245, n5246, n5247, n5248, n5249, n5250, n5251,
    n5252, n5253, n5254, n5255, n5256, n5257, n5258, n5259, n5260, n5261,
    n5262, n5263, n5264, n5265, n5266, n5267, n5268, n5269, n5270, n5271,
    n5272, n5273, n5274, n5275, n5276, n5277, n5278, n5279, n5280, n5281,
    n5282, n5283, n5284, n5285, n5286, n5287, n5288, n5289, n5290, n5291,
    n5292, n5293, n5294, n5295, n5296, n5297, n5298, n5299, n5300, n5301,
    n5302, n5303, n5304, n5305, n5306, n5307, n5308, n5309, n5310, n5311,
    n5313, n5314, n5315, n5316, n5317, n5318, n5319, n5320, n5321, n5322,
    n5323, n5324, n5325, n5326, n5327, n5328, n5329, n5330, n5331, n5332,
    n5333, n5334, n5335, n5336, n5337, n5338, n5339, n5340, n5341, n5342,
    n5343, n5344, n5345, n5346, n5347, n5348, n5349, n5350, n5351, n5352,
    n5353, n5354, n5355, n5356, n5357, n5358, n5359, n5360, n5361, n5362,
    n5363, n5364, n5365, n5366, n5367, n5368, n5369, n5370, n5371, n5372,
    n5373, n5374, n5375, n5376, n5377, n5378, n5379, n5380, n5381, n5382,
    n5383, n5384, n5385, n5386, n5387, n5388, n5389, n5390, n5391, n5392,
    n5393, n5394, n5395, n5396, n5397, n5398, n5399, n5400, n5401, n5402,
    n5403, n5404, n5405, n5406, n5407, n5408, n5409, n5410, n5411, n5412,
    n5413, n5414, n5415, n5416, n5417, n5418, n5419, n5420, n5421, n5422,
    n5423, n5424, n5425, n5426, n5427, n5428, n5429, n5430, n5431, n5432,
    n5433, n5434, n5435, n5436, n5437, n5438, n5439, n5440, n5441, n5442,
    n5443, n5444, n5445, n5446, n5447, n5448, n5449, n5450, n5451, n5452,
    n5453, n5454, n5455, n5456, n5457, n5458, n5459, n5460, n5461, n5462,
    n5463, n5464, n5465, n5466, n5467, n5468, n5469, n5470, n5471, n5472,
    n5473, n5474, n5475, n5476, n5477, n5478, n5479, n5480, n5481, n5482,
    n5483, n5484, n5485, n5486, n5487, n5488, n5489, n5490, n5491, n5492,
    n5493, n5494, n5495, n5496, n5497, n5498, n5499, n5500, n5501, n5502,
    n5503, n5504, n5505, n5506, n5507, n5508, n5509, n5510, n5511, n5512,
    n5513, n5514, n5515, n5516, n5517, n5518, n5519, n5520, n5521, n5522,
    n5523, n5524, n5525, n5526, n5527, n5528, n5529, n5530, n5531, n5532,
    n5533, n5534, n5535, n5536, n5537, n5538, n5539, n5540, n5541, n5542,
    n5543, n5544, n5545, n5546, n5547, n5548, n5549, n5550, n5551, n5552,
    n5553, n5554, n5555, n5556, n5557, n5558, n5559, n5560, n5561, n5562,
    n5563, n5564, n5565, n5566, n5567, n5568, n5569, n5570, n5571, n5572,
    n5573, n5574, n5575, n5576, n5577, n5578, n5579, n5580, n5581, n5582,
    n5583, n5584, n5585, n5586, n5587, n5588, n5589, n5590, n5591, n5592,
    n5593, n5594, n5595, n5596, n5597, n5598, n5599, n5600, n5601, n5602,
    n5603, n5604, n5605, n5606, n5607, n5608, n5609, n5610, n5611, n5612,
    n5613, n5614, n5615, n5616, n5617, n5618, n5619, n5620, n5621, n5622,
    n5623, n5624, n5625, n5626, n5627, n5628, n5629, n5630, n5631, n5632,
    n5633, n5634, n5635, n5636, n5637, n5638, n5639, n5640, n5641, n5642,
    n5643, n5644, n5645, n5646, n5647, n5648, n5649, n5650, n5651, n5652,
    n5653, n5654, n5655, n5656, n5657, n5658, n5659, n5660, n5661, n5662,
    n5663, n5664, n5665, n5666, n5667, n5668, n5669, n5670, n5671, n5672,
    n5673, n5674, n5675, n5676, n5677, n5678, n5679, n5680, n5681, n5682,
    n5683, n5684, n5685, n5686, n5687, n5688, n5689, n5690, n5691, n5692,
    n5693, n5694, n5695, n5696, n5697, n5698, n5699, n5700, n5701, n5702,
    n5703, n5704, n5705, n5706, n5707, n5708, n5709, n5710, n5711, n5712,
    n5713, n5714, n5715, n5716, n5717, n5718, n5719, n5720, n5721, n5722,
    n5723, n5724, n5725, n5726, n5727, n5728, n5729, n5730, n5731, n5732,
    n5733, n5734, n5735, n5736, n5737, n5738, n5739, n5740, n5741, n5742,
    n5743, n5744, n5745, n5746, n5747, n5748, n5749, n5750, n5751, n5752,
    n5753, n5754, n5755, n5756, n5757, n5758, n5759, n5760, n5761, n5762,
    n5763, n5764, n5765, n5766, n5767, n5768, n5769, n5770, n5771, n5772,
    n5773, n5774, n5775, n5776, n5777, n5778, n5779, n5780, n5781, n5782,
    n5783, n5784, n5785, n5786, n5787, n5788, n5789, n5790, n5791, n5792,
    n5793, n5794, n5795, n5796, n5797, n5798, n5799, n5800, n5801, n5802,
    n5803, n5804, n5805, n5806, n5807, n5808, n5809, n5810, n5811, n5812,
    n5813, n5814, n5815, n5816, n5817, n5818, n5819, n5820, n5821, n5822,
    n5823, n5824, n5825, n5826, n5827, n5828, n5829, n5830, n5831, n5832,
    n5833, n5834, n5835, n5836, n5837, n5838, n5839, n5840, n5841, n5842,
    n5843, n5844, n5845, n5846, n5847, n5848, n5849, n5850, n5851, n5852,
    n5853, n5854, n5855, n5856, n5857, n5858, n5859, n5860, n5861, n5862,
    n5863, n5864, n5865, n5866, n5867, n5868, n5869, n5870, n5871, n5872,
    n5873, n5874, n5875, n5876, n5877, n5878, n5879, n5880, n5881, n5882,
    n5883, n5884, n5885, n5886, n5887, n5888, n5889, n5890, n5891, n5892,
    n5893, n5894, n5895, n5896, n5897, n5898, n5899, n5900, n5901, n5902,
    n5903, n5904, n5905, n5906, n5907, n5908, n5909, n5910, n5911, n5912,
    n5913, n5914, n5915, n5916, n5917, n5918, n5919, n5920, n5921, n5922,
    n5923, n5924, n5925, n5926, n5927, n5928, n5929, n5930, n5931, n5932,
    n5933, n5934, n5935, n5936, n5937, n5938, n5939, n5940, n5941, n5942,
    n5943, n5944, n5945, n5946, n5947, n5948, n5949, n5950, n5951, n5952,
    n5953, n5954, n5955, n5956, n5957, n5958, n5959, n5960, n5961, n5962,
    n5963, n5964, n5965, n5966, n5967, n5968, n5969, n5970, n5971, n5972,
    n5973, n5974, n5975, n5976, n5977, n5978, n5979, n5980, n5981, n5982,
    n5983, n5984, n5985, n5986, n5987, n5988, n5989, n5990, n5991, n5992,
    n5993, n5994, n5995, n5996, n5997, n5998, n5999, n6000, n6001, n6002,
    n6003, n6004, n6005, n6006, n6007, n6008, n6009, n6010, n6011, n6012,
    n6013, n6014, n6015, n6016, n6017, n6018, n6019, n6020, n6021, n6022,
    n6023, n6024, n6025, n6026, n6027, n6028, n6029, n6030, n6031, n6032,
    n6033, n6034, n6035, n6036, n6037, n6038, n6039, n6040, n6041, n6042,
    n6043, n6044, n6045, n6046, n6047, n6048, n6049, n6050, n6051, n6052,
    n6053, n6054, n6055, n6056, n6057, n6058, n6059, n6060, n6061, n6062,
    n6063, n6064, n6065, n6066, n6067, n6068, n6069, n6070, n6071, n6072,
    n6073, n6074, n6075, n6076, n6077, n6078, n6079, n6080, n6081, n6082,
    n6083, n6084, n6085, n6086, n6087, n6088, n6089, n6090, n6091, n6092,
    n6093, n6094, n6095, n6096, n6097, n6098, n6099, n6100, n6101, n6102,
    n6103, n6104, n6105, n6106, n6107, n6108, n6109, n6110, n6111, n6112,
    n6113, n6114, n6115, n6116, n6117, n6118, n6119, n6120, n6121, n6122,
    n6123, n6124, n6125, n6126, n6127, n6128, n6129, n6130, n6131, n6132,
    n6133, n6134, n6135, n6136, n6137, n6138, n6139, n6140, n6141, n6142,
    n6143, n6144, n6145, n6146, n6147, n6148, n6149, n6150, n6151, n6152,
    n6153, n6154, n6155, n6156, n6157, n6158, n6159, n6160, n6161, n6162,
    n6163, n6164, n6165, n6166, n6167, n6168, n6169, n6170, n6171, n6172,
    n6173, n6174, n6175, n6176, n6177, n6178, n6179, n6180, n6181, n6182,
    n6183, n6184, n6185, n6186, n6187, n6188, n6189, n6190, n6191, n6192,
    n6193, n6194, n6195, n6196, n6197, n6198, n6199, n6200, n6201, n6202,
    n6203, n6204, n6205, n6206, n6207, n6208, n6209, n6210, n6211, n6212,
    n6213, n6214, n6215, n6216, n6217, n6218, n6219, n6220, n6221, n6222,
    n6223, n6224, n6225, n6226, n6227, n6228, n6229, n6230, n6231, n6232,
    n6233, n6234, n6235, n6236, n6237, n6238, n6239, n6240, n6241, n6242,
    n6243, n6244, n6245, n6246, n6247, n6248, n6249, n6250, n6251, n6252,
    n6253, n6254, n6255, n6256, n6257, n6258, n6259, n6260, n6261, n6262,
    n6263, n6264, n6265, n6266, n6267, n6268, n6269, n6270, n6271, n6272,
    n6273, n6274, n6275, n6276, n6277, n6278, n6279, n6280, n6281, n6282,
    n6283, n6284, n6285, n6286, n6287, n6288, n6289, n6290, n6291, n6292,
    n6293, n6294, n6295, n6296, n6297, n6298, n6299, n6300, n6301, n6302,
    n6303, n6304, n6305, n6306, n6307, n6308, n6309, n6310, n6311, n6312,
    n6313, n6314, n6315, n6316, n6317, n6318, n6319, n6320, n6321, n6322,
    n6323, n6324, n6325, n6326, n6327, n6328, n6329, n6330, n6331, n6332,
    n6333, n6334, n6335, n6336, n6337, n6338, n6340, n6341, n6342, n6343,
    n6344, n6345, n6346, n6347, n6348, n6349, n6350, n6351, n6352, n6353,
    n6354, n6355, n6356, n6357, n6358, n6359, n6360, n6361, n6362, n6363,
    n6364, n6365, n6366, n6367, n6368, n6369, n6370, n6371, n6372, n6373,
    n6374, n6375, n6376, n6377, n6378, n6379, n6380, n6381, n6382, n6383,
    n6384, n6385, n6386, n6387, n6388, n6389, n6390, n6391, n6392, n6393,
    n6394, n6395, n6396, n6397, n6398, n6399, n6400, n6401, n6402, n6403,
    n6404, n6405, n6406, n6407, n6408, n6409, n6410, n6411, n6412, n6413,
    n6414, n6415, n6416, n6417, n6418, n6419, n6420, n6421, n6422, n6423,
    n6424, n6425, n6426, n6427, n6428, n6429, n6430, n6431, n6432, n6433,
    n6434, n6435, n6436, n6437, n6438, n6439, n6440, n6441, n6442, n6443,
    n6444, n6445, n6446, n6447, n6448, n6449, n6450, n6451, n6452, n6453,
    n6454, n6455, n6456, n6457, n6458, n6459, n6460, n6461, n6462, n6463,
    n6464, n6465, n6466, n6467, n6468, n6469, n6470, n6471, n6472, n6473,
    n6474, n6475, n6476, n6477, n6478, n6479, n6480, n6481, n6482, n6483,
    n6484, n6485, n6486, n6487, n6488, n6489, n6490, n6491, n6492, n6493,
    n6494, n6495, n6496, n6497, n6498, n6499, n6500, n6501, n6502, n6503,
    n6504, n6505, n6506, n6507, n6508, n6509, n6510, n6511, n6512, n6513,
    n6514, n6515, n6516, n6517, n6518, n6519, n6520, n6521, n6522, n6523,
    n6524, n6525, n6526, n6527, n6528, n6529, n6530, n6531, n6532, n6533,
    n6534, n6535, n6536, n6537, n6538, n6539, n6540, n6541, n6542, n6543,
    n6544, n6545, n6546, n6547, n6548, n6549, n6550, n6551, n6552, n6553,
    n6554, n6555, n6556, n6557, n6558, n6559, n6560, n6561, n6562, n6563,
    n6564, n6565, n6566, n6567, n6568, n6569, n6570, n6571, n6572, n6573,
    n6574, n6575, n6576, n6577, n6578, n6579, n6580, n6581, n6582, n6583,
    n6584, n6585, n6586, n6587, n6588, n6589, n6590, n6591, n6592, n6593,
    n6594, n6595, n6596, n6597, n6598, n6599, n6600, n6601, n6602, n6603,
    n6604, n6605, n6606, n6607, n6608, n6609, n6610, n6611, n6612, n6613,
    n6614, n6615, n6616, n6617, n6618, n6619, n6620, n6621, n6622, n6623,
    n6624, n6625, n6626, n6627, n6628, n6629, n6630, n6631, n6632, n6633,
    n6634, n6635, n6636, n6637, n6638, n6639, n6640, n6641, n6642, n6643,
    n6644, n6645, n6646, n6647, n6648, n6649, n6650, n6651, n6652, n6653,
    n6654, n6655, n6656, n6657, n6658, n6659, n6660, n6661, n6662, n6663,
    n6664, n6665, n6666, n6667, n6668, n6669, n6670, n6671, n6672, n6673,
    n6674, n6675, n6676, n6677, n6678, n6679, n6680, n6681, n6682, n6683,
    n6684, n6685, n6686, n6687, n6688, n6689, n6690, n6691, n6692, n6693,
    n6694, n6695, n6696, n6697, n6698, n6699, n6700, n6701, n6702, n6703,
    n6704, n6705, n6706, n6707, n6708, n6709, n6710, n6711, n6712, n6713,
    n6714, n6715, n6716, n6717, n6718, n6719, n6720, n6721, n6722, n6723,
    n6724, n6725, n6726, n6727, n6728, n6729, n6730, n6731, n6732, n6733,
    n6734, n6735, n6736, n6737, n6738, n6739, n6740, n6741, n6742, n6743,
    n6744, n6745, n6746, n6747, n6748, n6749, n6750, n6751, n6752, n6753,
    n6754, n6755, n6756, n6757, n6758, n6759, n6760, n6761, n6762, n6763,
    n6764, n6765, n6766, n6767, n6768, n6769, n6770, n6771, n6772, n6773,
    n6774, n6775, n6776, n6777, n6778, n6779, n6780, n6781, n6782, n6783,
    n6784, n6785, n6786, n6787, n6788, n6789, n6790, n6791, n6792, n6793,
    n6795, n6796, n6797, n6798, n6799, n6800, n6801, n6802, n6803, n6804,
    n6805, n6806, n6807, n6808, n6809, n6810, n6811, n6812, n6813, n6814,
    n6815, n6816, n6817, n6818, n6819, n6820, n6821, n6822, n6823, n6824,
    n6825, n6826, n6827, n6828, n6829, n6830, n6831, n6832, n6833, n6834,
    n6835, n6836, n6837, n6838, n6839, n6840, n6841, n6842, n6843, n6844,
    n6845, n6846, n6847, n6848, n6849, n6850, n6851, n6852, n6853, n6854,
    n6855, n6856, n6857, n6858, n6859, n6860, n6861, n6862, n6863, n6864,
    n6865, n6866, n6867, n6868, n6869, n6870, n6871, n6872, n6873, n6874,
    n6875, n6876, n6877, n6878, n6879, n6880, n6881, n6882, n6883, n6884,
    n6885, n6886, n6887, n6888, n6889, n6890, n6891, n6892, n6893, n6894,
    n6895, n6896, n6897, n6898, n6899, n6900, n6901, n6902, n6903, n6904,
    n6905, n6906, n6907, n6908, n6909, n6910, n6911, n6912, n6913, n6914,
    n6915, n6916, n6917, n6918, n6919, n6920, n6921, n6922, n6923, n6924,
    n6925, n6926, n6927, n6928, n6929, n6930, n6931, n6932, n6933, n6934,
    n6935, n6936, n6937, n6938, n6939, n6940, n6941, n6942, n6943, n6944,
    n6945, n6946, n6947, n6948, n6949, n6950, n6951, n6952, n6953, n6954,
    n6955, n6956, n6957, n6958, n6959, n6960, n6961, n6962, n6963, n6964,
    n6965, n6966, n6967, n6968, n6969, n6970, n6971, n6972, n6973, n6974,
    n6975, n6976, n6977, n6978, n6979, n6980, n6981, n6982, n6983, n6984,
    n6985, n6986, n6987, n6988, n6989, n6990, n6991, n6992, n6993, n6994,
    n6995, n6996, n6997, n6998, n6999, n7000, n7001, n7002, n7003, n7004,
    n7005, n7006, n7007, n7008, n7009, n7010, n7011, n7012, n7013, n7014,
    n7015, n7016, n7017, n7018, n7019, n7020, n7021, n7022, n7023, n7024,
    n7025, n7026, n7027, n7028, n7029, n7030, n7031, n7032, n7033, n7034,
    n7035, n7036, n7037, n7038, n7039, n7040, n7041, n7042, n7043, n7044,
    n7045, n7046, n7047, n7048, n7049, n7050, n7051, n7052, n7053, n7054,
    n7055, n7056, n7057, n7058, n7059, n7060, n7061, n7062, n7063, n7064,
    n7065, n7066, n7067, n7068, n7069, n7070, n7071, n7072, n7073, n7074,
    n7075, n7076, n7077, n7078, n7079, n7080, n7081, n7082, n7083, n7084,
    n7085, n7086, n7087, n7088, n7089, n7090, n7091, n7092, n7093, n7094,
    n7095, n7096, n7097, n7098, n7099, n7100, n7101, n7102, n7103, n7104,
    n7105, n7106, n7107, n7108, n7109, n7110, n7111, n7112, n7113, n7114,
    n7115, n7116, n7117, n7118, n7119, n7120, n7121, n7122, n7123, n7124,
    n7125, n7126, n7127, n7128, n7129, n7130, n7131, n7132, n7133, n7134,
    n7135, n7136, n7137, n7138, n7139, n7140, n7141, n7142, n7143, n7144,
    n7145, n7146, n7147, n7148, n7149, n7150, n7151, n7152, n7153, n7154,
    n7155, n7156, n7157, n7158, n7159, n7160, n7161, n7162, n7163, n7164,
    n7165, n7166, n7167, n7168, n7169, n7170, n7171, n7172, n7173, n7174,
    n7175, n7176, n7177, n7178, n7179, n7180, n7181, n7182, n7183, n7184,
    n7185, n7186, n7187, n7188, n7189, n7190, n7191, n7192, n7193, n7194,
    n7195, n7196, n7197, n7198, n7199, n7200, n7201, n7202, n7203, n7204,
    n7205, n7207, n7208, n7209, n7210, n7211, n7212, n7213, n7214, n7215,
    n7216, n7217, n7218, n7219, n7220, n7221, n7222, n7223, n7224, n7225,
    n7226, n7227, n7228, n7229, n7230, n7231, n7232, n7233, n7234, n7235,
    n7236, n7237, n7238, n7239, n7240, n7241, n7242, n7243, n7244, n7245,
    n7246, n7247, n7248, n7249, n7250, n7251, n7252, n7253, n7254, n7255,
    n7256, n7257, n7258, n7259, n7260, n7261, n7262, n7263, n7264, n7265,
    n7266, n7267, n7268, n7269, n7270, n7271, n7272, n7273, n7274, n7275,
    n7276, n7277, n7278, n7279, n7280, n7281, n7282, n7283, n7284, n7285,
    n7286, n7287, n7288, n7289, n7290, n7291, n7292, n7293, n7294, n7295,
    n7296, n7297, n7298, n7299, n7300, n7301, n7302, n7303, n7304, n7305,
    n7306, n7307, n7308, n7309, n7310, n7311, n7312, n7313, n7314, n7315,
    n7316, n7317, n7318, n7319, n7320, n7321, n7322, n7323, n7324, n7325,
    n7326, n7327, n7328, n7329, n7330, n7331, n7332, n7333, n7334, n7335,
    n7336, n7337, n7338, n7339, n7340, n7341, n7342, n7343, n7344, n7345,
    n7346, n7347, n7348, n7349, n7350, n7351, n7352, n7353, n7354, n7355,
    n7356, n7357, n7358, n7359, n7360, n7361, n7362, n7363, n7364, n7365,
    n7366, n7367, n7368, n7369, n7370, n7371, n7372, n7373, n7374, n7375,
    n7376, n7377, n7378, n7379, n7380, n7381, n7382, n7383, n7384, n7385,
    n7386, n7387, n7388, n7389, n7390, n7391, n7392, n7393, n7394, n7395,
    n7396, n7397, n7398, n7399, n7400, n7401, n7402, n7403, n7404, n7405,
    n7406, n7407, n7408, n7409, n7410, n7411, n7412, n7413, n7414, n7415,
    n7416, n7417, n7418, n7419, n7420, n7421, n7422, n7423, n7424, n7425,
    n7426, n7427, n7428, n7429, n7430, n7431, n7432, n7433, n7434, n7435,
    n7436, n7437, n7438, n7439, n7440, n7441, n7442, n7443, n7444, n7445,
    n7446, n7447, n7448, n7449, n7450, n7451, n7452, n7453, n7454, n7455,
    n7456, n7457, n7458, n7459, n7460, n7461, n7462, n7463, n7464, n7465,
    n7466, n7467, n7468, n7469, n7470, n7471, n7472, n7473, n7474, n7475,
    n7476, n7477, n7478, n7479, n7480, n7481, n7482, n7483, n7484, n7485,
    n7486, n7487, n7488, n7489, n7490, n7491, n7492, n7493, n7494, n7495,
    n7496, n7497, n7498, n7499, n7500, n7501, n7502, n7503, n7504, n7505,
    n7506, n7507, n7508, n7509, n7510, n7511, n7512, n7513, n7514, n7516,
    n7517, n7518, n7519, n7520, n7521, n7522, n7523, n7524, n7525, n7526,
    n7527, n7528, n7529, n7530, n7531, n7532, n7533, n7534, n7535, n7536,
    n7537, n7538, n7539, n7540, n7541, n7542, n7543, n7544, n7545, n7546,
    n7547, n7548, n7549, n7550, n7551, n7552, n7553, n7554, n7555, n7556,
    n7557, n7558, n7559, n7560, n7561, n7562, n7563, n7564, n7565, n7566,
    n7567, n7568, n7569, n7570, n7571, n7572, n7573, n7574, n7575, n7576,
    n7577, n7578, n7579, n7580, n7581, n7582, n7583, n7584, n7585, n7586,
    n7587, n7588, n7589, n7590, n7591, n7592, n7593, n7594, n7595, n7596,
    n7597, n7598, n7599, n7600, n7601, n7602, n7603, n7604, n7605, n7606,
    n7607, n7608, n7609, n7610, n7611, n7612, n7613, n7614, n7615, n7616,
    n7617, n7618, n7619, n7620, n7621, n7622, n7623, n7624, n7625, n7626,
    n7627, n7628, n7629, n7630, n7631, n7632, n7633, n7634, n7635, n7636,
    n7637, n7638, n7639, n7640, n7641, n7642, n7643, n7644, n7645, n7646,
    n7647, n7648, n7649, n7650, n7651, n7652, n7653, n7654, n7655, n7656,
    n7657, n7658, n7659, n7660, n7661, n7662, n7663, n7664, n7665, n7666,
    n7667, n7668, n7669, n7670, n7671, n7672, n7673, n7674, n7675, n7676,
    n7677, n7678, n7679, n7680, n7681, n7682, n7683, n7684, n7685, n7686,
    n7687, n7688, n7689, n7690, n7691, n7692, n7693, n7694, n7695, n7696,
    n7697, n7698, n7699, n7700, n7701, n7702, n7703, n7704, n7705, n7706,
    n7707, n7709, n7710, n7711, n7712, n7713, n7714, n7715, n7716, n7717,
    n7718, n7719, n7720, n7721, n7722, n7723, n7724, n7725, n7726, n7727,
    n7728, n7729, n7730, n7731, n7732, n7733, n7734, n7735, n7736, n7737,
    n7738, n7739, n7740, n7741, n7742, n7743, n7744, n7745, n7746, n7747,
    n7748, n7749, n7750, n7751, n7752, n7753, n7754, n7755, n7756, n7757,
    n7758, n7759, n7760, n7761, n7762, n7763, n7764, n7765, n7766, n7767,
    n7768, n7769, n7770, n7771, n7772, n7773, n7774, n7775, n7776, n7777,
    n7778, n7779, n7780, n7781, n7782, n7783, n7784, n7785, n7786, n7787,
    n7788, n7789, n7790, n7791, n7792, n7793, n7794, n7795, n7796, n7797,
    n7798, n7799, n7800, n7801, n7802, n7803, n7804, n7805, n7806, n7807,
    n7808, n7809, n7810, n7811, n7812, n7813, n7814, n7815, n7816, n7817,
    n7818, n7819, n7820, n7821, n7822, n7823, n7824, n7825, n7826, n7827,
    n7828, n7829, n7830, n7831, n7832, n7833, n7834, n7835, n7836, n7837,
    n7838, n7839, n7840, n7841, n7842, n7843, n7844, n7845, n7846, n7847,
    n7848, n7849, n7850, n7851, n7852, n7853, n7854, n7855, n7856, n7857,
    n7858, n7859, n7860, n7861, n7862, n7863, n7864, n7865, n7866, n7867,
    n7868, n7869, n7870, n7871, n7872, n7873, n7874, n7875, n7876, n7877,
    n7878, n7879, n7880, n7881, n7882, n7883, n7884, n7885, n7886, n7887,
    n7888, n7889, n7890, n7891, n7892, n7893, n7894, n7895, n7896, n7897,
    n7898, n7899, n7900, n7901, n7903, n7904, n7905, n7906, n7907, n7908,
    n7909, n7910, n7911, n7912, n7913, n7914, n7915, n7916, n7917, n7918,
    n7919, n7920, n7921, n7922, n7923, n7924, n7925, n7926, n7927, n7928,
    n7929, n7930, n7931, n7932, n7933, n7934, n7935, n7936, n7937, n7938,
    n7939, n7940, n7941, n7942, n7943, n7944, n7945, n7946, n7947, n7948,
    n7949, n7950, n7951, n7952, n7953, n7954, n7955, n7956, n7957, n7958,
    n7959, n7960, n7961, n7962, n7963, n7964, n7965, n7966, n7967, n7968,
    n7969, n7970, n7971, n7972, n7973, n7974, n7975, n7976, n7977, n7978,
    n7979, n7980, n7981, n7982, n7983, n7984, n7985, n7986, n7987, n7988,
    n7989, n7990, n7991, n7992, n7993, n7994, n7995, n7996, n7998, n7999,
    n8001, n8002, n8003, n8004, n8005, n8006, n8007, n8008, n8009, n8010,
    n8011, n8012, n8013, n8014, n8015, n8016, n8017, n8018, n8019, n8020,
    n8021, n8022, n8023, n8025, n8026, n8027, n8028, n8029, n8030, n8031,
    n8032, n8033, n8034, n8035, n8036, n8037, n8038, n8039, n8040, n8041,
    n8042, n8043, n8044, n8045, n8046, n8047, n8048, n8049, n8050, n8051,
    n8052, n8053, n8054, n8055, n8056, n8057, n8058, n8059, n8060, n8061,
    n8062, n8063, n8064, n8065, n8066, n8067, n8068, n8069, n8070, n8071,
    n8072, n8073, n8074, n8075, n8076, n8077, n8078, n8079, n8080, n8081,
    n8082, n8083, n8084, n8085, n8086, n8087, n8088, n8089, n8090, n8091,
    n8092, n8093, n8094, n8095, n8096, n8097, n8098, n8099, n8100, n8101,
    n8102, n8103, n8104, n8105, n8106, n8107, n8108, n8109, n8110, n8111,
    n8112, n8113, n8114, n8115, n8116, n8117, n8118, n8119, n8120, n8121,
    n8122, n8123, n8124, n8125, n8126, n8127, n8128, n8129, n8130, n8131,
    n8132, n8133, n8134, n8135, n8136, n8137, n8138, n8139, n8140, n8141,
    n8142, n8143, n8144, n8145, n8146, n8147, n8148, n8149, n8150, n8151,
    n8152, n8153, n8154, n8155, n8156, n8157, n8158, n8159, n8160, n8161,
    n8162, n8163, n8164, n8165, n8166, n8167, n8168, n8169, n8170, n8171,
    n8172, n8173, n8174, n8175, n8176, n8177, n8178, n8179, n8180, n8181,
    n8182, n8183, n8184, n8185, n8186, n8187, n8188, n8189, n8190, n8191,
    n8192, n8193, n8194, n8195, n8196, n8197, n8198, n8199, n8200, n8201,
    n8202, n8203, n8204, n8205, n8206, n8207, n8208, n8209, n8210, n8211,
    n8212, n8213, n8214, n8215, n8216, n8217, n8218, n8219, n8220, n8221,
    n8222, n8223, n8224, n8225, n8226, n8227, n8228, n8229, n8230, n8231,
    n8232, n8233, n8234, n8235, n8236, n8237, n8238, n8239, n8240, n8241,
    n8242, n8243, n8244, n8245, n8246, n8247, n8248, n8249, n8250, n8251,
    n8252, n8253, n8254, n8255, n8256, n8257, n8258, n8259, n8260, n8261,
    n8262, n8263, n8264, n8265, n8266, n8267, n8268, n8269, n8270, n8271,
    n8273, n8274, n8276, n8277, n8278, n8279, n8280, n8281, n8282, n8283,
    n8284, n8285, n8286, n8287, n8288, n8289, n8290, n8291, n8292, n8293,
    n8294, n8295, n8296, n8297, n8298, n8300, n8301, n8302, n8303, n8304,
    n8305, n8306, n8307, n8308, n8309, n8310, n8311, n8312, n8313, n8314,
    n8315, n8316, n8317, n8318, n8319, n8320, n8321, n8322, n8323, n8324,
    n8325, n8326, n8327, n8328, n8329, n8330, n8331, n8332, n8333, n8334,
    n8335, n8336, n8337, n8338, n8339, n8340, n8341, n8342, n8343, n8344,
    n8345, n8346, n8347, n8348, n8349, n8350, n8351, n8352, n8353, n8354,
    n8355, n8356, n8357, n8358, n8359, n8360, n8361, n8362, n8363, n8364,
    n8365, n8366, n8367, n8368, n8369, n8370, n8371, n8372, n8373, n8374,
    n8375, n8376, n8377, n8378, n8379, n8380, n8381, n8382, n8383, n8384,
    n8385, n8386, n8387, n8388, n8389, n8390, n8391, n8392, n8393, n8394,
    n8395, n8396, n8397, n8398, n8399, n8400, n8401, n8402, n8403, n8404,
    n8405, n8406, n8407, n8408, n8409, n8410, n8411, n8412, n8413, n8414,
    n8415, n8416, n8417, n8418, n8419, n8420, n8421, n8422, n8423, n8424,
    n8425, n8426, n8427, n8428, n8429, n8430, n8431, n8432, n8433, n8434,
    n8435, n8436, n8437, n8438, n8439, n8440, n8441, n8442, n8443, n8444,
    n8445, n8446, n8447, n8448, n8449, n8450, n8451, n8452, n8453, n8454,
    n8455, n8456, n8457, n8458, n8459, n8460, n8461, n8462, n8463, n8464,
    n8465, n8466, n8467, n8468, n8469, n8470, n8471, n8472, n8473, n8474,
    n8475, n8476, n8477, n8478, n8479, n8480, n8481, n8482, n8483, n8484,
    n8485, n8486, n8487, n8488, n8489, n8490, n8491, n8492, n8493, n8494,
    n8495, n8496, n8497, n8498, n8499, n8500, n8501, n8502, n8503, n8504,
    n8505, n8506, n8507, n8508, n8509, n8510, n8511, n8512, n8513, n8514,
    n8515, n8516, n8517, n8518, n8519, n8520, n8521, n8522, n8523, n8524,
    n8525, n8526, n8527, n8528, n8529, n8530, n8531, n8532, n8533, n8534,
    n8535, n8536, n8537, n8538, n8539, n8540, n8541, n8542, n8543, n8544,
    n8545, n8546, n8547, n8548, n8549, n8550, n8551, n8552, n8553, n8554,
    n8555, n8556, n8557, n8558, n8559, n8560, n8561, n8562, n8563, n8564,
    n8565, n8566, n8567, n8568, n8569, n8570, n8571, n8572, n8573, n8574,
    n8575, n8576, n8577, n8578, n8579, n8580, n8581, n8582, n8583, n8584,
    n8585, n8586, n8587, n8588, n8589, n8590, n8591, n8592, n8593, n8594,
    n8595, n8596, n8597, n8598, n8599, n8600, n8601, n8602, n8603, n8604,
    n8605, n8606, n8607, n8608, n8609, n8610, n8611, n8612, n8613, n8614,
    n8615, n8616, n8617, n8618, n8619, n8620, n8621, n8622, n8623, n8624,
    n8625, n8626, n8627, n8628, n8629, n8630, n8631, n8632, n8633, n8634,
    n8635, n8636, n8637, n8638, n8639, n8640, n8641, n8642, n8643, n8644,
    n8645, n8646, n8647, n8648, n8649, n8650, n8651, n8652, n8653, n8654,
    n8655, n8656, n8657, n8658, n8659, n8660, n8661, n8662, n8663, n8664,
    n8665, n8666, n8667, n8668, n8669, n8670, n8671, n8672, n8673, n8674,
    n8675, n8676, n8677, n8678, n8679, n8680, n8681, n8682, n8683, n8684,
    n8685, n8686, n8687, n8688, n8689, n8690, n8691, n8692, n8693, n8694,
    n8695, n8696, n8697, n8698, n8699, n8700, n8701, n8702, n8703, n8704,
    n8705, n8706, n8707, n8708, n8709, n8710, n8711, n8712, n8713, n8714,
    n8715, n8716, n8717, n8718, n8719, n8720, n8721, n8722, n8723, n8724,
    n8725, n8726, n8727, n8728, n8729, n8730, n8731, n8732, n8733, n8734,
    n8735, n8736, n8737, n8738, n8739, n8740, n8741, n8742, n8743, n8744,
    n8745, n8746, n8747, n8748, n8749, n8750, n8751, n8752, n8753, n8754,
    n8755, n8756, n8757, n8758, n8759, n8760, n8761, n8762, n8763, n8764,
    n8765, n8766, n8767, n8768, n8769, n8770, n8771, n8772, n8773, n8774,
    n8775, n8776, n8777, n8778, n8779, n8780, n8781, n8782, n8783, n8784,
    n8785, n8786, n8787, n8788, n8789, n8790, n8791, n8792, n8793, n8794,
    n8795, n8796, n8797, n8798, n8799, n8800, n8801, n8802, n8803, n8804,
    n8805, n8806, n8807, n8808, n8809, n8810, n8811, n8812, n8813, n8814,
    n8815, n8816, n8817, n8818, n8819, n8820, n8821, n8822, n8823, n8824,
    n8825, n8826, n8827, n8828, n8829, n8830, n8831, n8832, n8833, n8834,
    n8835, n8836, n8837, n8838, n8839, n8840, n8841, n8842, n8843, n8844,
    n8845, n8846, n8847, n8848, n8849, n8850, n8851, n8852, n8853, n8854,
    n8855, n8856, n8857, n8858, n8859, n8860, n8861, n8862, n8863, n8864,
    n8865, n8866, n8867, n8868, n8869, n8870, n8871, n8872, n8873, n8874,
    n8875, n8876, n8877, n8878, n8879, n8880, n8881, n8882, n8883, n8884,
    n8885, n8886, n8887, n8888, n8889, n8890, n8891, n8892, n8893, n8894,
    n8895, n8896, n8897, n8898, n8899, n8900, n8901, n8902, n8903, n8904,
    n8905, n8906, n8907, n8908, n8909, n8910, n8911, n8912, n8913, n8914,
    n8915, n8916, n8917, n8918, n8919, n8920, n8921, n8922, n8923, n8924,
    n8925, n8926, n8927, n8928, n8929, n8930, n8931, n8932, n8933, n8934,
    n8935, n8936, n8937, n8938, n8939, n8940, n8941, n8942, n8943, n8944,
    n8945, n8946, n8947, n8948, n8949, n8950, n8951, n8952, n8953, n8954,
    n8955, n8956, n8957, n8958, n8959, n8960, n8961, n8962, n8963, n8964,
    n8965, n8966, n8967, n8968, n8969, n8970, n8971, n8972, n8973, n8974,
    n8975, n8976, n8977, n8978, n8979, n8980, n8981, n8982, n8983, n8984,
    n8985, n8986, n8987, n8988, n8989, n8990, n8991, n8992, n8993, n8994,
    n8995, n8996, n8997, n8998, n8999, n9000, n9001, n9002, n9003, n9004,
    n9005, n9006, n9007, n9008, n9009, n9010, n9011, n9012, n9013, n9014,
    n9015, n9016, n9017, n9018, n9019, n9020, n9021, n9022, n9023, n9024,
    n9025, n9026, n9027, n9028, n9029, n9030, n9031, n9032, n9033, n9034,
    n9035, n9036, n9037, n9038, n9039, n9040, n9041, n9042, n9043, n9044,
    n9045, n9046, n9047, n9048, n9049, n9050, n9051, n9052, n9053, n9054,
    n9055, n9056, n9057, n9058, n9059, n9060, n9061, n9062, n9063, n9064,
    n9066, n9067, n9068, n9069, n9070, n9071, n9072, n9073, n9074, n9075,
    n9076, n9077, n9078, n9079, n9080, n9081, n9082, n9083, n9084, n9085,
    n9086, n9087, n9088, n9089, n9090, n9091, n9092, n9093, n9094, n9095,
    n9096, n9097, n9098, n9099, n9100, n9101, n9102, n9103, n9104, n9105,
    n9106, n9107, n9108, n9109, n9110, n9111, n9112, n9113, n9114, n9115,
    n9116, n9117, n9118, n9119, n9120, n9121, n9122, n9123, n9124, n9125,
    n9126, n9127, n9128, n9129, n9130, n9131, n9132, n9133, n9134, n9135,
    n9136, n9137, n9138, n9139, n9140, n9141, n9142, n9143, n9144, n9145,
    n9146, n9147, n9148, n9149, n9150, n9151, n9152, n9153, n9154, n9155,
    n9156, n9157, n9158, n9159, n9160, n9161, n9162, n9163, n9164, n9165,
    n9166, n9167, n9168, n9169, n9170, n9172, n9173, n9175, n9176, n9177,
    n9178, n9179, n9180, n9181, n9182, n9183, n9184, n9185, n9186, n9187,
    n9188, n9189, n9190, n9191, n9192, n9193, n9194, n9195, n9196, n9197,
    n9198, n9199, n9200, n9201, n9202, n9203, n9204, n9205, n9206, n9207,
    n9208, n9209, n9210, n9211, n9212, n9213, n9214, n9215, n9216, n9217,
    n9218, n9219, n9220, n9221, n9222, n9223, n9224, n9225, n9226, n9227,
    n9228, n9229, n9230, n9231, n9232, n9233, n9234, n9235, n9236, n9237,
    n9238, n9239, n9240, n9241, n9242, n9243, n9244, n9245, n9246, n9247,
    n9248, n9249, n9250, n9251, n9252, n9253, n9254, n9255, n9256, n9257,
    n9258, n9259, n9260, n9261, n9262, n9263, n9264, n9265, n9266, n9267,
    n9268, n9269, n9270, n9271, n9272, n9273, n9274, n9275, n9276, n9277,
    n9278, n9279, n9280, n9281, n9282, n9283, n9284, n9285, n9286, n9287,
    n9288, n9289, n9290, n9291, n9292, n9293, n9294, n9295, n9296, n9297,
    n9298, n9299, n9300, n9301, n9302, n9303, n9304, n9305, n9306, n9307,
    n9308, n9309, n9310, n9311, n9312, n9313, n9314, n9315, n9316, n9317,
    n9318, n9319, n9320, n9321, n9322, n9323, n9324, n9325, n9326, n9327,
    n9328, n9329, n9330, n9331, n9332, n9333, n9334, n9335, n9336, n9337,
    n9338, n9339, n9340, n9341, n9342, n9343, n9344, n9345, n9346, n9347,
    n9348, n9349, n9350, n9351, n9352, n9353, n9354, n9355, n9356, n9357,
    n9358, n9359, n9360, n9361, n9362, n9363, n9364, n9365, n9366, n9367,
    n9368, n9369, n9370, n9371, n9372, n9373, n9374, n9375, n9376, n9377,
    n9378, n9379, n9380, n9381, n9382, n9383, n9384, n9385, n9386, n9387,
    n9388, n9389, n9390, n9391, n9392, n9393, n9394, n9395, n9396, n9397,
    n9398, n9399, n9400, n9401, n9402, n9403, n9404, n9405, n9406, n9407,
    n9408, n9409, n9410, n9411, n9412, n9413, n9414, n9415, n9416, n9417,
    n9418, n9419, n9420, n9421, n9422, n9423, n9424, n9425, n9426, n9427,
    n9428, n9429, n9430, n9431, n9432, n9433, n9434, n9435, n9436, n9437,
    n9438, n9439, n9440, n9441, n9442, n9443, n9444, n9445, n9446, n9447,
    n9448, n9449, n9450, n9451, n9452, n9453, n9454, n9455, n9456, n9457,
    n9458, n9459, n9460, n9461, n9462, n9463, n9464, n9465, n9467, n9468,
    n9469, n9470, n9471, n9472, n9473, n9474, n9475, n9476, n9477, n9478,
    n9479, n9480, n9481, n9482, n9483, n9484, n9485, n9486, n9487, n9488,
    n9489, n9490, n9491, n9492, n9493, n9494, n9495, n9496, n9497, n9498,
    n9499, n9500, n9501, n9502, n9503, n9504, n9505, n9506, n9507, n9508,
    n9509, n9510, n9511, n9512, n9513, n9514, n9515, n9516, n9517, n9518,
    n9519, n9520, n9521, n9522, n9523, n9524, n9525, n9526, n9527, n9528,
    n9529, n9530, n9531, n9532, n9533, n9534, n9535, n9536, n9537, n9538,
    n9539, n9540, n9541, n9542, n9543, n9544, n9545, n9546, n9547, n9548,
    n9549, n9550, n9551, n9552, n9553, n9554, n9555, n9556, n9557, n9558,
    n9559, n9560, n9561, n9562, n9563, n9564, n9565, n9566, n9567, n9568,
    n9569, n9570, n9572, n9573, n9574, n9575, n9576, n9577, n9578, n9579,
    n9580, n9581, n9582, n9583, n9584, n9585, n9586, n9587, n9588, n9589,
    n9590, n9591, n9592, n9593, n9594, n9595, n9596, n9597, n9598, n9599,
    n9600, n9601, n9602, n9603, n9604, n9605, n9606, n9607, n9608, n9609,
    n9610, n9611, n9612, n9613, n9614, n9615, n9616, n9617, n9618, n9619,
    n9620, n9621, n9622, n9623, n9624, n9625, n9626, n9627, n9628, n9629,
    n9630, n9631, n9632, n9633, n9634, n9635, n9636, n9637, n9638, n9639,
    n9640, n9641, n9642, n9643, n9644, n9645, n9646, n9647, n9648, n9649,
    n9650, n9651, n9652, n9653, n9654, n9655, n9656, n9657, n9658, n9659,
    n9660, n9661, n9662, n9663, n9664, n9665, n9666, n9667, n9668, n9669,
    n9670, n9671, n9672, n9673, n9674, n9675, n9676, n9677, n9678, n9679,
    n9680, n9681, n9682, n9684, n9685, n9686, n9687, n9688, n9689, n9690,
    n9691, n9692, n9693, n9694, n9695, n9696, n9697, n9698, n9699, n9700,
    n9701, n9702, n9703, n9704, n9705, n9706, n9707, n9708, n9709, n9710,
    n9711, n9712, n9713, n9714, n9715, n9716, n9717, n9718, n9719, n9720,
    n9721, n9722, n9723, n9724, n9725, n9726, n9727, n9728, n9729, n9730,
    n9731, n9732, n9733, n9734, n9735, n9736, n9737, n9738, n9739, n9740,
    n9741, n9742, n9743, n9744, n9745, n9746, n9747, n9748, n9749, n9750,
    n9751, n9752, n9753, n9754, n9755, n9756, n9757, n9758, n9759, n9760,
    n9761, n9762, n9763, n9764, n9765, n9766, n9767, n9768, n9769, n9770,
    n9771, n9772, n9773, n9774, n9775, n9776, n9777, n9778, n9779, n9780,
    n9781, n9782, n9783, n9784, n9785, n9786, n9787, n9788, n9789, n9791,
    n9792, n9793, n9794, n9795, n9796, n9797, n9798, n9799, n9800, n9801,
    n9802, n9803, n9804, n9805, n9806, n9807, n9808, n9809, n9810, n9811,
    n9812, n9813, n9814, n9815, n9816, n9817, n9818, n9819, n9820, n9821,
    n9822, n9823, n9824, n9825, n9826, n9827, n9828, n9829, n9830, n9831,
    n9832, n9833, n9834, n9835, n9836, n9837, n9838, n9839, n9840, n9841,
    n9842, n9843, n9844, n9845, n9846, n9847, n9848, n9849, n9850, n9851,
    n9852, n9853, n9854, n9855, n9856, n9857, n9858, n9859, n9860, n9861,
    n9862, n9863, n9864, n9865, n9866, n9867, n9868, n9869, n9870, n9871,
    n9872, n9873, n9874, n9875, n9876, n9877, n9878, n9879, n9880, n9881,
    n9882, n9883, n9884, n9885, n9886, n9887, n9888, n9889, n9890, n9891,
    n9892, n9893, n9894, n9895, n9896, n9897, n9898, n9899, n9900, n9901,
    n9902, n9903, n9904, n9905, n9906, n9907, n9909, n9910, n9911, n9912,
    n9913, n9914, n9915, n9916, n9917, n9918, n9919, n9920, n9921, n9922,
    n9923, n9924, n9925, n9926, n9927, n9928, n9929, n9930, n9931, n9932,
    n9933, n9934, n9935, n9936, n9937, n9938, n9939, n9940, n9941, n9942,
    n9943, n9944, n9945, n9946, n9947, n9948, n9949, n9950, n9951, n9952,
    n9953, n9954, n9955, n9956, n9957, n9958, n9959, n9960, n9961, n9962,
    n9963, n9964, n9965, n9966, n9967, n9968, n9969, n9970, n9971, n9972,
    n9973, n9974, n9975, n9976, n9977, n9978, n9979, n9980, n9981, n9982,
    n9983, n9984, n9985, n9986, n9987, n9988, n9989, n9990, n9991, n9992,
    n9993, n9994, n9995, n9996, n9997, n9998, n9999, n10000, n10001,
    n10002, n10003, n10004, n10005, n10006, n10007, n10008, n10009, n10010,
    n10011, n10012, n10013, n10014, n10015, n10016, n10017, n10018, n10019,
    n10020, n10021, n10022, n10023, n10024, n10025, n10026, n10027, n10028,
    n10029, n10030, n10031, n10032, n10033, n10034, n10035, n10036, n10037,
    n10038, n10039, n10040, n10041, n10042, n10043, n10044, n10045, n10046,
    n10047, n10048, n10049, n10050, n10051, n10052, n10053, n10054, n10055,
    n10056, n10057, n10058, n10059, n10060, n10061, n10062, n10063, n10064,
    n10065, n10066, n10067, n10068, n10069, n10070, n10071, n10072, n10073,
    n10074, n10075, n10076, n10077, n10078, n10079, n10080, n10081, n10082,
    n10083, n10084, n10085, n10086, n10087, n10088, n10089, n10090, n10091,
    n10092, n10093, n10094, n10095, n10096, n10097, n10098, n10099, n10100,
    n10101, n10102, n10103, n10104, n10105, n10106, n10107, n10108, n10109,
    n10110, n10111, n10112, n10113, n10114, n10115, n10116, n10117, n10118,
    n10119, n10120, n10121, n10122, n10123, n10124, n10125, n10126, n10127,
    n10128, n10129, n10130, n10131, n10132, n10133, n10134, n10135, n10136,
    n10137, n10138, n10139, n10140, n10141, n10142, n10143, n10144, n10145,
    n10146, n10147, n10148, n10149, n10150, n10151, n10152, n10153, n10154,
    n10155, n10156, n10157, n10158, n10159, n10160, n10161, n10162, n10163,
    n10164, n10165, n10166, n10167, n10168, n10169, n10170, n10171, n10172,
    n10173, n10174, n10175, n10176, n10177, n10178, n10179, n10180, n10181,
    n10182, n10183, n10184, n10185, n10186, n10187, n10188, n10189, n10190,
    n10191, n10192, n10193, n10194, n10195, n10196, n10197, n10198, n10199,
    n10200, n10201, n10202, n10203, n10204, n10205, n10206, n10207, n10208,
    n10209, n10210, n10211, n10212, n10213, n10214, n10215, n10216, n10217,
    n10218, n10219, n10220, n10221, n10222, n10223, n10224, n10225, n10226,
    n10227, n10228, n10229, n10230, n10231, n10232, n10233, n10234, n10235,
    n10236, n10237, n10238, n10239, n10240, n10241, n10242, n10243, n10244,
    n10245, n10246, n10247, n10248, n10249, n10250, n10251, n10252, n10253,
    n10254, n10255, n10256, n10257, n10258, n10259, n10260, n10261, n10262,
    n10263, n10264, n10265, n10266, n10267, n10268, n10269, n10270, n10271,
    n10272, n10273, n10274, n10275, n10276, n10277, n10278, n10279, n10280,
    n10281, n10282, n10283, n10284, n10285, n10286, n10287, n10288, n10289,
    n10290, n10291, n10292, n10293, n10294, n10295, n10296, n10297, n10298,
    n10299, n10300, n10301, n10302, n10303, n10304, n10305, n10306, n10307,
    n10308, n10309, n10310, n10311, n10312, n10313, n10314, n10315, n10316,
    n10317, n10318, n10319, n10320, n10321, n10322, n10323, n10324, n10325,
    n10326, n10327, n10328, n10329, n10330, n10331, n10332, n10333, n10334,
    n10335, n10336, n10337, n10338, n10339, n10340, n10341, n10342, n10343,
    n10344, n10345, n10346, n10347, n10348, n10349, n10350, n10351, n10352,
    n10353, n10354, n10355, n10356, n10357, n10358, n10359, n10360, n10361,
    n10362, n10364, n10365, n10366, n10367, n10368, n10369, n10370, n10371,
    n10372, n10373, n10374, n10375, n10376, n10377, n10378, n10379, n10380,
    n10381, n10382, n10383, n10384, n10385, n10386, n10387, n10388, n10389,
    n10390, n10391, n10392, n10393, n10394, n10395, n10396, n10397, n10398,
    n10399, n10400, n10401, n10402, n10403, n10404, n10405, n10406, n10407,
    n10408, n10409, n10410, n10411, n10412, n10413, n10414, n10415, n10416,
    n10417, n10418, n10419, n10420, n10421, n10422, n10423, n10424, n10425,
    n10426, n10427, n10428, n10429, n10430, n10431, n10432, n10433, n10434,
    n10435, n10436, n10437, n10438, n10439, n10440, n10441, n10442, n10443,
    n10444, n10445, n10446, n10447, n10448, n10449, n10450, n10451, n10452,
    n10453, n10454, n10455, n10456, n10457, n10458, n10459, n10460, n10461,
    n10462, n10463, n10464, n10465, n10466, n10468, n10469, n10470, n10471,
    n10472, n10473, n10474, n10475, n10476, n10477, n10478, n10479, n10480,
    n10481, n10482, n10483, n10484, n10485, n10486, n10487, n10488, n10489,
    n10490, n10491, n10492, n10493, n10494, n10495, n10496, n10497, n10498,
    n10499, n10500, n10501, n10502, n10503, n10504, n10505, n10506, n10507,
    n10508, n10509, n10510, n10511, n10512, n10513, n10514, n10515, n10516,
    n10517, n10518, n10519, n10520, n10521, n10522, n10523, n10524, n10525,
    n10526, n10527, n10528, n10529, n10530, n10531, n10532, n10533, n10534,
    n10535, n10536, n10537, n10538, n10539, n10540, n10541, n10542, n10543,
    n10544, n10545, n10546, n10547, n10548, n10549, n10550, n10551, n10552,
    n10553, n10554, n10555, n10556, n10557, n10558, n10559, n10560, n10561,
    n10562, n10563, n10564, n10565, n10566, n10567, n10568, n10569, n10570,
    n10571, n10572, n10573, n10574, n10575, n10576, n10577, n10578, n10579,
    n10580, n10582, n10583, n10584, n10585, n10586, n10587, n10588, n10589,
    n10590, n10591, n10592, n10593, n10594, n10595, n10596, n10597, n10598,
    n10599, n10600, n10601, n10602, n10603, n10604, n10605, n10606, n10607,
    n10608, n10609, n10610, n10611, n10612, n10613, n10614, n10615, n10616,
    n10617, n10618, n10619, n10620, n10621, n10622, n10623, n10624, n10625,
    n10626, n10627, n10628, n10629, n10630, n10631, n10632, n10633, n10634,
    n10635, n10636, n10637, n10638, n10639, n10640, n10641, n10642, n10643,
    n10644, n10645, n10646, n10647, n10648, n10649, n10650, n10651, n10652,
    n10653, n10654, n10655, n10656, n10657, n10658, n10659, n10660, n10661,
    n10662, n10663, n10664, n10665, n10666, n10667, n10668, n10669, n10670,
    n10671, n10672, n10673, n10674, n10675, n10676, n10677, n10678, n10679,
    n10680, n10681, n10682, n10683, n10684, n10685, n10686, n10687, n10688,
    n10689, n10690, n10691, n10692, n10693, n10694, n10695, n10696, n10697,
    n10698, n10699, n10700, n10701, n10702, n10703, n10704, n10705, n10706,
    n10707, n10708, n10709, n10710, n10711, n10712, n10713, n10714, n10715,
    n10716, n10717, n10718, n10719, n10720, n10721, n10722, n10723, n10724,
    n10725, n10726, n10727, n10728, n10729, n10730, n10731, n10732, n10733,
    n10734, n10735, n10736, n10737, n10738, n10739, n10740, n10741, n10742,
    n10743, n10744, n10745, n10746, n10747, n10748, n10749, n10750, n10751,
    n10752, n10753, n10754, n10755, n10756, n10757, n10758, n10759, n10760,
    n10761, n10762, n10763, n10764, n10765, n10766, n10767, n10768, n10769,
    n10770, n10771, n10772, n10773, n10774, n10775, n10776, n10777, n10778,
    n10779, n10780, n10781, n10782, n10783, n10784, n10785, n10786, n10787,
    n10788, n10789, n10790, n10791, n10792, n10793, n10794, n10795, n10796,
    n10797, n10798, n10799, n10800, n10801, n10802, n10803, n10804, n10805,
    n10806, n10807, n10808, n10809, n10810, n10811, n10812, n10813, n10814,
    n10815, n10816, n10817, n10818, n10819, n10820, n10821, n10822, n10823,
    n10824, n10825, n10826, n10827, n10828, n10829, n10830, n10831, n10832,
    n10833, n10834, n10835, n10836, n10837, n10838, n10839, n10840, n10841,
    n10842, n10843, n10844, n10845, n10846, n10847, n10848, n10849, n10850,
    n10851, n10852, n10853, n10854, n10855, n10856, n10857, n10858, n10859,
    n10860, n10861, n10862, n10863, n10864, n10865, n10866, n10867, n10868,
    n10869, n10871, n10872, n10873, n10874, n10875, n10876, n10877, n10878,
    n10879, n10880, n10881, n10882, n10883, n10884, n10885, n10886, n10887,
    n10888, n10889, n10890, n10891, n10892, n10893, n10894, n10895, n10896,
    n10897, n10898, n10899, n10900, n10901, n10902, n10903, n10904, n10905,
    n10906, n10907, n10908, n10909, n10910, n10911, n10912, n10913, n10914,
    n10915, n10916, n10917, n10918, n10919, n10920, n10921, n10922, n10923,
    n10924, n10925, n10926, n10927, n10928, n10929, n10930, n10931, n10932,
    n10933, n10934, n10935, n10936, n10937, n10938, n10939, n10940, n10941,
    n10942, n10943, n10944, n10945, n10946, n10947, n10948, n10949, n10950,
    n10951, n10952, n10953, n10954, n10955, n10956, n10957, n10958, n10959,
    n10960, n10961, n10962, n10963, n10964, n10965, n10966, n10967, n10968,
    n10969, n10970, n10971, n10972, n10973, n10974, n10976, n10977, n10978,
    n10979, n10980, n10981, n10982, n10983, n10984, n10985, n10986, n10987,
    n10988, n10989, n10990, n10991, n10992, n10993, n10994, n10995, n10996,
    n10997, n10998, n10999, n11000, n11001, n11002, n11003, n11004, n11005,
    n11006, n11007, n11008, n11009, n11010, n11011, n11012, n11013, n11014,
    n11015, n11016, n11017, n11018, n11019, n11020, n11021, n11022, n11023,
    n11024, n11025, n11026, n11027, n11028, n11029, n11030, n11031, n11032,
    n11033, n11034, n11035, n11036, n11037, n11038, n11039, n11040, n11041,
    n11042, n11043, n11044, n11045, n11046, n11047, n11048, n11049, n11050,
    n11051, n11052, n11053, n11054, n11055, n11056, n11057, n11058, n11059,
    n11060, n11061, n11062, n11063, n11064, n11065, n11066, n11067, n11068,
    n11069, n11070, n11071, n11072, n11073, n11074, n11075, n11076, n11077,
    n11078, n11079, n11080, n11081, n11082, n11083, n11084, n11085, n11086,
    n11087, n11088, n11089, n11091, n11092, n11093, n11094, n11095, n11096,
    n11097, n11098, n11099, n11100, n11101, n11102, n11103, n11104, n11105,
    n11106, n11107, n11108, n11109, n11110, n11111, n11112, n11113, n11114,
    n11115, n11116, n11117, n11118, n11119, n11120, n11121, n11122, n11123,
    n11124, n11125, n11126, n11127, n11128, n11129, n11130, n11131, n11132,
    n11133, n11134, n11135, n11136, n11137, n11138, n11139, n11140, n11141,
    n11142, n11143, n11144, n11145, n11146, n11147, n11148, n11149, n11150,
    n11151, n11152, n11153, n11154, n11155, n11156, n11157, n11158, n11159,
    n11160, n11161, n11162, n11163, n11164, n11165, n11166, n11167, n11168,
    n11169, n11170, n11171, n11172, n11173, n11174, n11175, n11176, n11177,
    n11178, n11179, n11180, n11181, n11182, n11183, n11184, n11185, n11186,
    n11187, n11188, n11189, n11190, n11191, n11192, n11193, n11194, n11195,
    n11196, n11197, n11199, n11200, n11201, n11202, n11203, n11204, n11205,
    n11206, n11207, n11208, n11209, n11210, n11211, n11212, n11213, n11214,
    n11215, n11216, n11217, n11218, n11219, n11220, n11221, n11223, n11224,
    n11225, n11226, n11227, n11228, n11229, n11230, n11231, n11232, n11233,
    n11234, n11235, n11236, n11237, n11238, n11239, n11240, n11241, n11242,
    n11243, n11244, n11245, n11246, n11247, n11248, n11249, n11250, n11251,
    n11252, n11253, n11254, n11255, n11256, n11257, n11258, n11259, n11260,
    n11261, n11262, n11263, n11264, n11265, n11266, n11267, n11268, n11269,
    n11270, n11271, n11272, n11273, n11274, n11275, n11276, n11277, n11278,
    n11279, n11280, n11281, n11282, n11283, n11284, n11285, n11286, n11287,
    n11288, n11289, n11290, n11291, n11292, n11293, n11294, n11295, n11296,
    n11297, n11298, n11299, n11300, n11301, n11302, n11303, n11304, n11305,
    n11306, n11307, n11308, n11309, n11310, n11311, n11312, n11313, n11314,
    n11315, n11316, n11317, n11318, n11319, n11320, n11321, n11323, n11324,
    n11325, n11326, n11327, n11328, n11329, n11330, n11331, n11332, n11333,
    n11334, n11335, n11336, n11337, n11338, n11339, n11340, n11341, n11342,
    n11344, n11345, n11346, n11347, n11348, n11349, n11350, n11351, n11352,
    n11353, n11354, n11355, n11356, n11357, n11358, n11359, n11360, n11361,
    n11362, n11363, n11364, n11365, n11366, n11367, n11368, n11369, n11370,
    n11371, n11372, n11373, n11374, n11375, n11376, n11377, n11378, n11379,
    n11380, n11381, n11382, n11383, n11384, n11385, n11386, n11387, n11388,
    n11389, n11390, n11391, n11392, n11393, n11394, n11395, n11396, n11397,
    n11398, n11399, n11400, n11401, n11402, n11403, n11404, n11405, n11406,
    n11407, n11408, n11409, n11410, n11411, n11412, n11413, n11414, n11415,
    n11416, n11417, n11418, n11419, n11420, n11421, n11422, n11423, n11424,
    n11425, n11426, n11427, n11428, n11429, n11430, n11431, n11432, n11433,
    n11434, n11435, n11436, n11437, n11438, n11439, n11440, n11441, n11442,
    n11443, n11444, n11445, n11446, n11447, n11448, n11449, n11450, n11451,
    n11452, n11453, n11454, n11455, n11456, n11457, n11458, n11459, n11460,
    n11461, n11462, n11463, n11464, n11465, n11466, n11467, n11468, n11469,
    n11470, n11471, n11472, n11473, n11474, n11475, n11476, n11477, n11478,
    n11479, n11480, n11481, n11482, n11483, n11484, n11485, n11486, n11487,
    n11488, n11489, n11490, n11491, n11492, n11493, n11494, n11495, n11496,
    n11497, n11498, n11499, n11500, n11501, n11502, n11503, n11504, n11505,
    n11506, n11507, n11508, n11509, n11510, n11511, n11512, n11513, n11514,
    n11515, n11516, n11517, n11518, n11519, n11520, n11521, n11522, n11523,
    n11524, n11525, n11526, n11527, n11528, n11529, n11530, n11531, n11532,
    n11533, n11534, n11535, n11536, n11537, n11538, n11539, n11540, n11541,
    n11542, n11543, n11544, n11545, n11546, n11547, n11548, n11549, n11550,
    n11551, n11552, n11553, n11554, n11555, n11556, n11557, n11558, n11559,
    n11560, n11561, n11562, n11563, n11564, n11565, n11566, n11567, n11568,
    n11569, n11570, n11571, n11572, n11573, n11574, n11575, n11576, n11577,
    n11578, n11579, n11580, n11581, n11582, n11583, n11584, n11585, n11586,
    n11587, n11588, n11589, n11590, n11591, n11592, n11593, n11594, n11595,
    n11596, n11597, n11598, n11599, n11600, n11601, n11602, n11603, n11604,
    n11605, n11606, n11607, n11608, n11609, n11610, n11611, n11612, n11613,
    n11614, n11615, n11616, n11617, n11618, n11619, n11620, n11621, n11622,
    n11623, n11624, n11625, n11626, n11627, n11628, n11629, n11630, n11631,
    n11632, n11633, n11634, n11635, n11636, n11637, n11638, n11639, n11640,
    n11641, n11642, n11643, n11644, n11645, n11646, n11647, n11648, n11649,
    n11650, n11651, n11652, n11653, n11654, n11655, n11656, n11657, n11658,
    n11659, n11660, n11661, n11662, n11663, n11664, n11665, n11666, n11667,
    n11668, n11669, n11670, n11671, n11672, n11673, n11674, n11675, n11676,
    n11677, n11678, n11679, n11680, n11681, n11682, n11683, n11684, n11685,
    n11686, n11687, n11688, n11689, n11690, n11691, n11692, n11693, n11694,
    n11695, n11696, n11697, n11698, n11699, n11700, n11701, n11702, n11703,
    n11704, n11705, n11706, n11707, n11708, n11709, n11710, n11711, n11712,
    n11713, n11714, n11715, n11716, n11717, n11718, n11719, n11720, n11721,
    n11722, n11723, n11724, n11725, n11726, n11727, n11728, n11729, n11730,
    n11731, n11732, n11733, n11734, n11735, n11736, n11737, n11738, n11739,
    n11740, n11741, n11742, n11743, n11744, n11745, n11746, n11747, n11748,
    n11749, n11750, n11751, n11752, n11753, n11754, n11755, n11756, n11757,
    n11758, n11759, n11760, n11761, n11762, n11763, n11764, n11765, n11766,
    n11767, n11768, n11769, n11770, n11771, n11772, n11773, n11774, n11775,
    n11776, n11777, n11778, n11779, n11780, n11781, n11782, n11783, n11784,
    n11785, n11786, n11787, n11788, n11789, n11790, n11791, n11792, n11793,
    n11794, n11795, n11796, n11797, n11798, n11799, n11800, n11801, n11802,
    n11803, n11804, n11805, n11806, n11807, n11808, n11809, n11810, n11811,
    n11812, n11813, n11814, n11815, n11816, n11817, n11818, n11819, n11820,
    n11821, n11822, n11823, n11824, n11825, n11826, n11827, n11828, n11829,
    n11830, n11831, n11832, n11833, n11834, n11835, n11836, n11837, n11838,
    n11839, n11840, n11841, n11842, n11843, n11844, n11845, n11846, n11847,
    n11848, n11849, n11850, n11851, n11852, n11853, n11854, n11855, n11856,
    n11857, n11858, n11859, n11860, n11861, n11862, n11863, n11864, n11865,
    n11866, n11867, n11868, n11869, n11870, n11871, n11872, n11873, n11874,
    n11875, n11876, n11877, n11878, n11879, n11880, n11881, n11882, n11883,
    n11884, n11885, n11886, n11887, n11888, n11889, n11890, n11891, n11892,
    n11893, n11894, n11895, n11896, n11897, n11898, n11899, n11900, n11901,
    n11902, n11903, n11904, n11905, n11906, n11907, n11908, n11909, n11910,
    n11911, n11912, n11913, n11914, n11915, n11916, n11917, n11918, n11919,
    n11920, n11921, n11922, n11923, n11924, n11925, n11926, n11927, n11928,
    n11929, n11930, n11931, n11932, n11933, n11934, n11935, n11936, n11937,
    n11938, n11939, n11940, n11941, n11942, n11943, n11944, n11945, n11946,
    n11947, n11948, n11949, n11950, n11951, n11952, n11953, n11954, n11955,
    n11956, n11957, n11958, n11959, n11960, n11961, n11962, n11963, n11965,
    n11966, n11967, n11968, n11969, n11970, n11971, n11972, n11973, n11974,
    n11975, n11976, n11977, n11978, n11979, n11980, n11981, n11982, n11983,
    n11984, n11985, n11986, n11987, n11988, n11989, n11990, n11991, n11992,
    n11993, n11994, n11995, n11996, n11997, n11998, n11999, n12000, n12001,
    n12002, n12003, n12004, n12005, n12006, n12007, n12008, n12009, n12010,
    n12011, n12012, n12013, n12014, n12015, n12016, n12017, n12018, n12019,
    n12020, n12021, n12022, n12023, n12024, n12025, n12026, n12027, n12028,
    n12029, n12030, n12031, n12032, n12033, n12034, n12035, n12036, n12037,
    n12038, n12039, n12040, n12041, n12042, n12043, n12044, n12045, n12046,
    n12047, n12048, n12049, n12050, n12051, n12052, n12053, n12054, n12055,
    n12056, n12057, n12058, n12059, n12060, n12061, n12062, n12063, n12064,
    n12065, n12066, n12067, n12068, n12069, n12070, n12071, n12072, n12073,
    n12074, n12075, n12076, n12077, n12078, n12079, n12080, n12081, n12082,
    n12083, n12084, n12085, n12086, n12087, n12088, n12089, n12090, n12091,
    n12092, n12093, n12094, n12095, n12096, n12097, n12098, n12099, n12100,
    n12101, n12102, n12103, n12104, n12105, n12106, n12107, n12108, n12109,
    n12110, n12111, n12112, n12113, n12114, n12115, n12116, n12117, n12118,
    n12119, n12120, n12121, n12122, n12123, n12124, n12125, n12126, n12127,
    n12128, n12129, n12130, n12131, n12132, n12133, n12134, n12135, n12136,
    n12137, n12138, n12139, n12140, n12141, n12142, n12143, n12144, n12145,
    n12146, n12147, n12148, n12149, n12150, n12151, n12152, n12153, n12154,
    n12155, n12156, n12157, n12158, n12159, n12160, n12161, n12162, n12163,
    n12164, n12165, n12166, n12167, n12168, n12169, n12170, n12171, n12172,
    n12173, n12174, n12175, n12176, n12177, n12178, n12179, n12180, n12181,
    n12182, n12183, n12184, n12185, n12186, n12187, n12188, n12189, n12190,
    n12191, n12192, n12193, n12194, n12195, n12196, n12197, n12198, n12199,
    n12200, n12201, n12202, n12203, n12204, n12205, n12206, n12207, n12208,
    n12209, n12210, n12211, n12212, n12213, n12214, n12215, n12216, n12217,
    n12218, n12219, n12220, n12221, n12222, n12223, n12224, n12225, n12226,
    n12227, n12228, n12229, n12230, n12231, n12232, n12233, n12234, n12235,
    n12236, n12237, n12238, n12239, n12240, n12241, n12242, n12243, n12244,
    n12245, n12246, n12247, n12248, n12249, n12250, n12251, n12252, n12253,
    n12254, n12255, n12256, n12257, n12258, n12259, n12260, n12261, n12262,
    n12263, n12264, n12265, n12267, n12268, n12269, n12270, n12271, n12272,
    n12273, n12274, n12275, n12276, n12277, n12278, n12279, n12280, n12281,
    n12282, n12283, n12284, n12285, n12286, n12287, n12288, n12289, n12290,
    n12291, n12292, n12293, n12294, n12295, n12296, n12297, n12298, n12299,
    n12300, n12301, n12302, n12303, n12304, n12305, n12306, n12307, n12308,
    n12309, n12310, n12311, n12312, n12313, n12314, n12315, n12316, n12317,
    n12318, n12319, n12320, n12321, n12322, n12323, n12324, n12325, n12326,
    n12327, n12328, n12329, n12330, n12331, n12332, n12333, n12334, n12335,
    n12336, n12337, n12338, n12339, n12340, n12341, n12342, n12343, n12344,
    n12345, n12346, n12347, n12348, n12349, n12350, n12351, n12352, n12353,
    n12354, n12355, n12356, n12357, n12358, n12359, n12360, n12361, n12362,
    n12363, n12364, n12365, n12366, n12367, n12368, n12369, n12370, n12371,
    n12372, n12373, n12374, n12375, n12376, n12377, n12378, n12379, n12380,
    n12381, n12382, n12383, n12384, n12385, n12386, n12387, n12388, n12389,
    n12390, n12391, n12392, n12393, n12394, n12395, n12396, n12397, n12398,
    n12399, n12400, n12401, n12402, n12403, n12404, n12405, n12406, n12407,
    n12408, n12409, n12410, n12411, n12412, n12413, n12414, n12415, n12416,
    n12417, n12418, n12419, n12420, n12421, n12422, n12423, n12424, n12425,
    n12426, n12427, n12428, n12429, n12430, n12431, n12432, n12433, n12434,
    n12435, n12436, n12437, n12438, n12439, n12440, n12441, n12442, n12443,
    n12444, n12445, n12446, n12447, n12448, n12449, n12450, n12451, n12452,
    n12453, n12454, n12455, n12456, n12457, n12458, n12459, n12460, n12461,
    n12462, n12463, n12464, n12465, n12466, n12467, n12468, n12469, n12470,
    n12471, n12472, n12473, n12474, n12475, n12476, n12477, n12478, n12479,
    n12480, n12481, n12482, n12483, n12484, n12485, n12486, n12487, n12488,
    n12489, n12490, n12491, n12492, n12493, n12494, n12495, n12496, n12497,
    n12498, n12499, n12500, n12501, n12502, n12503, n12504, n12505, n12506,
    n12507, n12508, n12509, n12510, n12511, n12512, n12513, n12514, n12515,
    n12516, n12517, n12518, n12519, n12520, n12521, n12522, n12523, n12524,
    n12525, n12526, n12527, n12528, n12529, n12530, n12531, n12532, n12533,
    n12534, n12535, n12536, n12537, n12538, n12539, n12540, n12541, n12542,
    n12543, n12544, n12545, n12546, n12547, n12548, n12549, n12550, n12551,
    n12552, n12553, n12554, n12555, n12556, n12557, n12558, n12559, n12560,
    n12561, n12562, n12563, n12564, n12565, n12566, n12567, n12569, n12570,
    n12571, n12572, n12573, n12574, n12575, n12576, n12577, n12578, n12579,
    n12580, n12581, n12582, n12583, n12584, n12585, n12586, n12587, n12588,
    n12589, n12590, n12591, n12592, n12593, n12594, n12595, n12596, n12597,
    n12598, n12599, n12600, n12601, n12602, n12603, n12604, n12605, n12606,
    n12607, n12608, n12609, n12610, n12611, n12612, n12613, n12614, n12615,
    n12616, n12617, n12618, n12619, n12620, n12621, n12622, n12623, n12624,
    n12625, n12626, n12627, n12628, n12629, n12630, n12631, n12632, n12633,
    n12634, n12635, n12636, n12637, n12638, n12639, n12640, n12641, n12642,
    n12643, n12644, n12645, n12646, n12647, n12648, n12649, n12650, n12651,
    n12652, n12653, n12654, n12655, n12656, n12657, n12658, n12659, n12660,
    n12661, n12662, n12663, n12664, n12665, n12666, n12667, n12668, n12669,
    n12670, n12671, n12672, n12673, n12674, n12675, n12676, n12677, n12678,
    n12679, n12680, n12681, n12682, n12683, n12685, n12686, n12687, n12688,
    n12689, n12690, n12691, n12692, n12693, n12694, n12695, n12696, n12697,
    n12698, n12699, n12700, n12701, n12702, n12703, n12704, n12705, n12706,
    n12707, n12708, n12709, n12710, n12711, n12712, n12713, n12714, n12715,
    n12716, n12717, n12718, n12719, n12720, n12721, n12722, n12723, n12724,
    n12725, n12726, n12727, n12728, n12729, n12730, n12731, n12732, n12733,
    n12734, n12735, n12736, n12737, n12738, n12739, n12740, n12741, n12742,
    n12743, n12744, n12745, n12746, n12747, n12748, n12749, n12750, n12751,
    n12752, n12753, n12754, n12755, n12756, n12757, n12758, n12759, n12760,
    n12761, n12762, n12763, n12764, n12765, n12766, n12767, n12768, n12769,
    n12770, n12771, n12772, n12773, n12774, n12775, n12776, n12777, n12778,
    n12779, n12780, n12781, n12782, n12783, n12784, n12785, n12786, n12787,
    n12788, n12789, n12790, n12791, n12792, n12793, n12794, n12795, n12796,
    n12797, n12798, n12799, n12800, n12801, n12802, n12803, n12804, n12805,
    n12806, n12807, n12808, n12809, n12810, n12811, n12812, n12813, n12814,
    n12815, n12816, n12817, n12818, n12819, n12820, n12821, n12822, n12823,
    n12824, n12825, n12826, n12827, n12828, n12829, n12830, n12831, n12832,
    n12833, n12834, n12835, n12836, n12837, n12838, n12839, n12840, n12841,
    n12842, n12843, n12844, n12845, n12846, n12847, n12848, n12849, n12850,
    n12851, n12852, n12853, n12854, n12855, n12856, n12857, n12858, n12859,
    n12860, n12861, n12862, n12863, n12864, n12865, n12866, n12867, n12868,
    n12869, n12870, n12871, n12872, n12873, n12874, n12875, n12877, n12878,
    n12879, n12880, n12881, n12882, n12883, n12884, n12885, n12886, n12887,
    n12888, n12889, n12890, n12891, n12892, n12893, n12894, n12895, n12896,
    n12897, n12898, n12899, n12900, n12901, n12902, n12903, n12904, n12905,
    n12906, n12907, n12908, n12909, n12910, n12911, n12912, n12913, n12914,
    n12915, n12916, n12917, n12918, n12919, n12920, n12921, n12922, n12923,
    n12924, n12925, n12926, n12927, n12928, n12929, n12930, n12931, n12932,
    n12933, n12934, n12935, n12936, n12937, n12938, n12939, n12940, n12941,
    n12942, n12943, n12944, n12945, n12946, n12947, n12948, n12949, n12950,
    n12951, n12952, n12953, n12954, n12955, n12956, n12957, n12958, n12959,
    n12960, n12961, n12962, n12963, n12964, n12965, n12966, n12967, n12968,
    n12969, n12970, n12971, n12972, n12973, n12974, n12975, n12976, n12977,
    n12978, n12980, n12981, n12982, n12983, n12984, n12985, n12986, n12987,
    n12988, n12989, n12990, n12991, n12992, n12993, n12994, n12995, n12996,
    n12997, n12998, n12999, n13000, n13001, n13002, n13003, n13004, n13005,
    n13006, n13007, n13008, n13009, n13010, n13011, n13012, n13013, n13014,
    n13015, n13016, n13017, n13018, n13019, n13020, n13021, n13022, n13023,
    n13024, n13025, n13026, n13027, n13028, n13029, n13030, n13031, n13032,
    n13033, n13034, n13035, n13036, n13037, n13038, n13039, n13040, n13041,
    n13042, n13043, n13044, n13045, n13046, n13047, n13048, n13049, n13050,
    n13051, n13052, n13053, n13054, n13055, n13056, n13057, n13058, n13059,
    n13060, n13061, n13062, n13063, n13064, n13065, n13066, n13067, n13068,
    n13069, n13070, n13071, n13072, n13073, n13074, n13075, n13076, n13077,
    n13078, n13079, n13080, n13081, n13082, n13083, n13084, n13085, n13087,
    n13088, n13089, n13090, n13091, n13092, n13093, n13094, n13095, n13096,
    n13097, n13098, n13099, n13100, n13101, n13102, n13103, n13104, n13105,
    n13106, n13108, n13109, n13110, n13111, n13112, n13113, n13114, n13115,
    n13116, n13117, n13118, n13119, n13120, n13121, n13122, n13123, n13124,
    n13125, n13126, n13127, n13128, n13129, n13130, n13131, n13132, n13133,
    n13134, n13135, n13136, n13137, n13138, n13139, n13140, n13141, n13142,
    n13143, n13144, n13145, n13146, n13147, n13148, n13149, n13150, n13151,
    n13152, n13153, n13154, n13155, n13156, n13157, n13158, n13159, n13160,
    n13161, n13162, n13163, n13164, n13165, n13166, n13167, n13168, n13169,
    n13170, n13171, n13172, n13173, n13174, n13175, n13176, n13177, n13178,
    n13179, n13180, n13181, n13182, n13183, n13184, n13185, n13186, n13187,
    n13188, n13189, n13190, n13191, n13192, n13193, n13194, n13195, n13196,
    n13197, n13198, n13199, n13200, n13201, n13202, n13203, n13204, n13205,
    n13206, n13207, n13208, n13209, n13210, n13211, n13212, n13213, n13214,
    n13215, n13216, n13217, n13218, n13219, n13220, n13221, n13222, n13223,
    n13224, n13225, n13226, n13228, n13229, n13230, n13231, n13232, n13233,
    n13234, n13235, n13236, n13237, n13238, n13239, n13240, n13241, n13242,
    n13243, n13244, n13245, n13246, n13247, n13248, n13249, n13250, n13251,
    n13252, n13253, n13255, n13256, n13257, n13258, n13259, n13260, n13261,
    n13262, n13263, n13264, n13265, n13266, n13267, n13268, n13269, n13270,
    n13271, n13272, n13273, n13274, n13275, n13276, n13277, n13278, n13279,
    n13280, n13281, n13282, n13283, n13284, n13285, n13286, n13287, n13288,
    n13289, n13290, n13291, n13292, n13293, n13294, n13295, n13296, n13297,
    n13298, n13299, n13300, n13301, n13302, n13303, n13304, n13305, n13306,
    n13307, n13308, n13309, n13310, n13311, n13312, n13313, n13314, n13315,
    n13316, n13317, n13318, n13319, n13320, n13321, n13322, n13323, n13324,
    n13325, n13326, n13327, n13328, n13329, n13330, n13331, n13332, n13333,
    n13334, n13335, n13336, n13337, n13338, n13339, n13340, n13341, n13342,
    n13343, n13344, n13345, n13346, n13347, n13348, n13349, n13350, n13351,
    n13352, n13353, n13354, n13355, n13356, n13357, n13358, n13359, n13360,
    n13361, n13362, n13363, n13364, n13365, n13366, n13367, n13368, n13369,
    n13370, n13371, n13372, n13373, n13374, n13375, n13376, n13377, n13378,
    n13379, n13380, n13381, n13382, n13383, n13384, n13385, n13386, n13387,
    n13388, n13389, n13390, n13391, n13392, n13393, n13394, n13395, n13396,
    n13397, n13398, n13399, n13400, n13401, n13402, n13403, n13404, n13405,
    n13406, n13407, n13408, n13409, n13410, n13411, n13412, n13413, n13414,
    n13415, n13416, n13417, n13418, n13419, n13420, n13421, n13422, n13423,
    n13424, n13425, n13426, n13427, n13428, n13429, n13430, n13431, n13432,
    n13433, n13434, n13435, n13436, n13437, n13438, n13439, n13440, n13441,
    n13442, n13443, n13444, n13445, n13446, n13447, n13448, n13449, n13450,
    n13451, n13452, n13453, n13454, n13455, n13456, n13457, n13458, n13459,
    n13460, n13461, n13462, n13463, n13464, n13465, n13466, n13467, n13468,
    n13469, n13470, n13471, n13472, n13473, n13474, n13475, n13476, n13477,
    n13478, n13479, n13480, n13481, n13482, n13483, n13484, n13485, n13486,
    n13487, n13488, n13489, n13490, n13491, n13492, n13493, n13494, n13495,
    n13496, n13497, n13498, n13499, n13500, n13501, n13502, n13503, n13504,
    n13505, n13506, n13507, n13508, n13509, n13510, n13511, n13512, n13513,
    n13514, n13515, n13516, n13517, n13518, n13519, n13520, n13521, n13522,
    n13523, n13524, n13525, n13526, n13527, n13528, n13529, n13530, n13531,
    n13532, n13533, n13534, n13535, n13536, n13537, n13538, n13539, n13540,
    n13541, n13542, n13543, n13544, n13545, n13546, n13547, n13548, n13549,
    n13550, n13551, n13552, n13553, n13554, n13555, n13556, n13557, n13558,
    n13559, n13560, n13561, n13562, n13563, n13564, n13565, n13566, n13567,
    n13568, n13569, n13570, n13571, n13572, n13573, n13574, n13575, n13576,
    n13577, n13578, n13579, n13580, n13581, n13582, n13583, n13584, n13585,
    n13586, n13587, n13588, n13589, n13590, n13591, n13592, n13593, n13594,
    n13595, n13596, n13597, n13598, n13599, n13600, n13601, n13602, n13603,
    n13604, n13605, n13606, n13607, n13608, n13609, n13610, n13611, n13612,
    n13613, n13614, n13615, n13616, n13617, n13618, n13619, n13620, n13621,
    n13622, n13623, n13624, n13625, n13626, n13627, n13628, n13629, n13630,
    n13631, n13632, n13633, n13634, n13635, n13636, n13637, n13638, n13639,
    n13640, n13641, n13643, n13644, n13645, n13646, n13647, n13648, n13649,
    n13650, n13651, n13652, n13653, n13654, n13655, n13656, n13657, n13658,
    n13659, n13660, n13661, n13662, n13663, n13664, n13665, n13666, n13667,
    n13668, n13669, n13670, n13671, n13672, n13673, n13674, n13675, n13676,
    n13677, n13678, n13679, n13680, n13681, n13682, n13683, n13684, n13685,
    n13686, n13687, n13688, n13689, n13690, n13691, n13692, n13693, n13694,
    n13695, n13696, n13697, n13698, n13699, n13700, n13701, n13702, n13703,
    n13704, n13705, n13706, n13707, n13708, n13709, n13710, n13711, n13712,
    n13713, n13714, n13715, n13716, n13717, n13718, n13719, n13720, n13721,
    n13722, n13723, n13724, n13725, n13726, n13727, n13728, n13729, n13730,
    n13731, n13732, n13733, n13734, n13735, n13736, n13737, n13738, n13739,
    n13740, n13741, n13742, n13743, n13744, n13745, n13746, n13747, n13748,
    n13749, n13750, n13751, n13752, n13753, n13754, n13755, n13756, n13757,
    n13758, n13759, n13760, n13761, n13762, n13763, n13764, n13765, n13766,
    n13767, n13768, n13769, n13770, n13771, n13772, n13773, n13774, n13775,
    n13776, n13777, n13778, n13779, n13780, n13781, n13782, n13783, n13784,
    n13785, n13786, n13787, n13788, n13789, n13790, n13791, n13792, n13793,
    n13794, n13795, n13796, n13797, n13798, n13799, n13800, n13801, n13802,
    n13803, n13804, n13805, n13806, n13807, n13808, n13809, n13810, n13811,
    n13812, n13813, n13814, n13815, n13816, n13817, n13818, n13819, n13820,
    n13821, n13822, n13823, n13824, n13825, n13826, n13827, n13828, n13829,
    n13830, n13831, n13832, n13833, n13834, n13835, n13836, n13837, n13838,
    n13839, n13840, n13841, n13842, n13843, n13844, n13845, n13846, n13847,
    n13848, n13849, n13850, n13851, n13852, n13853, n13854, n13855, n13856,
    n13857, n13858, n13859, n13860, n13861, n13862, n13863, n13864, n13865,
    n13866, n13867, n13868, n13869, n13870, n13871, n13872, n13873, n13874,
    n13875, n13876, n13877, n13878, n13879, n13880, n13881, n13882, n13883,
    n13884, n13885, n13886, n13887, n13888, n13889, n13890, n13891, n13892,
    n13893, n13894, n13895, n13896, n13897, n13898, n13899, n13900, n13901,
    n13902, n13903, n13904, n13905, n13906, n13907, n13908, n13909, n13910,
    n13911, n13912, n13913, n13914, n13915, n13916, n13917, n13918, n13919,
    n13920, n13921, n13922, n13923, n13924, n13925, n13926, n13927, n13928,
    n13929, n13930, n13931, n13932, n13933, n13934, n13935, n13936, n13937,
    n13938, n13939, n13940, n13941, n13942, n13943, n13944, n13945, n13946,
    n13947, n13948, n13949, n13950, n13951, n13952, n13953, n13954, n13955,
    n13956, n13957, n13958, n13959, n13960, n13961, n13962, n13963, n13964,
    n13965, n13966, n13967, n13968, n13969, n13970, n13971, n13972, n13973,
    n13974, n13975, n13976, n13977, n13978, n13979, n13980, n13981, n13982,
    n13983, n13984, n13985, n13986, n13987, n13988, n13989, n13990, n13991,
    n13992, n13993, n13994, n13995, n13996, n13997, n13998, n13999, n14000,
    n14001, n14003, n14004, n14005, n14006, n14007, n14008, n14009, n14010,
    n14011, n14012, n14013, n14014, n14015, n14016, n14017, n14018, n14019,
    n14020, n14021, n14022, n14023, n14024, n14025, n14026, n14027, n14028,
    n14029, n14030, n14031, n14032, n14033, n14034, n14035, n14036, n14037,
    n14038, n14039, n14040, n14041, n14042, n14043, n14044, n14045, n14046,
    n14047, n14048, n14049, n14050, n14051, n14052, n14053, n14054, n14055,
    n14056, n14057, n14058, n14059, n14060, n14061, n14062, n14063, n14064,
    n14065, n14066, n14067, n14068, n14069, n14070, n14071, n14072, n14073,
    n14074, n14075, n14076, n14077, n14078, n14079, n14080, n14081, n14082,
    n14083, n14084, n14085, n14086, n14087, n14088, n14089, n14090, n14091,
    n14092, n14093, n14094, n14095, n14096, n14097, n14098, n14099, n14100,
    n14101, n14102, n14103, n14104, n14105, n14106, n14107, n14108, n14109,
    n14110, n14111, n14112, n14113, n14114, n14115, n14116, n14117, n14118,
    n14119, n14120, n14121, n14122, n14123, n14124, n14125, n14126, n14127,
    n14128, n14129, n14130, n14131, n14132, n14133, n14134, n14135, n14136,
    n14137, n14138, n14139, n14140, n14141, n14142, n14143, n14144, n14145,
    n14146, n14147, n14148, n14149, n14150, n14151, n14152, n14153, n14154,
    n14155, n14156, n14157, n14158, n14159, n14160, n14161, n14162, n14163,
    n14164, n14165, n14166, n14167, n14168, n14169, n14170, n14171, n14172,
    n14173, n14174, n14175, n14176, n14177, n14178, n14179, n14180, n14181,
    n14182, n14183, n14184, n14185, n14187, n14188, n14189, n14190, n14191,
    n14192, n14193, n14194, n14195, n14196, n14197, n14198, n14199, n14200,
    n14201, n14202, n14203, n14204, n14206, n14207, n14208, n14209, n14210,
    n14211, n14212, n14213, n14214, n14215, n14216, n14217, n14218, n14219,
    n14220, n14221, n14222, n14224, n14225, n14226, n14227, n14228, n14229,
    n14230, n14231, n14232, n14233, n14234, n14235, n14236, n14237, n14238,
    n14239, n14240, n14241, n14242, n14243, n14244, n14245, n14246, n14247,
    n14248, n14249, n14250, n14251, n14252, n14253, n14254, n14255, n14256,
    n14257, n14258, n14259, n14260, n14261, n14262, n14263, n14264, n14265,
    n14266, n14267, n14268, n14269, n14270, n14271, n14272, n14273, n14274,
    n14275, n14276, n14277, n14278, n14279, n14280, n14281, n14282, n14283,
    n14284, n14285, n14286, n14287, n14288, n14289, n14290, n14291, n14292,
    n14293, n14294, n14295, n14296, n14297, n14298, n14299, n14300, n14301,
    n14302, n14303, n14304, n14305, n14306, n14307, n14308, n14309, n14310,
    n14311, n14312, n14313, n14314, n14315, n14316, n14317, n14318, n14319,
    n14320, n14321, n14322, n14323, n14324, n14325, n14326, n14327, n14328,
    n14329, n14330, n14331, n14332, n14333, n14334, n14335, n14336, n14337,
    n14338, n14339, n14340, n14341, n14342, n14343, n14344, n14345, n14346,
    n14347, n14348, n14349, n14350, n14351, n14352, n14353, n14354, n14355,
    n14356, n14357, n14358, n14359, n14360, n14361, n14362, n14363, n14364,
    n14365, n14366, n14367, n14368, n14369, n14370, n14371, n14372, n14373,
    n14374, n14375, n14376, n14377, n14378, n14379, n14380, n14381, n14382,
    n14383, n14384, n14385, n14386, n14387, n14388, n14389, n14390, n14391,
    n14392, n14393, n14394, n14395, n14396, n14397, n14398, n14399, n14400,
    n14401, n14402, n14403, n14404, n14405, n14406, n14407, n14408, n14409,
    n14410, n14411, n14412, n14413, n14414, n14415, n14416, n14417, n14418,
    n14419, n14420, n14421, n14422, n14423, n14424, n14425, n14426, n14427,
    n14428, n14429, n14430, n14431, n14432, n14433, n14434, n14435, n14436,
    n14437, n14438, n14439, n14440, n14441, n14442, n14443, n14444, n14445,
    n14446, n14447, n14448, n14449, n14450, n14451, n14452, n14453, n14454,
    n14455, n14456, n14457, n14458, n14459, n14460, n14461, n14462, n14463,
    n14464, n14465, n14466, n14467, n14468, n14469, n14470, n14471, n14472,
    n14473, n14474, n14475, n14476, n14477, n14478, n14479, n14480, n14481,
    n14482, n14483, n14484, n14485, n14486, n14487, n14488, n14489, n14490,
    n14491, n14492, n14493, n14494, n14495, n14496, n14497, n14498, n14499,
    n14500, n14501, n14502, n14503, n14504, n14505, n14506, n14507, n14508,
    n14509, n14510, n14511, n14512, n14513, n14514, n14515, n14516, n14517,
    n14518, n14519, n14520, n14521, n14522, n14523, n14524, n14525, n14526,
    n14527, n14528, n14529, n14530, n14531, n14532, n14533, n14534, n14535,
    n14536, n14537, n14538, n14539, n14540, n14541, n14542, n14543, n14544,
    n14545, n14546, n14547, n14548, n14549, n14550, n14551, n14552, n14553,
    n14554, n14555, n14556, n14557, n14558, n14559, n14560, n14561, n14562,
    n14563, n14564, n14565, n14566, n14567, n14568, n14569, n14570, n14571,
    n14572, n14573, n14574, n14575, n14576, n14577, n14578, n14579, n14580,
    n14581, n14582, n14583, n14584, n14585, n14586, n14587, n14588, n14589,
    n14590, n14591, n14592, n14593, n14594, n14595, n14596, n14597, n14598,
    n14599, n14600, n14601, n14602, n14603, n14604, n14605, n14606, n14607,
    n14608, n14609, n14610, n14611, n14612, n14613, n14614, n14615, n14616,
    n14617, n14618, n14619, n14620, n14621, n14622, n14623, n14624, n14625,
    n14626, n14627, n14628, n14629, n14630, n14631, n14632, n14633, n14634,
    n14635, n14636, n14637, n14638, n14639, n14640, n14641, n14642, n14643,
    n14644, n14645, n14646, n14647, n14648, n14649, n14650, n14651, n14652,
    n14653, n14654, n14655, n14656, n14657, n14658, n14659, n14660, n14661,
    n14662, n14663, n14664, n14665, n14666, n14667, n14668, n14669, n14670,
    n14671, n14672, n14673, n14674, n14676, n14677, n14678, n14679, n14680,
    n14681, n14682, n14683, n14684, n14685, n14686, n14687, n14688, n14689,
    n14690, n14691, n14692, n14693, n14694, n14695, n14696, n14697, n14698,
    n14699, n14700, n14701, n14702, n14703, n14704, n14705, n14706, n14707,
    n14708, n14709, n14710, n14711, n14712, n14713, n14714, n14715, n14716,
    n14717, n14718, n14719, n14720, n14721, n14722, n14723, n14724, n14725,
    n14726, n14727, n14728, n14729, n14730, n14731, n14732, n14733, n14734,
    n14735, n14736, n14737, n14738, n14739, n14740, n14741, n14742, n14743,
    n14744, n14745, n14746, n14747, n14748, n14749, n14750, n14751, n14752,
    n14753, n14754, n14755, n14756, n14757, n14758, n14759, n14760, n14761,
    n14762, n14763, n14764, n14765, n14766, n14767, n14768, n14769, n14770,
    n14771, n14772, n14773, n14774, n14775, n14776, n14777, n14778, n14779,
    n14780, n14781, n14782, n14783, n14784, n14785, n14786, n14787, n14788,
    n14789, n14790, n14791, n14792, n14793, n14794, n14795, n14796, n14797,
    n14798, n14799, n14800, n14801, n14802, n14803, n14804, n14805, n14806,
    n14807, n14808, n14809, n14810, n14811, n14812, n14813, n14814, n14815,
    n14816, n14817, n14818, n14819, n14820, n14821, n14822, n14823, n14824,
    n14825, n14826, n14827, n14828, n14829, n14830, n14831, n14832, n14833,
    n14834, n14835, n14836, n14837, n14838, n14839, n14840, n14841, n14842,
    n14843, n14844, n14845, n14846, n14847, n14848, n14849, n14850, n14851,
    n14852, n14853, n14854, n14855, n14856, n14857, n14858, n14859, n14860,
    n14862, n14863, n14864, n14865, n14866, n14867, n14868, n14869, n14870,
    n14871, n14872, n14873, n14874, n14875, n14876, n14877, n14878, n14879,
    n14880, n14881, n14882, n14883, n14884, n14885, n14886, n14887, n14888,
    n14889, n14890, n14891, n14892, n14893, n14894, n14895, n14896, n14897,
    n14898, n14899, n14900, n14901, n14902, n14903, n14904, n14905, n14906,
    n14907, n14908, n14909, n14910, n14911, n14912, n14913, n14914, n14915,
    n14916, n14917, n14918, n14919, n14920, n14921, n14922, n14923, n14924,
    n14925, n14926, n14927, n14928, n14929, n14930, n14931, n14932, n14933,
    n14934, n14935, n14936, n14937, n14938, n14939, n14940, n14941, n14942,
    n14943, n14944, n14945, n14946, n14947, n14948, n14949, n14950, n14951,
    n14952, n14953, n14954, n14955, n14956, n14957, n14958, n14959, n14960,
    n14961, n14962, n14963, n14964, n14965, n14966, n14967, n14968, n14969,
    n14970, n14971, n14972, n14973, n14974, n14976, n14977, n14978, n14979,
    n14980, n14981, n14982, n14983, n14984, n14985, n14986, n14987, n14988,
    n14989, n14990, n14991, n14992, n14993, n14994, n14995, n14996, n14997,
    n14998, n15000, n15001, n15002, n15003, n15004, n15005, n15006, n15007,
    n15008, n15009, n15010, n15011, n15012, n15013, n15014, n15015, n15016,
    n15018, n15019, n15020, n15021, n15022, n15023, n15024, n15025, n15026,
    n15027, n15028, n15029, n15030, n15031, n15032, n15033, n15034, n15036,
    n15037, n15038, n15039, n15040, n15041, n15042, n15043, n15044, n15045,
    n15046, n15047, n15048, n15049, n15050, n15051, n15052, n15053, n15054,
    n15055, n15056, n15057, n15058, n15059, n15060, n15061, n15062, n15063,
    n15064, n15065, n15066, n15067, n15068, n15069, n15070, n15071, n15072,
    n15073, n15074, n15075, n15076, n15077, n15078, n15079, n15080, n15081,
    n15082, n15083, n15084, n15085, n15086, n15087, n15088, n15089, n15090,
    n15091, n15092, n15093, n15094, n15095, n15096, n15097, n15098, n15099,
    n15100, n15101, n15102, n15103, n15104, n15105, n15106, n15107, n15108,
    n15109, n15110, n15111, n15112, n15113, n15114, n15115, n15116, n15117,
    n15118, n15119, n15120, n15121, n15122, n15123, n15124, n15125, n15126,
    n15127, n15128, n15129, n15130, n15131, n15132, n15133, n15134, n15135,
    n15136, n15137, n15138, n15139, n15140, n15141, n15142, n15144, n15145,
    n15146, n15147, n15148, n15149, n15150, n15151, n15152, n15153, n15154,
    n15155, n15156, n15157, n15158, n15159, n15160, n15161, n15162, n15163,
    n15165, n15166, n15167, n15168, n15169, n15170, n15171, n15172, n15173,
    n15174, n15175, n15176, n15177, n15178, n15179, n15180, n15181, n15183,
    n15184, n15185, n15186, n15187, n15188, n15189, n15190, n15191, n15192,
    n15193, n15194, n15195, n15196, n15197, n15198, n15199, n15200, n15201,
    n15202, n15203, n15204, n15205, n15206, n15207, n15208, n15209, n15210,
    n15211, n15212, n15213, n15214, n15215, n15216, n15217, n15218, n15219,
    n15220, n15221, n15222, n15223, n15224, n15225, n15226, n15227, n15228,
    n15229, n15230, n15231, n15232, n15233, n15234, n15235, n15236, n15237,
    n15238, n15239, n15240, n15241, n15242, n15243, n15244, n15245, n15246,
    n15247, n15248, n15249, n15250, n15251, n15252, n15253, n15254, n15255,
    n15256, n15257, n15258, n15259, n15260, n15261, n15262, n15263, n15264,
    n15265, n15266, n15267, n15268, n15269, n15270, n15271, n15272, n15273,
    n15274, n15275, n15276, n15277, n15278, n15279, n15280, n15281, n15282,
    n15283, n15284, n15285, n15286, n15287, n15288, n15290, n15291, n15292,
    n15293, n15294, n15295, n15296, n15297, n15298, n15299, n15300, n15301,
    n15302, n15303, n15304, n15305, n15306, n15307, n15308, n15309, n15311,
    n15312, n15313, n15314, n15315, n15316, n15317, n15318, n15319, n15320,
    n15321, n15322, n15323, n15324, n15325, n15326, n15327, n15329, n15330,
    n15331, n15332, n15333, n15334, n15335, n15336, n15337, n15338, n15339,
    n15340, n15341, n15342, n15343, n15344, n15345, n15346, n15347, n15348,
    n15349, n15350, n15351, n15352, n15353, n15354, n15356, n15357, n15358,
    n15359, n15360, n15361, n15362, n15363, n15364, n15365, n15366, n15367,
    n15368, n15369, n15370, n15371, n15372, n15373, n15374, n15375, n15376,
    n15377, n15378, n15379, n15380, n15381, n15383, n15384, n15385, n15386,
    n15387, n15388, n15389, n15390, n15391, n15392, n15393, n15394, n15395,
    n15396, n15397, n15398, n15399, n15400, n15401, n15402, n15404, n15405,
    n15406, n15407, n15408, n15409, n15410, n15411, n15412, n15413, n15414,
    n15415, n15416, n15417, n15418, n15419, n15420, n15421, n15422, n15423,
    n15424, n15425, n15426, n15427, n15428, n15429, n15430, n15431, n15432,
    n15433, n15434, n15435, n15436, n15437, n15438, n15439, n15440, n15441,
    n15442, n15443, n15444, n15445, n15446, n15447, n15448, n15449, n15450,
    n15451, n15452, n15453, n15454, n15455, n15456, n15457, n15458, n15459,
    n15460, n15461, n15462, n15463, n15464, n15465, n15466, n15467, n15468,
    n15469, n15470, n15471, n15472, n15473, n15474, n15475, n15476, n15477,
    n15478, n15479, n15480, n15481, n15482, n15483, n15484, n15485, n15486,
    n15487, n15488, n15489, n15490, n15491, n15492, n15493, n15494, n15495,
    n15496, n15497, n15498, n15499, n15500, n15501, n15502, n15503, n15504,
    n15505, n15506, n15507, n15508, n15509, n15510, n15511, n15512, n15513,
    n15514, n15515, n15516, n15517, n15518, n15519, n15520, n15521, n15522,
    n15523, n15524, n15525, n15526, n15527, n15528, n15529, n15530, n15531,
    n15532, n15533, n15534, n15535, n15536, n15537, n15538, n15539, n15540,
    n15541, n15542, n15543, n15544, n15545, n15546, n15547, n15548, n15549,
    n15550, n15551, n15552, n15553, n15554, n15555, n15556, n15557, n15558,
    n15559, n15560, n15561, n15562, n15563, n15564, n15565, n15566, n15567,
    n15568, n15569, n15570, n15571, n15572, n15573, n15574, n15575, n15576,
    n15577, n15578, n15579, n15580, n15581, n15582, n15583, n15584, n15585,
    n15586, n15587, n15588, n15589, n15590, n15591, n15592, n15593, n15594,
    n15595, n15596, n15597, n15598, n15599, n15600, n15601, n15602, n15603,
    n15604, n15605, n15606, n15607, n15608, n15609, n15610, n15611, n15612,
    n15613, n15614, n15615, n15616, n15617, n15618, n15619, n15620, n15621,
    n15622, n15623, n15624, n15625, n15626, n15627, n15628, n15629, n15630,
    n15631, n15632, n15633, n15634, n15635, n15636, n15637, n15638, n15639,
    n15640, n15641, n15642, n15643, n15644, n15645, n15646, n15647, n15648,
    n15649, n15650, n15651, n15652, n15653, n15654, n15655, n15656, n15657,
    n15658, n15659, n15660, n15662, n15663, n15664, n15665, n15666, n15667,
    n15668, n15669, n15670, n15671, n15672, n15673, n15674, n15675, n15676,
    n15677, n15678, n15679, n15680, n15681, n15682, n15683, n15684, n15685,
    n15686, n15687, n15688, n15689, n15690, n15691, n15692, n15693, n15694,
    n15695, n15696, n15697, n15698, n15699, n15700, n15701, n15702, n15703,
    n15704, n15705, n15706, n15707, n15708, n15709, n15710, n15711, n15712,
    n15713, n15714, n15715, n15716, n15717, n15718, n15719, n15720, n15721,
    n15722, n15723, n15724, n15725, n15726, n15727, n15728, n15729, n15730,
    n15731, n15732, n15733, n15734, n15735, n15736, n15737, n15738, n15739,
    n15740, n15741, n15742, n15743, n15744, n15745, n15746, n15747, n15748,
    n15749, n15750, n15751, n15752, n15753, n15754, n15755, n15756, n15757,
    n15758, n15759, n15760, n15761, n15762, n15763, n15765, n15766, n15767,
    n15768, n15769, n15770, n15771, n15772, n15773, n15774, n15775, n15776,
    n15777, n15778, n15779, n15780, n15781, n15782, n15783, n15784, n15786,
    n15787, n15788, n15789, n15790, n15791, n15792, n15793, n15794, n15795,
    n15796, n15797, n15798, n15799, n15800, n15801, n15802, n15804, n15805,
    n15806, n15807, n15808, n15809, n15810, n15811, n15812, n15813, n15814,
    n15815, n15816, n15817, n15818, n15819, n15820, n15821, n15822, n15823,
    n15824, n15825, n15826, n15827, n15828, n15829, n15830, n15832, n15833,
    n15834, n15835, n15836, n15837, n15838, n15839, n15840, n15841, n15842,
    n15843, n15844, n15845, n15846, n15847, n15848, n15849, n15850, n15851,
    n15852, n15853, n15854, n15855, n15856, n15857, n15858, n15859, n15860,
    n15861, n15862, n15863, n15864, n15865, n15866, n15867, n15868, n15869,
    n15870, n15871, n15872, n15873, n15874, n15875, n15876, n15877, n15878,
    n15879, n15880, n15881, n15882, n15883, n15884, n15885, n15886, n15887,
    n15888, n15889, n15890, n15891, n15892, n15893, n15894, n15895, n15896,
    n15897, n15898, n15899, n15900, n15901, n15902, n15903, n15904, n15905,
    n15906, n15907, n15908, n15909, n15910, n15911, n15912, n15913, n15914,
    n15915, n15916, n15917, n15918, n15919, n15920, n15921, n15922, n15923,
    n15924, n15925, n15926, n15927, n15928, n15929, n15930, n15931, n15932,
    n15933, n15935, n15936, n15937, n15938, n15939, n15940, n15941, n15942,
    n15943, n15944, n15945, n15946, n15947, n15948, n15949, n15950, n15951,
    n15952, n15953, n15954, n15955, n15956, n15957, n15958, n15959, n15960,
    n15961, n15962, n15963, n15964, n15965, n15966, n15967, n15968, n15969,
    n15970, n15971, n15972, n15973, n15974, n15975, n15976, n15977, n15978,
    n15979, n15980, n15981, n15982, n15983, n15984, n15985, n15986, n15987,
    n15988, n15989, n15990, n15991, n15992, n15993, n15994, n15995, n15996,
    n15997, n15998, n15999, n16000, n16001, n16002, n16003, n16004, n16005,
    n16006, n16007, n16008, n16009, n16010, n16011, n16012, n16013, n16014,
    n16015, n16016, n16017, n16018, n16019, n16020, n16021, n16022, n16023,
    n16024, n16025, n16026, n16027, n16028, n16029, n16030, n16031, n16032,
    n16033, n16034, n16035, n16036, n16037, n16038, n16039, n16040, n16042,
    n16043, n16044, n16045, n16046, n16047, n16048, n16049, n16050, n16051,
    n16052, n16053, n16054, n16055, n16056, n16057, n16058, n16059, n16060,
    n16061, n16063, n16064, n16065, n16066, n16067, n16068, n16069, n16070,
    n16071, n16072, n16073, n16074, n16075, n16076, n16077, n16078, n16079,
    n16080, n16081, n16082, n16084, n16085, n16086, n16087, n16088, n16089,
    n16090, n16091, n16092, n16093, n16094, n16095, n16096, n16097, n16098,
    n16099, n16100, n16101, n16102, n16103, n16105, n16106, n16107, n16108,
    n16109, n16110, n16111, n16112, n16113, n16114, n16115, n16116, n16117,
    n16118, n16119, n16120, n16121, n16122, n16123, n16124, n16125, n16126,
    n16127, n16129, n16130, n16131, n16132, n16133, n16134, n16135, n16136,
    n16137, n16138, n16139, n16140, n16141, n16142, n16143, n16144, n16145,
    n16147, n16148, n16149, n16150, n16151, n16152, n16153, n16154, n16155,
    n16156, n16157, n16158, n16159, n16160, n16161, n16162, n16163, n16164,
    n16165, n16166, n16168, n16169, n16170, n16171, n16172, n16173, n16174,
    n16175, n16176, n16177, n16178, n16179, n16180, n16181, n16182, n16183,
    n16184, n16185, n16186, n16187, n16188, n16189, n16190, n16191, n16192,
    n16193, n16194, n16195, n16196, n16197, n16198, n16199, n16200, n16201,
    n16202, n16203, n16204, n16205, n16206, n16207, n16208, n16209, n16210,
    n16211, n16212, n16213, n16214, n16215, n16216, n16217, n16218, n16219,
    n16220, n16221, n16222, n16223, n16224, n16225, n16226, n16227, n16228,
    n16229, n16230, n16231, n16232, n16233, n16234, n16235, n16236, n16237,
    n16238, n16239, n16240, n16241, n16242, n16243, n16244, n16245, n16246,
    n16247, n16248, n16249, n16250, n16251, n16252, n16253, n16254, n16255,
    n16256, n16257, n16258, n16259, n16260, n16261, n16262, n16263, n16264,
    n16265, n16266, n16267, n16268, n16269, n16270, n16271, n16272, n16273,
    n16275, n16276, n16277, n16278, n16279, n16280, n16281, n16282, n16283,
    n16284, n16285, n16286, n16287, n16288, n16289, n16290, n16291, n16292,
    n16293, n16294, n16296, n16297, n16298, n16299, n16300, n16301, n16302,
    n16303, n16304, n16305, n16306, n16307, n16308, n16309, n16310, n16311,
    n16312, n16313, n16314, n16315, n16316, n16317, n16318, n16319, n16320,
    n16321, n16323, n16324, n16325, n16326, n16327, n16328, n16329, n16330,
    n16331, n16332, n16333, n16334, n16335, n16336, n16337, n16338, n16339,
    n16340, n16341, n16342, n16343, n16344, n16345, n16346, n16347, n16348,
    n16349, n16350, n16351, n16352, n16353, n16354, n16355, n16356, n16357,
    n16358, n16359, n16360, n16361, n16362, n16363, n16364, n16365, n16366,
    n16367, n16368, n16369, n16370, n16371, n16372, n16373, n16374, n16375,
    n16376, n16377, n16378, n16379, n16380, n16381, n16382, n16383, n16384,
    n16385, n16386, n16387, n16388, n16389, n16390, n16391, n16392, n16393,
    n16394, n16395, n16396, n16397, n16398, n16399, n16400, n16401, n16402,
    n16403, n16404, n16405, n16406, n16407, n16408, n16409, n16410, n16411,
    n16412, n16413, n16414, n16415, n16416, n16417, n16418, n16419, n16420,
    n16422, n16423, n16424, n16425, n16426, n16427, n16428, n16429, n16430,
    n16431, n16432, n16433, n16434, n16435, n16436, n16437, n16438, n16439,
    n16440, n16441, n16443, n16444, n16445, n16446, n16447, n16448, n16449,
    n16450, n16451, n16452, n16453, n16454, n16455, n16456, n16457, n16458,
    n16459, n16460, n16461, n16462, n16464, n16465, n16466, n16467, n16468,
    n16469, n16470, n16471, n16472, n16473, n16474, n16475, n16476, n16477,
    n16478, n16479, n16480, n16481, n16482, n16483, n16484, n16486, n16487,
    n16488, n16489, n16490, n16491, n16492, n16493, n16494, n16495, n16496,
    n16497, n16498, n16499, n16500, n16501, n16502, n16504, n16505, n16506,
    n16507, n16508, n16509, n16510, n16511, n16512, n16513, n16514, n16515,
    n16516, n16517, n16518, n16519, n16520, n16522, n16523, n16524, n16525,
    n16526, n16527, n16528, n16529, n16530, n16531, n16532, n16533, n16534,
    n16535, n16536, n16537, n16538, n16540, n16541, n16542, n16543, n16544,
    n16545, n16546, n16547, n16548, n16549, n16550, n16551, n16552, n16553,
    n16554, n16555, n16556, n16558, n16559, n16560, n16561, n16562, n16563,
    n16564, n16565, n16566, n16567, n16568, n16569, n16570, n16571, n16572,
    n16573, n16574, n16575, n16576, n16577, n16579, n16580, n16581, n16582,
    n16583, n16584, n16585, n16586, n16587, n16588, n16589, n16590, n16591,
    n16592, n16593, n16594, n16595, n16597, n16598, n16599, n16600, n16601,
    n16602, n16603, n16604, n16605, n16606, n16607, n16608, n16609, n16610,
    n16611, n16612, n16613, n16615, n16616, n16617, n16618, n16619, n16620,
    n16621, n16622, n16623, n16624, n16625, n16626, n16627, n16628, n16629,
    n16630, n16631, n16632, n16633, n16634, n16635, n16636, n16637, n16639,
    n16640, n16641, n16642, n16643, n16644, n16645, n16646, n16647, n16648,
    n16649, n16650, n16651, n16652, n16653, n16654, n16655, n16656, n16657,
    n16658, n16660, n16661, n16662, n16663, n16664, n16665, n16666, n16667,
    n16668, n16669, n16670, n16671, n16672, n16673, n16674, n16675, n16676,
    n16677, n16678, n16679, n16680, n16682, n16683, n16684, n16685, n16686,
    n16687, n16688, n16689, n16690, n16691, n16692, n16693, n16694, n16695,
    n16696, n16697, n16698, n16700, n16701, n16702, n16703, n16704, n16705,
    n16706, n16707, n16708, n16709, n16710, n16711, n16712, n16713, n16714,
    n16715, n16716, n16718, n16719, n16720, n16721, n16722, n16723, n16724,
    n16725, n16726, n16727, n16728, n16729, n16730, n16731, n16732, n16733,
    n16734, n16735, n16736, n16737, n16739, n16740, n16741, n16742, n16743,
    n16744, n16745, n16746, n16747, n16748, n16749, n16750, n16751, n16752,
    n16753, n16754, n16755, n16757, n16758, n16759, n16760, n16761, n16762,
    n16763, n16764, n16765, n16766, n16767, n16768, n16769, n16770, n16771,
    n16772, n16773, n16774, n16775, n16776, n16778, n16779, n16780, n16781,
    n16782, n16783, n16784, n16785, n16786, n16787, n16788, n16789, n16790,
    n16791, n16792, n16793, n16794, n16795, n16796, n16797, n16799, n16800,
    n16801, n16802, n16803, n16804, n16805, n16806, n16807, n16808, n16809,
    n16810, n16811, n16812, n16813, n16814, n16815, n16817, n16818, n16819,
    n16820, n16821, n16822, n16823, n16824, n16825, n16826, n16827, n16828,
    n16829, n16830, n16831, n16832, n16833, n16835, n16836, n16837, n16838,
    n16839, n16840, n16841, n16842, n16843, n16844, n16845, n16846, n16847,
    n16848, n16849, n16850, n16851, n16852, n16853, n16854, n16856, n16857,
    n16858, n16859, n16860, n16861, n16862, n16863, n16864, n16865, n16866,
    n16867, n16868, n16869, n16870, n16871, n16872, n16874, n16875, n16876,
    n16877, n16878, n16879, n16880, n16881, n16882, n16883, n16884, n16885,
    n16886, n16887, n16888, n16889, n16890, n16891, n16892, n16893, n16895,
    n16896, n16897, n16898, n16899, n16900, n16901, n16902, n16903, n16904,
    n16905, n16906, n16907, n16908, n16909, n16910, n16911, n16912, n16913,
    n16914, n16916, n16917, n16918, n16919, n16920, n16921, n16922, n16923,
    n16924, n16925, n16926, n16927, n16928, n16929, n16930, n16931, n16932,
    n16933, n16934, n16935, n16936, n16937, n16938, n16939, n16940, n16941,
    n16943, n16944, n16945, n16946, n16947, n16948, n16949, n16950, n16951,
    n16952, n16953, n16954, n16955, n16956, n16957, n16958, n16959, n16960,
    n16961, n16962, n16963, n16965, n16966, n16967, n16968, n16969, n16970,
    n16971, n16972, n16973, n16974, n16975, n16976, n16977, n16978, n16979,
    n16980, n16981, n16983, n16984, n16985, n16986, n16987, n16988, n16989,
    n16990, n16991, n16992, n16993, n16994, n16995, n16996, n16997, n16998,
    n16999, n17001, n17002, n17003, n17004, n17005, n17006, n17007, n17008,
    n17009, n17010, n17011, n17012, n17013, n17014, n17015, n17016, n17017,
    n17018, n17019, n17020, n17022, n17023, n17024, n17025, n17026, n17027,
    n17028, n17029, n17030, n17031, n17032, n17033, n17034, n17035, n17036,
    n17037, n17038, n17040, n17041, n17042, n17043, n17044, n17045, n17046,
    n17047, n17048, n17049, n17050, n17051, n17052, n17053, n17054, n17055,
    n17056, n17057, n17058, n17059, n17061, n17062, n17063, n17064, n17065,
    n17066, n17067, n17068, n17069, n17070, n17071, n17072, n17073, n17074,
    n17075, n17076, n17077, n17079, n17080, n17081, n17082, n17083, n17084,
    n17085, n17086, n17087, n17088, n17089, n17090, n17091, n17092, n17093,
    n17094, n17095, n17096, n17097, n17098, n17100, n17101, n17102, n17103,
    n17104, n17105, n17106, n17107, n17108, n17109, n17110, n17111, n17112,
    n17113, n17114, n17115, n17116, n17118, n17119, n17120, n17121, n17122,
    n17123, n17124, n17125, n17126, n17127, n17128, n17129, n17130, n17131,
    n17132, n17133, n17134, n17135, n17136, n17137, n17138, n17140, n17141,
    n17142, n17143, n17144, n17145, n17146, n17147, n17148, n17149, n17150,
    n17151, n17152, n17153, n17154, n17155, n17156, n17158, n17159, n17160,
    n17161, n17162, n17163, n17164, n17165, n17166, n17167, n17168, n17169,
    n17170, n17171, n17172, n17173, n17174, n17175, n17176, n17177, n17179,
    n17180, n17181, n17182, n17183, n17184, n17185, n17186, n17187, n17188,
    n17189, n17190, n17191, n17192, n17193, n17194, n17195, n17197, n17198,
    n17199, n17200, n17201, n17202, n17203, n17204, n17205, n17206, n17207,
    n17208, n17209, n17210, n17211, n17212, n17213, n17215, n17216, n17217,
    n17218, n17219, n17220, n17221, n17222, n17223, n17224, n17225, n17226,
    n17227, n17228, n17229, n17230, n17231, n17232, n17233, n17234, n17236,
    n17237, n17238, n17239, n17240, n17241, n17242, n17243, n17244, n17245,
    n17246, n17247, n17248, n17249, n17250, n17251, n17252, n17253, n17254,
    n17255, n17257, n17258, n17259, n17260, n17261, n17262, n17263, n17264,
    n17265, n17266, n17267, n17268, n17269, n17270, n17271, n17272, n17273,
    n17275, n17276, n17277, n17278, n17279, n17280, n17281, n17282, n17283,
    n17284, n17285, n17286, n17287, n17288, n17289, n17290, n17291, n17292,
    n17293, n17294, n17295, n17296, n17297, n17298, n17299, n17300, n17301,
    n17302, n17303, n17304, n17305, n17306, n17307, n17308, n17309, n17310,
    n17311, n17312, n17313, n17314, n17315, n17316, n17317, n17318, n17319,
    n17320, n17321, n17322, n17323, n17324, n17325, n17326, n17327, n17328,
    n17329, n17330, n17331, n17332, n17333, n17334, n17335, n17336, n17337,
    n17338, n17339, n17340, n17341, n17342, n17343, n17344, n17345, n17346,
    n17347, n17348, n17349, n17350, n17351, n17352, n17353, n17354, n17355,
    n17356, n17357, n17358, n17359, n17360, n17361, n17362, n17363, n17364,
    n17365, n17366, n17367, n17368, n17369, n17370, n17371, n17372, n17373,
    n17374, n17375, n17376, n17377, n17378, n17379, n17380, n17381, n17382,
    n17383, n17384, n17385, n17386, n17387, n17388, n17389, n17390, n17391,
    n17392, n17393, n17394, n17395, n17396, n17397, n17398, n17399, n17400,
    n17401, n17402, n17403, n17404, n17405, n17406, n17407, n17408, n17409,
    n17410, n17411, n17412, n17413, n17414, n17415, n17416, n17417, n17418,
    n17419, n17420, n17421, n17422, n17423, n17424, n17425, n17426, n17427,
    n17428, n17429, n17430, n17431, n17432, n17433, n17434, n17435, n17436,
    n17437, n17438, n17439, n17440, n17441, n17442, n17443, n17444, n17445,
    n17446, n17447, n17448, n17449, n17450, n17451, n17453, n17454, n17455,
    n17456, n17457, n17458, n17459, n17460, n17461, n17462, n17463, n17464,
    n17465, n17466, n17467, n17468, n17469, n17470, n17471, n17472, n17474,
    n17475, n17476, n17477, n17478, n17479, n17480, n17481, n17482, n17483,
    n17484, n17485, n17486, n17487, n17488, n17489, n17490, n17491, n17492,
    n17493, n17495, n17496, n17497, n17498, n17499, n17500, n17501, n17502,
    n17503, n17504, n17505, n17506, n17507, n17508, n17509, n17510, n17511,
    n17513, n17514, n17515, n17516, n17517, n17518, n17519, n17520, n17521,
    n17522, n17523, n17524, n17525, n17526, n17527, n17528, n17529, n17530,
    n17531, n17532, n17534, n17535, n17536, n17537, n17538, n17539, n17540,
    n17541, n17542, n17543, n17544, n17545, n17546, n17547, n17548, n17549,
    n17550, n17552, n17553, n17554, n17555, n17556, n17557, n17558, n17559,
    n17560, n17561, n17562, n17563, n17564, n17565, n17566, n17567, n17568,
    n17569, n17570, n17571, n17573, n17574, n17575, n17576, n17577, n17578,
    n17579, n17580, n17581, n17582, n17583, n17584, n17585, n17586, n17587,
    n17588, n17589, n17591, n17592, n17593, n17594, n17595, n17596, n17597,
    n17598, n17599, n17600, n17601, n17602, n17603, n17604, n17605, n17606,
    n17607, n17608, n17609, n17610, n17611, n17612, n17613, n17614, n17615,
    n17616, n17617, n17618, n17619, n17620, n17621, n17622, n17623, n17624,
    n17625, n17626, n17627, n17628, n17629, n17630, n17631, n17632, n17633,
    n17634, n17635, n17636, n17637, n17638, n17639, n17640, n17641, n17642,
    n17643, n17644, n17645, n17646, n17647, n17648, n17649, n17650, n17651,
    n17652, n17653, n17654, n17655, n17656, n17657, n17658, n17659, n17660,
    n17661, n17662, n17663, n17664, n17665, n17666, n17667, n17668, n17669,
    n17670, n17671, n17672, n17673, n17674, n17675, n17676, n17677, n17678,
    n17679, n17680, n17681, n17682, n17683, n17684, n17685, n17686, n17687,
    n17688, n17689, n17690, n17691, n17692, n17693, n17694, n17695, n17696,
    n17697, n17698, n17699, n17700, n17701, n17702, n17703, n17704, n17705,
    n17706, n17707, n17708, n17709, n17710, n17711, n17712, n17713, n17714,
    n17715, n17716, n17717, n17718, n17719, n17720, n17721, n17722, n17723,
    n17724, n17725, n17726, n17727, n17728, n17729, n17730, n17731, n17732,
    n17733, n17734, n17735, n17736, n17737, n17738, n17739, n17740, n17741,
    n17742, n17743, n17744, n17745, n17746, n17747, n17748, n17749, n17750,
    n17751, n17752, n17753, n17754, n17755, n17756, n17757, n17758, n17759,
    n17760, n17761, n17762, n17763, n17764, n17765, n17766, n17767, n17768,
    n17769, n17770, n17771, n17772, n17773, n17774, n17775, n17776, n17777,
    n17778, n17779, n17780, n17781, n17782, n17783, n17784, n17785, n17787,
    n17788, n17789, n17790, n17791, n17793, n17794, n17795, n17796, n17797,
    n17798, n17799, n17800, n17802, n17803, n17804, n17805, n17806, n17807,
    n17808, n17809, n17810, n17811, n17812, n17813, n17814, n17815, n17817,
    n17818, n17819, n17820, n17821, n17822, n17823, n17824, n17825, n17826,
    n17827, n17828, n17829, n17830, n17831, n17832, n17833, n17834, n17835,
    n17836, n17837, n17838, n17839, n17840, n17841, n17842, n17843, n17844,
    n17845, n17846, n17847, n17848, n17849, n17850, n17851, n17852, n17853,
    n17854, n17855, n17856, n17857, n17858, n17859, n17860, n17861, n17862,
    n17863, n17864, n17865, n17866, n17867, n17868, n17869, n17870, n17871,
    n17872, n17873, n17874, n17875, n17876, n17877, n17878, n17879, n17880,
    n17881, n17882, n17883, n17884, n17885, n17886, n17887, n17888, n17889,
    n17890, n17891, n17892, n17893, n17894, n17895, n17896, n17897, n17898,
    n17899, n17900, n17901, n17902, n17903, n17904, n17905, n17906, n17907,
    n17908, n17909, n17910, n17911, n17912, n17913, n17914, n17915, n17916,
    n17917, n17918, n17919, n17920, n17921, n17922, n17923, n17924, n17925,
    n17926, n17927, n17928, n17929, n17930, n17931, n17932, n17933, n17934,
    n17935, n17936, n17937, n17938, n17939, n17940, n17941, n17942, n17943,
    n17944, n17945, n17946, n17947, n17948, n17949, n17950, n17951, n17952,
    n17954, n17955, n17956, n17957, n17958, n17959, n17960, n17961, n17962,
    n17963, n17964, n17965, n17966, n17967, n17968, n17969, n17970, n17971,
    n17972, n17973, n17974, n17975, n17976, n17977, n17978, n17979, n17980,
    n17981, n17982, n17983, n17984, n17985, n17986, n17987, n17988, n17989,
    n17990, n17991, n17992, n17993, n17994, n17995, n17996, n17997, n17998,
    n17999, n18000, n18001, n18002, n18003, n18004, n18005, n18006, n18007,
    n18008, n18009, n18010, n18011, n18012, n18013, n18014, n18015, n18016,
    n18017, n18018, n18019, n18020, n18021, n18022, n18023, n18024, n18025,
    n18026, n18027, n18028, n18029, n18030, n18031, n18032, n18033, n18034,
    n18035, n18036, n18037, n18038, n18039, n18040, n18041, n18042, n18043,
    n18044, n18045, n18046, n18047, n18048, n18049, n18050, n18051, n18052,
    n18053, n18054, n18055, n18056, n18057, n18058, n18059, n18060, n18061,
    n18062, n18063, n18064, n18065, n18066, n18067, n18068, n18069, n18070,
    n18071, n18072, n18073, n18074, n18075, n18076, n18077, n18079, n18080,
    n18081, n18082, n18083, n18084, n18085, n18086, n18087, n18088, n18089,
    n18091, n18092, n18093, n18094, n18095, n18096, n18097, n18098, n18099,
    n18100, n18101, n18102, n18103, n18104, n18106, n18107, n18108, n18109,
    n18110, n18111, n18112, n18113, n18114, n18115, n18116, n18117, n18118,
    n18119, n18120, n18121, n18122, n18123, n18124, n18125, n18126, n18127,
    n18128, n18129, n18130, n18131, n18132, n18133, n18134, n18135, n18136,
    n18137, n18138, n18139, n18140, n18141, n18142, n18143, n18144, n18145,
    n18146, n18147, n18148, n18149, n18150, n18151, n18152, n18153, n18154,
    n18155, n18156, n18157, n18158, n18159, n18160, n18161, n18162, n18163,
    n18164, n18165, n18166, n18167, n18168, n18169, n18170, n18171, n18172,
    n18173, n18174, n18175, n18176, n18177, n18178, n18179, n18180, n18181,
    n18182, n18183, n18184, n18185, n18186, n18187, n18188, n18189, n18190,
    n18191, n18192, n18193, n18194, n18195, n18196, n18197, n18198, n18199,
    n18200, n18201, n18202, n18203, n18204, n18205, n18206, n18207, n18208,
    n18209, n18210, n18211, n18212, n18213, n18214, n18215, n18216, n18217,
    n18218, n18219, n18220, n18221, n18222, n18223, n18224, n18225, n18226,
    n18227, n18228, n18229, n18230, n18231, n18232, n18233, n18234, n18235,
    n18236, n18237, n18238, n18239, n18240, n18241, n18242, n18243, n18244,
    n18245, n18246, n18247, n18248, n18249, n18250, n18251, n18252, n18253,
    n18254, n18255, n18256, n18257, n18258, n18259, n18260, n18261, n18262,
    n18263, n18264, n18265, n18266, n18267, n18268, n18269, n18270, n18271,
    n18272, n18273, n18274, n18275, n18276, n18277, n18278, n18279, n18280,
    n18281, n18282, n18284, n18285, n18286, n18287, n18288, n18289, n18290,
    n18291, n18292, n18293, n18294, n18295, n18296, n18297, n18299, n18300,
    n18301, n18302, n18303, n18304, n18305, n18306, n18307, n18308, n18309,
    n18310, n18311, n18312, n18313, n18314, n18315, n18316, n18317, n18318,
    n18319, n18320, n18321, n18322, n18323, n18324, n18325, n18326, n18327,
    n18328, n18329, n18330, n18331, n18332, n18333, n18334, n18335, n18336,
    n18337, n18338, n18339, n18340, n18341, n18342, n18343, n18344, n18345,
    n18346, n18347, n18348, n18349, n18350, n18351, n18352, n18353, n18354,
    n18355, n18356, n18357, n18358, n18359, n18360, n18361, n18362, n18363,
    n18364, n18365, n18366, n18367, n18368, n18369, n18370, n18371, n18372,
    n18373, n18374, n18375, n18376, n18377, n18378, n18379, n18380, n18381,
    n18382, n18383, n18384, n18385, n18386, n18387, n18388, n18389, n18390,
    n18391, n18392, n18393, n18394, n18395, n18396, n18397, n18398, n18399,
    n18400, n18401, n18402, n18403, n18404, n18405, n18406, n18407, n18408,
    n18409, n18410, n18411, n18412, n18413, n18414, n18416, n18417, n18418,
    n18419, n18420, n18421, n18422, n18423, n18424, n18425, n18426, n18427,
    n18428, n18429, n18431, n18432, n18433, n18434, n18435, n18436, n18437,
    n18438, n18440, n18441, n18442, n18443, n18444, n18445, n18446, n18447,
    n18448, n18449, n18450, n18451, n18452, n18453, n18454, n18455, n18456,
    n18457, n18458, n18459, n18460, n18461, n18462, n18463, n18464, n18465,
    n18466, n18467, n18468, n18469, n18470, n18471, n18472, n18473, n18474,
    n18475, n18476, n18477, n18478, n18479, n18480, n18481, n18482, n18483,
    n18484, n18485, n18486, n18487, n18488, n18489, n18490, n18491, n18492,
    n18493, n18494, n18495, n18496, n18497, n18498, n18499, n18500, n18501,
    n18502, n18503, n18504, n18505, n18506, n18507, n18508, n18509, n18510,
    n18511, n18512, n18513, n18514, n18515, n18516, n18517, n18518, n18519,
    n18520, n18521, n18522, n18523, n18524, n18525, n18526, n18527, n18528,
    n18529, n18530, n18531, n18532, n18533, n18534, n18535, n18536, n18537,
    n18538, n18539, n18540, n18541, n18542, n18543, n18544, n18545, n18546,
    n18547, n18548, n18549, n18550, n18551, n18552, n18553, n18554, n18555,
    n18556, n18557, n18558, n18559, n18560, n18561, n18562, n18563, n18564,
    n18565, n18566, n18567, n18568, n18569, n18570, n18571, n18572, n18573,
    n18574, n18575, n18576, n18577, n18578, n18579, n18580, n18581, n18582,
    n18583, n18584, n18585, n18586, n18587, n18588, n18589, n18590, n18591,
    n18592, n18593, n18594, n18595, n18596, n18597, n18598, n18599, n18600,
    n18601, n18602, n18603, n18604, n18605, n18606, n18607, n18608, n18609,
    n18610, n18611, n18612, n18613, n18614, n18615, n18616, n18617, n18618,
    n18619, n18620, n18621, n18622, n18623, n18624, n18625, n18627, n18628,
    n18629, n18630, n18631, n18632, n18633, n18634, n18635, n18636, n18637,
    n18638, n18639, n18640, n18641, n18642, n18643, n18644, n18645, n18646,
    n18647, n18648, n18649, n18650, n18651, n18652, n18653, n18654, n18655,
    n18656, n18657, n18658, n18659, n18660, n18661, n18662, n18663, n18664,
    n18665, n18666, n18667, n18668, n18669, n18670, n18671, n18672, n18673,
    n18674, n18675, n18676, n18677, n18678, n18679, n18680, n18681, n18682,
    n18683, n18684, n18685, n18686, n18687, n18688, n18689, n18690, n18691,
    n18692, n18693, n18694, n18695, n18696, n18697, n18698, n18699, n18700,
    n18701, n18702, n18703, n18704, n18705, n18706, n18707, n18708, n18709,
    n18710, n18711, n18712, n18713, n18714, n18715, n18716, n18717, n18718,
    n18719, n18720, n18721, n18722, n18723, n18724, n18725, n18726, n18727,
    n18728, n18729, n18730, n18731, n18732, n18733, n18734, n18735, n18736,
    n18737, n18738, n18739, n18740, n18741, n18742, n18743, n18744, n18745,
    n18746, n18747, n18748, n18749, n18750, n18751, n18752, n18753, n18755,
    n18756, n18757, n18758, n18759, n18761, n18762, n18763, n18764, n18765,
    n18766, n18767, n18768, n18769, n18770, n18771, n18772, n18773, n18774,
    n18775, n18776, n18777, n18778, n18779, n18780, n18781, n18782, n18783,
    n18784, n18785, n18786, n18787, n18788, n18789, n18790, n18791, n18792,
    n18793, n18794, n18795, n18796, n18797, n18798, n18799, n18800, n18801,
    n18802, n18803, n18804, n18805, n18806, n18807, n18808, n18809, n18810,
    n18811, n18812, n18813, n18814, n18815, n18816, n18817, n18818, n18819,
    n18820, n18821, n18822, n18823, n18824, n18825, n18826, n18827, n18828,
    n18829, n18830, n18831, n18832, n18833, n18834, n18835, n18836, n18837,
    n18838, n18839, n18840, n18841, n18842, n18843, n18844, n18845, n18846,
    n18847, n18848, n18849, n18850, n18851, n18852, n18853, n18854, n18855,
    n18856, n18857, n18858, n18859, n18861, n18862, n18863, n18864, n18865,
    n18866, n18867, n18868, n18869, n18870, n18871, n18873, n18874, n18875,
    n18876, n18877, n18878, n18879, n18880, n18881, n18882, n18883, n18884,
    n18885, n18886, n18888, n18889, n18890, n18891, n18892, n18894, n18895,
    n18896, n18897, n18898, n18899, n18900, n18901, n18903, n18904, n18905,
    n18906, n18907, n18908, n18909, n18910, n18911, n18912, n18913, n18914,
    n18915, n18916, n18917, n18918, n18919, n18920, n18921, n18922, n18923,
    n18924, n18925, n18926, n18927, n18928, n18929, n18930, n18931, n18932,
    n18933, n18934, n18935, n18936, n18937, n18938, n18939, n18940, n18941,
    n18942, n18943, n18944, n18945, n18946, n18947, n18948, n18949, n18950,
    n18951, n18952, n18953, n18954, n18955, n18956, n18957, n18958, n18959,
    n18960, n18961, n18962, n18963, n18964, n18965, n18966, n18967, n18968,
    n18969, n18970, n18971, n18972, n18973, n18974, n18975, n18976, n18977,
    n18978, n18979, n18980, n18981, n18982, n18983, n18984, n18985, n18986,
    n18987, n18988, n18989, n18990, n18991, n18992, n18993, n18994, n18995,
    n18996, n18997, n18998, n18999, n19000, n19001, n19002, n19003, n19004,
    n19005, n19006, n19007, n19008, n19009, n19010, n19011, n19012, n19014,
    n19015, n19016, n19017, n19018, n19019, n19020, n19021, n19022, n19023,
    n19024, n19025, n19026, n19027, n19028, n19029, n19030, n19031, n19032,
    n19033, n19034, n19035, n19036, n19037, n19038, n19039, n19040, n19041,
    n19042, n19043, n19044, n19045, n19046, n19047, n19048, n19049, n19050,
    n19051, n19052, n19053, n19054, n19055, n19056, n19057, n19058, n19059,
    n19060, n19061, n19062, n19063, n19064, n19065, n19066, n19067, n19068,
    n19069, n19070, n19071, n19072, n19073, n19074, n19075, n19076, n19077,
    n19078, n19079, n19080, n19081, n19082, n19083, n19084, n19085, n19086,
    n19087, n19088, n19089, n19090, n19091, n19092, n19093, n19094, n19095,
    n19096, n19097, n19098, n19099, n19100, n19101, n19102, n19103, n19104,
    n19105, n19106, n19107, n19108, n19109, n19110, n19111, n19112, n19113,
    n19114, n19115, n19116, n19117, n19118, n19119, n19120, n19121, n19122,
    n19123, n19124, n19125, n19126, n19127, n19128, n19129, n19130, n19131,
    n19132, n19134, n19135, n19136, n19137, n19138, n19139, n19140, n19141,
    n19142, n19143, n19144, n19145, n19146, n19147, n19148, n19149, n19150,
    n19151, n19152, n19153, n19154, n19155, n19156, n19157, n19158, n19159,
    n19160, n19161, n19162, n19163, n19164, n19165, n19166, n19167, n19168,
    n19169, n19170, n19171, n19172, n19173, n19174, n19175, n19176, n19177,
    n19178, n19179, n19180, n19181, n19182, n19183, n19184, n19185, n19186,
    n19187, n19188, n19189, n19190, n19191, n19192, n19193, n19194, n19195,
    n19196, n19197, n19198, n19199, n19200, n19201, n19202, n19203, n19204,
    n19205, n19206, n19207, n19208, n19209, n19210, n19211, n19212, n19213,
    n19214, n19215, n19216, n19217, n19218, n19219, n19220, n19221, n19222,
    n19223, n19224, n19225, n19226, n19227, n19228, n19229, n19230, n19231,
    n19232, n19233, n19234, n19235, n19236, n19237, n19238, n19239, n19240,
    n19241, n19242, n19243, n19244, n19245, n19246, n19247, n19248, n19249,
    n19251, n19252, n19253, n19254, n19255, n19256, n19257, n19258, n19259,
    n19260, n19261, n19262, n19263, n19264, n19266, n19267, n19268, n19269,
    n19270, n19271, n19272, n19273, n19274, n19275, n19276, n19277, n19278,
    n19279, n19280, n19281, n19282, n19283, n19284, n19285, n19286, n19287,
    n19288, n19289, n19290, n19291, n19292, n19293, n19294, n19295, n19296,
    n19297, n19298, n19299, n19300, n19301, n19302, n19303, n19304, n19305,
    n19306, n19307, n19308, n19309, n19310, n19311, n19312, n19313, n19314,
    n19315, n19316, n19317, n19318, n19319, n19320, n19321, n19322, n19323,
    n19324, n19325, n19326, n19327, n19328, n19329, n19330, n19331, n19332,
    n19333, n19334, n19335, n19336, n19337, n19338, n19339, n19340, n19341,
    n19342, n19343, n19344, n19345, n19346, n19347, n19348, n19349, n19350,
    n19351, n19352, n19353, n19354, n19355, n19356, n19357, n19358, n19359,
    n19360, n19361, n19362, n19363, n19364, n19365, n19366, n19367, n19368,
    n19369, n19370, n19371, n19372, n19373, n19374, n19375, n19377, n19378,
    n19379, n19380, n19381, n19382, n19383, n19384, n19385, n19386, n19387,
    n19388, n19389, n19390, n19391, n19392, n19393, n19394, n19395, n19396,
    n19397, n19398, n19399, n19400, n19401, n19402, n19403, n19404, n19405,
    n19406, n19407, n19408, n19409, n19410, n19411, n19412, n19413, n19414,
    n19415, n19416, n19417, n19418, n19419, n19420, n19421, n19422, n19423,
    n19424, n19425, n19426, n19427, n19428, n19429, n19430, n19431, n19432,
    n19433, n19434, n19435, n19436, n19437, n19438, n19439, n19440, n19441,
    n19442, n19443, n19444, n19445, n19446, n19447, n19448, n19449, n19450,
    n19451, n19452, n19453, n19454, n19455, n19456, n19457, n19458, n19459,
    n19460, n19461, n19462, n19463, n19464, n19465, n19466, n19467, n19468,
    n19469, n19470, n19471, n19472, n19473, n19474, n19475, n19476, n19477,
    n19478, n19479, n19480, n19482, n19483, n19484, n19485, n19486, n19487,
    n19488, n19489, n19490, n19491, n19492, n19493, n19494, n19495, n19496,
    n19497, n19498, n19499, n19500, n19501, n19502, n19503, n19504, n19505,
    n19506, n19507, n19508, n19509, n19510, n19511, n19512, n19513, n19514,
    n19515, n19516, n19517, n19518, n19519, n19520, n19521, n19522, n19523,
    n19524, n19525, n19526, n19527, n19528, n19529, n19530, n19531, n19532,
    n19533, n19534, n19535, n19536, n19537, n19538, n19539, n19540, n19541,
    n19542, n19543, n19544, n19545, n19546, n19547, n19548, n19549, n19550,
    n19551, n19552, n19553, n19554, n19555, n19556, n19557, n19558, n19559,
    n19560, n19561, n19562, n19563, n19564, n19565, n19566, n19567, n19568,
    n19569, n19570, n19571, n19572, n19573, n19574, n19575, n19576, n19577,
    n19578, n19579, n19580, n19581, n19582, n19583, n19584, n19585, n19586,
    n19587, n19588, n19589, n19590, n19591, n19592, n19593, n19594, n19595,
    n19596, n19597, n19599, n19600, n19601, n19602, n19603, n19604, n19605,
    n19606, n19607, n19608, n19609, n19610, n19611, n19612, n19614, n19615,
    n19617, n19618, n19619, n19620, n19621, n19622, n19623, n19624, n19625,
    n19626, n19627, n19628, n19629, n19630, n19631, n19632, n19633, n19634,
    n19635, n19636, n19637, n19638, n19639, n19640, n19641, n19642, n19643,
    n19644, n19645, n19646, n19647, n19648, n19649, n19650, n19651, n19652,
    n19653, n19654, n19655, n19656, n19657, n19658, n19659, n19660, n19661,
    n19662, n19663, n19664, n19665, n19666, n19667, n19668, n19669, n19670,
    n19671, n19672, n19673, n19674, n19675, n19676, n19677, n19678, n19679,
    n19680, n19681, n19682, n19683, n19684, n19685, n19686, n19687, n19688,
    n19689, n19690, n19691, n19692, n19693, n19694, n19695, n19696, n19697,
    n19698, n19699, n19700, n19701, n19702, n19703, n19704, n19705, n19706,
    n19707, n19708, n19709, n19710, n19711, n19713, n19714, n19715, n19716,
    n19717, n19718, n19719, n19720, n19722, n19723, n19724, n19725, n19726,
    n19727, n19728, n19729, n19730, n19731, n19732, n19733, n19734, n19735,
    n19736, n19737, n19738, n19739, n19740, n19741, n19742, n19743, n19744,
    n19745, n19746, n19747, n19748, n19749, n19750, n19751, n19752, n19753,
    n19754, n19755, n19756, n19757, n19758, n19759, n19760, n19761, n19762,
    n19763, n19764, n19765, n19766, n19767, n19768, n19769, n19770, n19771,
    n19772, n19773, n19774, n19775, n19776, n19777, n19778, n19779, n19780,
    n19781, n19782, n19783, n19784, n19785, n19786, n19787, n19788, n19789,
    n19790, n19791, n19792, n19793, n19794, n19795, n19796, n19797, n19798,
    n19799, n19800, n19801, n19802, n19803, n19804, n19805, n19806, n19807,
    n19808, n19809, n19810, n19811, n19812, n19813, n19814, n19815, n19816,
    n19817, n19818, n19819, n19820, n19821, n19822, n19823, n19824, n19825,
    n19826, n19827, n19828, n19829, n19831, n19832, n19833, n19834, n19835,
    n19837, n19838, n19839, n19840, n19841, n19842, n19843, n19844, n19845,
    n19846, n19847, n19849, n19850, n19851, n19852, n19853, n19854, n19855,
    n19856, n19857, n19858, n19859, n19860, n19861, n19862, n19864, n19865,
    n19866, n19867, n19868, n19869, n19870, n19871, n19872, n19873, n19874,
    n19875, n19876, n19877, n19879, n19880, n19881, n19882, n19883, n19884,
    n19885, n19886, n19887, n19888, n19889, n19890, n19891, n19892, n19894,
    n19895, n19896, n19897, n19898, n19900, n19901, n19902, n19903, n19904,
    n19905, n19906, n19907, n19908, n19909, n19910, n19911, n19912, n19913,
    n19914, n19915, n19916, n19917, n19918, n19919, n19920, n19921, n19922,
    n19923, n19924, n19925, n19926, n19927, n19928, n19929, n19930, n19931,
    n19932, n19933, n19934, n19935, n19936, n19937, n19938, n19939, n19940,
    n19941, n19942, n19943, n19944, n19945, n19946, n19947, n19948, n19949,
    n19950, n19951, n19952, n19953, n19954, n19955, n19956, n19957, n19958,
    n19959, n19960, n19961, n19962, n19963, n19964, n19965, n19966, n19967,
    n19968, n19969, n19970, n19971, n19972, n19973, n19974, n19975, n19976,
    n19977, n19978, n19979, n19980, n19981, n19982, n19983, n19984, n19985,
    n19986, n19987, n19988, n19989, n19990, n19991, n19992, n19993, n19994,
    n19995, n19996, n19997, n19998, n19999, n20000, n20001, n20003, n20004,
    n20005, n20006, n20007, n20008, n20009, n20010, n20011, n20012, n20013,
    n20014, n20015, n20016, n20017, n20018, n20019, n20020, n20021, n20022,
    n20023, n20024, n20025, n20026, n20027, n20028, n20029, n20030, n20031,
    n20032, n20033, n20034, n20035, n20036, n20037, n20038, n20039, n20040,
    n20041, n20042, n20043, n20044, n20045, n20046, n20047, n20048, n20049,
    n20050, n20051, n20052, n20053, n20054, n20055, n20056, n20057, n20058,
    n20059, n20060, n20061, n20062, n20063, n20064, n20065, n20066, n20067,
    n20068, n20069, n20070, n20071, n20072, n20073, n20074, n20075, n20076,
    n20077, n20078, n20079, n20080, n20081, n20082, n20083, n20084, n20085,
    n20086, n20087, n20088, n20089, n20090, n20091, n20092, n20093, n20094,
    n20095, n20096, n20097, n20098, n20099, n20100, n20101, n20102, n20103,
    n20104, n20105, n20107, n20108, n20109, n20110, n20111, n20112, n20113,
    n20114, n20115, n20116, n20117, n20118, n20119, n20120, n20122, n20123,
    n20124, n20125, n20126, n20128, n20129, n20130, n20131, n20132, n20133,
    n20134, n20135, n20137, n20138, n20139, n20140, n20141, n20142, n20143,
    n20144, n20145, n20146, n20147, n20148, n20149, n20150, n20151, n20152,
    n20153, n20154, n20155, n20156, n20157, n20158, n20159, n20160, n20161,
    n20162, n20163, n20164, n20165, n20166, n20167, n20168, n20169, n20170,
    n20171, n20172, n20173, n20174, n20175, n20176, n20177, n20178, n20179,
    n20180, n20181, n20182, n20183, n20184, n20185, n20186, n20187, n20188,
    n20189, n20190, n20191, n20192, n20193, n20194, n20195, n20196, n20197,
    n20198, n20199, n20200, n20201, n20202, n20203, n20204, n20205, n20206,
    n20207, n20208, n20209, n20210, n20211, n20212, n20213, n20214, n20215,
    n20216, n20217, n20218, n20219, n20220, n20221, n20222, n20223, n20224,
    n20225, n20226, n20227, n20228, n20229, n20230, n20231, n20232, n20233,
    n20234, n20235, n20236, n20237, n20238, n20239, n20241, n20242, n20243,
    n20244, n20245, n20246, n20247, n20248, n20249, n20250, n20251, n20252,
    n20253, n20254, n20255, n20256, n20257, n20258, n20259, n20260, n20261,
    n20262, n20263, n20264, n20265, n20266, n20267, n20268, n20269, n20270,
    n20271, n20272, n20273, n20274, n20275, n20276, n20277, n20278, n20279,
    n20280, n20281, n20282, n20283, n20284, n20285, n20286, n20287, n20288,
    n20289, n20290, n20291, n20292, n20293, n20294, n20295, n20296, n20297,
    n20298, n20299, n20300, n20301, n20302, n20303, n20304, n20305, n20306,
    n20307, n20308, n20309, n20310, n20311, n20312, n20313, n20314, n20315,
    n20316, n20317, n20318, n20319, n20320, n20321, n20322, n20323, n20324,
    n20325, n20326, n20327, n20328, n20329, n20330, n20331, n20332, n20333,
    n20334, n20336, n20337, n20338, n20339, n20340, n20341, n20342, n20343,
    n20344, n20345, n20346, n20347, n20348, n20349, n20351, n20352, n20354,
    n20355, n20357, n20358, n20359, n20360, n20361, n20362, n20363, n20364,
    n20366, n20367, n20368, n20369, n20370, n20371, n20372, n20373, n20374,
    n20375, n20376, n20377, n20378, n20379, n20380, n20381, n20382, n20383,
    n20384, n20385, n20386, n20387, n20388, n20389, n20390, n20391, n20392,
    n20393, n20394, n20395, n20396, n20397, n20398, n20399, n20400, n20401,
    n20402, n20403, n20404, n20405, n20406, n20407, n20408, n20409, n20410,
    n20411, n20412, n20413, n20414, n20415, n20416, n20417, n20418, n20419,
    n20420, n20421, n20422, n20423, n20424, n20425, n20426, n20427, n20428,
    n20429, n20430, n20431, n20432, n20433, n20434, n20435, n20436, n20437,
    n20438, n20439, n20440, n20441, n20442, n20443, n20444, n20445, n20446,
    n20447, n20448, n20449, n20450, n20451, n20452, n20453, n20454, n20455,
    n20456, n20458, n20459, n20460, n20461, n20462, n20463, n20464, n20465,
    n20467, n20468, n20469, n20470, n20471, n20473, n20474, n20475, n20476,
    n20477, n20478, n20479, n20480, n20481, n20482, n20483, n20484, n20485,
    n20486, n20488, n20489, n20490, n20491, n20492, n20493, n20494, n20495,
    n20496, n20497, n20498, n20499, n20500, n20501, n20502, n20503, n20504,
    n20505, n20506, n20507, n20508, n20509, n20510, n20511, n20512, n20513,
    n20514, n20515, n20516, n20517, n20518, n20519, n20520, n20521, n20522,
    n20523, n20524, n20525, n20526, n20527, n20528, n20529, n20530, n20531,
    n20532, n20533, n20534, n20535, n20536, n20537, n20538, n20539, n20540,
    n20541, n20542, n20543, n20544, n20545, n20546, n20547, n20548, n20549,
    n20550, n20551, n20552, n20553, n20554, n20555, n20556, n20557, n20558,
    n20559, n20560, n20561, n20562, n20563, n20564, n20565, n20566, n20567,
    n20568, n20569, n20570, n20571, n20572, n20573, n20574, n20575, n20576,
    n20577, n20578, n20579, n20580, n20581, n20582, n20583, n20584, n20585,
    n20586, n20587, n20588, n20589, n20590, n20592, n20593, n20594, n20595,
    n20596, n20597, n20598, n20599, n20600, n20601, n20602, n20603, n20604,
    n20605, n20606, n20607, n20608, n20609, n20610, n20611, n20612, n20613,
    n20614, n20615, n20616, n20617, n20618, n20619, n20620, n20621, n20622,
    n20623, n20624, n20625, n20626, n20627, n20628, n20629, n20630, n20631,
    n20632, n20633, n20634, n20635, n20636, n20637, n20638, n20639, n20640,
    n20641, n20642, n20643, n20644, n20645, n20646, n20647, n20648, n20649,
    n20650, n20651, n20652, n20653, n20654, n20655, n20656, n20657, n20658,
    n20659, n20660, n20661, n20662, n20663, n20664, n20665, n20666, n20667,
    n20668, n20669, n20670, n20671, n20672, n20673, n20674, n20675, n20676,
    n20677, n20678, n20679, n20680, n20681, n20682, n20683, n20684, n20685,
    n20686, n20688, n20689, n20690, n20691, n20692, n20693, n20694, n20695,
    n20696, n20697, n20698, n20699, n20700, n20701, n20703, n20704, n20706,
    n20707, n20708, n20709, n20710, n20712, n20713, n20715, n20716, n20717,
    n20718, n20719, n20721, n20722, n20723, n20724, n20725, n20726, n20727,
    n20728, n20730, n20731, n20732, n20733, n20734, n20735, n20736, n20737,
    n20738, n20739, n20740, n20741, n20742, n20743, n20745, n20746, n20747,
    n20748, n20749, n20750, n20751, n20752, n20754, n20755, n20756, n20757,
    n20758, n20759, n20760, n20761, n20762, n20763, n20764, n20765, n20766,
    n20767, n20769, n20770, n20772, n20773, n20775, n20776, n20778, n20779,
    n20781, n20782, n20784, n20785, n20787, n20788, n20790, n20791, n20793,
    n20794, n20796, n20797, n20799, n20800, n20802, n20803, n20805, n20806,
    n20808, n20809, n20810, n20811, n20812, n20813, n20814, n20815, n20816,
    n20817, n20818, n20819, n20820, n20821, n20822, n20823, n20824, n20825,
    n20826, n20827, n20828, n20829, n20830, n20831, n20832, n20833, n20834,
    n20835, n20836, n20837, n20838, n20839, n20840, n20841, n20842, n20843,
    n20844, n20845, n20846, n20847, n20848, n20849, n20850, n20851, n20852,
    n20853, n20854, n20855, n20856, n20857, n20858, n20859, n20860, n20861,
    n20862, n20863, n20864, n20865, n20866, n20867, n20868, n20869, n20870,
    n20871, n20872, n20873, n20874, n20875, n20876, n20877, n20878, n20879,
    n20880, n20881, n20882, n20883, n20884, n20885, n20886, n20887, n20888,
    n20889, n20890, n20891, n20892, n20893, n20894, n20895, n20896, n20897,
    n20898, n20899, n20900, n20901, n20902, n20903, n20904, n20905, n20906,
    n20908, n20909, n20910, n20911, n20912, n20913, n20914, n20915, n20917,
    n20918, n20919, n20920, n20921, n20922, n20923, n20924, n20925, n20926,
    n20927, n20928, n20929, n20930, n20932, n20933, n20934, n20935, n20936,
    n20937, n20938, n20939, n20941, n20942, n20944, n20945, n20947, n20948,
    n20950, n20951, n20953, n20954, n20955, n20956, n20957, n20958, n20959,
    n20960, n20961, n20962, n20963, n20964, n20965, n20966, n20968, n20969,
    n20971, n20972, n20973, n20974, n20975, n20976, n20977, n20978, n20979,
    n20980, n20981, n20982, n20983, n20984, n20985, n20986, n20987, n20988,
    n20989, n20990, n20991, n20992, n20993, n20994, n20995, n20996, n20997,
    n20998, n20999, n21000, n21001, n21002, n21003, n21004, n21005, n21006,
    n21007, n21008, n21009, n21010, n21011, n21012, n21013, n21014, n21015,
    n21016, n21017, n21018, n21019, n21020, n21021, n21022, n21023, n21024,
    n21025, n21026, n21027, n21028, n21029, n21030, n21031, n21032, n21033,
    n21034, n21035, n21036, n21037, n21038, n21039, n21040, n21041, n21042,
    n21043, n21044, n21045, n21046, n21047, n21048, n21049, n21050, n21051,
    n21052, n21053, n21054, n21055, n21056, n21057, n21058, n21059, n21060,
    n21061, n21062, n21063, n21065, n21066, n21067, n21068, n21069, n21070,
    n21071, n21072, n21073, n21074, n21075, n21076, n21077, n21078, n21079,
    n21080, n21081, n21082, n21083, n21084, n21085, n21086, n21087, n21088,
    n21089, n21090, n21091, n21092, n21093, n21094, n21095, n21096, n21097,
    n21098, n21099, n21100, n21101, n21102, n21103, n21104, n21105, n21106,
    n21107, n21108, n21109, n21110, n21111, n21112, n21113, n21114, n21115,
    n21116, n21117, n21118, n21119, n21120, n21121, n21122, n21123, n21124,
    n21125, n21126, n21127, n21128, n21129, n21130, n21131, n21132, n21133,
    n21134, n21135, n21136, n21137, n21138, n21139, n21140, n21141, n21142,
    n21143, n21144, n21145, n21146, n21147, n21148, n21149, n21150, n21151,
    n21152, n21153, n21154, n21155, n21156, n21157, n21159, n21160, n21161,
    n21162, n21163, n21164, n21165, n21166, n21167, n21168, n21169, n21170,
    n21171, n21172, n21173, n21174, n21175, n21176, n21177, n21178, n21179,
    n21180, n21181, n21182, n21183, n21184, n21185, n21186, n21187, n21188,
    n21189, n21190, n21191, n21192, n21193, n21194, n21195, n21196, n21197,
    n21198, n21199, n21200, n21201, n21202, n21203, n21204, n21205, n21206,
    n21207, n21208, n21209, n21210, n21211, n21212, n21213, n21214, n21215,
    n21216, n21217, n21218, n21219, n21220, n21221, n21222, n21223, n21224,
    n21225, n21226, n21227, n21228, n21229, n21230, n21231, n21232, n21233,
    n21234, n21235, n21236, n21237, n21238, n21239, n21240, n21241, n21242,
    n21243, n21244, n21245, n21246, n21247, n21248, n21249, n21250, n21251,
    n21252, n21253, n21254, n21255, n21256, n21257, n21258, n21259, n21260,
    n21261, n21263, n21264, n21265, n21266, n21267, n21268, n21269, n21270,
    n21271, n21272, n21273, n21274, n21275, n21276, n21277, n21278, n21279,
    n21280, n21281, n21282, n21283, n21284, n21285, n21286, n21287, n21288,
    n21289, n21290, n21291, n21292, n21293, n21294, n21295, n21296, n21297,
    n21298, n21299, n21300, n21301, n21302, n21303, n21304, n21305, n21306,
    n21307, n21308, n21309, n21310, n21311, n21312, n21313, n21314, n21315,
    n21316, n21317, n21318, n21319, n21320, n21321, n21322, n21323, n21324,
    n21325, n21326, n21327, n21328, n21329, n21330, n21331, n21332, n21333,
    n21334, n21335, n21336, n21337, n21338, n21339, n21340, n21341, n21342,
    n21343, n21344, n21345, n21346, n21347, n21348, n21349, n21350, n21351,
    n21352, n21353, n21354, n21356, n21357, n21358, n21359, n21360, n21361,
    n21362, n21363, n21364, n21365, n21366, n21367, n21368, n21369, n21371,
    n21372, n21373, n21374, n21375, n21377, n21378, n21379, n21380, n21381,
    n21383, n21384, n21385, n21386, n21387, n21389, n21390, n21391, n21392,
    n21393, n21395, n21396, n21397, n21398, n21399, n21400, n21401, n21402,
    n21404, n21405, n21406, n21407, n21408, n21409, n21410, n21411, n21413,
    n21414, n21415, n21416, n21417, n21418, n21419, n21420, n21422, n21423,
    n21424, n21425, n21426, n21427, n21428, n21429, n21431, n21432, n21433,
    n21434, n21435, n21436, n21437, n21438, n21440, n21441, n21442, n21443,
    n21444, n21445, n21446, n21447, n21448, n21449, n21450, n21451, n21452,
    n21453, n21455, n21456, n21457, n21458, n21459, n21460, n21461, n21462,
    n21463, n21464, n21465, n21466, n21467, n21468, n21470, n21471, n21472,
    n21473, n21474, n21475, n21476, n21477, n21478, n21479, n21480, n21481,
    n21482, n21483, n21485, n21486, n21487, n21488, n21489, n21490, n21491,
    n21492, n21493, n21494, n21495, n21496, n21497, n21498, n21500, n21501,
    n21503, n21504, n21506, n21507, n21509, n21510, n21512, n21513, n21515,
    n21516, n21518, n21519, n21521, n21522, n21524, n21525, n21527, n21528,
    n21530, n21531, n21533, n21534, n21536, n21537, n21539, n21540, n21542,
    n21543, n21545, n21546, n21548, n21549, n21551, n21552, n21554, n21555,
    n21557, n21558, n21560, n21561, n21562, n21563, n21564, n21565, n21566,
    n21567, n21569, n21570, n21571, n21572, n21573, n21575, n21576, n21577,
    n21578, n21579, n21580, n21581, n21582, n21583, n21584, n21585, n21586,
    n21587, n21588, n21589, n21590, n21591, n21592, n21593, n21594, n21595,
    n21596, n21597, n21598, n21599, n21600, n21601, n21602, n21603, n21604,
    n21605, n21606, n21607, n21608, n21609, n21610, n21611, n21612, n21613,
    n21614, n21615, n21616, n21617, n21618, n21619, n21620, n21621, n21622,
    n21623, n21624, n21625, n21626, n21627, n21628, n21629, n21630, n21631,
    n21632, n21633, n21634, n21635, n21636, n21637, n21638, n21639, n21640,
    n21641, n21642, n21643, n21644, n21645, n21646, n21647, n21648, n21649,
    n21650, n21651, n21652, n21653, n21654, n21655, n21656, n21657, n21658,
    n21659, n21660, n21661, n21662, n21663, n21664, n21665, n21666, n21667,
    n21668, n21669, n21670, n21672, n21673, n21674, n21675, n21676, n21677,
    n21678, n21679, n21680, n21681, n21682, n21683, n21684, n21685, n21686,
    n21687, n21688, n21689, n21690, n21691, n21692, n21693, n21694, n21695,
    n21696, n21697, n21698, n21699, n21700, n21701, n21702, n21703, n21704,
    n21705, n21706, n21707, n21708, n21709, n21710, n21711, n21712, n21713,
    n21714, n21715, n21716, n21717, n21718, n21719, n21720, n21721, n21722,
    n21723, n21724, n21725, n21726, n21727, n21728, n21729, n21730, n21731,
    n21732, n21733, n21734, n21735, n21736, n21737, n21738, n21739, n21740,
    n21741, n21742, n21743, n21744, n21745, n21746, n21747, n21748, n21749,
    n21750, n21751, n21752, n21753, n21754, n21755, n21756, n21757, n21758,
    n21759, n21760, n21761, n21762, n21763, n21764, n21765, n21766, n21767,
    n21768, n21769, n21770, n21771, n21773, n21774, n21776, n21777, n21779,
    n21780, n21782, n21783, n21785, n21786, n21788, n21789, n21791, n21792,
    n21794, n21795, n21797, n21798, n21799, n21800, n21801, n21802, n21803,
    n21804, n21805, n21806, n21807, n21808, n21809, n21810, n21811, n21812,
    n21813, n21814, n21815, n21816, n21817, n21818, n21819, n21820, n21821,
    n21822, n21823, n21824, n21825, n21826, n21827, n21828, n21829, n21830,
    n21831, n21832, n21833, n21834, n21835, n21836, n21837, n21838, n21839,
    n21840, n21841, n21842, n21843, n21844, n21845, n21846, n21847, n21848,
    n21849, n21850, n21851, n21852, n21853, n21854, n21855, n21856, n21857,
    n21858, n21859, n21860, n21861, n21862, n21863, n21864, n21865, n21866,
    n21867, n21868, n21869, n21870, n21871, n21872, n21873, n21874, n21875,
    n21876, n21877, n21878, n21879, n21880, n21881, n21882, n21883, n21884,
    n21885, n21886, n21887, n21888, n21889, n21890, n21891, n21892, n21894,
    n21895, n21896, n21897, n21898, n21899, n21900, n21901, n21902, n21903,
    n21904, n21906, n21907, n21908, n21909, n21910, n21912, n21913, n21914,
    n21915, n21916, n21917, n21918, n21919, n21920, n21921, n21922, n21923,
    n21924, n21925, n21927, n21928, n21929, n21930, n21931, n21933, n21934,
    n21935, n21936, n21937, n21939, n21940, n21941, n21942, n21943, n21944,
    n21945, n21946, n21948, n21949, n21950, n21951, n21952, n21953, n21954,
    n21955, n21957, n21958, n21959, n21960, n21961, n21962, n21963, n21964,
    n21965, n21966, n21967, n21968, n21969, n21970, n21972, n21973, n21974,
    n21975, n21976, n21977, n21978, n21979, n21980, n21981, n21982, n21983,
    n21984, n21985, n21987, n21988, n21990, n21991, n21992, n21993, n21994,
    n21996, n21997, n21999, n22000, n22001, n22002, n22003, n22005, n22006,
    n22007, n22008, n22009, n22010, n22011, n22012, n22014, n22015, n22017,
    n22018, n22019, n22020, n22021, n22022, n22023, n22024, n22026, n22027,
    n22028, n22029, n22030, n22031, n22032, n22033, n22034, n22035, n22036,
    n22037, n22038, n22039, n22041, n22042, n22043, n22044, n22045, n22046,
    n22047, n22048, n22049, n22050, n22051, n22052, n22053, n22054, n22056,
    n22057, n22059, n22060, n22062, n22063, n22065, n22066, n22068, n22069,
    n22071, n22072, n22074, n22075, n22077, n22078, n22080, n22081, n22083,
    n22084, n22086, n22087, n22089, n22090, n22092, n22093, n22095, n22096,
    n22098, n22099, n22101, n22102, n22103, n22104, n22105, n22106, n22107,
    n22108, n22110, n22111, n22112, n22113, n22114, n22115, n22116, n22117,
    n22118, n22119, n22120, n22121, n22122, n22123, n22125, n22126, n22127,
    n22128, n22129, n22130, n22131, n22132, n22134, n22135, n22137, n22138,
    n22140, n22141, n22143, n22144, n22146, n22147, n22149, n22150, n22152,
    n22153, n22155, n22156, n22158, n22159, n22161, n22162, n22164, n22165,
    n22167, n22168, n22170, n22171, n22173, n22174, n22176, n22177, n22179,
    n22180, n22181, n22182, n22183, n22185, n22186, n22187, n22188, n22189,
    n22190, n22191, n22192, n22194, n22195, n22196, n22197, n22198, n22199,
    n22200, n22201, n22202, n22203, n22204, n22205, n22206, n22207, n22209,
    n22210, n22212, n22213, n22215, n22216, n22218, n22219, n22221, n22222,
    n22224, n22225, n22227, n22228, n22230, n22231, n22233, n22234, n22236,
    n22237, n22239, n22240, n22242, n22243, n22245, n22246, n22248, n22249,
    n22251, n22252, n22254, n22255, n22257, n22258, n22260, n22261, n22263,
    n22264, n22266, n22267, n22269, n22270, n22271, n22272, n22273, n22274,
    n22275, n22276, n22277, n22278, n22279, n22280, n22281, n22282, n22284,
    n22285, n22287, n22288, n22290, n22291, n22293, n22294, n22295, n22296,
    n22297, n22298, n22299, n22300, n22302, n22303, n22305, n22306, n22307,
    n22308, n22309, n22310, n22311, n22312, n22314, n22315, n22316, n22317,
    n22318, n22320, n22321, n22322, n22323, n22324, n22325, n22326, n22327,
    n22329, n22330, n22331, n22332, n22333, n22334, n22335, n22336, n22337,
    n22338, n22339, n22340, n22341, n22342, n22344, n22345, n22346, n22347,
    n22348, n22349, n22350, n22351, n22352, n22353, n22354, n22355, n22356,
    n22357, n22359, n22360, n22361, n22362, n22363, n22365, n22366, n22367,
    n22368, n22369, n22370, n22371, n22372, n22373, n22374, n22375, n22376,
    n22377, n22378, n22380, n22381, n22383, n22384, n22385, n22386, n22387,
    n22389, n22390, n22391, n22392, n22393, n22394, n22395, n22396, n22398,
    n22399, n22400, n22401, n22402, n22403, n22404, n22405, n22406, n22407,
    n22408, n22409, n22410, n22411, n22413, n22414, n22416, n22417, n22419,
    n22420, n22422, n22423, n22425, n22426, n22428, n22429, n22431, n22432,
    n22434, n22435, n22437, n22438, n22440, n22441, n22443, n22444, n22446,
    n22447, n22448, n22449, n22450, n22452, n22453, n22454, n22455, n22456,
    n22458, n22459, n22460, n22461, n22462, n22463, n22464, n22465, n22466,
    n22467, n22468, n22469, n22470, n22471, n22473, n22474, n22475, n22476,
    n22477, n22478, n22479, n22480, n22482, n22483, n22485, n22486, n22487,
    n22488, n22489, n22490, n22491, n22492, n22494, n22495, n22496, n22497,
    n22498, n22500, n22501, n22503, n22504, n22506, n22507, n22509, n22510,
    n22512, n22513, n22515, n22516, n22518, n22519, n22521, n22522, n22523,
    n22524, n22525, n22526, n22527, n22528, n22529, n22530, n22531, n22532,
    n22533, n22534, n22535, n22537, n22538, n22539, n22540, n22541, n22543,
    n22544, n22545, n22547, n22548, n22549, n22550, n22551, n22552, n22553,
    n22554, n22555, n22556, n22557, n22560, n22562, n22563, n22564, n22566,
    n22567, n22568, n22569, n22570, n22573, n22575, n22577, n22578, n22579,
    n22580, n22581, n22582, n22584, n22585, n22587, n22588, n22589, n22590,
    n22593, n22594, n22596, n22597, n22599, n22600, n22602, n22603, n22605,
    n22606, n22608, n22609, n22611, n22612, n22614, n22615, n22617, n22618,
    n22620, n22621, n22623, n22624, n22626, n22627, n22629, n22630, n22632,
    n22633, n22635, n22636, n22638, n22639, n22641, n22642, n22644, n22645,
    n22647, n22648, n22650, n22651, n22653, n22654, n22656, n22657, n22659,
    n22660, n22662, n22663, n22665, n22666, n22668, n22669, n22671, n22672,
    n22674, n22675, n22677, n22678, n22680, n22681, n22683, n22684, n22686,
    n22687, n22689, n22690, n22692, n22693, n22695, n22696, n22698, n22699,
    n22701, n22702, n22704, n22705, n22707, n22708, n22710, n22711, n22713,
    n22714, n22716, n22717, n22719, n22720, n22722, n22723, n22725, n22726,
    n22728, n22729, n22731, n22732, n22734, n22735, n22737, n22738, n22740,
    n22741, n22743, n22744, n22746, n22747, n22749, n22750, n22752, n22753,
    n22755, n22756, n22758, n22759, n22761, n22762, n22764, n22765, n22767,
    n22768, n22770, n22771, n22773, n22774, n22776, n22777, n22779, n22780,
    n22782, n22783, n22785, n22786, n22788, n22789, n22791, n22792, n22794,
    n22795, n22797, n22798, n22800, n22801, n22803, n22804, n22806, n22807,
    n22809, n22810, n22812, n22813, n22815, n22816, n22818, n22819, n22821,
    n22822, n22824, n22825, n22827, n22828, n22830, n22831, n22833, n22834,
    n22836, n22837, n22839, n22840, n22842, n22843, n22845, n22846, n22849,
    n22850, n22852, n22853, n22855, n22856, n22858, n22859, n22861, n22862,
    n22864, n22865, n22867, n22868, n22870, n22871, n22873, n22874, n22876,
    n22877, n22879, n22880, n22882, n22883, n22885, n22886, n22888, n22889,
    n22891, n22892, n22894, n22895, n22897, n22898, n22900, n22901, n22903,
    n22904, n22906, n22907, n22909, n22910, n22912, n22913, n22915, n22916,
    n22918, n22919, n22921, n22922, n22924, n22925, n22927, n22928, n22930,
    n22931, n22933, n22934, n22936, n22937, n22939, n22940, n22942, n22943,
    n22945, n22946, n22948, n22949, n22951, n22952, n22954, n22955, n22957,
    n22958, n22960, n22961, n22963, n22964, n22966, n22967, n22969, n22970,
    n22972, n22973, n22975, n22976, n22978, n22979;
  assign n1459 = ~pi159 & pi490;
  assign n1460 = pi159 & ~pi490;
  assign n1461 = ~n1459 & ~n1460;
  assign n1462 = pi529 & ~n1461;
  assign n1463 = pi072 & ~pi108;
  assign n1464 = ~pi107 & n1463;
  assign n1465 = ~pi014 & n1464;
  assign n1466 = pi082 & pi108;
  assign n1467 = pi072 & n1466;
  assign n1468 = ~pi014 & n1467;
  assign n1469 = ~n1465 & ~n1468;
  assign n1470 = ~pi083 & ~n1469;
  assign n1471 = ~pi072 & pi108;
  assign n1472 = ~pi107 & n1471;
  assign n1473 = pi014 & n1472;
  assign n1474 = ~pi083 & n1473;
  assign n1475 = ~n1470 & ~n1474;
  assign n1476 = pi072 & pi108;
  assign n1477 = pi107 & n1476;
  assign n1478 = ~pi014 & n1477;
  assign n1479 = n1475 & ~n1478;
  assign n1480 = ~pi040 & ~n1479;
  assign n1481 = pi082 & ~pi108;
  assign n1482 = pi072 & n1481;
  assign n1483 = ~pi107 & n1482;
  assign n1484 = ~pi014 & n1483;
  assign n1485 = ~pi082 & ~pi108;
  assign n1486 = ~pi072 & n1485;
  assign n1487 = pi107 & n1486;
  assign n1488 = pi014 & n1487;
  assign n1489 = ~n1484 & ~n1488;
  assign n1490 = ~pi083 & ~n1489;
  assign n1491 = ~pi040 & pi083;
  assign n1492 = ~pi072 & n1466;
  assign n1493 = pi107 & n1492;
  assign n1494 = pi014 & n1493;
  assign n1495 = pi072 & pi082;
  assign n1496 = pi107 & n1495;
  assign n1497 = ~pi014 & n1496;
  assign n1498 = ~n1494 & ~n1497;
  assign n1499 = pi014 & n1486;
  assign n1500 = n1498 & ~n1499;
  assign n1501 = n1491 & ~n1500;
  assign n1502 = ~n1490 & ~n1501;
  assign n1503 = ~n1480 & n1502;
  assign n1504 = pi107 & n1482;
  assign n1505 = pi014 & n1504;
  assign n1506 = ~n1487 & ~n1505;
  assign n1507 = ~pi083 & ~n1506;
  assign n1508 = pi014 & pi083;
  assign n1509 = pi072 & n1485;
  assign n1510 = pi107 & n1509;
  assign n1511 = pi107 & n1467;
  assign n1512 = ~n1510 & ~n1511;
  assign n1513 = n1508 & ~n1512;
  assign n1514 = ~pi107 & n1486;
  assign n1515 = n1508 & n1514;
  assign n1516 = ~n1513 & ~n1515;
  assign n1517 = ~pi014 & pi083;
  assign n1518 = ~pi072 & pi082;
  assign n1519 = pi107 & n1518;
  assign n1520 = n1517 & n1519;
  assign n1521 = pi014 & ~pi082;
  assign n1522 = pi107 & n1521;
  assign n1523 = ~pi072 & n1481;
  assign n1524 = pi014 & n1523;
  assign n1525 = ~n1522 & ~n1524;
  assign n1526 = ~pi083 & ~n1525;
  assign n1527 = ~n1520 & ~n1526;
  assign n1528 = ~pi082 & pi108;
  assign n1529 = pi072 & n1528;
  assign n1530 = pi014 & n1529;
  assign n1531 = n1527 & ~n1530;
  assign n1532 = ~pi014 & pi107;
  assign n1533 = n1492 & n1532;
  assign n1534 = n1531 & ~n1533;
  assign n1535 = pi040 & ~n1534;
  assign n1536 = ~n1470 & ~n1535;
  assign n1537 = n1516 & n1536;
  assign n1538 = ~n1507 & n1537;
  assign n1539 = ~pi107 & pi108;
  assign n1540 = ~pi083 & n1539;
  assign n1541 = ~pi107 & n1476;
  assign n1542 = pi014 & n1541;
  assign n1543 = ~n1540 & ~n1542;
  assign n1544 = ~pi040 & ~n1543;
  assign n1545 = pi107 & n1471;
  assign n1546 = n1508 & n1545;
  assign n1547 = pi083 & n1486;
  assign n1548 = ~n1546 & ~n1547;
  assign n1549 = ~pi040 & ~n1548;
  assign n1550 = ~n1544 & ~n1549;
  assign n1551 = n1538 & n1550;
  assign n1552 = ~pi078 & ~n1551;
  assign n1553 = pi107 & n1481;
  assign n1554 = ~pi014 & n1553;
  assign n1555 = ~pi083 & n1554;
  assign n1556 = ~pi072 & ~pi082;
  assign n1557 = pi107 & n1556;
  assign n1558 = ~n1496 & ~n1557;
  assign n1559 = ~n1553 & n1558;
  assign n1560 = ~pi083 & ~n1559;
  assign n1561 = ~pi083 & n1482;
  assign n1562 = ~pi014 & n1472;
  assign n1563 = pi083 & n1562;
  assign n1564 = ~pi014 & n1481;
  assign n1565 = ~pi083 & n1564;
  assign n1566 = ~n1563 & ~n1565;
  assign n1567 = ~n1561 & n1566;
  assign n1568 = ~n1560 & n1567;
  assign n1569 = pi072 & ~pi082;
  assign n1570 = ~pi107 & n1569;
  assign n1571 = pi014 & n1570;
  assign n1572 = ~n1554 & ~n1571;
  assign n1573 = n1568 & n1572;
  assign n1574 = ~pi040 & ~n1573;
  assign n1575 = ~pi107 & n1518;
  assign n1576 = n1508 & n1575;
  assign n1577 = ~pi107 & n1466;
  assign n1578 = ~pi014 & n1577;
  assign n1579 = pi107 & n1569;
  assign n1580 = ~pi014 & n1579;
  assign n1581 = ~n1578 & ~n1580;
  assign n1582 = ~n1504 & n1581;
  assign n1583 = pi083 & ~n1582;
  assign n1584 = ~n1576 & ~n1583;
  assign n1585 = n1463 & n1532;
  assign n1586 = n1584 & ~n1585;
  assign n1587 = pi040 & pi083;
  assign n1588 = ~pi014 & n1485;
  assign n1589 = ~n1557 & ~n1588;
  assign n1590 = pi014 & n1481;
  assign n1591 = pi082 & ~pi107;
  assign n1592 = ~n1590 & ~n1591;
  assign n1593 = n1589 & n1592;
  assign n1594 = n1587 & ~n1593;
  assign n1595 = ~pi014 & ~pi083;
  assign n1596 = ~pi072 & n1528;
  assign n1597 = n1595 & n1596;
  assign n1598 = ~n1494 & ~n1597;
  assign n1599 = pi040 & ~n1598;
  assign n1600 = ~n1594 & ~n1599;
  assign n1601 = n1586 & n1600;
  assign n1602 = ~n1574 & n1601;
  assign n1603 = ~n1555 & n1602;
  assign n1604 = pi078 & ~n1603;
  assign n1605 = ~pi107 & n1523;
  assign n1606 = ~pi107 & n1467;
  assign n1607 = ~n1605 & ~n1606;
  assign n1608 = ~n1579 & n1607;
  assign n1609 = pi014 & ~n1608;
  assign n1610 = pi014 & n1509;
  assign n1611 = ~n1609 & ~n1610;
  assign n1612 = ~pi083 & ~n1611;
  assign n1613 = pi014 & n1482;
  assign n1614 = ~pi107 & n1492;
  assign n1615 = ~n1613 & ~n1614;
  assign n1616 = ~pi107 & n1509;
  assign n1617 = ~n1577 & ~n1616;
  assign n1618 = pi107 & n1596;
  assign n1619 = n1617 & ~n1618;
  assign n1620 = ~pi014 & ~n1619;
  assign n1621 = n1615 & ~n1620;
  assign n1622 = pi083 & ~n1621;
  assign n1623 = ~n1612 & ~n1622;
  assign n1624 = pi040 & ~n1623;
  assign n1625 = ~n1604 & ~n1624;
  assign n1626 = ~n1552 & n1625;
  assign n1627 = n1503 & n1626;
  assign n1628 = pi014 & n1467;
  assign n1629 = pi107 & n1529;
  assign n1630 = ~pi014 & n1629;
  assign n1631 = ~n1628 & ~n1630;
  assign n1632 = ~n1562 & n1631;
  assign n1633 = ~pi083 & ~n1632;
  assign n1634 = ~pi072 & ~pi083;
  assign n1635 = ~pi108 & n1634;
  assign n1636 = ~pi082 & n1635;
  assign n1637 = ~pi014 & n1569;
  assign n1638 = ~n1529 & ~n1637;
  assign n1639 = ~n1545 & n1638;
  assign n1640 = pi083 & ~n1639;
  assign n1641 = pi014 & n1492;
  assign n1642 = ~n1640 & ~n1641;
  assign n1643 = ~n1636 & n1642;
  assign n1644 = ~n1629 & n1643;
  assign n1645 = ~n1478 & ~n1565;
  assign n1646 = n1644 & n1645;
  assign n1647 = pi040 & ~n1646;
  assign n1648 = pi014 & ~pi107;
  assign n1649 = n1482 & n1648;
  assign n1650 = ~n1647 & ~n1649;
  assign n1651 = ~n1633 & n1650;
  assign n1652 = pi014 & n1618;
  assign n1653 = ~pi014 & n1492;
  assign n1654 = ~n1524 & ~n1653;
  assign n1655 = ~pi083 & ~n1654;
  assign n1656 = pi014 & n1596;
  assign n1657 = pi083 & n1656;
  assign n1658 = pi083 & n1482;
  assign n1659 = pi083 & n1464;
  assign n1660 = ~n1658 & ~n1659;
  assign n1661 = ~n1657 & n1660;
  assign n1662 = ~n1655 & n1661;
  assign n1663 = ~pi107 & n1485;
  assign n1664 = ~pi014 & n1663;
  assign n1665 = ~pi014 & ~pi107;
  assign n1666 = n1495 & n1665;
  assign n1667 = ~n1664 & ~n1666;
  assign n1668 = n1662 & n1667;
  assign n1669 = ~n1652 & n1668;
  assign n1670 = ~pi040 & ~n1669;
  assign n1671 = n1651 & ~n1670;
  assign n1672 = pi014 & n1528;
  assign n1673 = pi107 & n1672;
  assign n1674 = ~n1523 & ~n1596;
  assign n1675 = pi107 & ~n1674;
  assign n1676 = ~n1673 & ~n1675;
  assign n1677 = pi083 & ~n1676;
  assign n1678 = n1671 & ~n1677;
  assign n1679 = pi078 & ~n1678;
  assign n1680 = pi107 & n1523;
  assign n1681 = pi014 & n1680;
  assign n1682 = pi014 & n1577;
  assign n1683 = ~pi040 & ~pi083;
  assign n1684 = n1682 & n1683;
  assign n1685 = ~n1681 & ~n1684;
  assign n1686 = n1508 & n1614;
  assign n1687 = pi083 & n1652;
  assign n1688 = ~n1686 & ~n1687;
  assign n1689 = n1495 & n1648;
  assign n1690 = ~n1641 & ~n1689;
  assign n1691 = pi083 & ~n1690;
  assign n1692 = ~pi107 & n1596;
  assign n1693 = pi014 & ~pi083;
  assign n1694 = n1692 & n1693;
  assign n1695 = pi083 & pi107;
  assign n1696 = pi072 & n1695;
  assign n1697 = n1528 & n1696;
  assign n1698 = ~n1694 & ~n1697;
  assign n1699 = ~pi107 & n1529;
  assign n1700 = ~n1557 & ~n1699;
  assign n1701 = ~pi107 & n1481;
  assign n1702 = n1700 & ~n1701;
  assign n1703 = n1595 & ~n1702;
  assign n1704 = n1698 & ~n1703;
  assign n1705 = ~n1691 & n1704;
  assign n1706 = pi040 & ~n1705;
  assign n1707 = ~pi014 & n1487;
  assign n1708 = pi083 & n1707;
  assign n1709 = n1517 & n1605;
  assign n1710 = ~n1708 & ~n1709;
  assign n1711 = ~pi040 & ~n1710;
  assign n1712 = ~n1706 & ~n1711;
  assign n1713 = n1688 & n1712;
  assign n1714 = n1685 & n1713;
  assign n1715 = ~pi083 & n1699;
  assign n1716 = ~pi014 & n1504;
  assign n1717 = ~pi072 & ~pi108;
  assign n1718 = ~pi107 & n1717;
  assign n1719 = ~n1716 & ~n1718;
  assign n1720 = pi083 & ~n1719;
  assign n1721 = ~pi014 & n1606;
  assign n1722 = ~n1656 & ~n1721;
  assign n1723 = pi014 & n1511;
  assign n1724 = n1722 & ~n1723;
  assign n1725 = ~n1720 & n1724;
  assign n1726 = ~n1715 & n1725;
  assign n1727 = pi040 & ~n1726;
  assign n1728 = pi083 & n1606;
  assign n1729 = n1508 & n1718;
  assign n1730 = ~pi014 & n1511;
  assign n1731 = pi014 & n1553;
  assign n1732 = ~n1730 & ~n1731;
  assign n1733 = ~pi083 & ~n1732;
  assign n1734 = ~pi014 & n1605;
  assign n1735 = ~n1733 & ~n1734;
  assign n1736 = ~n1729 & n1735;
  assign n1737 = ~n1728 & n1736;
  assign n1738 = n1629 & n1693;
  assign n1739 = ~n1487 & ~n1562;
  assign n1740 = ~n1466 & ~n1476;
  assign n1741 = n1517 & ~n1740;
  assign n1742 = pi107 & n1485;
  assign n1743 = pi083 & n1742;
  assign n1744 = ~n1741 & ~n1743;
  assign n1745 = n1739 & n1744;
  assign n1746 = ~n1738 & n1745;
  assign n1747 = ~pi040 & ~n1746;
  assign n1748 = n1737 & ~n1747;
  assign n1749 = ~n1727 & n1748;
  assign n1750 = ~pi078 & ~n1749;
  assign n1751 = n1714 & ~n1750;
  assign n1752 = ~n1679 & n1751;
  assign n1753 = ~n1627 & n1752;
  assign n1754 = n1627 & ~n1752;
  assign n1755 = ~n1753 & ~n1754;
  assign n1756 = pi021 & pi098;
  assign n1757 = ~pi054 & n1756;
  assign n1758 = pi007 & n1757;
  assign n1759 = ~pi013 & n1758;
  assign n1760 = ~pi114 & n1759;
  assign n1761 = pi021 & ~pi054;
  assign n1762 = ~pi007 & n1761;
  assign n1763 = ~pi013 & n1762;
  assign n1764 = ~pi021 & ~pi098;
  assign n1765 = ~pi054 & n1764;
  assign n1766 = pi007 & n1765;
  assign n1767 = pi013 & n1766;
  assign n1768 = ~n1763 & ~n1767;
  assign n1769 = pi114 & ~n1768;
  assign n1770 = pi021 & ~pi098;
  assign n1771 = pi007 & n1770;
  assign n1772 = pi013 & n1771;
  assign n1773 = pi001 & n1772;
  assign n1774 = ~pi021 & pi098;
  assign n1775 = ~pi054 & n1774;
  assign n1776 = ~pi007 & n1775;
  assign n1777 = pi054 & n1774;
  assign n1778 = pi007 & n1777;
  assign n1779 = ~pi013 & n1777;
  assign n1780 = ~n1778 & ~n1779;
  assign n1781 = ~n1776 & n1780;
  assign n1782 = pi001 & ~pi114;
  assign n1783 = ~n1781 & n1782;
  assign n1784 = ~n1773 & ~n1783;
  assign n1785 = pi021 & pi054;
  assign n1786 = pi007 & n1785;
  assign n1787 = pi114 & n1786;
  assign n1788 = pi114 & n1765;
  assign n1789 = ~n1787 & ~n1788;
  assign n1790 = ~pi001 & ~n1789;
  assign n1791 = ~pi013 & ~pi114;
  assign n1792 = pi054 & n1770;
  assign n1793 = n1791 & n1792;
  assign n1794 = ~pi007 & n1764;
  assign n1795 = pi013 & n1794;
  assign n1796 = ~n1793 & ~n1795;
  assign n1797 = ~pi001 & ~n1796;
  assign n1798 = ~n1790 & ~n1797;
  assign n1799 = n1784 & n1798;
  assign n1800 = ~n1769 & n1799;
  assign n1801 = ~n1760 & n1800;
  assign n1802 = ~pi007 & ~pi013;
  assign n1803 = pi054 & n1764;
  assign n1804 = n1802 & n1803;
  assign n1805 = ~pi013 & pi114;
  assign n1806 = ~pi054 & pi098;
  assign n1807 = pi007 & n1806;
  assign n1808 = n1805 & n1807;
  assign n1809 = pi114 & n1792;
  assign n1810 = ~n1808 & ~n1809;
  assign n1811 = pi001 & ~n1810;
  assign n1812 = ~n1804 & ~n1811;
  assign n1813 = n1801 & n1812;
  assign n1814 = ~pi029 & ~n1813;
  assign n1815 = ~pi013 & n1771;
  assign n1816 = pi114 & n1815;
  assign n1817 = pi013 & n1803;
  assign n1818 = pi114 & n1817;
  assign n1819 = pi013 & n1758;
  assign n1820 = ~n1818 & ~n1819;
  assign n1821 = ~n1761 & ~n1806;
  assign n1822 = pi013 & ~n1821;
  assign n1823 = pi054 & n1756;
  assign n1824 = ~pi007 & n1823;
  assign n1825 = ~pi013 & n1824;
  assign n1826 = ~n1822 & ~n1825;
  assign n1827 = n1765 & n1802;
  assign n1828 = n1826 & ~n1827;
  assign n1829 = ~pi114 & ~n1828;
  assign n1830 = pi013 & n1776;
  assign n1831 = ~n1829 & ~n1830;
  assign n1832 = n1820 & n1831;
  assign n1833 = ~n1816 & n1832;
  assign n1834 = pi001 & ~n1833;
  assign n1835 = ~pi021 & pi054;
  assign n1836 = ~pi007 & n1835;
  assign n1837 = pi013 & n1836;
  assign n1838 = pi007 & pi013;
  assign n1839 = ~n1802 & ~n1838;
  assign n1840 = n1775 & ~n1839;
  assign n1841 = pi013 & n1792;
  assign n1842 = ~pi013 & n1803;
  assign n1843 = ~n1841 & ~n1842;
  assign n1844 = ~n1840 & n1843;
  assign n1845 = ~n1837 & n1844;
  assign n1846 = pi114 & ~n1845;
  assign n1847 = pi007 & n1792;
  assign n1848 = pi013 & n1847;
  assign n1849 = pi007 & n1761;
  assign n1850 = ~pi013 & n1849;
  assign n1851 = pi013 & n1824;
  assign n1852 = ~n1850 & ~n1851;
  assign n1853 = ~pi013 & n1757;
  assign n1854 = n1852 & ~n1853;
  assign n1855 = ~pi114 & ~n1854;
  assign n1856 = ~n1848 & ~n1855;
  assign n1857 = ~n1846 & n1856;
  assign n1858 = ~n1804 & n1857;
  assign n1859 = ~pi001 & ~n1858;
  assign n1860 = ~n1834 & ~n1859;
  assign n1861 = ~n1814 & n1860;
  assign n1862 = ~pi054 & n1770;
  assign n1863 = ~pi007 & n1862;
  assign n1864 = ~pi114 & n1863;
  assign n1865 = ~n1787 & ~n1864;
  assign n1866 = pi013 & ~n1865;
  assign n1867 = ~pi007 & n1774;
  assign n1868 = pi114 & n1867;
  assign n1869 = ~pi007 & n1803;
  assign n1870 = pi013 & n1869;
  assign n1871 = ~pi007 & n1770;
  assign n1872 = pi007 & n1775;
  assign n1873 = ~n1871 & ~n1872;
  assign n1874 = ~pi114 & ~n1873;
  assign n1875 = ~n1870 & ~n1874;
  assign n1876 = ~n1868 & n1875;
  assign n1877 = pi007 & ~pi013;
  assign n1878 = n1765 & n1877;
  assign n1879 = n1876 & ~n1878;
  assign n1880 = pi001 & ~n1879;
  assign n1881 = pi013 & n1775;
  assign n1882 = pi013 & ~pi021;
  assign n1883 = ~pi007 & n1882;
  assign n1884 = ~n1881 & ~n1883;
  assign n1885 = ~pi013 & ~pi098;
  assign n1886 = pi007 & n1885;
  assign n1887 = ~n1824 & ~n1886;
  assign n1888 = n1884 & n1887;
  assign n1889 = pi114 & ~n1888;
  assign n1890 = pi013 & n1757;
  assign n1891 = pi013 & n1871;
  assign n1892 = ~n1827 & ~n1891;
  assign n1893 = ~n1890 & n1892;
  assign n1894 = ~pi114 & ~n1893;
  assign n1895 = ~n1889 & ~n1894;
  assign n1896 = pi054 & pi098;
  assign n1897 = ~pi007 & n1896;
  assign n1898 = ~pi114 & n1897;
  assign n1899 = ~pi007 & n1756;
  assign n1900 = pi013 & n1899;
  assign n1901 = pi007 & n1764;
  assign n1902 = pi013 & n1901;
  assign n1903 = ~pi114 & n1902;
  assign n1904 = pi013 & n1896;
  assign n1905 = ~n1903 & ~n1904;
  assign n1906 = ~n1900 & n1905;
  assign n1907 = ~n1898 & n1906;
  assign n1908 = pi114 & n1778;
  assign n1909 = n1907 & ~n1908;
  assign n1910 = ~pi001 & ~n1909;
  assign n1911 = n1895 & ~n1910;
  assign n1912 = ~n1880 & n1911;
  assign n1913 = pi029 & ~n1912;
  assign n1914 = ~n1866 & ~n1913;
  assign n1915 = n1861 & n1914;
  assign n1916 = ~pi023 & ~pi027;
  assign n1917 = ~pi047 & ~pi093;
  assign n1918 = pi111 & n1917;
  assign n1919 = n1916 & n1918;
  assign n1920 = pi047 & ~pi111;
  assign n1921 = ~pi023 & n1920;
  assign n1922 = ~pi027 & n1921;
  assign n1923 = ~pi111 & n1917;
  assign n1924 = pi023 & n1923;
  assign n1925 = pi027 & n1924;
  assign n1926 = ~n1922 & ~n1925;
  assign n1927 = pi123 & ~n1926;
  assign n1928 = ~pi047 & pi093;
  assign n1929 = ~pi111 & n1928;
  assign n1930 = ~pi023 & n1929;
  assign n1931 = pi111 & n1928;
  assign n1932 = pi023 & n1931;
  assign n1933 = ~n1930 & ~n1932;
  assign n1934 = ~pi027 & n1931;
  assign n1935 = n1933 & ~n1934;
  assign n1936 = ~pi123 & ~n1935;
  assign n1937 = pi047 & ~pi093;
  assign n1938 = pi111 & n1937;
  assign n1939 = pi123 & n1938;
  assign n1940 = pi023 & n1937;
  assign n1941 = pi027 & n1940;
  assign n1942 = ~n1939 & ~n1941;
  assign n1943 = ~pi027 & pi123;
  assign n1944 = pi093 & ~pi111;
  assign n1945 = pi023 & n1944;
  assign n1946 = n1943 & n1945;
  assign n1947 = n1942 & ~n1946;
  assign n1948 = ~n1936 & n1947;
  assign n1949 = pi048 & ~n1948;
  assign n1950 = pi047 & pi093;
  assign n1951 = ~pi111 & n1950;
  assign n1952 = pi023 & n1951;
  assign n1953 = ~pi027 & n1952;
  assign n1954 = ~pi123 & n1953;
  assign n1955 = ~pi023 & n1917;
  assign n1956 = pi027 & n1955;
  assign n1957 = pi123 & n1923;
  assign n1958 = ~n1956 & ~n1957;
  assign n1959 = pi047 & pi111;
  assign n1960 = pi023 & n1959;
  assign n1961 = pi123 & n1960;
  assign n1962 = ~pi027 & n1938;
  assign n1963 = ~pi123 & n1962;
  assign n1964 = ~n1961 & ~n1963;
  assign n1965 = n1958 & n1964;
  assign n1966 = ~pi048 & ~n1965;
  assign n1967 = ~n1954 & ~n1966;
  assign n1968 = ~n1949 & n1967;
  assign n1969 = ~n1927 & n1968;
  assign n1970 = ~n1919 & n1969;
  assign n1971 = ~pi020 & ~n1970;
  assign n1972 = pi023 & pi027;
  assign n1973 = pi123 & n1959;
  assign n1974 = n1972 & n1973;
  assign n1975 = pi027 & ~pi123;
  assign n1976 = ~pi111 & n1937;
  assign n1977 = ~pi023 & n1976;
  assign n1978 = n1975 & n1977;
  assign n1979 = ~n1974 & ~n1978;
  assign n1980 = ~pi027 & n1940;
  assign n1981 = pi123 & n1980;
  assign n1982 = pi027 & pi123;
  assign n1983 = pi111 & n1982;
  assign n1984 = n1917 & n1983;
  assign n1985 = ~n1981 & ~n1984;
  assign n1986 = pi048 & ~n1985;
  assign n1987 = n1979 & ~n1986;
  assign n1988 = pi027 & n1930;
  assign n1989 = ~n1920 & ~n1944;
  assign n1990 = pi027 & ~n1989;
  assign n1991 = pi111 & n1950;
  assign n1992 = ~pi023 & n1991;
  assign n1993 = ~pi027 & n1992;
  assign n1994 = ~n1990 & ~n1993;
  assign n1995 = ~pi023 & n1923;
  assign n1996 = ~pi027 & n1995;
  assign n1997 = n1994 & ~n1996;
  assign n1998 = ~pi123 & ~n1997;
  assign n1999 = ~n1988 & ~n1998;
  assign n2000 = pi027 & n1952;
  assign n2001 = n1999 & ~n2000;
  assign n2002 = pi048 & ~n2001;
  assign n2003 = pi023 & n1938;
  assign n2004 = pi027 & n2003;
  assign n2005 = pi023 & n1929;
  assign n2006 = pi027 & n2005;
  assign n2007 = ~pi111 & n1916;
  assign n2008 = n1928 & n2007;
  assign n2009 = ~n2006 & ~n2008;
  assign n2010 = pi027 & n1938;
  assign n2011 = ~pi027 & n1918;
  assign n2012 = ~pi047 & pi111;
  assign n2013 = ~pi023 & n2012;
  assign n2014 = pi027 & n2013;
  assign n2015 = ~n2011 & ~n2014;
  assign n2016 = ~n2010 & n2015;
  assign n2017 = n2009 & n2016;
  assign n2018 = pi123 & ~n2017;
  assign n2019 = pi023 & n1920;
  assign n2020 = ~pi027 & n2019;
  assign n2021 = pi027 & n1992;
  assign n2022 = ~n2020 & ~n2021;
  assign n2023 = ~pi027 & n1951;
  assign n2024 = n2022 & ~n2023;
  assign n2025 = ~pi123 & ~n2024;
  assign n2026 = ~n2018 & ~n2025;
  assign n2027 = ~n2004 & n2026;
  assign n2028 = ~n1919 & n2027;
  assign n2029 = ~pi048 & ~n2028;
  assign n2030 = ~n2002 & ~n2029;
  assign n2031 = pi027 & n1929;
  assign n2032 = ~pi023 & pi027;
  assign n2033 = ~pi047 & n2032;
  assign n2034 = ~n2031 & ~n2033;
  assign n2035 = pi123 & ~n2034;
  assign n2036 = n1917 & n1972;
  assign n2037 = ~pi123 & n2036;
  assign n2038 = pi093 & pi111;
  assign n2039 = pi027 & n2038;
  assign n2040 = ~n2037 & ~n2039;
  assign n2041 = ~pi023 & n2038;
  assign n2042 = ~pi123 & n2041;
  assign n2043 = ~pi023 & n1950;
  assign n2044 = pi027 & n2043;
  assign n2045 = ~n2042 & ~n2044;
  assign n2046 = n2040 & n2045;
  assign n2047 = pi123 & n1932;
  assign n2048 = n2046 & ~n2047;
  assign n2049 = ~pi048 & ~n2048;
  assign n2050 = ~pi027 & n1924;
  assign n2051 = ~pi023 & n1918;
  assign n2052 = pi027 & n2051;
  assign n2053 = ~n2050 & ~n2052;
  assign n2054 = ~pi023 & n1928;
  assign n2055 = pi123 & n2054;
  assign n2056 = ~pi023 & n1937;
  assign n2057 = ~n2005 & ~n2056;
  assign n2058 = ~pi123 & ~n2057;
  assign n2059 = ~n2055 & ~n2058;
  assign n2060 = n2053 & n2059;
  assign n2061 = pi048 & ~n2060;
  assign n2062 = ~n2049 & ~n2061;
  assign n2063 = ~pi027 & ~pi093;
  assign n2064 = pi023 & n2063;
  assign n2065 = ~n1992 & ~n2064;
  assign n2066 = pi123 & ~n2065;
  assign n2067 = pi027 & n2056;
  assign n2068 = pi027 & n1951;
  assign n2069 = ~n2067 & ~n2068;
  assign n2070 = ~n1996 & n2069;
  assign n2071 = ~pi123 & ~n2070;
  assign n2072 = ~n2066 & ~n2071;
  assign n2073 = n2062 & n2072;
  assign n2074 = ~n2035 & n2073;
  assign n2075 = pi020 & ~n2074;
  assign n2076 = n2030 & ~n2075;
  assign n2077 = n1987 & n2076;
  assign n2078 = ~n1971 & n2077;
  assign n2079 = ~n1915 & n2078;
  assign n2080 = n1915 & ~n2078;
  assign n2081 = ~n2079 & ~n2080;
  assign n2082 = ~n1755 & n2081;
  assign n2083 = n1755 & ~n2081;
  assign n2084 = ~n2082 & ~n2083;
  assign n2085 = pi063 & ~pi126;
  assign n2086 = ~pi033 & n2085;
  assign n2087 = ~pi127 & n2086;
  assign n2088 = pi069 & n2087;
  assign n2089 = ~pi104 & n2088;
  assign n2090 = pi069 & pi104;
  assign n2091 = pi033 & pi063;
  assign n2092 = pi127 & n2091;
  assign n2093 = n2090 & n2092;
  assign n2094 = ~n2089 & ~n2093;
  assign n2095 = ~pi063 & ~pi126;
  assign n2096 = pi033 & n2095;
  assign n2097 = ~pi069 & n2096;
  assign n2098 = ~pi127 & n2097;
  assign n2099 = ~pi126 & n2091;
  assign n2100 = pi127 & n2099;
  assign n2101 = pi069 & n2100;
  assign n2102 = ~n2098 & ~n2101;
  assign n2103 = ~pi063 & pi126;
  assign n2104 = ~pi033 & n2103;
  assign n2105 = ~pi069 & ~pi127;
  assign n2106 = pi069 & pi127;
  assign n2107 = ~n2105 & ~n2106;
  assign n2108 = n2104 & ~n2107;
  assign n2109 = pi033 & ~pi063;
  assign n2110 = ~pi127 & n2109;
  assign n2111 = pi069 & n2110;
  assign n2112 = pi069 & n2099;
  assign n2113 = ~n2111 & ~n2112;
  assign n2114 = ~n2108 & n2113;
  assign n2115 = ~n2097 & n2114;
  assign n2116 = pi104 & ~n2115;
  assign n2117 = ~pi033 & pi063;
  assign n2118 = pi127 & n2117;
  assign n2119 = ~pi069 & n2118;
  assign n2120 = pi063 & pi126;
  assign n2121 = pi033 & n2120;
  assign n2122 = ~pi127 & n2121;
  assign n2123 = pi069 & n2122;
  assign n2124 = ~n2119 & ~n2123;
  assign n2125 = ~pi033 & n2120;
  assign n2126 = ~pi069 & n2125;
  assign n2127 = n2124 & ~n2126;
  assign n2128 = ~pi104 & ~n2127;
  assign n2129 = ~n2116 & ~n2128;
  assign n2130 = n2102 & n2129;
  assign n2131 = ~pi102 & ~n2130;
  assign n2132 = pi127 & n2125;
  assign n2133 = ~pi104 & n2132;
  assign n2134 = ~pi069 & n2133;
  assign n2135 = ~pi069 & ~pi104;
  assign n2136 = ~pi126 & n2135;
  assign n2137 = n2091 & n2136;
  assign n2138 = ~pi127 & n2095;
  assign n2139 = pi069 & n2138;
  assign n2140 = ~pi033 & n2095;
  assign n2141 = pi104 & n2140;
  assign n2142 = ~n2139 & ~n2141;
  assign n2143 = pi104 & n2092;
  assign n2144 = n2142 & ~n2143;
  assign n2145 = ~n2137 & n2144;
  assign n2146 = ~pi102 & ~n2145;
  assign n2147 = ~n2098 & ~n2146;
  assign n2148 = pi033 & n2103;
  assign n2149 = ~pi069 & n2148;
  assign n2150 = ~pi127 & n2104;
  assign n2151 = ~n2149 & ~n2150;
  assign n2152 = pi127 & n2148;
  assign n2153 = n2151 & ~n2152;
  assign n2154 = ~pi104 & ~n2153;
  assign n2155 = pi104 & n2099;
  assign n2156 = pi127 & n2085;
  assign n2157 = pi069 & n2156;
  assign n2158 = ~n2155 & ~n2157;
  assign n2159 = ~pi069 & pi104;
  assign n2160 = ~pi033 & pi126;
  assign n2161 = pi127 & n2160;
  assign n2162 = n2159 & n2161;
  assign n2163 = n2158 & ~n2162;
  assign n2164 = ~n2154 & n2163;
  assign n2165 = pi102 & ~n2164;
  assign n2166 = n2106 & n2140;
  assign n2167 = ~pi127 & n2117;
  assign n2168 = ~pi069 & n2167;
  assign n2169 = ~n2166 & ~n2168;
  assign n2170 = pi104 & ~n2169;
  assign n2171 = ~n2165 & ~n2170;
  assign n2172 = n2147 & n2171;
  assign n2173 = ~n2134 & n2172;
  assign n2174 = ~pi012 & ~n2173;
  assign n2175 = ~n2131 & ~n2174;
  assign n2176 = n2094 & n2175;
  assign n2177 = ~n2117 & ~n2160;
  assign n2178 = pi069 & ~n2177;
  assign n2179 = ~pi069 & n2122;
  assign n2180 = ~n2178 & ~n2179;
  assign n2181 = n2105 & n2140;
  assign n2182 = n2180 & ~n2181;
  assign n2183 = ~pi104 & ~n2182;
  assign n2184 = pi069 & n2150;
  assign n2185 = ~pi069 & n2156;
  assign n2186 = pi104 & n2185;
  assign n2187 = ~n2184 & ~n2186;
  assign n2188 = ~n2183 & n2187;
  assign n2189 = pi069 & n2096;
  assign n2190 = pi104 & n2189;
  assign n2191 = pi069 & n2132;
  assign n2192 = ~n2190 & ~n2191;
  assign n2193 = n2188 & n2192;
  assign n2194 = pi102 & ~n2193;
  assign n2195 = pi069 & ~pi127;
  assign n2196 = ~pi063 & n2195;
  assign n2197 = pi069 & n2104;
  assign n2198 = ~n2196 & ~n2197;
  assign n2199 = pi104 & ~n2198;
  assign n2200 = ~pi069 & pi127;
  assign n2201 = ~pi126 & n2200;
  assign n2202 = ~n2122 & ~n2201;
  assign n2203 = pi104 & ~n2202;
  assign n2204 = ~n2199 & ~n2203;
  assign n2205 = pi127 & n2140;
  assign n2206 = ~pi069 & n2205;
  assign n2207 = ~pi127 & n2096;
  assign n2208 = pi069 & n2207;
  assign n2209 = ~n2206 & ~n2208;
  assign n2210 = ~pi127 & n2103;
  assign n2211 = pi104 & n2210;
  assign n2212 = ~pi127 & n2085;
  assign n2213 = pi127 & n2104;
  assign n2214 = ~n2212 & ~n2213;
  assign n2215 = ~pi104 & ~n2214;
  assign n2216 = ~n2211 & ~n2215;
  assign n2217 = n2209 & n2216;
  assign n2218 = pi102 & ~n2217;
  assign n2219 = pi069 & n2212;
  assign n2220 = pi069 & n2125;
  assign n2221 = ~n2219 & ~n2220;
  assign n2222 = ~n2181 & n2221;
  assign n2223 = ~pi104 & ~n2222;
  assign n2224 = n2095 & n2106;
  assign n2225 = ~pi104 & n2224;
  assign n2226 = pi033 & pi126;
  assign n2227 = pi069 & n2226;
  assign n2228 = ~n2225 & ~n2227;
  assign n2229 = ~pi127 & n2226;
  assign n2230 = ~pi104 & n2229;
  assign n2231 = ~pi127 & n2120;
  assign n2232 = pi069 & n2231;
  assign n2233 = ~n2230 & ~n2232;
  assign n2234 = n2228 & n2233;
  assign n2235 = pi104 & n2152;
  assign n2236 = n2234 & ~n2235;
  assign n2237 = ~pi102 & ~n2236;
  assign n2238 = ~n2223 & ~n2237;
  assign n2239 = ~n2218 & n2238;
  assign n2240 = n2204 & n2239;
  assign n2241 = pi012 & ~n2240;
  assign n2242 = ~n2194 & ~n2241;
  assign n2243 = n2176 & n2242;
  assign n2244 = pi159 & n2243;
  assign n2245 = ~pi159 & ~n2243;
  assign n2246 = ~n2244 & ~n2245;
  assign n2247 = ~pi127 & n2160;
  assign n2248 = n2159 & n2247;
  assign n2249 = ~pi104 & n2099;
  assign n2250 = ~pi033 & ~pi063;
  assign n2251 = pi127 & n2250;
  assign n2252 = ~n2092 & ~n2251;
  assign n2253 = ~n2156 & n2252;
  assign n2254 = ~pi104 & ~n2253;
  assign n2255 = ~pi069 & n2085;
  assign n2256 = ~pi104 & n2255;
  assign n2257 = ~n2254 & ~n2256;
  assign n2258 = ~n2249 & n2257;
  assign n2259 = ~n2248 & n2258;
  assign n2260 = ~n2111 & ~n2185;
  assign n2261 = n2259 & n2260;
  assign n2262 = ~pi102 & ~n2261;
  assign n2263 = n2104 & n2135;
  assign n2264 = ~n2191 & ~n2263;
  assign n2265 = pi102 & ~n2264;
  assign n2266 = pi102 & pi104;
  assign n2267 = ~pi069 & n2095;
  assign n2268 = ~n2251 & ~n2267;
  assign n2269 = pi069 & n2085;
  assign n2270 = pi063 & ~pi127;
  assign n2271 = ~n2269 & ~n2270;
  assign n2272 = n2268 & n2271;
  assign n2273 = n2266 & ~n2272;
  assign n2274 = ~n2265 & ~n2273;
  assign n2275 = ~pi104 & n2185;
  assign n2276 = n2090 & n2167;
  assign n2277 = pi033 & ~pi126;
  assign n2278 = n2200 & n2277;
  assign n2279 = ~n2276 & ~n2278;
  assign n2280 = ~n2275 & n2279;
  assign n2281 = ~pi069 & n2231;
  assign n2282 = pi127 & n2109;
  assign n2283 = ~pi069 & n2282;
  assign n2284 = ~n2281 & ~n2283;
  assign n2285 = ~n2100 & n2284;
  assign n2286 = pi104 & ~n2285;
  assign n2287 = n2280 & ~n2286;
  assign n2288 = n2274 & n2287;
  assign n2289 = ~n2262 & n2288;
  assign n2290 = pi012 & ~n2289;
  assign n2291 = ~n2087 & ~n2122;
  assign n2292 = ~n2282 & n2291;
  assign n2293 = pi069 & ~n2292;
  assign n2294 = ~n2189 & ~n2293;
  assign n2295 = pi102 & ~pi104;
  assign n2296 = ~n2294 & n2295;
  assign n2297 = ~pi127 & n2125;
  assign n2298 = ~n2112 & ~n2297;
  assign n2299 = ~n2207 & ~n2231;
  assign n2300 = ~n2213 & n2299;
  assign n2301 = ~pi069 & ~n2300;
  assign n2302 = n2298 & ~n2301;
  assign n2303 = n2266 & ~n2302;
  assign n2304 = ~n2296 & ~n2303;
  assign n2305 = pi069 & n2247;
  assign n2306 = ~pi104 & n2305;
  assign n2307 = ~pi127 & n2277;
  assign n2308 = ~pi069 & n2307;
  assign n2309 = ~pi069 & n2121;
  assign n2310 = ~n2308 & ~n2309;
  assign n2311 = ~pi104 & ~n2310;
  assign n2312 = ~n2306 & ~n2311;
  assign n2313 = pi127 & n2226;
  assign n2314 = ~pi069 & n2313;
  assign n2315 = n2312 & ~n2314;
  assign n2316 = ~pi102 & ~n2315;
  assign n2317 = n2099 & n2105;
  assign n2318 = ~n2166 & ~n2317;
  assign n2319 = ~pi104 & ~n2318;
  assign n2320 = pi069 & n2140;
  assign n2321 = ~pi069 & n2092;
  assign n2322 = ~n2191 & ~n2321;
  assign n2323 = ~n2320 & n2322;
  assign n2324 = ~pi102 & pi104;
  assign n2325 = ~n2323 & n2324;
  assign n2326 = ~n2319 & ~n2325;
  assign n2327 = ~n2316 & n2326;
  assign n2328 = n2304 & n2327;
  assign n2329 = n2090 & n2161;
  assign n2330 = ~n2141 & ~n2329;
  assign n2331 = ~pi102 & ~n2330;
  assign n2332 = ~n2101 & ~n2205;
  assign n2333 = ~pi104 & ~n2332;
  assign n2334 = ~n2311 & ~n2333;
  assign n2335 = ~pi104 & ~pi127;
  assign n2336 = pi126 & n2335;
  assign n2337 = pi069 & n2229;
  assign n2338 = ~n2336 & ~n2337;
  assign n2339 = ~pi102 & ~n2338;
  assign n2340 = pi127 & n2096;
  assign n2341 = pi127 & n2121;
  assign n2342 = ~n2340 & ~n2341;
  assign n2343 = n2090 & ~n2342;
  assign n2344 = ~pi127 & n2090;
  assign n2345 = ~pi033 & n2344;
  assign n2346 = n2095 & n2345;
  assign n2347 = ~n2343 & ~n2346;
  assign n2348 = ~n2339 & n2347;
  assign n2349 = n2334 & n2348;
  assign n2350 = ~n2331 & n2349;
  assign n2351 = ~pi069 & n2132;
  assign n2352 = pi069 & n2148;
  assign n2353 = ~n2351 & ~n2352;
  assign n2354 = n2118 & n2159;
  assign n2355 = ~pi063 & n2106;
  assign n2356 = pi069 & n2086;
  assign n2357 = ~n2355 & ~n2356;
  assign n2358 = ~pi104 & ~n2357;
  assign n2359 = ~n2354 & ~n2358;
  assign n2360 = n2353 & n2359;
  assign n2361 = pi102 & ~n2360;
  assign n2362 = n2350 & ~n2361;
  assign n2363 = ~pi012 & ~n2362;
  assign n2364 = n2328 & ~n2363;
  assign n2365 = ~n2290 & n2364;
  assign n2366 = ~pi069 & n2247;
  assign n2367 = pi069 & n2121;
  assign n2368 = ~pi069 & n2152;
  assign n2369 = ~n2367 & ~n2368;
  assign n2370 = ~n2366 & n2369;
  assign n2371 = ~pi104 & ~n2370;
  assign n2372 = ~pi127 & n2099;
  assign n2373 = pi069 & n2372;
  assign n2374 = ~pi069 & n2109;
  assign n2375 = ~n2148 & ~n2374;
  assign n2376 = ~n2161 & n2375;
  assign n2377 = pi104 & ~n2376;
  assign n2378 = ~pi104 & n2140;
  assign n2379 = ~n2152 & ~n2220;
  assign n2380 = ~n2378 & n2379;
  assign n2381 = ~n2377 & n2380;
  assign n2382 = ~n2256 & ~n2314;
  assign n2383 = n2381 & n2382;
  assign n2384 = pi102 & ~n2383;
  assign n2385 = ~n2373 & ~n2384;
  assign n2386 = ~n2371 & n2385;
  assign n2387 = pi104 & n2307;
  assign n2388 = pi069 & ~pi104;
  assign n2389 = n2086 & n2388;
  assign n2390 = pi104 & n2197;
  assign n2391 = ~n2155 & ~n2390;
  assign n2392 = ~n2389 & n2391;
  assign n2393 = ~n2387 & n2392;
  assign n2394 = n2125 & n2135;
  assign n2395 = n2104 & n2106;
  assign n2396 = ~pi069 & n2138;
  assign n2397 = n2091 & n2105;
  assign n2398 = ~n2396 & ~n2397;
  assign n2399 = ~n2395 & n2398;
  assign n2400 = ~n2394 & n2399;
  assign n2401 = n2393 & n2400;
  assign n2402 = ~pi102 & ~n2401;
  assign n2403 = n2386 & ~n2402;
  assign n2404 = pi069 & n2103;
  assign n2405 = pi127 & n2404;
  assign n2406 = ~n2086 & ~n2104;
  assign n2407 = pi127 & ~n2406;
  assign n2408 = ~n2405 & ~n2407;
  assign n2409 = pi104 & ~n2408;
  assign n2410 = n2403 & ~n2409;
  assign n2411 = pi012 & ~n2410;
  assign n2412 = ~pi127 & n2148;
  assign n2413 = ~pi104 & n2412;
  assign n2414 = ~n2179 & ~n2197;
  assign n2415 = ~pi033 & ~pi126;
  assign n2416 = ~pi127 & n2415;
  assign n2417 = ~pi069 & n2100;
  assign n2418 = ~n2416 & ~n2417;
  assign n2419 = pi104 & ~n2418;
  assign n2420 = pi069 & n2341;
  assign n2421 = ~n2419 & ~n2420;
  assign n2422 = n2414 & n2421;
  assign n2423 = ~n2413 & n2422;
  assign n2424 = pi102 & ~n2423;
  assign n2425 = n2152 & n2388;
  assign n2426 = ~n2205 & ~n2366;
  assign n2427 = pi127 & n2095;
  assign n2428 = pi104 & n2427;
  assign n2429 = ~n2120 & ~n2226;
  assign n2430 = n2159 & ~n2429;
  assign n2431 = ~n2428 & ~n2430;
  assign n2432 = n2426 & n2431;
  assign n2433 = ~n2425 & n2432;
  assign n2434 = ~pi102 & ~n2433;
  assign n2435 = ~n2424 & ~n2434;
  assign n2436 = ~pi069 & n2087;
  assign n2437 = ~pi069 & n2341;
  assign n2438 = ~n2157 & ~n2437;
  assign n2439 = ~pi104 & ~n2438;
  assign n2440 = pi104 & n2122;
  assign n2441 = n2090 & n2416;
  assign n2442 = ~n2440 & ~n2441;
  assign n2443 = ~n2439 & n2442;
  assign n2444 = ~n2436 & n2443;
  assign n2445 = n2435 & n2444;
  assign n2446 = ~pi012 & ~n2445;
  assign n2447 = n2091 & n2195;
  assign n2448 = ~n2220 & ~n2447;
  assign n2449 = pi104 & ~n2448;
  assign n2450 = ~n2212 & ~n2412;
  assign n2451 = ~n2251 & n2450;
  assign n2452 = n2135 & ~n2451;
  assign n2453 = ~n2449 & ~n2452;
  assign n2454 = ~pi104 & n2184;
  assign n2455 = n2453 & ~n2454;
  assign n2456 = ~n2235 & n2455;
  assign n2457 = pi102 & ~n2456;
  assign n2458 = n2090 & n2297;
  assign n2459 = pi104 & n2395;
  assign n2460 = ~n2458 & ~n2459;
  assign n2461 = pi127 & n2086;
  assign n2462 = pi069 & n2461;
  assign n2463 = n2460 & ~n2462;
  assign n2464 = ~pi104 & n2232;
  assign n2465 = ~pi102 & n2464;
  assign n2466 = n2463 & ~n2465;
  assign n2467 = ~n2457 & n2466;
  assign n2468 = pi104 & n2206;
  assign n2469 = n2087 & n2159;
  assign n2470 = ~n2468 & ~n2469;
  assign n2471 = ~pi102 & ~n2470;
  assign n2472 = n2467 & ~n2471;
  assign n2473 = ~n2446 & n2472;
  assign n2474 = ~n2411 & n2473;
  assign n2475 = ~n2365 & n2474;
  assign n2476 = n2365 & ~n2474;
  assign n2477 = ~n2475 & ~n2476;
  assign n2478 = ~n2246 & ~n2477;
  assign n2479 = n2246 & n2477;
  assign n2480 = ~n2478 & ~n2479;
  assign n2481 = ~n2084 & n2480;
  assign n2482 = n2084 & ~n2480;
  assign n2483 = ~n2481 & ~n2482;
  assign n2484 = ~pi529 & n2483;
  assign po130 = n1462 | n2484;
  assign n2486 = pi267 & pi503;
  assign n2487 = ~pi267 & ~pi503;
  assign n2488 = ~n2486 & ~n2487;
  assign n2489 = pi529 & n2488;
  assign n2490 = ~n2092 & ~n2297;
  assign n2491 = pi069 & ~n2490;
  assign n2492 = ~n2351 & ~n2491;
  assign n2493 = n2266 & ~n2492;
  assign n2494 = ~n2459 & ~n2493;
  assign n2495 = ~n2346 & n2494;
  assign n2496 = ~pi069 & n2104;
  assign n2497 = ~n2437 & ~n2496;
  assign n2498 = ~n2396 & n2497;
  assign n2499 = n2324 & ~n2498;
  assign n2500 = n2495 & ~n2499;
  assign n2501 = pi104 & n2126;
  assign n2502 = ~n2118 & ~n2247;
  assign n2503 = pi069 & n2120;
  assign n2504 = n2502 & ~n2503;
  assign n2505 = pi104 & ~n2504;
  assign n2506 = ~n2420 & ~n2505;
  assign n2507 = ~n2297 & n2506;
  assign n2508 = pi102 & ~n2507;
  assign n2509 = ~n2501 & ~n2508;
  assign n2510 = ~pi069 & n2340;
  assign n2511 = ~pi069 & n2099;
  assign n2512 = ~n2352 & ~n2511;
  assign n2513 = ~n2087 & ~n2340;
  assign n2514 = n2512 & n2513;
  assign n2515 = ~pi104 & ~n2514;
  assign n2516 = ~pi069 & n2412;
  assign n2517 = ~pi104 & n2404;
  assign n2518 = ~n2516 & ~n2517;
  assign n2519 = n2106 & n2277;
  assign n2520 = ~n2087 & ~n2519;
  assign n2521 = ~n2405 & n2520;
  assign n2522 = n2518 & n2521;
  assign n2523 = ~pi102 & ~n2522;
  assign n2524 = ~n2351 & ~n2523;
  assign n2525 = ~n2515 & n2524;
  assign n2526 = ~n2510 & n2525;
  assign n2527 = n2509 & n2526;
  assign n2528 = pi012 & ~n2527;
  assign n2529 = n2135 & n2152;
  assign n2530 = ~pi104 & n2123;
  assign n2531 = ~n2529 & ~n2530;
  assign n2532 = pi104 & n2220;
  assign n2533 = ~pi033 & n2105;
  assign n2534 = n2120 & n2533;
  assign n2535 = ~n2461 & ~n2534;
  assign n2536 = ~pi104 & ~n2535;
  assign n2537 = ~n2123 & ~n2536;
  assign n2538 = n2099 & n2159;
  assign n2539 = ~n2462 & ~n2538;
  assign n2540 = n2537 & n2539;
  assign n2541 = ~n2532 & n2540;
  assign n2542 = ~pi102 & ~n2541;
  assign n2543 = ~n2219 & ~n2320;
  assign n2544 = ~n2112 & n2543;
  assign n2545 = ~n2309 & ~n2313;
  assign n2546 = pi104 & ~n2545;
  assign n2547 = ~pi069 & ~n2103;
  assign n2548 = pi069 & ~n2118;
  assign n2549 = ~n2547 & ~n2548;
  assign n2550 = ~pi127 & n2250;
  assign n2551 = ~n2549 & ~n2550;
  assign n2552 = ~pi104 & ~n2551;
  assign n2553 = ~n2546 & ~n2552;
  assign n2554 = n2544 & n2553;
  assign n2555 = pi102 & ~n2554;
  assign n2556 = ~n2542 & ~n2555;
  assign n2557 = ~n2396 & n2556;
  assign n2558 = n2531 & n2557;
  assign n2559 = ~pi069 & n2140;
  assign n2560 = ~pi126 & n2105;
  assign n2561 = ~n2559 & ~n2560;
  assign n2562 = pi104 & ~n2561;
  assign n2563 = pi069 & n2340;
  assign n2564 = pi104 & n2563;
  assign n2565 = ~n2562 & ~n2564;
  assign n2566 = n2558 & n2565;
  assign n2567 = ~pi012 & ~n2566;
  assign n2568 = ~pi127 & n2140;
  assign n2569 = ~n2372 & ~n2568;
  assign n2570 = ~pi069 & n2110;
  assign n2571 = ~n2097 & ~n2570;
  assign n2572 = n2569 & n2571;
  assign n2573 = ~pi104 & ~n2572;
  assign n2574 = n2140 & n2388;
  assign n2575 = ~n2573 & ~n2574;
  assign n2576 = pi102 & ~n2575;
  assign n2577 = ~n2337 & ~n2356;
  assign n2578 = ~n2206 & n2577;
  assign n2579 = ~pi104 & ~n2578;
  assign n2580 = ~n2395 & ~n2579;
  assign n2581 = ~n2563 & n2580;
  assign n2582 = ~pi102 & ~n2581;
  assign n2583 = ~n2576 & ~n2582;
  assign n2584 = ~n2567 & n2583;
  assign n2585 = ~n2528 & n2584;
  assign n2586 = n2500 & n2585;
  assign n2587 = ~pi267 & ~n2586;
  assign n2588 = pi267 & n2586;
  assign n2589 = ~n2587 & ~n2588;
  assign n2590 = pi014 & n1510;
  assign n2591 = ~n1652 & ~n2590;
  assign n2592 = ~n1524 & ~n1542;
  assign n2593 = ~n1707 & n2592;
  assign n2594 = ~pi083 & ~n2593;
  assign n2595 = n2591 & ~n2594;
  assign n2596 = ~pi040 & ~n2595;
  assign n2597 = ~pi014 & n1596;
  assign n2598 = ~n1730 & ~n2597;
  assign n2599 = ~n1664 & n2598;
  assign n2600 = n1491 & ~n2599;
  assign n2601 = ~n2596 & ~n2600;
  assign n2602 = ~n1515 & ~n1687;
  assign n2603 = ~n1496 & ~n1614;
  assign n2604 = pi014 & ~n2603;
  assign n2605 = ~n1533 & ~n2604;
  assign n2606 = n1587 & ~n2605;
  assign n2607 = ~pi014 & n1570;
  assign n2608 = ~pi014 & n1509;
  assign n2609 = ~n1483 & ~n1514;
  assign n2610 = ~n2608 & n2609;
  assign n2611 = ~n2607 & n2610;
  assign n2612 = ~pi083 & ~n2611;
  assign n2613 = n1486 & n1693;
  assign n2614 = ~n2612 & ~n2613;
  assign n2615 = pi040 & ~n2614;
  assign n2616 = ~n2606 & ~n2615;
  assign n2617 = n2602 & n2616;
  assign n2618 = pi083 & n2590;
  assign n2619 = ~n1468 & ~n1477;
  assign n2620 = pi083 & ~n2619;
  assign n2621 = ~pi014 & ~n1528;
  assign n2622 = pi014 & ~n1519;
  assign n2623 = ~n2621 & ~n2622;
  assign n2624 = ~pi107 & n1556;
  assign n2625 = ~n2623 & ~n2624;
  assign n2626 = ~pi083 & ~n2625;
  assign n2627 = ~n2620 & ~n2626;
  assign n2628 = pi014 & n1701;
  assign n2629 = ~n1613 & ~n2628;
  assign n2630 = ~n1499 & n2629;
  assign n2631 = n2627 & n2630;
  assign n2632 = pi040 & ~n2631;
  assign n2633 = ~pi014 & n1486;
  assign n2634 = ~pi107 & ~pi108;
  assign n2635 = ~pi014 & n2634;
  assign n2636 = ~n2633 & ~n2635;
  assign n2637 = pi083 & ~n2636;
  assign n2638 = ~n2632 & ~n2637;
  assign n2639 = ~n2618 & n2638;
  assign n2640 = pi083 & n1641;
  assign n2641 = pi014 & n1606;
  assign n2642 = ~pi072 & n1665;
  assign n2643 = n1466 & n2642;
  assign n2644 = ~n1680 & ~n2643;
  assign n2645 = ~pi083 & ~n2644;
  assign n2646 = ~n2641 & ~n2645;
  assign n2647 = n1482 & n1517;
  assign n2648 = ~n1681 & ~n2647;
  assign n2649 = n2646 & n2648;
  assign n2650 = ~n2640 & n2649;
  assign n2651 = ~pi040 & ~n2650;
  assign n2652 = ~n1630 & ~n2641;
  assign n2653 = ~pi083 & ~n2652;
  assign n2654 = ~n2651 & ~n2653;
  assign n2655 = ~n1664 & n2654;
  assign n2656 = n2639 & n2655;
  assign n2657 = ~pi078 & ~n2656;
  assign n2658 = pi083 & n1653;
  assign n2659 = pi014 & pi107;
  assign n2660 = n1463 & n2659;
  assign n2661 = ~n1605 & ~n2660;
  assign n2662 = ~n1673 & n2661;
  assign n2663 = ~pi014 & n1699;
  assign n2664 = ~pi083 & n1672;
  assign n2665 = ~n2663 & ~n2664;
  assign n2666 = n2662 & n2665;
  assign n2667 = ~pi040 & ~n2666;
  assign n2668 = ~pi014 & n1482;
  assign n2669 = ~n1530 & ~n2668;
  assign n2670 = ~n1605 & n2669;
  assign n2671 = ~n1510 & n2670;
  assign n2672 = ~pi083 & ~n2671;
  assign n2673 = ~pi014 & n1510;
  assign n2674 = ~n2672 & ~n2673;
  assign n2675 = ~n2667 & n2674;
  assign n2676 = ~n2658 & n2675;
  assign n2677 = ~n1533 & n2676;
  assign n2678 = ~n1614 & ~n1723;
  assign n2679 = ~n1472 & ~n1519;
  assign n2680 = pi014 & n1466;
  assign n2681 = n2679 & ~n2680;
  assign n2682 = pi083 & ~n2681;
  assign n2683 = n2678 & ~n2682;
  assign n2684 = pi040 & ~n2683;
  assign n2685 = n2677 & ~n2684;
  assign n2686 = pi078 & ~n2685;
  assign n2687 = ~n2657 & ~n2686;
  assign n2688 = n2617 & n2687;
  assign n2689 = n2601 & n2688;
  assign n2690 = pi123 & n2006;
  assign n2691 = n1982 & n1995;
  assign n2692 = ~n2690 & ~n2691;
  assign n2693 = ~pi048 & pi123;
  assign n2694 = ~pi027 & n1955;
  assign n2695 = ~pi027 & n1929;
  assign n2696 = ~n2694 & ~n2695;
  assign n2697 = pi023 & n1991;
  assign n2698 = ~pi027 & n2697;
  assign n2699 = n2696 & ~n2698;
  assign n2700 = n2693 & ~n2699;
  assign n2701 = pi023 & n1918;
  assign n2702 = pi027 & n2701;
  assign n2703 = ~n2006 & ~n2702;
  assign n2704 = pi027 & n1976;
  assign n2705 = pi027 & n2041;
  assign n2706 = ~n2704 & ~n2705;
  assign n2707 = ~n2050 & n2706;
  assign n2708 = ~pi123 & ~n2707;
  assign n2709 = n2703 & ~n2708;
  assign n2710 = ~pi048 & ~n2709;
  assign n2711 = ~n2700 & ~n2710;
  assign n2712 = n2692 & n2711;
  assign n2713 = ~pi027 & n2013;
  assign n2714 = ~pi023 & n1938;
  assign n2715 = ~n1995 & ~n2714;
  assign n2716 = ~n2011 & n2715;
  assign n2717 = ~n2713 & n2716;
  assign n2718 = ~pi123 & ~n2717;
  assign n2719 = pi048 & n2718;
  assign n2720 = pi048 & pi123;
  assign n2721 = ~pi023 & n1951;
  assign n2722 = ~n1960 & ~n2721;
  assign n2723 = pi027 & ~n2722;
  assign n2724 = ~n1953 & ~n2723;
  assign n2725 = n2720 & ~n2724;
  assign n2726 = pi027 & pi048;
  assign n2727 = ~pi123 & n1923;
  assign n2728 = n2726 & n2727;
  assign n2729 = ~n2725 & ~n2728;
  assign n2730 = ~n2719 & n2729;
  assign n2731 = ~n2010 & ~n2067;
  assign n2732 = pi027 & n1923;
  assign n2733 = n2731 & ~n2732;
  assign n2734 = ~pi027 & ~n1928;
  assign n2735 = pi027 & ~n2019;
  assign n2736 = ~n2734 & ~n2735;
  assign n2737 = ~pi047 & ~pi111;
  assign n2738 = ~pi023 & n2737;
  assign n2739 = ~n2736 & ~n2738;
  assign n2740 = ~pi123 & ~n2739;
  assign n2741 = pi023 & n2038;
  assign n2742 = ~pi027 & n1991;
  assign n2743 = ~n2741 & ~n2742;
  assign n2744 = pi123 & ~n2743;
  assign n2745 = ~n2740 & ~n2744;
  assign n2746 = n2733 & n2745;
  assign n2747 = pi048 & ~n2746;
  assign n2748 = pi023 & n1976;
  assign n2749 = ~pi027 & n2721;
  assign n2750 = ~n2748 & ~n2749;
  assign n2751 = ~pi123 & ~n2750;
  assign n2752 = n1972 & n1976;
  assign n2753 = pi123 & n2068;
  assign n2754 = ~n2752 & ~n2753;
  assign n2755 = ~n2021 & n2754;
  assign n2756 = ~n2751 & n2755;
  assign n2757 = pi123 & n1962;
  assign n2758 = n2756 & ~n2757;
  assign n2759 = ~pi048 & ~n2758;
  assign n2760 = n1982 & n2701;
  assign n2761 = ~pi023 & ~pi093;
  assign n2762 = ~pi027 & n2761;
  assign n2763 = ~pi027 & n1923;
  assign n2764 = ~n2762 & ~n2763;
  assign n2765 = pi123 & ~n2764;
  assign n2766 = ~pi027 & n1932;
  assign n2767 = ~n2021 & ~n2766;
  assign n2768 = ~pi123 & ~n2767;
  assign n2769 = ~n2765 & ~n2768;
  assign n2770 = ~n2694 & n2769;
  assign n2771 = ~n2760 & n2770;
  assign n2772 = ~n2759 & n2771;
  assign n2773 = ~n2747 & n2772;
  assign n2774 = ~pi020 & ~n2773;
  assign n2775 = ~pi027 & n2701;
  assign n2776 = pi027 & n1931;
  assign n2777 = ~n1962 & ~n2776;
  assign n2778 = ~n1977 & ~n2701;
  assign n2779 = n2777 & n2778;
  assign n2780 = ~pi123 & ~n2779;
  assign n2781 = ~pi023 & n1931;
  assign n2782 = ~pi027 & n2781;
  assign n2783 = pi027 & n1928;
  assign n2784 = ~pi123 & n2783;
  assign n2785 = ~n2782 & ~n2784;
  assign n2786 = pi023 & n2783;
  assign n2787 = ~pi093 & pi111;
  assign n2788 = n1972 & n2787;
  assign n2789 = ~n1977 & ~n2788;
  assign n2790 = ~n2786 & n2789;
  assign n2791 = n2785 & n2790;
  assign n2792 = ~pi048 & ~n2791;
  assign n2793 = ~n1953 & ~n2792;
  assign n2794 = ~n2780 & n2793;
  assign n2795 = ~n2775 & n2794;
  assign n2796 = pi123 & n2023;
  assign n2797 = pi027 & n2697;
  assign n2798 = ~n2721 & ~n2797;
  assign n2799 = ~pi023 & n1944;
  assign n2800 = ~n2019 & ~n2799;
  assign n2801 = pi027 & n1950;
  assign n2802 = n2800 & ~n2801;
  assign n2803 = pi123 & ~n2802;
  assign n2804 = n2798 & ~n2803;
  assign n2805 = pi048 & ~n2804;
  assign n2806 = ~n2796 & ~n2805;
  assign n2807 = n2795 & n2806;
  assign n2808 = pi020 & ~n2807;
  assign n2809 = ~n2774 & ~n2808;
  assign n2810 = n2730 & n2809;
  assign n2811 = n2712 & n2810;
  assign n2812 = ~n2689 & n2811;
  assign n2813 = n2689 & ~n2811;
  assign n2814 = ~n2812 & ~n2813;
  assign n2815 = ~n2589 & n2814;
  assign n2816 = n2589 & ~n2814;
  assign n2817 = ~n2815 & ~n2816;
  assign n2818 = ~n1766 & ~n1848;
  assign n2819 = ~pi114 & ~n2818;
  assign n2820 = pi054 & ~pi098;
  assign n2821 = ~pi007 & n2820;
  assign n2822 = ~pi013 & n2821;
  assign n2823 = ~pi013 & n1823;
  assign n2824 = ~n2822 & ~n2823;
  assign n2825 = ~pi114 & ~n2824;
  assign n2826 = ~n2819 & ~n2825;
  assign n2827 = pi013 & pi114;
  assign n2828 = ~pi007 & n1765;
  assign n2829 = n2827 & n2828;
  assign n2830 = pi007 & n1803;
  assign n2831 = pi007 & n1823;
  assign n2832 = ~n2830 & ~n2831;
  assign n2833 = n2827 & ~n2832;
  assign n2834 = ~n2829 & ~n2833;
  assign n2835 = ~pi007 & pi098;
  assign n2836 = ~pi114 & n2835;
  assign n2837 = pi013 & n1897;
  assign n2838 = ~n2836 & ~n2837;
  assign n2839 = ~pi001 & ~n2838;
  assign n2840 = n1807 & n2827;
  assign n2841 = ~n1788 & ~n2840;
  assign n2842 = ~pi001 & ~n2841;
  assign n2843 = ~n2839 & ~n2842;
  assign n2844 = n2834 & n2843;
  assign n2845 = pi013 & n1777;
  assign n2846 = ~n1759 & ~n2845;
  assign n2847 = pi007 & n1882;
  assign n2848 = pi013 & n1862;
  assign n2849 = ~n2847 & ~n2848;
  assign n2850 = ~pi114 & ~n2849;
  assign n2851 = n1805 & n1849;
  assign n2852 = ~n2850 & ~n2851;
  assign n2853 = n2846 & n2852;
  assign n2854 = pi001 & ~n2853;
  assign n2855 = n2844 & ~n2854;
  assign n2856 = n2826 & n2855;
  assign n2857 = ~pi029 & n2856;
  assign n2858 = ~pi114 & n1815;
  assign n2859 = ~pi013 & n1899;
  assign n2860 = pi007 & n1835;
  assign n2861 = ~pi013 & n2860;
  assign n2862 = ~n2859 & ~n2861;
  assign n2863 = ~n1847 & n2862;
  assign n2864 = pi114 & ~n2863;
  assign n2865 = n1877 & n2820;
  assign n2866 = n1762 & n2827;
  assign n2867 = ~n2865 & ~n2866;
  assign n2868 = ~n2864 & n2867;
  assign n2869 = ~pi021 & ~pi054;
  assign n2870 = pi007 & n2869;
  assign n2871 = ~n1786 & ~n2870;
  assign n2872 = ~n1771 & n2871;
  assign n2873 = ~pi114 & ~n2872;
  assign n2874 = ~pi114 & n1792;
  assign n2875 = ~pi007 & n1806;
  assign n2876 = ~pi013 & n2875;
  assign n2877 = pi114 & n2876;
  assign n2878 = ~pi013 & n1770;
  assign n2879 = ~pi114 & n2878;
  assign n2880 = ~n2877 & ~n2879;
  assign n2881 = ~n2874 & n2880;
  assign n2882 = ~n2873 & n2881;
  assign n2883 = ~n1815 & ~n1837;
  assign n2884 = n2882 & n2883;
  assign n2885 = ~pi001 & ~n2884;
  assign n2886 = pi001 & pi114;
  assign n2887 = ~pi013 & n1764;
  assign n2888 = ~n2870 & ~n2887;
  assign n2889 = pi013 & n1770;
  assign n2890 = ~pi007 & pi021;
  assign n2891 = ~n2889 & ~n2890;
  assign n2892 = n2888 & n2891;
  assign n2893 = n2886 & ~n2892;
  assign n2894 = n1775 & n1791;
  assign n2895 = ~n1819 & ~n2894;
  assign n2896 = pi001 & ~n2895;
  assign n2897 = ~n2893 & ~n2896;
  assign n2898 = ~n2885 & n2897;
  assign n2899 = n2868 & n2898;
  assign n2900 = ~n2858 & n2899;
  assign n2901 = pi029 & n2900;
  assign n2902 = ~n2857 & ~n2901;
  assign n2903 = pi054 & n1802;
  assign n2904 = n1770 & n2903;
  assign n2905 = ~n1767 & ~n2904;
  assign n2906 = ~pi114 & ~n2905;
  assign n2907 = pi013 & n2875;
  assign n2908 = ~pi114 & n2907;
  assign n2909 = ~n2825 & ~n2908;
  assign n2910 = pi007 & n1896;
  assign n2911 = ~pi013 & n2910;
  assign n2912 = n2909 & ~n2911;
  assign n2913 = ~pi001 & ~n2912;
  assign n2914 = ~pi001 & pi114;
  assign n2915 = ~pi013 & n1786;
  assign n2916 = ~n1819 & ~n2915;
  assign n2917 = pi013 & n1765;
  assign n2918 = n2916 & ~n2917;
  assign n2919 = n2914 & ~n2918;
  assign n2920 = ~n2913 & ~n2919;
  assign n2921 = ~n2906 & n2920;
  assign n2922 = ~pi007 & n1757;
  assign n2923 = ~n1841 & ~n2922;
  assign n2924 = ~n1869 & ~n1899;
  assign n2925 = ~n1872 & n2924;
  assign n2926 = ~pi013 & ~n2925;
  assign n2927 = n2923 & ~n2926;
  assign n2928 = pi114 & ~n2927;
  assign n2929 = ~n1824 & ~n1863;
  assign n2930 = ~n2860 & n2929;
  assign n2931 = pi013 & ~n2930;
  assign n2932 = ~n1817 & ~n2931;
  assign n2933 = ~pi114 & ~n2932;
  assign n2934 = ~n2928 & ~n2933;
  assign n2935 = pi001 & ~n2934;
  assign n2936 = n2921 & ~n2935;
  assign n2937 = ~n2902 & n2936;
  assign n2938 = ~pi013 & ~n2929;
  assign n2939 = ~n1903 & ~n2938;
  assign n2940 = ~pi001 & ~n2939;
  assign n2941 = ~pi013 & n1896;
  assign n2942 = ~n1777 & ~n2941;
  assign n2943 = n2914 & ~n2942;
  assign n2944 = ~n2940 & ~n2943;
  assign n2945 = ~pi007 & pi013;
  assign n2946 = ~n1761 & ~n1803;
  assign n2947 = n2945 & ~n2946;
  assign n2948 = pi114 & n2947;
  assign n2949 = pi114 & n1841;
  assign n2950 = n1791 & n1806;
  assign n2951 = ~n1794 & ~n2887;
  assign n2952 = pi013 & n1756;
  assign n2953 = pi007 & n2952;
  assign n2954 = n2951 & ~n2953;
  assign n2955 = ~n2950 & n2954;
  assign n2956 = ~n2949 & n2955;
  assign n2957 = pi001 & ~n2956;
  assign n2958 = ~pi007 & n2869;
  assign n2959 = ~pi013 & n2958;
  assign n2960 = pi013 & n1823;
  assign n2961 = ~pi013 & n1778;
  assign n2962 = ~n2960 & ~n2961;
  assign n2963 = ~n2959 & n2962;
  assign n2964 = ~pi114 & ~n2963;
  assign n2965 = ~n2957 & ~n2964;
  assign n2966 = ~n2948 & n2965;
  assign n2967 = n2944 & n2966;
  assign n2968 = ~pi029 & ~n2967;
  assign n2969 = ~pi013 & n1792;
  assign n2970 = ~n1830 & ~n2969;
  assign n2971 = ~n2831 & ~n2865;
  assign n2972 = ~pi114 & ~n2971;
  assign n2973 = pi054 & n1838;
  assign n2974 = n1764 & n2973;
  assign n2975 = ~n2961 & ~n2974;
  assign n2976 = ~n2837 & n2975;
  assign n2977 = ~n1776 & n2976;
  assign n2978 = pi114 & ~n2977;
  assign n2979 = ~pi114 & n1765;
  assign n2980 = pi007 & n1862;
  assign n2981 = ~pi114 & n1785;
  assign n2982 = ~n2980 & ~n2981;
  assign n2983 = ~n2979 & n2982;
  assign n2984 = pi001 & ~n2983;
  assign n2985 = ~pi013 & n1765;
  assign n2986 = ~n1847 & ~n2985;
  assign n2987 = ~n1758 & n2986;
  assign n2988 = pi114 & ~n2987;
  assign n2989 = pi013 & n1867;
  assign n2990 = pi013 & ~pi054;
  assign n2991 = ~pi007 & n2990;
  assign n2992 = ~n2822 & ~n2991;
  assign n2993 = ~n2989 & n2992;
  assign n2994 = n1791 & n1872;
  assign n2995 = n2993 & ~n2994;
  assign n2996 = ~n2988 & n2995;
  assign n2997 = ~pi001 & ~n2996;
  assign n2998 = ~pi007 & ~pi098;
  assign n2999 = pi013 & n2998;
  assign n3000 = pi013 & n1761;
  assign n3001 = ~n2999 & ~n3000;
  assign n3002 = ~pi114 & ~n3001;
  assign n3003 = ~n2997 & ~n3002;
  assign n3004 = ~n2984 & n3003;
  assign n3005 = ~n2978 & n3004;
  assign n3006 = ~n2972 & n3005;
  assign n3007 = n2970 & n3006;
  assign n3008 = pi029 & ~n3007;
  assign n3009 = ~n2968 & ~n3008;
  assign n3010 = pi114 & ~n2904;
  assign n3011 = ~pi114 & ~n2953;
  assign n3012 = ~n3010 & ~n3011;
  assign n3013 = pi114 & n1881;
  assign n3014 = n1862 & n1877;
  assign n3015 = pi114 & ~n3014;
  assign n3016 = ~pi114 & ~n2911;
  assign n3017 = ~n3015 & ~n3016;
  assign n3018 = ~n1870 & ~n3017;
  assign n3019 = ~n3013 & n3018;
  assign n3020 = ~n1827 & n3019;
  assign n3021 = pi001 & ~n3020;
  assign n3022 = ~n3012 & ~n3021;
  assign n3023 = ~pi013 & n1862;
  assign n3024 = ~n1804 & ~n3023;
  assign n3025 = ~n1815 & n3024;
  assign n3026 = ~pi114 & ~n3025;
  assign n3027 = ~pi114 & n2945;
  assign n3028 = pi054 & n3027;
  assign n3029 = n1770 & n3028;
  assign n3030 = pi114 & n2974;
  assign n3031 = n1775 & n1802;
  assign n3032 = n1785 & n1802;
  assign n3033 = ~n3031 & ~n3032;
  assign n3034 = pi114 & ~n3033;
  assign n3035 = ~n3030 & ~n3034;
  assign n3036 = ~n3029 & n3035;
  assign n3037 = ~n3026 & n3036;
  assign n3038 = ~pi001 & ~n3037;
  assign n3039 = n3022 & ~n3038;
  assign n3040 = n3009 & n3039;
  assign n3041 = ~n2937 & n3040;
  assign n3042 = n2937 & ~n3040;
  assign n3043 = ~n3041 & ~n3042;
  assign n3044 = ~n1918 & ~n1920;
  assign n3045 = n2032 & ~n3044;
  assign n3046 = pi123 & n3045;
  assign n3047 = ~pi027 & n2038;
  assign n3048 = ~n1931 & ~n3047;
  assign n3049 = n2693 & ~n3048;
  assign n3050 = ~n3046 & ~n3049;
  assign n3051 = ~pi027 & ~pi123;
  assign n3052 = n1944 & n3051;
  assign n3053 = n1950 & n1972;
  assign n3054 = pi123 & n2010;
  assign n3055 = ~n3053 & ~n3054;
  assign n3056 = ~n3052 & n3055;
  assign n3057 = ~pi027 & n1917;
  assign n3058 = ~n1955 & ~n3057;
  assign n3059 = n3056 & n3058;
  assign n3060 = pi048 & ~n3059;
  assign n3061 = n3050 & ~n3060;
  assign n3062 = ~n1977 & ~n1992;
  assign n3063 = ~pi027 & ~n3062;
  assign n3064 = ~n2037 & ~n3063;
  assign n3065 = ~pi048 & ~n3064;
  assign n3066 = ~pi027 & n2738;
  assign n3067 = ~n2766 & ~n3066;
  assign n3068 = pi027 & n1991;
  assign n3069 = n3067 & ~n3068;
  assign n3070 = ~pi123 & ~n3069;
  assign n3071 = ~n3065 & ~n3070;
  assign n3072 = n3061 & n3071;
  assign n3073 = ~pi020 & ~n3072;
  assign n3074 = ~n1962 & ~n1988;
  assign n3075 = ~n2702 & ~n2705;
  assign n3076 = ~n2766 & n3075;
  assign n3077 = ~n1930 & n3076;
  assign n3078 = pi123 & ~n3077;
  assign n3079 = pi023 & ~pi027;
  assign n3080 = n2787 & n3079;
  assign n3081 = ~n2697 & ~n3080;
  assign n3082 = ~pi123 & ~n3081;
  assign n3083 = ~n3078 & ~n3082;
  assign n3084 = pi027 & n1920;
  assign n3085 = pi027 & n2761;
  assign n3086 = ~n3084 & ~n3085;
  assign n3087 = ~pi123 & ~n3086;
  assign n3088 = pi027 & ~pi111;
  assign n3089 = ~pi023 & n3088;
  assign n3090 = pi027 & n2054;
  assign n3091 = ~n3089 & ~n3090;
  assign n3092 = ~pi023 & n2787;
  assign n3093 = ~pi027 & n3092;
  assign n3094 = n3091 & ~n3093;
  assign n3095 = n2005 & n3051;
  assign n3096 = ~n2003 & ~n2763;
  assign n3097 = ~n1952 & n3096;
  assign n3098 = pi123 & ~n3097;
  assign n3099 = ~n3095 & ~n3098;
  assign n3100 = n3094 & n3099;
  assign n3101 = ~pi048 & ~n3100;
  assign n3102 = ~n3087 & ~n3101;
  assign n3103 = ~pi123 & n1959;
  assign n3104 = ~n2727 & ~n3103;
  assign n3105 = ~n2748 & n3104;
  assign n3106 = pi048 & ~n3105;
  assign n3107 = n3102 & ~n3106;
  assign n3108 = n3083 & n3107;
  assign n3109 = n3074 & n3108;
  assign n3110 = pi020 & ~n3109;
  assign n3111 = ~pi027 & n2714;
  assign n3112 = pi123 & n3111;
  assign n3113 = ~pi123 & n3053;
  assign n3114 = n1916 & n1959;
  assign n3115 = ~n2008 & ~n3114;
  assign n3116 = n2693 & ~n3115;
  assign n3117 = ~n3113 & ~n3116;
  assign n3118 = ~n3112 & n3117;
  assign n3119 = ~pi027 & n1976;
  assign n3120 = ~n1919 & ~n3119;
  assign n3121 = ~n1980 & n3120;
  assign n3122 = ~pi123 & ~n3121;
  assign n3123 = pi027 & n2714;
  assign n3124 = ~pi123 & n3123;
  assign n3125 = ~n3122 & ~n3124;
  assign n3126 = ~n2760 & n3125;
  assign n3127 = ~pi048 & ~n3126;
  assign n3128 = ~n1996 & ~n2052;
  assign n3129 = pi123 & n3079;
  assign n3130 = n1976 & n3129;
  assign n3131 = pi123 & n2031;
  assign n3132 = ~pi027 & n2741;
  assign n3133 = ~pi123 & n3132;
  assign n3134 = ~n3131 & ~n3133;
  assign n3135 = ~n3130 & n3134;
  assign n3136 = n3128 & n3135;
  assign n3137 = pi048 & ~n3136;
  assign n3138 = ~n3127 & ~n3137;
  assign n3139 = n3118 & n3138;
  assign n3140 = ~n3110 & n3139;
  assign n3141 = ~n3073 & n3140;
  assign n3142 = ~n2742 & ~n3093;
  assign n3143 = ~pi123 & ~n3142;
  assign n3144 = ~n1924 & ~n2004;
  assign n3145 = ~pi123 & ~n3144;
  assign n3146 = ~n3143 & ~n3145;
  assign n3147 = n1945 & n1982;
  assign n3148 = ~n1957 & ~n3147;
  assign n3149 = ~pi048 & ~n3148;
  assign n3150 = ~n2697 & ~n2701;
  assign n3151 = n1982 & ~n3150;
  assign n3152 = ~n3149 & ~n3151;
  assign n3153 = ~n2691 & n3152;
  assign n3154 = ~pi023 & pi093;
  assign n3155 = ~pi123 & n3154;
  assign n3156 = ~n2705 & ~n3155;
  assign n3157 = ~pi048 & ~n3156;
  assign n3158 = n3153 & ~n3157;
  assign n3159 = ~n1953 & ~n2776;
  assign n3160 = ~pi047 & n1972;
  assign n3161 = ~n2704 & ~n3160;
  assign n3162 = ~pi123 & ~n3161;
  assign n3163 = n1943 & n2019;
  assign n3164 = ~n3162 & ~n3163;
  assign n3165 = n3159 & n3164;
  assign n3166 = pi048 & ~n3165;
  assign n3167 = n3158 & ~n3166;
  assign n3168 = n3146 & n3167;
  assign n3169 = ~pi020 & n3168;
  assign n3170 = ~pi123 & n1938;
  assign n3171 = ~pi027 & n2799;
  assign n3172 = pi123 & n3171;
  assign n3173 = ~pi027 & n1937;
  assign n3174 = ~pi123 & n3173;
  assign n3175 = ~n3172 & ~n3174;
  assign n3176 = ~n3170 & n3175;
  assign n3177 = pi023 & n2737;
  assign n3178 = ~n1960 & ~n3177;
  assign n3179 = ~n1940 & n3178;
  assign n3180 = ~pi123 & ~n3179;
  assign n3181 = n3176 & ~n3180;
  assign n3182 = ~n1980 & ~n2014;
  assign n3183 = n3181 & n3182;
  assign n3184 = ~pi048 & ~n3183;
  assign n3185 = ~pi023 & pi047;
  assign n3186 = pi027 & n1937;
  assign n3187 = ~n3057 & ~n3177;
  assign n3188 = ~n3186 & n3187;
  assign n3189 = ~n3185 & n3188;
  assign n3190 = n2720 & ~n3189;
  assign n3191 = ~n3080 & ~n3190;
  assign n3192 = pi020 & n3191;
  assign n3193 = ~pi123 & n1980;
  assign n3194 = n3192 & ~n3193;
  assign n3195 = n1921 & n1982;
  assign n3196 = pi023 & n2012;
  assign n3197 = ~pi027 & n3196;
  assign n3198 = ~pi027 & n2043;
  assign n3199 = ~n2003 & ~n3198;
  assign n3200 = ~n3197 & n3199;
  assign n3201 = pi123 & ~n3200;
  assign n3202 = ~n3195 & ~n3201;
  assign n3203 = n1929 & n3051;
  assign n3204 = ~n2000 & ~n3203;
  assign n3205 = pi048 & ~n3204;
  assign n3206 = n3202 & ~n3205;
  assign n3207 = n3194 & n3206;
  assign n3208 = ~n3184 & n3207;
  assign n3209 = ~n3169 & ~n3208;
  assign n3210 = ~n1925 & ~n3111;
  assign n3211 = ~pi123 & ~n3210;
  assign n3212 = pi027 & n2799;
  assign n3213 = ~pi123 & n3212;
  assign n3214 = ~n3143 & ~n3213;
  assign n3215 = ~n3132 & n3214;
  assign n3216 = ~pi048 & ~n3215;
  assign n3217 = ~pi027 & n1960;
  assign n3218 = ~n2000 & ~n3217;
  assign n3219 = ~n2732 & n3218;
  assign n3220 = n2693 & ~n3219;
  assign n3221 = ~n3216 & ~n3220;
  assign n3222 = ~n3211 & n3221;
  assign n3223 = ~n2010 & ~n2721;
  assign n3224 = ~n2005 & ~n2051;
  assign n3225 = ~n2043 & n3224;
  assign n3226 = ~pi027 & ~n3225;
  assign n3227 = n3223 & ~n3226;
  assign n3228 = pi123 & ~n3227;
  assign n3229 = pi027 & n1918;
  assign n3230 = ~n1977 & ~n3196;
  assign n3231 = ~n1992 & n3230;
  assign n3232 = pi027 & ~n3231;
  assign n3233 = ~n3229 & ~n3232;
  assign n3234 = ~pi123 & ~n3233;
  assign n3235 = ~n3228 & ~n3234;
  assign n3236 = pi048 & ~n3235;
  assign n3237 = n3222 & ~n3236;
  assign n3238 = ~n3209 & n3237;
  assign n3239 = ~n3141 & n3238;
  assign n3240 = n3141 & ~n3238;
  assign n3241 = ~n3239 & ~n3240;
  assign n3242 = ~n3043 & n3241;
  assign n3243 = n2937 & n3040;
  assign n3244 = ~n2937 & ~n3040;
  assign n3245 = ~n3243 & ~n3244;
  assign n3246 = ~n3241 & ~n3245;
  assign n3247 = ~n3242 & ~n3246;
  assign n3248 = n2817 & n3247;
  assign n3249 = ~n2817 & ~n3247;
  assign n3250 = ~n3248 & ~n3249;
  assign n3251 = ~pi529 & n3250;
  assign po131 = n2489 | n3251;
  assign n3253 = ~pi268 & pi527;
  assign n3254 = pi268 & ~pi527;
  assign n3255 = ~n3253 & ~n3254;
  assign n3256 = pi529 & n3255;
  assign n3257 = pi073 & pi080;
  assign n3258 = pi042 & pi110;
  assign n3259 = ~pi071 & n3258;
  assign n3260 = pi075 & n3259;
  assign n3261 = ~pi079 & n3260;
  assign n3262 = ~pi075 & n3259;
  assign n3263 = pi042 & pi071;
  assign n3264 = pi075 & n3263;
  assign n3265 = ~n3262 & ~n3264;
  assign n3266 = pi079 & ~n3265;
  assign n3267 = ~n3261 & ~n3266;
  assign n3268 = n3257 & ~n3267;
  assign n3269 = ~pi042 & ~pi110;
  assign n3270 = ~pi071 & n3269;
  assign n3271 = ~pi075 & n3270;
  assign n3272 = ~pi110 & n3263;
  assign n3273 = ~pi075 & n3272;
  assign n3274 = ~n3271 & ~n3273;
  assign n3275 = ~pi042 & pi071;
  assign n3276 = ~pi075 & n3275;
  assign n3277 = ~pi079 & n3276;
  assign n3278 = pi071 & n3269;
  assign n3279 = ~pi079 & n3278;
  assign n3280 = ~n3277 & ~n3279;
  assign n3281 = n3274 & n3280;
  assign n3282 = ~pi080 & ~n3281;
  assign n3283 = pi079 & ~pi080;
  assign n3284 = n3270 & n3283;
  assign n3285 = ~n3282 & ~n3284;
  assign n3286 = pi073 & ~n3285;
  assign n3287 = ~n3268 & ~n3286;
  assign n3288 = pi079 & pi080;
  assign n3289 = n3271 & n3288;
  assign n3290 = ~pi073 & pi080;
  assign n3291 = ~pi075 & n3269;
  assign n3292 = ~pi079 & n3291;
  assign n3293 = pi071 & n3258;
  assign n3294 = pi075 & n3293;
  assign n3295 = ~pi079 & n3294;
  assign n3296 = ~pi042 & pi110;
  assign n3297 = ~pi071 & n3296;
  assign n3298 = ~pi079 & n3297;
  assign n3299 = ~n3295 & ~n3298;
  assign n3300 = ~n3292 & n3299;
  assign n3301 = n3290 & ~n3300;
  assign n3302 = pi075 & pi079;
  assign n3303 = n3297 & n3302;
  assign n3304 = pi080 & n3303;
  assign n3305 = ~n3301 & ~n3304;
  assign n3306 = ~n3289 & n3305;
  assign n3307 = pi075 & n3278;
  assign n3308 = pi079 & n3307;
  assign n3309 = pi042 & ~pi110;
  assign n3310 = ~pi071 & n3309;
  assign n3311 = pi079 & n3310;
  assign n3312 = pi071 & pi110;
  assign n3313 = ~pi075 & n3312;
  assign n3314 = pi079 & n3313;
  assign n3315 = ~n3311 & ~n3314;
  assign n3316 = pi075 & n3270;
  assign n3317 = ~pi079 & n3316;
  assign n3318 = n3315 & ~n3317;
  assign n3319 = ~pi080 & ~n3318;
  assign n3320 = ~n3303 & ~n3319;
  assign n3321 = ~n3308 & n3320;
  assign n3322 = ~pi073 & ~n3321;
  assign n3323 = n3306 & ~n3322;
  assign n3324 = ~pi079 & n3307;
  assign n3325 = ~pi079 & n3272;
  assign n3326 = pi110 & n3275;
  assign n3327 = pi079 & n3326;
  assign n3328 = ~n3325 & ~n3327;
  assign n3329 = ~pi075 & n3310;
  assign n3330 = ~n3307 & ~n3329;
  assign n3331 = n3328 & n3330;
  assign n3332 = ~pi080 & ~n3331;
  assign n3333 = ~pi075 & n3326;
  assign n3334 = ~pi079 & n3333;
  assign n3335 = pi079 & n3296;
  assign n3336 = ~pi080 & n3335;
  assign n3337 = ~n3334 & ~n3336;
  assign n3338 = pi075 & n3335;
  assign n3339 = pi071 & ~pi110;
  assign n3340 = n3302 & n3339;
  assign n3341 = ~n3329 & ~n3340;
  assign n3342 = ~n3338 & n3341;
  assign n3343 = n3337 & n3342;
  assign n3344 = ~pi073 & ~n3343;
  assign n3345 = ~n3261 & ~n3344;
  assign n3346 = ~n3332 & n3345;
  assign n3347 = ~n3324 & n3346;
  assign n3348 = ~pi079 & n3259;
  assign n3349 = pi080 & n3348;
  assign n3350 = pi042 & ~pi071;
  assign n3351 = pi075 & n3350;
  assign n3352 = ~pi071 & pi110;
  assign n3353 = ~pi075 & n3352;
  assign n3354 = ~n3351 & ~n3353;
  assign n3355 = pi079 & n3258;
  assign n3356 = n3354 & ~n3355;
  assign n3357 = pi080 & ~n3356;
  assign n3358 = pi079 & n3294;
  assign n3359 = ~n3357 & ~n3358;
  assign n3360 = ~n3262 & n3359;
  assign n3361 = pi073 & ~n3360;
  assign n3362 = ~n3349 & ~n3361;
  assign n3363 = n3347 & n3362;
  assign n3364 = pi015 & ~n3363;
  assign n3365 = pi075 & n3326;
  assign n3366 = ~pi079 & ~pi080;
  assign n3367 = n3365 & n3366;
  assign n3368 = ~pi075 & n3293;
  assign n3369 = pi079 & n3368;
  assign n3370 = ~pi080 & n3369;
  assign n3371 = ~n3367 & ~n3370;
  assign n3372 = pi079 & n3272;
  assign n3373 = pi079 & n3270;
  assign n3374 = ~pi075 & n3309;
  assign n3375 = pi079 & n3374;
  assign n3376 = ~n3373 & ~n3375;
  assign n3377 = ~n3372 & n3376;
  assign n3378 = pi075 & n3312;
  assign n3379 = ~pi079 & n3293;
  assign n3380 = ~n3378 & ~n3379;
  assign n3381 = pi080 & ~n3380;
  assign n3382 = ~pi079 & ~n3296;
  assign n3383 = pi079 & ~n3351;
  assign n3384 = ~n3382 & ~n3383;
  assign n3385 = ~pi042 & ~pi071;
  assign n3386 = ~pi075 & n3385;
  assign n3387 = ~n3384 & ~n3386;
  assign n3388 = ~pi080 & ~n3387;
  assign n3389 = ~n3381 & ~n3388;
  assign n3390 = n3377 & n3389;
  assign n3391 = pi073 & ~n3390;
  assign n3392 = pi079 & n3259;
  assign n3393 = pi080 & n3392;
  assign n3394 = pi075 & n3310;
  assign n3395 = ~pi075 & ~pi079;
  assign n3396 = ~pi071 & n3395;
  assign n3397 = n3258 & n3396;
  assign n3398 = ~n3394 & ~n3397;
  assign n3399 = ~pi080 & ~n3398;
  assign n3400 = ~n3369 & ~n3399;
  assign n3401 = ~pi079 & pi080;
  assign n3402 = n3272 & n3401;
  assign n3403 = pi079 & n3394;
  assign n3404 = ~n3402 & ~n3403;
  assign n3405 = n3400 & n3404;
  assign n3406 = ~n3393 & n3405;
  assign n3407 = ~pi073 & ~n3406;
  assign n3408 = ~n3391 & ~n3407;
  assign n3409 = ~n3292 & n3408;
  assign n3410 = n3371 & n3409;
  assign n3411 = ~pi079 & n3270;
  assign n3412 = ~pi110 & n3395;
  assign n3413 = ~n3411 & ~n3412;
  assign n3414 = pi080 & ~n3413;
  assign n3415 = pi080 & n3308;
  assign n3416 = ~n3414 & ~n3415;
  assign n3417 = n3410 & n3416;
  assign n3418 = ~pi015 & ~n3417;
  assign n3419 = ~n3364 & ~n3418;
  assign n3420 = n3323 & n3419;
  assign n3421 = n3287 & n3420;
  assign n3422 = pi268 & ~n3421;
  assign n3423 = ~pi268 & n3421;
  assign n3424 = ~n3422 & ~n3423;
  assign n3425 = ~pi046 & pi050;
  assign n3426 = ~pi087 & n3425;
  assign n3427 = pi085 & n3426;
  assign n3428 = pi028 & n3427;
  assign n3429 = pi092 & n3428;
  assign n3430 = ~pi046 & ~pi050;
  assign n3431 = ~pi087 & n3430;
  assign n3432 = ~pi085 & n3431;
  assign n3433 = pi028 & pi092;
  assign n3434 = n3432 & n3433;
  assign n3435 = ~n3429 & ~n3434;
  assign n3436 = ~pi028 & ~pi085;
  assign n3437 = ~pi050 & n3436;
  assign n3438 = ~pi046 & n3437;
  assign n3439 = pi046 & pi050;
  assign n3440 = pi087 & n3439;
  assign n3441 = pi085 & n3440;
  assign n3442 = ~pi028 & n3441;
  assign n3443 = ~pi028 & n3426;
  assign n3444 = ~n3442 & ~n3443;
  assign n3445 = ~n3438 & n3444;
  assign n3446 = ~pi089 & pi092;
  assign n3447 = ~n3445 & n3446;
  assign n3448 = n3435 & ~n3447;
  assign n3449 = pi087 & n3430;
  assign n3450 = pi085 & n3449;
  assign n3451 = pi028 & n3450;
  assign n3452 = ~n3428 & ~n3451;
  assign n3453 = pi046 & ~pi050;
  assign n3454 = ~pi087 & n3453;
  assign n3455 = pi028 & n3454;
  assign n3456 = pi050 & pi087;
  assign n3457 = ~pi085 & n3456;
  assign n3458 = pi028 & n3457;
  assign n3459 = ~n3455 & ~n3458;
  assign n3460 = pi085 & n3431;
  assign n3461 = ~pi028 & n3460;
  assign n3462 = n3459 & ~n3461;
  assign n3463 = ~pi092 & ~n3462;
  assign n3464 = n3452 & ~n3463;
  assign n3465 = ~pi089 & ~n3464;
  assign n3466 = n3448 & ~n3465;
  assign n3467 = ~pi087 & n3439;
  assign n3468 = ~pi028 & pi085;
  assign n3469 = n3467 & n3468;
  assign n3470 = ~pi085 & n3467;
  assign n3471 = pi046 & pi087;
  assign n3472 = pi085 & n3471;
  assign n3473 = ~n3470 & ~n3472;
  assign n3474 = pi028 & ~n3473;
  assign n3475 = ~n3469 & ~n3474;
  assign n3476 = pi089 & pi092;
  assign n3477 = ~n3475 & n3476;
  assign n3478 = ~pi046 & pi087;
  assign n3479 = ~pi085 & n3478;
  assign n3480 = ~pi028 & n3479;
  assign n3481 = ~pi028 & n3449;
  assign n3482 = pi087 & n3453;
  assign n3483 = ~pi085 & n3482;
  assign n3484 = ~n3432 & ~n3483;
  assign n3485 = ~n3481 & n3484;
  assign n3486 = ~n3480 & n3485;
  assign n3487 = ~pi092 & ~n3486;
  assign n3488 = pi028 & ~pi092;
  assign n3489 = n3431 & n3488;
  assign n3490 = ~n3487 & ~n3489;
  assign n3491 = pi089 & ~n3490;
  assign n3492 = ~n3477 & ~n3491;
  assign n3493 = ~pi085 & n3440;
  assign n3494 = pi028 & n3493;
  assign n3495 = pi087 & n3425;
  assign n3496 = pi085 & n3495;
  assign n3497 = ~pi028 & n3496;
  assign n3498 = ~n3494 & ~n3497;
  assign n3499 = ~pi092 & ~n3498;
  assign n3500 = pi028 & n3467;
  assign n3501 = pi092 & n3500;
  assign n3502 = pi085 & n3454;
  assign n3503 = ~pi028 & n3467;
  assign n3504 = ~pi085 & n3503;
  assign n3505 = ~n3502 & ~n3504;
  assign n3506 = ~pi092 & ~n3505;
  assign n3507 = ~n3494 & ~n3506;
  assign n3508 = ~pi028 & pi092;
  assign n3509 = n3482 & n3508;
  assign n3510 = pi028 & n3502;
  assign n3511 = ~n3509 & ~n3510;
  assign n3512 = n3507 & n3511;
  assign n3513 = ~n3501 & n3512;
  assign n3514 = ~pi089 & ~n3513;
  assign n3515 = ~pi085 & n3453;
  assign n3516 = pi028 & n3515;
  assign n3517 = pi028 & n3482;
  assign n3518 = ~n3516 & ~n3517;
  assign n3519 = pi028 & n3431;
  assign n3520 = n3518 & ~n3519;
  assign n3521 = pi085 & n3456;
  assign n3522 = ~pi028 & n3440;
  assign n3523 = ~n3521 & ~n3522;
  assign n3524 = pi092 & ~n3523;
  assign n3525 = ~pi028 & ~n3425;
  assign n3526 = pi046 & ~pi087;
  assign n3527 = pi085 & n3526;
  assign n3528 = pi028 & ~n3527;
  assign n3529 = ~n3525 & ~n3528;
  assign n3530 = ~pi046 & ~pi087;
  assign n3531 = ~pi085 & n3530;
  assign n3532 = ~n3529 & ~n3531;
  assign n3533 = ~pi092 & ~n3532;
  assign n3534 = ~n3524 & ~n3533;
  assign n3535 = n3520 & n3534;
  assign n3536 = pi089 & ~n3535;
  assign n3537 = ~n3514 & ~n3536;
  assign n3538 = ~n3438 & n3537;
  assign n3539 = ~n3499 & n3538;
  assign n3540 = ~pi028 & ~pi087;
  assign n3541 = ~pi050 & n3540;
  assign n3542 = ~pi046 & n3541;
  assign n3543 = ~pi050 & ~pi085;
  assign n3544 = ~pi028 & n3543;
  assign n3545 = ~n3542 & ~n3544;
  assign n3546 = pi092 & ~n3545;
  assign n3547 = pi092 & n3451;
  assign n3548 = ~n3546 & ~n3547;
  assign n3549 = n3539 & n3548;
  assign n3550 = ~pi053 & ~n3549;
  assign n3551 = pi028 & n3425;
  assign n3552 = pi085 & n3551;
  assign n3553 = ~pi085 & n3454;
  assign n3554 = pi028 & pi085;
  assign n3555 = ~pi050 & pi087;
  assign n3556 = n3554 & n3555;
  assign n3557 = ~n3553 & ~n3556;
  assign n3558 = ~n3552 & n3557;
  assign n3559 = ~pi085 & n3495;
  assign n3560 = ~pi028 & n3559;
  assign n3561 = ~pi092 & n3551;
  assign n3562 = ~n3560 & ~n3561;
  assign n3563 = n3558 & n3562;
  assign n3564 = ~pi089 & ~n3563;
  assign n3565 = ~pi028 & n3482;
  assign n3566 = pi028 & n3495;
  assign n3567 = ~n3565 & ~n3566;
  assign n3568 = ~n3553 & n3567;
  assign n3569 = ~n3450 & n3568;
  assign n3570 = ~pi092 & ~n3569;
  assign n3571 = ~pi028 & n3450;
  assign n3572 = ~n3570 & ~n3571;
  assign n3573 = pi028 & n3441;
  assign n3574 = ~n3470 & ~n3573;
  assign n3575 = pi050 & ~pi087;
  assign n3576 = ~pi085 & n3575;
  assign n3577 = ~n3527 & ~n3576;
  assign n3578 = pi028 & n3439;
  assign n3579 = n3577 & ~n3578;
  assign n3580 = pi092 & ~n3579;
  assign n3581 = n3574 & ~n3580;
  assign n3582 = pi089 & ~n3581;
  assign n3583 = pi092 & n3503;
  assign n3584 = ~n3469 & ~n3583;
  assign n3585 = ~n3582 & n3584;
  assign n3586 = n3572 & n3585;
  assign n3587 = ~n3564 & n3586;
  assign n3588 = pi053 & ~n3587;
  assign n3589 = ~n3550 & ~n3588;
  assign n3590 = n3492 & n3589;
  assign n3591 = n3466 & n3590;
  assign n3592 = ~pi026 & pi115;
  assign n3593 = ~pi056 & ~pi099;
  assign n3594 = ~pi059 & n3593;
  assign n3595 = ~pi008 & n3594;
  assign n3596 = ~pi056 & pi099;
  assign n3597 = ~pi095 & n3596;
  assign n3598 = ~pi008 & n3597;
  assign n3599 = ~n3595 & ~n3598;
  assign n3600 = pi056 & pi099;
  assign n3601 = pi095 & n3600;
  assign n3602 = pi059 & n3601;
  assign n3603 = ~pi008 & n3602;
  assign n3604 = n3599 & ~n3603;
  assign n3605 = n3592 & ~n3604;
  assign n3606 = pi059 & n3597;
  assign n3607 = pi008 & n3606;
  assign n3608 = pi115 & n3607;
  assign n3609 = pi008 & pi115;
  assign n3610 = ~pi056 & ~pi095;
  assign n3611 = ~pi099 & n3610;
  assign n3612 = ~pi059 & n3611;
  assign n3613 = n3609 & n3612;
  assign n3614 = ~n3608 & ~n3613;
  assign n3615 = ~n3605 & n3614;
  assign n3616 = pi095 & n3593;
  assign n3617 = pi059 & n3616;
  assign n3618 = ~pi008 & n3617;
  assign n3619 = pi056 & ~pi099;
  assign n3620 = pi095 & n3619;
  assign n3621 = ~pi008 & n3620;
  assign n3622 = pi095 & n3596;
  assign n3623 = pi008 & n3622;
  assign n3624 = ~n3621 & ~n3623;
  assign n3625 = ~pi095 & n3619;
  assign n3626 = ~pi059 & n3625;
  assign n3627 = ~n3617 & ~n3626;
  assign n3628 = n3624 & n3627;
  assign n3629 = ~pi115 & ~n3628;
  assign n3630 = ~pi095 & n3600;
  assign n3631 = pi059 & n3630;
  assign n3632 = ~pi008 & n3631;
  assign n3633 = ~pi059 & n3622;
  assign n3634 = ~pi008 & n3633;
  assign n3635 = pi008 & n3596;
  assign n3636 = ~pi115 & n3635;
  assign n3637 = ~n3634 & ~n3636;
  assign n3638 = pi059 & n3635;
  assign n3639 = pi008 & pi059;
  assign n3640 = pi095 & ~pi099;
  assign n3641 = n3639 & n3640;
  assign n3642 = ~n3638 & ~n3641;
  assign n3643 = ~n3626 & n3642;
  assign n3644 = n3637 & n3643;
  assign n3645 = ~pi026 & ~n3644;
  assign n3646 = ~n3632 & ~n3645;
  assign n3647 = ~n3629 & n3646;
  assign n3648 = ~n3618 & n3647;
  assign n3649 = ~pi008 & n3630;
  assign n3650 = pi115 & n3649;
  assign n3651 = ~pi059 & n3630;
  assign n3652 = pi008 & n3602;
  assign n3653 = ~n3651 & ~n3652;
  assign n3654 = pi056 & ~pi095;
  assign n3655 = pi059 & n3654;
  assign n3656 = ~pi095 & pi099;
  assign n3657 = ~pi059 & n3656;
  assign n3658 = ~n3655 & ~n3657;
  assign n3659 = pi008 & n3600;
  assign n3660 = n3658 & ~n3659;
  assign n3661 = pi115 & ~n3660;
  assign n3662 = n3653 & ~n3661;
  assign n3663 = pi026 & ~n3662;
  assign n3664 = ~n3650 & ~n3663;
  assign n3665 = n3648 & n3664;
  assign n3666 = pi030 & ~n3665;
  assign n3667 = pi059 & n3625;
  assign n3668 = ~pi008 & n3651;
  assign n3669 = ~n3667 & ~n3668;
  assign n3670 = ~pi115 & ~n3669;
  assign n3671 = ~pi059 & n3601;
  assign n3672 = pi008 & n3671;
  assign n3673 = n3625 & n3639;
  assign n3674 = pi008 & n3630;
  assign n3675 = pi115 & n3674;
  assign n3676 = ~n3673 & ~n3675;
  assign n3677 = ~n3672 & n3676;
  assign n3678 = ~n3670 & n3677;
  assign n3679 = pi115 & n3621;
  assign n3680 = n3678 & ~n3679;
  assign n3681 = ~pi026 & ~n3680;
  assign n3682 = ~pi059 & n3619;
  assign n3683 = pi008 & n3682;
  assign n3684 = pi008 & n3620;
  assign n3685 = ~n3683 & ~n3684;
  assign n3686 = pi008 & n3611;
  assign n3687 = n3685 & ~n3686;
  assign n3688 = ~pi008 & ~n3596;
  assign n3689 = pi008 & ~n3655;
  assign n3690 = ~n3688 & ~n3689;
  assign n3691 = ~pi059 & n3610;
  assign n3692 = ~n3690 & ~n3691;
  assign n3693 = ~pi115 & ~n3692;
  assign n3694 = pi095 & pi099;
  assign n3695 = pi059 & n3694;
  assign n3696 = ~pi008 & n3601;
  assign n3697 = ~n3695 & ~n3696;
  assign n3698 = pi115 & ~n3697;
  assign n3699 = ~n3693 & ~n3698;
  assign n3700 = n3687 & n3699;
  assign n3701 = pi026 & ~n3700;
  assign n3702 = ~n3681 & ~n3701;
  assign n3703 = pi059 & n3622;
  assign n3704 = ~pi008 & n3703;
  assign n3705 = ~n3672 & ~n3704;
  assign n3706 = ~pi115 & ~n3705;
  assign n3707 = ~n3595 & ~n3706;
  assign n3708 = n3609 & n3617;
  assign n3709 = ~pi059 & ~pi099;
  assign n3710 = ~pi008 & n3709;
  assign n3711 = ~pi008 & n3611;
  assign n3712 = ~n3710 & ~n3711;
  assign n3713 = pi115 & ~n3712;
  assign n3714 = ~n3708 & ~n3713;
  assign n3715 = n3707 & n3714;
  assign n3716 = n3702 & n3715;
  assign n3717 = ~pi030 & ~n3716;
  assign n3718 = ~pi056 & pi095;
  assign n3719 = ~pi059 & n3718;
  assign n3720 = ~pi008 & n3719;
  assign n3721 = ~pi008 & n3616;
  assign n3722 = ~pi059 & n3620;
  assign n3723 = ~n3612 & ~n3722;
  assign n3724 = ~n3721 & n3723;
  assign n3725 = ~n3720 & n3724;
  assign n3726 = ~pi115 & ~n3725;
  assign n3727 = pi026 & n3726;
  assign n3728 = pi026 & pi115;
  assign n3729 = pi056 & pi095;
  assign n3730 = pi059 & n3729;
  assign n3731 = ~n3651 & ~n3730;
  assign n3732 = pi008 & ~n3731;
  assign n3733 = ~n3632 & ~n3732;
  assign n3734 = n3728 & ~n3733;
  assign n3735 = pi008 & pi026;
  assign n3736 = ~pi115 & n3611;
  assign n3737 = n3735 & n3736;
  assign n3738 = ~n3734 & ~n3737;
  assign n3739 = ~n3727 & n3738;
  assign n3740 = pi008 & n3617;
  assign n3741 = ~n3607 & ~n3740;
  assign n3742 = pi008 & n3625;
  assign n3743 = ~pi059 & n3694;
  assign n3744 = pi008 & n3743;
  assign n3745 = ~n3742 & ~n3744;
  assign n3746 = pi059 & n3611;
  assign n3747 = ~pi008 & n3746;
  assign n3748 = n3745 & ~n3747;
  assign n3749 = ~pi115 & ~n3748;
  assign n3750 = n3741 & ~n3749;
  assign n3751 = ~pi026 & ~n3750;
  assign n3752 = n3739 & ~n3751;
  assign n3753 = ~n3717 & n3752;
  assign n3754 = ~n3666 & n3753;
  assign n3755 = n3615 & n3754;
  assign n3756 = ~n3591 & n3755;
  assign n3757 = n3591 & ~n3755;
  assign n3758 = ~n3756 & ~n3757;
  assign n3759 = ~n3424 & n3758;
  assign n3760 = n3424 & ~n3758;
  assign n3761 = ~n3759 & ~n3760;
  assign n3762 = pi064 & ~pi105;
  assign n3763 = ~pi032 & n3762;
  assign n3764 = ~pi067 & n3763;
  assign n3765 = pi061 & pi105;
  assign n3766 = pi064 & n3765;
  assign n3767 = ~pi067 & n3766;
  assign n3768 = ~n3764 & ~n3767;
  assign n3769 = ~pi117 & ~n3768;
  assign n3770 = ~pi064 & pi105;
  assign n3771 = ~pi032 & n3770;
  assign n3772 = pi067 & n3771;
  assign n3773 = ~pi117 & n3772;
  assign n3774 = ~n3769 & ~n3773;
  assign n3775 = pi064 & pi105;
  assign n3776 = pi032 & n3775;
  assign n3777 = ~pi067 & n3776;
  assign n3778 = n3774 & ~n3777;
  assign n3779 = ~pi002 & ~n3778;
  assign n3780 = ~pi002 & pi117;
  assign n3781 = ~pi061 & ~pi105;
  assign n3782 = ~pi064 & n3781;
  assign n3783 = pi067 & n3782;
  assign n3784 = ~pi064 & n3765;
  assign n3785 = pi032 & n3784;
  assign n3786 = pi067 & n3785;
  assign n3787 = pi061 & pi064;
  assign n3788 = pi032 & n3787;
  assign n3789 = ~pi067 & n3788;
  assign n3790 = ~n3786 & ~n3789;
  assign n3791 = ~n3783 & n3790;
  assign n3792 = n3780 & ~n3791;
  assign n3793 = pi061 & ~pi105;
  assign n3794 = pi064 & n3793;
  assign n3795 = ~pi067 & n3794;
  assign n3796 = ~pi032 & n3795;
  assign n3797 = pi032 & n3782;
  assign n3798 = pi067 & n3797;
  assign n3799 = ~n3796 & ~n3798;
  assign n3800 = ~pi117 & ~n3799;
  assign n3801 = ~n3792 & ~n3800;
  assign n3802 = ~n3779 & n3801;
  assign n3803 = ~pi061 & pi064;
  assign n3804 = pi032 & n3803;
  assign n3805 = ~pi064 & n3793;
  assign n3806 = ~pi032 & n3805;
  assign n3807 = ~pi032 & n3766;
  assign n3808 = ~n3806 & ~n3807;
  assign n3809 = ~n3804 & n3808;
  assign n3810 = pi067 & ~n3809;
  assign n3811 = pi064 & n3781;
  assign n3812 = pi067 & n3811;
  assign n3813 = ~n3810 & ~n3812;
  assign n3814 = ~pi117 & ~n3813;
  assign n3815 = pi067 & n3794;
  assign n3816 = ~pi032 & n3784;
  assign n3817 = ~n3815 & ~n3816;
  assign n3818 = ~pi032 & n3765;
  assign n3819 = ~pi032 & n3811;
  assign n3820 = ~n3818 & ~n3819;
  assign n3821 = ~pi061 & pi105;
  assign n3822 = ~pi064 & n3821;
  assign n3823 = pi032 & n3822;
  assign n3824 = n3820 & ~n3823;
  assign n3825 = ~pi067 & ~n3824;
  assign n3826 = n3817 & ~n3825;
  assign n3827 = pi117 & ~n3826;
  assign n3828 = ~n3814 & ~n3827;
  assign n3829 = pi002 & ~n3828;
  assign n3830 = pi032 & n3793;
  assign n3831 = ~pi067 & n3830;
  assign n3832 = ~pi117 & n3831;
  assign n3833 = ~pi061 & ~pi064;
  assign n3834 = pi032 & n3833;
  assign n3835 = ~n3788 & ~n3834;
  assign n3836 = ~n3830 & n3835;
  assign n3837 = ~pi117 & ~n3836;
  assign n3838 = ~pi117 & n3794;
  assign n3839 = ~pi067 & n3771;
  assign n3840 = pi117 & n3839;
  assign n3841 = ~pi067 & n3793;
  assign n3842 = ~pi117 & n3841;
  assign n3843 = ~n3840 & ~n3842;
  assign n3844 = ~n3838 & n3843;
  assign n3845 = ~n3837 & n3844;
  assign n3846 = ~pi032 & n3803;
  assign n3847 = pi067 & n3846;
  assign n3848 = ~n3831 & ~n3847;
  assign n3849 = n3845 & n3848;
  assign n3850 = ~pi002 & ~n3849;
  assign n3851 = ~pi067 & n3818;
  assign n3852 = ~pi067 & n3804;
  assign n3853 = ~n3851 & ~n3852;
  assign n3854 = pi032 & n3794;
  assign n3855 = n3853 & ~n3854;
  assign n3856 = pi117 & ~n3855;
  assign n3857 = pi032 & ~pi067;
  assign n3858 = n3762 & n3857;
  assign n3859 = pi061 & ~pi064;
  assign n3860 = ~pi032 & n3859;
  assign n3861 = pi067 & pi117;
  assign n3862 = n3860 & n3861;
  assign n3863 = ~n3858 & ~n3862;
  assign n3864 = ~n3856 & n3863;
  assign n3865 = pi002 & pi117;
  assign n3866 = ~pi067 & n3781;
  assign n3867 = ~n3834 & ~n3866;
  assign n3868 = pi067 & n3793;
  assign n3869 = ~pi032 & pi061;
  assign n3870 = ~n3868 & ~n3869;
  assign n3871 = n3867 & n3870;
  assign n3872 = n3865 & ~n3871;
  assign n3873 = ~pi067 & ~pi117;
  assign n3874 = n3822 & n3873;
  assign n3875 = ~n3786 & ~n3874;
  assign n3876 = pi002 & ~n3875;
  assign n3877 = ~n3872 & ~n3876;
  assign n3878 = n3864 & n3877;
  assign n3879 = ~n3850 & n3878;
  assign n3880 = ~n3832 & n3879;
  assign n3881 = pi036 & ~n3880;
  assign n3882 = pi032 & n3811;
  assign n3883 = pi032 & n3766;
  assign n3884 = ~n3882 & ~n3883;
  assign n3885 = n3861 & ~n3884;
  assign n3886 = ~pi032 & n3782;
  assign n3887 = n3861 & n3886;
  assign n3888 = ~pi067 & n3785;
  assign n3889 = pi064 & n3821;
  assign n3890 = pi067 & n3889;
  assign n3891 = ~n3888 & ~n3890;
  assign n3892 = ~pi061 & pi067;
  assign n3893 = pi032 & n3892;
  assign n3894 = pi067 & n3805;
  assign n3895 = ~n3893 & ~n3894;
  assign n3896 = ~pi117 & ~n3895;
  assign n3897 = ~pi067 & pi117;
  assign n3898 = pi032 & n3859;
  assign n3899 = n3897 & n3898;
  assign n3900 = ~n3896 & ~n3899;
  assign n3901 = n3891 & n3900;
  assign n3902 = pi002 & ~n3901;
  assign n3903 = pi067 & n3854;
  assign n3904 = ~n3797 & ~n3903;
  assign n3905 = ~pi117 & ~n3904;
  assign n3906 = ~n3769 & ~n3905;
  assign n3907 = ~n3902 & n3906;
  assign n3908 = ~n3887 & n3907;
  assign n3909 = ~n3885 & n3908;
  assign n3910 = ~pi032 & pi105;
  assign n3911 = ~pi117 & n3910;
  assign n3912 = ~pi032 & n3775;
  assign n3913 = pi067 & n3912;
  assign n3914 = ~n3911 & ~n3913;
  assign n3915 = ~pi002 & ~n3914;
  assign n3916 = pi032 & n3770;
  assign n3917 = n3861 & n3916;
  assign n3918 = pi117 & n3782;
  assign n3919 = ~n3917 & ~n3918;
  assign n3920 = ~pi002 & ~n3919;
  assign n3921 = ~n3915 & ~n3920;
  assign n3922 = n3909 & n3921;
  assign n3923 = ~pi036 & ~n3922;
  assign n3924 = ~n3881 & ~n3923;
  assign n3925 = ~n3829 & n3924;
  assign n3926 = n3802 & n3925;
  assign n3927 = ~pi032 & n3833;
  assign n3928 = ~pi067 & n3927;
  assign n3929 = pi032 & n3889;
  assign n3930 = ~pi067 & n3929;
  assign n3931 = pi067 & n3766;
  assign n3932 = ~n3930 & ~n3931;
  assign n3933 = ~n3928 & n3932;
  assign n3934 = ~pi117 & ~n3933;
  assign n3935 = ~pi032 & pi067;
  assign n3936 = ~n3811 & ~n3859;
  assign n3937 = n3935 & ~n3936;
  assign n3938 = pi117 & n3937;
  assign n3939 = ~pi067 & ~n3808;
  assign n3940 = pi032 & n3781;
  assign n3941 = pi067 & n3940;
  assign n3942 = ~pi117 & n3941;
  assign n3943 = ~n3939 & ~n3942;
  assign n3944 = ~pi002 & ~n3943;
  assign n3945 = ~pi067 & n3775;
  assign n3946 = ~n3889 & ~n3945;
  assign n3947 = n3780 & ~n3946;
  assign n3948 = ~n3944 & ~n3947;
  assign n3949 = pi064 & n3861;
  assign n3950 = n3793 & n3949;
  assign n3951 = n3770 & n3873;
  assign n3952 = ~pi032 & n3781;
  assign n3953 = ~n3866 & ~n3952;
  assign n3954 = pi067 & n3765;
  assign n3955 = pi032 & n3954;
  assign n3956 = n3953 & ~n3955;
  assign n3957 = ~n3951 & n3956;
  assign n3958 = ~n3950 & n3957;
  assign n3959 = pi002 & ~n3958;
  assign n3960 = n3948 & ~n3959;
  assign n3961 = ~n3938 & n3960;
  assign n3962 = ~n3934 & n3961;
  assign n3963 = ~pi036 & ~n3962;
  assign n3964 = ~pi032 & n3822;
  assign n3965 = pi067 & n3964;
  assign n3966 = ~n3795 & ~n3965;
  assign n3967 = ~n3858 & ~n3883;
  assign n3968 = ~pi117 & ~n3967;
  assign n3969 = ~pi117 & n3782;
  assign n3970 = pi032 & n3805;
  assign n3971 = ~pi117 & n3787;
  assign n3972 = ~n3970 & ~n3971;
  assign n3973 = ~n3969 & n3972;
  assign n3974 = pi002 & ~n3973;
  assign n3975 = pi032 & pi067;
  assign n3976 = pi064 & n3975;
  assign n3977 = n3781 & n3976;
  assign n3978 = ~n3930 & ~n3977;
  assign n3979 = ~n3913 & n3978;
  assign n3980 = ~n3964 & n3979;
  assign n3981 = pi117 & ~n3980;
  assign n3982 = ~pi032 & n3821;
  assign n3983 = pi067 & n3982;
  assign n3984 = ~pi064 & pi067;
  assign n3985 = ~pi032 & n3984;
  assign n3986 = ~n3764 & ~n3985;
  assign n3987 = ~n3983 & n3986;
  assign n3988 = ~pi067 & n3782;
  assign n3989 = ~n3854 & ~n3988;
  assign n3990 = ~n3785 & n3989;
  assign n3991 = pi117 & ~n3990;
  assign n3992 = n3823 & n3873;
  assign n3993 = ~n3991 & ~n3992;
  assign n3994 = n3987 & n3993;
  assign n3995 = ~pi002 & ~n3994;
  assign n3996 = ~pi032 & ~pi105;
  assign n3997 = pi067 & n3996;
  assign n3998 = pi067 & n3859;
  assign n3999 = ~n3997 & ~n3998;
  assign n4000 = ~pi117 & ~n3999;
  assign n4001 = ~n3995 & ~n4000;
  assign n4002 = ~n3981 & n4001;
  assign n4003 = ~n3974 & n4002;
  assign n4004 = ~n3968 & n4003;
  assign n4005 = n3966 & n4004;
  assign n4006 = pi036 & ~n4005;
  assign n4007 = ~n3963 & ~n4006;
  assign n4008 = pi067 & n3822;
  assign n4009 = pi117 & n4008;
  assign n4010 = pi067 & n3819;
  assign n4011 = n3805 & n3857;
  assign n4012 = pi117 & ~n4011;
  assign n4013 = ~pi117 & ~n3777;
  assign n4014 = ~n4012 & ~n4013;
  assign n4015 = ~n4010 & ~n4014;
  assign n4016 = ~n4009 & n4015;
  assign n4017 = ~pi032 & ~pi067;
  assign n4018 = n3782 & n4017;
  assign n4019 = n4016 & ~n4018;
  assign n4020 = pi002 & ~n4019;
  assign n4021 = ~pi067 & n3805;
  assign n4022 = n3811 & n4017;
  assign n4023 = ~n4021 & ~n4022;
  assign n4024 = ~n3831 & n4023;
  assign n4025 = ~pi117 & ~n4024;
  assign n4026 = ~pi117 & n3935;
  assign n4027 = n3794 & n4026;
  assign n4028 = pi117 & n3977;
  assign n4029 = n3822 & n4017;
  assign n4030 = n3787 & n4017;
  assign n4031 = ~n4029 & ~n4030;
  assign n4032 = pi117 & ~n4031;
  assign n4033 = ~n4028 & ~n4032;
  assign n4034 = ~n4027 & n4033;
  assign n4035 = ~n4025 & n4034;
  assign n4036 = ~pi002 & ~n4035;
  assign n4037 = ~n4020 & ~n4036;
  assign n4038 = n4007 & n4037;
  assign n4039 = pi117 & ~n3796;
  assign n4040 = ~pi117 & ~n3955;
  assign n4041 = ~n4039 & ~n4040;
  assign n4042 = n4038 & ~n4041;
  assign n4043 = ~n3926 & n4042;
  assign n4044 = n3926 & ~n4042;
  assign n4045 = ~n4043 & ~n4044;
  assign n4046 = ~pi008 & n3694;
  assign n4047 = ~n3622 & ~n4046;
  assign n4048 = n3592 & ~n4047;
  assign n4049 = ~pi008 & ~pi115;
  assign n4050 = n3656 & n4049;
  assign n4051 = n3600 & n3639;
  assign n4052 = pi115 & n3684;
  assign n4053 = ~n4051 & ~n4052;
  assign n4054 = ~n4050 & n4053;
  assign n4055 = ~pi008 & n3593;
  assign n4056 = ~n3594 & ~n4055;
  assign n4057 = n4054 & n4056;
  assign n4058 = pi026 & ~n4057;
  assign n4059 = ~n3616 & ~n3654;
  assign n4060 = pi008 & ~pi059;
  assign n4061 = ~n4059 & n4060;
  assign n4062 = pi115 & n4061;
  assign n4063 = ~n4058 & ~n4062;
  assign n4064 = ~n4048 & n4063;
  assign n4065 = ~pi008 & n3691;
  assign n4066 = ~n3704 & ~n4065;
  assign n4067 = pi008 & n3601;
  assign n4068 = n4066 & ~n4067;
  assign n4069 = ~pi115 & ~n4068;
  assign n4070 = ~n3626 & ~n3671;
  assign n4071 = ~pi008 & ~n4070;
  assign n4072 = n3593 & n3639;
  assign n4073 = ~pi115 & n4072;
  assign n4074 = ~n4071 & ~n4073;
  assign n4075 = ~pi026 & ~n4074;
  assign n4076 = ~n4069 & ~n4075;
  assign n4077 = n4064 & n4076;
  assign n4078 = ~pi030 & ~n4077;
  assign n4079 = ~pi059 & n3597;
  assign n4080 = pi008 & n4079;
  assign n4081 = ~n3621 & ~n4080;
  assign n4082 = ~n3740 & ~n3744;
  assign n4083 = ~n3704 & n4082;
  assign n4084 = ~n4079 & n4083;
  assign n4085 = pi115 & ~n4084;
  assign n4086 = ~pi008 & pi059;
  assign n4087 = n3640 & n4086;
  assign n4088 = ~n3602 & ~n4087;
  assign n4089 = ~pi115 & ~n4088;
  assign n4090 = ~n4085 & ~n4089;
  assign n4091 = pi008 & n3654;
  assign n4092 = pi008 & n3709;
  assign n4093 = ~n4091 & ~n4092;
  assign n4094 = ~pi115 & ~n4093;
  assign n4095 = pi008 & ~pi095;
  assign n4096 = ~pi059 & n4095;
  assign n4097 = ~pi059 & n3596;
  assign n4098 = pi008 & n4097;
  assign n4099 = ~n4096 & ~n4098;
  assign n4100 = ~pi059 & n3640;
  assign n4101 = ~pi008 & n4100;
  assign n4102 = n4099 & ~n4101;
  assign n4103 = n3606 & n4049;
  assign n4104 = pi059 & n3620;
  assign n4105 = ~n3711 & ~n4104;
  assign n4106 = ~n3631 & n4105;
  assign n4107 = pi115 & ~n4106;
  assign n4108 = ~n4103 & ~n4107;
  assign n4109 = n4102 & n4108;
  assign n4110 = ~pi026 & ~n4109;
  assign n4111 = ~n4094 & ~n4110;
  assign n4112 = ~pi115 & n3729;
  assign n4113 = ~n3736 & ~n4112;
  assign n4114 = ~n3667 & n4113;
  assign n4115 = pi026 & ~n4114;
  assign n4116 = n4111 & ~n4115;
  assign n4117 = n4090 & n4116;
  assign n4118 = n4081 & n4117;
  assign n4119 = pi030 & ~n4118;
  assign n4120 = ~pi008 & n4079;
  assign n4121 = ~pi008 & ~pi059;
  assign n4122 = n3729 & n4121;
  assign n4123 = ~n4120 & ~n4122;
  assign n4124 = n3592 & ~n4123;
  assign n4125 = pi095 & n4121;
  assign n4126 = n3619 & n4125;
  assign n4127 = pi115 & n4126;
  assign n4128 = ~pi115 & n4051;
  assign n4129 = ~n4127 & ~n4128;
  assign n4130 = ~n4124 & n4129;
  assign n4131 = ~pi008 & n3625;
  assign n4132 = n3616 & n4121;
  assign n4133 = ~n4131 & ~n4132;
  assign n4134 = pi059 & n3619;
  assign n4135 = ~pi008 & n4134;
  assign n4136 = n4133 & ~n4135;
  assign n4137 = ~pi115 & ~n4136;
  assign n4138 = pi008 & n3722;
  assign n4139 = ~pi115 & n4138;
  assign n4140 = ~n4137 & ~n4139;
  assign n4141 = ~n3708 & n4140;
  assign n4142 = ~pi026 & ~n4141;
  assign n4143 = pi115 & n4086;
  assign n4144 = n3625 & n4143;
  assign n4145 = pi008 & n3597;
  assign n4146 = pi115 & n4145;
  assign n4147 = ~pi115 & n3695;
  assign n4148 = ~pi008 & n4147;
  assign n4149 = ~n4146 & ~n4148;
  assign n4150 = ~n4144 & n4149;
  assign n4151 = ~pi059 & n3616;
  assign n4152 = pi008 & n4151;
  assign n4153 = ~pi095 & n4121;
  assign n4154 = n3593 & n4153;
  assign n4155 = ~n4152 & ~n4154;
  assign n4156 = n4150 & n4155;
  assign n4157 = pi026 & ~n4156;
  assign n4158 = ~n4142 & ~n4157;
  assign n4159 = n4130 & n4158;
  assign n4160 = ~n4119 & n4159;
  assign n4161 = ~n4078 & n4160;
  assign n4162 = pi059 & n3718;
  assign n4163 = n4070 & ~n4162;
  assign n4164 = pi008 & ~n4163;
  assign n4165 = pi008 & n3616;
  assign n4166 = ~n4164 & ~n4165;
  assign n4167 = ~pi115 & ~n4166;
  assign n4168 = ~n3651 & ~n3684;
  assign n4169 = ~pi059 & n3600;
  assign n4170 = ~n4151 & ~n4169;
  assign n4171 = ~n3606 & n4170;
  assign n4172 = ~pi008 & ~n4171;
  assign n4173 = n4168 & ~n4172;
  assign n4174 = pi115 & ~n4173;
  assign n4175 = ~n4167 & ~n4174;
  assign n4176 = pi026 & ~n4175;
  assign n4177 = pi008 & n3746;
  assign n4178 = ~n4126 & ~n4177;
  assign n4179 = ~pi115 & ~n4178;
  assign n4180 = pi008 & n3631;
  assign n4181 = ~pi008 & n3730;
  assign n4182 = ~n4180 & ~n4181;
  assign n4183 = ~n3686 & n4182;
  assign n4184 = n3592 & ~n4183;
  assign n4185 = ~n3696 & ~n4101;
  assign n4186 = ~pi115 & ~n4185;
  assign n4187 = pi008 & n3657;
  assign n4188 = ~pi115 & n4187;
  assign n4189 = ~n4186 & ~n4188;
  assign n4190 = ~pi008 & n3695;
  assign n4191 = n4189 & ~n4190;
  assign n4192 = ~pi026 & ~n4191;
  assign n4193 = ~n4184 & ~n4192;
  assign n4194 = ~n4179 & n4193;
  assign n4195 = ~pi115 & n4135;
  assign n4196 = pi059 & n3610;
  assign n4197 = ~n3730 & ~n4196;
  assign n4198 = ~n4134 & n4197;
  assign n4199 = ~pi115 & ~n4198;
  assign n4200 = ~pi115 & n3620;
  assign n4201 = ~pi008 & n3657;
  assign n4202 = pi115 & n4201;
  assign n4203 = ~pi008 & n3619;
  assign n4204 = ~pi115 & n4203;
  assign n4205 = ~n4202 & ~n4204;
  assign n4206 = ~n4200 & n4205;
  assign n4207 = ~n4199 & n4206;
  assign n4208 = pi008 & n3719;
  assign n4209 = ~n4135 & ~n4208;
  assign n4210 = n4207 & n4209;
  assign n4211 = ~pi026 & ~n4210;
  assign n4212 = ~pi059 & n3654;
  assign n4213 = n3609 & n4212;
  assign n4214 = ~pi008 & n4169;
  assign n4215 = ~pi008 & n4162;
  assign n4216 = ~n4214 & ~n4215;
  assign n4217 = ~n4104 & n4216;
  assign n4218 = pi115 & ~n4217;
  assign n4219 = ~n4213 & ~n4218;
  assign n4220 = ~n4087 & n4219;
  assign n4221 = ~n4055 & ~n4196;
  assign n4222 = pi008 & n3619;
  assign n4223 = pi056 & ~pi059;
  assign n4224 = ~n4222 & ~n4223;
  assign n4225 = n4221 & n4224;
  assign n4226 = n3728 & ~n4225;
  assign n4227 = n3597 & n4049;
  assign n4228 = ~n4180 & ~n4227;
  assign n4229 = pi026 & ~n4228;
  assign n4230 = ~n4226 & ~n4229;
  assign n4231 = n4220 & n4230;
  assign n4232 = ~n4211 & n4231;
  assign n4233 = ~n4195 & n4232;
  assign n4234 = pi030 & ~n4233;
  assign n4235 = pi059 & n3656;
  assign n4236 = n3609 & n4235;
  assign n4237 = pi115 & n3611;
  assign n4238 = ~n4236 & ~n4237;
  assign n4239 = ~pi026 & ~n4238;
  assign n4240 = ~n3602 & ~n3617;
  assign n4241 = n3609 & ~n4240;
  assign n4242 = ~n3613 & ~n4241;
  assign n4243 = ~n4239 & n4242;
  assign n4244 = ~pi059 & pi099;
  assign n4245 = ~pi115 & n4244;
  assign n4246 = ~n3744 & ~n4245;
  assign n4247 = ~pi026 & ~n4246;
  assign n4248 = n4243 & ~n4247;
  assign n4249 = pi008 & n4104;
  assign n4250 = ~n3746 & ~n4249;
  assign n4251 = ~pi115 & ~n4250;
  assign n4252 = ~n4186 & ~n4251;
  assign n4253 = n4248 & n4252;
  assign n4254 = ~n3623 & ~n3632;
  assign n4255 = ~pi056 & n3639;
  assign n4256 = ~n3742 & ~n4255;
  assign n4257 = ~pi115 & ~n4256;
  assign n4258 = ~pi008 & pi115;
  assign n4259 = n3655 & n4258;
  assign n4260 = ~n4257 & ~n4259;
  assign n4261 = n4254 & n4260;
  assign n4262 = pi026 & ~n4261;
  assign n4263 = n4253 & ~n4262;
  assign n4264 = ~pi030 & ~n4263;
  assign n4265 = ~n4234 & ~n4264;
  assign n4266 = n4194 & n4265;
  assign n4267 = ~n4176 & n4266;
  assign n4268 = ~n4161 & n4267;
  assign n4269 = n4161 & ~n4267;
  assign n4270 = ~n4268 & ~n4269;
  assign n4271 = ~n4045 & n4270;
  assign n4272 = n3926 & n4042;
  assign n4273 = ~n3926 & ~n4042;
  assign n4274 = ~n4272 & ~n4273;
  assign n4275 = ~n4270 & ~n4274;
  assign n4276 = ~n4271 & ~n4275;
  assign n4277 = n3761 & n4276;
  assign n4278 = ~n3761 & ~n4276;
  assign n4279 = ~n4277 & ~n4278;
  assign n4280 = ~pi529 & n4279;
  assign po132 = n3256 | n4280;
  assign n4282 = pi303 & pi478;
  assign n4283 = ~pi303 & ~pi478;
  assign n4284 = ~n4282 & ~n4283;
  assign n4285 = pi529 & n4284;
  assign n4286 = ~pi051 & ~pi112;
  assign n4287 = pi086 & n4286;
  assign n4288 = pi049 & n4287;
  assign n4289 = pi019 & n4288;
  assign n4290 = pi019 & pi049;
  assign n4291 = pi051 & ~pi112;
  assign n4292 = ~pi086 & n4291;
  assign n4293 = n4290 & n4292;
  assign n4294 = ~pi051 & pi112;
  assign n4295 = ~pi086 & n4294;
  assign n4296 = pi019 & n4295;
  assign n4297 = ~pi086 & n4286;
  assign n4298 = pi049 & n4297;
  assign n4299 = ~pi019 & n4298;
  assign n4300 = ~n4296 & ~n4299;
  assign n4301 = pi051 & pi086;
  assign n4302 = ~pi049 & n4301;
  assign n4303 = pi019 & n4302;
  assign n4304 = n4300 & ~n4303;
  assign n4305 = ~pi090 & ~n4304;
  assign n4306 = ~n4293 & ~n4305;
  assign n4307 = ~n4289 & n4306;
  assign n4308 = ~pi088 & ~n4307;
  assign n4309 = pi051 & pi112;
  assign n4310 = ~pi086 & n4309;
  assign n4311 = pi049 & n4310;
  assign n4312 = ~pi019 & n4311;
  assign n4313 = ~pi049 & n4310;
  assign n4314 = pi086 & pi112;
  assign n4315 = pi049 & n4314;
  assign n4316 = ~n4313 & ~n4315;
  assign n4317 = pi019 & ~n4316;
  assign n4318 = ~n4312 & ~n4317;
  assign n4319 = pi088 & pi090;
  assign n4320 = ~n4318 & n4319;
  assign n4321 = ~n4308 & ~n4320;
  assign n4322 = pi019 & pi090;
  assign n4323 = ~pi049 & n4322;
  assign n4324 = ~pi086 & n4323;
  assign n4325 = n4286 & n4324;
  assign n4326 = pi090 & n4293;
  assign n4327 = ~n4325 & ~n4326;
  assign n4328 = pi019 & ~pi090;
  assign n4329 = n4297 & n4328;
  assign n4330 = ~pi019 & n4287;
  assign n4331 = pi086 & n4294;
  assign n4332 = ~pi049 & n4331;
  assign n4333 = ~n4330 & ~n4332;
  assign n4334 = pi086 & ~pi112;
  assign n4335 = ~pi049 & n4334;
  assign n4336 = ~pi019 & n4335;
  assign n4337 = ~pi049 & n4297;
  assign n4338 = ~n4336 & ~n4337;
  assign n4339 = n4333 & n4338;
  assign n4340 = ~pi090 & ~n4339;
  assign n4341 = ~n4329 & ~n4340;
  assign n4342 = pi088 & ~n4341;
  assign n4343 = ~pi088 & pi090;
  assign n4344 = ~pi049 & n4286;
  assign n4345 = ~pi019 & n4344;
  assign n4346 = ~pi019 & n4292;
  assign n4347 = pi086 & n4309;
  assign n4348 = pi049 & n4347;
  assign n4349 = ~pi019 & n4348;
  assign n4350 = ~n4346 & ~n4349;
  assign n4351 = ~n4345 & n4350;
  assign n4352 = n4343 & ~n4351;
  assign n4353 = ~n4342 & ~n4352;
  assign n4354 = n4327 & n4353;
  assign n4355 = n4321 & n4354;
  assign n4356 = ~pi049 & n4347;
  assign n4357 = pi019 & n4356;
  assign n4358 = ~pi090 & n4357;
  assign n4359 = pi086 & n4291;
  assign n4360 = pi049 & n4359;
  assign n4361 = ~pi090 & n4360;
  assign n4362 = ~pi019 & n4361;
  assign n4363 = ~n4358 & ~n4362;
  assign n4364 = ~n4345 & n4363;
  assign n4365 = ~pi019 & n4310;
  assign n4366 = ~pi049 & n4365;
  assign n4367 = pi049 & n4295;
  assign n4368 = ~n4366 & ~n4367;
  assign n4369 = ~pi090 & ~n4368;
  assign n4370 = n4290 & n4295;
  assign n4371 = pi019 & n4310;
  assign n4372 = pi090 & n4371;
  assign n4373 = ~n4370 & ~n4372;
  assign n4374 = ~n4357 & n4373;
  assign n4375 = ~n4369 & n4374;
  assign n4376 = ~pi019 & n4331;
  assign n4377 = pi090 & n4376;
  assign n4378 = n4375 & ~n4377;
  assign n4379 = ~pi088 & ~n4378;
  assign n4380 = n4364 & ~n4379;
  assign n4381 = pi090 & n4289;
  assign n4382 = ~pi019 & ~n4291;
  assign n4383 = ~pi086 & pi112;
  assign n4384 = pi049 & n4383;
  assign n4385 = pi019 & ~n4384;
  assign n4386 = ~n4382 & ~n4385;
  assign n4387 = ~pi086 & ~pi112;
  assign n4388 = ~pi049 & n4387;
  assign n4389 = ~n4386 & ~n4388;
  assign n4390 = ~pi090 & ~n4389;
  assign n4391 = pi019 & n4297;
  assign n4392 = pi019 & n4331;
  assign n4393 = ~pi049 & n4294;
  assign n4394 = pi019 & n4393;
  assign n4395 = ~n4392 & ~n4394;
  assign n4396 = ~n4391 & n4395;
  assign n4397 = ~pi019 & n4347;
  assign n4398 = pi049 & n4301;
  assign n4399 = ~n4397 & ~n4398;
  assign n4400 = pi090 & ~n4399;
  assign n4401 = n4396 & ~n4400;
  assign n4402 = ~n4390 & n4401;
  assign n4403 = pi088 & ~n4402;
  assign n4404 = ~pi019 & n4297;
  assign n4405 = ~pi049 & ~pi051;
  assign n4406 = ~pi019 & n4405;
  assign n4407 = ~n4404 & ~n4406;
  assign n4408 = pi090 & ~n4407;
  assign n4409 = ~n4403 & ~n4408;
  assign n4410 = ~n4381 & n4409;
  assign n4411 = n4380 & n4410;
  assign n4412 = ~pi006 & ~n4411;
  assign n4413 = ~pi019 & n4288;
  assign n4414 = pi019 & n4359;
  assign n4415 = ~pi049 & ~pi086;
  assign n4416 = n4294 & n4415;
  assign n4417 = ~n4288 & ~n4376;
  assign n4418 = ~n4416 & n4417;
  assign n4419 = ~n4414 & n4418;
  assign n4420 = ~pi090 & ~n4419;
  assign n4421 = ~n4413 & ~n4420;
  assign n4422 = pi090 & n4365;
  assign n4423 = pi019 & n4348;
  assign n4424 = pi019 & n4309;
  assign n4425 = pi051 & ~pi086;
  assign n4426 = ~pi049 & n4425;
  assign n4427 = ~n4424 & ~n4426;
  assign n4428 = ~n4384 & n4427;
  assign n4429 = pi090 & ~n4428;
  assign n4430 = ~n4313 & ~n4429;
  assign n4431 = ~n4423 & n4430;
  assign n4432 = pi088 & ~n4431;
  assign n4433 = ~n4422 & ~n4432;
  assign n4434 = pi019 & n4291;
  assign n4435 = ~pi090 & n4434;
  assign n4436 = ~pi049 & n4359;
  assign n4437 = ~pi019 & n4436;
  assign n4438 = ~n4435 & ~n4437;
  assign n4439 = ~pi051 & pi086;
  assign n4440 = n4290 & n4439;
  assign n4441 = ~n4416 & ~n4440;
  assign n4442 = pi049 & n4434;
  assign n4443 = n4441 & ~n4442;
  assign n4444 = n4438 & n4443;
  assign n4445 = ~pi088 & ~n4444;
  assign n4446 = n4433 & ~n4445;
  assign n4447 = ~n4312 & n4446;
  assign n4448 = n4421 & n4447;
  assign n4449 = pi006 & ~n4448;
  assign n4450 = ~n4412 & ~n4449;
  assign n4451 = n4355 & n4450;
  assign n4452 = ~pi303 & ~n4451;
  assign n4453 = pi303 & n4451;
  assign n4454 = ~n4452 & ~n4453;
  assign n4455 = ~pi057 & ~pi097;
  assign n4456 = pi022 & n4455;
  assign n4457 = pi000 & n4456;
  assign n4458 = pi011 & n4457;
  assign n4459 = ~pi057 & pi097;
  assign n4460 = ~pi022 & n4459;
  assign n4461 = pi000 & n4460;
  assign n4462 = pi011 & n4461;
  assign n4463 = ~n4458 & ~n4462;
  assign n4464 = pi057 & ~pi097;
  assign n4465 = ~pi022 & n4464;
  assign n4466 = pi011 & n4465;
  assign n4467 = pi022 & pi097;
  assign n4468 = ~pi000 & n4467;
  assign n4469 = pi011 & n4468;
  assign n4470 = ~n4466 & ~n4469;
  assign n4471 = ~pi022 & n4455;
  assign n4472 = pi000 & n4471;
  assign n4473 = ~pi011 & n4472;
  assign n4474 = n4470 & ~n4473;
  assign n4475 = ~pi116 & ~n4474;
  assign n4476 = n4463 & ~n4475;
  assign n4477 = ~pi058 & ~n4476;
  assign n4478 = ~pi022 & ~pi057;
  assign n4479 = ~pi097 & n4478;
  assign n4480 = ~pi000 & n4479;
  assign n4481 = pi011 & pi116;
  assign n4482 = n4480 & n4481;
  assign n4483 = pi116 & n4462;
  assign n4484 = pi011 & ~pi116;
  assign n4485 = n4471 & n4484;
  assign n4486 = pi022 & ~pi057;
  assign n4487 = ~pi000 & n4486;
  assign n4488 = ~pi011 & n4487;
  assign n4489 = ~pi011 & n4456;
  assign n4490 = pi022 & n4464;
  assign n4491 = ~pi000 & n4490;
  assign n4492 = ~n4480 & ~n4491;
  assign n4493 = ~n4489 & n4492;
  assign n4494 = ~n4488 & n4493;
  assign n4495 = ~pi116 & ~n4494;
  assign n4496 = ~n4485 & ~n4495;
  assign n4497 = pi058 & ~n4496;
  assign n4498 = pi057 & pi097;
  assign n4499 = ~pi022 & n4498;
  assign n4500 = pi000 & ~pi011;
  assign n4501 = n4499 & n4500;
  assign n4502 = ~pi000 & n4499;
  assign n4503 = pi022 & pi057;
  assign n4504 = pi000 & n4503;
  assign n4505 = ~n4502 & ~n4504;
  assign n4506 = pi011 & ~n4505;
  assign n4507 = ~n4501 & ~n4506;
  assign n4508 = pi058 & pi116;
  assign n4509 = ~n4507 & n4508;
  assign n4510 = ~n4497 & ~n4509;
  assign n4511 = ~pi058 & pi116;
  assign n4512 = ~pi000 & ~pi011;
  assign n4513 = ~pi097 & n4512;
  assign n4514 = ~pi057 & n4513;
  assign n4515 = ~pi011 & n4460;
  assign n4516 = ~n4514 & ~n4515;
  assign n4517 = pi022 & n4498;
  assign n4518 = pi000 & n4517;
  assign n4519 = ~pi011 & n4518;
  assign n4520 = n4516 & ~n4519;
  assign n4521 = n4511 & ~n4520;
  assign n4522 = n4510 & ~n4521;
  assign n4523 = ~n4483 & n4522;
  assign n4524 = ~n4482 & n4523;
  assign n4525 = ~pi000 & n4517;
  assign n4526 = pi011 & n4525;
  assign n4527 = pi022 & n4459;
  assign n4528 = pi000 & n4527;
  assign n4529 = ~pi011 & n4528;
  assign n4530 = ~n4526 & ~n4529;
  assign n4531 = ~pi116 & ~n4530;
  assign n4532 = pi011 & n4499;
  assign n4533 = pi116 & n4532;
  assign n4534 = pi000 & n4465;
  assign n4535 = ~pi011 & n4499;
  assign n4536 = ~pi000 & n4535;
  assign n4537 = ~n4534 & ~n4536;
  assign n4538 = ~pi116 & ~n4537;
  assign n4539 = ~n4526 & ~n4538;
  assign n4540 = ~pi011 & pi116;
  assign n4541 = n4490 & n4540;
  assign n4542 = pi011 & n4534;
  assign n4543 = ~n4541 & ~n4542;
  assign n4544 = n4539 & n4543;
  assign n4545 = ~n4533 & n4544;
  assign n4546 = ~pi058 & ~n4545;
  assign n4547 = ~pi000 & n4464;
  assign n4548 = pi011 & n4547;
  assign n4549 = pi011 & n4490;
  assign n4550 = ~n4548 & ~n4549;
  assign n4551 = pi011 & n4471;
  assign n4552 = n4550 & ~n4551;
  assign n4553 = pi000 & n4467;
  assign n4554 = ~pi011 & n4517;
  assign n4555 = ~n4553 & ~n4554;
  assign n4556 = pi116 & ~n4555;
  assign n4557 = ~pi011 & ~n4459;
  assign n4558 = ~pi022 & pi057;
  assign n4559 = pi000 & n4558;
  assign n4560 = pi011 & ~n4559;
  assign n4561 = ~n4557 & ~n4560;
  assign n4562 = ~pi000 & n4478;
  assign n4563 = ~n4561 & ~n4562;
  assign n4564 = ~pi116 & ~n4563;
  assign n4565 = ~n4556 & ~n4564;
  assign n4566 = n4552 & n4565;
  assign n4567 = pi058 & ~n4566;
  assign n4568 = ~n4546 & ~n4567;
  assign n4569 = ~n4514 & n4568;
  assign n4570 = ~n4531 & n4569;
  assign n4571 = ~pi000 & ~pi097;
  assign n4572 = ~pi011 & n4571;
  assign n4573 = ~pi011 & n4471;
  assign n4574 = ~n4572 & ~n4573;
  assign n4575 = pi116 & ~n4574;
  assign n4576 = pi116 & n4458;
  assign n4577 = ~n4575 & ~n4576;
  assign n4578 = n4570 & n4577;
  assign n4579 = ~pi060 & ~n4578;
  assign n4580 = pi011 & n4459;
  assign n4581 = pi000 & n4580;
  assign n4582 = ~pi000 & n4465;
  assign n4583 = pi000 & pi011;
  assign n4584 = pi022 & ~pi097;
  assign n4585 = n4583 & n4584;
  assign n4586 = ~n4582 & ~n4585;
  assign n4587 = ~n4581 & n4586;
  assign n4588 = ~pi000 & n4527;
  assign n4589 = ~pi011 & n4588;
  assign n4590 = ~pi116 & n4580;
  assign n4591 = ~n4589 & ~n4590;
  assign n4592 = n4587 & n4591;
  assign n4593 = ~pi058 & ~n4592;
  assign n4594 = ~pi011 & n4490;
  assign n4595 = pi011 & n4527;
  assign n4596 = ~n4594 & ~n4595;
  assign n4597 = ~n4582 & n4596;
  assign n4598 = ~n4457 & n4597;
  assign n4599 = ~pi116 & ~n4598;
  assign n4600 = ~pi011 & n4457;
  assign n4601 = ~n4599 & ~n4600;
  assign n4602 = ~pi022 & pi097;
  assign n4603 = ~pi000 & n4602;
  assign n4604 = ~n4559 & ~n4603;
  assign n4605 = pi011 & n4498;
  assign n4606 = n4604 & ~n4605;
  assign n4607 = pi116 & ~n4606;
  assign n4608 = pi011 & n4518;
  assign n4609 = ~n4502 & ~n4608;
  assign n4610 = ~n4607 & n4609;
  assign n4611 = pi058 & ~n4610;
  assign n4612 = pi116 & n4535;
  assign n4613 = ~n4501 & ~n4612;
  assign n4614 = ~n4611 & n4613;
  assign n4615 = n4601 & n4614;
  assign n4616 = ~n4593 & n4615;
  assign n4617 = pi060 & ~n4616;
  assign n4618 = ~n4579 & ~n4617;
  assign n4619 = n4524 & n4618;
  assign n4620 = ~n4477 & n4619;
  assign n4621 = ~pi034 & pi118;
  assign n4622 = ~pi062 & ~pi119;
  assign n4623 = ~pi103 & n4622;
  assign n4624 = ~pi066 & n4623;
  assign n4625 = pi062 & pi119;
  assign n4626 = pi101 & n4625;
  assign n4627 = pi103 & n4626;
  assign n4628 = ~pi066 & n4627;
  assign n4629 = ~pi062 & pi119;
  assign n4630 = ~pi101 & n4629;
  assign n4631 = ~pi066 & n4630;
  assign n4632 = ~n4628 & ~n4631;
  assign n4633 = ~n4624 & n4632;
  assign n4634 = n4621 & ~n4633;
  assign n4635 = pi062 & ~pi119;
  assign n4636 = ~pi101 & n4635;
  assign n4637 = pi066 & n4636;
  assign n4638 = pi101 & pi119;
  assign n4639 = ~pi103 & n4638;
  assign n4640 = pi066 & n4639;
  assign n4641 = ~n4637 & ~n4640;
  assign n4642 = ~pi101 & n4622;
  assign n4643 = pi103 & n4642;
  assign n4644 = ~pi066 & n4643;
  assign n4645 = n4641 & ~n4644;
  assign n4646 = ~pi118 & ~n4645;
  assign n4647 = pi103 & n4630;
  assign n4648 = pi066 & n4647;
  assign n4649 = pi101 & n4622;
  assign n4650 = pi103 & n4649;
  assign n4651 = pi066 & n4650;
  assign n4652 = ~n4648 & ~n4651;
  assign n4653 = ~n4646 & n4652;
  assign n4654 = ~pi034 & ~n4653;
  assign n4655 = ~n4634 & ~n4654;
  assign n4656 = ~pi101 & n4625;
  assign n4657 = ~pi066 & n4656;
  assign n4658 = pi118 & n4657;
  assign n4659 = ~pi062 & pi101;
  assign n4660 = pi119 & n4659;
  assign n4661 = ~pi103 & n4660;
  assign n4662 = ~pi066 & n4661;
  assign n4663 = pi066 & n4629;
  assign n4664 = ~pi118 & n4663;
  assign n4665 = ~n4662 & ~n4664;
  assign n4666 = pi103 & n4663;
  assign n4667 = ~pi103 & n4636;
  assign n4668 = pi066 & pi103;
  assign n4669 = pi101 & ~pi119;
  assign n4670 = n4668 & n4669;
  assign n4671 = ~n4667 & ~n4670;
  assign n4672 = ~n4666 & n4671;
  assign n4673 = n4665 & n4672;
  assign n4674 = ~pi034 & ~n4673;
  assign n4675 = pi101 & n4635;
  assign n4676 = ~pi066 & n4675;
  assign n4677 = pi066 & n4660;
  assign n4678 = ~n4676 & ~n4677;
  assign n4679 = ~n4650 & ~n4667;
  assign n4680 = n4678 & n4679;
  assign n4681 = ~pi118 & ~n4680;
  assign n4682 = ~n4674 & ~n4681;
  assign n4683 = ~n4658 & n4682;
  assign n4684 = pi103 & n4656;
  assign n4685 = ~pi066 & n4684;
  assign n4686 = ~pi103 & n4656;
  assign n4687 = pi062 & ~pi101;
  assign n4688 = pi103 & n4687;
  assign n4689 = ~pi101 & pi119;
  assign n4690 = ~pi103 & n4689;
  assign n4691 = ~n4688 & ~n4690;
  assign n4692 = pi066 & n4625;
  assign n4693 = n4691 & ~n4692;
  assign n4694 = pi118 & ~n4693;
  assign n4695 = pi066 & n4627;
  assign n4696 = ~n4694 & ~n4695;
  assign n4697 = ~n4686 & n4696;
  assign n4698 = pi034 & ~n4697;
  assign n4699 = ~pi066 & n4650;
  assign n4700 = ~n4698 & ~n4699;
  assign n4701 = ~n4685 & n4700;
  assign n4702 = n4683 & n4701;
  assign n4703 = pi038 & ~n4702;
  assign n4704 = ~pi103 & n4626;
  assign n4705 = pi066 & n4704;
  assign n4706 = pi103 & n4660;
  assign n4707 = ~pi066 & n4706;
  assign n4708 = ~n4705 & ~n4707;
  assign n4709 = ~pi118 & ~n4708;
  assign n4710 = pi103 & n4636;
  assign n4711 = ~pi066 & n4686;
  assign n4712 = ~n4710 & ~n4711;
  assign n4713 = ~pi118 & ~n4712;
  assign n4714 = n4636 & n4668;
  assign n4715 = pi066 & n4656;
  assign n4716 = pi118 & n4715;
  assign n4717 = ~n4705 & ~n4716;
  assign n4718 = ~n4714 & n4717;
  assign n4719 = ~n4713 & n4718;
  assign n4720 = pi118 & n4676;
  assign n4721 = n4719 & ~n4720;
  assign n4722 = ~pi034 & ~n4721;
  assign n4723 = ~pi103 & n4635;
  assign n4724 = pi066 & n4723;
  assign n4725 = pi066 & n4675;
  assign n4726 = ~n4724 & ~n4725;
  assign n4727 = pi066 & n4642;
  assign n4728 = n4726 & ~n4727;
  assign n4729 = ~pi066 & ~n4629;
  assign n4730 = pi066 & ~n4688;
  assign n4731 = ~n4729 & ~n4730;
  assign n4732 = ~pi062 & ~pi101;
  assign n4733 = ~pi103 & n4732;
  assign n4734 = ~n4731 & ~n4733;
  assign n4735 = ~pi118 & ~n4734;
  assign n4736 = pi103 & n4638;
  assign n4737 = ~pi066 & n4626;
  assign n4738 = ~n4736 & ~n4737;
  assign n4739 = pi118 & ~n4738;
  assign n4740 = ~n4735 & ~n4739;
  assign n4741 = n4728 & n4740;
  assign n4742 = pi034 & ~n4741;
  assign n4743 = ~n4722 & ~n4742;
  assign n4744 = ~n4624 & n4743;
  assign n4745 = ~n4709 & n4744;
  assign n4746 = ~pi103 & ~pi119;
  assign n4747 = ~pi066 & n4746;
  assign n4748 = ~pi101 & ~pi119;
  assign n4749 = ~pi066 & n4748;
  assign n4750 = ~pi062 & n4749;
  assign n4751 = ~n4747 & ~n4750;
  assign n4752 = pi118 & ~n4751;
  assign n4753 = pi066 & pi118;
  assign n4754 = n4650 & n4753;
  assign n4755 = ~n4752 & ~n4754;
  assign n4756 = n4745 & n4755;
  assign n4757 = ~pi038 & ~n4756;
  assign n4758 = pi118 & n4648;
  assign n4759 = ~pi103 & n4642;
  assign n4760 = n4753 & n4759;
  assign n4761 = ~n4758 & ~n4760;
  assign n4762 = pi034 & pi118;
  assign n4763 = pi062 & pi101;
  assign n4764 = pi103 & n4763;
  assign n4765 = ~n4686 & ~n4764;
  assign n4766 = pi066 & ~n4765;
  assign n4767 = ~n4685 & ~n4766;
  assign n4768 = n4762 & ~n4767;
  assign n4769 = n4761 & ~n4768;
  assign n4770 = pi034 & pi066;
  assign n4771 = ~pi118 & n4642;
  assign n4772 = n4770 & n4771;
  assign n4773 = ~pi066 & n4649;
  assign n4774 = ~pi103 & n4675;
  assign n4775 = ~pi103 & n4659;
  assign n4776 = ~pi066 & n4775;
  assign n4777 = ~n4774 & ~n4776;
  assign n4778 = ~n4759 & n4777;
  assign n4779 = ~n4773 & n4778;
  assign n4780 = ~pi118 & ~n4779;
  assign n4781 = pi034 & n4780;
  assign n4782 = ~n4772 & ~n4781;
  assign n4783 = n4769 & n4782;
  assign n4784 = ~n4757 & n4783;
  assign n4785 = ~n4703 & n4784;
  assign n4786 = n4655 & n4785;
  assign n4787 = ~n4620 & n4786;
  assign n4788 = n4620 & ~n4786;
  assign n4789 = ~n4787 & ~n4788;
  assign n4790 = ~n4454 & n4789;
  assign n4791 = n4454 & ~n4789;
  assign n4792 = ~n4790 & ~n4791;
  assign n4793 = ~pi045 & pi081;
  assign n4794 = pi041 & n4793;
  assign n4795 = pi074 & n4794;
  assign n4796 = pi045 & pi081;
  assign n4797 = ~pi041 & n4796;
  assign n4798 = ~pi016 & n4797;
  assign n4799 = ~n4795 & ~n4798;
  assign n4800 = ~pi016 & n4796;
  assign n4801 = ~pi045 & ~pi081;
  assign n4802 = pi041 & n4801;
  assign n4803 = ~pi016 & n4802;
  assign n4804 = ~n4800 & ~n4803;
  assign n4805 = pi045 & ~pi081;
  assign n4806 = ~pi041 & n4805;
  assign n4807 = pi016 & n4806;
  assign n4808 = n4804 & ~n4807;
  assign n4809 = ~pi074 & ~n4808;
  assign n4810 = n4799 & ~n4809;
  assign n4811 = pi120 & ~n4810;
  assign n4812 = pi041 & ~pi081;
  assign n4813 = pi016 & n4812;
  assign n4814 = ~pi041 & n4793;
  assign n4815 = ~pi016 & n4814;
  assign n4816 = pi041 & n4796;
  assign n4817 = ~pi016 & n4816;
  assign n4818 = ~n4815 & ~n4817;
  assign n4819 = ~n4813 & n4818;
  assign n4820 = pi074 & ~n4819;
  assign n4821 = pi074 & n4802;
  assign n4822 = ~n4820 & ~n4821;
  assign n4823 = ~pi120 & ~n4822;
  assign n4824 = ~n4811 & ~n4823;
  assign n4825 = pi003 & ~n4824;
  assign n4826 = pi016 & n4797;
  assign n4827 = pi074 & n4826;
  assign n4828 = ~pi041 & n4801;
  assign n4829 = pi074 & n4828;
  assign n4830 = pi041 & pi081;
  assign n4831 = pi016 & n4830;
  assign n4832 = ~pi074 & n4831;
  assign n4833 = ~n4829 & ~n4832;
  assign n4834 = ~n4827 & n4833;
  assign n4835 = ~pi003 & pi120;
  assign n4836 = ~n4834 & n4835;
  assign n4837 = pi041 & ~pi045;
  assign n4838 = ~pi016 & n4837;
  assign n4839 = ~pi074 & n4838;
  assign n4840 = ~pi074 & n4816;
  assign n4841 = ~n4839 & ~n4840;
  assign n4842 = ~pi120 & ~n4841;
  assign n4843 = pi041 & pi045;
  assign n4844 = pi016 & n4843;
  assign n4845 = ~pi074 & n4844;
  assign n4846 = ~pi041 & pi045;
  assign n4847 = ~pi016 & n4846;
  assign n4848 = pi074 & n4847;
  assign n4849 = ~pi120 & n4848;
  assign n4850 = ~n4845 & ~n4849;
  assign n4851 = ~n4842 & n4850;
  assign n4852 = ~pi003 & ~n4851;
  assign n4853 = ~n4836 & ~n4852;
  assign n4854 = ~pi016 & n4794;
  assign n4855 = ~pi074 & n4854;
  assign n4856 = pi016 & n4828;
  assign n4857 = pi074 & n4856;
  assign n4858 = ~n4855 & ~n4857;
  assign n4859 = ~pi120 & ~n4858;
  assign n4860 = n4853 & ~n4859;
  assign n4861 = pi016 & n4793;
  assign n4862 = ~pi074 & n4861;
  assign n4863 = ~pi120 & n4862;
  assign n4864 = ~pi041 & ~pi081;
  assign n4865 = pi016 & n4864;
  assign n4866 = ~n4831 & ~n4865;
  assign n4867 = ~n4861 & n4866;
  assign n4868 = ~pi120 & ~n4867;
  assign n4869 = ~pi120 & n4794;
  assign n4870 = ~pi074 & n4847;
  assign n4871 = pi120 & n4870;
  assign n4872 = ~pi074 & n4793;
  assign n4873 = ~pi120 & n4872;
  assign n4874 = ~n4871 & ~n4873;
  assign n4875 = ~n4869 & n4874;
  assign n4876 = ~n4868 & n4875;
  assign n4877 = ~pi016 & n4812;
  assign n4878 = pi074 & n4877;
  assign n4879 = ~n4862 & ~n4878;
  assign n4880 = n4876 & n4879;
  assign n4881 = ~pi003 & ~n4880;
  assign n4882 = pi003 & pi120;
  assign n4883 = ~pi074 & n4801;
  assign n4884 = ~n4865 & ~n4883;
  assign n4885 = pi074 & n4793;
  assign n4886 = ~pi016 & pi081;
  assign n4887 = ~n4885 & ~n4886;
  assign n4888 = n4884 & n4887;
  assign n4889 = n4882 & ~n4888;
  assign n4890 = ~pi074 & ~pi120;
  assign n4891 = n4806 & n4890;
  assign n4892 = ~n4827 & ~n4891;
  assign n4893 = pi003 & ~n4892;
  assign n4894 = ~n4889 & ~n4893;
  assign n4895 = ~pi074 & n4800;
  assign n4896 = ~pi074 & n4813;
  assign n4897 = ~n4895 & ~n4896;
  assign n4898 = pi016 & n4794;
  assign n4899 = n4897 & ~n4898;
  assign n4900 = pi120 & ~n4899;
  assign n4901 = pi016 & ~pi074;
  assign n4902 = n4837 & n4901;
  assign n4903 = ~pi041 & pi081;
  assign n4904 = ~pi016 & n4903;
  assign n4905 = pi074 & pi120;
  assign n4906 = n4904 & n4905;
  assign n4907 = ~n4902 & ~n4906;
  assign n4908 = ~n4900 & n4907;
  assign n4909 = n4894 & n4908;
  assign n4910 = ~n4881 & n4909;
  assign n4911 = ~n4863 & n4910;
  assign n4912 = pi044 & ~n4911;
  assign n4913 = pi016 & n4802;
  assign n4914 = pi016 & n4816;
  assign n4915 = ~n4913 & ~n4914;
  assign n4916 = n4905 & ~n4915;
  assign n4917 = ~pi016 & n4828;
  assign n4918 = n4905 & n4917;
  assign n4919 = ~pi074 & n4826;
  assign n4920 = pi041 & n4805;
  assign n4921 = pi074 & n4920;
  assign n4922 = ~n4919 & ~n4921;
  assign n4923 = pi074 & ~pi081;
  assign n4924 = pi016 & n4923;
  assign n4925 = pi074 & n4814;
  assign n4926 = ~n4924 & ~n4925;
  assign n4927 = ~pi120 & ~n4926;
  assign n4928 = ~pi074 & pi120;
  assign n4929 = pi016 & n4903;
  assign n4930 = n4928 & n4929;
  assign n4931 = ~n4927 & ~n4930;
  assign n4932 = n4922 & n4931;
  assign n4933 = pi003 & ~n4932;
  assign n4934 = pi074 & n4898;
  assign n4935 = ~n4856 & ~n4934;
  assign n4936 = ~pi120 & ~n4935;
  assign n4937 = ~n4842 & ~n4936;
  assign n4938 = ~n4933 & n4937;
  assign n4939 = ~n4918 & n4938;
  assign n4940 = ~n4916 & n4939;
  assign n4941 = ~pi016 & pi045;
  assign n4942 = ~pi120 & n4941;
  assign n4943 = ~pi016 & n4843;
  assign n4944 = pi074 & n4943;
  assign n4945 = ~n4942 & ~n4944;
  assign n4946 = ~pi003 & ~n4945;
  assign n4947 = pi016 & n4846;
  assign n4948 = n4905 & n4947;
  assign n4949 = pi120 & n4828;
  assign n4950 = ~n4948 & ~n4949;
  assign n4951 = ~pi003 & ~n4950;
  assign n4952 = ~n4946 & ~n4951;
  assign n4953 = n4940 & n4952;
  assign n4954 = ~pi044 & ~n4953;
  assign n4955 = ~n4912 & ~n4954;
  assign n4956 = n4860 & n4955;
  assign n4957 = ~n4825 & n4956;
  assign n4958 = ~pi074 & ~n4818;
  assign n4959 = pi016 & n4801;
  assign n4960 = pi074 & n4959;
  assign n4961 = ~pi120 & n4960;
  assign n4962 = ~n4958 & ~n4961;
  assign n4963 = ~pi003 & ~n4962;
  assign n4964 = ~pi074 & n4843;
  assign n4965 = ~n4920 & ~n4964;
  assign n4966 = n4835 & ~n4965;
  assign n4967 = ~n4963 & ~n4966;
  assign n4968 = ~n4802 & ~n4903;
  assign n4969 = ~pi016 & pi074;
  assign n4970 = ~n4968 & n4969;
  assign n4971 = pi120 & n4970;
  assign n4972 = ~pi016 & n4864;
  assign n4973 = ~pi074 & n4972;
  assign n4974 = pi074 & n4816;
  assign n4975 = pi016 & n4920;
  assign n4976 = ~pi074 & n4975;
  assign n4977 = ~n4974 & ~n4976;
  assign n4978 = ~n4973 & n4977;
  assign n4979 = ~pi120 & ~n4978;
  assign n4980 = pi041 & n4905;
  assign n4981 = n4793 & n4980;
  assign n4982 = n4846 & n4890;
  assign n4983 = ~pi016 & n4801;
  assign n4984 = ~n4883 & ~n4983;
  assign n4985 = pi074 & n4796;
  assign n4986 = pi016 & n4985;
  assign n4987 = n4984 & ~n4986;
  assign n4988 = ~n4982 & n4987;
  assign n4989 = ~n4981 & n4988;
  assign n4990 = pi003 & ~n4989;
  assign n4991 = ~n4979 & ~n4990;
  assign n4992 = ~n4971 & n4991;
  assign n4993 = n4967 & n4992;
  assign n4994 = ~pi044 & ~n4993;
  assign n4995 = ~pi016 & n4806;
  assign n4996 = pi074 & n4995;
  assign n4997 = ~pi074 & n4794;
  assign n4998 = ~n4996 & ~n4997;
  assign n4999 = ~n4902 & ~n4914;
  assign n5000 = ~pi120 & ~n4999;
  assign n5001 = ~pi120 & n4828;
  assign n5002 = pi016 & n4814;
  assign n5003 = ~pi120 & n4830;
  assign n5004 = ~n5002 & ~n5003;
  assign n5005 = ~n5001 & n5004;
  assign n5006 = pi003 & ~n5005;
  assign n5007 = pi016 & pi074;
  assign n5008 = pi041 & n5007;
  assign n5009 = n4801 & n5008;
  assign n5010 = ~n4976 & ~n5009;
  assign n5011 = ~n4944 & n5010;
  assign n5012 = ~n4995 & n5011;
  assign n5013 = pi120 & ~n5012;
  assign n5014 = ~pi074 & n4828;
  assign n5015 = ~n4898 & ~n5014;
  assign n5016 = ~n4826 & n5015;
  assign n5017 = pi120 & ~n5016;
  assign n5018 = ~pi016 & n4805;
  assign n5019 = pi074 & n5018;
  assign n5020 = ~pi041 & pi074;
  assign n5021 = ~pi016 & n5020;
  assign n5022 = ~n4839 & ~n5021;
  assign n5023 = ~n5019 & n5022;
  assign n5024 = n4807 & n4890;
  assign n5025 = n5023 & ~n5024;
  assign n5026 = ~n5017 & n5025;
  assign n5027 = ~pi003 & ~n5026;
  assign n5028 = ~pi016 & ~pi045;
  assign n5029 = pi074 & n5028;
  assign n5030 = pi074 & n4903;
  assign n5031 = ~n5029 & ~n5030;
  assign n5032 = ~pi120 & ~n5031;
  assign n5033 = ~n5027 & ~n5032;
  assign n5034 = ~n5013 & n5033;
  assign n5035 = ~n5006 & n5034;
  assign n5036 = ~n5000 & n5035;
  assign n5037 = n4998 & n5036;
  assign n5038 = pi044 & ~n5037;
  assign n5039 = ~n4994 & ~n5038;
  assign n5040 = pi120 & ~n4855;
  assign n5041 = ~pi120 & ~n4986;
  assign n5042 = ~n5040 & ~n5041;
  assign n5043 = pi074 & n4806;
  assign n5044 = pi120 & n5043;
  assign n5045 = pi074 & n4803;
  assign n5046 = n4814 & n4901;
  assign n5047 = pi120 & ~n5046;
  assign n5048 = ~pi120 & ~n4845;
  assign n5049 = ~n5047 & ~n5048;
  assign n5050 = ~n5045 & ~n5049;
  assign n5051 = ~n5044 & n5050;
  assign n5052 = ~pi016 & ~pi074;
  assign n5053 = n4828 & n5052;
  assign n5054 = n5051 & ~n5053;
  assign n5055 = pi003 & ~n5054;
  assign n5056 = ~n5042 & ~n5055;
  assign n5057 = ~pi074 & n4814;
  assign n5058 = n4802 & n5052;
  assign n5059 = ~n5057 & ~n5058;
  assign n5060 = ~n4862 & n5059;
  assign n5061 = ~pi120 & ~n5060;
  assign n5062 = ~pi120 & n4969;
  assign n5063 = n4794 & n5062;
  assign n5064 = pi120 & n5009;
  assign n5065 = n4806 & n5052;
  assign n5066 = n4830 & n5052;
  assign n5067 = ~n5065 & ~n5066;
  assign n5068 = pi120 & ~n5067;
  assign n5069 = ~n5064 & ~n5068;
  assign n5070 = ~n5063 & n5069;
  assign n5071 = ~n5061 & n5070;
  assign n5072 = ~pi003 & ~n5071;
  assign n5073 = n5056 & ~n5072;
  assign n5074 = n5039 & n5073;
  assign n5075 = ~n4957 & n5074;
  assign n5076 = n4957 & ~n5074;
  assign n5077 = ~n5075 & ~n5076;
  assign n5078 = ~pi066 & ~pi103;
  assign n5079 = ~pi101 & n5078;
  assign n5080 = n4629 & n5079;
  assign n5081 = n4763 & n5078;
  assign n5082 = ~n5080 & ~n5081;
  assign n5083 = n4621 & ~n5082;
  assign n5084 = n4625 & n4668;
  assign n5085 = ~pi118 & n5084;
  assign n5086 = ~pi066 & n4774;
  assign n5087 = pi118 & n5086;
  assign n5088 = ~n5085 & ~n5087;
  assign n5089 = ~n5083 & n5088;
  assign n5090 = ~pi066 & ~pi118;
  assign n5091 = n4689 & n5090;
  assign n5092 = pi118 & n4725;
  assign n5093 = ~n5084 & ~n5092;
  assign n5094 = ~n5091 & n5093;
  assign n5095 = ~pi066 & n4622;
  assign n5096 = ~n4623 & ~n5095;
  assign n5097 = n5094 & n5096;
  assign n5098 = pi034 & ~n5097;
  assign n5099 = ~pi066 & n4638;
  assign n5100 = ~n4660 & ~n5099;
  assign n5101 = n4621 & ~n5100;
  assign n5102 = ~n4649 & ~n4687;
  assign n5103 = pi066 & ~pi103;
  assign n5104 = ~n5102 & n5103;
  assign n5105 = pi118 & n5104;
  assign n5106 = ~n5101 & ~n5105;
  assign n5107 = ~n5098 & n5106;
  assign n5108 = ~n4667 & ~n4704;
  assign n5109 = ~pi066 & ~n5108;
  assign n5110 = n4622 & n4668;
  assign n5111 = ~pi118 & n5110;
  assign n5112 = ~n5109 & ~n5111;
  assign n5113 = ~pi034 & ~n5112;
  assign n5114 = ~pi066 & n4733;
  assign n5115 = ~n4707 & ~n5114;
  assign n5116 = pi066 & n4626;
  assign n5117 = n5115 & ~n5116;
  assign n5118 = ~pi118 & ~n5117;
  assign n5119 = ~n5113 & ~n5118;
  assign n5120 = n5107 & n5119;
  assign n5121 = ~pi038 & ~n5120;
  assign n5122 = ~pi103 & n4630;
  assign n5123 = pi066 & n5122;
  assign n5124 = ~n4676 & ~n5123;
  assign n5125 = ~n4640 & ~n4651;
  assign n5126 = ~n4707 & n5125;
  assign n5127 = ~n5122 & n5126;
  assign n5128 = pi118 & ~n5127;
  assign n5129 = ~pi066 & pi103;
  assign n5130 = n4669 & n5129;
  assign n5131 = ~n4627 & ~n5130;
  assign n5132 = ~pi118 & ~n5131;
  assign n5133 = ~n5128 & ~n5132;
  assign n5134 = pi066 & n4687;
  assign n5135 = pi066 & n4746;
  assign n5136 = ~n5134 & ~n5135;
  assign n5137 = ~pi118 & ~n5136;
  assign n5138 = pi066 & ~pi101;
  assign n5139 = ~pi103 & n5138;
  assign n5140 = ~pi103 & n4629;
  assign n5141 = pi066 & n5140;
  assign n5142 = ~n5139 & ~n5141;
  assign n5143 = ~pi103 & n4669;
  assign n5144 = ~pi066 & n5143;
  assign n5145 = n5142 & ~n5144;
  assign n5146 = n4647 & n5090;
  assign n5147 = pi103 & n4675;
  assign n5148 = ~n4750 & ~n5147;
  assign n5149 = ~n4684 & n5148;
  assign n5150 = pi118 & ~n5149;
  assign n5151 = ~n5146 & ~n5150;
  assign n5152 = n5145 & n5151;
  assign n5153 = ~pi034 & ~n5152;
  assign n5154 = ~n5137 & ~n5153;
  assign n5155 = ~pi118 & n4763;
  assign n5156 = ~n4771 & ~n5155;
  assign n5157 = ~n4710 & n5156;
  assign n5158 = pi034 & ~n5157;
  assign n5159 = n5154 & ~n5158;
  assign n5160 = n5133 & n5159;
  assign n5161 = n5124 & n5160;
  assign n5162 = pi038 & ~n5161;
  assign n5163 = ~pi103 & n4649;
  assign n5164 = pi066 & n5163;
  assign n5165 = ~pi066 & n4759;
  assign n5166 = ~n5164 & ~n5165;
  assign n5167 = pi118 & n5129;
  assign n5168 = n4636 & n5167;
  assign n5169 = pi066 & n4630;
  assign n5170 = pi118 & n5169;
  assign n5171 = ~pi066 & n4736;
  assign n5172 = ~pi118 & n5171;
  assign n5173 = ~n5170 & ~n5172;
  assign n5174 = ~n5168 & n5173;
  assign n5175 = n5166 & n5174;
  assign n5176 = pi034 & ~n5175;
  assign n5177 = ~pi066 & n4636;
  assign n5178 = n4649 & n5078;
  assign n5179 = ~n5177 & ~n5178;
  assign n5180 = pi103 & n4635;
  assign n5181 = ~pi066 & n5180;
  assign n5182 = n5179 & ~n5181;
  assign n5183 = ~pi118 & ~n5182;
  assign n5184 = pi066 & n4774;
  assign n5185 = ~pi118 & n5184;
  assign n5186 = ~n5183 & ~n5185;
  assign n5187 = ~n4754 & n5186;
  assign n5188 = ~pi034 & ~n5187;
  assign n5189 = ~n5176 & ~n5188;
  assign n5190 = ~n5162 & n5189;
  assign n5191 = ~n5121 & n5190;
  assign n5192 = n5089 & n5191;
  assign n5193 = pi103 & n4659;
  assign n5194 = n5108 & ~n5193;
  assign n5195 = pi066 & ~n5194;
  assign n5196 = pi066 & n4649;
  assign n5197 = ~n5195 & ~n5196;
  assign n5198 = ~pi118 & ~n5197;
  assign n5199 = ~n4686 & ~n4725;
  assign n5200 = ~pi103 & n4625;
  assign n5201 = ~n5163 & ~n5200;
  assign n5202 = ~n4647 & n5201;
  assign n5203 = ~pi066 & ~n5202;
  assign n5204 = n5199 & ~n5203;
  assign n5205 = pi118 & ~n5204;
  assign n5206 = ~n5198 & ~n5205;
  assign n5207 = pi034 & ~n5206;
  assign n5208 = pi066 & n4643;
  assign n5209 = ~n5086 & ~n5208;
  assign n5210 = ~pi118 & ~n5209;
  assign n5211 = pi066 & n4684;
  assign n5212 = ~pi066 & n4764;
  assign n5213 = ~n5211 & ~n5212;
  assign n5214 = ~n4727 & n5213;
  assign n5215 = n4621 & ~n5214;
  assign n5216 = ~n4737 & ~n5144;
  assign n5217 = ~pi118 & ~n5216;
  assign n5218 = pi066 & n4690;
  assign n5219 = ~pi118 & n5218;
  assign n5220 = ~n5217 & ~n5219;
  assign n5221 = ~n5171 & n5220;
  assign n5222 = ~pi034 & ~n5221;
  assign n5223 = ~n5215 & ~n5222;
  assign n5224 = ~n5210 & n5223;
  assign n5225 = pi103 & n4689;
  assign n5226 = n4753 & n5225;
  assign n5227 = pi118 & n4642;
  assign n5228 = ~n5226 & ~n5227;
  assign n5229 = ~pi034 & ~n5228;
  assign n5230 = ~n4627 & ~n4650;
  assign n5231 = n4753 & ~n5230;
  assign n5232 = ~n4760 & ~n5231;
  assign n5233 = ~n5229 & n5232;
  assign n5234 = ~pi103 & pi119;
  assign n5235 = ~pi118 & n5234;
  assign n5236 = ~n4640 & ~n5235;
  assign n5237 = ~pi034 & ~n5236;
  assign n5238 = n5233 & ~n5237;
  assign n5239 = n4635 & n4668;
  assign n5240 = pi101 & n5239;
  assign n5241 = ~n4643 & ~n5240;
  assign n5242 = ~pi118 & ~n5241;
  assign n5243 = ~n5217 & ~n5242;
  assign n5244 = n5238 & n5243;
  assign n5245 = ~n4677 & ~n4685;
  assign n5246 = ~pi062 & n4668;
  assign n5247 = ~n4637 & ~n5246;
  assign n5248 = ~pi118 & ~n5247;
  assign n5249 = ~pi066 & pi118;
  assign n5250 = n4688 & n5249;
  assign n5251 = ~n5248 & ~n5250;
  assign n5252 = n5245 & n5251;
  assign n5253 = pi034 & ~n5252;
  assign n5254 = n5244 & ~n5253;
  assign n5255 = ~pi038 & ~n5254;
  assign n5256 = ~pi103 & n4687;
  assign n5257 = n4753 & n5256;
  assign n5258 = ~n5130 & ~n5257;
  assign n5259 = ~pi118 & n5181;
  assign n5260 = n5258 & ~n5259;
  assign n5261 = ~pi066 & n5200;
  assign n5262 = ~pi066 & n5193;
  assign n5263 = ~n5261 & ~n5262;
  assign n5264 = ~n5147 & n5263;
  assign n5265 = pi118 & ~n5264;
  assign n5266 = n5260 & ~n5265;
  assign n5267 = pi103 & n4732;
  assign n5268 = ~n4764 & ~n5267;
  assign n5269 = ~n5180 & n5268;
  assign n5270 = ~pi118 & ~n5269;
  assign n5271 = ~pi118 & n4675;
  assign n5272 = ~pi066 & n4690;
  assign n5273 = pi118 & n5272;
  assign n5274 = ~pi066 & n4635;
  assign n5275 = ~pi118 & n5274;
  assign n5276 = ~n5273 & ~n5275;
  assign n5277 = ~n5271 & n5276;
  assign n5278 = ~n5270 & n5277;
  assign n5279 = pi066 & n4775;
  assign n5280 = ~n5181 & ~n5279;
  assign n5281 = n5278 & n5280;
  assign n5282 = ~pi034 & ~n5281;
  assign n5283 = n4630 & n5090;
  assign n5284 = ~n5211 & ~n5283;
  assign n5285 = pi034 & ~n5284;
  assign n5286 = ~n5095 & ~n5267;
  assign n5287 = pi066 & n4635;
  assign n5288 = pi062 & ~pi103;
  assign n5289 = ~n5287 & ~n5288;
  assign n5290 = n5286 & n5289;
  assign n5291 = n4762 & ~n5290;
  assign n5292 = ~n5285 & ~n5291;
  assign n5293 = ~n5282 & n5292;
  assign n5294 = n5266 & n5293;
  assign n5295 = pi038 & ~n5294;
  assign n5296 = ~n5255 & ~n5295;
  assign n5297 = n5224 & n5296;
  assign n5298 = ~n5207 & n5297;
  assign n5299 = ~n5192 & n5298;
  assign n5300 = n5192 & ~n5298;
  assign n5301 = ~n5299 & ~n5300;
  assign n5302 = ~n5077 & n5301;
  assign n5303 = n4957 & n5074;
  assign n5304 = ~n4957 & ~n5074;
  assign n5305 = ~n5303 & ~n5304;
  assign n5306 = ~n5301 & ~n5305;
  assign n5307 = ~n5302 & ~n5306;
  assign n5308 = n4792 & n5307;
  assign n5309 = ~n4792 & ~n5307;
  assign n5310 = ~n5308 & ~n5309;
  assign n5311 = ~pi529 & n5310;
  assign po133 = n4285 | n5311;
  assign n5313 = ~pi185 & pi444;
  assign n5314 = pi185 & ~pi444;
  assign n5315 = ~n5313 & ~n5314;
  assign n5316 = pi529 & ~n5315;
  assign n5317 = pi077 & ~pi109;
  assign n5318 = ~pi043 & ~pi076;
  assign n5319 = pi070 & n5318;
  assign n5320 = n5317 & n5319;
  assign n5321 = ~pi077 & ~pi109;
  assign n5322 = ~pi070 & n5321;
  assign n5323 = pi076 & n5322;
  assign n5324 = pi043 & n5323;
  assign n5325 = ~n5320 & ~n5324;
  assign n5326 = ~pi122 & ~n5325;
  assign n5327 = pi070 & ~pi109;
  assign n5328 = ~pi076 & n5327;
  assign n5329 = ~pi043 & n5328;
  assign n5330 = pi077 & pi109;
  assign n5331 = pi070 & n5330;
  assign n5332 = ~pi043 & n5331;
  assign n5333 = ~n5329 & ~n5332;
  assign n5334 = ~pi122 & ~n5333;
  assign n5335 = pi070 & pi109;
  assign n5336 = pi076 & n5335;
  assign n5337 = ~pi043 & n5336;
  assign n5338 = ~pi070 & pi109;
  assign n5339 = ~pi076 & n5338;
  assign n5340 = pi043 & n5339;
  assign n5341 = ~pi122 & n5340;
  assign n5342 = ~n5337 & ~n5341;
  assign n5343 = ~n5334 & n5342;
  assign n5344 = ~pi039 & ~n5343;
  assign n5345 = ~pi070 & n5330;
  assign n5346 = pi076 & n5345;
  assign n5347 = pi043 & n5346;
  assign n5348 = pi043 & n5322;
  assign n5349 = pi070 & pi077;
  assign n5350 = pi076 & n5349;
  assign n5351 = ~pi043 & n5350;
  assign n5352 = ~n5348 & ~n5351;
  assign n5353 = ~n5347 & n5352;
  assign n5354 = ~pi039 & pi122;
  assign n5355 = ~n5353 & n5354;
  assign n5356 = ~n5344 & ~n5355;
  assign n5357 = ~n5326 & n5356;
  assign n5358 = ~pi043 & n5346;
  assign n5359 = ~pi077 & n5335;
  assign n5360 = pi043 & n5359;
  assign n5361 = ~n5358 & ~n5360;
  assign n5362 = ~pi043 & pi122;
  assign n5363 = ~pi070 & pi077;
  assign n5364 = pi076 & n5363;
  assign n5365 = n5362 & n5364;
  assign n5366 = pi043 & pi076;
  assign n5367 = ~pi077 & n5366;
  assign n5368 = ~pi070 & n5317;
  assign n5369 = pi043 & n5368;
  assign n5370 = ~n5367 & ~n5369;
  assign n5371 = ~pi122 & ~n5370;
  assign n5372 = ~n5365 & ~n5371;
  assign n5373 = n5361 & n5372;
  assign n5374 = pi039 & ~n5373;
  assign n5375 = pi070 & n5317;
  assign n5376 = pi076 & n5375;
  assign n5377 = pi043 & n5376;
  assign n5378 = ~n5323 & ~n5377;
  assign n5379 = ~pi122 & ~n5378;
  assign n5380 = ~n5334 & ~n5379;
  assign n5381 = pi043 & pi122;
  assign n5382 = ~pi070 & ~pi109;
  assign n5383 = ~pi076 & n5382;
  assign n5384 = ~pi077 & n5383;
  assign n5385 = n5381 & n5384;
  assign n5386 = pi076 & n5338;
  assign n5387 = n5381 & n5386;
  assign n5388 = pi122 & n5322;
  assign n5389 = ~n5387 & ~n5388;
  assign n5390 = ~pi039 & ~n5389;
  assign n5391 = pi070 & n5321;
  assign n5392 = pi076 & n5391;
  assign n5393 = pi076 & n5331;
  assign n5394 = ~n5392 & ~n5393;
  assign n5395 = n5381 & ~n5394;
  assign n5396 = ~n5390 & ~n5395;
  assign n5397 = ~n5385 & n5396;
  assign n5398 = ~pi076 & pi109;
  assign n5399 = ~pi122 & n5398;
  assign n5400 = ~pi076 & n5335;
  assign n5401 = pi043 & n5400;
  assign n5402 = ~n5399 & ~n5401;
  assign n5403 = ~pi039 & ~n5402;
  assign n5404 = n5397 & ~n5403;
  assign n5405 = n5380 & n5404;
  assign n5406 = ~n5374 & n5405;
  assign n5407 = ~pi017 & ~n5406;
  assign n5408 = n5357 & ~n5407;
  assign n5409 = pi076 & n5317;
  assign n5410 = ~pi043 & n5409;
  assign n5411 = ~pi122 & n5410;
  assign n5412 = ~pi070 & ~pi077;
  assign n5413 = pi076 & n5412;
  assign n5414 = ~n5350 & ~n5413;
  assign n5415 = ~n5409 & n5414;
  assign n5416 = ~pi122 & ~n5415;
  assign n5417 = ~pi122 & n5375;
  assign n5418 = ~pi043 & n5339;
  assign n5419 = pi122 & n5418;
  assign n5420 = ~pi043 & n5317;
  assign n5421 = ~pi122 & n5420;
  assign n5422 = ~n5419 & ~n5421;
  assign n5423 = ~n5417 & n5422;
  assign n5424 = ~n5416 & n5423;
  assign n5425 = pi070 & ~pi077;
  assign n5426 = ~pi076 & n5425;
  assign n5427 = pi043 & n5426;
  assign n5428 = ~n5410 & ~n5427;
  assign n5429 = n5424 & n5428;
  assign n5430 = ~pi039 & ~n5429;
  assign n5431 = pi076 & n5425;
  assign n5432 = ~pi043 & n5431;
  assign n5433 = ~pi076 & n5330;
  assign n5434 = ~pi043 & n5433;
  assign n5435 = ~n5376 & ~n5434;
  assign n5436 = ~n5432 & n5435;
  assign n5437 = pi122 & ~n5436;
  assign n5438 = ~pi043 & pi076;
  assign n5439 = n5327 & n5438;
  assign n5440 = ~pi076 & n5363;
  assign n5441 = n5381 & n5440;
  assign n5442 = ~n5439 & ~n5441;
  assign n5443 = ~n5437 & n5442;
  assign n5444 = ~pi043 & ~pi122;
  assign n5445 = ~pi077 & pi109;
  assign n5446 = ~pi070 & n5445;
  assign n5447 = n5444 & n5446;
  assign n5448 = ~n5347 & ~n5447;
  assign n5449 = pi039 & ~n5448;
  assign n5450 = ~pi076 & pi077;
  assign n5451 = pi043 & n5317;
  assign n5452 = ~pi043 & n5321;
  assign n5453 = ~n5413 & ~n5452;
  assign n5454 = ~n5451 & n5453;
  assign n5455 = ~n5450 & n5454;
  assign n5456 = pi039 & pi122;
  assign n5457 = ~n5455 & n5456;
  assign n5458 = ~n5449 & ~n5457;
  assign n5459 = n5443 & n5458;
  assign n5460 = ~n5430 & n5459;
  assign n5461 = ~n5411 & n5460;
  assign n5462 = pi017 & ~n5461;
  assign n5463 = pi043 & n5375;
  assign n5464 = ~pi076 & n5345;
  assign n5465 = ~n5463 & ~n5464;
  assign n5466 = pi076 & n5446;
  assign n5467 = ~pi076 & n5391;
  assign n5468 = ~n5466 & ~n5467;
  assign n5469 = ~n5433 & n5468;
  assign n5470 = ~pi043 & ~n5469;
  assign n5471 = n5465 & ~n5470;
  assign n5472 = pi122 & ~n5471;
  assign n5473 = pi043 & n5391;
  assign n5474 = ~pi076 & n5331;
  assign n5475 = ~pi076 & n5368;
  assign n5476 = ~n5431 & ~n5475;
  assign n5477 = ~n5474 & n5476;
  assign n5478 = pi043 & ~n5477;
  assign n5479 = ~n5473 & ~n5478;
  assign n5480 = ~pi122 & ~n5479;
  assign n5481 = ~n5472 & ~n5480;
  assign n5482 = pi039 & ~n5481;
  assign n5483 = ~n5462 & ~n5482;
  assign n5484 = n5408 & n5483;
  assign n5485 = pi043 & n5331;
  assign n5486 = pi076 & n5359;
  assign n5487 = ~pi043 & n5486;
  assign n5488 = ~n5485 & ~n5487;
  assign n5489 = ~n5418 & n5488;
  assign n5490 = ~pi122 & ~n5489;
  assign n5491 = ~pi076 & n5375;
  assign n5492 = pi043 & n5491;
  assign n5493 = pi043 & n5345;
  assign n5494 = ~pi122 & n5322;
  assign n5495 = ~pi043 & n5425;
  assign n5496 = ~n5359 & ~n5495;
  assign n5497 = ~n5386 & n5496;
  assign n5498 = pi122 & ~n5497;
  assign n5499 = ~n5494 & ~n5498;
  assign n5500 = ~n5493 & n5499;
  assign n5501 = ~n5486 & n5500;
  assign n5502 = ~n5337 & ~n5421;
  assign n5503 = n5501 & n5502;
  assign n5504 = pi039 & ~n5503;
  assign n5505 = ~n5492 & ~n5504;
  assign n5506 = ~n5490 & n5505;
  assign n5507 = ~pi043 & n5345;
  assign n5508 = ~n5369 & ~n5507;
  assign n5509 = ~pi122 & ~n5508;
  assign n5510 = pi122 & n5375;
  assign n5511 = n5318 & n5349;
  assign n5512 = ~pi076 & n5321;
  assign n5513 = ~pi043 & n5512;
  assign n5514 = ~n5511 & ~n5513;
  assign n5515 = ~n5510 & n5514;
  assign n5516 = pi043 & n5466;
  assign n5517 = pi043 & n5446;
  assign n5518 = pi122 & n5517;
  assign n5519 = ~n5516 & ~n5518;
  assign n5520 = n5515 & n5519;
  assign n5521 = pi122 & n5328;
  assign n5522 = n5520 & ~n5521;
  assign n5523 = ~n5509 & n5522;
  assign n5524 = ~pi039 & ~n5523;
  assign n5525 = n5506 & ~n5524;
  assign n5526 = pi043 & n5445;
  assign n5527 = pi076 & n5526;
  assign n5528 = ~n5368 & ~n5446;
  assign n5529 = pi076 & ~n5528;
  assign n5530 = ~n5527 & ~n5529;
  assign n5531 = pi122 & ~n5530;
  assign n5532 = n5525 & ~n5531;
  assign n5533 = pi017 & ~n5532;
  assign n5534 = ~pi043 & n5393;
  assign n5535 = pi043 & n5409;
  assign n5536 = ~n5534 & ~n5535;
  assign n5537 = ~pi122 & ~n5536;
  assign n5538 = pi043 & ~pi122;
  assign n5539 = n5486 & n5538;
  assign n5540 = ~n5330 & ~n5335;
  assign n5541 = n5362 & ~n5540;
  assign n5542 = pi122 & n5321;
  assign n5543 = pi076 & n5542;
  assign n5544 = ~n5541 & ~n5543;
  assign n5545 = ~n5323 & ~n5418;
  assign n5546 = n5544 & n5545;
  assign n5547 = ~n5539 & n5546;
  assign n5548 = ~pi039 & ~n5547;
  assign n5549 = n5381 & n5383;
  assign n5550 = ~pi043 & n5475;
  assign n5551 = pi122 & n5474;
  assign n5552 = ~n5550 & ~n5551;
  assign n5553 = ~n5549 & n5552;
  assign n5554 = ~n5548 & n5553;
  assign n5555 = ~n5537 & n5554;
  assign n5556 = ~pi076 & n5359;
  assign n5557 = ~pi122 & n5556;
  assign n5558 = pi043 & n5393;
  assign n5559 = ~n5517 & ~n5558;
  assign n5560 = ~pi043 & n5474;
  assign n5561 = n5559 & ~n5560;
  assign n5562 = ~pi043 & n5376;
  assign n5563 = ~n5383 & ~n5562;
  assign n5564 = pi122 & ~n5563;
  assign n5565 = n5561 & ~n5564;
  assign n5566 = ~n5557 & n5565;
  assign n5567 = pi039 & ~n5566;
  assign n5568 = n5555 & ~n5567;
  assign n5569 = ~pi017 & ~n5568;
  assign n5570 = n5366 & n5368;
  assign n5571 = ~pi043 & n5323;
  assign n5572 = pi122 & n5571;
  assign n5573 = n5362 & n5475;
  assign n5574 = ~n5572 & ~n5573;
  assign n5575 = ~pi039 & ~n5574;
  assign n5576 = n5381 & n5464;
  assign n5577 = pi122 & n5516;
  assign n5578 = ~n5576 & ~n5577;
  assign n5579 = ~n5575 & n5578;
  assign n5580 = ~n5570 & n5579;
  assign n5581 = pi122 & n5486;
  assign n5582 = ~pi076 & n5317;
  assign n5583 = ~n5556 & ~n5582;
  assign n5584 = ~n5413 & n5583;
  assign n5585 = n5444 & ~n5584;
  assign n5586 = ~pi076 & n5446;
  assign n5587 = pi043 & n5586;
  assign n5588 = ~pi122 & n5587;
  assign n5589 = ~n5585 & ~n5588;
  assign n5590 = ~n5581 & n5589;
  assign n5591 = pi039 & ~n5590;
  assign n5592 = pi043 & n5433;
  assign n5593 = ~pi039 & ~pi122;
  assign n5594 = n5592 & n5593;
  assign n5595 = ~n5591 & ~n5594;
  assign n5596 = pi043 & ~pi076;
  assign n5597 = n5349 & n5596;
  assign n5598 = ~n5493 & ~n5597;
  assign n5599 = n5456 & ~n5598;
  assign n5600 = n5595 & ~n5599;
  assign n5601 = n5580 & n5600;
  assign n5602 = ~n5569 & n5601;
  assign n5603 = ~n5533 & n5602;
  assign n5604 = n5484 & n5603;
  assign n5605 = ~n5484 & ~n5603;
  assign n5606 = ~n5604 & ~n5605;
  assign n5607 = pi005 & pi091;
  assign n5608 = ~pi052 & ~pi084;
  assign n5609 = ~pi094 & n5608;
  assign n5610 = ~pi004 & n5609;
  assign n5611 = n5607 & n5610;
  assign n5612 = pi084 & ~pi094;
  assign n5613 = ~pi004 & n5612;
  assign n5614 = ~pi005 & n5613;
  assign n5615 = pi052 & pi094;
  assign n5616 = pi084 & n5615;
  assign n5617 = ~pi005 & n5616;
  assign n5618 = ~n5614 & ~n5617;
  assign n5619 = ~pi091 & ~n5618;
  assign n5620 = pi052 & ~pi094;
  assign n5621 = pi084 & n5620;
  assign n5622 = pi004 & n5621;
  assign n5623 = pi005 & n5622;
  assign n5624 = pi004 & n5609;
  assign n5625 = ~n5623 & ~n5624;
  assign n5626 = ~pi091 & ~n5625;
  assign n5627 = ~n5619 & ~n5626;
  assign n5628 = ~pi004 & pi094;
  assign n5629 = ~pi091 & n5628;
  assign n5630 = pi084 & pi094;
  assign n5631 = ~pi004 & n5630;
  assign n5632 = pi005 & n5631;
  assign n5633 = ~n5629 & ~n5632;
  assign n5634 = ~pi024 & ~n5633;
  assign n5635 = ~pi052 & ~pi094;
  assign n5636 = pi084 & n5635;
  assign n5637 = pi004 & n5636;
  assign n5638 = pi004 & n5616;
  assign n5639 = ~n5637 & ~n5638;
  assign n5640 = n5607 & ~n5639;
  assign n5641 = ~pi018 & ~n5640;
  assign n5642 = ~n5634 & n5641;
  assign n5643 = ~pi084 & pi094;
  assign n5644 = pi004 & n5643;
  assign n5645 = n5607 & n5644;
  assign n5646 = pi091 & n5609;
  assign n5647 = ~n5645 & ~n5646;
  assign n5648 = ~pi024 & ~n5647;
  assign n5649 = n5642 & ~n5648;
  assign n5650 = ~pi084 & n5615;
  assign n5651 = pi004 & n5650;
  assign n5652 = ~pi005 & n5651;
  assign n5653 = ~pi052 & pi094;
  assign n5654 = pi084 & n5653;
  assign n5655 = pi005 & n5654;
  assign n5656 = ~n5652 & ~n5655;
  assign n5657 = pi005 & ~pi052;
  assign n5658 = pi004 & n5657;
  assign n5659 = ~pi084 & n5620;
  assign n5660 = pi005 & n5659;
  assign n5661 = ~n5658 & ~n5660;
  assign n5662 = ~pi091 & ~n5661;
  assign n5663 = ~pi005 & pi091;
  assign n5664 = pi052 & ~pi084;
  assign n5665 = pi004 & n5664;
  assign n5666 = n5663 & n5665;
  assign n5667 = ~n5662 & ~n5666;
  assign n5668 = n5656 & n5667;
  assign n5669 = pi024 & ~n5668;
  assign n5670 = n5649 & ~n5669;
  assign n5671 = n5627 & n5670;
  assign n5672 = ~n5611 & n5671;
  assign n5673 = pi004 & n5620;
  assign n5674 = ~pi005 & n5673;
  assign n5675 = ~pi091 & n5674;
  assign n5676 = pi004 & n5608;
  assign n5677 = pi052 & pi084;
  assign n5678 = pi004 & n5677;
  assign n5679 = ~n5676 & ~n5678;
  assign n5680 = ~n5673 & n5679;
  assign n5681 = ~pi091 & ~n5680;
  assign n5682 = ~pi091 & n5621;
  assign n5683 = ~pi004 & n5643;
  assign n5684 = ~pi005 & n5683;
  assign n5685 = pi091 & n5684;
  assign n5686 = ~pi091 & n5620;
  assign n5687 = ~pi005 & n5686;
  assign n5688 = ~n5685 & ~n5687;
  assign n5689 = ~n5682 & n5688;
  assign n5690 = ~n5681 & n5689;
  assign n5691 = ~pi052 & pi084;
  assign n5692 = ~pi004 & n5691;
  assign n5693 = pi005 & n5692;
  assign n5694 = ~n5674 & ~n5693;
  assign n5695 = n5690 & n5694;
  assign n5696 = ~pi024 & ~n5695;
  assign n5697 = pi024 & pi091;
  assign n5698 = ~pi005 & n5635;
  assign n5699 = ~n5676 & ~n5698;
  assign n5700 = pi005 & n5620;
  assign n5701 = ~pi004 & pi052;
  assign n5702 = ~n5700 & ~n5701;
  assign n5703 = n5699 & n5702;
  assign n5704 = n5697 & ~n5703;
  assign n5705 = ~pi005 & ~pi091;
  assign n5706 = ~pi084 & n5653;
  assign n5707 = n5705 & n5706;
  assign n5708 = pi005 & n5651;
  assign n5709 = ~n5707 & ~n5708;
  assign n5710 = pi024 & ~n5709;
  assign n5711 = ~n5704 & ~n5710;
  assign n5712 = ~pi004 & n5615;
  assign n5713 = ~pi005 & n5712;
  assign n5714 = pi004 & n5691;
  assign n5715 = ~pi005 & n5714;
  assign n5716 = ~n5713 & ~n5715;
  assign n5717 = ~n5622 & n5716;
  assign n5718 = pi091 & ~n5717;
  assign n5719 = pi004 & ~pi005;
  assign n5720 = n5612 & n5719;
  assign n5721 = ~pi004 & n5664;
  assign n5722 = n5607 & n5721;
  assign n5723 = ~n5720 & ~n5722;
  assign n5724 = ~n5718 & n5723;
  assign n5725 = n5711 & n5724;
  assign n5726 = ~n5696 & n5725;
  assign n5727 = ~n5675 & n5726;
  assign n5728 = pi018 & n5727;
  assign n5729 = ~n5672 & ~n5728;
  assign n5730 = ~pi004 & ~pi005;
  assign n5731 = pi084 & n5730;
  assign n5732 = n5620 & n5731;
  assign n5733 = pi005 & n5624;
  assign n5734 = ~n5732 & ~n5733;
  assign n5735 = ~pi091 & ~n5734;
  assign n5736 = ~pi024 & pi091;
  assign n5737 = ~pi005 & n5678;
  assign n5738 = ~n5708 & ~n5737;
  assign n5739 = pi005 & n5609;
  assign n5740 = n5738 & ~n5739;
  assign n5741 = n5736 & ~n5740;
  assign n5742 = pi005 & n5683;
  assign n5743 = ~pi091 & n5742;
  assign n5744 = ~n5619 & ~n5743;
  assign n5745 = pi004 & n5630;
  assign n5746 = ~pi005 & n5745;
  assign n5747 = n5744 & ~n5746;
  assign n5748 = ~pi024 & ~n5747;
  assign n5749 = ~n5741 & ~n5748;
  assign n5750 = ~n5735 & n5749;
  assign n5751 = pi005 & n5621;
  assign n5752 = ~pi004 & n5650;
  assign n5753 = ~n5751 & ~n5752;
  assign n5754 = ~pi004 & n5636;
  assign n5755 = ~n5712 & ~n5754;
  assign n5756 = pi004 & n5706;
  assign n5757 = n5755 & ~n5756;
  assign n5758 = ~pi005 & ~n5757;
  assign n5759 = n5753 & ~n5758;
  assign n5760 = pi091 & ~n5759;
  assign n5761 = ~pi004 & n5659;
  assign n5762 = ~pi004 & n5616;
  assign n5763 = ~n5761 & ~n5762;
  assign n5764 = ~n5714 & n5763;
  assign n5765 = pi005 & ~n5764;
  assign n5766 = pi005 & n5636;
  assign n5767 = ~n5765 & ~n5766;
  assign n5768 = ~pi091 & ~n5767;
  assign n5769 = ~n5760 & ~n5768;
  assign n5770 = pi024 & ~n5769;
  assign n5771 = n5750 & ~n5770;
  assign n5772 = ~n5729 & n5771;
  assign n5773 = pi004 & n5654;
  assign n5774 = pi005 & n5650;
  assign n5775 = ~n5773 & ~n5774;
  assign n5776 = ~pi005 & n5691;
  assign n5777 = ~n5654 & ~n5776;
  assign n5778 = ~n5644 & n5777;
  assign n5779 = pi091 & ~n5778;
  assign n5780 = n5775 & ~n5779;
  assign n5781 = ~pi091 & n5609;
  assign n5782 = n5780 & ~n5781;
  assign n5783 = ~n5687 & ~n5746;
  assign n5784 = n5782 & n5783;
  assign n5785 = pi024 & ~n5784;
  assign n5786 = ~pi005 & n5773;
  assign n5787 = ~n5684 & ~n5786;
  assign n5788 = pi005 & n5616;
  assign n5789 = n5787 & ~n5788;
  assign n5790 = ~pi091 & ~n5789;
  assign n5791 = pi091 & n5613;
  assign n5792 = pi091 & n5621;
  assign n5793 = ~n5791 & ~n5792;
  assign n5794 = pi005 & n5706;
  assign n5795 = pi091 & n5794;
  assign n5796 = pi004 & pi005;
  assign n5797 = n5706 & n5796;
  assign n5798 = ~pi005 & n5650;
  assign n5799 = ~n5660 & ~n5798;
  assign n5800 = ~pi091 & ~n5799;
  assign n5801 = ~n5797 & ~n5800;
  assign n5802 = ~n5795 & n5801;
  assign n5803 = n5793 & n5802;
  assign n5804 = ~pi004 & ~pi052;
  assign n5805 = ~pi094 & n5804;
  assign n5806 = ~pi005 & n5805;
  assign n5807 = n5677 & n5730;
  assign n5808 = ~n5806 & ~n5807;
  assign n5809 = n5803 & n5808;
  assign n5810 = ~pi024 & ~n5809;
  assign n5811 = ~pi004 & pi005;
  assign n5812 = n5621 & n5811;
  assign n5813 = ~n5810 & ~n5812;
  assign n5814 = ~n5790 & n5813;
  assign n5815 = ~n5785 & n5814;
  assign n5816 = ~n5659 & ~n5706;
  assign n5817 = pi004 & ~n5816;
  assign n5818 = pi005 & n5653;
  assign n5819 = pi004 & n5818;
  assign n5820 = ~n5817 & ~n5819;
  assign n5821 = pi091 & ~n5820;
  assign n5822 = n5815 & ~n5821;
  assign n5823 = pi018 & ~n5822;
  assign n5824 = ~pi005 & n5761;
  assign n5825 = ~pi005 & n5638;
  assign n5826 = pi005 & n5673;
  assign n5827 = ~n5825 & ~n5826;
  assign n5828 = ~pi091 & ~n5827;
  assign n5829 = pi091 & n5762;
  assign n5830 = ~pi084 & ~pi094;
  assign n5831 = ~pi004 & n5830;
  assign n5832 = n5607 & n5831;
  assign n5833 = ~n5829 & ~n5832;
  assign n5834 = ~n5828 & n5833;
  assign n5835 = ~n5824 & n5834;
  assign n5836 = pi005 & ~pi091;
  assign n5837 = n5773 & n5836;
  assign n5838 = ~n5624 & ~n5684;
  assign n5839 = pi004 & n5635;
  assign n5840 = pi091 & n5839;
  assign n5841 = ~n5615 & ~n5630;
  assign n5842 = n5663 & ~n5841;
  assign n5843 = ~n5840 & ~n5842;
  assign n5844 = n5838 & n5843;
  assign n5845 = ~n5837 & n5844;
  assign n5846 = ~pi024 & ~n5845;
  assign n5847 = n5835 & ~n5846;
  assign n5848 = ~pi005 & n5762;
  assign n5849 = ~n5794 & ~n5848;
  assign n5850 = ~pi004 & n5654;
  assign n5851 = ~pi091 & n5850;
  assign n5852 = ~pi005 & n5622;
  assign n5853 = ~n5831 & ~n5852;
  assign n5854 = pi091 & ~n5853;
  assign n5855 = ~n5851 & ~n5854;
  assign n5856 = pi005 & n5638;
  assign n5857 = n5855 & ~n5856;
  assign n5858 = n5849 & n5857;
  assign n5859 = pi024 & ~n5858;
  assign n5860 = n5847 & ~n5859;
  assign n5861 = ~pi018 & ~n5860;
  assign n5862 = ~n5823 & ~n5861;
  assign n5863 = ~pi024 & ~pi091;
  assign n5864 = pi005 & n5712;
  assign n5865 = n5863 & n5864;
  assign n5866 = ~pi004 & n5706;
  assign n5867 = pi005 & n5866;
  assign n5868 = ~pi091 & n5867;
  assign n5869 = pi091 & n5773;
  assign n5870 = ~n5868 & ~n5869;
  assign n5871 = ~n5676 & ~n5850;
  assign n5872 = ~pi004 & n5620;
  assign n5873 = n5871 & ~n5872;
  assign n5874 = n5705 & ~n5873;
  assign n5875 = n5870 & ~n5874;
  assign n5876 = pi024 & ~n5875;
  assign n5877 = ~n5865 & ~n5876;
  assign n5878 = n5677 & n5811;
  assign n5879 = ~n5774 & ~n5878;
  assign n5880 = n5697 & ~n5879;
  assign n5881 = n5877 & ~n5880;
  assign n5882 = n5609 & n5719;
  assign n5883 = pi091 & n5882;
  assign n5884 = n5663 & n5761;
  assign n5885 = ~n5883 & ~n5884;
  assign n5886 = ~pi024 & ~n5885;
  assign n5887 = n5607 & n5756;
  assign n5888 = pi005 & n5752;
  assign n5889 = pi091 & n5888;
  assign n5890 = ~n5887 & ~n5889;
  assign n5891 = n5659 & n5796;
  assign n5892 = n5890 & ~n5891;
  assign n5893 = ~n5886 & n5892;
  assign n5894 = n5881 & n5893;
  assign n5895 = n5862 & n5894;
  assign n5896 = n5772 & ~n5895;
  assign n5897 = ~n5772 & n5895;
  assign n5898 = ~n5896 & ~n5897;
  assign n5899 = n5606 & n5898;
  assign n5900 = ~n5606 & ~n5898;
  assign n5901 = ~n5899 & ~n5900;
  assign n5902 = pi055 & ~pi124;
  assign n5903 = pi125 & n5902;
  assign n5904 = ~pi009 & n5903;
  assign n5905 = pi113 & n5904;
  assign n5906 = ~pi025 & pi055;
  assign n5907 = ~pi025 & pi124;
  assign n5908 = ~n5906 & ~n5907;
  assign n5909 = pi009 & ~n5908;
  assign n5910 = pi055 & pi124;
  assign n5911 = pi025 & n5910;
  assign n5912 = ~pi125 & n5911;
  assign n5913 = ~pi009 & n5912;
  assign n5914 = ~n5909 & ~n5913;
  assign n5915 = ~pi055 & ~pi124;
  assign n5916 = ~pi025 & n5915;
  assign n5917 = ~pi009 & ~pi125;
  assign n5918 = n5916 & n5917;
  assign n5919 = n5914 & ~n5918;
  assign n5920 = ~pi113 & ~n5919;
  assign n5921 = pi025 & n5915;
  assign n5922 = pi009 & n5921;
  assign n5923 = pi113 & n5922;
  assign n5924 = ~pi025 & n5910;
  assign n5925 = pi125 & n5924;
  assign n5926 = pi009 & n5925;
  assign n5927 = ~n5923 & ~n5926;
  assign n5928 = ~pi055 & pi124;
  assign n5929 = ~pi025 & n5928;
  assign n5930 = ~pi125 & n5929;
  assign n5931 = pi009 & n5930;
  assign n5932 = n5927 & ~n5931;
  assign n5933 = ~n5920 & n5932;
  assign n5934 = ~n5905 & n5933;
  assign n5935 = pi096 & ~n5934;
  assign n5936 = pi025 & pi055;
  assign n5937 = pi125 & n5936;
  assign n5938 = pi009 & pi113;
  assign n5939 = n5937 & n5938;
  assign n5940 = ~pi025 & n5902;
  assign n5941 = ~pi125 & n5940;
  assign n5942 = pi009 & n5941;
  assign n5943 = ~pi113 & n5942;
  assign n5944 = ~n5939 & ~n5943;
  assign n5945 = ~n5935 & n5944;
  assign n5946 = ~pi113 & n5925;
  assign n5947 = ~pi009 & n5946;
  assign n5948 = pi025 & n5928;
  assign n5949 = ~pi009 & n5948;
  assign n5950 = ~n5930 & ~n5949;
  assign n5951 = pi125 & n5948;
  assign n5952 = n5950 & ~n5951;
  assign n5953 = ~pi113 & ~n5952;
  assign n5954 = ~pi124 & n5936;
  assign n5955 = pi113 & n5954;
  assign n5956 = pi009 & n5903;
  assign n5957 = ~n5955 & ~n5956;
  assign n5958 = ~pi009 & pi113;
  assign n5959 = pi125 & n5907;
  assign n5960 = n5958 & n5959;
  assign n5961 = n5957 & ~n5960;
  assign n5962 = ~n5953 & n5961;
  assign n5963 = pi096 & ~n5962;
  assign n5964 = ~pi125 & n5921;
  assign n5965 = ~pi009 & n5964;
  assign n5966 = ~pi009 & ~pi113;
  assign n5967 = ~pi124 & n5966;
  assign n5968 = n5936 & n5967;
  assign n5969 = ~pi125 & n5915;
  assign n5970 = pi009 & n5969;
  assign n5971 = pi113 & n5916;
  assign n5972 = ~n5970 & ~n5971;
  assign n5973 = pi113 & n5937;
  assign n5974 = n5972 & ~n5973;
  assign n5975 = ~n5968 & n5974;
  assign n5976 = ~pi096 & ~n5975;
  assign n5977 = ~n5965 & ~n5976;
  assign n5978 = pi009 & pi125;
  assign n5979 = n5916 & n5978;
  assign n5980 = ~pi125 & n5906;
  assign n5981 = ~pi009 & n5980;
  assign n5982 = ~n5979 & ~n5981;
  assign n5983 = pi113 & ~n5982;
  assign n5984 = n5977 & ~n5983;
  assign n5985 = ~n5963 & n5984;
  assign n5986 = ~n5947 & n5985;
  assign n5987 = pi010 & ~n5986;
  assign n5988 = n5945 & ~n5987;
  assign n5989 = pi009 & ~pi125;
  assign n5990 = ~pi055 & n5989;
  assign n5991 = pi009 & n5929;
  assign n5992 = ~n5990 & ~n5991;
  assign n5993 = pi113 & ~n5992;
  assign n5994 = ~pi009 & pi125;
  assign n5995 = ~pi124 & n5994;
  assign n5996 = ~n5912 & ~n5995;
  assign n5997 = pi113 & ~n5996;
  assign n5998 = ~n5993 & ~n5997;
  assign n5999 = pi125 & n5916;
  assign n6000 = ~pi009 & n5999;
  assign n6001 = pi009 & n5964;
  assign n6002 = ~n6000 & ~n6001;
  assign n6003 = ~pi125 & n5902;
  assign n6004 = pi125 & n5929;
  assign n6005 = ~n6003 & ~n6004;
  assign n6006 = ~pi113 & ~n6005;
  assign n6007 = ~pi125 & n5928;
  assign n6008 = pi113 & n6007;
  assign n6009 = ~n6006 & ~n6008;
  assign n6010 = n6002 & n6009;
  assign n6011 = pi096 & ~n6010;
  assign n6012 = pi025 & pi124;
  assign n6013 = ~pi125 & n6012;
  assign n6014 = ~pi113 & n6013;
  assign n6015 = ~pi125 & n5910;
  assign n6016 = pi009 & n6015;
  assign n6017 = n5915 & n5978;
  assign n6018 = ~pi113 & n6017;
  assign n6019 = pi009 & n6012;
  assign n6020 = ~n6018 & ~n6019;
  assign n6021 = ~n6016 & n6020;
  assign n6022 = ~n6014 & n6021;
  assign n6023 = pi113 & n5951;
  assign n6024 = n6022 & ~n6023;
  assign n6025 = ~pi096 & ~n6024;
  assign n6026 = pi009 & n6003;
  assign n6027 = pi009 & n5924;
  assign n6028 = ~n6026 & ~n6027;
  assign n6029 = ~n5918 & n6028;
  assign n6030 = ~pi113 & ~n6029;
  assign n6031 = ~n6025 & ~n6030;
  assign n6032 = ~n6011 & n6031;
  assign n6033 = n5998 & n6032;
  assign n6034 = ~pi010 & ~n6033;
  assign n6035 = ~pi009 & n5921;
  assign n6036 = ~n5917 & ~n5978;
  assign n6037 = n5929 & ~n6036;
  assign n6038 = pi025 & ~pi055;
  assign n6039 = ~pi125 & n6038;
  assign n6040 = pi009 & n6039;
  assign n6041 = pi009 & n5954;
  assign n6042 = ~n6040 & ~n6041;
  assign n6043 = ~n6037 & n6042;
  assign n6044 = ~n6035 & n6043;
  assign n6045 = pi113 & ~n6044;
  assign n6046 = pi125 & n5954;
  assign n6047 = pi009 & n6046;
  assign n6048 = ~n5965 & ~n6047;
  assign n6049 = pi125 & n5906;
  assign n6050 = ~pi009 & n6049;
  assign n6051 = pi009 & n5912;
  assign n6052 = ~n6050 & ~n6051;
  assign n6053 = ~pi009 & n5924;
  assign n6054 = n6052 & ~n6053;
  assign n6055 = ~pi113 & ~n6054;
  assign n6056 = n6048 & ~n6055;
  assign n6057 = ~n6045 & n6056;
  assign n6058 = ~pi096 & ~n6057;
  assign n6059 = ~n6034 & ~n6058;
  assign n6060 = n5988 & n6059;
  assign n6061 = ~pi185 & ~n6060;
  assign n6062 = pi185 & n6060;
  assign n6063 = ~n6061 & ~n6062;
  assign n6064 = pi122 & n5410;
  assign n6065 = pi122 & n5473;
  assign n6066 = ~n6064 & ~n6065;
  assign n6067 = pi039 & n6066;
  assign n6068 = ~pi070 & n5318;
  assign n6069 = n5445 & n6068;
  assign n6070 = ~n5516 & ~n6069;
  assign n6071 = ~pi043 & n5391;
  assign n6072 = ~n5427 & ~n6071;
  assign n6073 = ~n5463 & n6072;
  assign n6074 = n6070 & n6073;
  assign n6075 = pi122 & ~n6074;
  assign n6076 = ~pi043 & n5364;
  assign n6077 = pi043 & n5474;
  assign n6078 = ~n6076 & ~n6077;
  assign n6079 = ~n5507 & n6078;
  assign n6080 = ~pi122 & ~n6079;
  assign n6081 = ~n5377 & ~n6080;
  assign n6082 = ~n6075 & n6081;
  assign n6083 = n5318 & n5391;
  assign n6084 = ~pi039 & ~n6083;
  assign n6085 = n6082 & n6084;
  assign n6086 = ~n6067 & ~n6085;
  assign n6087 = ~n5486 & ~n5586;
  assign n6088 = ~pi043 & n5359;
  assign n6089 = n6087 & ~n6088;
  assign n6090 = ~pi122 & ~n6089;
  assign n6091 = ~n5510 & ~n5535;
  assign n6092 = n5362 & n5386;
  assign n6093 = n6091 & ~n6092;
  assign n6094 = ~n6090 & n6093;
  assign n6095 = pi039 & ~n6094;
  assign n6096 = ~pi122 & n5358;
  assign n6097 = pi043 & n5512;
  assign n6098 = ~n5388 & ~n6097;
  assign n6099 = pi122 & n5350;
  assign n6100 = ~pi043 & n5375;
  assign n6101 = ~pi122 & n6100;
  assign n6102 = ~n6099 & ~n6101;
  assign n6103 = n6098 & n6102;
  assign n6104 = ~pi039 & ~n6103;
  assign n6105 = ~n6096 & ~n6104;
  assign n6106 = ~n6095 & n6105;
  assign n6107 = ~pi043 & n5440;
  assign n6108 = ~n5324 & ~n6107;
  assign n6109 = pi122 & ~n6108;
  assign n6110 = ~n6083 & ~n6109;
  assign n6111 = n6106 & n6110;
  assign n6112 = ~pi017 & ~n6111;
  assign n6113 = ~n5338 & ~n5363;
  assign n6114 = pi043 & ~n6113;
  assign n6115 = ~n5560 & ~n6114;
  assign n6116 = n5321 & n6068;
  assign n6117 = n6115 & ~n6116;
  assign n6118 = ~pi122 & ~n6117;
  assign n6119 = ~n5587 & ~n6118;
  assign n6120 = ~n5347 & n6119;
  assign n6121 = pi039 & ~n6120;
  assign n6122 = ~n6112 & ~n6121;
  assign n6123 = ~n6086 & n6122;
  assign n6124 = pi122 & n5349;
  assign n6125 = n5366 & n6124;
  assign n6126 = n5475 & n5538;
  assign n6127 = ~n6125 & ~n6126;
  assign n6128 = ~pi077 & n5596;
  assign n6129 = ~n5517 & ~n6128;
  assign n6130 = pi122 & ~n6129;
  assign n6131 = n5321 & n5366;
  assign n6132 = ~pi122 & n6131;
  assign n6133 = pi043 & n5335;
  assign n6134 = ~n6132 & ~n6133;
  assign n6135 = ~pi122 & n5400;
  assign n6136 = ~n5592 & ~n6135;
  assign n6137 = n6134 & n6136;
  assign n6138 = ~n5581 & n6137;
  assign n6139 = ~pi039 & ~n6138;
  assign n6140 = pi043 & n5467;
  assign n6141 = ~n5571 & ~n6140;
  assign n6142 = ~pi076 & n5445;
  assign n6143 = pi122 & n6142;
  assign n6144 = ~n5466 & ~n5582;
  assign n6145 = ~pi122 & ~n6144;
  assign n6146 = ~n6143 & ~n6145;
  assign n6147 = n6141 & n6146;
  assign n6148 = pi039 & ~n6147;
  assign n6149 = ~n6139 & ~n6148;
  assign n6150 = ~pi043 & ~pi109;
  assign n6151 = pi076 & n6150;
  assign n6152 = ~n5474 & ~n6151;
  assign n6153 = pi122 & ~n6152;
  assign n6154 = pi043 & n5582;
  assign n6155 = ~n5493 & ~n6154;
  assign n6156 = ~n6116 & n6155;
  assign n6157 = ~pi122 & ~n6156;
  assign n6158 = ~n6153 & ~n6157;
  assign n6159 = n6149 & n6158;
  assign n6160 = ~n6130 & n6159;
  assign n6161 = pi017 & ~n6160;
  assign n6162 = n6127 & ~n6161;
  assign n6163 = n6123 & n6162;
  assign n6164 = pi031 & ~pi035;
  assign n6165 = pi100 & pi128;
  assign n6166 = ~pi037 & n6165;
  assign n6167 = n6164 & n6166;
  assign n6168 = ~pi106 & n6167;
  assign n6169 = ~pi100 & pi128;
  assign n6170 = pi037 & n6169;
  assign n6171 = ~pi035 & n6170;
  assign n6172 = ~pi037 & n6169;
  assign n6173 = ~pi031 & n6172;
  assign n6174 = ~n6171 & ~n6173;
  assign n6175 = pi031 & n6170;
  assign n6176 = n6174 & ~n6175;
  assign n6177 = ~pi106 & ~n6176;
  assign n6178 = pi100 & ~pi128;
  assign n6179 = pi037 & n6178;
  assign n6180 = pi106 & n6179;
  assign n6181 = pi031 & n6178;
  assign n6182 = pi035 & n6181;
  assign n6183 = ~n6180 & ~n6182;
  assign n6184 = ~pi035 & pi106;
  assign n6185 = ~pi037 & pi128;
  assign n6186 = pi031 & n6185;
  assign n6187 = n6184 & n6186;
  assign n6188 = n6183 & ~n6187;
  assign n6189 = ~n6177 & n6188;
  assign n6190 = pi065 & ~n6189;
  assign n6191 = ~pi100 & ~pi128;
  assign n6192 = pi037 & n6191;
  assign n6193 = ~pi031 & n6192;
  assign n6194 = ~pi035 & n6193;
  assign n6195 = ~pi031 & n6191;
  assign n6196 = pi035 & n6195;
  assign n6197 = ~pi037 & n6191;
  assign n6198 = pi106 & n6197;
  assign n6199 = ~n6196 & ~n6198;
  assign n6200 = ~pi035 & n6179;
  assign n6201 = ~pi106 & n6200;
  assign n6202 = pi037 & pi100;
  assign n6203 = pi031 & n6202;
  assign n6204 = pi106 & n6203;
  assign n6205 = ~n6201 & ~n6204;
  assign n6206 = n6199 & n6205;
  assign n6207 = ~pi065 & ~n6206;
  assign n6208 = ~n6194 & ~n6207;
  assign n6209 = ~pi037 & pi100;
  assign n6210 = ~pi031 & n6209;
  assign n6211 = ~pi035 & n6210;
  assign n6212 = pi031 & n6197;
  assign n6213 = pi035 & n6212;
  assign n6214 = ~n6211 & ~n6213;
  assign n6215 = pi106 & ~n6214;
  assign n6216 = n6208 & ~n6215;
  assign n6217 = ~n6190 & n6216;
  assign n6218 = ~n6168 & n6217;
  assign n6219 = ~pi068 & ~n6218;
  assign n6220 = pi031 & n6166;
  assign n6221 = pi035 & n6220;
  assign n6222 = pi035 & n6173;
  assign n6223 = ~n6221 & ~n6222;
  assign n6224 = ~n6185 & ~n6209;
  assign n6225 = pi035 & ~n6224;
  assign n6226 = pi037 & n6165;
  assign n6227 = ~pi035 & n6226;
  assign n6228 = ~pi031 & n6227;
  assign n6229 = ~n6225 & ~n6228;
  assign n6230 = ~pi031 & ~pi037;
  assign n6231 = ~pi035 & n6230;
  assign n6232 = n6191 & n6231;
  assign n6233 = n6229 & ~n6232;
  assign n6234 = ~pi106 & ~n6233;
  assign n6235 = ~pi035 & n6181;
  assign n6236 = pi106 & n6235;
  assign n6237 = pi035 & n6192;
  assign n6238 = pi106 & n6237;
  assign n6239 = ~n6236 & ~n6238;
  assign n6240 = ~n6234 & n6239;
  assign n6241 = n6223 & n6240;
  assign n6242 = pi065 & ~n6241;
  assign n6243 = ~n6219 & ~n6242;
  assign n6244 = pi037 & pi128;
  assign n6245 = pi035 & n6244;
  assign n6246 = pi031 & pi035;
  assign n6247 = ~pi106 & n6246;
  assign n6248 = n6191 & n6247;
  assign n6249 = pi106 & n6175;
  assign n6250 = ~pi031 & n6165;
  assign n6251 = pi035 & n6250;
  assign n6252 = ~pi031 & n6244;
  assign n6253 = ~pi106 & n6252;
  assign n6254 = ~n6251 & ~n6253;
  assign n6255 = ~n6249 & n6254;
  assign n6256 = ~n6248 & n6255;
  assign n6257 = ~n6245 & n6256;
  assign n6258 = ~pi065 & ~n6257;
  assign n6259 = ~pi031 & n6169;
  assign n6260 = pi106 & n6259;
  assign n6261 = ~pi035 & n6212;
  assign n6262 = ~pi031 & n6178;
  assign n6263 = pi031 & n6172;
  assign n6264 = ~n6262 & ~n6263;
  assign n6265 = ~pi106 & ~n6264;
  assign n6266 = ~n6261 & ~n6265;
  assign n6267 = ~n6260 & n6266;
  assign n6268 = ~pi031 & pi035;
  assign n6269 = n6192 & n6268;
  assign n6270 = n6267 & ~n6269;
  assign n6271 = pi065 & ~n6270;
  assign n6272 = ~pi035 & ~pi128;
  assign n6273 = pi031 & n6272;
  assign n6274 = ~pi031 & n6226;
  assign n6275 = ~n6273 & ~n6274;
  assign n6276 = pi106 & ~n6275;
  assign n6277 = pi035 & ~pi100;
  assign n6278 = ~pi031 & n6277;
  assign n6279 = pi035 & n6172;
  assign n6280 = ~n6278 & ~n6279;
  assign n6281 = pi106 & ~n6280;
  assign n6282 = ~n6276 & ~n6281;
  assign n6283 = pi035 & n6262;
  assign n6284 = pi035 & n6166;
  assign n6285 = ~n6232 & ~n6284;
  assign n6286 = ~n6283 & n6285;
  assign n6287 = ~pi106 & ~n6286;
  assign n6288 = n6282 & ~n6287;
  assign n6289 = ~n6271 & n6288;
  assign n6290 = ~n6258 & n6289;
  assign n6291 = pi068 & ~n6290;
  assign n6292 = n6243 & ~n6291;
  assign n6293 = pi037 & ~pi100;
  assign n6294 = ~pi031 & n6293;
  assign n6295 = pi035 & n6294;
  assign n6296 = ~pi031 & ~pi035;
  assign n6297 = ~pi037 & n6296;
  assign n6298 = n6169 & n6297;
  assign n6299 = ~n6295 & ~n6298;
  assign n6300 = ~pi035 & n6192;
  assign n6301 = pi035 & n6179;
  assign n6302 = pi035 & n6263;
  assign n6303 = ~n6301 & ~n6302;
  assign n6304 = ~n6300 & n6303;
  assign n6305 = n6299 & n6304;
  assign n6306 = pi106 & ~n6305;
  assign n6307 = pi031 & n6179;
  assign n6308 = pi035 & n6307;
  assign n6309 = ~n6194 & ~n6308;
  assign n6310 = pi035 & n6274;
  assign n6311 = ~pi035 & n6166;
  assign n6312 = pi031 & n6209;
  assign n6313 = ~pi035 & n6312;
  assign n6314 = ~n6311 & ~n6313;
  assign n6315 = ~n6310 & n6314;
  assign n6316 = ~pi106 & ~n6315;
  assign n6317 = n6309 & ~n6316;
  assign n6318 = ~n6306 & n6317;
  assign n6319 = ~pi065 & ~n6318;
  assign n6320 = pi035 & pi106;
  assign n6321 = n6203 & n6320;
  assign n6322 = ~pi037 & n6178;
  assign n6323 = ~pi031 & n6322;
  assign n6324 = pi035 & n6323;
  assign n6325 = ~pi106 & n6324;
  assign n6326 = ~n6321 & ~n6325;
  assign n6327 = ~n6319 & n6326;
  assign n6328 = n6292 & n6327;
  assign n6329 = ~n6163 & n6328;
  assign n6330 = n6163 & ~n6328;
  assign n6331 = ~n6329 & ~n6330;
  assign n6332 = ~n6063 & ~n6331;
  assign n6333 = n6063 & n6331;
  assign n6334 = ~n6332 & ~n6333;
  assign n6335 = ~n5901 & n6334;
  assign n6336 = n5901 & ~n6334;
  assign n6337 = ~n6335 & ~n6336;
  assign n6338 = ~pi529 & n6337;
  assign po134 = n5316 | n6338;
  assign n6340 = ~pi138 & pi517;
  assign n6341 = pi138 & ~pi517;
  assign n6342 = ~n6340 & ~n6341;
  assign n6343 = pi529 & ~n6342;
  assign n6344 = pi076 & n5381;
  assign n6345 = n5345 & n6344;
  assign n6346 = pi043 & n5330;
  assign n6347 = ~n5383 & ~n6346;
  assign n6348 = pi043 & n5363;
  assign n6349 = n6347 & ~n6348;
  assign n6350 = ~pi122 & ~n6349;
  assign n6351 = ~n5360 & ~n6350;
  assign n6352 = ~n5452 & ~n6154;
  assign n6353 = pi122 & ~n6352;
  assign n6354 = n6351 & ~n6353;
  assign n6355 = pi039 & ~n6354;
  assign n6356 = ~pi122 & n6140;
  assign n6357 = ~n5486 & ~n6356;
  assign n6358 = n5327 & n5538;
  assign n6359 = ~n5337 & ~n6358;
  assign n6360 = ~pi039 & ~n6359;
  assign n6361 = n6357 & ~n6360;
  assign n6362 = ~n6355 & n6361;
  assign n6363 = ~n6345 & n6362;
  assign n6364 = ~pi017 & ~n6363;
  assign n6365 = pi122 & n5475;
  assign n6366 = pi039 & pi043;
  assign n6367 = n6365 & n6366;
  assign n6368 = ~n5338 & ~n5391;
  assign n6369 = n5318 & ~n6368;
  assign n6370 = pi122 & n6369;
  assign n6371 = ~n5588 & ~n6370;
  assign n6372 = ~pi043 & n5398;
  assign n6373 = ~n5346 & ~n6372;
  assign n6374 = n5456 & ~n6373;
  assign n6375 = n6371 & ~n6374;
  assign n6376 = ~pi122 & n5558;
  assign n6377 = n5438 & n5445;
  assign n6378 = ~n5464 & ~n6377;
  assign n6379 = ~pi122 & ~n6378;
  assign n6380 = ~n6376 & ~n6379;
  assign n6381 = ~n5507 & n6380;
  assign n6382 = pi039 & ~n6381;
  assign n6383 = n6375 & ~n6382;
  assign n6384 = ~n6367 & n6383;
  assign n6385 = pi122 & n5420;
  assign n6386 = ~pi122 & n5513;
  assign n6387 = ~n6143 & ~n6386;
  assign n6388 = ~n5510 & n6387;
  assign n6389 = ~n6385 & n6388;
  assign n6390 = ~pi122 & n5346;
  assign n6391 = ~n5329 & ~n6071;
  assign n6392 = ~n5592 & n6391;
  assign n6393 = ~n6390 & n6392;
  assign n6394 = n6389 & n6393;
  assign n6395 = ~pi039 & ~n6394;
  assign n6396 = pi122 & n6100;
  assign n6397 = ~n6069 & ~n6396;
  assign n6398 = ~n6395 & n6397;
  assign n6399 = pi122 & n5512;
  assign n6400 = pi077 & n5438;
  assign n6401 = ~n5413 & ~n6400;
  assign n6402 = ~pi122 & ~n6401;
  assign n6403 = ~n6399 & ~n6402;
  assign n6404 = ~pi122 & n5492;
  assign n6405 = n6403 & ~n6404;
  assign n6406 = pi039 & ~n6405;
  assign n6407 = pi076 & n5368;
  assign n6408 = ~n5392 & ~n6407;
  assign n6409 = ~n5331 & n6408;
  assign n6410 = n5381 & ~n6409;
  assign n6411 = ~n6083 & ~n6410;
  assign n6412 = ~n6406 & n6411;
  assign n6413 = n6398 & n6412;
  assign n6414 = pi017 & ~n6413;
  assign n6415 = pi043 & n5413;
  assign n6416 = pi043 & n5412;
  assign n6417 = ~n6077 & ~n6416;
  assign n6418 = ~n5337 & n6417;
  assign n6419 = pi122 & ~n6418;
  assign n6420 = ~n5377 & ~n5467;
  assign n6421 = ~n5527 & n6420;
  assign n6422 = ~pi122 & ~n6421;
  assign n6423 = n5391 & n5444;
  assign n6424 = ~n6422 & ~n6423;
  assign n6425 = ~n6419 & n6424;
  assign n6426 = ~n6415 & n6425;
  assign n6427 = ~n5586 & n6426;
  assign n6428 = ~pi039 & ~n6427;
  assign n6429 = ~n6414 & ~n6428;
  assign n6430 = n6384 & n6429;
  assign n6431 = ~n6364 & n6430;
  assign n6432 = n5484 & n6431;
  assign n6433 = ~n5484 & ~n6431;
  assign n6434 = ~n6432 & ~n6433;
  assign n6435 = ~pi091 & n5856;
  assign n6436 = n5653 & n5719;
  assign n6437 = ~n5752 & ~n6436;
  assign n6438 = ~pi091 & ~n6437;
  assign n6439 = ~n6435 & ~n6438;
  assign n6440 = ~n5798 & n6439;
  assign n6441 = pi024 & ~n6440;
  assign n6442 = n5607 & n5761;
  assign n6443 = pi024 & n6442;
  assign n6444 = ~n6441 & ~n6443;
  assign n6445 = ~n5636 & ~n5643;
  assign n6446 = n5730 & ~n6445;
  assign n6447 = pi091 & n6446;
  assign n6448 = ~n5868 & ~n6447;
  assign n6449 = ~pi005 & n5628;
  assign n6450 = ~n5651 & ~n6449;
  assign n6451 = n5697 & ~n6450;
  assign n6452 = n6448 & ~n6451;
  assign n6453 = n6444 & n6452;
  assign n6454 = pi005 & n5676;
  assign n6455 = ~n5623 & ~n5754;
  assign n6456 = ~n5819 & n6455;
  assign n6457 = ~pi091 & ~n6456;
  assign n6458 = pi005 & n5762;
  assign n6459 = pi005 & n5608;
  assign n6460 = ~n6458 & ~n6459;
  assign n6461 = ~n5746 & n6460;
  assign n6462 = pi091 & ~n6461;
  assign n6463 = ~pi005 & n5636;
  assign n6464 = ~pi091 & n6463;
  assign n6465 = ~n6462 & ~n6464;
  assign n6466 = ~n6457 & n6465;
  assign n6467 = ~n6454 & n6466;
  assign n6468 = ~n5866 & n6467;
  assign n6469 = ~pi024 & ~n6468;
  assign n6470 = n5706 & n5730;
  assign n6471 = n5636 & n5730;
  assign n6472 = ~n6470 & ~n6471;
  assign n6473 = n5621 & n5663;
  assign n6474 = ~n5616 & ~n5637;
  assign n6475 = pi004 & n5659;
  assign n6476 = n6474 & ~n6475;
  assign n6477 = n5607 & ~n6476;
  assign n6478 = ~n6473 & ~n6477;
  assign n6479 = ~pi091 & n5811;
  assign n6480 = n5621 & n6479;
  assign n6481 = ~pi005 & pi052;
  assign n6482 = pi004 & n6481;
  assign n6483 = ~n5676 & ~n6482;
  assign n6484 = ~pi091 & ~n6483;
  assign n6485 = ~pi004 & n5635;
  assign n6486 = pi091 & n6485;
  assign n6487 = ~n6484 & ~n6486;
  assign n6488 = ~n6480 & n6487;
  assign n6489 = pi024 & ~n6488;
  assign n6490 = ~pi005 & n5620;
  assign n6491 = pi091 & n6490;
  assign n6492 = ~pi091 & n5806;
  assign n6493 = ~pi004 & n5653;
  assign n6494 = pi091 & n6493;
  assign n6495 = ~n6492 & ~n6494;
  assign n6496 = ~n5792 & n6495;
  assign n6497 = ~n6491 & n6496;
  assign n6498 = ~pi091 & n5651;
  assign n6499 = ~n5614 & ~n6463;
  assign n6500 = ~n5864 & n6499;
  assign n6501 = ~n6498 & n6500;
  assign n6502 = n6497 & n6501;
  assign n6503 = ~pi024 & ~n6502;
  assign n6504 = ~n6489 & ~n6503;
  assign n6505 = n6478 & n6504;
  assign n6506 = n6472 & n6505;
  assign n6507 = pi018 & ~n6506;
  assign n6508 = pi004 & n5607;
  assign n6509 = n5650 & n6508;
  assign n6510 = pi005 & n5615;
  assign n6511 = ~n5831 & ~n6510;
  assign n6512 = pi005 & n5664;
  assign n6513 = n6511 & ~n6512;
  assign n6514 = ~pi091 & ~n6513;
  assign n6515 = ~n5655 & ~n6514;
  assign n6516 = pi005 & n5872;
  assign n6517 = ~n5698 & ~n6516;
  assign n6518 = pi091 & ~n6517;
  assign n6519 = n6515 & ~n6518;
  assign n6520 = pi024 & ~n6519;
  assign n6521 = pi005 & n5754;
  assign n6522 = ~pi091 & n6521;
  assign n6523 = ~n5773 & ~n6522;
  assign n6524 = n5612 & n5836;
  assign n6525 = ~n5746 & ~n6524;
  assign n6526 = ~pi024 & ~n6525;
  assign n6527 = n6523 & ~n6526;
  assign n6528 = ~n6520 & n6527;
  assign n6529 = ~n6509 & n6528;
  assign n6530 = ~pi018 & ~n6529;
  assign n6531 = ~n6507 & ~n6530;
  assign n6532 = ~n6469 & n6531;
  assign n6533 = n6453 & n6532;
  assign n6534 = ~n5772 & n6533;
  assign n6535 = n5772 & ~n6533;
  assign n6536 = ~n6534 & ~n6535;
  assign n6537 = n6434 & n6536;
  assign n6538 = ~n6434 & ~n6536;
  assign n6539 = ~n6537 & ~n6538;
  assign n6540 = pi031 & n6322;
  assign n6541 = pi035 & n6540;
  assign n6542 = pi106 & n6302;
  assign n6543 = ~pi031 & n6166;
  assign n6544 = n6320 & n6543;
  assign n6545 = ~n6542 & ~n6544;
  assign n6546 = ~n6541 & n6545;
  assign n6547 = n6184 & n6323;
  assign n6548 = pi106 & n6261;
  assign n6549 = ~n6547 & ~n6548;
  assign n6550 = ~pi065 & ~n6549;
  assign n6551 = n6546 & ~n6550;
  assign n6552 = ~pi031 & n6179;
  assign n6553 = pi035 & n6552;
  assign n6554 = ~pi031 & n6185;
  assign n6555 = ~pi035 & n6554;
  assign n6556 = ~pi035 & n6175;
  assign n6557 = pi035 & n6226;
  assign n6558 = ~n6556 & ~n6557;
  assign n6559 = ~n6555 & n6558;
  assign n6560 = ~pi106 & ~n6559;
  assign n6561 = pi106 & n6279;
  assign n6562 = pi035 & n6322;
  assign n6563 = ~n6311 & ~n6562;
  assign n6564 = ~pi106 & ~n6563;
  assign n6565 = n6202 & n6296;
  assign n6566 = ~pi035 & n6195;
  assign n6567 = ~n6565 & ~n6566;
  assign n6568 = ~n6564 & n6567;
  assign n6569 = ~n6561 & n6568;
  assign n6570 = pi037 & ~pi128;
  assign n6571 = ~pi031 & n6570;
  assign n6572 = pi106 & n6571;
  assign n6573 = ~n6180 & ~n6572;
  assign n6574 = ~n6302 & n6573;
  assign n6575 = n6569 & n6574;
  assign n6576 = ~pi065 & ~n6575;
  assign n6577 = ~pi106 & n6197;
  assign n6578 = ~pi035 & n6178;
  assign n6579 = ~pi106 & n6578;
  assign n6580 = ~pi035 & n6293;
  assign n6581 = ~n6186 & ~n6580;
  assign n6582 = ~n6170 & n6581;
  assign n6583 = pi106 & ~n6582;
  assign n6584 = pi031 & n6244;
  assign n6585 = ~pi035 & n6584;
  assign n6586 = ~n6583 & ~n6585;
  assign n6587 = ~n6579 & n6586;
  assign n6588 = ~n6577 & n6587;
  assign n6589 = ~n6175 & ~n6284;
  assign n6590 = n6588 & n6589;
  assign n6591 = pi065 & ~n6590;
  assign n6592 = ~n6576 & ~n6591;
  assign n6593 = ~n6560 & n6592;
  assign n6594 = ~n6553 & n6593;
  assign n6595 = ~n6172 & ~n6322;
  assign n6596 = pi031 & ~n6595;
  assign n6597 = pi035 & n6169;
  assign n6598 = pi031 & n6597;
  assign n6599 = ~n6596 & ~n6598;
  assign n6600 = pi106 & ~n6599;
  assign n6601 = n6594 & ~n6600;
  assign n6602 = pi068 & ~n6601;
  assign n6603 = ~pi031 & n6170;
  assign n6604 = ~pi106 & n6603;
  assign n6605 = pi031 & n6226;
  assign n6606 = pi035 & n6605;
  assign n6607 = ~n6279 & ~n6606;
  assign n6608 = ~pi035 & n6307;
  assign n6609 = ~pi037 & ~pi128;
  assign n6610 = ~pi031 & n6609;
  assign n6611 = ~n6608 & ~n6610;
  assign n6612 = pi106 & ~n6611;
  assign n6613 = ~n6228 & ~n6612;
  assign n6614 = n6607 & n6613;
  assign n6615 = ~n6604 & n6614;
  assign n6616 = pi065 & ~n6615;
  assign n6617 = pi035 & ~pi106;
  assign n6618 = n6175 & n6617;
  assign n6619 = ~n6212 & ~n6555;
  assign n6620 = ~n6165 & ~n6244;
  assign n6621 = n6184 & ~n6620;
  assign n6622 = pi031 & pi106;
  assign n6623 = n6191 & n6622;
  assign n6624 = ~n6621 & ~n6623;
  assign n6625 = n6619 & n6624;
  assign n6626 = ~n6618 & n6625;
  assign n6627 = ~pi065 & ~n6626;
  assign n6628 = ~n6616 & ~n6627;
  assign n6629 = ~pi035 & n6323;
  assign n6630 = ~pi035 & n6605;
  assign n6631 = ~n6182 & ~n6630;
  assign n6632 = ~pi106 & ~n6631;
  assign n6633 = pi106 & n6274;
  assign n6634 = n6320 & n6610;
  assign n6635 = ~n6633 & ~n6634;
  assign n6636 = ~n6632 & n6635;
  assign n6637 = ~n6629 & n6636;
  assign n6638 = n6628 & n6637;
  assign n6639 = ~pi068 & ~n6638;
  assign n6640 = n6202 & n6268;
  assign n6641 = ~n6284 & ~n6640;
  assign n6642 = pi106 & ~n6641;
  assign n6643 = n6173 & n6617;
  assign n6644 = ~n6249 & ~n6643;
  assign n6645 = ~pi035 & ~pi106;
  assign n6646 = ~n6262 & ~n6603;
  assign n6647 = ~pi037 & ~pi100;
  assign n6648 = pi031 & n6647;
  assign n6649 = n6646 & ~n6648;
  assign n6650 = n6645 & ~n6649;
  assign n6651 = n6644 & ~n6650;
  assign n6652 = ~n6642 & n6651;
  assign n6653 = pi065 & ~n6652;
  assign n6654 = ~pi065 & ~pi106;
  assign n6655 = n6251 & n6654;
  assign n6656 = ~n6653 & ~n6655;
  assign n6657 = ~n6639 & n6656;
  assign n6658 = ~n6602 & n6657;
  assign n6659 = n6551 & n6658;
  assign n6660 = ~n5603 & n6659;
  assign n6661 = n5603 & ~n6659;
  assign n6662 = ~n6660 & ~n6661;
  assign n6663 = ~pi125 & n5907;
  assign n6664 = ~pi009 & n6663;
  assign n6665 = pi009 & n5911;
  assign n6666 = ~pi009 & n5951;
  assign n6667 = ~n6665 & ~n6666;
  assign n6668 = ~n6664 & n6667;
  assign n6669 = ~pi113 & ~n6668;
  assign n6670 = ~pi125 & n5936;
  assign n6671 = ~pi124 & n6670;
  assign n6672 = pi009 & n6671;
  assign n6673 = pi009 & n5928;
  assign n6674 = pi125 & n6673;
  assign n6675 = ~n5929 & ~n5940;
  assign n6676 = pi125 & ~n6675;
  assign n6677 = ~n6674 & ~n6676;
  assign n6678 = pi113 & ~n6677;
  assign n6679 = ~n6672 & ~n6678;
  assign n6680 = n5929 & n5978;
  assign n6681 = pi025 & ~pi124;
  assign n6682 = ~pi125 & n6681;
  assign n6683 = pi113 & n6682;
  assign n6684 = pi113 & n5991;
  assign n6685 = pi009 & ~pi113;
  assign n6686 = n5940 & n6685;
  assign n6687 = ~n5955 & ~n6686;
  assign n6688 = ~n6684 & n6687;
  assign n6689 = ~n6683 & n6688;
  assign n6690 = ~n6680 & n6689;
  assign n6691 = ~pi009 & n5969;
  assign n6692 = n5917 & n5936;
  assign n6693 = ~n6691 & ~n6692;
  assign n6694 = n5924 & n5966;
  assign n6695 = n6693 & ~n6694;
  assign n6696 = n6690 & n6695;
  assign n6697 = ~pi096 & ~n6696;
  assign n6698 = ~pi009 & n6038;
  assign n6699 = ~n5948 & ~n6698;
  assign n6700 = ~n5959 & n6699;
  assign n6701 = pi113 & ~n6700;
  assign n6702 = ~pi113 & n5916;
  assign n6703 = ~n5951 & ~n6027;
  assign n6704 = ~n6702 & n6703;
  assign n6705 = ~n6701 & n6704;
  assign n6706 = ~pi009 & n5902;
  assign n6707 = ~pi113 & n6706;
  assign n6708 = pi125 & n6012;
  assign n6709 = ~pi009 & n6708;
  assign n6710 = ~n6707 & ~n6709;
  assign n6711 = n6705 & n6710;
  assign n6712 = pi096 & ~n6711;
  assign n6713 = ~n6697 & ~n6712;
  assign n6714 = n6679 & n6713;
  assign n6715 = ~n6669 & n6714;
  assign n6716 = ~pi010 & ~n6715;
  assign n6717 = ~pi025 & ~pi124;
  assign n6718 = ~pi125 & n6717;
  assign n6719 = n5938 & n6718;
  assign n6720 = pi113 & n5912;
  assign n6721 = ~n6719 & ~n6720;
  assign n6722 = pi125 & n5911;
  assign n6723 = ~pi009 & n6722;
  assign n6724 = ~n5956 & ~n6723;
  assign n6725 = ~pi113 & ~n6724;
  assign n6726 = ~pi009 & n5941;
  assign n6727 = ~n6725 & ~n6726;
  assign n6728 = n6721 & n6727;
  assign n6729 = ~n5913 & ~n5991;
  assign n6730 = ~pi125 & n5948;
  assign n6731 = ~pi113 & n6730;
  assign n6732 = pi009 & n6722;
  assign n6733 = pi096 & ~n6732;
  assign n6734 = ~pi009 & n6046;
  assign n6735 = ~n6718 & ~n6734;
  assign n6736 = pi113 & ~n6735;
  assign n6737 = n6733 & ~n6736;
  assign n6738 = ~n6731 & n6737;
  assign n6739 = n6729 & n6738;
  assign n6740 = n5951 & n6685;
  assign n6741 = ~pi096 & ~n6740;
  assign n6742 = ~n5999 & ~n6664;
  assign n6743 = pi125 & n5915;
  assign n6744 = pi113 & n6743;
  assign n6745 = ~n5910 & ~n6012;
  assign n6746 = n5958 & ~n6745;
  assign n6747 = ~n6744 & ~n6746;
  assign n6748 = n6742 & n6747;
  assign n6749 = n6741 & n6748;
  assign n6750 = ~n6739 & ~n6749;
  assign n6751 = n6728 & ~n6750;
  assign n6752 = pi010 & ~n6751;
  assign n6753 = n5936 & n5989;
  assign n6754 = ~n6027 & ~n6753;
  assign n6755 = pi113 & ~n6754;
  assign n6756 = ~pi025 & ~pi055;
  assign n6757 = pi125 & n6756;
  assign n6758 = ~n6003 & ~n6730;
  assign n6759 = ~n6757 & n6758;
  assign n6760 = n5966 & ~n6759;
  assign n6761 = ~n6755 & ~n6760;
  assign n6762 = ~pi113 & n5931;
  assign n6763 = n6761 & ~n6762;
  assign n6764 = ~n6023 & n6763;
  assign n6765 = pi096 & ~n6764;
  assign n6766 = ~pi125 & n5924;
  assign n6767 = n5938 & n6766;
  assign n6768 = pi113 & n6680;
  assign n6769 = ~n6767 & ~n6768;
  assign n6770 = pi125 & n5940;
  assign n6771 = pi009 & n6770;
  assign n6772 = n6769 & ~n6771;
  assign n6773 = ~pi096 & ~pi113;
  assign n6774 = n6016 & n6773;
  assign n6775 = n6772 & ~n6774;
  assign n6776 = ~n6765 & n6775;
  assign n6777 = pi113 & n6000;
  assign n6778 = n5941 & n5958;
  assign n6779 = ~n6777 & ~n6778;
  assign n6780 = ~pi096 & ~n6779;
  assign n6781 = n6776 & ~n6780;
  assign n6782 = ~n6752 & n6781;
  assign n6783 = ~n6716 & n6782;
  assign n6784 = ~pi138 & ~n6783;
  assign n6785 = pi138 & n6783;
  assign n6786 = ~n6784 & ~n6785;
  assign n6787 = n6662 & n6786;
  assign n6788 = ~n6662 & ~n6786;
  assign n6789 = ~n6787 & ~n6788;
  assign n6790 = ~n6539 & n6789;
  assign n6791 = n6539 & ~n6789;
  assign n6792 = ~n6790 & ~n6791;
  assign n6793 = ~pi529 & n6792;
  assign po135 = n6343 | n6793;
  assign n6795 = pi191 & pi405;
  assign n6796 = ~pi191 & ~pi405;
  assign n6797 = ~n6795 & ~n6796;
  assign n6798 = pi529 & n6797;
  assign n6799 = n5938 & n5959;
  assign n6800 = ~n5971 & ~n6799;
  assign n6801 = ~pi096 & ~n6800;
  assign n6802 = ~pi009 & n6682;
  assign n6803 = ~pi009 & n5911;
  assign n6804 = ~n6802 & ~n6803;
  assign n6805 = ~pi113 & ~n6804;
  assign n6806 = ~n5999 & ~n6047;
  assign n6807 = ~pi113 & ~n6806;
  assign n6808 = ~n6805 & ~n6807;
  assign n6809 = ~pi113 & ~pi125;
  assign n6810 = pi124 & n6809;
  assign n6811 = pi009 & n6013;
  assign n6812 = ~n6810 & ~n6811;
  assign n6813 = ~pi096 & ~n6812;
  assign n6814 = pi125 & n5921;
  assign n6815 = ~n6722 & ~n6814;
  assign n6816 = n5938 & ~n6815;
  assign n6817 = ~pi125 & n5938;
  assign n6818 = ~pi025 & n6817;
  assign n6819 = n5915 & n6818;
  assign n6820 = ~n6816 & ~n6819;
  assign n6821 = ~n6813 & n6820;
  assign n6822 = n6808 & n6821;
  assign n6823 = ~n6801 & n6822;
  assign n6824 = n5958 & n6049;
  assign n6825 = pi009 & n5948;
  assign n6826 = ~pi055 & n5978;
  assign n6827 = pi009 & n5940;
  assign n6828 = ~n6826 & ~n6827;
  assign n6829 = ~pi113 & ~n6828;
  assign n6830 = ~pi009 & n5925;
  assign n6831 = ~n6829 & ~n6830;
  assign n6832 = ~n6825 & n6831;
  assign n6833 = ~n6824 & n6832;
  assign n6834 = pi096 & ~n6833;
  assign n6835 = n6823 & ~n6834;
  assign n6836 = pi010 & ~n6835;
  assign n6837 = ~n6041 & ~n6766;
  assign n6838 = ~n5964 & ~n6004;
  assign n6839 = ~n6015 & n6838;
  assign n6840 = ~pi009 & ~n6839;
  assign n6841 = n6837 & ~n6840;
  assign n6842 = pi096 & pi113;
  assign n6843 = ~n6841 & n6842;
  assign n6844 = n5917 & n5954;
  assign n6845 = ~n5979 & ~n6844;
  assign n6846 = ~pi113 & ~n6845;
  assign n6847 = ~n6843 & ~n6846;
  assign n6848 = pi009 & n5916;
  assign n6849 = ~pi009 & n5937;
  assign n6850 = ~n5926 & ~n6849;
  assign n6851 = ~n6848 & n6850;
  assign n6852 = ~pi096 & pi113;
  assign n6853 = ~n6851 & n6852;
  assign n6854 = pi096 & ~pi113;
  assign n6855 = pi125 & n6038;
  assign n6856 = ~n5912 & ~n5941;
  assign n6857 = ~n6855 & n6856;
  assign n6858 = pi009 & ~n6857;
  assign n6859 = ~n5922 & ~n6858;
  assign n6860 = n6854 & ~n6859;
  assign n6861 = pi009 & n6663;
  assign n6862 = ~pi113 & n6861;
  assign n6863 = ~n6805 & ~n6862;
  assign n6864 = ~n6709 & n6863;
  assign n6865 = ~pi096 & ~n6864;
  assign n6866 = ~n6860 & ~n6865;
  assign n6867 = ~n6853 & n6866;
  assign n6868 = n6847 & n6867;
  assign n6869 = ~pi009 & n6015;
  assign n6870 = ~pi009 & n6855;
  assign n6871 = ~n6869 & ~n6870;
  assign n6872 = ~n6046 & n6871;
  assign n6873 = pi113 & ~n6872;
  assign n6874 = n5938 & n5980;
  assign n6875 = n5994 & n6681;
  assign n6876 = ~n6874 & ~n6875;
  assign n6877 = ~n6873 & n6876;
  assign n6878 = ~n5937 & ~n6757;
  assign n6879 = ~n5903 & n6878;
  assign n6880 = ~pi113 & ~n6879;
  assign n6881 = ~pi113 & n5954;
  assign n6882 = n5958 & n6663;
  assign n6883 = ~n6707 & ~n6882;
  assign n6884 = ~n6881 & n6883;
  assign n6885 = ~n6880 & n6884;
  assign n6886 = ~n5904 & ~n6040;
  assign n6887 = n6885 & n6886;
  assign n6888 = ~pi096 & ~n6887;
  assign n6889 = n6877 & ~n6888;
  assign n6890 = n5929 & n5966;
  assign n6891 = ~n5926 & ~n6890;
  assign n6892 = pi096 & ~n6891;
  assign n6893 = ~pi113 & n5904;
  assign n6894 = ~pi009 & n5915;
  assign n6895 = ~n6757 & ~n6894;
  assign n6896 = pi009 & n5902;
  assign n6897 = pi055 & ~pi125;
  assign n6898 = ~n6896 & ~n6897;
  assign n6899 = n6895 & n6898;
  assign n6900 = n6842 & ~n6899;
  assign n6901 = ~n6893 & ~n6900;
  assign n6902 = ~n6892 & n6901;
  assign n6903 = n6889 & n6902;
  assign n6904 = ~pi010 & ~n6903;
  assign n6905 = n6868 & ~n6904;
  assign n6906 = ~n6836 & n6905;
  assign n6907 = pi191 & n6906;
  assign n6908 = ~pi191 & ~n6906;
  assign n6909 = ~n6907 & ~n6908;
  assign n6910 = ~pi005 & ~n5763;
  assign n6911 = pi005 & n5839;
  assign n6912 = ~pi091 & n6911;
  assign n6913 = ~n6910 & ~n6912;
  assign n6914 = ~pi024 & ~n6913;
  assign n6915 = ~pi005 & n5630;
  assign n6916 = ~n5654 & ~n6915;
  assign n6917 = n5736 & ~n6916;
  assign n6918 = ~n6914 & ~n6917;
  assign n6919 = ~n5636 & ~n5664;
  assign n6920 = n5811 & ~n6919;
  assign n6921 = pi091 & n6920;
  assign n6922 = ~pi004 & n5608;
  assign n6923 = ~pi005 & n6922;
  assign n6924 = ~n5786 & ~n5788;
  assign n6925 = ~n6923 & n6924;
  assign n6926 = ~pi091 & ~n6925;
  assign n6927 = n5643 & n5705;
  assign n6928 = pi004 & n6510;
  assign n6929 = pi091 & n5751;
  assign n6930 = ~n6928 & ~n6929;
  assign n6931 = ~n6927 & n6930;
  assign n6932 = ~n5698 & ~n6485;
  assign n6933 = n6931 & n6932;
  assign n6934 = pi024 & ~n6933;
  assign n6935 = ~n6926 & ~n6934;
  assign n6936 = ~n6921 & n6935;
  assign n6937 = n6918 & n6936;
  assign n6938 = ~pi018 & ~n6937;
  assign n6939 = ~pi004 & ~pi094;
  assign n6940 = pi005 & n6939;
  assign n6941 = ~n6512 & ~n6940;
  assign n6942 = ~pi091 & ~n6941;
  assign n6943 = pi005 & n6493;
  assign n6944 = pi005 & ~pi084;
  assign n6945 = ~pi004 & n6944;
  assign n6946 = ~n5614 & ~n6945;
  assign n6947 = ~n6943 & n6946;
  assign n6948 = n5705 & n5756;
  assign n6949 = ~pi005 & n5609;
  assign n6950 = ~n5622 & ~n6949;
  assign n6951 = ~n5651 & n6950;
  assign n6952 = pi091 & ~n6951;
  assign n6953 = ~n6948 & ~n6952;
  assign n6954 = n6947 & n6953;
  assign n6955 = ~pi024 & ~n6954;
  assign n6956 = ~n6942 & ~n6955;
  assign n6957 = pi005 & n5637;
  assign n6958 = ~n5786 & ~n6957;
  assign n6959 = ~n5632 & n6958;
  assign n6960 = ~n5866 & n6959;
  assign n6961 = pi091 & ~n6960;
  assign n6962 = ~n5638 & ~n5720;
  assign n6963 = ~pi091 & ~n6962;
  assign n6964 = ~n6961 & ~n6963;
  assign n6965 = ~pi005 & n5621;
  assign n6966 = ~n5867 & ~n6965;
  assign n6967 = ~pi091 & n5677;
  assign n6968 = ~n6475 & ~n6967;
  assign n6969 = ~n5781 & n6968;
  assign n6970 = pi024 & ~n6969;
  assign n6971 = n6966 & ~n6970;
  assign n6972 = n6964 & n6971;
  assign n6973 = n6956 & n6972;
  assign n6974 = pi018 & ~n6973;
  assign n6975 = ~n6938 & ~n6974;
  assign n6976 = n5659 & n5719;
  assign n6977 = pi091 & n6976;
  assign n6978 = ~pi091 & n5746;
  assign n6979 = ~n6977 & ~n6978;
  assign n6980 = n5609 & n5730;
  assign n6981 = ~n6521 & ~n6980;
  assign n6982 = ~n5795 & n6981;
  assign n6983 = n6979 & n6982;
  assign n6984 = pi024 & ~n6983;
  assign n6985 = ~pi005 & n5659;
  assign n6986 = ~n6471 & ~n6985;
  assign n6987 = ~n5674 & n6986;
  assign n6988 = ~pi091 & ~n6987;
  assign n6989 = pi091 & n6957;
  assign n6990 = ~n5807 & ~n6470;
  assign n6991 = pi091 & ~n6990;
  assign n6992 = ~n6989 & ~n6991;
  assign n6993 = ~n6480 & n6992;
  assign n6994 = ~n6988 & n6993;
  assign n6995 = ~pi024 & ~n6994;
  assign n6996 = ~n6984 & ~n6995;
  assign n6997 = ~pi091 & n6928;
  assign n6998 = pi091 & n5732;
  assign n6999 = ~n6997 & ~n6998;
  assign n7000 = n6996 & n6999;
  assign n7001 = n6975 & n7000;
  assign n7002 = ~n5772 & n7001;
  assign n7003 = n5772 & ~n7001;
  assign n7004 = ~n7002 & ~n7003;
  assign n7005 = ~pi031 & n6647;
  assign n7006 = ~pi035 & n7005;
  assign n7007 = n6558 & ~n7006;
  assign n7008 = ~pi106 & ~n7007;
  assign n7009 = ~pi065 & pi106;
  assign n7010 = ~pi035 & n6244;
  assign n7011 = ~n6170 & ~n7010;
  assign n7012 = n7009 & ~n7011;
  assign n7013 = ~n6274 & ~n6323;
  assign n7014 = ~pi035 & ~n7013;
  assign n7015 = ~n6248 & ~n7014;
  assign n7016 = ~pi065 & ~n7015;
  assign n7017 = ~n7012 & ~n7016;
  assign n7018 = ~n7008 & n7017;
  assign n7019 = n6185 & n6645;
  assign n7020 = ~pi035 & n6191;
  assign n7021 = pi106 & n6301;
  assign n7022 = ~n7020 & ~n7021;
  assign n7023 = ~n7019 & n7022;
  assign n7024 = pi035 & n6165;
  assign n7025 = pi031 & n7024;
  assign n7026 = ~n6195 & ~n7025;
  assign n7027 = n7023 & n7026;
  assign n7028 = pi065 & ~n7027;
  assign n7029 = ~n6192 & ~n6209;
  assign n7030 = ~pi031 & ~n7029;
  assign n7031 = n6320 & n7030;
  assign n7032 = ~n7028 & ~n7031;
  assign n7033 = n7018 & n7032;
  assign n7034 = ~pi068 & ~n7033;
  assign n7035 = n6164 & n6570;
  assign n7036 = ~n6605 & ~n7035;
  assign n7037 = ~pi106 & ~n7036;
  assign n7038 = ~n6173 & ~n6556;
  assign n7039 = pi031 & n6192;
  assign n7040 = pi035 & n7039;
  assign n7041 = pi035 & n6252;
  assign n7042 = ~n7040 & ~n7041;
  assign n7043 = n7038 & n7042;
  assign n7044 = pi106 & ~n7043;
  assign n7045 = ~n7037 & ~n7044;
  assign n7046 = ~n6200 & ~n6222;
  assign n7047 = n7045 & n7046;
  assign n7048 = ~pi128 & n6268;
  assign n7049 = pi035 & n6209;
  assign n7050 = ~n7048 & ~n7049;
  assign n7051 = ~pi106 & ~n7050;
  assign n7052 = ~pi037 & n6268;
  assign n7053 = pi035 & n6259;
  assign n7054 = ~n7052 & ~n7053;
  assign n7055 = ~pi035 & n6571;
  assign n7056 = n7054 & ~n7055;
  assign n7057 = n6263 & n6645;
  assign n7058 = ~pi035 & ~pi037;
  assign n7059 = ~pi100 & n7058;
  assign n7060 = ~pi128 & n7059;
  assign n7061 = ~n6307 & ~n7060;
  assign n7062 = ~n6220 & n7061;
  assign n7063 = pi106 & ~n7062;
  assign n7064 = ~n7057 & ~n7063;
  assign n7065 = n7056 & n7064;
  assign n7066 = ~pi065 & ~n7065;
  assign n7067 = ~n7051 & ~n7066;
  assign n7068 = ~pi106 & n6202;
  assign n7069 = ~n6577 & ~n7068;
  assign n7070 = ~n6540 & n7069;
  assign n7071 = pi065 & ~n7070;
  assign n7072 = n7067 & ~n7071;
  assign n7073 = n7047 & n7072;
  assign n7074 = pi068 & ~n7073;
  assign n7075 = ~pi035 & n6552;
  assign n7076 = pi106 & n7075;
  assign n7077 = ~pi106 & n7025;
  assign n7078 = ~n7076 & ~n7077;
  assign n7079 = n6164 & n6322;
  assign n7080 = pi106 & ~n7079;
  assign n7081 = ~pi106 & ~n6585;
  assign n7082 = ~n7080 & ~n7081;
  assign n7083 = ~n6232 & ~n7082;
  assign n7084 = ~n6561 & n7083;
  assign n7085 = ~n6269 & n7084;
  assign n7086 = pi065 & ~n7085;
  assign n7087 = n7078 & ~n7086;
  assign n7088 = ~pi106 & n6553;
  assign n7089 = ~pi035 & n6322;
  assign n7090 = ~n6235 & ~n7089;
  assign n7091 = ~n6194 & n7090;
  assign n7092 = ~pi106 & ~n7091;
  assign n7093 = ~n6298 & ~n6565;
  assign n7094 = pi106 & ~n7093;
  assign n7095 = ~n7092 & ~n7094;
  assign n7096 = ~n7088 & n7095;
  assign n7097 = n6320 & n7039;
  assign n7098 = n7096 & ~n7097;
  assign n7099 = ~pi065 & ~n7098;
  assign n7100 = n7087 & ~n7099;
  assign n7101 = ~n7074 & n7100;
  assign n7102 = ~n7034 & n7101;
  assign n7103 = pi122 & n5320;
  assign n7104 = n5330 & n5366;
  assign n7105 = ~pi122 & n7104;
  assign n7106 = ~n7103 & ~n7105;
  assign n7107 = ~pi043 & n5335;
  assign n7108 = ~n5359 & ~n7107;
  assign n7109 = n5354 & ~n7108;
  assign n7110 = ~n5474 & ~n5475;
  assign n7111 = ~pi043 & ~n7110;
  assign n7112 = ~n6132 & ~n7111;
  assign n7113 = ~pi039 & ~n7112;
  assign n7114 = n5338 & n5444;
  assign n7115 = pi122 & n5463;
  assign n7116 = ~n7104 & ~n7115;
  assign n7117 = ~n7114 & n7116;
  assign n7118 = ~n5452 & ~n5512;
  assign n7119 = n7117 & n7118;
  assign n7120 = pi039 & ~n7119;
  assign n7121 = ~n5363 & ~n5391;
  assign n7122 = n5596 & ~n7121;
  assign n7123 = pi122 & n7122;
  assign n7124 = ~n7120 & ~n7123;
  assign n7125 = ~n7113 & n7124;
  assign n7126 = ~n7109 & n7125;
  assign n7127 = ~pi076 & n5412;
  assign n7128 = ~pi043 & n7127;
  assign n7129 = ~n5487 & ~n7128;
  assign n7130 = ~n5485 & n7129;
  assign n7131 = ~pi122 & ~n7130;
  assign n7132 = n7126 & ~n7131;
  assign n7133 = ~pi017 & ~n7132;
  assign n7134 = ~n5587 & ~n6100;
  assign n7135 = pi043 & n5392;
  assign n7136 = ~n5401 & ~n7135;
  assign n7137 = ~n5487 & n7136;
  assign n7138 = ~n5586 & n7137;
  assign n7139 = pi122 & ~n7138;
  assign n7140 = ~n5393 & ~n5439;
  assign n7141 = ~pi122 & ~n7140;
  assign n7142 = ~n7139 & ~n7141;
  assign n7143 = ~pi076 & ~pi109;
  assign n7144 = pi043 & n7143;
  assign n7145 = ~n6348 & ~n7144;
  assign n7146 = ~pi122 & ~n7145;
  assign n7147 = pi043 & n6142;
  assign n7148 = pi043 & ~pi070;
  assign n7149 = ~pi076 & n7148;
  assign n7150 = ~n5329 & ~n7149;
  assign n7151 = ~n7147 & n7150;
  assign n7152 = n5444 & n5466;
  assign n7153 = ~pi043 & n5322;
  assign n7154 = ~n5376 & ~n7153;
  assign n7155 = ~n5346 & n7154;
  assign n7156 = pi122 & ~n7155;
  assign n7157 = ~n7152 & ~n7156;
  assign n7158 = n7151 & n7157;
  assign n7159 = ~pi039 & ~n7158;
  assign n7160 = ~n7146 & ~n7159;
  assign n7161 = ~pi122 & n5349;
  assign n7162 = ~n5494 & ~n7161;
  assign n7163 = ~n6407 & n7162;
  assign n7164 = pi039 & ~n7163;
  assign n7165 = n7160 & ~n7164;
  assign n7166 = n7142 & n7165;
  assign n7167 = n7134 & n7166;
  assign n7168 = pi017 & ~n7167;
  assign n7169 = ~n6116 & ~n6140;
  assign n7170 = pi122 & n5438;
  assign n7171 = n5368 & n7170;
  assign n7172 = ~pi122 & n5336;
  assign n7173 = ~pi043 & n7172;
  assign n7174 = ~n5518 & ~n7173;
  assign n7175 = ~n7171 & n7174;
  assign n7176 = n7169 & n7175;
  assign n7177 = pi039 & ~n7176;
  assign n7178 = ~n5511 & ~n6069;
  assign n7179 = n5354 & ~n7178;
  assign n7180 = ~pi043 & n5368;
  assign n7181 = ~n5410 & ~n7180;
  assign n7182 = ~n6083 & n7181;
  assign n7183 = ~pi122 & ~n7182;
  assign n7184 = ~n6404 & ~n7183;
  assign n7185 = n5381 & n5392;
  assign n7186 = n7184 & ~n7185;
  assign n7187 = ~pi039 & ~n7186;
  assign n7188 = ~n7179 & ~n7187;
  assign n7189 = ~n7177 & n7188;
  assign n7190 = ~n7168 & n7189;
  assign n7191 = ~n7133 & n7190;
  assign n7192 = n7106 & n7191;
  assign n7193 = n7102 & ~n7192;
  assign n7194 = ~n7102 & n7192;
  assign n7195 = ~n7193 & ~n7194;
  assign n7196 = ~n7004 & n7195;
  assign n7197 = n5772 & n7001;
  assign n7198 = ~n5772 & ~n7001;
  assign n7199 = ~n7197 & ~n7198;
  assign n7200 = ~n7195 & ~n7199;
  assign n7201 = ~n7196 & ~n7200;
  assign n7202 = n6909 & n7201;
  assign n7203 = ~n6909 & ~n7201;
  assign n7204 = ~n7202 & ~n7203;
  assign n7205 = ~pi529 & n7204;
  assign po136 = n6798 | n7205;
  assign n7207 = ~pi221 & pi432;
  assign n7208 = pi221 & ~pi432;
  assign n7209 = ~n7207 & ~n7208;
  assign n7210 = pi529 & ~n7209;
  assign n7211 = ~pi027 & n2012;
  assign n7212 = ~n1931 & ~n7211;
  assign n7213 = ~n1945 & n7212;
  assign n7214 = pi123 & ~n7213;
  assign n7215 = ~n2068 & ~n7214;
  assign n7216 = ~n2727 & n7215;
  assign n7217 = ~n1932 & n7216;
  assign n7218 = ~n3132 & ~n3174;
  assign n7219 = n7217 & n7218;
  assign n7220 = pi048 & ~n7219;
  assign n7221 = ~n2766 & ~n3068;
  assign n7222 = ~n3171 & n7221;
  assign n7223 = ~pi123 & ~n7222;
  assign n7224 = ~n3123 & ~n7223;
  assign n7225 = ~n7220 & n7224;
  assign n7226 = ~n2694 & ~n3114;
  assign n7227 = ~n2023 & ~n2704;
  assign n7228 = ~pi123 & ~n7227;
  assign n7229 = pi123 & n3092;
  assign n7230 = ~n1939 & ~n7229;
  assign n7231 = ~n3131 & n7230;
  assign n7232 = ~n7228 & n7231;
  assign n7233 = n7226 & n7232;
  assign n7234 = ~n2006 & n7233;
  assign n7235 = ~pi048 & ~n7234;
  assign n7236 = n7225 & ~n7235;
  assign n7237 = ~n1929 & ~n1976;
  assign n7238 = pi023 & ~n7237;
  assign n7239 = ~n2786 & ~n7238;
  assign n7240 = pi123 & ~n7239;
  assign n7241 = n7236 & ~n7240;
  assign n7242 = pi020 & ~n7241;
  assign n7243 = ~n1924 & ~n3171;
  assign n7244 = n1932 & n1975;
  assign n7245 = ~n1950 & ~n2038;
  assign n7246 = n1943 & ~n7245;
  assign n7247 = pi123 & n1917;
  assign n7248 = pi023 & n7247;
  assign n7249 = ~n7246 & ~n7248;
  assign n7250 = ~n7244 & n7249;
  assign n7251 = n7243 & n7250;
  assign n7252 = ~pi048 & ~n7251;
  assign n7253 = ~n1993 & ~n2031;
  assign n7254 = ~pi027 & n2003;
  assign n7255 = ~pi093 & ~pi111;
  assign n7256 = ~pi023 & n7255;
  assign n7257 = ~n7254 & ~n7256;
  assign n7258 = pi123 & ~n7257;
  assign n7259 = n7253 & ~n7258;
  assign n7260 = ~pi123 & n2781;
  assign n7261 = n7259 & ~n7260;
  assign n7262 = ~n2797 & n7261;
  assign n7263 = pi048 & ~n7262;
  assign n7264 = ~n7252 & ~n7263;
  assign n7265 = n1982 & n7256;
  assign n7266 = pi123 & n1992;
  assign n7267 = ~n7265 & ~n7266;
  assign n7268 = ~pi027 & n1977;
  assign n7269 = ~n1941 & ~n2698;
  assign n7270 = ~pi123 & ~n7269;
  assign n7271 = ~n7268 & ~n7270;
  assign n7272 = n7267 & n7271;
  assign n7273 = n7264 & n7272;
  assign n7274 = ~pi020 & ~n7273;
  assign n7275 = pi123 & n2050;
  assign n7276 = n1943 & n1977;
  assign n7277 = ~n7275 & ~n7276;
  assign n7278 = ~pi048 & ~n7277;
  assign n7279 = n1982 & n2721;
  assign n7280 = ~n2690 & ~n7279;
  assign n7281 = ~n7278 & n7280;
  assign n7282 = ~n2752 & n7281;
  assign n7283 = ~n2056 & ~n2781;
  assign n7284 = ~n3177 & n7283;
  assign n7285 = n3051 & ~n7284;
  assign n7286 = ~pi123 & n1988;
  assign n7287 = ~n7285 & ~n7286;
  assign n7288 = ~n2047 & n7287;
  assign n7289 = pi048 & ~n7288;
  assign n7290 = ~pi048 & ~pi123;
  assign n7291 = n2044 & n7290;
  assign n7292 = ~n7289 & ~n7291;
  assign n7293 = n1959 & n2032;
  assign n7294 = ~n2068 & ~n7293;
  assign n7295 = n2720 & ~n7294;
  assign n7296 = n7292 & ~n7295;
  assign n7297 = n7282 & n7296;
  assign n7298 = ~n7274 & n7297;
  assign n7299 = ~n7242 & n7298;
  assign n7300 = n3238 & n7299;
  assign n7301 = ~n3238 & ~n7299;
  assign n7302 = ~n7300 & ~n7301;
  assign n7303 = n1792 & n2945;
  assign n7304 = ~pi013 & n1835;
  assign n7305 = ~n1777 & ~n7304;
  assign n7306 = ~n1807 & n7305;
  assign n7307 = pi114 & ~n7306;
  assign n7308 = ~n1778 & ~n1890;
  assign n7309 = ~n2979 & n7308;
  assign n7310 = ~n7307 & n7309;
  assign n7311 = ~n2879 & ~n2911;
  assign n7312 = n7310 & n7311;
  assign n7313 = pi001 & ~n7312;
  assign n7314 = ~n1775 & ~n1862;
  assign n7315 = pi007 & ~n7314;
  assign n7316 = pi013 & n1774;
  assign n7317 = pi007 & n7316;
  assign n7318 = ~n7315 & ~n7317;
  assign n7319 = pi114 & ~n7318;
  assign n7320 = ~n2876 & ~n2961;
  assign n7321 = ~n2960 & n7320;
  assign n7322 = ~pi114 & ~n7321;
  assign n7323 = ~n7319 & ~n7322;
  assign n7324 = pi114 & n2821;
  assign n7325 = ~n1809 & ~n7324;
  assign n7326 = n1775 & n1838;
  assign n7327 = ~n1853 & ~n2848;
  assign n7328 = ~pi114 & ~n7327;
  assign n7329 = ~n3013 & ~n7328;
  assign n7330 = ~n7326 & n7329;
  assign n7331 = n7325 & n7330;
  assign n7332 = ~pi013 & n1794;
  assign n7333 = ~n3032 & ~n7332;
  assign n7334 = n7331 & n7333;
  assign n7335 = ~pi001 & ~n7334;
  assign n7336 = n7323 & ~n7335;
  assign n7337 = ~n7313 & n7336;
  assign n7338 = ~n7303 & n7337;
  assign n7339 = pi029 & ~n7338;
  assign n7340 = ~pi001 & ~pi114;
  assign n7341 = n1900 & n7340;
  assign n7342 = ~pi114 & n1830;
  assign n7343 = ~n1908 & ~n7342;
  assign n7344 = ~pi007 & n1777;
  assign n7345 = ~n2870 & ~n7344;
  assign n7346 = ~n1871 & n7345;
  assign n7347 = n1791 & ~n7346;
  assign n7348 = n7343 & ~n7347;
  assign n7349 = pi001 & ~n7348;
  assign n7350 = ~n7341 & ~n7349;
  assign n7351 = n1785 & n2945;
  assign n7352 = ~n1890 & ~n7351;
  assign n7353 = n2886 & ~n7352;
  assign n7354 = n1805 & n1863;
  assign n7355 = pi114 & n1878;
  assign n7356 = ~n7354 & ~n7355;
  assign n7357 = ~pi001 & ~n7356;
  assign n7358 = n1872 & n2827;
  assign n7359 = pi013 & n2922;
  assign n7360 = pi114 & n7359;
  assign n7361 = ~n7358 & ~n7360;
  assign n7362 = n1838 & n1862;
  assign n7363 = n7361 & ~n7362;
  assign n7364 = ~n7357 & n7363;
  assign n7365 = ~n7353 & n7364;
  assign n7366 = n7350 & n7365;
  assign n7367 = ~n1766 & ~n2876;
  assign n7368 = ~n1756 & ~n1896;
  assign n7369 = n1805 & ~n7368;
  assign n7370 = pi114 & n1901;
  assign n7371 = ~n7369 & ~n7370;
  assign n7372 = pi013 & ~pi114;
  assign n7373 = n1778 & n7372;
  assign n7374 = n7371 & ~n7373;
  assign n7375 = n7367 & n7374;
  assign n7376 = ~pi001 & ~n7375;
  assign n7377 = ~pi013 & n1863;
  assign n7378 = ~pi013 & n2831;
  assign n7379 = ~n1772 & ~n7378;
  assign n7380 = ~pi114 & ~n7379;
  assign n7381 = pi114 & n1824;
  assign n7382 = ~pi054 & ~pi098;
  assign n7383 = ~pi007 & n7382;
  assign n7384 = n2827 & n7383;
  assign n7385 = ~n7381 & ~n7384;
  assign n7386 = ~n7380 & n7385;
  assign n7387 = ~n7377 & n7386;
  assign n7388 = ~n7376 & n7387;
  assign n7389 = ~pi114 & n7344;
  assign n7390 = ~pi013 & n1847;
  assign n7391 = ~n7383 & ~n7390;
  assign n7392 = pi114 & ~n7391;
  assign n7393 = ~n1825 & ~n1881;
  assign n7394 = pi013 & n2831;
  assign n7395 = n7393 & ~n7394;
  assign n7396 = ~n7392 & n7395;
  assign n7397 = ~n7389 & n7396;
  assign n7398 = pi001 & ~n7397;
  assign n7399 = n7388 & ~n7398;
  assign n7400 = ~pi029 & ~n7399;
  assign n7401 = n7366 & ~n7400;
  assign n7402 = ~n7339 & n7401;
  assign n7403 = ~n2937 & n7402;
  assign n7404 = n2937 & ~n7402;
  assign n7405 = ~n7403 & ~n7404;
  assign n7406 = n7302 & n7405;
  assign n7407 = ~n7302 & ~n7405;
  assign n7408 = ~n7406 & ~n7407;
  assign n7409 = ~pi221 & ~n2243;
  assign n7410 = pi221 & n2243;
  assign n7411 = ~n7409 & ~n7410;
  assign n7412 = pi014 & n1605;
  assign n7413 = ~pi083 & n7412;
  assign n7414 = n1496 & n1508;
  assign n7415 = ~n7413 & ~n7414;
  assign n7416 = n1509 & n1665;
  assign n7417 = ~pi083 & n1533;
  assign n7418 = ~pi014 & n1529;
  assign n7419 = ~n1692 & ~n7418;
  assign n7420 = ~n1629 & n7419;
  assign n7421 = ~pi083 & ~n7420;
  assign n7422 = ~n1658 & ~n1731;
  assign n7423 = n1517 & n1545;
  assign n7424 = n7422 & ~n7423;
  assign n7425 = ~n7421 & n7424;
  assign n7426 = pi040 & ~n7425;
  assign n7427 = pi014 & n1663;
  assign n7428 = ~n1547 & ~n7427;
  assign n7429 = pi083 & n1496;
  assign n7430 = ~pi083 & n2668;
  assign n7431 = ~n7429 & ~n7430;
  assign n7432 = n7428 & n7431;
  assign n7433 = ~pi040 & ~n7432;
  assign n7434 = ~pi014 & n1575;
  assign n7435 = ~n1488 & ~n7434;
  assign n7436 = pi083 & ~n7435;
  assign n7437 = ~n7433 & ~n7436;
  assign n7438 = ~n7426 & n7437;
  assign n7439 = ~n7417 & n7438;
  assign n7440 = ~n7416 & n7439;
  assign n7441 = ~pi078 & ~n7440;
  assign n7442 = ~pi107 & n1521;
  assign n7443 = ~n1656 & ~n7442;
  assign n7444 = ~pi014 & ~pi108;
  assign n7445 = pi107 & n7444;
  assign n7446 = ~n1606 & ~n7445;
  assign n7447 = n7443 & n7446;
  assign n7448 = pi083 & ~n7447;
  assign n7449 = n1486 & n1665;
  assign n7450 = ~n2628 & ~n7449;
  assign n7451 = ~n1641 & n7450;
  assign n7452 = ~pi083 & ~n7451;
  assign n7453 = ~n7448 & ~n7452;
  assign n7454 = pi014 & n1616;
  assign n7455 = ~n1707 & ~n7454;
  assign n7456 = ~n1618 & ~n1701;
  assign n7457 = ~pi083 & ~n7456;
  assign n7458 = ~pi107 & n1528;
  assign n7459 = pi083 & n7458;
  assign n7460 = ~n7457 & ~n7459;
  assign n7461 = n7455 & n7460;
  assign n7462 = pi040 & ~n7461;
  assign n7463 = n1693 & n1742;
  assign n7464 = pi014 & n1476;
  assign n7465 = ~n7463 & ~n7464;
  assign n7466 = ~pi083 & n1541;
  assign n7467 = ~n1682 & ~n7466;
  assign n7468 = n7465 & n7467;
  assign n7469 = ~n1697 & n7468;
  assign n7470 = ~pi040 & ~n7469;
  assign n7471 = ~n7462 & ~n7470;
  assign n7472 = n7453 & n7471;
  assign n7473 = pi078 & ~n7472;
  assign n7474 = ~pi014 & n1519;
  assign n7475 = ~n2641 & ~n7474;
  assign n7476 = ~n1653 & n7475;
  assign n7477 = ~pi083 & ~n7476;
  assign n7478 = n1596 & n1665;
  assign n7479 = ~n1652 & ~n7478;
  assign n7480 = ~n1571 & ~n2608;
  assign n7481 = ~n1613 & n7480;
  assign n7482 = n7479 & n7481;
  assign n7483 = pi083 & ~n7482;
  assign n7484 = ~n1505 & ~n7416;
  assign n7485 = ~n7483 & n7484;
  assign n7486 = ~n7477 & n7485;
  assign n7487 = ~pi040 & ~n7486;
  assign n7488 = ~n7473 & ~n7487;
  assign n7489 = pi083 & n1554;
  assign n7490 = ~n1471 & ~n1518;
  assign n7491 = pi014 & ~n7490;
  assign n7492 = ~n1721 & ~n7491;
  assign n7493 = ~n7449 & n7492;
  assign n7494 = ~pi083 & ~n7493;
  assign n7495 = pi083 & n1610;
  assign n7496 = ~n1494 & ~n7495;
  assign n7497 = pi014 & n1692;
  assign n7498 = n7496 & ~n7497;
  assign n7499 = ~n7494 & n7498;
  assign n7500 = ~n7489 & n7499;
  assign n7501 = pi040 & ~n7500;
  assign n7502 = n7488 & ~n7501;
  assign n7503 = ~n7441 & n7502;
  assign n7504 = n7415 & n7503;
  assign n7505 = n2078 & n7504;
  assign n7506 = ~n2078 & ~n7504;
  assign n7507 = ~n7505 & ~n7506;
  assign n7508 = ~n7411 & n7507;
  assign n7509 = n7411 & ~n7507;
  assign n7510 = ~n7508 & ~n7509;
  assign n7511 = ~n7408 & n7510;
  assign n7512 = n7408 & ~n7510;
  assign n7513 = ~n7511 & ~n7512;
  assign n7514 = ~pi529 & n7513;
  assign po137 = n7210 | n7514;
  assign n7516 = ~pi121 & pi441;
  assign n7517 = pi121 & ~pi441;
  assign n7518 = ~n7516 & ~n7517;
  assign n7519 = pi529 & ~n7518;
  assign n7520 = pi107 & n1508;
  assign n7521 = n1492 & n7520;
  assign n7522 = ~n1718 & ~n2680;
  assign n7523 = pi014 & n1518;
  assign n7524 = n7522 & ~n7523;
  assign n7525 = ~pi083 & ~n7524;
  assign n7526 = ~n1530 & ~n7525;
  assign n7527 = ~n1588 & ~n2628;
  assign n7528 = pi083 & ~n7527;
  assign n7529 = n7526 & ~n7528;
  assign n7530 = pi040 & ~n7529;
  assign n7531 = ~pi083 & n7454;
  assign n7532 = ~n1629 & ~n7531;
  assign n7533 = n1463 & n1693;
  assign n7534 = ~n1478 & ~n7533;
  assign n7535 = ~pi040 & ~n7534;
  assign n7536 = n7532 & ~n7535;
  assign n7537 = ~n7530 & n7536;
  assign n7538 = ~n7521 & n7537;
  assign n7539 = ~pi078 & ~n7538;
  assign n7540 = ~n1471 & ~n1509;
  assign n7541 = n1665 & ~n7540;
  assign n7542 = pi083 & n7541;
  assign n7543 = ~n1694 & ~n7542;
  assign n7544 = n1587 & n7412;
  assign n7545 = n7543 & ~n7544;
  assign n7546 = ~pi014 & n1539;
  assign n7547 = ~n1493 & ~n7546;
  assign n7548 = n1587 & ~n7547;
  assign n7549 = n7545 & ~n7548;
  assign n7550 = ~n7539 & n7549;
  assign n7551 = ~pi083 & n1723;
  assign n7552 = n1528 & n1532;
  assign n7553 = ~n1614 & ~n7552;
  assign n7554 = ~pi083 & ~n7553;
  assign n7555 = ~n7551 & ~n7554;
  assign n7556 = ~n1653 & n7555;
  assign n7557 = pi040 & ~n7556;
  assign n7558 = pi014 & n1557;
  assign n7559 = ~n1505 & ~n1616;
  assign n7560 = ~n1673 & n7559;
  assign n7561 = ~pi083 & ~n7560;
  assign n7562 = pi014 & n1556;
  assign n7563 = ~n2641 & ~n7562;
  assign n7564 = ~n1478 & n7563;
  assign n7565 = pi083 & ~n7564;
  assign n7566 = n1509 & n1595;
  assign n7567 = ~n7565 & ~n7566;
  assign n7568 = ~n7561 & n7567;
  assign n7569 = ~n7558 & n7568;
  assign n7570 = ~n1692 & n7569;
  assign n7571 = ~pi040 & ~n7570;
  assign n7572 = ~n7557 & ~n7571;
  assign n7573 = ~pi083 & n1648;
  assign n7574 = n1482 & n7573;
  assign n7575 = pi083 & n1663;
  assign n7576 = ~pi014 & pi082;
  assign n7577 = pi107 & n7576;
  assign n7578 = ~n1557 & ~n7577;
  assign n7579 = ~pi083 & ~n7578;
  assign n7580 = ~n7575 & ~n7579;
  assign n7581 = ~n7574 & n7580;
  assign n7582 = pi040 & ~n7581;
  assign n7583 = ~n1467 & ~n1510;
  assign n7584 = ~n1680 & n7583;
  assign n7585 = n1508 & ~n7584;
  assign n7586 = ~n7416 & ~n7478;
  assign n7587 = ~n2647 & n7586;
  assign n7588 = ~n7585 & n7587;
  assign n7589 = ~pi107 & n1595;
  assign n7590 = n1485 & n7589;
  assign n7591 = pi083 & n1564;
  assign n7592 = ~n7459 & ~n7591;
  assign n7593 = ~n1658 & n7592;
  assign n7594 = ~n7590 & n7593;
  assign n7595 = ~pi083 & n1493;
  assign n7596 = ~n1465 & ~n2608;
  assign n7597 = ~n1682 & n7596;
  assign n7598 = ~n7595 & n7597;
  assign n7599 = n7594 & n7598;
  assign n7600 = ~pi040 & ~n7599;
  assign n7601 = n7588 & ~n7600;
  assign n7602 = ~n7582 & n7601;
  assign n7603 = pi078 & ~n7602;
  assign n7604 = n7572 & ~n7603;
  assign n7605 = n7550 & n7604;
  assign n7606 = n3238 & ~n7605;
  assign n7607 = ~n3238 & n7605;
  assign n7608 = ~n7606 & ~n7607;
  assign n7609 = ~pi027 & n3154;
  assign n7610 = ~n1952 & ~n7609;
  assign n7611 = n2720 & ~n7610;
  assign n7612 = ~pi123 & n2797;
  assign n7613 = n1928 & n3079;
  assign n7614 = ~n2721 & ~n7613;
  assign n7615 = ~pi123 & ~n7614;
  assign n7616 = ~n7612 & ~n7615;
  assign n7617 = ~n2023 & n7616;
  assign n7618 = pi048 & ~n7617;
  assign n7619 = pi123 & n1977;
  assign n7620 = n2726 & n7619;
  assign n7621 = ~n1918 & ~n1944;
  assign n7622 = n1916 & ~n7621;
  assign n7623 = pi123 & n7622;
  assign n7624 = ~n7286 & ~n7623;
  assign n7625 = ~n7620 & n7624;
  assign n7626 = ~n7618 & n7625;
  assign n7627 = ~n7611 & n7626;
  assign n7628 = pi027 & n3177;
  assign n7629 = pi027 & n2737;
  assign n7630 = ~n2021 & ~n7629;
  assign n7631 = ~n3132 & n7630;
  assign n7632 = pi123 & ~n7631;
  assign n7633 = ~n2004 & ~n2051;
  assign n7634 = ~n2786 & n7633;
  assign n7635 = ~pi123 & ~n7634;
  assign n7636 = n1918 & n3051;
  assign n7637 = ~n7635 & ~n7636;
  assign n7638 = ~n7632 & n7637;
  assign n7639 = ~n7628 & n7638;
  assign n7640 = ~n1930 & n7639;
  assign n7641 = ~pi048 & ~n7640;
  assign n7642 = pi123 & n3173;
  assign n7643 = ~pi123 & n1916;
  assign n7644 = n1917 & n7643;
  assign n7645 = ~n2055 & ~n7644;
  assign n7646 = ~n1939 & n7645;
  assign n7647 = ~n7642 & n7646;
  assign n7648 = ~pi123 & n1952;
  assign n7649 = ~n2011 & ~n3093;
  assign n7650 = ~n2044 & n7649;
  assign n7651 = ~n7648 & n7650;
  assign n7652 = n7647 & n7651;
  assign n7653 = ~pi048 & ~n7652;
  assign n7654 = pi123 & n1955;
  assign n7655 = pi047 & n3079;
  assign n7656 = ~n3177 & ~n7655;
  assign n7657 = ~pi123 & ~n7656;
  assign n7658 = ~n7654 & ~n7657;
  assign n7659 = ~n3124 & n7658;
  assign n7660 = pi048 & ~n7659;
  assign n7661 = ~n7653 & ~n7660;
  assign n7662 = ~n2701 & ~n2748;
  assign n7663 = ~n1991 & n7662;
  assign n7664 = n1982 & ~n7663;
  assign n7665 = ~n2008 & ~n2757;
  assign n7666 = ~n7664 & n7665;
  assign n7667 = ~n1919 & n7666;
  assign n7668 = n7661 & n7667;
  assign n7669 = pi020 & ~n7668;
  assign n7670 = pi023 & n1982;
  assign n7671 = n1951 & n7670;
  assign n7672 = ~n2801 & ~n7256;
  assign n7673 = ~n3084 & n7672;
  assign n7674 = ~pi123 & ~n7673;
  assign n7675 = ~n2776 & ~n7674;
  assign n7676 = ~n2067 & ~n3057;
  assign n7677 = pi123 & ~n7676;
  assign n7678 = n7675 & ~n7677;
  assign n7679 = pi048 & ~n7678;
  assign n7680 = ~pi123 & n2052;
  assign n7681 = ~n1932 & ~n7680;
  assign n7682 = n1975 & n2787;
  assign n7683 = ~n3132 & ~n7682;
  assign n7684 = ~pi048 & ~n7683;
  assign n7685 = n7681 & ~n7684;
  assign n7686 = ~n7679 & n7685;
  assign n7687 = ~n7671 & n7686;
  assign n7688 = ~pi020 & ~n7687;
  assign n7689 = ~n7669 & ~n7688;
  assign n7690 = ~n7641 & n7689;
  assign n7691 = n7627 & n7690;
  assign n7692 = n7402 & ~n7691;
  assign n7693 = ~n7402 & n7691;
  assign n7694 = ~n7692 & ~n7693;
  assign n7695 = ~n7608 & n7694;
  assign n7696 = n7608 & ~n7694;
  assign n7697 = ~n7695 & ~n7696;
  assign n7698 = ~pi121 & n2474;
  assign n7699 = pi121 & ~n2474;
  assign n7700 = ~n7698 & ~n7699;
  assign n7701 = ~n1755 & n7700;
  assign n7702 = n1755 & ~n7700;
  assign n7703 = ~n7701 & ~n7702;
  assign n7704 = ~n7697 & n7703;
  assign n7705 = n7697 & ~n7703;
  assign n7706 = ~n7704 & ~n7705;
  assign n7707 = ~pi529 & n7706;
  assign po138 = n7519 | n7707;
  assign n7709 = ~pi143 & pi412;
  assign n7710 = pi143 & ~pi412;
  assign n7711 = ~n7709 & ~n7710;
  assign n7712 = pi529 & ~n7711;
  assign n7713 = ~pi143 & ~n2365;
  assign n7714 = pi143 & n2365;
  assign n7715 = ~n7713 & ~n7714;
  assign n7716 = pi104 & ~pi127;
  assign n7717 = ~pi069 & n7716;
  assign n7718 = ~n2096 & ~n2160;
  assign n7719 = n7717 & ~n7718;
  assign n7720 = ~n2454 & ~n7719;
  assign n7721 = pi069 & n2251;
  assign n7722 = ~n2101 & ~n2207;
  assign n7723 = ~n2405 & n7722;
  assign n7724 = ~pi104 & ~n7723;
  assign n7725 = pi069 & n2250;
  assign n7726 = ~n2314 & ~n7725;
  assign n7727 = ~n2123 & n7726;
  assign n7728 = pi104 & ~n7727;
  assign n7729 = n2096 & n2135;
  assign n7730 = ~n7728 & ~n7729;
  assign n7731 = ~n7724 & n7730;
  assign n7732 = ~n7721 & n7731;
  assign n7733 = ~n2150 & n7732;
  assign n7734 = ~pi102 & ~n7733;
  assign n7735 = ~pi104 & n2420;
  assign n7736 = n2103 & n2200;
  assign n7737 = ~n2297 & ~n7736;
  assign n7738 = ~pi104 & ~n7737;
  assign n7739 = pi104 & n2088;
  assign n7740 = ~n2126 & ~n7739;
  assign n7741 = ~n7738 & n7740;
  assign n7742 = ~n7735 & n7741;
  assign n7743 = pi126 & n2105;
  assign n7744 = ~n2132 & ~n7743;
  assign n7745 = pi104 & ~n7744;
  assign n7746 = n7742 & ~n7745;
  assign n7747 = pi102 & ~n7746;
  assign n7748 = ~n7734 & ~n7747;
  assign n7749 = n7720 & n7748;
  assign n7750 = n2104 & n2105;
  assign n7751 = ~n2538 & ~n7750;
  assign n7752 = pi012 & n7751;
  assign n7753 = pi104 & n2138;
  assign n7754 = pi063 & n2200;
  assign n7755 = ~n2251 & ~n7754;
  assign n7756 = ~pi104 & ~n7755;
  assign n7757 = ~n7753 & ~n7756;
  assign n7758 = ~pi104 & n2373;
  assign n7759 = n7757 & ~n7758;
  assign n7760 = pi102 & ~n7759;
  assign n7761 = ~n2340 & ~n2461;
  assign n7762 = ~n2121 & n7761;
  assign n7763 = n2090 & ~n7762;
  assign n7764 = ~n2098 & ~n7763;
  assign n7765 = ~pi104 & n2396;
  assign n7766 = pi104 & n2255;
  assign n7767 = ~n2155 & ~n7766;
  assign n7768 = ~n2211 & n7767;
  assign n7769 = ~n2133 & ~n2232;
  assign n7770 = n7768 & n7769;
  assign n7771 = ~n7765 & n7770;
  assign n7772 = ~n2097 & ~n2308;
  assign n7773 = n7771 & n7772;
  assign n7774 = ~pi102 & ~n7773;
  assign n7775 = n7764 & ~n7774;
  assign n7776 = ~n7760 & n7775;
  assign n7777 = n7752 & n7776;
  assign n7778 = pi069 & n2117;
  assign n7779 = ~n2503 & ~n7778;
  assign n7780 = ~n2416 & n7779;
  assign n7781 = ~pi104 & ~n7780;
  assign n7782 = ~n2352 & ~n7781;
  assign n7783 = ~n2219 & ~n2267;
  assign n7784 = pi104 & ~n7783;
  assign n7785 = n7782 & ~n7784;
  assign n7786 = pi102 & ~n7785;
  assign n7787 = n2277 & n2388;
  assign n7788 = ~n2314 & ~n7787;
  assign n7789 = ~pi102 & ~n7788;
  assign n7790 = pi104 & n2191;
  assign n7791 = ~n7789 & ~n7790;
  assign n7792 = ~n7786 & n7791;
  assign n7793 = ~pi104 & n2208;
  assign n7794 = ~n2152 & ~n7793;
  assign n7795 = ~pi012 & n7794;
  assign n7796 = n7792 & n7795;
  assign n7797 = ~n7777 & ~n7796;
  assign n7798 = n7749 & ~n7797;
  assign n7799 = ~n1752 & n7798;
  assign n7800 = n1752 & ~n7798;
  assign n7801 = ~n7799 & ~n7800;
  assign n7802 = ~n7715 & n7801;
  assign n7803 = n7715 & ~n7801;
  assign n7804 = ~n7802 & ~n7803;
  assign n7805 = pi001 & n2827;
  assign n7806 = n1863 & n7805;
  assign n7807 = ~pi114 & n7394;
  assign n7808 = n1774 & n1877;
  assign n7809 = ~n2922 & ~n7808;
  assign n7810 = ~pi114 & ~n7809;
  assign n7811 = ~n7807 & ~n7810;
  assign n7812 = ~n1853 & n7811;
  assign n7813 = pi001 & ~n7812;
  assign n7814 = ~pi013 & n2835;
  assign n7815 = ~n1758 & ~n7814;
  assign n7816 = n2886 & ~n7815;
  assign n7817 = ~n1803 & ~n1806;
  assign n7818 = n1802 & ~n7817;
  assign n7819 = pi114 & n7818;
  assign n7820 = ~n7816 & ~n7819;
  assign n7821 = ~n7813 & n7820;
  assign n7822 = ~n7342 & n7821;
  assign n7823 = ~n7806 & n7822;
  assign n7824 = pi013 & n2870;
  assign n7825 = ~n1848 & ~n1869;
  assign n7826 = ~n7317 & n7825;
  assign n7827 = ~pi114 & ~n7826;
  assign n7828 = pi013 & n2869;
  assign n7829 = ~n1851 & ~n7828;
  assign n7830 = ~n2911 & n7829;
  assign n7831 = pi114 & ~n7830;
  assign n7832 = ~pi114 & n1842;
  assign n7833 = ~n7831 & ~n7832;
  assign n7834 = ~n7827 & n7833;
  assign n7835 = ~n7824 & n7834;
  assign n7836 = ~n1776 & n7835;
  assign n7837 = ~pi001 & ~n7836;
  assign n7838 = pi007 & n2827;
  assign n7839 = n1757 & n7838;
  assign n7840 = ~n2952 & ~n7383;
  assign n7841 = ~n3000 & n7840;
  assign n7842 = ~pi114 & ~n7841;
  assign n7843 = ~n2845 & ~n7842;
  assign n7844 = ~n1891 & ~n2887;
  assign n7845 = pi114 & ~n7844;
  assign n7846 = n7843 & ~n7845;
  assign n7847 = pi001 & ~n7846;
  assign n7848 = ~pi114 & n1870;
  assign n7849 = ~n1778 & ~n7848;
  assign n7850 = n2820 & n7372;
  assign n7851 = ~n2911 & ~n7850;
  assign n7852 = ~pi001 & ~n7851;
  assign n7853 = n7849 & ~n7852;
  assign n7854 = ~n7847 & n7853;
  assign n7855 = ~n7839 & n7854;
  assign n7856 = ~pi029 & ~n7855;
  assign n7857 = pi114 & n2878;
  assign n7858 = ~pi114 & n7332;
  assign n7859 = ~n1868 & ~n7858;
  assign n7860 = ~n1809 & n7859;
  assign n7861 = ~n7857 & n7860;
  assign n7862 = ~pi114 & n1758;
  assign n7863 = ~n1842 & ~n2822;
  assign n7864 = ~n1900 & n7863;
  assign n7865 = ~n7862 & n7864;
  assign n7866 = n7861 & n7865;
  assign n7867 = ~pi001 & ~n7866;
  assign n7868 = pi114 & n1794;
  assign n7869 = ~pi013 & pi021;
  assign n7870 = pi007 & n7869;
  assign n7871 = ~n2870 & ~n7870;
  assign n7872 = ~pi114 & ~n7871;
  assign n7873 = ~n7868 & ~n7872;
  assign n7874 = ~n3029 & n7873;
  assign n7875 = pi001 & ~n7874;
  assign n7876 = ~n7867 & ~n7875;
  assign n7877 = ~n1823 & ~n2830;
  assign n7878 = ~n2980 & n7877;
  assign n7879 = n2827 & ~n7878;
  assign n7880 = ~n1804 & ~n3031;
  assign n7881 = n1792 & n1805;
  assign n7882 = n7880 & ~n7881;
  assign n7883 = ~n7879 & n7882;
  assign n7884 = n7876 & n7883;
  assign n7885 = pi029 & ~n7884;
  assign n7886 = ~n7856 & ~n7885;
  assign n7887 = ~n7837 & n7886;
  assign n7888 = n7823 & n7887;
  assign n7889 = ~n2937 & n7888;
  assign n7890 = n2937 & ~n7888;
  assign n7891 = ~n7889 & ~n7890;
  assign n7892 = ~n7299 & n7402;
  assign n7893 = n7299 & ~n7402;
  assign n7894 = ~n7892 & ~n7893;
  assign n7895 = n7891 & n7894;
  assign n7896 = ~n7891 & ~n7894;
  assign n7897 = ~n7895 & ~n7896;
  assign n7898 = ~n7804 & n7897;
  assign n7899 = n7804 & ~n7897;
  assign n7900 = ~n7898 & ~n7899;
  assign n7901 = ~pi529 & n7900;
  assign po139 = n7712 | n7901;
  assign n7903 = ~pi150 & n2365;
  assign n7904 = pi150 & ~n2365;
  assign n7905 = ~n7903 & ~n7904;
  assign n7906 = ~pi014 & ~n1607;
  assign n7907 = ~n7463 & ~n7906;
  assign n7908 = ~pi040 & ~n7907;
  assign n7909 = ~pi014 & n1476;
  assign n7910 = ~n1529 & ~n7909;
  assign n7911 = n1491 & ~n7910;
  assign n7912 = ~n7908 & ~n7911;
  assign n7913 = ~n1509 & ~n1518;
  assign n7914 = n1648 & ~n7913;
  assign n7915 = pi083 & n7914;
  assign n7916 = ~pi014 & n2624;
  assign n7917 = n1631 & ~n7916;
  assign n7918 = ~pi083 & ~n7917;
  assign n7919 = pi072 & n1508;
  assign n7920 = n1481 & n7919;
  assign n7921 = n1471 & n1595;
  assign n7922 = ~n1588 & ~n1663;
  assign n7923 = pi107 & n2680;
  assign n7924 = n7922 & ~n7923;
  assign n7925 = ~n7921 & n7924;
  assign n7926 = ~n7920 & n7925;
  assign n7927 = pi040 & ~n7926;
  assign n7928 = ~n7918 & ~n7927;
  assign n7929 = ~n7915 & n7928;
  assign n7930 = n7912 & n7929;
  assign n7931 = ~pi078 & ~n7930;
  assign n7932 = ~n2668 & ~n7497;
  assign n7933 = ~n1511 & ~n1585;
  assign n7934 = ~pi083 & ~n7933;
  assign n7935 = ~n1630 & ~n2590;
  assign n7936 = ~n1542 & n7935;
  assign n7937 = ~n1692 & n7936;
  assign n7938 = pi083 & ~n7937;
  assign n7939 = ~n1504 & ~n2633;
  assign n7940 = ~n1493 & n7939;
  assign n7941 = pi083 & ~n7940;
  assign n7942 = pi014 & ~pi072;
  assign n7943 = ~pi107 & n7942;
  assign n7944 = pi014 & n7458;
  assign n7945 = ~n7943 & ~n7944;
  assign n7946 = ~n1465 & n7945;
  assign n7947 = n1595 & n1618;
  assign n7948 = n7946 & ~n7947;
  assign n7949 = ~n7941 & n7948;
  assign n7950 = ~pi040 & ~n7949;
  assign n7951 = pi014 & n2634;
  assign n7952 = ~n7523 & ~n7951;
  assign n7953 = ~pi083 & ~n7952;
  assign n7954 = ~n7950 & ~n7953;
  assign n7955 = ~pi083 & n1495;
  assign n7956 = ~n1680 & ~n7955;
  assign n7957 = ~n1636 & n7956;
  assign n7958 = pi040 & ~n7957;
  assign n7959 = n7954 & ~n7958;
  assign n7960 = ~n7938 & n7959;
  assign n7961 = ~n7934 & n7960;
  assign n7962 = n7932 & n7961;
  assign n7963 = pi078 & ~n7962;
  assign n7964 = ~n7931 & ~n7963;
  assign n7965 = n1523 & n1532;
  assign n7966 = pi083 & ~n7965;
  assign n7967 = ~pi083 & ~n1478;
  assign n7968 = ~n7966 & ~n7967;
  assign n7969 = ~n7454 & ~n7968;
  assign n7970 = ~n1657 & n7969;
  assign n7971 = ~n7449 & n7970;
  assign n7972 = pi040 & ~n7971;
  assign n7973 = ~n1666 & ~n7478;
  assign n7974 = pi083 & ~n7973;
  assign n7975 = ~pi014 & n1523;
  assign n7976 = ~n7416 & ~n7975;
  assign n7977 = ~n1554 & n7976;
  assign n7978 = ~pi083 & ~n7977;
  assign n7979 = ~n7974 & ~n7978;
  assign n7980 = ~n7574 & n7979;
  assign n7981 = ~n2618 & n7980;
  assign n7982 = ~pi040 & ~n7981;
  assign n7983 = ~n7972 & ~n7982;
  assign n7984 = n7964 & n7983;
  assign n7985 = pi083 & ~n1484;
  assign n7986 = ~pi083 & ~n7923;
  assign n7987 = ~n7985 & ~n7986;
  assign n7988 = n7984 & ~n7987;
  assign n7989 = ~n3141 & n7988;
  assign n7990 = n3141 & ~n7988;
  assign n7991 = ~n7989 & ~n7990;
  assign n7992 = ~n3043 & n7991;
  assign n7993 = ~n3245 & ~n7991;
  assign n7994 = ~n7992 & ~n7993;
  assign n7995 = ~n7905 & n7994;
  assign n7996 = n7905 & ~n7994;
  assign po141 = ~n7995 & ~n7996;
  assign n7998 = ~pi150 & pi483;
  assign n7999 = pi150 & ~pi483;
  assign po143 = n7998 | n7999;
  assign n8001 = ~pi137 & pi495;
  assign n8002 = pi137 & ~pi495;
  assign n8003 = ~n8001 & ~n8002;
  assign n8004 = pi529 & ~n8003;
  assign n8005 = ~n1627 & n7605;
  assign n8006 = n1627 & ~n7605;
  assign n8007 = ~n8005 & ~n8006;
  assign n8008 = n7894 & ~n8007;
  assign n8009 = ~n7894 & n8007;
  assign n8010 = ~n8008 & ~n8009;
  assign n8011 = ~n2365 & n7798;
  assign n8012 = n2365 & ~n7798;
  assign n8013 = ~n8011 & ~n8012;
  assign n8014 = ~pi137 & n2474;
  assign n8015 = pi137 & ~n2474;
  assign n8016 = ~n8014 & ~n8015;
  assign n8017 = ~n8013 & n8016;
  assign n8018 = n8013 & ~n8016;
  assign n8019 = ~n8017 & ~n8018;
  assign n8020 = ~n8010 & n8019;
  assign n8021 = n8010 & ~n8019;
  assign n8022 = ~n8020 & ~n8021;
  assign n8023 = ~pi529 & n8022;
  assign po144 = n8004 | n8023;
  assign n8025 = pi075 & n3385;
  assign n8026 = ~pi079 & n3269;
  assign n8027 = ~n8025 & ~n8026;
  assign n8028 = pi079 & n3309;
  assign n8029 = pi042 & ~pi075;
  assign n8030 = ~n8028 & ~n8029;
  assign n8031 = n8027 & n8030;
  assign n8032 = n3257 & ~n8031;
  assign n8033 = pi075 & n3309;
  assign n8034 = ~pi079 & n8033;
  assign n8035 = ~pi080 & n8034;
  assign n8036 = ~n8032 & ~n8035;
  assign n8037 = ~pi080 & n3272;
  assign n8038 = ~pi079 & n3309;
  assign n8039 = ~pi080 & n8038;
  assign n8040 = ~n8037 & ~n8039;
  assign n8041 = pi079 & n3276;
  assign n8042 = ~n8034 & ~n8041;
  assign n8043 = n8040 & n8042;
  assign n8044 = ~n3264 & ~n8025;
  assign n8045 = ~n8033 & n8044;
  assign n8046 = ~pi080 & ~n8045;
  assign n8047 = n3353 & n3401;
  assign n8048 = ~n8046 & ~n8047;
  assign n8049 = n8043 & n8048;
  assign n8050 = ~pi073 & ~n8049;
  assign n8051 = pi075 & n3272;
  assign n8052 = ~pi075 & n3258;
  assign n8053 = ~pi079 & n8052;
  assign n8054 = pi075 & n3275;
  assign n8055 = ~pi079 & n8054;
  assign n8056 = ~n8053 & ~n8055;
  assign n8057 = ~n8051 & n8056;
  assign n8058 = pi080 & ~n8057;
  assign n8059 = ~pi075 & n3350;
  assign n8060 = n3288 & n8059;
  assign n8061 = pi075 & ~pi079;
  assign n8062 = n3339 & n8061;
  assign n8063 = ~n8060 & ~n8062;
  assign n8064 = ~n8058 & n8063;
  assign n8065 = pi079 & n3260;
  assign n8066 = n3297 & n3366;
  assign n8067 = ~n8065 & ~n8066;
  assign n8068 = pi073 & ~n8067;
  assign n8069 = n8064 & ~n8068;
  assign n8070 = ~n8050 & n8069;
  assign n8071 = n8036 & n8070;
  assign n8072 = pi015 & ~n8071;
  assign n8073 = pi075 & n3352;
  assign n8074 = n3288 & n8073;
  assign n8075 = pi080 & n3270;
  assign n8076 = ~n8074 & ~n8075;
  assign n8077 = ~pi073 & ~n8076;
  assign n8078 = ~pi075 & n3339;
  assign n8079 = ~pi079 & n8078;
  assign n8080 = ~n3379 & ~n8079;
  assign n8081 = ~pi080 & ~n8080;
  assign n8082 = pi079 & n8051;
  assign n8083 = ~n3316 & ~n8082;
  assign n8084 = ~pi080 & ~n8083;
  assign n8085 = ~n8081 & ~n8084;
  assign n8086 = ~pi075 & ~pi080;
  assign n8087 = pi110 & n8086;
  assign n8088 = ~n3314 & ~n8087;
  assign n8089 = ~pi073 & ~n8088;
  assign n8090 = ~n3294 & ~n3307;
  assign n8091 = n3288 & ~n8090;
  assign n8092 = ~n3289 & ~n8091;
  assign n8093 = ~n8089 & n8092;
  assign n8094 = n8085 & n8093;
  assign n8095 = ~n8077 & n8094;
  assign n8096 = ~n3261 & ~n3327;
  assign n8097 = n3351 & n3401;
  assign n8098 = ~pi042 & n3302;
  assign n8099 = ~n3311 & ~n8098;
  assign n8100 = ~pi080 & ~n8099;
  assign n8101 = ~n8097 & ~n8100;
  assign n8102 = n8096 & n8101;
  assign n8103 = pi073 & ~n8102;
  assign n8104 = n8095 & ~n8103;
  assign n8105 = ~pi015 & ~n8104;
  assign n8106 = pi079 & n3353;
  assign n8107 = ~pi080 & n8106;
  assign n8108 = ~n8081 & ~n8107;
  assign n8109 = ~pi079 & n3378;
  assign n8110 = n8108 & ~n8109;
  assign n8111 = ~pi073 & ~n8110;
  assign n8112 = pi079 & n3278;
  assign n8113 = ~n3329 & ~n3368;
  assign n8114 = ~n8054 & n8113;
  assign n8115 = pi079 & ~n8114;
  assign n8116 = ~n8112 & ~n8115;
  assign n8117 = pi073 & ~pi080;
  assign n8118 = ~n8116 & n8117;
  assign n8119 = ~n8111 & ~n8118;
  assign n8120 = n3270 & n3302;
  assign n8121 = n3272 & n3395;
  assign n8122 = ~n8120 & ~n8121;
  assign n8123 = ~pi080 & ~n8122;
  assign n8124 = ~pi079 & n3264;
  assign n8125 = ~n8065 & ~n8124;
  assign n8126 = ~n3373 & n8125;
  assign n8127 = n3290 & ~n8126;
  assign n8128 = ~n8123 & ~n8127;
  assign n8129 = ~n3262 & ~n3372;
  assign n8130 = ~pi075 & n3278;
  assign n8131 = ~n8052 & ~n8130;
  assign n8132 = pi075 & n3297;
  assign n8133 = n8131 & ~n8132;
  assign n8134 = ~pi079 & ~n8133;
  assign n8135 = n8129 & ~n8134;
  assign n8136 = n3257 & ~n8135;
  assign n8137 = n8128 & ~n8136;
  assign n8138 = n8119 & n8137;
  assign n8139 = ~n8105 & n8138;
  assign n8140 = ~n8072 & n8139;
  assign n8141 = pi190 & n8140;
  assign n8142 = ~pi190 & ~n8140;
  assign n8143 = ~n8141 & ~n8142;
  assign n8144 = ~pi085 & n3426;
  assign n8145 = pi028 & n8144;
  assign n8146 = ~n3565 & ~n8145;
  assign n8147 = n3468 & n3555;
  assign n8148 = ~n3441 & ~n8147;
  assign n8149 = ~pi092 & ~n8148;
  assign n8150 = ~n3451 & ~n3497;
  assign n8151 = ~n3458 & n8150;
  assign n8152 = ~n8144 & n8151;
  assign n8153 = pi092 & ~n8152;
  assign n8154 = ~pi087 & ~pi092;
  assign n8155 = ~pi050 & n8154;
  assign n8156 = ~pi046 & n8155;
  assign n8157 = ~pi092 & n3471;
  assign n8158 = ~n3502 & ~n8157;
  assign n8159 = ~n8156 & n8158;
  assign n8160 = pi089 & ~n8159;
  assign n8161 = pi085 & n3467;
  assign n8162 = pi085 & n3482;
  assign n8163 = ~n3542 & ~n8162;
  assign n8164 = ~n8161 & n8163;
  assign n8165 = pi092 & ~n8164;
  assign n8166 = pi028 & ~pi087;
  assign n8167 = ~pi085 & n8166;
  assign n8168 = ~pi085 & n3425;
  assign n8169 = pi028 & n8168;
  assign n8170 = ~n8167 & ~n8169;
  assign n8171 = ~pi085 & n3555;
  assign n8172 = ~pi028 & n8171;
  assign n8173 = n8170 & ~n8172;
  assign n8174 = ~pi028 & ~pi092;
  assign n8175 = n3427 & n8174;
  assign n8176 = n8173 & ~n8175;
  assign n8177 = ~n8165 & n8176;
  assign n8178 = ~pi089 & ~n8177;
  assign n8179 = pi028 & n3543;
  assign n8180 = pi028 & n3526;
  assign n8181 = ~n8179 & ~n8180;
  assign n8182 = ~pi092 & ~n8181;
  assign n8183 = ~n8178 & ~n8182;
  assign n8184 = ~n8160 & n8183;
  assign n8185 = ~n8153 & n8184;
  assign n8186 = ~n8149 & n8185;
  assign n8187 = n8146 & n8186;
  assign n8188 = pi053 & ~n8187;
  assign n8189 = pi085 & n3430;
  assign n8190 = n3488 & n8189;
  assign n8191 = ~n3493 & ~n3553;
  assign n8192 = ~pi028 & ~n8191;
  assign n8193 = ~n8190 & ~n8192;
  assign n8194 = ~pi089 & ~n8193;
  assign n8195 = ~pi028 & n3456;
  assign n8196 = ~n3495 & ~n8195;
  assign n8197 = n3446 & ~n8196;
  assign n8198 = ~n8194 & ~n8197;
  assign n8199 = pi028 & ~pi085;
  assign n8200 = ~n3449 & ~n3526;
  assign n8201 = n8199 & ~n8200;
  assign n8202 = pi092 & n8201;
  assign n8203 = ~pi087 & n3436;
  assign n8204 = ~pi046 & n8203;
  assign n8205 = pi028 & n3440;
  assign n8206 = ~n3497 & ~n8205;
  assign n8207 = ~n8204 & n8206;
  assign n8208 = ~pi092 & ~n8207;
  assign n8209 = pi087 & n3433;
  assign n8210 = n3453 & n8209;
  assign n8211 = n3575 & n8174;
  assign n8212 = ~pi085 & n3430;
  assign n8213 = ~pi028 & n3430;
  assign n8214 = ~n8212 & ~n8213;
  assign n8215 = pi085 & n3578;
  assign n8216 = n8214 & ~n8215;
  assign n8217 = ~n8211 & n8216;
  assign n8218 = ~n8210 & n8217;
  assign n8219 = pi089 & ~n8218;
  assign n8220 = ~n8208 & ~n8219;
  assign n8221 = ~n8202 & n8220;
  assign n8222 = n8198 & n8221;
  assign n8223 = ~pi053 & ~n8222;
  assign n8224 = ~pi085 & n3565;
  assign n8225 = pi092 & ~n8224;
  assign n8226 = ~pi092 & ~n8215;
  assign n8227 = ~n8225 & ~n8226;
  assign n8228 = ~n8223 & ~n8227;
  assign n8229 = ~n8188 & n8228;
  assign n8230 = pi028 & n3426;
  assign n8231 = pi092 & n8230;
  assign n8232 = ~pi085 & n3449;
  assign n8233 = pi028 & n8232;
  assign n8234 = n3454 & n3468;
  assign n8235 = pi092 & ~n8234;
  assign n8236 = ~pi028 & n3521;
  assign n8237 = ~pi092 & ~n8236;
  assign n8238 = ~n8235 & ~n8237;
  assign n8239 = ~n8233 & ~n8238;
  assign n8240 = ~n8231 & n8239;
  assign n8241 = n3431 & n3436;
  assign n8242 = n8240 & ~n8241;
  assign n8243 = pi089 & ~n8242;
  assign n8244 = ~pi092 & n8199;
  assign n8245 = pi087 & n8244;
  assign n8246 = n3453 & n8245;
  assign n8247 = n3426 & n3436;
  assign n8248 = n3436 & n3471;
  assign n8249 = ~n8247 & ~n8248;
  assign n8250 = pi092 & ~n8249;
  assign n8251 = ~pi028 & n3454;
  assign n8252 = n3436 & n3449;
  assign n8253 = ~n8251 & ~n8252;
  assign n8254 = pi085 & n3453;
  assign n8255 = ~pi028 & n8254;
  assign n8256 = n8253 & ~n8255;
  assign n8257 = ~pi092 & ~n8256;
  assign n8258 = ~n8250 & ~n8257;
  assign n8259 = ~n8246 & n8258;
  assign n8260 = ~n3547 & n8259;
  assign n8261 = ~pi089 & ~n8260;
  assign n8262 = ~n8243 & ~n8261;
  assign n8263 = n8229 & n8262;
  assign n8264 = ~n4161 & n8263;
  assign n8265 = n4161 & ~n8263;
  assign n8266 = ~n8264 & ~n8265;
  assign n8267 = ~n4045 & n8266;
  assign n8268 = ~n4274 & ~n8266;
  assign n8269 = ~n8267 & ~n8268;
  assign n8270 = ~n8143 & n8269;
  assign n8271 = n8143 & ~n8269;
  assign po145 = ~n8270 & ~n8271;
  assign n8273 = pi190 & pi410;
  assign n8274 = ~pi190 & ~pi410;
  assign po146 = n8273 | n8274;
  assign n8276 = ~pi136 & pi438;
  assign n8277 = pi136 & ~pi438;
  assign n8278 = ~n8276 & ~n8277;
  assign n8279 = pi529 & ~n8278;
  assign n8280 = n3238 & n7691;
  assign n8281 = ~n3238 & ~n7691;
  assign n8282 = ~n8280 & ~n8281;
  assign n8283 = n7891 & n8282;
  assign n8284 = ~n7891 & ~n8282;
  assign n8285 = ~n8283 & ~n8284;
  assign n8286 = n1752 & ~n7299;
  assign n8287 = ~n1752 & n7299;
  assign n8288 = ~n8286 & ~n8287;
  assign n8289 = ~pi136 & ~n2474;
  assign n8290 = pi136 & n2474;
  assign n8291 = ~n8289 & ~n8290;
  assign n8292 = n8288 & n8291;
  assign n8293 = ~n8288 & ~n8291;
  assign n8294 = ~n8292 & ~n8293;
  assign n8295 = ~n8285 & n8294;
  assign n8296 = n8285 & ~n8294;
  assign n8297 = ~n8295 & ~n8296;
  assign n8298 = ~pi529 & n8297;
  assign po147 = n8279 | n8298;
  assign n8300 = ~pi171 & pi443;
  assign n8301 = pi171 & ~pi443;
  assign n8302 = ~n8300 & ~n8301;
  assign n8303 = pi529 & ~n8302;
  assign n8304 = ~pi019 & pi049;
  assign n8305 = n4439 & n8304;
  assign n8306 = pi049 & n4331;
  assign n8307 = ~pi049 & n4309;
  assign n8308 = ~pi019 & n8307;
  assign n8309 = pi049 & n4334;
  assign n8310 = ~pi019 & n8309;
  assign n8311 = ~n8308 & ~n8310;
  assign n8312 = ~n8306 & n8311;
  assign n8313 = pi090 & ~n8312;
  assign n8314 = ~pi049 & n4383;
  assign n8315 = n4322 & n8314;
  assign n8316 = ~n8313 & ~n8315;
  assign n8317 = ~n8305 & n8316;
  assign n8318 = pi049 & n4387;
  assign n8319 = pi049 & n4294;
  assign n8320 = ~n8318 & ~n8319;
  assign n8321 = ~n4315 & n8320;
  assign n8322 = ~pi090 & ~n8321;
  assign n8323 = ~pi090 & n4331;
  assign n8324 = ~pi019 & pi090;
  assign n8325 = n4426 & n8324;
  assign n8326 = ~pi019 & n4294;
  assign n8327 = ~pi090 & n8326;
  assign n8328 = ~n8325 & ~n8327;
  assign n8329 = ~n8323 & n8328;
  assign n8330 = ~n8322 & n8329;
  assign n8331 = pi019 & n4335;
  assign n8332 = ~pi019 & n8319;
  assign n8333 = ~n8331 & ~n8332;
  assign n8334 = n8330 & n8333;
  assign n8335 = ~pi088 & ~n8334;
  assign n8336 = n8317 & ~n8335;
  assign n8337 = ~pi019 & n4286;
  assign n8338 = ~n8318 & ~n8337;
  assign n8339 = pi019 & n4294;
  assign n8340 = ~pi049 & pi112;
  assign n8341 = ~n8339 & ~n8340;
  assign n8342 = n8338 & n8341;
  assign n8343 = n4319 & ~n8342;
  assign n8344 = pi019 & n4311;
  assign n8345 = ~pi019 & ~pi090;
  assign n8346 = n4292 & n8345;
  assign n8347 = ~n8344 & ~n8346;
  assign n8348 = pi088 & ~n8347;
  assign n8349 = ~n8343 & ~n8348;
  assign n8350 = ~pi090 & n8332;
  assign n8351 = n8349 & ~n8350;
  assign n8352 = n8336 & n8351;
  assign n8353 = pi006 & ~n8352;
  assign n8354 = ~n4313 & ~n4392;
  assign n8355 = pi049 & n4292;
  assign n8356 = ~n8307 & ~n8355;
  assign n8357 = ~pi049 & n4287;
  assign n8358 = n8356 & ~n8357;
  assign n8359 = ~pi019 & ~n8358;
  assign n8360 = n8354 & ~n8359;
  assign n8361 = n4319 & ~n8360;
  assign n8362 = n4290 & n4297;
  assign n8363 = ~pi019 & ~pi049;
  assign n8364 = n4331 & n8363;
  assign n8365 = ~n8362 & ~n8364;
  assign n8366 = ~pi090 & ~n8365;
  assign n8367 = ~n8361 & ~n8366;
  assign n8368 = ~pi019 & n4315;
  assign n8369 = ~n4391 & ~n8368;
  assign n8370 = ~n8344 & n8369;
  assign n8371 = n4343 & ~n8370;
  assign n8372 = ~pi049 & n4439;
  assign n8373 = ~pi019 & n8372;
  assign n8374 = ~n4397 & ~n8373;
  assign n8375 = ~pi090 & ~n8374;
  assign n8376 = pi019 & n4426;
  assign n8377 = ~pi090 & n8376;
  assign n8378 = ~n8375 & ~n8377;
  assign n8379 = ~pi019 & n4398;
  assign n8380 = n8378 & ~n8379;
  assign n8381 = ~pi088 & ~n8380;
  assign n8382 = ~n4356 & ~n4416;
  assign n8383 = ~n8309 & n8382;
  assign n8384 = pi019 & ~n8383;
  assign n8385 = pi019 & n4287;
  assign n8386 = ~n8384 & ~n8385;
  assign n8387 = pi088 & ~pi090;
  assign n8388 = ~n8386 & n8387;
  assign n8389 = ~n8381 & ~n8388;
  assign n8390 = ~n8371 & n8389;
  assign n8391 = n8367 & n8390;
  assign n8392 = ~n4312 & ~n4414;
  assign n8393 = n4384 & n8324;
  assign n8394 = pi019 & ~pi112;
  assign n8395 = pi049 & n8394;
  assign n8396 = ~n4296 & ~n8395;
  assign n8397 = ~pi090 & ~n8396;
  assign n8398 = ~n8393 & ~n8397;
  assign n8399 = n8392 & n8398;
  assign n8400 = pi088 & ~n8399;
  assign n8401 = pi049 & n4425;
  assign n8402 = n4322 & n8401;
  assign n8403 = pi090 & n4297;
  assign n8404 = ~n8402 & ~n8403;
  assign n8405 = ~pi088 & ~n8404;
  assign n8406 = ~pi049 & pi051;
  assign n8407 = ~pi090 & n8406;
  assign n8408 = ~n4303 & ~n8407;
  assign n8409 = ~pi088 & ~n8408;
  assign n8410 = ~n8405 & ~n8409;
  assign n8411 = ~n8400 & n8410;
  assign n8412 = pi019 & n8306;
  assign n8413 = ~n4298 & ~n8412;
  assign n8414 = ~pi090 & ~n8413;
  assign n8415 = ~n8375 & ~n8414;
  assign n8416 = ~n4288 & ~n4348;
  assign n8417 = n4322 & ~n8416;
  assign n8418 = ~n4325 & ~n8417;
  assign n8419 = n8415 & n8418;
  assign n8420 = n8411 & n8419;
  assign n8421 = ~pi006 & ~n8420;
  assign n8422 = n8391 & ~n8421;
  assign n8423 = ~n8353 & n8422;
  assign n8424 = ~n4287 & ~n4425;
  assign n8425 = n8363 & ~n8424;
  assign n8426 = pi090 & n8425;
  assign n8427 = ~pi049 & n4292;
  assign n8428 = n4328 & n8427;
  assign n8429 = ~n8426 & ~n8428;
  assign n8430 = pi019 & n4416;
  assign n8431 = pi090 & n8430;
  assign n8432 = n4291 & n8304;
  assign n8433 = ~n4313 & ~n8432;
  assign n8434 = ~pi090 & ~n8433;
  assign n8435 = ~pi090 & n4423;
  assign n8436 = ~n4365 & ~n8435;
  assign n8437 = ~n8434 & n8436;
  assign n8438 = ~n8431 & n8437;
  assign n8439 = ~pi019 & n8406;
  assign n8440 = ~n4311 & ~n8439;
  assign n8441 = pi090 & ~n8440;
  assign n8442 = n8438 & ~n8441;
  assign n8443 = pi088 & ~n8442;
  assign n8444 = n8429 & ~n8443;
  assign n8445 = ~pi049 & n8345;
  assign n8446 = n4286 & n8445;
  assign n8447 = pi090 & n8326;
  assign n8448 = ~pi049 & n4291;
  assign n8449 = pi090 & n8448;
  assign n8450 = ~n8447 & ~n8449;
  assign n8451 = pi090 & n4331;
  assign n8452 = n8450 & ~n8451;
  assign n8453 = ~pi090 & n4311;
  assign n8454 = n8452 & ~n8453;
  assign n8455 = ~n4330 & n8454;
  assign n8456 = ~n8446 & n8455;
  assign n8457 = pi019 & n8307;
  assign n8458 = ~n8373 & ~n8457;
  assign n8459 = n8456 & n8458;
  assign n8460 = ~pi088 & ~n8459;
  assign n8461 = pi019 & ~pi049;
  assign n8462 = ~pi090 & n8461;
  assign n8463 = n4331 & n8462;
  assign n8464 = ~pi019 & pi112;
  assign n8465 = pi049 & n8464;
  assign n8466 = ~n8318 & ~n8465;
  assign n8467 = ~pi090 & ~n8466;
  assign n8468 = pi090 & n4344;
  assign n8469 = ~n8467 & ~n8468;
  assign n8470 = ~n8463 & n8469;
  assign n8471 = pi088 & ~n8470;
  assign n8472 = ~n8460 & ~n8471;
  assign n8473 = n4292 & n8363;
  assign n8474 = ~pi019 & n8357;
  assign n8475 = ~n4288 & ~n4367;
  assign n8476 = ~n4347 & n8475;
  assign n8477 = n4322 & ~n8476;
  assign n8478 = ~n4377 & ~n8477;
  assign n8479 = ~n8474 & n8478;
  assign n8480 = ~n8473 & n8479;
  assign n8481 = pi006 & n8480;
  assign n8482 = n8472 & n8481;
  assign n8483 = n4328 & n4439;
  assign n8484 = ~n8379 & ~n8483;
  assign n8485 = ~pi088 & ~n8484;
  assign n8486 = pi019 & n8357;
  assign n8487 = ~pi090 & n8486;
  assign n8488 = ~n4360 & ~n8487;
  assign n8489 = pi049 & n4322;
  assign n8490 = n4310 & n8489;
  assign n8491 = n8488 & ~n8490;
  assign n8492 = ~pi051 & n4415;
  assign n8493 = ~n4424 & ~n8492;
  assign n8494 = pi019 & n4383;
  assign n8495 = n8493 & ~n8494;
  assign n8496 = ~pi090 & ~n8495;
  assign n8497 = ~n4414 & ~n8496;
  assign n8498 = ~n4394 & ~n8337;
  assign n8499 = pi090 & ~n8498;
  assign n8500 = n8497 & ~n8499;
  assign n8501 = pi088 & ~n8500;
  assign n8502 = n8491 & ~n8501;
  assign n8503 = ~n8485 & n8502;
  assign n8504 = ~pi006 & n8503;
  assign n8505 = ~n8482 & ~n8504;
  assign n8506 = pi019 & n8318;
  assign n8507 = ~n4442 & ~n8357;
  assign n8508 = ~n8412 & n8507;
  assign n8509 = ~pi090 & ~n8508;
  assign n8510 = ~n8506 & ~n8509;
  assign n8511 = n4287 & n8345;
  assign n8512 = pi019 & n4387;
  assign n8513 = ~n8379 & ~n8512;
  assign n8514 = ~n4357 & n8513;
  assign n8515 = pi090 & ~n8514;
  assign n8516 = ~n8427 & ~n8515;
  assign n8517 = ~n8511 & n8516;
  assign n8518 = n8510 & n8517;
  assign n8519 = ~pi088 & ~n8518;
  assign n8520 = ~n8505 & ~n8519;
  assign n8521 = n8444 & n8520;
  assign n8522 = ~n8423 & n8521;
  assign n8523 = n8423 & ~n8521;
  assign n8524 = ~n8522 & ~n8523;
  assign n8525 = n4416 & n8324;
  assign n8526 = pi090 & n4299;
  assign n8527 = ~n8525 & ~n8526;
  assign n8528 = ~pi088 & ~n8527;
  assign n8529 = n4313 & n4322;
  assign n8530 = ~n4370 & ~n8529;
  assign n8531 = ~n8528 & n8530;
  assign n8532 = ~n4393 & ~n8318;
  assign n8533 = ~n4436 & n8532;
  assign n8534 = n8345 & ~n8533;
  assign n8535 = ~n8428 & ~n8534;
  assign n8536 = n4314 & n8461;
  assign n8537 = ~n4371 & ~n8536;
  assign n8538 = pi090 & ~n8537;
  assign n8539 = pi090 & n4360;
  assign n8540 = ~n8538 & ~n8539;
  assign n8541 = n8535 & n8540;
  assign n8542 = pi088 & ~n8541;
  assign n8543 = ~pi088 & ~pi090;
  assign n8544 = n8457 & n8543;
  assign n8545 = ~n4326 & ~n8544;
  assign n8546 = ~n8542 & n8545;
  assign n8547 = n4331 & n8461;
  assign n8548 = ~pi090 & n4297;
  assign n8549 = ~pi019 & n4334;
  assign n8550 = ~n4359 & ~n8549;
  assign n8551 = ~n8401 & n8550;
  assign n8552 = pi090 & ~n8551;
  assign n8553 = ~n8327 & ~n8552;
  assign n8554 = ~n8379 & n8553;
  assign n8555 = ~n8548 & n8554;
  assign n8556 = ~n4360 & ~n4371;
  assign n8557 = n8555 & n8556;
  assign n8558 = pi088 & ~n8557;
  assign n8559 = n4295 & n4328;
  assign n8560 = pi090 & n8372;
  assign n8561 = n4292 & n4322;
  assign n8562 = ~n8560 & ~n8561;
  assign n8563 = ~n8451 & n8562;
  assign n8564 = ~pi086 & n8345;
  assign n8565 = n4309 & n8564;
  assign n8566 = n8563 & ~n8565;
  assign n8567 = ~n4345 & n8566;
  assign n8568 = ~n8559 & n8567;
  assign n8569 = n4314 & n8363;
  assign n8570 = ~n4293 & ~n8569;
  assign n8571 = n8568 & n8570;
  assign n8572 = ~pi088 & ~n8571;
  assign n8573 = ~pi019 & n4426;
  assign n8574 = pi019 & n4347;
  assign n8575 = ~n8573 & ~n8574;
  assign n8576 = ~pi019 & n4360;
  assign n8577 = n8575 & ~n8576;
  assign n8578 = ~pi090 & ~n8577;
  assign n8579 = ~n8572 & ~n8578;
  assign n8580 = ~n8558 & n8579;
  assign n8581 = ~n8547 & n8580;
  assign n8582 = ~n4292 & ~n4295;
  assign n8583 = pi049 & ~n8582;
  assign n8584 = ~n4442 & ~n8583;
  assign n8585 = pi090 & ~n8584;
  assign n8586 = n8581 & ~n8585;
  assign n8587 = pi006 & ~n8586;
  assign n8588 = n4328 & n4360;
  assign n8589 = ~n4301 & ~n4309;
  assign n8590 = n8324 & ~n8589;
  assign n8591 = pi049 & pi090;
  assign n8592 = n4286 & n8591;
  assign n8593 = ~n8590 & ~n8592;
  assign n8594 = ~n4298 & ~n8573;
  assign n8595 = n8593 & n8594;
  assign n8596 = ~n8588 & n8595;
  assign n8597 = ~pi088 & ~n8596;
  assign n8598 = n4331 & n8304;
  assign n8599 = ~n8492 & ~n8598;
  assign n8600 = pi090 & ~n8599;
  assign n8601 = ~pi090 & n4436;
  assign n8602 = pi019 & n4292;
  assign n8603 = n4347 & n8363;
  assign n8604 = ~n8602 & ~n8603;
  assign n8605 = ~n8601 & n8604;
  assign n8606 = ~n8600 & n8605;
  assign n8607 = ~n4423 & n8606;
  assign n8608 = pi088 & ~n8607;
  assign n8609 = ~n8597 & ~n8608;
  assign n8610 = ~pi019 & n4416;
  assign n8611 = pi019 & n8319;
  assign n8612 = ~n4349 & ~n8611;
  assign n8613 = ~pi090 & ~n8612;
  assign n8614 = pi090 & n4356;
  assign n8615 = n4322 & n8492;
  assign n8616 = ~n8614 & ~n8615;
  assign n8617 = ~n8613 & n8616;
  assign n8618 = ~n8610 & n8617;
  assign n8619 = n8609 & n8618;
  assign n8620 = ~pi006 & ~n8619;
  assign n8621 = ~n8587 & ~n8620;
  assign n8622 = n8546 & n8621;
  assign n8623 = n8531 & n8622;
  assign n8624 = ~pi171 & ~n8623;
  assign n8625 = pi171 & n8623;
  assign n8626 = ~n8624 & ~n8625;
  assign n8627 = ~n8524 & n8626;
  assign n8628 = n8524 & ~n8626;
  assign n8629 = ~n8627 & ~n8628;
  assign n8630 = ~n4502 & ~n4549;
  assign n8631 = ~pi000 & n4498;
  assign n8632 = ~pi000 & n4456;
  assign n8633 = ~n8631 & ~n8632;
  assign n8634 = ~n4461 & n8633;
  assign n8635 = ~pi011 & ~n8634;
  assign n8636 = n8630 & ~n8635;
  assign n8637 = pi116 & ~n8636;
  assign n8638 = pi000 & n4486;
  assign n8639 = ~n4525 & ~n4582;
  assign n8640 = ~n8638 & n8639;
  assign n8641 = pi011 & ~n8640;
  assign n8642 = pi011 & n4456;
  assign n8643 = ~n8641 & ~n8642;
  assign n8644 = ~pi116 & ~n8643;
  assign n8645 = ~n8637 & ~n8644;
  assign n8646 = pi058 & ~n8645;
  assign n8647 = pi022 & n4512;
  assign n8648 = n4464 & n8647;
  assign n8649 = pi011 & n4472;
  assign n8650 = ~n8648 & ~n8649;
  assign n8651 = ~pi116 & ~n8650;
  assign n8652 = pi000 & n4499;
  assign n8653 = pi011 & n8652;
  assign n8654 = ~pi011 & n4504;
  assign n8655 = ~n8653 & ~n8654;
  assign n8656 = ~n4551 & n8655;
  assign n8657 = n4511 & ~n8656;
  assign n8658 = ~pi000 & n4584;
  assign n8659 = ~pi011 & n8658;
  assign n8660 = ~n4554 & ~n8659;
  assign n8661 = ~pi116 & ~n8660;
  assign n8662 = ~pi011 & n4553;
  assign n8663 = pi011 & n4603;
  assign n8664 = ~pi116 & n8663;
  assign n8665 = ~n8662 & ~n8664;
  assign n8666 = ~n8661 & n8665;
  assign n8667 = ~pi058 & ~n8666;
  assign n8668 = ~n8657 & ~n8667;
  assign n8669 = ~n8651 & n8668;
  assign n8670 = ~pi000 & n4558;
  assign n8671 = n4481 & n8670;
  assign n8672 = ~pi011 & n8631;
  assign n8673 = ~pi011 & n8638;
  assign n8674 = ~n8672 & ~n8673;
  assign n8675 = pi000 & n4490;
  assign n8676 = n8674 & ~n8675;
  assign n8677 = pi116 & ~n8676;
  assign n8678 = ~n8671 & ~n8677;
  assign n8679 = n4500 & n4584;
  assign n8680 = n8678 & ~n8679;
  assign n8681 = pi000 & n4464;
  assign n8682 = ~pi011 & n8681;
  assign n8683 = ~pi116 & n8682;
  assign n8684 = pi000 & n4478;
  assign n8685 = ~n4504 & ~n8684;
  assign n8686 = ~n8681 & n8685;
  assign n8687 = ~pi116 & ~n8686;
  assign n8688 = ~pi116 & n4490;
  assign n8689 = ~pi011 & n4603;
  assign n8690 = pi116 & n8689;
  assign n8691 = ~pi011 & n4464;
  assign n8692 = ~pi116 & n8691;
  assign n8693 = ~n8690 & ~n8692;
  assign n8694 = ~n8688 & n8693;
  assign n8695 = ~n8687 & n8694;
  assign n8696 = pi011 & n4487;
  assign n8697 = ~n8682 & ~n8696;
  assign n8698 = n8695 & n8697;
  assign n8699 = ~pi058 & ~n8698;
  assign n8700 = ~pi011 & n4455;
  assign n8701 = ~n8684 & ~n8700;
  assign n8702 = pi011 & n4464;
  assign n8703 = ~pi000 & pi057;
  assign n8704 = ~n8702 & ~n8703;
  assign n8705 = n8701 & n8704;
  assign n8706 = n4508 & ~n8705;
  assign n8707 = ~pi011 & ~pi116;
  assign n8708 = n4460 & n8707;
  assign n8709 = ~n8653 & ~n8708;
  assign n8710 = pi058 & ~n8709;
  assign n8711 = ~n8706 & ~n8710;
  assign n8712 = ~n8699 & n8711;
  assign n8713 = ~n8683 & n8712;
  assign n8714 = n8680 & n8713;
  assign n8715 = pi060 & ~n8714;
  assign n8716 = pi011 & n8675;
  assign n8717 = ~n4472 & ~n8716;
  assign n8718 = ~pi116 & ~n8717;
  assign n8719 = ~n4457 & ~n4518;
  assign n8720 = n4481 & ~n8719;
  assign n8721 = ~n4482 & ~n8720;
  assign n8722 = n4540 & n4559;
  assign n8723 = pi011 & ~pi057;
  assign n8724 = pi000 & n8723;
  assign n8725 = ~n4466 & ~n8724;
  assign n8726 = ~pi116 & ~n8725;
  assign n8727 = ~n8722 & ~n8726;
  assign n8728 = ~n4595 & n8727;
  assign n8729 = ~n4501 & n8728;
  assign n8730 = pi058 & ~n8729;
  assign n8731 = ~n8661 & ~n8730;
  assign n8732 = n8721 & n8731;
  assign n8733 = ~n8718 & n8732;
  assign n8734 = ~pi000 & pi097;
  assign n8735 = ~pi116 & n8734;
  assign n8736 = ~n4469 & ~n8735;
  assign n8737 = ~pi058 & ~n8736;
  assign n8738 = pi000 & n4602;
  assign n8739 = n4481 & n8738;
  assign n8740 = pi116 & n4471;
  assign n8741 = ~n8739 & ~n8740;
  assign n8742 = ~pi058 & ~n8741;
  assign n8743 = ~n8737 & ~n8742;
  assign n8744 = n8733 & n8743;
  assign n8745 = ~pi060 & ~n8744;
  assign n8746 = ~n8715 & ~n8745;
  assign n8747 = n8669 & n8746;
  assign n8748 = ~n8646 & n8747;
  assign n8749 = ~pi000 & pi011;
  assign n8750 = ~pi116 & n8749;
  assign n8751 = pi022 & n8750;
  assign n8752 = n4464 & n8751;
  assign n8753 = ~pi000 & n4455;
  assign n8754 = pi116 & n8753;
  assign n8755 = ~pi011 & pi057;
  assign n8756 = pi000 & n8755;
  assign n8757 = ~n8684 & ~n8756;
  assign n8758 = ~pi116 & ~n8757;
  assign n8759 = ~n8754 & ~n8758;
  assign n8760 = ~n8752 & n8759;
  assign n8761 = pi058 & ~n8760;
  assign n8762 = ~n4457 & ~n4517;
  assign n8763 = ~n4534 & n8762;
  assign n8764 = n4481 & ~n8763;
  assign n8765 = n4460 & n4512;
  assign n8766 = n4456 & n4512;
  assign n8767 = ~n8765 & ~n8766;
  assign n8768 = ~n4541 & n8767;
  assign n8769 = ~n8764 & n8768;
  assign n8770 = pi116 & n8691;
  assign n8771 = pi116 & n4490;
  assign n8772 = ~pi116 & n4514;
  assign n8773 = ~pi000 & n4459;
  assign n8774 = pi116 & n8773;
  assign n8775 = ~n8772 & ~n8774;
  assign n8776 = ~n8771 & n8775;
  assign n8777 = ~n8770 & n8776;
  assign n8778 = ~pi116 & n8652;
  assign n8779 = ~n4489 & ~n8659;
  assign n8780 = pi011 & n8631;
  assign n8781 = n8779 & ~n8780;
  assign n8782 = ~n8778 & n8781;
  assign n8783 = n8777 & n8782;
  assign n8784 = ~pi058 & ~n8783;
  assign n8785 = n8769 & ~n8784;
  assign n8786 = ~n8761 & n8785;
  assign n8787 = pi060 & ~n8786;
  assign n8788 = pi000 & n4481;
  assign n8789 = n4499 & n8788;
  assign n8790 = ~pi022 & ~pi097;
  assign n8791 = ~pi000 & n8790;
  assign n8792 = ~n4605 & ~n8791;
  assign n8793 = pi011 & n4558;
  assign n8794 = n8792 & ~n8793;
  assign n8795 = ~pi116 & ~n8794;
  assign n8796 = ~n4595 & ~n8795;
  assign n8797 = ~n4548 & ~n8700;
  assign n8798 = pi116 & ~n8797;
  assign n8799 = n8796 & ~n8798;
  assign n8800 = pi058 & ~n8799;
  assign n8801 = pi011 & n8632;
  assign n8802 = ~pi116 & n8801;
  assign n8803 = ~n4528 & ~n8802;
  assign n8804 = n4484 & n4584;
  assign n8805 = ~n8662 & ~n8804;
  assign n8806 = ~pi058 & ~n8805;
  assign n8807 = n8803 & ~n8806;
  assign n8808 = ~n8800 & n8807;
  assign n8809 = ~n8789 & n8808;
  assign n8810 = ~pi060 & ~n8809;
  assign n8811 = ~n8787 & ~n8810;
  assign n8812 = pi011 & n4582;
  assign n8813 = n4508 & n8812;
  assign n8814 = ~pi011 & n8734;
  assign n8815 = ~n8652 & ~n8814;
  assign n8816 = n4508 & ~n8815;
  assign n8817 = ~pi116 & n4608;
  assign n8818 = n4459 & n4500;
  assign n8819 = ~n4502 & ~n8818;
  assign n8820 = ~pi116 & ~n8819;
  assign n8821 = ~n8817 & ~n8820;
  assign n8822 = ~n4535 & n8821;
  assign n8823 = pi058 & ~n8822;
  assign n8824 = ~pi000 & n4460;
  assign n8825 = n4484 & n8824;
  assign n8826 = ~n4456 & ~n4602;
  assign n8827 = n4512 & ~n8826;
  assign n8828 = pi116 & n8827;
  assign n8829 = ~n8825 & ~n8828;
  assign n8830 = ~n8823 & n8829;
  assign n8831 = ~n8816 & n8830;
  assign n8832 = pi011 & n8684;
  assign n8833 = ~n8632 & ~n8716;
  assign n8834 = ~n4581 & n8833;
  assign n8835 = ~pi116 & ~n8834;
  assign n8836 = pi011 & n4478;
  assign n8837 = ~n4526 & ~n8836;
  assign n8838 = ~n8662 & n8837;
  assign n8839 = pi116 & ~n8838;
  assign n8840 = n4456 & n8707;
  assign n8841 = ~n8839 & ~n8840;
  assign n8842 = ~n8835 & n8841;
  assign n8843 = ~n8832 & n8842;
  assign n8844 = ~n8824 & n8843;
  assign n8845 = ~pi058 & ~n8844;
  assign n8846 = n8831 & ~n8845;
  assign n8847 = ~n8813 & n8846;
  assign n8848 = n8811 & n8847;
  assign n8849 = ~n8748 & n8848;
  assign n8850 = n8748 & ~n8848;
  assign n8851 = ~n8849 & ~n8850;
  assign n8852 = ~n4624 & ~n5081;
  assign n8853 = ~n4637 & ~n4657;
  assign n8854 = ~pi118 & ~n8853;
  assign n8855 = pi118 & n4675;
  assign n8856 = pi118 & n5143;
  assign n8857 = ~n5170 & ~n8856;
  assign n8858 = ~n8855 & n8857;
  assign n8859 = ~n8854 & n8858;
  assign n8860 = n8852 & n8859;
  assign n8861 = ~n4648 & n8860;
  assign n8862 = ~pi034 & ~n8861;
  assign n8863 = ~n4630 & ~n4636;
  assign n8864 = pi103 & ~n8863;
  assign n8865 = ~n4666 & ~n8864;
  assign n8866 = pi118 & ~n8865;
  assign n8867 = ~pi066 & n4659;
  assign n8868 = ~n4660 & ~n8867;
  assign n8869 = ~n5225 & n8868;
  assign n8870 = pi118 & ~n8869;
  assign n8871 = ~n5171 & ~n5275;
  assign n8872 = ~n4715 & n8871;
  assign n8873 = ~n8870 & n8872;
  assign n8874 = ~n4706 & ~n4771;
  assign n8875 = n8873 & n8874;
  assign n8876 = pi034 & ~n8875;
  assign n8877 = ~n4707 & ~n5272;
  assign n8878 = ~n5116 & n8877;
  assign n8879 = ~pi118 & ~n8878;
  assign n8880 = ~n8876 & ~n8879;
  assign n8881 = ~n5184 & n8880;
  assign n8882 = ~n8866 & n8881;
  assign n8883 = ~n8862 & n8882;
  assign n8884 = pi038 & ~n8883;
  assign n8885 = ~pi066 & n4704;
  assign n8886 = ~n5169 & ~n8885;
  assign n8887 = ~pi066 & n5147;
  assign n8888 = ~pi103 & n4748;
  assign n8889 = ~n8887 & ~n8888;
  assign n8890 = pi118 & ~n8889;
  assign n8891 = ~n4695 & ~n8890;
  assign n8892 = ~pi118 & n4661;
  assign n8893 = n8891 & ~n8892;
  assign n8894 = n8886 & n8893;
  assign n8895 = pi034 & ~n8894;
  assign n8896 = pi066 & ~pi118;
  assign n8897 = n4706 & n8896;
  assign n8898 = ~n4643 & ~n5272;
  assign n8899 = ~n4625 & ~n4638;
  assign n8900 = n5249 & ~n8899;
  assign n8901 = pi118 & n4622;
  assign n8902 = pi103 & n8901;
  assign n8903 = ~n8900 & ~n8902;
  assign n8904 = n8898 & n8903;
  assign n8905 = ~n8897 & n8904;
  assign n8906 = ~pi034 & ~n8905;
  assign n8907 = ~n8895 & ~n8906;
  assign n8908 = ~pi066 & n4667;
  assign n8909 = pi066 & n5180;
  assign n8910 = ~n4628 & ~n8909;
  assign n8911 = ~pi118 & ~n8910;
  assign n8912 = ~n8908 & ~n8911;
  assign n8913 = pi118 & n4704;
  assign n8914 = n4753 & n8888;
  assign n8915 = ~n8913 & ~n8914;
  assign n8916 = n8912 & n8915;
  assign n8917 = n8907 & n8916;
  assign n8918 = ~pi038 & ~n8917;
  assign n8919 = n4667 & n5249;
  assign n8920 = pi118 & n4644;
  assign n8921 = ~n8919 & ~n8920;
  assign n8922 = ~pi034 & ~n8921;
  assign n8923 = n4686 & n4753;
  assign n8924 = ~n4758 & ~n8923;
  assign n8925 = ~n8922 & n8924;
  assign n8926 = ~n4714 & n8925;
  assign n8927 = pi118 & n4706;
  assign n8928 = ~pi118 & n5123;
  assign n8929 = ~n8927 & ~n8928;
  assign n8930 = ~n4661 & ~n4723;
  assign n8931 = ~n5267 & n8930;
  assign n8932 = n5090 & ~n8931;
  assign n8933 = n8929 & ~n8932;
  assign n8934 = pi034 & ~n8933;
  assign n8935 = pi066 & n5200;
  assign n8936 = ~pi034 & ~pi118;
  assign n8937 = n8935 & n8936;
  assign n8938 = ~n8934 & ~n8937;
  assign n8939 = n4763 & n5103;
  assign n8940 = ~n4715 & ~n8939;
  assign n8941 = n4762 & ~n8940;
  assign n8942 = n8938 & ~n8941;
  assign n8943 = n8926 & n8942;
  assign n8944 = ~n8918 & n8943;
  assign n8945 = ~n8884 & n8944;
  assign n8946 = n4828 & n4901;
  assign n8947 = pi120 & n8946;
  assign n8948 = n4815 & n4928;
  assign n8949 = ~n8947 & ~n8948;
  assign n8950 = ~pi003 & ~n8949;
  assign n8951 = n4807 & n4905;
  assign n8952 = pi074 & n4798;
  assign n8953 = pi120 & n8952;
  assign n8954 = ~n8951 & ~n8953;
  assign n8955 = n4814 & n5007;
  assign n8956 = n8954 & ~n8955;
  assign n8957 = ~n8950 & n8956;
  assign n8958 = ~pi041 & ~pi045;
  assign n8959 = ~pi016 & n8958;
  assign n8960 = n4905 & n8959;
  assign n8961 = ~pi074 & n4914;
  assign n8962 = pi074 & n4861;
  assign n8963 = ~n8961 & ~n8962;
  assign n8964 = ~pi120 & ~n8963;
  assign n8965 = ~pi074 & n4815;
  assign n8966 = ~n8964 & ~n8965;
  assign n8967 = pi074 & ~pi120;
  assign n8968 = n4975 & n8967;
  assign n8969 = ~n4856 & ~n4870;
  assign n8970 = ~n4796 & ~n4843;
  assign n8971 = n4928 & ~n8970;
  assign n8972 = pi120 & n4959;
  assign n8973 = ~n8971 & ~n8972;
  assign n8974 = n8969 & n8973;
  assign n8975 = ~n8968 & n8974;
  assign n8976 = ~pi003 & ~n8975;
  assign n8977 = pi120 & n4817;
  assign n8978 = ~n8976 & ~n8977;
  assign n8979 = n8966 & n8978;
  assign n8980 = ~n8960 & n8979;
  assign n8981 = ~pi074 & n4817;
  assign n8982 = ~n5043 & ~n8981;
  assign n8983 = ~pi016 & n4920;
  assign n8984 = ~pi120 & n8983;
  assign n8985 = ~pi074 & n4898;
  assign n8986 = ~n8959 & ~n8985;
  assign n8987 = pi120 & ~n8986;
  assign n8988 = ~n8984 & ~n8987;
  assign n8989 = pi074 & n4914;
  assign n8990 = n8988 & ~n8989;
  assign n8991 = n8982 & n8990;
  assign n8992 = pi003 & ~n8991;
  assign n8993 = n8980 & ~n8992;
  assign n8994 = ~pi044 & ~n8993;
  assign n8995 = ~pi074 & n4812;
  assign n8996 = ~n4920 & ~n8995;
  assign n8997 = ~n4947 & n8996;
  assign n8998 = pi120 & ~n8997;
  assign n8999 = pi074 & n4797;
  assign n9000 = ~n8998 & ~n8999;
  assign n9001 = ~n5001 & n9000;
  assign n9002 = ~n4975 & n9001;
  assign n9003 = ~n4845 & ~n4873;
  assign n9004 = n9002 & n9003;
  assign n9005 = pi003 & ~n9004;
  assign n9006 = ~n4870 & ~n4976;
  assign n9007 = ~n4974 & n9006;
  assign n9008 = ~pi120 & ~n9007;
  assign n9009 = pi120 & n4838;
  assign n9010 = pi120 & n4794;
  assign n9011 = ~n9009 & ~n9010;
  assign n9012 = n4806 & n5007;
  assign n9013 = ~pi074 & n4797;
  assign n9014 = ~n4925 & ~n9013;
  assign n9015 = ~pi120 & ~n9014;
  assign n9016 = ~n9012 & ~n9015;
  assign n9017 = ~n5044 & n9016;
  assign n9018 = n9011 & n9017;
  assign n9019 = ~pi074 & n4983;
  assign n9020 = ~n5066 & ~n9019;
  assign n9021 = n9018 & n9020;
  assign n9022 = ~pi003 & ~n9021;
  assign n9023 = n4794 & n4969;
  assign n9024 = ~n9022 & ~n9023;
  assign n9025 = ~n9008 & n9024;
  assign n9026 = ~n9005 & n9025;
  assign n9027 = ~n4806 & ~n4814;
  assign n9028 = pi016 & ~n9027;
  assign n9029 = pi074 & n4805;
  assign n9030 = pi016 & n9029;
  assign n9031 = ~n9028 & ~n9030;
  assign n9032 = pi120 & ~n9031;
  assign n9033 = n9026 & ~n9032;
  assign n9034 = pi044 & ~n9033;
  assign n9035 = ~pi003 & ~pi120;
  assign n9036 = pi074 & n4800;
  assign n9037 = n9035 & n9036;
  assign n9038 = ~pi120 & n4996;
  assign n9039 = pi120 & n4975;
  assign n9040 = ~n9038 & ~n9039;
  assign n9041 = ~n4865 & ~n8983;
  assign n9042 = ~pi016 & n4793;
  assign n9043 = n9041 & ~n9042;
  assign n9044 = n4890 & ~n9043;
  assign n9045 = n9040 & ~n9044;
  assign n9046 = pi003 & ~n9045;
  assign n9047 = ~n9037 & ~n9046;
  assign n9048 = n4830 & n4969;
  assign n9049 = ~n8999 & ~n9048;
  assign n9050 = n4882 & ~n9049;
  assign n9051 = n9047 & ~n9050;
  assign n9052 = ~n9034 & n9051;
  assign n9053 = ~n8994 & n9052;
  assign n9054 = n8957 & n9053;
  assign n9055 = ~n8945 & n9054;
  assign n9056 = n8945 & ~n9054;
  assign n9057 = ~n9055 & ~n9056;
  assign n9058 = ~n8851 & n9057;
  assign n9059 = n8851 & ~n9057;
  assign n9060 = ~n9058 & ~n9059;
  assign n9061 = n8629 & n9060;
  assign n9062 = ~n8629 & ~n9060;
  assign n9063 = ~n9061 & ~n9062;
  assign n9064 = ~pi529 & n9063;
  assign po148 = n8303 | n9064;
  assign n9066 = ~pi187 & n8423;
  assign n9067 = pi187 & ~n8423;
  assign n9068 = ~n9066 & ~n9067;
  assign n9069 = pi000 & n4455;
  assign n9070 = n4484 & n9069;
  assign n9071 = ~pi011 & ~n8639;
  assign n9072 = ~n9070 & ~n9071;
  assign n9073 = ~pi058 & ~n9072;
  assign n9074 = ~pi011 & n4467;
  assign n9075 = ~n4527 & ~n9074;
  assign n9076 = n4511 & ~n9075;
  assign n9077 = ~n9073 & ~n9076;
  assign n9078 = ~n4456 & ~n4558;
  assign n9079 = n8749 & ~n9078;
  assign n9080 = pi116 & n9079;
  assign n9081 = ~pi011 & n4562;
  assign n9082 = pi011 & n4517;
  assign n9083 = ~n4529 & ~n9082;
  assign n9084 = ~n9081 & n9083;
  assign n9085 = ~pi116 & ~n9084;
  assign n9086 = n4602 & n8707;
  assign n9087 = pi000 & n4605;
  assign n9088 = pi116 & n4549;
  assign n9089 = ~n9087 & ~n9088;
  assign n9090 = ~n9086 & n9089;
  assign n9091 = ~n8700 & ~n8753;
  assign n9092 = n9090 & n9091;
  assign n9093 = pi058 & ~n9092;
  assign n9094 = ~n9085 & ~n9093;
  assign n9095 = ~n9080 & n9094;
  assign n9096 = n9077 & n9095;
  assign n9097 = ~pi060 & ~n9096;
  assign n9098 = n4503 & n4512;
  assign n9099 = ~n8765 & ~n9098;
  assign n9100 = pi116 & ~n9099;
  assign n9101 = ~pi011 & n4465;
  assign n9102 = ~n8766 & ~n9101;
  assign n9103 = ~n8682 & n9102;
  assign n9104 = ~pi116 & ~n9103;
  assign n9105 = ~n9100 & ~n9104;
  assign n9106 = ~n8752 & n9105;
  assign n9107 = ~n4576 & n9106;
  assign n9108 = ~pi058 & ~n9107;
  assign n9109 = ~n9097 & ~n9108;
  assign n9110 = pi011 & n4571;
  assign n9111 = ~n8793 & ~n9110;
  assign n9112 = ~pi116 & ~n9111;
  assign n9113 = pi011 & n8773;
  assign n9114 = pi011 & ~pi022;
  assign n9115 = ~pi000 & n9114;
  assign n9116 = ~n8659 & ~n9115;
  assign n9117 = ~n9113 & n9116;
  assign n9118 = n4461 & n8707;
  assign n9119 = ~n4573 & ~n8675;
  assign n9120 = ~n8652 & n9119;
  assign n9121 = pi116 & ~n9120;
  assign n9122 = ~n9118 & ~n9121;
  assign n9123 = n9117 & n9122;
  assign n9124 = ~pi058 & ~n9123;
  assign n9125 = ~n9112 & ~n9124;
  assign n9126 = ~n4529 & ~n8824;
  assign n9127 = ~n4469 & n9126;
  assign n9128 = ~n4458 & n9127;
  assign n9129 = pi116 & ~n9128;
  assign n9130 = ~n4518 & ~n8679;
  assign n9131 = ~pi116 & ~n9130;
  assign n9132 = ~n9129 & ~n9131;
  assign n9133 = pi011 & n8824;
  assign n9134 = ~n4594 & ~n9133;
  assign n9135 = ~pi116 & n4503;
  assign n9136 = ~pi022 & ~pi116;
  assign n9137 = ~pi097 & n9136;
  assign n9138 = ~pi057 & n9137;
  assign n9139 = ~n9135 & ~n9138;
  assign n9140 = ~n4534 & n9139;
  assign n9141 = pi058 & ~n9140;
  assign n9142 = n9134 & ~n9141;
  assign n9143 = n9132 & n9142;
  assign n9144 = n9125 & n9143;
  assign n9145 = pi060 & ~n9144;
  assign n9146 = ~pi116 & n8662;
  assign n9147 = n4465 & n4500;
  assign n9148 = pi116 & n9147;
  assign n9149 = pi011 & n4460;
  assign n9150 = pi116 & n9149;
  assign n9151 = ~n8801 & ~n9150;
  assign n9152 = ~n9148 & n9151;
  assign n9153 = ~n9146 & n9152;
  assign n9154 = n4471 & n4512;
  assign n9155 = n9153 & ~n9154;
  assign n9156 = pi058 & ~n9155;
  assign n9157 = ~n9145 & ~n9156;
  assign n9158 = n9109 & n9157;
  assign n9159 = pi116 & ~n8648;
  assign n9160 = ~pi116 & ~n9087;
  assign n9161 = ~n9159 & ~n9160;
  assign n9162 = n9158 & ~n9161;
  assign n9163 = ~n5192 & n9162;
  assign n9164 = n5192 & ~n9162;
  assign n9165 = ~n9163 & ~n9164;
  assign n9166 = ~n5077 & n9165;
  assign n9167 = ~n5305 & ~n9165;
  assign n9168 = ~n9166 & ~n9167;
  assign n9169 = ~n9068 & n9168;
  assign n9170 = n9068 & ~n9168;
  assign po149 = ~n9169 & ~n9170;
  assign n9172 = ~pi187 & pi439;
  assign n9173 = pi187 & ~pi439;
  assign po150 = n9172 | n9173;
  assign n9175 = ~pi255 & pi505;
  assign n9176 = pi255 & ~pi505;
  assign n9177 = ~n9175 & ~n9176;
  assign n9178 = pi529 & ~n9177;
  assign n9179 = n4957 & ~n9054;
  assign n9180 = ~n4957 & n9054;
  assign n9181 = ~n9179 & ~n9180;
  assign n9182 = n5298 & n8945;
  assign n9183 = ~n5298 & ~n8945;
  assign n9184 = ~n9182 & ~n9183;
  assign n9185 = n9181 & n9184;
  assign n9186 = ~n9181 & ~n9184;
  assign n9187 = ~n9185 & ~n9186;
  assign n9188 = ~pi090 & n4312;
  assign n9189 = ~n8451 & ~n8611;
  assign n9190 = ~pi019 & n4359;
  assign n9191 = ~n8427 & ~n9190;
  assign n9192 = ~n4360 & n9191;
  assign n9193 = ~pi090 & ~n9192;
  assign n9194 = n8324 & n8401;
  assign n9195 = ~n9193 & ~n9194;
  assign n9196 = n9189 & n9195;
  assign n9197 = pi088 & ~n9196;
  assign n9198 = pi090 & n4315;
  assign n9199 = pi019 & n4344;
  assign n9200 = ~n8403 & ~n9199;
  assign n9201 = ~pi090 & n4376;
  assign n9202 = n9200 & ~n9201;
  assign n9203 = ~n9198 & n9202;
  assign n9204 = ~pi088 & ~n9203;
  assign n9205 = ~n8474 & ~n9204;
  assign n9206 = ~pi019 & n8314;
  assign n9207 = ~n8362 & ~n9206;
  assign n9208 = pi090 & ~n9207;
  assign n9209 = n9205 & ~n9208;
  assign n9210 = ~n9197 & n9209;
  assign n9211 = ~n9188 & n9210;
  assign n9212 = ~pi006 & ~n9211;
  assign n9213 = pi090 & n8332;
  assign n9214 = n4287 & n4322;
  assign n9215 = ~n8344 & ~n9214;
  assign n9216 = n4297 & n8363;
  assign n9217 = ~n4383 & ~n4425;
  assign n9218 = pi019 & ~n9217;
  assign n9219 = ~n8603 & ~n9218;
  assign n9220 = ~n9216 & n9219;
  assign n9221 = ~pi090 & ~n9220;
  assign n9222 = pi019 & n8427;
  assign n9223 = ~n9221 & ~n9222;
  assign n9224 = n9215 & n9223;
  assign n9225 = ~n9213 & n9224;
  assign n9226 = pi088 & ~n9225;
  assign n9227 = ~n9212 & ~n9226;
  assign n9228 = ~n8412 & ~n8474;
  assign n9229 = ~n4293 & ~n4392;
  assign n9230 = ~n8331 & n9229;
  assign n9231 = ~n4330 & n9230;
  assign n9232 = ~n8473 & n9231;
  assign n9233 = pi090 & ~n9232;
  assign n9234 = ~pi019 & n4384;
  assign n9235 = ~n4357 & ~n9234;
  assign n9236 = ~n4365 & n9235;
  assign n9237 = ~pi090 & ~n9236;
  assign n9238 = ~n9233 & ~n9237;
  assign n9239 = n9228 & n9238;
  assign n9240 = ~pi088 & ~n9239;
  assign n9241 = ~pi090 & n8430;
  assign n9242 = n4315 & n4322;
  assign n9243 = ~n9241 & ~n9242;
  assign n9244 = ~n4393 & ~n8355;
  assign n9245 = ~pi090 & ~n9244;
  assign n9246 = ~n4299 & ~n8486;
  assign n9247 = ~n8449 & n9246;
  assign n9248 = ~n9245 & n9247;
  assign n9249 = pi088 & ~n9248;
  assign n9250 = pi019 & n4301;
  assign n9251 = ~pi090 & n4302;
  assign n9252 = ~n9250 & ~n9251;
  assign n9253 = n4286 & n4290;
  assign n9254 = ~pi090 & n9253;
  assign n9255 = ~n8457 & ~n9254;
  assign n9256 = ~n8539 & n9255;
  assign n9257 = n9252 & n9256;
  assign n9258 = ~pi088 & ~n9257;
  assign n9259 = ~n9249 & ~n9258;
  assign n9260 = ~pi051 & n8304;
  assign n9261 = ~pi049 & n8394;
  assign n9262 = ~n8602 & ~n9261;
  assign n9263 = ~n4356 & n9262;
  assign n9264 = ~n9260 & n9263;
  assign n9265 = pi090 & ~n9264;
  assign n9266 = ~n4394 & ~n9216;
  assign n9267 = ~n4371 & n9266;
  assign n9268 = ~pi090 & ~n9267;
  assign n9269 = ~n9265 & ~n9268;
  assign n9270 = n9259 & n9269;
  assign n9271 = pi006 & ~n9270;
  assign n9272 = n9243 & ~n9271;
  assign n9273 = ~n9240 & n9272;
  assign n9274 = n9227 & n9273;
  assign n9275 = ~pi255 & ~n9274;
  assign n9276 = pi255 & n9274;
  assign n9277 = ~n9275 & ~n9276;
  assign n9278 = ~n4687 & ~n4689;
  assign n9279 = pi066 & ~n9278;
  assign n9280 = ~n8885 & ~n9279;
  assign n9281 = ~n5165 & n9280;
  assign n9282 = ~pi118 & ~n9281;
  assign n9283 = ~n5123 & ~n9282;
  assign n9284 = ~n5211 & n9283;
  assign n9285 = pi034 & ~n9284;
  assign n9286 = ~n4648 & ~n5080;
  assign n9287 = ~n4773 & ~n5279;
  assign n9288 = ~n4725 & n9287;
  assign n9289 = n9286 & n9288;
  assign n9290 = pi118 & ~n9289;
  assign n9291 = ~pi066 & n4688;
  assign n9292 = ~n4705 & ~n9291;
  assign n9293 = ~n4657 & n9292;
  assign n9294 = ~pi118 & ~n9293;
  assign n9295 = ~n5240 & ~n9294;
  assign n9296 = ~n9290 & n9295;
  assign n9297 = ~n5178 & n9296;
  assign n9298 = ~pi034 & ~n9297;
  assign n9299 = ~pi066 & n5256;
  assign n9300 = ~n5208 & ~n9299;
  assign n9301 = pi118 & ~n9300;
  assign n9302 = ~n4706 & ~n5122;
  assign n9303 = ~pi066 & n4660;
  assign n9304 = n9302 & ~n9303;
  assign n9305 = ~pi118 & ~n9304;
  assign n9306 = ~n8855 & ~n8909;
  assign n9307 = n5225 & n5249;
  assign n9308 = n9306 & ~n9307;
  assign n9309 = ~n9305 & n9308;
  assign n9310 = pi034 & ~n9309;
  assign n9311 = ~pi118 & n4676;
  assign n9312 = pi066 & n4623;
  assign n9313 = ~n5227 & ~n9312;
  assign n9314 = pi118 & n4764;
  assign n9315 = n9313 & ~n9314;
  assign n9316 = ~n9311 & n9315;
  assign n9317 = ~pi034 & ~n9316;
  assign n9318 = ~pi118 & n4685;
  assign n9319 = ~n9317 & ~n9318;
  assign n9320 = ~n9310 & n9319;
  assign n9321 = ~n9301 & n9320;
  assign n9322 = ~n5178 & n9321;
  assign n9323 = ~pi038 & ~n9322;
  assign n9324 = pi118 & n5181;
  assign n9325 = pi101 & n4753;
  assign n9326 = n4622 & n9325;
  assign n9327 = ~n9324 & ~n9326;
  assign n9328 = pi034 & ~n9327;
  assign n9329 = ~n9323 & ~n9328;
  assign n9330 = ~n9298 & n9329;
  assign n9331 = ~n9285 & n9330;
  assign n9332 = pi118 & n4763;
  assign n9333 = n4668 & n9332;
  assign n9334 = n4667 & n8896;
  assign n9335 = ~n9333 & ~n9334;
  assign n9336 = ~pi062 & n5103;
  assign n9337 = ~n5169 & ~n9336;
  assign n9338 = pi118 & ~n9337;
  assign n9339 = ~pi118 & n4639;
  assign n9340 = pi066 & n4638;
  assign n9341 = ~n5111 & ~n9340;
  assign n9342 = ~n8935 & n9341;
  assign n9343 = ~n9339 & n9342;
  assign n9344 = ~n8927 & n9343;
  assign n9345 = ~pi034 & ~n9344;
  assign n9346 = pi118 & n5140;
  assign n9347 = ~n4647 & ~n4723;
  assign n9348 = ~pi118 & ~n9347;
  assign n9349 = ~n9346 & ~n9348;
  assign n9350 = ~n4644 & n9349;
  assign n9351 = ~n5164 & n9350;
  assign n9352 = pi034 & ~n9351;
  assign n9353 = ~n9345 & ~n9352;
  assign n9354 = ~pi066 & ~pi119;
  assign n9355 = pi103 & n9354;
  assign n9356 = ~n4704 & ~n9355;
  assign n9357 = pi118 & ~n9356;
  assign n9358 = ~n4715 & ~n4724;
  assign n9359 = ~n5165 & n9358;
  assign n9360 = ~pi118 & ~n9359;
  assign n9361 = ~n9357 & ~n9360;
  assign n9362 = n9353 & n9361;
  assign n9363 = ~n9338 & n9362;
  assign n9364 = pi038 & ~n9363;
  assign n9365 = n9335 & ~n9364;
  assign n9366 = n9331 & n9365;
  assign n9367 = pi116 & n8682;
  assign n9368 = ~n4558 & ~n4602;
  assign n9369 = pi011 & ~n9368;
  assign n9370 = ~pi011 & n4525;
  assign n9371 = ~n9369 & ~n9370;
  assign n9372 = ~n9154 & n9371;
  assign n9373 = ~pi116 & ~n9372;
  assign n9374 = pi116 & n8642;
  assign n9375 = ~n8653 & ~n9374;
  assign n9376 = ~n9133 & n9375;
  assign n9377 = ~n9373 & n9376;
  assign n9378 = ~n9367 & n9377;
  assign n9379 = pi058 & ~n9378;
  assign n9380 = ~n4548 & ~n9154;
  assign n9381 = ~n4532 & n9380;
  assign n9382 = ~pi116 & ~n9381;
  assign n9383 = ~pi116 & n4468;
  assign n9384 = ~n8780 & ~n9383;
  assign n9385 = pi000 & pi116;
  assign n9386 = pi022 & n9385;
  assign n9387 = n4459 & n9386;
  assign n9388 = pi011 & n4467;
  assign n9389 = ~n9070 & ~n9388;
  assign n9390 = ~n9387 & n9389;
  assign n9391 = n9384 & n9390;
  assign n9392 = ~pi058 & ~n9391;
  assign n9393 = ~pi000 & n8723;
  assign n9394 = ~pi011 & ~pi097;
  assign n9395 = pi000 & n9394;
  assign n9396 = ~n4525 & ~n9395;
  assign n9397 = ~n9149 & n9396;
  assign n9398 = ~n9393 & n9397;
  assign n9399 = pi116 & ~n9398;
  assign n9400 = ~n4461 & ~n4547;
  assign n9401 = ~pi116 & ~n9400;
  assign n9402 = ~n4473 & ~n8801;
  assign n9403 = ~n8774 & n9402;
  assign n9404 = ~n9401 & n9403;
  assign n9405 = pi058 & ~n9404;
  assign n9406 = ~n9399 & ~n9405;
  assign n9407 = ~n9392 & n9406;
  assign n9408 = ~n9382 & n9407;
  assign n9409 = pi060 & ~n9408;
  assign n9410 = ~pi116 & n8812;
  assign n9411 = n4481 & n4504;
  assign n9412 = ~n9410 & ~n9411;
  assign n9413 = ~pi011 & n4559;
  assign n9414 = ~n4526 & ~n9413;
  assign n9415 = ~n4535 & n9414;
  assign n9416 = ~pi116 & ~n9415;
  assign n9417 = ~n4462 & ~n8765;
  assign n9418 = ~n4489 & ~n8696;
  assign n9419 = ~n4549 & n9418;
  assign n9420 = n9417 & n9419;
  assign n9421 = pi116 & ~n9420;
  assign n9422 = ~n8716 & ~n8766;
  assign n9423 = ~n9421 & n9422;
  assign n9424 = ~n9416 & n9423;
  assign n9425 = ~pi058 & ~n9424;
  assign n9426 = n9412 & ~n9425;
  assign n9427 = ~pi116 & n4501;
  assign n9428 = ~pi011 & n4527;
  assign n9429 = ~n8824 & ~n9428;
  assign n9430 = ~n4528 & n9429;
  assign n9431 = ~pi116 & ~n9430;
  assign n9432 = pi011 & n8681;
  assign n9433 = ~n8771 & ~n9432;
  assign n9434 = n4540 & n8738;
  assign n9435 = n9433 & ~n9434;
  assign n9436 = ~n9431 & n9435;
  assign n9437 = pi058 & ~n9436;
  assign n9438 = pi011 & n8753;
  assign n9439 = ~n8740 & ~n9438;
  assign n9440 = pi116 & n4504;
  assign n9441 = ~pi116 & n4594;
  assign n9442 = ~n9440 & ~n9441;
  assign n9443 = n9439 & n9442;
  assign n9444 = ~pi058 & ~n9443;
  assign n9445 = ~pi011 & n8670;
  assign n9446 = ~n8649 & ~n9445;
  assign n9447 = pi116 & ~n9446;
  assign n9448 = ~n9444 & ~n9447;
  assign n9449 = ~n9437 & n9448;
  assign n9450 = ~n9427 & n9449;
  assign n9451 = ~n8766 & n9450;
  assign n9452 = ~pi060 & ~n9451;
  assign n9453 = n9426 & ~n9452;
  assign n9454 = ~n9409 & n9453;
  assign n9455 = ~n9379 & n9454;
  assign n9456 = n9366 & n9455;
  assign n9457 = ~n9366 & ~n9455;
  assign n9458 = ~n9456 & ~n9457;
  assign n9459 = ~n9277 & n9458;
  assign n9460 = n9277 & ~n9458;
  assign n9461 = ~n9459 & ~n9460;
  assign n9462 = ~n9187 & n9461;
  assign n9463 = n9187 & ~n9461;
  assign n9464 = ~n9462 & ~n9463;
  assign n9465 = ~pi529 & n9464;
  assign po151 = n9178 | n9465;
  assign n9467 = pi189 & pi496;
  assign n9468 = ~pi189 & ~pi496;
  assign n9469 = ~n9467 & ~n9468;
  assign n9470 = pi529 & n9469;
  assign n9471 = ~pi090 & n8379;
  assign n9472 = ~pi019 & n4367;
  assign n9473 = pi090 & n9472;
  assign n9474 = ~n8486 & ~n8561;
  assign n9475 = ~n9473 & n9474;
  assign n9476 = ~n9471 & n9475;
  assign n9477 = ~n9216 & n9476;
  assign n9478 = pi088 & ~n9477;
  assign n9479 = pi090 & n8364;
  assign n9480 = ~n9478 & ~n9479;
  assign n9481 = ~n4381 & ~n8463;
  assign n9482 = ~pi019 & n4295;
  assign n9483 = ~n8332 & ~n9482;
  assign n9484 = ~n8474 & n9483;
  assign n9485 = ~pi090 & ~n9484;
  assign n9486 = ~n8473 & ~n8569;
  assign n9487 = pi090 & ~n9486;
  assign n9488 = ~n9485 & ~n9487;
  assign n9489 = n9481 & n9488;
  assign n9490 = ~pi088 & ~n9489;
  assign n9491 = n9480 & ~n9490;
  assign n9492 = ~n4348 & ~n8305;
  assign n9493 = ~pi090 & ~n9492;
  assign n9494 = ~pi090 & n4314;
  assign n9495 = ~n4367 & ~n9494;
  assign n9496 = ~n8548 & n9495;
  assign n9497 = pi088 & ~n9496;
  assign n9498 = ~n8427 & ~n8576;
  assign n9499 = ~n4289 & ~n4303;
  assign n9500 = n9498 & n9499;
  assign n9501 = pi090 & ~n9500;
  assign n9502 = pi019 & n4405;
  assign n9503 = ~n8494 & ~n9502;
  assign n9504 = ~pi090 & ~n9503;
  assign n9505 = ~n4376 & ~n9504;
  assign n9506 = ~n9501 & n9505;
  assign n9507 = ~n9497 & n9506;
  assign n9508 = ~n9493 & n9507;
  assign n9509 = n8345 & n8355;
  assign n9510 = ~n4311 & ~n4404;
  assign n9511 = ~n8306 & n9510;
  assign n9512 = pi090 & ~n9511;
  assign n9513 = ~n9509 & ~n9512;
  assign n9514 = pi019 & n8448;
  assign n9515 = pi019 & n4415;
  assign n9516 = ~n8373 & ~n9515;
  assign n9517 = ~n9514 & n9516;
  assign n9518 = n9513 & n9517;
  assign n9519 = ~pi088 & ~n9518;
  assign n9520 = ~n9222 & ~n9519;
  assign n9521 = n9508 & n9520;
  assign n9522 = pi006 & ~n9521;
  assign n9523 = n9491 & ~n9522;
  assign n9524 = pi019 & pi112;
  assign n9525 = pi049 & pi051;
  assign n9526 = n9524 & n9525;
  assign n9527 = ~pi090 & n9526;
  assign n9528 = ~pi019 & n4301;
  assign n9529 = ~n4359 & ~n9528;
  assign n9530 = n4343 & ~n9529;
  assign n9531 = ~n4287 & ~n4383;
  assign n9532 = n8461 & ~n9531;
  assign n9533 = pi090 & n9532;
  assign n9534 = n4387 & n8363;
  assign n9535 = ~n8574 & ~n9534;
  assign n9536 = ~pi090 & ~n9535;
  assign n9537 = ~n9533 & ~n9536;
  assign n9538 = ~n4362 & n9537;
  assign n9539 = ~pi019 & ~n8382;
  assign n9540 = ~n9254 & ~n9539;
  assign n9541 = ~pi088 & ~n9540;
  assign n9542 = n4425 & n8345;
  assign n9543 = pi090 & n4392;
  assign n9544 = ~n4344 & ~n8337;
  assign n9545 = ~n9526 & n9544;
  assign n9546 = ~n9543 & n9545;
  assign n9547 = ~n9542 & n9546;
  assign n9548 = pi088 & ~n9547;
  assign n9549 = ~n9541 & ~n9548;
  assign n9550 = n9538 & n9549;
  assign n9551 = ~n9530 & n9550;
  assign n9552 = ~pi006 & ~n9551;
  assign n9553 = ~n9527 & ~n9552;
  assign n9554 = n9523 & n9553;
  assign n9555 = ~pi189 & ~n9554;
  assign n9556 = pi189 & n9554;
  assign n9557 = ~n9555 & ~n9556;
  assign n9558 = ~n8748 & n9162;
  assign n9559 = n8748 & ~n9162;
  assign n9560 = ~n9558 & ~n9559;
  assign n9561 = ~n5074 & n5298;
  assign n9562 = n5074 & ~n5298;
  assign n9563 = ~n9561 & ~n9562;
  assign n9564 = ~n9560 & n9563;
  assign n9565 = n9560 & ~n9563;
  assign n9566 = ~n9564 & ~n9565;
  assign n9567 = n9557 & n9566;
  assign n9568 = ~n9557 & ~n9566;
  assign n9569 = ~n9567 & ~n9568;
  assign n9570 = ~pi529 & n9569;
  assign po152 = n9470 | n9570;
  assign n9572 = pi139 & pi418;
  assign n9573 = ~pi139 & ~pi418;
  assign n9574 = ~n9572 & ~n9573;
  assign n9575 = pi529 & n9574;
  assign n9576 = pi009 & n6814;
  assign n9577 = ~n6811 & ~n9576;
  assign n9578 = ~n6666 & n9577;
  assign n9579 = ~n5930 & n9578;
  assign n9580 = pi113 & ~n9579;
  assign n9581 = n5966 & n6004;
  assign n9582 = ~pi009 & n5916;
  assign n9583 = ~n5925 & ~n6046;
  assign n9584 = ~n9582 & n9583;
  assign n9585 = pi113 & ~n9584;
  assign n9586 = ~n9581 & ~n9585;
  assign n9587 = pi009 & n6007;
  assign n9588 = ~pi025 & n5989;
  assign n9589 = ~n6802 & ~n9588;
  assign n9590 = ~n9587 & n9589;
  assign n9591 = n9586 & n9590;
  assign n9592 = ~pi096 & ~n9591;
  assign n9593 = ~pi009 & n5954;
  assign n9594 = pi009 & n5906;
  assign n9595 = ~pi124 & n5989;
  assign n9596 = ~n9594 & ~n9595;
  assign n9597 = ~pi113 & ~n9596;
  assign n9598 = ~n6722 & ~n6875;
  assign n9599 = ~pi113 & ~n9598;
  assign n9600 = ~n9597 & ~n9599;
  assign n9601 = ~n9593 & n9600;
  assign n9602 = ~pi113 & n5936;
  assign n9603 = ~n6702 & ~n9602;
  assign n9604 = ~n6770 & n9603;
  assign n9605 = pi096 & ~n9604;
  assign n9606 = n9601 & ~n9605;
  assign n9607 = ~n9592 & n9606;
  assign n9608 = ~n9580 & n9607;
  assign n9609 = ~n5931 & n9608;
  assign n9610 = ~pi010 & ~n9609;
  assign n9611 = n5910 & n5978;
  assign n9612 = ~pi113 & n9611;
  assign n9613 = ~n9610 & ~n9612;
  assign n9614 = pi113 & n5917;
  assign n9615 = ~pi124 & n9614;
  assign n9616 = n5936 & n9615;
  assign n9617 = ~n5904 & ~n5965;
  assign n9618 = ~pi009 & n5940;
  assign n9619 = n9617 & ~n9618;
  assign n9620 = ~pi113 & ~n9619;
  assign n9621 = ~pi113 & n6672;
  assign n9622 = pi113 & n9576;
  assign n9623 = ~n9621 & ~n9622;
  assign n9624 = n5917 & n5929;
  assign n9625 = ~n6692 & ~n9624;
  assign n9626 = pi113 & ~n9625;
  assign n9627 = n9623 & ~n9626;
  assign n9628 = ~n9620 & n9627;
  assign n9629 = ~pi096 & ~n9628;
  assign n9630 = ~pi113 & n6709;
  assign n9631 = ~pi009 & n6770;
  assign n9632 = pi113 & n9631;
  assign n9633 = ~n6001 & ~n6684;
  assign n9634 = ~n9632 & n9633;
  assign n9635 = ~n9630 & n9634;
  assign n9636 = ~n5918 & n9635;
  assign n9637 = pi096 & ~n9636;
  assign n9638 = ~n9629 & ~n9637;
  assign n9639 = n5907 & n5966;
  assign n9640 = pi113 & n6041;
  assign n9641 = ~n9611 & ~n9640;
  assign n9642 = ~n9639 & n9641;
  assign n9643 = ~n5969 & ~n6894;
  assign n9644 = n9642 & n9643;
  assign n9645 = pi096 & ~n9644;
  assign n9646 = ~pi009 & ~n6856;
  assign n9647 = ~n6018 & ~n9646;
  assign n9648 = ~pi096 & ~n9647;
  assign n9649 = n5917 & n6756;
  assign n9650 = ~n6665 & ~n9649;
  assign n9651 = ~pi113 & ~n9650;
  assign n9652 = n5951 & n5966;
  assign n9653 = ~n9651 & ~n9652;
  assign n9654 = pi113 & ~pi125;
  assign n9655 = ~n5906 & ~n5921;
  assign n9656 = n9654 & ~n9655;
  assign n9657 = pi009 & n9656;
  assign n9658 = n9653 & ~n9657;
  assign n9659 = ~pi009 & n6012;
  assign n9660 = ~n5948 & ~n9659;
  assign n9661 = n6852 & ~n9660;
  assign n9662 = n9658 & ~n9661;
  assign n9663 = ~n9648 & n9662;
  assign n9664 = ~n9645 & n9663;
  assign n9665 = pi010 & ~n9664;
  assign n9666 = n9638 & ~n9665;
  assign n9667 = ~n9616 & n9666;
  assign n9668 = n9613 & n9667;
  assign n9669 = ~pi139 & ~n9668;
  assign n9670 = pi139 & n9668;
  assign n9671 = ~n9669 & ~n9670;
  assign n9672 = n5484 & ~n5772;
  assign n9673 = ~n5484 & n5772;
  assign n9674 = ~n9672 & ~n9673;
  assign n9675 = ~n7195 & n9674;
  assign n9676 = ~n7193 & ~n9674;
  assign n9677 = ~n7194 & n9676;
  assign n9678 = ~n9675 & ~n9677;
  assign n9679 = n9671 & n9678;
  assign n9680 = ~n9671 & ~n9678;
  assign n9681 = ~n9679 & ~n9680;
  assign n9682 = ~pi529 & n9681;
  assign po153 = n9575 | n9682;
  assign n9684 = ~pi182 & pi436;
  assign n9685 = pi182 & ~pi436;
  assign n9686 = ~n9684 & ~n9685;
  assign n9687 = pi529 & ~n9686;
  assign n9688 = ~pi182 & ~n6906;
  assign n9689 = pi182 & n6906;
  assign n9690 = ~n9688 & ~n9689;
  assign n9691 = pi113 & n5926;
  assign n9692 = pi009 & n5910;
  assign n9693 = ~n9594 & ~n9692;
  assign n9694 = ~n6718 & n9693;
  assign n9695 = ~pi113 & ~n9694;
  assign n9696 = ~n6825 & ~n9695;
  assign n9697 = ~n6026 & ~n6894;
  assign n9698 = pi113 & ~n9697;
  assign n9699 = n9696 & ~n9698;
  assign n9700 = pi096 & ~n9699;
  assign n9701 = ~pi113 & n6001;
  assign n9702 = ~n5951 & ~n9701;
  assign n9703 = n6681 & n6685;
  assign n9704 = ~n6709 & ~n9703;
  assign n9705 = ~pi096 & ~n9704;
  assign n9706 = n9702 & ~n9705;
  assign n9707 = ~n9700 & n9706;
  assign n9708 = ~n9691 & n9707;
  assign n9709 = pi010 & ~n9708;
  assign n9710 = ~n5907 & ~n5921;
  assign n9711 = ~pi009 & n9654;
  assign n9712 = ~n9710 & n9711;
  assign n9713 = ~n6762 & ~n9712;
  assign n9714 = ~n9709 & n9713;
  assign n9715 = n5954 & n5958;
  assign n9716 = ~n9624 & ~n9715;
  assign n9717 = pi113 & ~n5969;
  assign n9718 = pi055 & n5994;
  assign n9719 = ~n6757 & ~n9718;
  assign n9720 = ~pi113 & n9719;
  assign n9721 = ~n9717 & ~n9720;
  assign n9722 = ~n9621 & ~n9721;
  assign n9723 = pi096 & ~n9722;
  assign n9724 = ~pi113 & n6691;
  assign n9725 = pi113 & n6706;
  assign n9726 = ~n5955 & ~n9725;
  assign n9727 = ~n6008 & n9726;
  assign n9728 = ~n5946 & ~n6016;
  assign n9729 = n9727 & n9728;
  assign n9730 = ~n9724 & n9729;
  assign n9731 = ~n6035 & ~n6802;
  assign n9732 = n9730 & n9731;
  assign n9733 = ~pi096 & ~n9732;
  assign n9734 = ~n6770 & ~n6814;
  assign n9735 = ~n5911 & n9734;
  assign n9736 = n5938 & ~n9735;
  assign n9737 = ~n5965 & ~n9736;
  assign n9738 = ~n9733 & n9737;
  assign n9739 = ~n9723 & n9738;
  assign n9740 = n9716 & n9739;
  assign n9741 = ~pi010 & ~n9740;
  assign n9742 = n9714 & ~n9741;
  assign n9743 = pi009 & n6757;
  assign n9744 = pi009 & n6756;
  assign n9745 = ~n6051 & ~n9744;
  assign n9746 = ~n6709 & n9745;
  assign n9747 = pi113 & ~n9746;
  assign n9748 = ~n5964 & ~n6047;
  assign n9749 = ~n6674 & n9748;
  assign n9750 = ~pi113 & ~n9749;
  assign n9751 = n5921 & n5966;
  assign n9752 = ~n9750 & ~n9751;
  assign n9753 = ~n9747 & n9752;
  assign n9754 = ~n9743 & n9753;
  assign n9755 = ~n5930 & n9754;
  assign n9756 = ~pi096 & ~n9755;
  assign n9757 = ~pi113 & n6732;
  assign n9758 = n5928 & n5994;
  assign n9759 = ~n6766 & ~n9758;
  assign n9760 = ~pi113 & ~n9759;
  assign n9761 = pi113 & n5942;
  assign n9762 = ~n6053 & ~n9761;
  assign n9763 = ~n9760 & n9762;
  assign n9764 = ~n9757 & n9763;
  assign n9765 = pi124 & n5917;
  assign n9766 = ~n5925 & ~n9765;
  assign n9767 = pi113 & ~n9766;
  assign n9768 = n9764 & ~n9767;
  assign n9769 = pi096 & ~n9768;
  assign n9770 = ~n9756 & ~n9769;
  assign n9771 = n9742 & n9770;
  assign n9772 = ~n6659 & n9771;
  assign n9773 = n6659 & ~n9771;
  assign n9774 = ~n9772 & ~n9773;
  assign n9775 = ~n9690 & n9774;
  assign n9776 = n9690 & ~n9774;
  assign n9777 = ~n9775 & ~n9776;
  assign n9778 = ~n5823 & n5894;
  assign n9779 = ~n5861 & n9778;
  assign n9780 = n5603 & ~n9779;
  assign n9781 = ~n5603 & n9779;
  assign n9782 = ~n9780 & ~n9781;
  assign n9783 = n6536 & n9782;
  assign n9784 = ~n6536 & ~n9782;
  assign n9785 = ~n9783 & ~n9784;
  assign n9786 = ~n9777 & n9785;
  assign n9787 = n9777 & ~n9785;
  assign n9788 = ~n9786 & ~n9787;
  assign n9789 = ~pi529 & n9788;
  assign po154 = n9687 | n9789;
  assign n9791 = pi193 & pi475;
  assign n9792 = ~pi193 & ~pi475;
  assign n9793 = ~n9791 & ~n9792;
  assign n9794 = pi529 & n9793;
  assign n9795 = ~pi193 & ~n9668;
  assign n9796 = pi193 & n9668;
  assign n9797 = ~n9795 & ~n9796;
  assign n9798 = n5484 & ~n7001;
  assign n9799 = ~n5484 & n7001;
  assign n9800 = ~n9798 & ~n9799;
  assign n9801 = ~n6301 & ~n6543;
  assign n9802 = ~n6193 & ~n6263;
  assign n9803 = ~n6250 & n9802;
  assign n9804 = ~pi035 & ~n9803;
  assign n9805 = n9801 & ~n9804;
  assign n9806 = pi106 & ~n9805;
  assign n9807 = pi031 & n6293;
  assign n9808 = n7013 & ~n9807;
  assign n9809 = pi035 & ~n9808;
  assign n9810 = ~n6237 & ~n9809;
  assign n9811 = ~pi106 & ~n9810;
  assign n9812 = ~n9806 & ~n9811;
  assign n9813 = pi065 & ~n9812;
  assign n9814 = pi031 & n6277;
  assign n9815 = ~n6562 & ~n9814;
  assign n9816 = ~pi106 & ~n9815;
  assign n9817 = pi035 & n6170;
  assign n9818 = n6184 & n6312;
  assign n9819 = ~n9817 & ~n9818;
  assign n9820 = ~n9816 & n9819;
  assign n9821 = ~n6167 & n9820;
  assign n9822 = pi065 & ~pi068;
  assign n9823 = ~n9821 & n9822;
  assign n9824 = pi035 & n6197;
  assign n9825 = ~pi035 & n6203;
  assign n9826 = ~n6221 & ~n9825;
  assign n9827 = ~n9824 & n9826;
  assign n9828 = n7009 & ~n9827;
  assign n9829 = ~n6213 & ~n7075;
  assign n9830 = ~pi106 & ~n9829;
  assign n9831 = ~n6227 & ~n7055;
  assign n9832 = ~pi106 & ~n9831;
  assign n9833 = pi035 & n6554;
  assign n9834 = ~pi106 & n9833;
  assign n9835 = ~n9832 & ~n9834;
  assign n9836 = ~n6585 & n9835;
  assign n9837 = ~pi065 & ~n9836;
  assign n9838 = ~n9830 & ~n9837;
  assign n9839 = ~n9828 & n9838;
  assign n9840 = n6186 & n6320;
  assign n9841 = ~n6198 & ~n9840;
  assign n9842 = ~pi065 & ~n9841;
  assign n9843 = ~n6212 & ~n6308;
  assign n9844 = ~pi106 & ~n9843;
  assign n9845 = ~n9832 & ~n9844;
  assign n9846 = ~pi106 & pi128;
  assign n9847 = ~pi031 & n9846;
  assign n9848 = ~n7041 & ~n9847;
  assign n9849 = ~pi065 & ~n9848;
  assign n9850 = ~n6605 & ~n7039;
  assign n9851 = n6320 & ~n9850;
  assign n9852 = ~pi031 & n6197;
  assign n9853 = n6320 & n9852;
  assign n9854 = ~n9851 & ~n9853;
  assign n9855 = ~n9849 & n9854;
  assign n9856 = n9845 & n9855;
  assign n9857 = ~n9842 & n9856;
  assign n9858 = ~pi068 & ~n9857;
  assign n9859 = n9839 & ~n9858;
  assign n9860 = ~pi035 & n6250;
  assign n9861 = ~pi035 & n9807;
  assign n9862 = ~n9860 & ~n9861;
  assign n9863 = ~n6307 & n9862;
  assign n9864 = pi106 & ~n9863;
  assign n9865 = ~n7035 & ~n9864;
  assign n9866 = n6210 & n6320;
  assign n9867 = pi035 & n6178;
  assign n9868 = ~pi031 & pi100;
  assign n9869 = ~n6648 & ~n9868;
  assign n9870 = ~n7020 & n9869;
  assign n9871 = ~n9867 & n9870;
  assign n9872 = pi065 & pi106;
  assign n9873 = ~n9871 & n9872;
  assign n9874 = ~n9866 & ~n9873;
  assign n9875 = n9865 & n9874;
  assign n9876 = n6172 & n6645;
  assign n9877 = ~n6221 & ~n9876;
  assign n9878 = pi065 & ~n9877;
  assign n9879 = ~pi106 & n6235;
  assign n9880 = ~n9878 & ~n9879;
  assign n9881 = n6184 & n6554;
  assign n9882 = ~n6181 & ~n6203;
  assign n9883 = ~n6648 & n9882;
  assign n9884 = ~pi106 & ~n9883;
  assign n9885 = ~pi106 & n6179;
  assign n9886 = ~n9884 & ~n9885;
  assign n9887 = ~n6579 & n9886;
  assign n9888 = ~n9881 & n9887;
  assign n9889 = ~n6235 & ~n6295;
  assign n9890 = n9888 & n9889;
  assign n9891 = ~pi065 & ~n9890;
  assign n9892 = n9880 & ~n9891;
  assign n9893 = n9875 & n9892;
  assign n9894 = pi068 & ~n9893;
  assign n9895 = n9859 & ~n9894;
  assign n9896 = ~n9823 & n9895;
  assign n9897 = ~n9813 & n9896;
  assign n9898 = ~n7102 & n9897;
  assign n9899 = n7102 & ~n9897;
  assign n9900 = ~n9898 & ~n9899;
  assign n9901 = ~n9800 & n9900;
  assign n9902 = n9800 & ~n9900;
  assign n9903 = ~n9901 & ~n9902;
  assign n9904 = n9797 & n9903;
  assign n9905 = ~n9797 & ~n9903;
  assign n9906 = ~n9904 & ~n9905;
  assign n9907 = ~pi529 & n9906;
  assign po155 = n9794 | n9907;
  assign n9909 = n2731 & ~n3092;
  assign n9910 = ~pi123 & ~n9909;
  assign n9911 = pi123 & n2698;
  assign n9912 = ~n7648 & ~n9911;
  assign n9913 = ~n3123 & n9912;
  assign n9914 = ~n9910 & n9913;
  assign n9915 = pi023 & n7255;
  assign n9916 = pi027 & pi111;
  assign n9917 = ~pi023 & n9916;
  assign n9918 = ~n2738 & ~n9917;
  assign n9919 = ~n9915 & n9918;
  assign n9920 = pi048 & ~n9919;
  assign n9921 = ~pi123 & n9920;
  assign n9922 = ~n2702 & ~n3090;
  assign n9923 = ~n2050 & ~n2766;
  assign n9924 = n9922 & n9923;
  assign n9925 = pi048 & ~n9924;
  assign n9926 = ~n9921 & ~n9925;
  assign n9927 = n9914 & n9926;
  assign n9928 = ~n2010 & ~n2698;
  assign n9929 = ~n1921 & ~n2036;
  assign n9930 = pi123 & ~n9929;
  assign n9931 = ~pi123 & n2031;
  assign n9932 = ~n9930 & ~n9931;
  assign n9933 = n9928 & n9932;
  assign n9934 = ~n3170 & n9933;
  assign n9935 = ~pi048 & ~n9934;
  assign n9936 = ~n7276 & ~n9935;
  assign n9937 = n9927 & n9936;
  assign n9938 = pi020 & ~n9937;
  assign n9939 = ~pi123 & n1932;
  assign n9940 = ~pi023 & ~pi123;
  assign n9941 = ~pi111 & n9940;
  assign n9942 = n1950 & n9941;
  assign n9943 = ~n9939 & ~n9942;
  assign n9944 = n1975 & n9915;
  assign n9945 = ~n1995 & ~n9944;
  assign n9946 = n9943 & n9945;
  assign n9947 = n1923 & n1943;
  assign n9948 = ~n1993 & ~n9947;
  assign n9949 = ~pi027 & n2005;
  assign n9950 = n1982 & n2738;
  assign n9951 = ~n9949 & ~n9950;
  assign n9952 = n9948 & n9951;
  assign n9953 = ~pi048 & ~n9952;
  assign n9954 = pi027 & n2741;
  assign n9955 = ~n1955 & ~n9954;
  assign n9956 = pi027 & n7256;
  assign n9957 = n1976 & n3079;
  assign n9958 = ~n9956 & ~n9957;
  assign n9959 = n9955 & n9958;
  assign n9960 = pi123 & ~n9959;
  assign n9961 = ~n2783 & ~n3197;
  assign n9962 = ~pi027 & n2056;
  assign n9963 = n9961 & ~n9962;
  assign n9964 = ~pi123 & ~n9963;
  assign n9965 = ~n2023 & ~n9954;
  assign n9966 = ~n2003 & ~n2039;
  assign n9967 = pi123 & ~n9966;
  assign n9968 = n9965 & ~n9967;
  assign n9969 = ~n9964 & n9968;
  assign n9970 = ~n2732 & ~n2781;
  assign n9971 = ~n3111 & n9970;
  assign n9972 = n9969 & n9971;
  assign n9973 = pi048 & ~n9972;
  assign n9974 = ~n9960 & ~n9973;
  assign n9975 = ~n9953 & n9974;
  assign n9976 = n9946 & n9975;
  assign n9977 = ~pi020 & ~n9976;
  assign n9978 = ~n9938 & ~n9977;
  assign n9979 = ~pi027 & n2041;
  assign n9980 = ~n2004 & ~n9979;
  assign n9981 = ~n1952 & n9980;
  assign n9982 = n7290 & ~n9981;
  assign n9983 = n1982 & n3196;
  assign n9984 = n3079 & ~n7237;
  assign n9985 = ~n2698 & ~n9984;
  assign n9986 = pi123 & ~n9985;
  assign n9987 = ~n9983 & ~n9986;
  assign n9988 = ~n2694 & n9987;
  assign n9989 = ~pi048 & ~n9988;
  assign n9990 = ~n2760 & ~n7680;
  assign n9991 = ~pi123 & n2023;
  assign n9992 = n9990 & ~n9991;
  assign n9993 = ~n9989 & n9992;
  assign n9994 = ~n9982 & n9993;
  assign n9995 = pi027 & n1995;
  assign n9996 = ~n9939 & ~n9995;
  assign n9997 = pi048 & ~n9996;
  assign n9998 = n2720 & n7254;
  assign n9999 = ~n9997 & ~n9998;
  assign n10000 = n9994 & n9999;
  assign n10001 = n9978 & n10000;
  assign n10002 = ~n1841 & ~n1891;
  assign n10003 = ~n2821 & n10002;
  assign n10004 = ~pi114 & ~n10003;
  assign n10005 = pi114 & n7378;
  assign n10006 = ~n7862 & ~n10005;
  assign n10007 = ~n7303 & n10006;
  assign n10008 = ~n10004 & n10007;
  assign n10009 = ~pi114 & n1881;
  assign n10010 = ~n1762 & ~n1902;
  assign n10011 = pi114 & ~n10010;
  assign n10012 = ~n1841 & ~n7378;
  assign n10013 = ~n2874 & n10012;
  assign n10014 = ~n10011 & n10013;
  assign n10015 = ~n10009 & n10014;
  assign n10016 = ~pi001 & ~n10015;
  assign n10017 = n10008 & ~n10016;
  assign n10018 = ~n1878 & ~n2961;
  assign n10019 = ~n2974 & ~n2989;
  assign n10020 = n10018 & n10019;
  assign n10021 = pi001 & ~n10020;
  assign n10022 = pi013 & pi054;
  assign n10023 = ~pi007 & n10022;
  assign n10024 = pi007 & n7382;
  assign n10025 = ~n10023 & ~n10024;
  assign n10026 = ~n2958 & n10025;
  assign n10027 = n1782 & ~n10026;
  assign n10028 = ~n7354 & ~n10027;
  assign n10029 = ~n10021 & n10028;
  assign n10030 = n10017 & n10029;
  assign n10031 = pi029 & ~n10030;
  assign n10032 = n2827 & n2860;
  assign n10033 = ~pi013 & n1897;
  assign n10034 = ~n1848 & ~n10033;
  assign n10035 = ~n1758 & n10034;
  assign n10036 = ~pi114 & ~n10035;
  assign n10037 = ~n10032 & ~n10036;
  assign n10038 = ~n7332 & n10037;
  assign n10039 = n1877 & ~n7314;
  assign n10040 = ~n7378 & ~n10039;
  assign n10041 = pi114 & ~n10040;
  assign n10042 = n10038 & ~n10041;
  assign n10043 = ~pi001 & ~n10042;
  assign n10044 = pi013 & n2828;
  assign n10045 = n1805 & n1847;
  assign n10046 = ~n10044 & ~n10045;
  assign n10047 = pi001 & ~n10046;
  assign n10048 = ~n1794 & ~n3014;
  assign n10049 = pi114 & ~n10048;
  assign n10050 = pi013 & n2910;
  assign n10051 = pi013 & n7383;
  assign n10052 = ~n10050 & ~n10051;
  assign n10053 = pi114 & ~n10052;
  assign n10054 = ~n10049 & ~n10053;
  assign n10055 = ~pi114 & n2922;
  assign n10056 = n7372 & n10024;
  assign n10057 = ~n2828 & ~n10056;
  assign n10058 = ~pi114 & n1778;
  assign n10059 = n10057 & ~n10058;
  assign n10060 = ~n10055 & n10059;
  assign n10061 = n10054 & n10060;
  assign n10062 = n1775 & n1877;
  assign n10063 = ~n1825 & ~n10062;
  assign n10064 = ~pi001 & ~n10063;
  assign n10065 = ~n2861 & ~n7316;
  assign n10066 = ~pi013 & n1871;
  assign n10067 = n10065 & ~n10066;
  assign n10068 = ~pi114 & ~n10067;
  assign n10069 = ~n1853 & ~n10050;
  assign n10070 = ~n1847 & ~n1904;
  assign n10071 = pi114 & ~n10070;
  assign n10072 = n10069 & ~n10071;
  assign n10073 = ~n10068 & n10072;
  assign n10074 = ~n2917 & ~n7344;
  assign n10075 = ~n2904 & n10074;
  assign n10076 = n10073 & n10075;
  assign n10077 = pi001 & ~n10076;
  assign n10078 = n2827 & n2958;
  assign n10079 = n1765 & n1805;
  assign n10080 = ~n10078 & ~n10079;
  assign n10081 = ~pi001 & ~n10080;
  assign n10082 = ~n10077 & ~n10081;
  assign n10083 = ~n10064 & n10082;
  assign n10084 = n10061 & n10083;
  assign n10085 = ~pi029 & ~n10084;
  assign n10086 = pi001 & n10058;
  assign n10087 = ~n10085 & ~n10086;
  assign n10088 = ~n10047 & n10087;
  assign n10089 = ~n10043 & n10088;
  assign n10090 = ~n10031 & n10089;
  assign n10091 = ~pi114 & n1853;
  assign n10092 = ~n3030 & ~n10091;
  assign n10093 = ~n7848 & n10092;
  assign n10094 = n10090 & n10093;
  assign n10095 = ~n10001 & ~n10094;
  assign n10096 = n10001 & n10094;
  assign n10097 = ~n10095 & ~n10096;
  assign n10098 = ~n2181 & ~n2425;
  assign n10099 = n2140 & n2159;
  assign n10100 = pi104 & n2462;
  assign n10101 = ~n10099 & ~n10100;
  assign n10102 = pi069 & n2412;
  assign n10103 = ~n2396 & ~n10102;
  assign n10104 = ~n2205 & n10103;
  assign n10105 = n2266 & ~n10104;
  assign n10106 = pi102 & n7793;
  assign n10107 = ~n10105 & ~n10106;
  assign n10108 = n10101 & n10107;
  assign n10109 = n10098 & n10108;
  assign n10110 = pi104 & n2139;
  assign n10111 = ~n2152 & ~n2352;
  assign n10112 = ~n2461 & n10111;
  assign n10113 = ~pi104 & ~n10112;
  assign n10114 = ~n2397 & ~n2440;
  assign n10115 = ~n2405 & n10114;
  assign n10116 = ~n10113 & n10115;
  assign n10117 = ~n10110 & n10116;
  assign n10118 = ~pi102 & ~n10117;
  assign n10119 = n10109 & ~n10118;
  assign n10120 = ~n2156 & ~n2412;
  assign n10121 = ~n2534 & n10120;
  assign n10122 = pi104 & ~n10121;
  assign n10123 = ~pi033 & pi127;
  assign n10124 = ~n2250 & ~n10123;
  assign n10125 = n2135 & ~n10124;
  assign n10126 = ~n2563 & ~n10125;
  assign n10127 = ~n2337 & n10126;
  assign n10128 = ~n10122 & n10127;
  assign n10129 = pi102 & ~n10128;
  assign n10130 = pi126 & n2106;
  assign n10131 = ~n2086 & ~n10130;
  assign n10132 = pi104 & ~n10131;
  assign n10133 = ~pi033 & n2335;
  assign n10134 = n2120 & n10133;
  assign n10135 = pi127 & n2415;
  assign n10136 = n2388 & n10135;
  assign n10137 = ~n7729 & ~n10136;
  assign n10138 = ~n2152 & n10137;
  assign n10139 = ~n10134 & n10138;
  assign n10140 = ~n10132 & n10139;
  assign n10141 = ~pi102 & ~n10140;
  assign n10142 = ~n10129 & ~n10141;
  assign n10143 = ~n2283 & ~n2372;
  assign n10144 = ~pi104 & ~n10143;
  assign n10145 = ~n2197 & ~n2437;
  assign n10146 = ~n2157 & ~n2568;
  assign n10147 = n10145 & n10146;
  assign n10148 = pi104 & ~n10147;
  assign n10149 = ~n10144 & ~n10148;
  assign n10150 = n10142 & n10149;
  assign n10151 = pi012 & ~n10150;
  assign n10152 = ~pi104 & n2568;
  assign n10153 = ~pi069 & n2416;
  assign n10154 = ~n2314 & ~n10153;
  assign n10155 = pi104 & ~n10154;
  assign n10156 = ~n10152 & ~n10155;
  assign n10157 = ~n2101 & n10156;
  assign n10158 = pi102 & ~n10157;
  assign n10159 = ~pi104 & n10130;
  assign n10160 = ~pi069 & n2210;
  assign n10161 = ~n10159 & ~n10160;
  assign n10162 = ~n2190 & ~n2305;
  assign n10163 = ~n2351 & ~n2372;
  assign n10164 = n10162 & n10163;
  assign n10165 = n10161 & n10164;
  assign n10166 = ~pi102 & ~n10165;
  assign n10167 = ~n10158 & ~n10166;
  assign n10168 = n2105 & n2250;
  assign n10169 = ~n2351 & ~n10168;
  assign n10170 = pi104 & ~n10169;
  assign n10171 = ~pi069 & n2251;
  assign n10172 = pi127 & n2511;
  assign n10173 = ~n2177 & n2195;
  assign n10174 = ~n10172 & ~n10173;
  assign n10175 = ~n2220 & n10174;
  assign n10176 = ~n10171 & n10175;
  assign n10177 = ~pi104 & ~n10176;
  assign n10178 = ~n10170 & ~n10177;
  assign n10179 = n10167 & n10178;
  assign n10180 = ~pi012 & ~n10179;
  assign n10181 = ~n10151 & ~n10180;
  assign n10182 = n10119 & n10181;
  assign n10183 = ~pi153 & ~n10182;
  assign n10184 = pi153 & n10182;
  assign n10185 = ~n10183 & ~n10184;
  assign n10186 = ~n1940 & ~n2781;
  assign n10187 = ~n2749 & n10186;
  assign n10188 = pi123 & ~n10187;
  assign n10189 = pi023 & ~pi111;
  assign n10190 = ~n2737 & ~n10189;
  assign n10191 = n3051 & ~n10190;
  assign n10192 = n3075 & ~n10191;
  assign n10193 = ~n10188 & n10192;
  assign n10194 = pi048 & ~n10193;
  assign n10195 = pi027 & pi093;
  assign n10196 = pi023 & n10195;
  assign n10197 = ~n1976 & ~n10196;
  assign n10198 = pi123 & ~n10197;
  assign n10199 = ~n1932 & ~n7636;
  assign n10200 = ~n9942 & n10199;
  assign n10201 = ~n9944 & n10200;
  assign n10202 = ~n10198 & n10201;
  assign n10203 = ~pi048 & ~n10202;
  assign n10204 = ~n10194 & ~n10203;
  assign n10205 = ~n2714 & ~n3197;
  assign n10206 = ~pi123 & ~n10205;
  assign n10207 = ~n2031 & ~n2698;
  assign n10208 = ~n1995 & n10207;
  assign n10209 = ~n1941 & n10208;
  assign n10210 = pi123 & ~n10209;
  assign n10211 = ~n10206 & ~n10210;
  assign n10212 = n10204 & n10211;
  assign n10213 = pi020 & ~n10212;
  assign n10214 = pi027 & n2781;
  assign n10215 = ~n2694 & ~n10214;
  assign n10216 = ~n1924 & n10215;
  assign n10217 = n2720 & ~n10216;
  assign n10218 = pi048 & n7680;
  assign n10219 = ~pi027 & n7256;
  assign n10220 = ~n3132 & ~n10219;
  assign n10221 = pi123 & ~n10220;
  assign n10222 = ~pi123 & n1995;
  assign n10223 = ~n2004 & ~n10222;
  assign n10224 = ~n10221 & n10223;
  assign n10225 = pi048 & ~n10224;
  assign n10226 = ~n1984 & ~n2714;
  assign n10227 = ~n1953 & n10226;
  assign n10228 = ~pi123 & n10196;
  assign n10229 = ~pi027 & n2054;
  assign n10230 = ~n10228 & ~n10229;
  assign n10231 = ~n3212 & n10230;
  assign n10232 = n10227 & n10231;
  assign n10233 = ~pi048 & ~n10232;
  assign n10234 = ~n10225 & ~n10233;
  assign n10235 = ~n1953 & ~n3066;
  assign n10236 = pi123 & ~n10235;
  assign n10237 = ~pi027 & n3177;
  assign n10238 = pi023 & n1962;
  assign n10239 = ~n10237 & ~n10238;
  assign n10240 = ~n1989 & n2032;
  assign n10241 = ~n2068 & ~n10240;
  assign n10242 = n10239 & n10241;
  assign n10243 = ~pi123 & ~n10242;
  assign n10244 = ~n10236 & ~n10243;
  assign n10245 = n10234 & n10244;
  assign n10246 = ~pi020 & ~n10245;
  assign n10247 = ~n10218 & ~n10246;
  assign n10248 = pi123 & n1956;
  assign n10249 = ~n1932 & ~n2776;
  assign n10250 = ~n2748 & n10249;
  assign n10251 = ~pi123 & ~n10250;
  assign n10252 = ~n3114 & ~n7266;
  assign n10253 = ~n2786 & n10252;
  assign n10254 = ~n10251 & n10253;
  assign n10255 = ~n10248 & n10254;
  assign n10256 = ~pi048 & ~n10255;
  assign n10257 = pi123 & n2752;
  assign n10258 = ~n10256 & ~n10257;
  assign n10259 = ~n1996 & ~n9947;
  assign n10260 = ~n7244 & n10259;
  assign n10261 = n10258 & n10260;
  assign n10262 = n10247 & n10261;
  assign n10263 = ~n10217 & n10262;
  assign n10264 = ~n10213 & n10263;
  assign n10265 = ~n1738 & ~n7449;
  assign n10266 = pi040 & n7531;
  assign n10267 = n10265 & ~n10266;
  assign n10268 = ~pi072 & pi107;
  assign n10269 = ~n1556 & ~n10268;
  assign n10270 = n1595 & ~n10269;
  assign n10271 = ~n1542 & ~n2590;
  assign n10272 = ~n10270 & n10271;
  assign n10273 = ~n1553 & ~n1699;
  assign n10274 = ~n2643 & n10273;
  assign n10275 = pi083 & ~n10274;
  assign n10276 = n10272 & ~n10275;
  assign n10277 = pi040 & ~n10276;
  assign n10278 = ~pi083 & n1614;
  assign n10279 = pi107 & n1717;
  assign n10280 = n1693 & n10279;
  assign n10281 = pi014 & pi108;
  assign n10282 = pi107 & n10281;
  assign n10283 = ~n1523 & ~n10282;
  assign n10284 = pi083 & ~n10283;
  assign n10285 = ~n1629 & ~n7566;
  assign n10286 = ~n10284 & n10285;
  assign n10287 = ~n10280 & n10286;
  assign n10288 = ~n10278 & n10287;
  assign n10289 = ~pi040 & ~n10288;
  assign n10290 = ~n10277 & ~n10289;
  assign n10291 = ~n1514 & ~n1731;
  assign n10292 = ~n1730 & n10291;
  assign n10293 = ~n1656 & n10292;
  assign n10294 = pi083 & ~n10293;
  assign n10295 = ~n1483 & ~n1580;
  assign n10296 = ~pi083 & ~n10295;
  assign n10297 = ~n10294 & ~n10296;
  assign n10298 = n10290 & n10297;
  assign n10299 = pi078 & ~n10298;
  assign n10300 = n10267 & ~n10299;
  assign n10301 = pi014 & n1699;
  assign n10302 = ~n1664 & ~n10301;
  assign n10303 = ~n1487 & n10302;
  assign n10304 = n1587 & ~n10303;
  assign n10305 = pi083 & n7427;
  assign n10306 = ~n1666 & ~n1728;
  assign n10307 = ~n1530 & ~n1629;
  assign n10308 = ~n1680 & n10307;
  assign n10309 = ~pi083 & ~n10308;
  assign n10310 = ~n1673 & ~n10309;
  assign n10311 = n10306 & n10310;
  assign n10312 = ~n10305 & n10311;
  assign n10313 = ~pi040 & ~n10312;
  assign n10314 = pi083 & n1681;
  assign n10315 = ~n10313 & ~n10314;
  assign n10316 = n1486 & n1517;
  assign n10317 = n10315 & ~n10316;
  assign n10318 = ~n10304 & n10317;
  assign n10319 = ~pi014 & n1718;
  assign n10320 = ~n1478 & ~n10319;
  assign n10321 = pi083 & ~n10320;
  assign n10322 = ~pi083 & n1514;
  assign n10323 = ~n10321 & ~n10322;
  assign n10324 = ~n1505 & n10323;
  assign n10325 = pi040 & ~n10324;
  assign n10326 = ~n1483 & ~n1533;
  assign n10327 = ~pi014 & n7458;
  assign n10328 = ~pi083 & n10282;
  assign n10329 = ~n10327 & ~n10328;
  assign n10330 = n10326 & n10329;
  assign n10331 = ~n7495 & n10330;
  assign n10332 = ~n1473 & n10331;
  assign n10333 = ~pi040 & ~n10332;
  assign n10334 = ~n10325 & ~n10333;
  assign n10335 = pi107 & n2668;
  assign n10336 = ~pi014 & n1557;
  assign n10337 = n1648 & ~n7490;
  assign n10338 = ~n10336 & ~n10337;
  assign n10339 = ~n10335 & n10338;
  assign n10340 = ~n1641 & n10339;
  assign n10341 = ~pi083 & ~n10340;
  assign n10342 = ~n1533 & ~n7916;
  assign n10343 = pi083 & ~n10342;
  assign n10344 = ~n10341 & ~n10343;
  assign n10345 = n10334 & n10344;
  assign n10346 = ~pi078 & ~n10345;
  assign n10347 = n10318 & ~n10346;
  assign n10348 = n10300 & n10347;
  assign n10349 = ~n10264 & n10348;
  assign n10350 = n10264 & ~n10348;
  assign n10351 = ~n10349 & ~n10350;
  assign n10352 = ~n10185 & n10351;
  assign n10353 = n10185 & ~n10351;
  assign n10354 = ~n10352 & ~n10353;
  assign n10355 = n10097 & n10354;
  assign n10356 = ~n10097 & ~n10354;
  assign n10357 = ~n10355 & ~n10356;
  assign n10358 = ~pi529 & ~n10357;
  assign n10359 = ~pi153 & pi515;
  assign n10360 = pi153 & ~pi515;
  assign n10361 = ~n10359 & ~n10360;
  assign n10362 = pi529 & ~n10361;
  assign po156 = n10358 | n10362;
  assign n10364 = pi179 & pi457;
  assign n10365 = ~pi179 & ~pi457;
  assign n10366 = ~n10364 & ~n10365;
  assign n10367 = pi529 & n10366;
  assign n10368 = pi033 & n2195;
  assign n10369 = ~n10135 & ~n10368;
  assign n10370 = ~n2550 & n10369;
  assign n10371 = n2295 & ~n10370;
  assign n10372 = ~n2206 & ~n2368;
  assign n10373 = pi069 & n2210;
  assign n10374 = ~n2563 & ~n10373;
  assign n10375 = n10372 & n10374;
  assign n10376 = pi102 & ~n10375;
  assign n10377 = pi104 & n2437;
  assign n10378 = ~n2112 & ~n2219;
  assign n10379 = ~n2307 & n10378;
  assign n10380 = ~pi104 & ~n10379;
  assign n10381 = ~n10377 & ~n10380;
  assign n10382 = ~n2373 & n10381;
  assign n10383 = ~n2133 & n10382;
  assign n10384 = ~n10376 & n10383;
  assign n10385 = ~n10371 & n10384;
  assign n10386 = ~n2112 & ~n2437;
  assign n10387 = ~n2167 & ~n2224;
  assign n10388 = pi104 & ~n10387;
  assign n10389 = ~pi104 & n2197;
  assign n10390 = ~n2249 & ~n10389;
  assign n10391 = ~n10388 & n10390;
  assign n10392 = n10386 & n10391;
  assign n10393 = ~pi102 & ~n10392;
  assign n10394 = ~n2469 & ~n10393;
  assign n10395 = n10385 & n10394;
  assign n10396 = pi012 & ~n10395;
  assign n10397 = ~pi069 & n2461;
  assign n10398 = pi069 & n2313;
  assign n10399 = ~n2138 & ~n10398;
  assign n10400 = pi069 & n2416;
  assign n10401 = n10399 & ~n10400;
  assign n10402 = ~n10397 & n10401;
  assign n10403 = pi104 & ~n10402;
  assign n10404 = ~n2179 & ~n10099;
  assign n10405 = ~pi069 & n2213;
  assign n10406 = n2090 & n2550;
  assign n10407 = ~n10405 & ~n10406;
  assign n10408 = n10404 & n10407;
  assign n10409 = ~pi102 & ~n10408;
  assign n10410 = ~n2100 & ~n2227;
  assign n10411 = pi104 & ~n10410;
  assign n10412 = ~n2283 & ~n2404;
  assign n10413 = ~pi069 & n2212;
  assign n10414 = n10412 & ~n10413;
  assign n10415 = ~pi104 & ~n10414;
  assign n10416 = ~n2317 & ~n2320;
  assign n10417 = ~n2412 & n10416;
  assign n10418 = ~n2126 & ~n10398;
  assign n10419 = n10417 & n10418;
  assign n10420 = ~n10415 & n10419;
  assign n10421 = ~n10411 & n10420;
  assign n10422 = pi102 & ~n10421;
  assign n10423 = ~n10409 & ~n10422;
  assign n10424 = ~n10403 & n10423;
  assign n10425 = ~pi104 & n2152;
  assign n10426 = ~n10136 & ~n10425;
  assign n10427 = ~n2568 & n10426;
  assign n10428 = ~n10134 & n10427;
  assign n10429 = n10424 & n10428;
  assign n10430 = ~pi012 & ~n10429;
  assign n10431 = pi069 & n2568;
  assign n10432 = ~n10425 & ~n10431;
  assign n10433 = pi102 & ~n10432;
  assign n10434 = n2266 & n2417;
  assign n10435 = ~n2394 & ~n10434;
  assign n10436 = ~n10433 & n10435;
  assign n10437 = ~n7793 & n10436;
  assign n10438 = ~n2564 & n10437;
  assign n10439 = ~pi069 & n2229;
  assign n10440 = ~n2101 & ~n10439;
  assign n10441 = ~n2132 & n10440;
  assign n10442 = ~pi104 & ~n10441;
  assign n10443 = n2200 & ~n2406;
  assign n10444 = ~n2437 & ~n10443;
  assign n10445 = pi104 & ~n10444;
  assign n10446 = n2090 & n2282;
  assign n10447 = ~n10445 & ~n10446;
  assign n10448 = ~n2396 & n10447;
  assign n10449 = ~n10442 & n10448;
  assign n10450 = ~pi102 & ~n10449;
  assign n10451 = n10438 & ~n10450;
  assign n10452 = ~n10430 & n10451;
  assign n10453 = ~n10396 & n10452;
  assign n10454 = ~pi179 & ~n10453;
  assign n10455 = pi179 & n10453;
  assign n10456 = ~n10454 & ~n10455;
  assign n10457 = ~n2243 & n10456;
  assign n10458 = n2243 & ~n10456;
  assign n10459 = ~n10457 & ~n10458;
  assign n10460 = ~n7504 & ~n10097;
  assign n10461 = n7504 & n10097;
  assign n10462 = ~n10460 & ~n10461;
  assign n10463 = n10459 & n10462;
  assign n10464 = ~n10459 & ~n10462;
  assign n10465 = ~n10463 & ~n10464;
  assign n10466 = ~pi529 & n10465;
  assign po157 = n10367 | n10466;
  assign n10468 = ~pi358 & pi481;
  assign n10469 = pi358 & ~pi481;
  assign n10470 = ~n10468 & ~n10469;
  assign n10471 = pi529 & ~n10470;
  assign n10472 = ~n5484 & n6659;
  assign n10473 = n5484 & ~n6659;
  assign n10474 = ~n10472 & ~n10473;
  assign n10475 = pi091 & n5674;
  assign n10476 = pi091 & n5766;
  assign n10477 = ~n5708 & ~n10476;
  assign n10478 = ~n5643 & ~n5664;
  assign n10479 = pi005 & ~n10478;
  assign n10480 = ~n5848 & ~n10479;
  assign n10481 = ~n6980 & n10480;
  assign n10482 = ~pi091 & ~n10481;
  assign n10483 = ~n5867 & ~n10482;
  assign n10484 = n10477 & n10483;
  assign n10485 = ~n10475 & n10484;
  assign n10486 = pi024 & ~n10485;
  assign n10487 = ~n5797 & ~n6470;
  assign n10488 = ~n6463 & n10487;
  assign n10489 = ~n5751 & n10488;
  assign n10490 = ~n5693 & n10489;
  assign n10491 = pi091 & ~n10490;
  assign n10492 = ~pi005 & n5665;
  assign n10493 = ~n6458 & ~n10492;
  assign n10494 = ~n5798 & n10493;
  assign n10495 = ~pi091 & ~n10494;
  assign n10496 = ~n5623 & ~n10495;
  assign n10497 = ~n10491 & n10496;
  assign n10498 = ~n6471 & n10497;
  assign n10499 = ~pi024 & ~n10498;
  assign n10500 = ~n10486 & ~n10499;
  assign n10501 = ~n5756 & ~n5872;
  assign n10502 = ~pi091 & ~n10501;
  assign n10503 = ~n6521 & ~n10502;
  assign n10504 = ~n6494 & n10503;
  assign n10505 = ~n5882 & n10504;
  assign n10506 = pi024 & ~n10505;
  assign n10507 = ~pi005 & ~pi094;
  assign n10508 = pi004 & n10507;
  assign n10509 = ~n5762 & ~n10508;
  assign n10510 = ~pi004 & n5657;
  assign n10511 = ~n5794 & ~n10510;
  assign n10512 = n10509 & n10511;
  assign n10513 = pi091 & ~n10512;
  assign n10514 = ~n6516 & ~n6980;
  assign n10515 = ~n5774 & n10514;
  assign n10516 = ~pi091 & ~n10515;
  assign n10517 = ~n10513 & ~n10516;
  assign n10518 = ~pi091 & n5631;
  assign n10519 = pi005 & n5630;
  assign n10520 = ~n6912 & ~n10519;
  assign n10521 = ~n5864 & n10520;
  assign n10522 = ~n10518 & n10521;
  assign n10523 = ~n5869 & n10522;
  assign n10524 = ~pi024 & ~n10523;
  assign n10525 = n10517 & ~n10524;
  assign n10526 = ~n10506 & n10525;
  assign n10527 = pi018 & ~n10526;
  assign n10528 = n10500 & ~n10527;
  assign n10529 = ~pi091 & n5761;
  assign n10530 = pi091 & n5678;
  assign n10531 = ~n10529 & ~n10530;
  assign n10532 = pi005 & ~n10531;
  assign n10533 = pi024 & n5826;
  assign n10534 = ~pi091 & n5652;
  assign n10535 = ~n10533 & ~n10534;
  assign n10536 = n5621 & n5705;
  assign n10537 = pi005 & n6485;
  assign n10538 = ~n10536 & ~n10537;
  assign n10539 = ~pi024 & ~n10538;
  assign n10540 = n10535 & ~n10539;
  assign n10541 = ~n5646 & ~n10530;
  assign n10542 = ~pi024 & ~n10541;
  assign n10543 = ~pi005 & n5654;
  assign n10544 = ~n5773 & ~n10543;
  assign n10545 = ~n5866 & n10544;
  assign n10546 = pi024 & ~pi091;
  assign n10547 = ~n10545 & n10546;
  assign n10548 = ~n10542 & ~n10547;
  assign n10549 = ~pi005 & n5721;
  assign n10550 = ~n5733 & ~n10549;
  assign n10551 = pi091 & ~n10550;
  assign n10552 = n10548 & ~n10551;
  assign n10553 = n10540 & n10552;
  assign n10554 = n5644 & n5663;
  assign n10555 = ~n5792 & ~n10554;
  assign n10556 = pi024 & ~n10555;
  assign n10557 = ~n6471 & ~n10556;
  assign n10558 = n10553 & n10557;
  assign n10559 = ~pi018 & ~n10558;
  assign n10560 = ~n10532 & ~n10559;
  assign n10561 = n10528 & n10560;
  assign n10562 = n5603 & n10561;
  assign n10563 = ~n5603 & ~n10561;
  assign n10564 = ~n10562 & ~n10563;
  assign n10565 = n10474 & n10564;
  assign n10566 = ~n10474 & ~n10564;
  assign n10567 = ~n10565 & ~n10566;
  assign n10568 = n6328 & ~n9897;
  assign n10569 = ~n6328 & n9897;
  assign n10570 = ~n10568 & ~n10569;
  assign n10571 = ~pi358 & ~n6060;
  assign n10572 = pi358 & n6060;
  assign n10573 = ~n10571 & ~n10572;
  assign n10574 = ~n10570 & n10573;
  assign n10575 = n10570 & ~n10573;
  assign n10576 = ~n10574 & ~n10575;
  assign n10577 = n10567 & n10576;
  assign n10578 = ~n10567 & ~n10576;
  assign n10579 = ~n10577 & ~n10578;
  assign n10580 = ~pi529 & n10579;
  assign po158 = n10471 | n10580;
  assign n10582 = pi302 & pi502;
  assign n10583 = ~pi302 & ~pi502;
  assign n10584 = ~n10582 & ~n10583;
  assign n10585 = pi529 & n10584;
  assign n10586 = ~pi043 & n5392;
  assign n10587 = ~pi043 & n5556;
  assign n10588 = ~pi122 & n5526;
  assign n10589 = ~n10587 & ~n10588;
  assign n10590 = n5327 & n5366;
  assign n10591 = ~n5475 & ~n10590;
  assign n10592 = ~n5527 & n10591;
  assign n10593 = n10589 & n10592;
  assign n10594 = ~pi039 & ~n10593;
  assign n10595 = pi122 & n5507;
  assign n10596 = ~n10594 & ~n10595;
  assign n10597 = ~n10586 & n10596;
  assign n10598 = ~n5358 & n10597;
  assign n10599 = ~n5360 & ~n6100;
  assign n10600 = ~n5392 & ~n5475;
  assign n10601 = n10599 & n10600;
  assign n10602 = ~pi122 & ~n10601;
  assign n10603 = ~n5464 & ~n5558;
  assign n10604 = ~n5339 & ~n5364;
  assign n10605 = ~n6346 & n10604;
  assign n10606 = pi122 & ~n10605;
  assign n10607 = n10603 & ~n10606;
  assign n10608 = pi039 & ~n10607;
  assign n10609 = ~n10602 & ~n10608;
  assign n10610 = n10598 & n10609;
  assign n10611 = pi017 & ~n10610;
  assign n10612 = ~n5487 & ~n6077;
  assign n10613 = ~pi122 & ~n10612;
  assign n10614 = ~pi043 & n5464;
  assign n10615 = ~n6407 & ~n10614;
  assign n10616 = ~pi122 & ~n10615;
  assign n10617 = pi122 & n5493;
  assign n10618 = ~n5570 & ~n10617;
  assign n10619 = ~n6077 & n10618;
  assign n10620 = ~n10616 & n10619;
  assign n10621 = ~n6396 & n10620;
  assign n10622 = ~pi039 & ~n10621;
  assign n10623 = ~pi043 & ~n5445;
  assign n10624 = pi043 & ~n5364;
  assign n10625 = ~n10623 & ~n10624;
  assign n10626 = ~n7127 & ~n10625;
  assign n10627 = ~pi122 & ~n10626;
  assign n10628 = ~n5332 & ~n5336;
  assign n10629 = pi122 & ~n10628;
  assign n10630 = ~n10627 & ~n10629;
  assign n10631 = ~n5463 & ~n6154;
  assign n10632 = ~n5348 & n10631;
  assign n10633 = n10630 & n10632;
  assign n10634 = pi039 & ~n10633;
  assign n10635 = ~n10622 & ~n10634;
  assign n10636 = ~n5513 & n10635;
  assign n10637 = ~n10613 & n10636;
  assign n10638 = ~pi043 & n7143;
  assign n10639 = ~n7153 & ~n10638;
  assign n10640 = pi122 & ~n10639;
  assign n10641 = ~n7185 & ~n10640;
  assign n10642 = n10637 & n10641;
  assign n10643 = ~pi017 & ~n10642;
  assign n10644 = ~pi043 & n5426;
  assign n10645 = ~n5384 & ~n5491;
  assign n10646 = ~n6071 & n10645;
  assign n10647 = ~n10644 & n10646;
  assign n10648 = ~pi122 & ~n10647;
  assign n10649 = pi039 & n10648;
  assign n10650 = ~n5350 & ~n5464;
  assign n10651 = pi043 & ~n10650;
  assign n10652 = ~n5358 & ~n10651;
  assign n10653 = n5456 & ~n10652;
  assign n10654 = n5494 & n6366;
  assign n10655 = ~n10653 & ~n10654;
  assign n10656 = ~n10649 & n10655;
  assign n10657 = ~n5385 & ~n5577;
  assign n10658 = ~pi043 & n5446;
  assign n10659 = ~n5534 & ~n10658;
  assign n10660 = ~n5513 & n10659;
  assign n10661 = n5354 & ~n10660;
  assign n10662 = ~n5516 & ~n7135;
  assign n10663 = ~n5369 & ~n5401;
  assign n10664 = ~n5571 & n10663;
  assign n10665 = ~pi122 & ~n10664;
  assign n10666 = n10662 & ~n10665;
  assign n10667 = ~pi039 & ~n10666;
  assign n10668 = ~n10661 & ~n10667;
  assign n10669 = n10657 & n10668;
  assign n10670 = n10656 & n10669;
  assign n10671 = ~n10643 & n10670;
  assign n10672 = ~n10611 & n10671;
  assign n10673 = ~n6542 & ~n9853;
  assign n10674 = ~pi035 & n6172;
  assign n10675 = ~n6630 & ~n10674;
  assign n10676 = ~n6566 & n10675;
  assign n10677 = n7009 & ~n10676;
  assign n10678 = ~n6302 & ~n7040;
  assign n10679 = ~n6562 & ~n7041;
  assign n10680 = ~n6261 & n10679;
  assign n10681 = ~pi106 & ~n10680;
  assign n10682 = n10678 & ~n10681;
  assign n10683 = ~pi065 & ~n10682;
  assign n10684 = ~n10677 & ~n10683;
  assign n10685 = n10673 & n10684;
  assign n10686 = ~n6203 & ~n6543;
  assign n10687 = pi035 & ~n10686;
  assign n10688 = ~n6167 & ~n10687;
  assign n10689 = n9872 & ~n10688;
  assign n10690 = ~pi035 & n6294;
  assign n10691 = ~n6552 & ~n9852;
  assign n10692 = ~n6300 & n10691;
  assign n10693 = ~n10690 & n10692;
  assign n10694 = ~pi106 & ~n10693;
  assign n10695 = n6197 & n6617;
  assign n10696 = ~n10694 & ~n10695;
  assign n10697 = pi065 & ~n10696;
  assign n10698 = ~n10689 & ~n10697;
  assign n10699 = ~pi031 & n6272;
  assign n10700 = ~n7060 & ~n10699;
  assign n10701 = pi106 & ~n10700;
  assign n10702 = ~n7097 & ~n10701;
  assign n10703 = ~n6310 & ~n6556;
  assign n10704 = ~pi106 & ~n10703;
  assign n10705 = ~n6566 & ~n10704;
  assign n10706 = ~pi035 & n6169;
  assign n10707 = pi035 & n6312;
  assign n10708 = ~n7005 & ~n10707;
  assign n10709 = ~n10706 & n10708;
  assign n10710 = ~pi106 & ~n10709;
  assign n10711 = ~n6283 & ~n6301;
  assign n10712 = ~n9824 & n10711;
  assign n10713 = ~n6227 & ~n6584;
  assign n10714 = pi106 & ~n10713;
  assign n10715 = n10712 & ~n10714;
  assign n10716 = ~n10710 & n10715;
  assign n10717 = pi065 & ~n10716;
  assign n10718 = n6165 & n6297;
  assign n10719 = ~n6540 & ~n10718;
  assign n10720 = ~pi106 & ~n10719;
  assign n10721 = pi106 & n6284;
  assign n10722 = ~n6541 & ~n10721;
  assign n10723 = ~n10720 & n10722;
  assign n10724 = ~n6310 & n10723;
  assign n10725 = pi106 & n6200;
  assign n10726 = n10724 & ~n10725;
  assign n10727 = ~pi065 & ~n10726;
  assign n10728 = ~n10717 & ~n10727;
  assign n10729 = n10705 & n10728;
  assign n10730 = n10702 & n10729;
  assign n10731 = ~pi068 & ~n10730;
  assign n10732 = n6246 & n6570;
  assign n10733 = ~n6323 & ~n10732;
  assign n10734 = ~n6598 & n10733;
  assign n10735 = ~pi106 & n6597;
  assign n10736 = ~pi035 & n6603;
  assign n10737 = ~n10735 & ~n10736;
  assign n10738 = n10734 & n10737;
  assign n10739 = ~pi065 & ~n10738;
  assign n10740 = ~n6200 & ~n9817;
  assign n10741 = ~n6323 & ~n7039;
  assign n10742 = n10740 & n10741;
  assign n10743 = ~pi106 & ~n10742;
  assign n10744 = ~pi035 & n7039;
  assign n10745 = ~n10743 & ~n10744;
  assign n10746 = pi106 & n6311;
  assign n10747 = n10745 & ~n10746;
  assign n10748 = ~n10739 & n10747;
  assign n10749 = ~n6167 & n10748;
  assign n10750 = ~n6543 & ~n6606;
  assign n10751 = ~n6554 & ~n7024;
  assign n10752 = ~n6312 & n10751;
  assign n10753 = pi106 & ~n10752;
  assign n10754 = n10750 & ~n10753;
  assign n10755 = pi065 & ~n10754;
  assign n10756 = n10749 & ~n10755;
  assign n10757 = pi068 & ~n10756;
  assign n10758 = ~n10731 & ~n10757;
  assign n10759 = n10698 & n10758;
  assign n10760 = n10685 & n10759;
  assign n10761 = ~n10672 & n10760;
  assign n10762 = n10672 & ~n10760;
  assign n10763 = ~n10761 & ~n10762;
  assign n10764 = ~pi009 & n5929;
  assign n10765 = ~n6723 & ~n10764;
  assign n10766 = ~n6691 & n10765;
  assign n10767 = n6852 & ~n10766;
  assign n10768 = ~n6000 & ~n6827;
  assign n10769 = ~n6811 & n10768;
  assign n10770 = ~pi113 & ~n10769;
  assign n10771 = ~n6680 & ~n10770;
  assign n10772 = ~n9576 & n10771;
  assign n10773 = ~pi096 & ~n10772;
  assign n10774 = ~n10767 & ~n10773;
  assign n10775 = ~pi009 & n6814;
  assign n10776 = ~n6825 & ~n9593;
  assign n10777 = ~n5941 & ~n6814;
  assign n10778 = n10776 & n10777;
  assign n10779 = ~pi113 & ~n10778;
  assign n10780 = ~pi009 & n6730;
  assign n10781 = ~pi113 & n6673;
  assign n10782 = ~n10780 & ~n10781;
  assign n10783 = n5978 & n6681;
  assign n10784 = ~n6674 & ~n10783;
  assign n10785 = ~n5941 & n10784;
  assign n10786 = n10782 & n10785;
  assign n10787 = ~pi096 & ~n10786;
  assign n10788 = ~n6830 & ~n10787;
  assign n10789 = ~n10779 & n10788;
  assign n10790 = ~n10775 & n10789;
  assign n10791 = pi113 & n6053;
  assign n10792 = ~n6732 & ~n6766;
  assign n10793 = ~n6049 & ~n6663;
  assign n10794 = ~n9692 & n10793;
  assign n10795 = pi113 & ~n10794;
  assign n10796 = n10792 & ~n10795;
  assign n10797 = pi096 & ~n10796;
  assign n10798 = ~n10791 & ~n10797;
  assign n10799 = n10790 & n10798;
  assign n10800 = ~pi010 & ~n10799;
  assign n10801 = ~n5937 & ~n6766;
  assign n10802 = pi009 & ~n10801;
  assign n10803 = ~n6830 & ~n10802;
  assign n10804 = n6842 & ~n10803;
  assign n10805 = ~n6768 & ~n6819;
  assign n10806 = ~n10804 & n10805;
  assign n10807 = n5916 & n6685;
  assign n10808 = ~pi125 & n5916;
  assign n10809 = ~n6671 & ~n10808;
  assign n10810 = ~pi009 & n6039;
  assign n10811 = ~n6035 & ~n10810;
  assign n10812 = n10809 & n10811;
  assign n10813 = ~pi113 & ~n10812;
  assign n10814 = ~n10807 & ~n10813;
  assign n10815 = pi096 & ~n10814;
  assign n10816 = n10806 & ~n10815;
  assign n10817 = ~pi113 & n6051;
  assign n10818 = ~n9652 & ~n10817;
  assign n10819 = ~n6691 & n10818;
  assign n10820 = pi113 & n6027;
  assign n10821 = ~pi025 & n5917;
  assign n10822 = n5910 & n10821;
  assign n10823 = ~n6770 & ~n10822;
  assign n10824 = ~pi113 & ~n10823;
  assign n10825 = ~n6051 & ~n10824;
  assign n10826 = ~n6771 & ~n9715;
  assign n10827 = n10825 & n10826;
  assign n10828 = ~n10820 & n10827;
  assign n10829 = ~pi096 & ~n10828;
  assign n10830 = ~n6026 & ~n6041;
  assign n10831 = ~n6848 & n10830;
  assign n10832 = ~n6708 & ~n6803;
  assign n10833 = pi113 & ~n10832;
  assign n10834 = ~pi009 & ~n5928;
  assign n10835 = pi009 & ~n6049;
  assign n10836 = ~n10834 & ~n10835;
  assign n10837 = ~pi125 & n6756;
  assign n10838 = ~n10836 & ~n10837;
  assign n10839 = ~pi113 & ~n10838;
  assign n10840 = ~n10833 & ~n10839;
  assign n10841 = n10831 & n10840;
  assign n10842 = pi096 & ~n10841;
  assign n10843 = ~n10829 & ~n10842;
  assign n10844 = n10819 & n10843;
  assign n10845 = ~pi124 & n5917;
  assign n10846 = ~n9582 & ~n10845;
  assign n10847 = pi113 & ~n10846;
  assign n10848 = ~n9622 & ~n10847;
  assign n10849 = n10844 & n10848;
  assign n10850 = pi010 & ~n10849;
  assign n10851 = n10816 & ~n10850;
  assign n10852 = ~n10800 & n10851;
  assign n10853 = n10774 & n10852;
  assign n10854 = ~pi302 & ~n10853;
  assign n10855 = pi302 & n10853;
  assign n10856 = ~n10854 & ~n10855;
  assign n10857 = ~n10763 & n10856;
  assign n10858 = n10763 & ~n10856;
  assign n10859 = ~n10857 & ~n10858;
  assign n10860 = n5484 & ~n7192;
  assign n10861 = ~n5484 & n7192;
  assign n10862 = ~n10860 & ~n10861;
  assign n10863 = ~n7004 & n10862;
  assign n10864 = ~n7199 & ~n10862;
  assign n10865 = ~n10863 & ~n10864;
  assign n10866 = n10859 & n10865;
  assign n10867 = ~n10859 & ~n10865;
  assign n10868 = ~n10866 & ~n10867;
  assign n10869 = ~pi529 & n10868;
  assign po159 = n10585 | n10869;
  assign n10871 = pi142 & pi400;
  assign n10872 = ~pi142 & ~pi400;
  assign n10873 = ~n10871 & ~n10872;
  assign n10874 = pi529 & n10873;
  assign n10875 = n1587 & n1716;
  assign n10876 = ~pi083 & n1653;
  assign n10877 = ~n2618 & ~n10876;
  assign n10878 = ~n7531 & n10877;
  assign n10879 = ~n10875 & n10878;
  assign n10880 = ~pi083 & n1629;
  assign n10881 = pi014 & n1514;
  assign n10882 = ~n10880 & ~n10881;
  assign n10883 = pi040 & ~n10882;
  assign n10884 = n10879 & ~n10883;
  assign n10885 = ~n1464 & n2629;
  assign n10886 = ~pi083 & ~n10885;
  assign n10887 = pi083 & n1730;
  assign n10888 = ~n10886 & ~n10887;
  assign n10889 = ~n1649 & n10888;
  assign n10890 = ~n7595 & n10889;
  assign n10891 = pi014 & pi072;
  assign n10892 = ~pi107 & n10891;
  assign n10893 = ~n2624 & ~n10892;
  assign n10894 = ~n10279 & n10893;
  assign n10895 = pi040 & ~n10894;
  assign n10896 = ~pi083 & n10895;
  assign n10897 = ~n1630 & ~n1707;
  assign n10898 = ~n2590 & ~n7944;
  assign n10899 = n10897 & n10898;
  assign n10900 = pi040 & ~n10899;
  assign n10901 = ~n10896 & ~n10900;
  assign n10902 = n10890 & n10901;
  assign n10903 = ~n1613 & ~n1730;
  assign n10904 = ~pi083 & n1656;
  assign n10905 = pi014 & n1742;
  assign n10906 = ~n1575 & ~n10905;
  assign n10907 = pi083 & ~n10906;
  assign n10908 = ~n10904 & ~n10907;
  assign n10909 = n10903 & n10908;
  assign n10910 = ~n1561 & n10909;
  assign n10911 = ~pi040 & ~n10910;
  assign n10912 = ~n1709 & ~n10911;
  assign n10913 = n10902 & n10912;
  assign n10914 = pi078 & n10913;
  assign n10915 = ~n1721 & ~n10316;
  assign n10916 = ~pi014 & n1618;
  assign n10917 = n1508 & n2624;
  assign n10918 = ~n10916 & ~n10917;
  assign n10919 = n10915 & n10918;
  assign n10920 = ~pi040 & ~n10919;
  assign n10921 = pi014 & n1477;
  assign n10922 = ~n1663 & ~n10921;
  assign n10923 = pi014 & n1718;
  assign n10924 = ~n7965 & ~n10923;
  assign n10925 = n10922 & n10924;
  assign n10926 = pi083 & ~n10925;
  assign n10927 = ~n10278 & ~n10880;
  assign n10928 = ~n1514 & n10927;
  assign n10929 = ~n10280 & n10928;
  assign n10930 = ~n10926 & n10929;
  assign n10931 = ~n1580 & ~n1672;
  assign n10932 = ~pi014 & n1701;
  assign n10933 = n10931 & ~n10932;
  assign n10934 = ~pi083 & ~n10933;
  assign n10935 = ~n1653 & ~n10921;
  assign n10936 = ~n1504 & ~n7464;
  assign n10937 = pi083 & ~n10936;
  assign n10938 = n10935 & ~n10937;
  assign n10939 = ~n10934 & n10938;
  assign n10940 = ~n1499 & ~n1699;
  assign n10941 = ~n1484 & n10940;
  assign n10942 = n10939 & n10941;
  assign n10943 = pi040 & ~n10942;
  assign n10944 = n10930 & ~n10943;
  assign n10945 = ~n10920 & n10944;
  assign n10946 = ~pi078 & n10945;
  assign n10947 = ~n10914 & ~n10946;
  assign n10948 = ~pi014 & n1541;
  assign n10949 = ~n1505 & ~n10948;
  assign n10950 = ~n1493 & n10949;
  assign n10951 = n1683 & ~n10950;
  assign n10952 = n1532 & ~n1674;
  assign n10953 = ~n1730 & ~n10952;
  assign n10954 = pi083 & ~n10953;
  assign n10955 = n1508 & n1579;
  assign n10956 = ~n1664 & ~n10955;
  assign n10957 = ~n10954 & n10956;
  assign n10958 = ~pi040 & ~n10957;
  assign n10959 = ~n10951 & ~n10958;
  assign n10960 = ~n10947 & n10959;
  assign n10961 = n10884 & n10960;
  assign n10962 = n2243 & ~n10961;
  assign n10963 = ~n2243 & n10961;
  assign n10964 = ~n10962 & ~n10963;
  assign n10965 = ~pi142 & n10964;
  assign n10966 = pi142 & ~n10964;
  assign n10967 = ~n10965 & ~n10966;
  assign n10968 = n1915 & n10097;
  assign n10969 = ~n1915 & ~n10097;
  assign n10970 = ~n10968 & ~n10969;
  assign n10971 = ~n10967 & n10970;
  assign n10972 = n10967 & ~n10970;
  assign n10973 = ~n10971 & ~n10972;
  assign n10974 = ~pi529 & n10973;
  assign po160 = n10874 | n10974;
  assign n10976 = pi173 & pi407;
  assign n10977 = ~pi173 & ~pi407;
  assign n10978 = ~n10976 & ~n10977;
  assign n10979 = pi529 & n10978;
  assign n10980 = pi013 & n1786;
  assign n10981 = ~n7359 & ~n10980;
  assign n10982 = ~n1759 & n10981;
  assign n10983 = n2886 & ~n10982;
  assign n10984 = pi001 & n1765;
  assign n10985 = n7372 & n10984;
  assign n10986 = ~n10983 & ~n10985;
  assign n10987 = ~n2829 & ~n7358;
  assign n10988 = ~pi013 & n1836;
  assign n10989 = ~pi007 & n1792;
  assign n10990 = ~n2828 & ~n10989;
  assign n10991 = ~n1842 & n10990;
  assign n10992 = ~n10988 & n10991;
  assign n10993 = n1782 & ~n10992;
  assign n10994 = ~n1878 & ~n2848;
  assign n10995 = ~n2837 & n10994;
  assign n10996 = n7340 & ~n10995;
  assign n10997 = ~pi013 & n1775;
  assign n10998 = ~n7332 & ~n10997;
  assign n10999 = ~n7378 & n10998;
  assign n11000 = n2914 & ~n10999;
  assign n11001 = ~n2974 & ~n7326;
  assign n11002 = ~pi001 & ~n11001;
  assign n11003 = ~n11000 & ~n11002;
  assign n11004 = ~n10996 & n11003;
  assign n11005 = ~n10993 & n11004;
  assign n11006 = n10987 & n11005;
  assign n11007 = n10986 & n11006;
  assign n11008 = ~pi114 & n7316;
  assign n11009 = n1838 & n2820;
  assign n11010 = ~pi013 & n7344;
  assign n11011 = ~n11009 & ~n11010;
  assign n11012 = ~n11008 & n11011;
  assign n11013 = ~n1863 & ~n7317;
  assign n11014 = n11012 & n11013;
  assign n11015 = ~pi001 & ~n11014;
  assign n11016 = ~n1849 & ~n2875;
  assign n11017 = ~n2952 & n11016;
  assign n11018 = n2886 & ~n11017;
  assign n11019 = ~n2922 & ~n7394;
  assign n11020 = pi001 & ~n11019;
  assign n11021 = ~n1759 & ~n11020;
  assign n11022 = ~n11018 & n11021;
  assign n11023 = ~pi013 & n2830;
  assign n11024 = ~n2845 & ~n2969;
  assign n11025 = ~n1863 & ~n2830;
  assign n11026 = n11024 & n11025;
  assign n11027 = ~pi114 & ~n11026;
  assign n11028 = ~n11023 & ~n11027;
  assign n11029 = n11022 & n11028;
  assign n11030 = pi114 & n1853;
  assign n11031 = n11029 & ~n11030;
  assign n11032 = ~n11015 & n11031;
  assign n11033 = pi029 & ~n11032;
  assign n11034 = pi114 & n1890;
  assign n11035 = ~n7881 & ~n11034;
  assign n11036 = ~pi001 & ~n11035;
  assign n11037 = ~pi013 & n2922;
  assign n11038 = ~n2980 & ~n11037;
  assign n11039 = ~pi114 & ~n11038;
  assign n11040 = ~n7362 & ~n11039;
  assign n11041 = ~n1851 & n11040;
  assign n11042 = ~pi001 & ~n11041;
  assign n11043 = ~n1851 & ~n2961;
  assign n11044 = ~pi114 & ~n11043;
  assign n11045 = ~n7332 & ~n11044;
  assign n11046 = ~n2823 & ~n2910;
  assign n11047 = n2886 & ~n11046;
  assign n11048 = n11045 & ~n11047;
  assign n11049 = ~n11042 & n11048;
  assign n11050 = ~n11036 & n11049;
  assign n11051 = ~pi013 & ~n1774;
  assign n11052 = pi013 & ~n1849;
  assign n11053 = ~n11051 & ~n11052;
  assign n11054 = ~n2958 & ~n11053;
  assign n11055 = ~pi114 & ~n11054;
  assign n11056 = n10002 & ~n11055;
  assign n11057 = ~n2917 & n11056;
  assign n11058 = pi001 & ~n11057;
  assign n11059 = ~pi013 & n2998;
  assign n11060 = ~n2985 & ~n11059;
  assign n11061 = pi114 & ~n11060;
  assign n11062 = ~n3030 & ~n11061;
  assign n11063 = ~n11058 & n11062;
  assign n11064 = n11050 & n11063;
  assign n11065 = ~pi029 & ~n11064;
  assign n11066 = ~n11033 & ~n11065;
  assign n11067 = n11007 & n11066;
  assign n11068 = ~n3141 & n11067;
  assign n11069 = n3141 & ~n11067;
  assign n11070 = ~n11068 & ~n11069;
  assign n11071 = n3238 & ~n7988;
  assign n11072 = ~n3238 & n7988;
  assign n11073 = ~n11071 & ~n11072;
  assign n11074 = ~n11070 & n11073;
  assign n11075 = n11070 & ~n11073;
  assign n11076 = ~n11074 & ~n11075;
  assign n11077 = ~pi173 & ~n2586;
  assign n11078 = pi173 & n2586;
  assign n11079 = ~n11077 & ~n11078;
  assign n11080 = n1627 & ~n2689;
  assign n11081 = ~n1627 & n2689;
  assign n11082 = ~n11080 & ~n11081;
  assign n11083 = ~n11079 & n11082;
  assign n11084 = n11079 & ~n11082;
  assign n11085 = ~n11083 & ~n11084;
  assign n11086 = n11076 & n11085;
  assign n11087 = ~n11076 & ~n11085;
  assign n11088 = ~n11086 & ~n11087;
  assign n11089 = ~pi529 & n11088;
  assign po161 = n10979 | n11089;
  assign n11091 = ~pi132 & pi447;
  assign n11092 = pi132 & ~pi447;
  assign n11093 = ~n11091 & ~n11092;
  assign n11094 = pi529 & ~n11093;
  assign n11095 = ~n6185 & ~n6192;
  assign n11096 = n6184 & ~n11095;
  assign n11097 = ~pi031 & n11096;
  assign n11098 = ~n6643 & ~n11097;
  assign n11099 = pi128 & n6296;
  assign n11100 = ~n6220 & ~n11099;
  assign n11101 = n9872 & ~n11100;
  assign n11102 = n6324 & n9872;
  assign n11103 = ~n11101 & ~n11102;
  assign n11104 = n11098 & n11103;
  assign n11105 = pi031 & n10706;
  assign n11106 = ~n6543 & ~n11105;
  assign n11107 = ~pi106 & ~n11106;
  assign n11108 = ~pi106 & n6606;
  assign n11109 = ~n11107 & ~n11108;
  assign n11110 = ~n6311 & n11109;
  assign n11111 = pi065 & ~n11110;
  assign n11112 = n11104 & ~n11111;
  assign n11113 = pi035 & n6648;
  assign n11114 = ~n6193 & ~n6598;
  assign n11115 = ~n6308 & n11114;
  assign n11116 = ~pi106 & ~n11115;
  assign n11117 = ~n11113 & ~n11116;
  assign n11118 = pi035 & n6647;
  assign n11119 = ~n6585 & ~n11118;
  assign n11120 = ~n6310 & n11119;
  assign n11121 = pi106 & ~n11120;
  assign n11122 = n6192 & n6645;
  assign n11123 = ~n6173 & ~n11122;
  assign n11124 = ~n11121 & n11123;
  assign n11125 = n11117 & n11124;
  assign n11126 = ~pi065 & ~n11125;
  assign n11127 = ~pi106 & n6566;
  assign n11128 = pi106 & n6578;
  assign n11129 = ~n6260 & ~n11128;
  assign n11130 = ~n6180 & n11129;
  assign n11131 = ~pi106 & n6220;
  assign n11132 = ~n6251 & ~n11131;
  assign n11133 = n11130 & n11132;
  assign n11134 = ~n11127 & n11133;
  assign n11135 = ~n6300 & ~n7055;
  assign n11136 = n11134 & n11135;
  assign n11137 = ~pi065 & ~n11136;
  assign n11138 = pi106 & n6195;
  assign n11139 = pi100 & n6164;
  assign n11140 = ~n6648 & ~n11139;
  assign n11141 = ~pi106 & ~n11140;
  assign n11142 = ~n7088 & ~n11141;
  assign n11143 = ~n11138 & n11142;
  assign n11144 = pi065 & ~n11143;
  assign n11145 = ~n11137 & ~n11144;
  assign n11146 = ~n6540 & ~n7039;
  assign n11147 = ~n6226 & n11146;
  assign n11148 = n6320 & ~n11147;
  assign n11149 = ~n6194 & ~n11148;
  assign n11150 = ~n10725 & n11149;
  assign n11151 = ~n6298 & n11150;
  assign n11152 = n11145 & n11151;
  assign n11153 = pi068 & ~n11152;
  assign n11154 = pi106 & n6221;
  assign n11155 = ~pi106 & n6268;
  assign n11156 = n6192 & n11155;
  assign n11157 = ~n6175 & ~n11156;
  assign n11158 = ~n7024 & ~n7049;
  assign n11159 = ~n6610 & n11158;
  assign n11160 = ~pi106 & ~n11159;
  assign n11161 = ~n9817 & ~n11160;
  assign n11162 = ~n6283 & ~n7020;
  assign n11163 = pi106 & ~n11162;
  assign n11164 = n11161 & ~n11163;
  assign n11165 = pi065 & ~n11164;
  assign n11166 = n6570 & n6617;
  assign n11167 = ~n6585 & ~n11166;
  assign n11168 = ~pi065 & ~n11167;
  assign n11169 = ~n11165 & ~n11168;
  assign n11170 = n11157 & n11169;
  assign n11171 = ~n11154 & n11170;
  assign n11172 = ~pi068 & ~n11171;
  assign n11173 = ~n11153 & ~n11172;
  assign n11174 = ~n11126 & n11173;
  assign n11175 = n11112 & n11174;
  assign n11176 = n5484 & ~n11175;
  assign n11177 = ~n5484 & n11175;
  assign n11178 = ~n11176 & ~n11177;
  assign n11179 = ~n6431 & n9779;
  assign n11180 = n6431 & ~n9779;
  assign n11181 = ~n11179 & ~n11180;
  assign n11182 = ~n11178 & n11181;
  assign n11183 = n11178 & ~n11181;
  assign n11184 = ~n11182 & ~n11183;
  assign n11185 = n6659 & ~n9897;
  assign n11186 = ~n6659 & n9897;
  assign n11187 = ~n11185 & ~n11186;
  assign n11188 = ~pi132 & ~n6783;
  assign n11189 = pi132 & n6783;
  assign n11190 = ~n11188 & ~n11189;
  assign n11191 = ~n11187 & n11190;
  assign n11192 = n11187 & ~n11190;
  assign n11193 = ~n11191 & ~n11192;
  assign n11194 = n11184 & n11193;
  assign n11195 = ~n11184 & ~n11193;
  assign n11196 = ~n11194 & ~n11195;
  assign n11197 = ~pi529 & n11196;
  assign po162 = n11094 | n11197;
  assign n11199 = ~pi175 & pi416;
  assign n11200 = pi175 & ~pi416;
  assign n11201 = ~n11199 & ~n11200;
  assign n11202 = pi529 & ~n11201;
  assign n11203 = ~n6906 & n9771;
  assign n11204 = n6906 & ~n9771;
  assign n11205 = ~n11203 & ~n11204;
  assign n11206 = ~pi175 & ~n6783;
  assign n11207 = pi175 & n6783;
  assign n11208 = ~n11206 & ~n11207;
  assign n11209 = ~n11205 & n11208;
  assign n11210 = n11205 & ~n11208;
  assign n11211 = ~n11209 & ~n11210;
  assign n11212 = n9897 & ~n11175;
  assign n11213 = ~n9897 & n11175;
  assign n11214 = ~n11212 & ~n11213;
  assign n11215 = n9782 & n11214;
  assign n11216 = ~n9782 & ~n11214;
  assign n11217 = ~n11215 & ~n11216;
  assign n11218 = ~n11211 & n11217;
  assign n11219 = n11211 & ~n11217;
  assign n11220 = ~n11218 & ~n11219;
  assign n11221 = ~pi529 & n11220;
  assign po163 = n11202 | n11221;
  assign n11223 = pi164 & pi448;
  assign n11224 = ~pi164 & ~pi448;
  assign n11225 = ~n11223 & ~n11224;
  assign n11226 = pi529 & n11225;
  assign n11227 = pi104 & n2091;
  assign n11228 = ~pi126 & n11227;
  assign n11229 = n2105 & n11228;
  assign n11230 = n2106 & n2120;
  assign n11231 = ~pi104 & n11230;
  assign n11232 = ~n11229 & ~n11231;
  assign n11233 = ~n2098 & ~n2185;
  assign n11234 = ~pi069 & n2086;
  assign n11235 = n11233 & ~n11234;
  assign n11236 = ~pi104 & ~n11235;
  assign n11237 = ~n2564 & ~n7758;
  assign n11238 = ~n2397 & ~n7750;
  assign n11239 = pi104 & ~n11238;
  assign n11240 = n11237 & ~n11239;
  assign n11241 = ~n11236 & n11240;
  assign n11242 = ~pi102 & ~n11241;
  assign n11243 = n11232 & ~n11242;
  assign n11244 = ~pi104 & n2091;
  assign n11245 = ~n2378 & ~n11244;
  assign n11246 = ~n2461 & n11245;
  assign n11247 = pi102 & ~n11246;
  assign n11248 = n2135 & n2213;
  assign n11249 = ~n2100 & ~n2132;
  assign n11250 = ~n2559 & n11249;
  assign n11251 = pi104 & ~n11250;
  assign n11252 = ~n11248 & ~n11251;
  assign n11253 = ~pi033 & n2195;
  assign n11254 = ~n2308 & ~n11253;
  assign n11255 = ~n10373 & n11254;
  assign n11256 = n11252 & n11255;
  assign n11257 = ~pi102 & ~n11256;
  assign n11258 = ~n2278 & ~n2341;
  assign n11259 = ~pi104 & ~n11258;
  assign n11260 = ~pi126 & n2195;
  assign n11261 = ~n7778 & ~n11260;
  assign n11262 = ~pi104 & ~n11261;
  assign n11263 = ~n11259 & ~n11262;
  assign n11264 = ~n2511 & n11263;
  assign n11265 = ~n2337 & ~n2563;
  assign n11266 = ~n2368 & n11265;
  assign n11267 = ~n2150 & n11266;
  assign n11268 = pi104 & ~n11267;
  assign n11269 = n11264 & ~n11268;
  assign n11270 = ~n11257 & n11269;
  assign n11271 = ~n11247 & n11270;
  assign n11272 = ~n2184 & n11271;
  assign n11273 = pi012 & ~n11272;
  assign n11274 = n2135 & n2160;
  assign n11275 = pi104 & n2112;
  assign n11276 = ~n11230 & ~n11275;
  assign n11277 = ~n11274 & n11276;
  assign n11278 = ~n2138 & ~n2267;
  assign n11279 = n11277 & n11278;
  assign n11280 = pi102 & ~n11279;
  assign n11281 = ~pi069 & ~n2291;
  assign n11282 = ~n2225 & ~n11281;
  assign n11283 = ~pi102 & ~n11282;
  assign n11284 = ~n2096 & ~n2117;
  assign n11285 = n7716 & ~n11284;
  assign n11286 = pi069 & n11285;
  assign n11287 = ~n2367 & ~n10168;
  assign n11288 = ~pi104 & ~n11287;
  assign n11289 = ~n11286 & ~n11288;
  assign n11290 = ~n2529 & n11289;
  assign n11291 = ~pi069 & n2226;
  assign n11292 = ~n2148 & ~n11291;
  assign n11293 = n2324 & ~n11292;
  assign n11294 = n11290 & ~n11293;
  assign n11295 = ~n11283 & n11294;
  assign n11296 = ~n11280 & n11295;
  assign n11297 = ~pi012 & ~n11296;
  assign n11298 = ~pi104 & n2314;
  assign n11299 = pi104 & n10397;
  assign n11300 = ~n2208 & ~n2390;
  assign n11301 = ~n11299 & n11300;
  assign n11302 = ~n11298 & n11301;
  assign n11303 = ~n2181 & n11302;
  assign n11304 = pi102 & ~n11303;
  assign n11305 = ~n11297 & ~n11304;
  assign n11306 = ~n11273 & n11305;
  assign n11307 = n11243 & n11306;
  assign n11308 = ~pi164 & ~n11307;
  assign n11309 = pi164 & n11307;
  assign n11310 = ~n11308 & ~n11309;
  assign n11311 = n2937 & ~n3238;
  assign n11312 = ~n2937 & n3238;
  assign n11313 = ~n11311 & ~n11312;
  assign n11314 = ~n7991 & n11313;
  assign n11315 = ~n7989 & ~n11313;
  assign n11316 = ~n7990 & n11315;
  assign n11317 = ~n11314 & ~n11316;
  assign n11318 = n11310 & n11317;
  assign n11319 = ~n11310 & ~n11317;
  assign n11320 = ~n11318 & ~n11319;
  assign n11321 = ~pi529 & n11320;
  assign po164 = n11226 | n11321;
  assign n11323 = pi154 & pi516;
  assign n11324 = ~pi154 & ~pi516;
  assign n11325 = ~n11323 & ~n11324;
  assign n11326 = pi529 & n11325;
  assign n11327 = ~pi154 & ~n11307;
  assign n11328 = pi154 & n11307;
  assign n11329 = ~n11327 & ~n11328;
  assign n11330 = ~n1627 & n7988;
  assign n11331 = n1627 & ~n7988;
  assign n11332 = ~n11330 & ~n11331;
  assign n11333 = ~n3040 & n3238;
  assign n11334 = n3040 & ~n3238;
  assign n11335 = ~n11333 & ~n11334;
  assign n11336 = ~n11332 & n11335;
  assign n11337 = n11332 & ~n11335;
  assign n11338 = ~n11336 & ~n11337;
  assign n11339 = n11329 & n11338;
  assign n11340 = ~n11329 & ~n11338;
  assign n11341 = ~n11339 & ~n11340;
  assign n11342 = ~pi529 & n11341;
  assign po165 = n11326 | n11342;
  assign n11344 = ~pi301 & pi512;
  assign n11345 = pi301 & ~pi512;
  assign n11346 = ~n11344 & ~n11345;
  assign n11347 = pi529 & ~n11346;
  assign n11348 = ~n3470 & ~n3517;
  assign n11349 = ~pi085 & n3439;
  assign n11350 = ~n8232 & ~n11349;
  assign n11351 = ~n3427 & n11350;
  assign n11352 = ~pi028 & ~n11351;
  assign n11353 = n11348 & ~n11352;
  assign n11354 = pi092 & ~n11353;
  assign n11355 = pi085 & n3478;
  assign n11356 = n8191 & ~n11355;
  assign n11357 = pi028 & ~n11356;
  assign n11358 = pi028 & n3449;
  assign n11359 = ~n11357 & ~n11358;
  assign n11360 = ~pi092 & ~n11359;
  assign n11361 = ~n11354 & ~n11360;
  assign n11362 = pi089 & ~n11361;
  assign n11363 = pi028 & n8161;
  assign n11364 = ~pi028 & n3472;
  assign n11365 = ~n11363 & ~n11364;
  assign n11366 = ~n3519 & n11365;
  assign n11367 = n3446 & ~n11366;
  assign n11368 = ~n3522 & ~n8172;
  assign n11369 = ~pi092 & ~n11368;
  assign n11370 = pi028 & n3576;
  assign n11371 = ~pi092 & n11370;
  assign n11372 = ~n11369 & ~n11371;
  assign n11373 = ~n8236 & n11372;
  assign n11374 = ~pi089 & ~n11373;
  assign n11375 = pi028 & n3460;
  assign n11376 = ~n8224 & ~n11375;
  assign n11377 = ~pi092 & ~n11376;
  assign n11378 = ~n11374 & ~n11377;
  assign n11379 = ~n11367 & n11378;
  assign n11380 = ~pi092 & n8255;
  assign n11381 = n3426 & n8174;
  assign n11382 = ~n11363 & ~n11381;
  assign n11383 = pi089 & ~n11382;
  assign n11384 = pi085 & n3530;
  assign n11385 = ~n8213 & ~n11384;
  assign n11386 = pi028 & n3453;
  assign n11387 = pi046 & ~pi085;
  assign n11388 = ~n11386 & ~n11387;
  assign n11389 = n11385 & n11388;
  assign n11390 = n3476 & ~n11389;
  assign n11391 = ~n11383 & ~n11390;
  assign n11392 = ~pi085 & n3526;
  assign n11393 = n3433 & n11392;
  assign n11394 = ~pi028 & n11349;
  assign n11395 = ~pi028 & n11355;
  assign n11396 = ~n11394 & ~n11395;
  assign n11397 = ~n8162 & n11396;
  assign n11398 = pi092 & ~n11397;
  assign n11399 = ~n11393 & ~n11398;
  assign n11400 = ~n8147 & n11399;
  assign n11401 = ~n3472 & ~n11384;
  assign n11402 = ~n8254 & n11401;
  assign n11403 = ~pi092 & ~n11402;
  assign n11404 = ~pi092 & n3482;
  assign n11405 = ~pi028 & n3576;
  assign n11406 = pi092 & n11405;
  assign n11407 = ~pi028 & n3453;
  assign n11408 = ~pi092 & n11407;
  assign n11409 = ~n11406 & ~n11408;
  assign n11410 = ~n11404 & n11409;
  assign n11411 = ~n11403 & n11410;
  assign n11412 = pi028 & n3479;
  assign n11413 = ~n8255 & ~n11412;
  assign n11414 = n11411 & n11413;
  assign n11415 = ~pi089 & ~n11414;
  assign n11416 = n11400 & ~n11415;
  assign n11417 = n11391 & n11416;
  assign n11418 = ~n11380 & n11417;
  assign n11419 = pi053 & ~n11418;
  assign n11420 = pi028 & n8162;
  assign n11421 = ~n3460 & ~n11420;
  assign n11422 = ~pi092 & ~n11421;
  assign n11423 = ~n3441 & ~n3450;
  assign n11424 = n3433 & ~n11423;
  assign n11425 = ~n3434 & ~n11424;
  assign n11426 = n3508 & n3527;
  assign n11427 = pi028 & ~pi046;
  assign n11428 = pi085 & n11427;
  assign n11429 = ~n3455 & ~n11428;
  assign n11430 = ~pi092 & ~n11429;
  assign n11431 = ~n11426 & ~n11430;
  assign n11432 = ~n3566 & n11431;
  assign n11433 = ~n3469 & n11432;
  assign n11434 = pi089 & ~n11433;
  assign n11435 = ~n11369 & ~n11434;
  assign n11436 = n11425 & n11435;
  assign n11437 = ~n11422 & n11436;
  assign n11438 = pi050 & ~pi085;
  assign n11439 = ~pi092 & n11438;
  assign n11440 = ~n3458 & ~n11439;
  assign n11441 = ~pi089 & ~n11440;
  assign n11442 = pi085 & n3575;
  assign n11443 = n3433 & n11442;
  assign n11444 = pi092 & n3431;
  assign n11445 = ~n11443 & ~n11444;
  assign n11446 = ~pi089 & ~n11445;
  assign n11447 = ~n11441 & ~n11446;
  assign n11448 = n11437 & n11447;
  assign n11449 = ~pi053 & ~n11448;
  assign n11450 = ~n11419 & ~n11449;
  assign n11451 = n11379 & n11450;
  assign n11452 = ~n11362 & n11451;
  assign n11453 = n8206 & ~n11405;
  assign n11454 = ~pi092 & ~n11453;
  assign n11455 = n3482 & n8199;
  assign n11456 = ~pi028 & n3478;
  assign n11457 = ~n3495 & ~n11456;
  assign n11458 = ~n11442 & n11457;
  assign n11459 = pi092 & ~n11458;
  assign n11460 = ~n3496 & ~n3500;
  assign n11461 = ~n8156 & n11460;
  assign n11462 = ~n11459 & n11461;
  assign n11463 = ~n8236 & ~n11408;
  assign n11464 = n11462 & n11463;
  assign n11465 = pi089 & ~n11464;
  assign n11466 = ~n11455 & ~n11465;
  assign n11467 = ~n11454 & n11466;
  assign n11468 = ~n3455 & ~n3503;
  assign n11469 = ~pi092 & ~n11468;
  assign n11470 = pi092 & n3482;
  assign n11471 = pi092 & n8171;
  assign n11472 = ~n11470 & ~n11471;
  assign n11473 = ~n8231 & n11472;
  assign n11474 = ~n11469 & n11473;
  assign n11475 = ~n3438 & ~n8248;
  assign n11476 = n11474 & n11475;
  assign n11477 = ~n3428 & n11476;
  assign n11478 = ~pi089 & ~n11477;
  assign n11479 = n11467 & ~n11478;
  assign n11480 = ~n3426 & ~n3454;
  assign n11481 = pi085 & ~n11480;
  assign n11482 = ~n3552 & ~n11481;
  assign n11483 = pi092 & ~n11482;
  assign n11484 = n11479 & ~n11483;
  assign n11485 = pi053 & ~n11484;
  assign n11486 = ~pi092 & n3559;
  assign n11487 = ~pi028 & n8162;
  assign n11488 = ~pi050 & ~pi087;
  assign n11489 = ~pi085 & n11488;
  assign n11490 = ~n11487 & ~n11489;
  assign n11491 = pi092 & ~n11490;
  assign n11492 = ~pi028 & n3493;
  assign n11493 = ~n8230 & ~n11492;
  assign n11494 = ~n3573 & n11493;
  assign n11495 = ~n11491 & n11494;
  assign n11496 = ~n11486 & n11495;
  assign n11497 = pi089 & ~n11496;
  assign n11498 = pi092 & n3493;
  assign n11499 = n3433 & n11489;
  assign n11500 = pi028 & n8254;
  assign n11501 = ~n3442 & ~n11500;
  assign n11502 = ~pi092 & ~n11501;
  assign n11503 = ~pi028 & n3553;
  assign n11504 = ~n11502 & ~n11503;
  assign n11505 = ~n11499 & n11504;
  assign n11506 = ~n11498 & n11505;
  assign n11507 = n3488 & n3496;
  assign n11508 = ~n3460 & ~n11405;
  assign n11509 = ~n3439 & ~n3456;
  assign n11510 = n3508 & ~n11509;
  assign n11511 = pi092 & n8189;
  assign n11512 = ~n11510 & ~n11511;
  assign n11513 = n11508 & n11512;
  assign n11514 = ~n11507 & n11513;
  assign n11515 = ~pi089 & ~n11514;
  assign n11516 = n11506 & ~n11515;
  assign n11517 = ~n11497 & n11516;
  assign n11518 = ~pi053 & ~n11517;
  assign n11519 = pi028 & n11349;
  assign n11520 = ~pi089 & ~pi092;
  assign n11521 = n11519 & n11520;
  assign n11522 = ~n3510 & ~n11521;
  assign n11523 = n3433 & n3470;
  assign n11524 = ~n3429 & ~n11523;
  assign n11525 = n3471 & n8199;
  assign n11526 = ~n3500 & ~n11525;
  assign n11527 = pi092 & ~n11526;
  assign n11528 = n3488 & n8144;
  assign n11529 = pi092 & n3496;
  assign n11530 = ~n11528 & ~n11529;
  assign n11531 = ~n3559 & ~n11384;
  assign n11532 = ~n3515 & n11531;
  assign n11533 = n8174 & ~n11532;
  assign n11534 = n11530 & ~n11533;
  assign n11535 = ~n11527 & n11534;
  assign n11536 = pi089 & ~n11535;
  assign n11537 = pi092 & n3461;
  assign n11538 = n3508 & n3553;
  assign n11539 = ~n11537 & ~n11538;
  assign n11540 = ~pi089 & ~n11539;
  assign n11541 = ~n11536 & ~n11540;
  assign n11542 = n11524 & n11541;
  assign n11543 = n11522 & n11542;
  assign n11544 = ~n11518 & n11543;
  assign n11545 = ~n11485 & n11544;
  assign n11546 = ~n11452 & n11545;
  assign n11547 = n11452 & ~n11545;
  assign n11548 = ~n11546 & ~n11547;
  assign n11549 = ~pi067 & n3860;
  assign n11550 = ~n3798 & ~n11549;
  assign n11551 = pi117 & ~n11550;
  assign n11552 = pi117 & n3788;
  assign n11553 = ~n3918 & ~n11552;
  assign n11554 = ~pi002 & ~n11553;
  assign n11555 = pi067 & n3830;
  assign n11556 = pi002 & n11555;
  assign n11557 = ~n4022 & ~n11556;
  assign n11558 = ~n11554 & n11557;
  assign n11559 = n3897 & n3916;
  assign n11560 = pi117 & n3794;
  assign n11561 = ~n11559 & ~n11560;
  assign n11562 = pi002 & ~n11561;
  assign n11563 = ~pi117 & n3888;
  assign n11564 = ~n11562 & ~n11563;
  assign n11565 = n11558 & n11564;
  assign n11566 = ~n11551 & n11565;
  assign n11567 = ~pi067 & n3889;
  assign n11568 = ~n3929 & ~n11567;
  assign n11569 = ~n3964 & n11568;
  assign n11570 = pi002 & ~pi117;
  assign n11571 = ~n11569 & n11570;
  assign n11572 = n3794 & n3873;
  assign n11573 = pi067 & n3952;
  assign n11574 = ~n11572 & ~n11573;
  assign n11575 = ~pi002 & ~n11574;
  assign n11576 = ~n11571 & ~n11575;
  assign n11577 = n11566 & n11576;
  assign n11578 = ~pi036 & ~n11577;
  assign n11579 = pi117 & n3831;
  assign n11580 = n3781 & n3949;
  assign n11581 = ~n3786 & ~n11580;
  assign n11582 = ~n3770 & ~n3859;
  assign n11583 = pi067 & ~n11582;
  assign n11584 = ~pi067 & n3807;
  assign n11585 = ~n11583 & ~n11584;
  assign n11586 = ~n4018 & n11585;
  assign n11587 = ~pi117 & ~n11586;
  assign n11588 = ~n3965 & ~n11587;
  assign n11589 = n11581 & n11588;
  assign n11590 = ~n11579 & n11589;
  assign n11591 = pi002 & ~n11590;
  assign n11592 = ~n3975 & ~n4017;
  assign n11593 = n3822 & ~n11592;
  assign n11594 = ~pi067 & n3811;
  assign n11595 = ~n11593 & ~n11594;
  assign n11596 = ~n3815 & n11595;
  assign n11597 = ~n3847 & n11596;
  assign n11598 = pi117 & ~n11597;
  assign n11599 = ~pi067 & n3898;
  assign n11600 = pi067 & n3807;
  assign n11601 = ~n11599 & ~n11600;
  assign n11602 = ~pi067 & n3784;
  assign n11603 = n11601 & ~n11602;
  assign n11604 = ~pi117 & ~n11603;
  assign n11605 = ~n3903 & ~n11604;
  assign n11606 = ~n11598 & n11605;
  assign n11607 = ~n4022 & n11606;
  assign n11608 = ~pi002 & ~n11607;
  assign n11609 = ~n11591 & ~n11608;
  assign n11610 = ~n11578 & n11609;
  assign n11611 = ~pi117 & n3806;
  assign n11612 = ~n11552 & ~n11611;
  assign n11613 = pi067 & ~n11612;
  assign n11614 = pi117 & n3982;
  assign n11615 = ~pi032 & n3793;
  assign n11616 = ~n3823 & ~n11615;
  assign n11617 = ~pi117 & ~n11616;
  assign n11618 = ~n4010 & ~n11617;
  assign n11619 = ~n11614 & n11618;
  assign n11620 = n3782 & n3857;
  assign n11621 = n11619 & ~n11620;
  assign n11622 = pi002 & ~n11621;
  assign n11623 = ~pi067 & ~pi105;
  assign n11624 = pi032 & n11623;
  assign n11625 = ~n3807 & ~n11624;
  assign n11626 = ~pi032 & n3892;
  assign n11627 = ~n4008 & ~n11626;
  assign n11628 = n11625 & n11627;
  assign n11629 = pi117 & ~n11628;
  assign n11630 = pi067 & n3784;
  assign n11631 = pi067 & n11615;
  assign n11632 = ~n4018 & ~n11631;
  assign n11633 = ~n11630 & n11632;
  assign n11634 = ~pi117 & ~n11633;
  assign n11635 = ~n11629 & ~n11634;
  assign n11636 = ~pi117 & n3912;
  assign n11637 = pi067 & n3818;
  assign n11638 = pi067 & n3775;
  assign n11639 = ~n3942 & ~n11638;
  assign n11640 = ~n11637 & n11639;
  assign n11641 = ~n11636 & n11640;
  assign n11642 = pi117 & n3929;
  assign n11643 = n11641 & ~n11642;
  assign n11644 = ~pi002 & ~n11643;
  assign n11645 = n11635 & ~n11644;
  assign n11646 = ~n11622 & n11645;
  assign n11647 = pi036 & ~n11646;
  assign n11648 = ~n11613 & ~n11647;
  assign n11649 = n11610 & n11648;
  assign n11650 = pi115 & n4135;
  assign n11651 = pi095 & n3609;
  assign n11652 = n3593 & n11651;
  assign n11653 = ~n11650 & ~n11652;
  assign n11654 = pi026 & ~n11653;
  assign n11655 = ~n3654 & ~n3656;
  assign n11656 = pi008 & ~n11655;
  assign n11657 = ~pi008 & n3671;
  assign n11658 = ~n11656 & ~n11657;
  assign n11659 = ~n4154 & n11658;
  assign n11660 = ~pi115 & ~n11659;
  assign n11661 = ~n4080 & ~n11660;
  assign n11662 = ~n4180 & n11661;
  assign n11663 = pi026 & ~n11662;
  assign n11664 = ~n3607 & ~n4120;
  assign n11665 = ~n3721 & ~n4208;
  assign n11666 = ~n3684 & n11665;
  assign n11667 = n11664 & n11666;
  assign n11668 = pi115 & ~n11667;
  assign n11669 = ~pi008 & n3655;
  assign n11670 = ~n3672 & ~n11669;
  assign n11671 = ~n3649 & n11670;
  assign n11672 = ~pi115 & ~n11671;
  assign n11673 = ~n11668 & ~n11672;
  assign n11674 = ~n4249 & n11673;
  assign n11675 = ~n4132 & n11674;
  assign n11676 = ~pi026 & ~n11675;
  assign n11677 = pi008 & n4134;
  assign n11678 = pi115 & n3620;
  assign n11679 = ~n11677 & ~n11678;
  assign n11680 = ~n3703 & ~n4079;
  assign n11681 = ~pi008 & n3622;
  assign n11682 = n11680 & ~n11681;
  assign n11683 = ~pi115 & ~n11682;
  assign n11684 = n4235 & n4258;
  assign n11685 = ~n11683 & ~n11684;
  assign n11686 = n11679 & n11685;
  assign n11687 = pi026 & ~n11686;
  assign n11688 = ~pi115 & n3632;
  assign n11689 = pi008 & n3594;
  assign n11690 = ~n4237 & ~n11689;
  assign n11691 = pi115 & n3730;
  assign n11692 = ~pi115 & n3621;
  assign n11693 = ~n11691 & ~n11692;
  assign n11694 = n11690 & n11693;
  assign n11695 = ~pi026 & ~n11694;
  assign n11696 = ~n11688 & ~n11695;
  assign n11697 = ~n11687 & n11696;
  assign n11698 = ~pi008 & n4212;
  assign n11699 = ~n4177 & ~n11698;
  assign n11700 = pi115 & ~n11699;
  assign n11701 = ~n4132 & ~n11700;
  assign n11702 = n11697 & n11701;
  assign n11703 = ~pi030 & ~n11702;
  assign n11704 = ~n11676 & ~n11703;
  assign n11705 = ~n11663 & n11704;
  assign n11706 = ~n11654 & n11705;
  assign n11707 = pi115 & n3729;
  assign n11708 = n3639 & n11707;
  assign n11709 = pi008 & ~pi115;
  assign n11710 = n3626 & n11709;
  assign n11711 = ~n11708 & ~n11710;
  assign n11712 = ~pi056 & n4060;
  assign n11713 = ~n4145 & ~n11712;
  assign n11714 = pi115 & ~n11713;
  assign n11715 = pi008 & n3694;
  assign n11716 = ~n4073 & ~n11715;
  assign n11717 = ~pi115 & n3743;
  assign n11718 = pi008 & n4169;
  assign n11719 = ~n11717 & ~n11718;
  assign n11720 = n11716 & n11719;
  assign n11721 = pi115 & n3703;
  assign n11722 = n11720 & ~n11721;
  assign n11723 = ~pi026 & ~n11722;
  assign n11724 = ~n3747 & ~n4152;
  assign n11725 = pi115 & n4097;
  assign n11726 = ~n3606 & ~n3682;
  assign n11727 = ~pi115 & ~n11726;
  assign n11728 = ~n11725 & ~n11727;
  assign n11729 = n11724 & n11728;
  assign n11730 = pi026 & ~n11729;
  assign n11731 = ~n11723 & ~n11730;
  assign n11732 = ~pi008 & ~pi099;
  assign n11733 = pi059 & n11732;
  assign n11734 = ~n3671 & ~n11733;
  assign n11735 = pi115 & ~n11734;
  assign n11736 = ~n3674 & ~n3683;
  assign n11737 = ~n4154 & n11736;
  assign n11738 = ~pi115 & ~n11737;
  assign n11739 = ~n11735 & ~n11738;
  assign n11740 = n11731 & n11739;
  assign n11741 = ~n11714 & n11740;
  assign n11742 = pi030 & ~n11741;
  assign n11743 = n11711 & ~n11742;
  assign n11744 = n11706 & n11743;
  assign n11745 = ~n11649 & n11744;
  assign n11746 = n11649 & ~n11744;
  assign n11747 = ~n11745 & ~n11746;
  assign n11748 = ~n11548 & n11747;
  assign n11749 = n11548 & ~n11747;
  assign n11750 = ~n11748 & ~n11749;
  assign n11751 = ~pi080 & n3261;
  assign n11752 = ~pi075 & n3279;
  assign n11753 = ~pi110 & n3366;
  assign n11754 = n3263 & n11753;
  assign n11755 = pi079 & n3291;
  assign n11756 = ~n8075 & ~n11755;
  assign n11757 = pi080 & n3264;
  assign n11758 = n11756 & ~n11757;
  assign n11759 = ~n11754 & n11758;
  assign n11760 = ~pi073 & ~n11759;
  assign n11761 = ~n11752 & ~n11760;
  assign n11762 = ~pi075 & n3297;
  assign n11763 = ~pi079 & n3326;
  assign n11764 = ~n11762 & ~n11763;
  assign n11765 = ~n3365 & n11764;
  assign n11766 = ~pi080 & ~n11765;
  assign n11767 = pi080 & n3272;
  assign n11768 = pi079 & n8033;
  assign n11769 = ~n11767 & ~n11768;
  assign n11770 = n3401 & n8073;
  assign n11771 = n11769 & ~n11770;
  assign n11772 = ~n11766 & n11771;
  assign n11773 = pi073 & ~n11772;
  assign n11774 = ~pi079 & n8059;
  assign n11775 = ~n8120 & ~n11774;
  assign n11776 = pi080 & ~n11775;
  assign n11777 = ~n11773 & ~n11776;
  assign n11778 = n11761 & n11777;
  assign n11779 = ~n11751 & n11778;
  assign n11780 = ~pi015 & ~n11779;
  assign n11781 = pi079 & n3329;
  assign n11782 = ~pi080 & n11781;
  assign n11783 = n3264 & n3288;
  assign n11784 = ~n11782 & ~n11783;
  assign n11785 = n3270 & n3395;
  assign n11786 = ~n3350 & ~n3352;
  assign n11787 = pi079 & ~n11786;
  assign n11788 = ~pi079 & n3368;
  assign n11789 = ~n11787 & ~n11788;
  assign n11790 = ~n11785 & n11789;
  assign n11791 = ~pi080 & ~n11790;
  assign n11792 = pi079 & n11762;
  assign n11793 = pi080 & n8034;
  assign n11794 = ~n11792 & ~n11793;
  assign n11795 = ~n11791 & n11794;
  assign n11796 = pi080 & n8112;
  assign n11797 = ~n8065 & ~n11796;
  assign n11798 = n11795 & n11797;
  assign n11799 = pi073 & ~n11798;
  assign n11800 = n11784 & ~n11799;
  assign n11801 = pi079 & n8130;
  assign n11802 = ~n3317 & ~n11801;
  assign n11803 = ~pi075 & n3296;
  assign n11804 = pi080 & n11803;
  assign n11805 = ~n3374 & ~n8132;
  assign n11806 = ~pi080 & ~n11805;
  assign n11807 = ~n11804 & ~n11806;
  assign n11808 = n11802 & n11807;
  assign n11809 = pi073 & ~n11808;
  assign n11810 = ~n3375 & ~n3392;
  assign n11811 = ~n11785 & n11810;
  assign n11812 = ~pi080 & ~n11811;
  assign n11813 = n3269 & n3302;
  assign n11814 = ~pi080 & n11813;
  assign n11815 = pi079 & n3312;
  assign n11816 = ~n11814 & ~n11815;
  assign n11817 = ~pi080 & n3313;
  assign n11818 = pi079 & n8052;
  assign n11819 = ~n11817 & ~n11818;
  assign n11820 = n11816 & n11819;
  assign n11821 = pi080 & n3365;
  assign n11822 = n11820 & ~n11821;
  assign n11823 = ~pi073 & ~n11822;
  assign n11824 = ~n11812 & ~n11823;
  assign n11825 = ~n11809 & n11824;
  assign n11826 = ~pi075 & pi079;
  assign n11827 = ~pi042 & n11826;
  assign n11828 = pi079 & n3297;
  assign n11829 = ~n11827 & ~n11828;
  assign n11830 = pi080 & ~n11829;
  assign n11831 = ~pi110 & n8061;
  assign n11832 = ~n3368 & ~n11831;
  assign n11833 = pi080 & ~n11832;
  assign n11834 = ~n11830 & ~n11833;
  assign n11835 = n11825 & n11834;
  assign n11836 = pi015 & ~n11835;
  assign n11837 = ~n3302 & ~n3395;
  assign n11838 = n3297 & ~n11837;
  assign n11839 = ~n3372 & ~n8041;
  assign n11840 = ~n11838 & n11839;
  assign n11841 = ~n3279 & n11840;
  assign n11842 = pi080 & ~n11841;
  assign n11843 = ~n8082 & ~n11752;
  assign n11844 = ~pi079 & n3351;
  assign n11845 = ~n3369 & ~n11844;
  assign n11846 = ~n3348 & n11845;
  assign n11847 = ~pi080 & ~n11846;
  assign n11848 = n11843 & ~n11847;
  assign n11849 = ~n11842 & n11848;
  assign n11850 = ~pi073 & ~n11849;
  assign n11851 = ~n11836 & ~n11850;
  assign n11852 = n11800 & n11851;
  assign n11853 = ~n11780 & n11852;
  assign n11854 = ~pi301 & ~n11853;
  assign n11855 = pi301 & n11853;
  assign n11856 = ~n11854 & ~n11855;
  assign n11857 = ~pi079 & n3353;
  assign n11858 = pi079 & n3293;
  assign n11859 = ~pi079 & n3365;
  assign n11860 = ~n11858 & ~n11859;
  assign n11861 = ~n11857 & n11860;
  assign n11862 = ~pi080 & ~n11861;
  assign n11863 = pi079 & n3273;
  assign n11864 = ~pi079 & n3275;
  assign n11865 = ~n3326 & ~n11864;
  assign n11866 = ~n8073 & n11865;
  assign n11867 = pi080 & ~n11866;
  assign n11868 = ~pi080 & n3270;
  assign n11869 = ~n3365 & ~n3392;
  assign n11870 = ~n11868 & n11869;
  assign n11871 = ~n11867 & n11870;
  assign n11872 = ~n8039 & ~n8109;
  assign n11873 = n11871 & n11872;
  assign n11874 = pi073 & ~n11873;
  assign n11875 = ~n11863 & ~n11874;
  assign n11876 = ~n11862 & n11875;
  assign n11877 = pi080 & n8078;
  assign n11878 = n3283 & n3310;
  assign n11879 = pi080 & n11828;
  assign n11880 = ~n11767 & ~n11879;
  assign n11881 = ~n11878 & n11880;
  assign n11882 = ~n11877 & n11881;
  assign n11883 = n3259 & n3366;
  assign n11884 = n3263 & n3395;
  assign n11885 = ~n3292 & ~n11884;
  assign n11886 = ~n3303 & n11885;
  assign n11887 = ~n11883 & n11886;
  assign n11888 = n11882 & n11887;
  assign n11889 = ~pi073 & ~n11888;
  assign n11890 = n11876 & ~n11889;
  assign n11891 = ~n3297 & ~n3310;
  assign n11892 = pi075 & ~n11891;
  assign n11893 = ~n3338 & ~n11892;
  assign n11894 = pi080 & ~n11893;
  assign n11895 = n11890 & ~n11894;
  assign n11896 = pi015 & ~n11895;
  assign n11897 = ~pi080 & n3333;
  assign n11898 = ~n11788 & ~n11828;
  assign n11899 = ~pi071 & ~pi110;
  assign n11900 = ~pi075 & n11899;
  assign n11901 = ~pi079 & n8051;
  assign n11902 = ~n11900 & ~n11901;
  assign n11903 = pi080 & ~n11902;
  assign n11904 = ~n3358 & ~n11903;
  assign n11905 = n11898 & n11904;
  assign n11906 = ~n11897 & n11905;
  assign n11907 = pi073 & ~n11906;
  assign n11908 = n3283 & n3365;
  assign n11909 = ~n3316 & ~n11857;
  assign n11910 = pi075 & n3269;
  assign n11911 = pi080 & n11910;
  assign n11912 = ~n3258 & ~n3312;
  assign n11913 = n3401 & ~n11912;
  assign n11914 = ~n11911 & ~n11913;
  assign n11915 = n11909 & n11914;
  assign n11916 = ~n11908 & n11915;
  assign n11917 = ~pi073 & ~n11916;
  assign n11918 = ~n11907 & ~n11917;
  assign n11919 = ~pi079 & n3329;
  assign n11920 = pi080 & n3368;
  assign n11921 = ~n3295 & ~n11768;
  assign n11922 = ~pi080 & ~n11921;
  assign n11923 = n3288 & n11900;
  assign n11924 = ~n11922 & ~n11923;
  assign n11925 = ~n11920 & n11924;
  assign n11926 = ~n11919 & n11925;
  assign n11927 = n11918 & n11926;
  assign n11928 = ~pi015 & ~n11927;
  assign n11929 = n3263 & n11826;
  assign n11930 = ~n3392 & ~n11929;
  assign n11931 = pi080 & ~n11930;
  assign n11932 = ~n3333 & ~n8025;
  assign n11933 = ~n3374 & n11932;
  assign n11934 = n3366 & ~n11933;
  assign n11935 = ~n11931 & ~n11934;
  assign n11936 = ~pi080 & n11792;
  assign n11937 = n11935 & ~n11936;
  assign n11938 = ~n11821 & n11937;
  assign n11939 = pi073 & ~n11938;
  assign n11940 = n3262 & n3288;
  assign n11941 = ~n3304 & ~n11940;
  assign n11942 = ~n3403 & n11941;
  assign n11943 = ~pi080 & n11818;
  assign n11944 = ~pi073 & n11943;
  assign n11945 = n11942 & ~n11944;
  assign n11946 = ~n11939 & n11945;
  assign n11947 = pi080 & n3317;
  assign n11948 = n3329 & n3401;
  assign n11949 = ~n11947 & ~n11948;
  assign n11950 = ~pi073 & ~n11949;
  assign n11951 = n11946 & ~n11950;
  assign n11952 = ~n11928 & n11951;
  assign n11953 = ~n11896 & n11952;
  assign n11954 = ~n8140 & n11953;
  assign n11955 = n8140 & ~n11953;
  assign n11956 = ~n11954 & ~n11955;
  assign n11957 = ~n11856 & ~n11956;
  assign n11958 = n11856 & n11956;
  assign n11959 = ~n11957 & ~n11958;
  assign n11960 = ~n11750 & n11959;
  assign n11961 = n11750 & ~n11959;
  assign n11962 = ~n11960 & ~n11961;
  assign n11963 = ~pi529 & n11962;
  assign po166 = n11347 | n11963;
  assign n11965 = pi184 & pi442;
  assign n11966 = ~pi184 & ~pi442;
  assign n11967 = ~n11965 & ~n11966;
  assign n11968 = pi529 & ~n11967;
  assign n11969 = ~n3597 & ~n3625;
  assign n11970 = pi059 & ~n11969;
  assign n11971 = ~n3638 & ~n11970;
  assign n11972 = pi115 & ~n11971;
  assign n11973 = ~n4138 & ~n11972;
  assign n11974 = ~n3704 & ~n4067;
  assign n11975 = ~n4201 & n11974;
  assign n11976 = ~pi115 & ~n11975;
  assign n11977 = ~pi008 & n3718;
  assign n11978 = ~n3622 & ~n11977;
  assign n11979 = ~n4235 & n11978;
  assign n11980 = pi115 & ~n11979;
  assign n11981 = ~n3736 & ~n11980;
  assign n11982 = ~n3674 & ~n4204;
  assign n11983 = ~n3703 & n11982;
  assign n11984 = ~n4190 & n11983;
  assign n11985 = n11981 & n11984;
  assign n11986 = pi026 & ~n11985;
  assign n11987 = ~n11976 & ~n11986;
  assign n11988 = n11973 & n11987;
  assign n11989 = ~n3649 & ~n3742;
  assign n11990 = ~pi115 & ~n11989;
  assign n11991 = pi115 & n4100;
  assign n11992 = ~n11678 & ~n11991;
  assign n11993 = ~n4146 & n11992;
  assign n11994 = ~n11990 & n11993;
  assign n11995 = ~n3595 & ~n4122;
  assign n11996 = n11994 & n11995;
  assign n11997 = ~n3607 & n11996;
  assign n11998 = ~pi026 & ~n11997;
  assign n11999 = n11988 & ~n11998;
  assign n12000 = pi030 & ~n11999;
  assign n12001 = ~pi115 & n3633;
  assign n12002 = ~n3652 & ~n12001;
  assign n12003 = ~n4145 & ~n11657;
  assign n12004 = ~pi008 & n4104;
  assign n12005 = ~pi095 & ~pi099;
  assign n12006 = ~pi059 & n12005;
  assign n12007 = ~n12004 & ~n12006;
  assign n12008 = pi115 & ~n12007;
  assign n12009 = n12003 & ~n12008;
  assign n12010 = n12002 & n12009;
  assign n12011 = pi026 & n12010;
  assign n12012 = pi115 & n3593;
  assign n12013 = pi059 & n12012;
  assign n12014 = ~n3600 & ~n3694;
  assign n12015 = n4258 & ~n12014;
  assign n12016 = ~n4201 & ~n12015;
  assign n12017 = ~n3746 & n12016;
  assign n12018 = n3703 & n11709;
  assign n12019 = n12017 & ~n12018;
  assign n12020 = ~n12013 & n12019;
  assign n12021 = ~pi026 & n12020;
  assign n12022 = ~n12011 & ~n12021;
  assign n12023 = ~n3603 & ~n11677;
  assign n12024 = ~pi115 & ~n12023;
  assign n12025 = ~pi008 & n3626;
  assign n12026 = ~n12024 & ~n12025;
  assign n12027 = pi115 & n3671;
  assign n12028 = n3609 & n12006;
  assign n12029 = ~n12027 & ~n12028;
  assign n12030 = n12026 & n12029;
  assign n12031 = ~n12022 & n12030;
  assign n12032 = ~pi030 & ~n12031;
  assign n12033 = pi115 & n3747;
  assign n12034 = n3626 & n4258;
  assign n12035 = ~n12033 & ~n12034;
  assign n12036 = ~pi026 & ~n12035;
  assign n12037 = n3609 & n3651;
  assign n12038 = ~n3608 & ~n12037;
  assign n12039 = ~n12036 & n12038;
  assign n12040 = ~n3673 & n12039;
  assign n12041 = ~pi026 & ~pi115;
  assign n12042 = n11718 & n12041;
  assign n12043 = ~pi115 & n4080;
  assign n12044 = ~n11721 & ~n12043;
  assign n12045 = ~n3633 & ~n3682;
  assign n12046 = ~n4196 & n12045;
  assign n12047 = n4049 & ~n12046;
  assign n12048 = n12044 & ~n12047;
  assign n12049 = pi026 & ~n12048;
  assign n12050 = ~n12042 & ~n12049;
  assign n12051 = n3729 & n4060;
  assign n12052 = ~n3674 & ~n12051;
  assign n12053 = n3728 & ~n12052;
  assign n12054 = n12050 & ~n12053;
  assign n12055 = n12040 & n12054;
  assign n12056 = ~n12032 & n12055;
  assign n12057 = ~n12000 & n12056;
  assign n12058 = n4267 & n12057;
  assign n12059 = ~n4267 & ~n12057;
  assign n12060 = ~n12058 & ~n12059;
  assign n12061 = n3794 & n3935;
  assign n12062 = ~pi067 & n3803;
  assign n12063 = ~n3889 & ~n12062;
  assign n12064 = ~n3916 & n12063;
  assign n12065 = pi117 & ~n12064;
  assign n12066 = ~n3929 & ~n11630;
  assign n12067 = ~n3969 & n12066;
  assign n12068 = ~n12065 & n12067;
  assign n12069 = ~n3777 & ~n3842;
  assign n12070 = n12068 & n12069;
  assign n12071 = pi002 & ~n12070;
  assign n12072 = ~n3839 & ~n3930;
  assign n12073 = ~n3931 & n12072;
  assign n12074 = ~pi117 & ~n12073;
  assign n12075 = ~n3805 & ~n3822;
  assign n12076 = pi032 & ~n12075;
  assign n12077 = pi067 & n3821;
  assign n12078 = pi032 & n12077;
  assign n12079 = ~n12076 & ~n12078;
  assign n12080 = pi117 & ~n12079;
  assign n12081 = ~n12074 & ~n12080;
  assign n12082 = pi117 & n3763;
  assign n12083 = ~n11560 & ~n12082;
  assign n12084 = ~n3894 & ~n11602;
  assign n12085 = ~pi117 & ~n12084;
  assign n12086 = n3822 & n3975;
  assign n12087 = ~n12085 & ~n12086;
  assign n12088 = ~n4009 & n12087;
  assign n12089 = n12083 & n12088;
  assign n12090 = ~pi067 & n3952;
  assign n12091 = ~n4030 & ~n12090;
  assign n12092 = n12089 & n12091;
  assign n12093 = ~pi002 & ~n12092;
  assign n12094 = n12081 & ~n12093;
  assign n12095 = ~n12071 & n12094;
  assign n12096 = ~n12061 & n12095;
  assign n12097 = pi036 & ~n12096;
  assign n12098 = ~pi002 & ~pi117;
  assign n12099 = n11637 & n12098;
  assign n12100 = ~pi117 & n3965;
  assign n12101 = ~n11642 & ~n12100;
  assign n12102 = ~pi032 & n3889;
  assign n12103 = ~n3834 & ~n12102;
  assign n12104 = ~n11615 & n12103;
  assign n12105 = n3873 & ~n12104;
  assign n12106 = n12101 & ~n12105;
  assign n12107 = pi002 & ~n12106;
  assign n12108 = ~n12099 & ~n12107;
  assign n12109 = pi117 & n11620;
  assign n12110 = n3806 & n3897;
  assign n12111 = ~n12109 & ~n12110;
  assign n12112 = ~pi002 & ~n12111;
  assign n12113 = n3823 & n3861;
  assign n12114 = pi067 & n3816;
  assign n12115 = pi117 & n12114;
  assign n12116 = ~n12113 & ~n12115;
  assign n12117 = n3805 & n3975;
  assign n12118 = n12116 & ~n12117;
  assign n12119 = n3787 & n3935;
  assign n12120 = ~n11630 & ~n12119;
  assign n12121 = n3865 & ~n12120;
  assign n12122 = n12118 & ~n12121;
  assign n12123 = ~n12112 & n12122;
  assign n12124 = n12108 & n12123;
  assign n12125 = ~n3797 & ~n3839;
  assign n12126 = ~n3765 & ~n3775;
  assign n12127 = n3897 & ~n12126;
  assign n12128 = pi117 & n3940;
  assign n12129 = ~n12127 & ~n12128;
  assign n12130 = pi067 & ~pi117;
  assign n12131 = n3929 & n12130;
  assign n12132 = n12129 & ~n12131;
  assign n12133 = n12125 & n12132;
  assign n12134 = ~pi002 & ~n12133;
  assign n12135 = ~pi067 & n3806;
  assign n12136 = ~pi067 & n3883;
  assign n12137 = ~n11555 & ~n12136;
  assign n12138 = ~pi117 & ~n12137;
  assign n12139 = pi117 & n3807;
  assign n12140 = ~pi064 & ~pi105;
  assign n12141 = ~pi032 & n12140;
  assign n12142 = n3861 & n12141;
  assign n12143 = ~n12139 & ~n12142;
  assign n12144 = ~n12138 & n12143;
  assign n12145 = ~n12135 & n12144;
  assign n12146 = ~n12134 & n12145;
  assign n12147 = ~pi117 & n12102;
  assign n12148 = ~pi067 & n3854;
  assign n12149 = ~n12141 & ~n12148;
  assign n12150 = pi117 & ~n12149;
  assign n12151 = ~n4008 & ~n11584;
  assign n12152 = pi067 & n3883;
  assign n12153 = n12151 & ~n12152;
  assign n12154 = ~n12150 & n12153;
  assign n12155 = ~n12147 & n12154;
  assign n12156 = pi002 & ~n12155;
  assign n12157 = n12146 & ~n12156;
  assign n12158 = ~pi036 & ~n12157;
  assign n12159 = n12124 & ~n12158;
  assign n12160 = ~n12097 & n12159;
  assign n12161 = ~n3926 & n12160;
  assign n12162 = n3926 & ~n12160;
  assign n12163 = ~n12161 & ~n12162;
  assign n12164 = n12060 & n12163;
  assign n12165 = ~n12060 & ~n12163;
  assign n12166 = ~n12164 & ~n12165;
  assign n12167 = pi092 & n8255;
  assign n12168 = ~n3526 & ~n3575;
  assign n12169 = pi028 & ~n12168;
  assign n12170 = ~n11492 & ~n12169;
  assign n12171 = ~n8241 & n12170;
  assign n12172 = ~pi092 & ~n12171;
  assign n12173 = pi092 & n11358;
  assign n12174 = ~n11363 & ~n12173;
  assign n12175 = ~n8145 & n12174;
  assign n12176 = ~n12172 & n12175;
  assign n12177 = ~n12167 & n12176;
  assign n12178 = pi089 & ~n12177;
  assign n12179 = ~pi092 & n3469;
  assign n12180 = ~pi028 & n3495;
  assign n12181 = ~n8144 & ~n12180;
  assign n12182 = ~n3496 & n12181;
  assign n12183 = ~pi092 & ~n12182;
  assign n12184 = ~n11470 & ~n11500;
  assign n12185 = n3508 & n11442;
  assign n12186 = n12184 & ~n12185;
  assign n12187 = ~n12183 & n12186;
  assign n12188 = pi089 & ~n12187;
  assign n12189 = pi028 & n8212;
  assign n12190 = ~n11444 & ~n12189;
  assign n12191 = pi092 & n3472;
  assign n12192 = ~pi092 & n3565;
  assign n12193 = ~n12191 & ~n12192;
  assign n12194 = n12190 & n12193;
  assign n12195 = ~pi089 & ~n12194;
  assign n12196 = ~pi028 & n11392;
  assign n12197 = ~n11375 & ~n12196;
  assign n12198 = pi092 & ~n12197;
  assign n12199 = ~n12195 & ~n12198;
  assign n12200 = ~n12188 & n12199;
  assign n12201 = ~n12179 & n12200;
  assign n12202 = ~n8252 & n12201;
  assign n12203 = ~pi053 & ~n12202;
  assign n12204 = ~n12178 & ~n12203;
  assign n12205 = ~pi028 & n3527;
  assign n12206 = ~n3494 & ~n12205;
  assign n12207 = ~n3503 & n12206;
  assign n12208 = ~pi092 & ~n12207;
  assign n12209 = ~n3428 & ~n8247;
  assign n12210 = ~n3481 & ~n11412;
  assign n12211 = ~n3517 & n12210;
  assign n12212 = n12209 & n12211;
  assign n12213 = pi092 & ~n12212;
  assign n12214 = ~n8252 & ~n11420;
  assign n12215 = ~n12213 & n12214;
  assign n12216 = ~n12208 & n12215;
  assign n12217 = ~pi089 & ~n12216;
  assign n12218 = n3433 & n3472;
  assign n12219 = pi028 & n3553;
  assign n12220 = ~pi092 & n12219;
  assign n12221 = ~n12218 & ~n12220;
  assign n12222 = ~n3461 & ~n8233;
  assign n12223 = ~n3427 & ~n3515;
  assign n12224 = ~pi092 & ~n12223;
  assign n12225 = pi092 & n8168;
  assign n12226 = ~n12224 & ~n12225;
  assign n12227 = n12222 & n12226;
  assign n12228 = pi089 & ~n12227;
  assign n12229 = ~n3516 & ~n8241;
  assign n12230 = ~n3500 & n12229;
  assign n12231 = ~pi092 & ~n12230;
  assign n12232 = ~pi085 & n11427;
  assign n12233 = ~n8230 & ~n12232;
  assign n12234 = ~pi028 & ~pi050;
  assign n12235 = pi085 & n12234;
  assign n12236 = ~n3493 & ~n12235;
  assign n12237 = n12233 & n12236;
  assign n12238 = pi092 & ~n12237;
  assign n12239 = ~n12231 & ~n12238;
  assign n12240 = pi028 & n3456;
  assign n12241 = ~n8190 & ~n12240;
  assign n12242 = ~pi092 & n3457;
  assign n12243 = ~n11519 & ~n12242;
  assign n12244 = n12241 & n12243;
  assign n12245 = ~n11529 & n12244;
  assign n12246 = ~pi089 & ~n12245;
  assign n12247 = n12239 & ~n12246;
  assign n12248 = ~n12228 & n12247;
  assign n12249 = pi053 & ~n12248;
  assign n12250 = n12221 & ~n12249;
  assign n12251 = ~n12217 & n12250;
  assign n12252 = n12204 & n12251;
  assign n12253 = n11744 & n12252;
  assign n12254 = ~n11744 & ~n12252;
  assign n12255 = ~n12253 & ~n12254;
  assign n12256 = pi184 & ~n11853;
  assign n12257 = ~pi184 & n11853;
  assign n12258 = ~n12256 & ~n12257;
  assign n12259 = ~n12255 & n12258;
  assign n12260 = n12255 & ~n12258;
  assign n12261 = ~n12259 & ~n12260;
  assign n12262 = ~n12166 & n12261;
  assign n12263 = n12166 & ~n12261;
  assign n12264 = ~n12262 & ~n12263;
  assign n12265 = ~pi529 & n12264;
  assign po167 = n11968 | n12265;
  assign n12267 = ~pi178 & pi450;
  assign n12268 = pi178 & ~pi450;
  assign n12269 = ~n12267 & ~n12268;
  assign n12270 = pi529 & n12269;
  assign n12271 = ~pi092 & n8233;
  assign n12272 = n3476 & n11487;
  assign n12273 = ~pi092 & n3503;
  assign n12274 = ~n12272 & ~n12273;
  assign n12275 = ~n3547 & n12274;
  assign n12276 = ~n12271 & n12275;
  assign n12277 = ~pi028 & n3457;
  assign n12278 = ~n11420 & ~n12277;
  assign n12279 = ~n8161 & n12278;
  assign n12280 = n11520 & ~n12279;
  assign n12281 = n3468 & ~n11480;
  assign n12282 = ~n3442 & ~n12281;
  assign n12283 = pi092 & ~n12282;
  assign n12284 = n3433 & n11355;
  assign n12285 = ~n3438 & ~n12284;
  assign n12286 = ~n12283 & n12285;
  assign n12287 = ~pi089 & ~n12286;
  assign n12288 = ~n12280 & ~n12287;
  assign n12289 = ~pi092 & n3496;
  assign n12290 = pi028 & n3432;
  assign n12291 = ~n12289 & ~n12290;
  assign n12292 = pi089 & ~n12291;
  assign n12293 = n12288 & ~n12292;
  assign n12294 = n3518 & ~n8171;
  assign n12295 = ~pi092 & ~n12294;
  assign n12296 = ~pi092 & n8161;
  assign n12297 = pi092 & n3442;
  assign n12298 = ~n12296 & ~n12297;
  assign n12299 = ~n11455 & n12298;
  assign n12300 = ~n12295 & n12299;
  assign n12301 = pi085 & n11488;
  assign n12302 = pi028 & pi087;
  assign n12303 = ~pi085 & n12302;
  assign n12304 = ~n3531 & ~n12303;
  assign n12305 = ~n12301 & n12304;
  assign n12306 = pi089 & ~n12305;
  assign n12307 = ~pi092 & n12306;
  assign n12308 = ~n3461 & ~n3497;
  assign n12309 = ~n3451 & ~n8169;
  assign n12310 = n12308 & n12309;
  assign n12311 = pi089 & ~n12310;
  assign n12312 = ~n12307 & ~n12311;
  assign n12313 = n12300 & n12312;
  assign n12314 = ~n3442 & ~n3517;
  assign n12315 = ~pi092 & n8230;
  assign n12316 = pi028 & n8189;
  assign n12317 = ~n11392 & ~n12316;
  assign n12318 = pi092 & ~n12317;
  assign n12319 = ~n12315 & ~n12318;
  assign n12320 = n12314 & n12319;
  assign n12321 = ~n11404 & n12320;
  assign n12322 = ~pi089 & ~n12321;
  assign n12323 = ~n11538 & ~n12322;
  assign n12324 = n12313 & n12323;
  assign n12325 = pi053 & ~n12324;
  assign n12326 = n3431 & n3508;
  assign n12327 = ~n11492 & ~n12326;
  assign n12328 = ~pi028 & n3427;
  assign n12329 = n3433 & n3531;
  assign n12330 = ~n12328 & ~n12329;
  assign n12331 = n12327 & n12330;
  assign n12332 = ~pi089 & ~n12331;
  assign n12333 = pi028 & n3521;
  assign n12334 = ~n8212 & ~n12333;
  assign n12335 = pi028 & n11489;
  assign n12336 = ~n8234 & ~n12335;
  assign n12337 = n12334 & n12336;
  assign n12338 = pi092 & ~n12337;
  assign n12339 = ~n3551 & ~n11395;
  assign n12340 = ~pi028 & n3515;
  assign n12341 = n12339 & ~n12340;
  assign n12342 = ~pi092 & ~n12341;
  assign n12343 = ~n3503 & ~n12333;
  assign n12344 = ~n8162 & ~n12240;
  assign n12345 = pi092 & ~n12344;
  assign n12346 = n12343 & ~n12345;
  assign n12347 = ~n12342 & n12346;
  assign n12348 = ~n3519 & ~n3559;
  assign n12349 = ~n8224 & n12348;
  assign n12350 = n12347 & n12349;
  assign n12351 = pi089 & ~n12350;
  assign n12352 = n3488 & n12301;
  assign n12353 = ~pi092 & n3470;
  assign n12354 = ~n12289 & ~n12353;
  assign n12355 = ~n3432 & n12354;
  assign n12356 = ~n12352 & n12355;
  assign n12357 = ~n12351 & n12356;
  assign n12358 = ~n12338 & n12357;
  assign n12359 = ~n12332 & n12358;
  assign n12360 = ~pi053 & ~n12359;
  assign n12361 = ~n12325 & ~n12360;
  assign n12362 = n12293 & n12361;
  assign n12363 = n12276 & n12362;
  assign n12364 = n11853 & ~n12363;
  assign n12365 = ~n11853 & n12363;
  assign n12366 = ~n12364 & ~n12365;
  assign n12367 = pi178 & n12366;
  assign n12368 = ~pi178 & ~n12366;
  assign n12369 = ~n12367 & ~n12368;
  assign n12370 = n3685 & ~n4100;
  assign n12371 = ~pi115 & ~n12370;
  assign n12372 = ~pi115 & n3631;
  assign n12373 = pi115 & n3603;
  assign n12374 = ~n12372 & ~n12373;
  assign n12375 = ~n4138 & n12374;
  assign n12376 = ~n12371 & n12375;
  assign n12377 = pi059 & n12005;
  assign n12378 = pi008 & pi095;
  assign n12379 = ~pi059 & n12378;
  assign n12380 = ~n3691 & ~n12379;
  assign n12381 = ~n12377 & n12380;
  assign n12382 = pi026 & ~n12381;
  assign n12383 = ~pi115 & n12382;
  assign n12384 = ~n3740 & ~n4098;
  assign n12385 = ~n3704 & ~n3747;
  assign n12386 = n12384 & n12385;
  assign n12387 = pi026 & ~n12386;
  assign n12388 = ~n12383 & ~n12387;
  assign n12389 = n12376 & n12388;
  assign n12390 = ~n3603 & ~n3684;
  assign n12391 = ~n4072 & ~n4212;
  assign n12392 = pi115 & ~n12391;
  assign n12393 = ~pi115 & n4145;
  assign n12394 = ~n12392 & ~n12393;
  assign n12395 = n12390 & n12394;
  assign n12396 = ~n4200 & n12395;
  assign n12397 = ~pi026 & ~n12396;
  assign n12398 = ~n12034 & ~n12397;
  assign n12399 = n12389 & n12398;
  assign n12400 = pi030 & ~n12399;
  assign n12401 = ~pi115 & n3703;
  assign n12402 = ~pi115 & n3651;
  assign n12403 = ~n12401 & ~n12402;
  assign n12404 = n11709 & n12377;
  assign n12405 = ~n3612 & ~n12404;
  assign n12406 = n12403 & n12405;
  assign n12407 = n3611 & n4258;
  assign n12408 = ~n11657 & ~n12407;
  assign n12409 = ~pi008 & n3606;
  assign n12410 = n3609 & n3691;
  assign n12411 = ~n12409 & ~n12410;
  assign n12412 = n12408 & n12411;
  assign n12413 = ~pi026 & ~n12412;
  assign n12414 = ~n3635 & ~n4215;
  assign n12415 = ~pi008 & n3682;
  assign n12416 = n12414 & ~n12415;
  assign n12417 = ~pi115 & ~n12416;
  assign n12418 = pi008 & n3695;
  assign n12419 = ~n3649 & ~n12418;
  assign n12420 = ~n4104 & ~n11715;
  assign n12421 = pi115 & ~n12420;
  assign n12422 = n12419 & ~n12421;
  assign n12423 = ~n12417 & n12422;
  assign n12424 = ~n3633 & ~n3686;
  assign n12425 = ~n4126 & n12424;
  assign n12426 = n12423 & n12425;
  assign n12427 = pi026 & ~n12426;
  assign n12428 = ~n3594 & ~n12418;
  assign n12429 = pi008 & n12006;
  assign n12430 = n3625 & n4086;
  assign n12431 = ~n12429 & ~n12430;
  assign n12432 = n12428 & n12431;
  assign n12433 = pi115 & ~n12432;
  assign n12434 = ~n12427 & ~n12433;
  assign n12435 = ~n12413 & n12434;
  assign n12436 = n12406 & n12435;
  assign n12437 = ~pi030 & ~n12436;
  assign n12438 = ~n12400 & ~n12437;
  assign n12439 = ~pi008 & n3743;
  assign n12440 = ~n4249 & ~n12439;
  assign n12441 = ~n3631 & n12440;
  assign n12442 = n12041 & ~n12441;
  assign n12443 = pi008 & n3612;
  assign n12444 = ~n12401 & ~n12443;
  assign n12445 = pi026 & ~n12444;
  assign n12446 = ~pi115 & n4152;
  assign n12447 = ~n3708 & ~n12446;
  assign n12448 = ~pi115 & n3649;
  assign n12449 = n12447 & ~n12448;
  assign n12450 = ~n12445 & n12449;
  assign n12451 = ~n12442 & n12450;
  assign n12452 = n3609 & n4162;
  assign n12453 = n4086 & ~n11969;
  assign n12454 = ~n3603 & ~n12453;
  assign n12455 = pi115 & ~n12454;
  assign n12456 = ~n12452 & ~n12455;
  assign n12457 = ~n3595 & n12456;
  assign n12458 = ~pi026 & ~n12457;
  assign n12459 = n3728 & n12004;
  assign n12460 = ~n12458 & ~n12459;
  assign n12461 = n12451 & n12460;
  assign n12462 = n12438 & n12461;
  assign n12463 = n3804 & n3861;
  assign n12464 = ~pi067 & n3912;
  assign n12465 = ~n3903 & ~n12464;
  assign n12466 = ~n3785 & n12465;
  assign n12467 = ~pi117 & ~n12466;
  assign n12468 = ~n12463 & ~n12467;
  assign n12469 = ~n12090 & n12468;
  assign n12470 = n3857 & ~n12075;
  assign n12471 = ~n12136 & ~n12470;
  assign n12472 = pi117 & ~n12471;
  assign n12473 = n12469 & ~n12472;
  assign n12474 = ~pi002 & ~n12473;
  assign n12475 = ~n3952 & ~n4011;
  assign n12476 = pi117 & ~n12475;
  assign n12477 = pi067 & n3776;
  assign n12478 = pi067 & n12141;
  assign n12479 = ~n12477 & ~n12478;
  assign n12480 = pi117 & ~n12479;
  assign n12481 = ~n12476 & ~n12480;
  assign n12482 = ~pi117 & n3816;
  assign n12483 = pi032 & n12140;
  assign n12484 = n12130 & n12483;
  assign n12485 = ~n3886 & ~n12484;
  assign n12486 = ~pi117 & n3929;
  assign n12487 = n12485 & ~n12486;
  assign n12488 = ~n12482 & n12487;
  assign n12489 = n12481 & n12488;
  assign n12490 = n3822 & n3857;
  assign n12491 = ~n11584 & ~n12490;
  assign n12492 = ~pi002 & ~n12491;
  assign n12493 = ~n3852 & ~n12077;
  assign n12494 = ~pi067 & n11615;
  assign n12495 = n12493 & ~n12494;
  assign n12496 = ~pi117 & ~n12495;
  assign n12497 = ~n11602 & ~n12477;
  assign n12498 = ~n3854 & ~n11638;
  assign n12499 = pi117 & ~n12498;
  assign n12500 = n12497 & ~n12499;
  assign n12501 = ~n12496 & n12500;
  assign n12502 = ~n3783 & ~n12102;
  assign n12503 = ~n3796 & n12502;
  assign n12504 = n12501 & n12503;
  assign n12505 = pi002 & ~n12504;
  assign n12506 = n3861 & n3927;
  assign n12507 = n3782 & n3897;
  assign n12508 = ~n12506 & ~n12507;
  assign n12509 = ~pi002 & ~n12508;
  assign n12510 = ~n12505 & ~n12509;
  assign n12511 = ~n12492 & n12510;
  assign n12512 = n12489 & n12511;
  assign n12513 = ~pi036 & ~n12512;
  assign n12514 = pi002 & n12486;
  assign n12515 = pi067 & n3886;
  assign n12516 = n3854 & n3897;
  assign n12517 = ~n12515 & ~n12516;
  assign n12518 = pi002 & ~n12517;
  assign n12519 = ~n12514 & ~n12518;
  assign n12520 = ~n12513 & n12519;
  assign n12521 = ~n12474 & n12520;
  assign n12522 = pi064 & pi067;
  assign n12523 = ~pi032 & n12522;
  assign n12524 = ~n12483 & ~n12523;
  assign n12525 = ~n3927 & n12524;
  assign n12526 = n11570 & ~n12525;
  assign n12527 = ~n12110 & ~n12526;
  assign n12528 = ~n3930 & ~n11620;
  assign n12529 = ~n3977 & ~n3983;
  assign n12530 = n12528 & n12529;
  assign n12531 = pi002 & ~n12530;
  assign n12532 = ~pi117 & n4008;
  assign n12533 = ~n3860 & ~n3941;
  assign n12534 = pi117 & ~n12533;
  assign n12535 = ~n3815 & ~n12136;
  assign n12536 = ~n3838 & n12535;
  assign n12537 = ~n12534 & n12536;
  assign n12538 = ~n12532 & n12537;
  assign n12539 = ~pi002 & ~n12538;
  assign n12540 = ~n12531 & ~n12539;
  assign n12541 = ~pi117 & n3785;
  assign n12542 = ~n12061 & ~n12541;
  assign n12543 = ~n3815 & ~n11631;
  assign n12544 = ~n3763 & n12543;
  assign n12545 = ~pi117 & ~n12544;
  assign n12546 = pi117 & n12136;
  assign n12547 = ~n12545 & ~n12546;
  assign n12548 = n12542 & n12547;
  assign n12549 = n12540 & n12548;
  assign n12550 = n12527 & n12549;
  assign n12551 = pi036 & ~n12550;
  assign n12552 = n12521 & ~n12551;
  assign n12553 = ~pi117 & n11602;
  assign n12554 = ~n4028 & ~n12553;
  assign n12555 = ~pi117 & n4010;
  assign n12556 = n12554 & ~n12555;
  assign n12557 = n12552 & n12556;
  assign n12558 = ~n12462 & n12557;
  assign n12559 = n12462 & ~n12557;
  assign n12560 = ~n12558 & ~n12559;
  assign n12561 = n11649 & ~n12560;
  assign n12562 = ~n11649 & n12560;
  assign n12563 = ~n12561 & ~n12562;
  assign n12564 = ~n12369 & n12563;
  assign n12565 = n12369 & ~n12563;
  assign n12566 = ~n12564 & ~n12565;
  assign n12567 = ~pi529 & n12566;
  assign po168 = n12270 | n12567;
  assign n12569 = pi281 & pi426;
  assign n12570 = ~pi281 & ~pi426;
  assign n12571 = ~n12569 & ~n12570;
  assign n12572 = pi529 & n12571;
  assign n12573 = pi067 & n3788;
  assign n12574 = ~n12114 & ~n12573;
  assign n12575 = ~n3888 & n12574;
  assign n12576 = n3865 & ~n12575;
  assign n12577 = pi002 & n3782;
  assign n12578 = n12130 & n12577;
  assign n12579 = ~n12576 & ~n12578;
  assign n12580 = ~pi067 & n3846;
  assign n12581 = ~pi032 & n3794;
  assign n12582 = ~n3886 & ~n12581;
  assign n12583 = ~n11594 & n12582;
  assign n12584 = ~n12580 & n12583;
  assign n12585 = n11570 & ~n12584;
  assign n12586 = ~n3894 & ~n11620;
  assign n12587 = ~n3913 & n12586;
  assign n12588 = n12098 & ~n12587;
  assign n12589 = ~n3977 & ~n12086;
  assign n12590 = ~pi002 & ~n12589;
  assign n12591 = ~pi067 & n3822;
  assign n12592 = ~n12090 & ~n12591;
  assign n12593 = ~n12136 & n12592;
  assign n12594 = n3780 & ~n12593;
  assign n12595 = ~n12590 & ~n12594;
  assign n12596 = ~n12588 & n12595;
  assign n12597 = ~n12585 & n12596;
  assign n12598 = ~n3887 & ~n12113;
  assign n12599 = n12597 & n12598;
  assign n12600 = n12579 & n12599;
  assign n12601 = ~n3771 & ~n3898;
  assign n12602 = ~n3954 & n12601;
  assign n12603 = n3865 & ~n12602;
  assign n12604 = ~n3816 & ~n12152;
  assign n12605 = pi002 & ~n12604;
  assign n12606 = ~n3888 & ~n12605;
  assign n12607 = ~n12603 & n12606;
  assign n12608 = ~pi067 & n3882;
  assign n12609 = ~n3795 & ~n3890;
  assign n12610 = ~n3806 & ~n3882;
  assign n12611 = n12609 & n12610;
  assign n12612 = ~pi117 & ~n12611;
  assign n12613 = ~n12608 & ~n12612;
  assign n12614 = n12607 & n12613;
  assign n12615 = ~pi117 & n12077;
  assign n12616 = n3762 & n3975;
  assign n12617 = ~pi067 & n12102;
  assign n12618 = ~n12616 & ~n12617;
  assign n12619 = ~n12615 & n12618;
  assign n12620 = ~n3806 & ~n12078;
  assign n12621 = n12619 & n12620;
  assign n12622 = ~pi002 & ~n12621;
  assign n12623 = pi117 & n11602;
  assign n12624 = ~n12622 & ~n12623;
  assign n12625 = n12614 & n12624;
  assign n12626 = pi036 & ~n12625;
  assign n12627 = n12600 & ~n12626;
  assign n12628 = ~pi067 & ~n3821;
  assign n12629 = pi067 & ~n3898;
  assign n12630 = ~n12628 & ~n12629;
  assign n12631 = ~n3927 & ~n12630;
  assign n12632 = ~pi117 & ~n12631;
  assign n12633 = n12543 & ~n12632;
  assign n12634 = ~n3783 & n12633;
  assign n12635 = pi002 & ~n12634;
  assign n12636 = ~n3930 & ~n11600;
  assign n12637 = ~pi117 & ~n12636;
  assign n12638 = ~n12090 & ~n12637;
  assign n12639 = ~n3767 & ~n3776;
  assign n12640 = n3865 & ~n12639;
  assign n12641 = n12638 & ~n12640;
  assign n12642 = ~n12635 & n12641;
  assign n12643 = ~pi067 & n3816;
  assign n12644 = ~n3970 & ~n12643;
  assign n12645 = ~pi117 & ~n12644;
  assign n12646 = ~n12117 & ~n12645;
  assign n12647 = ~n11600 & n12646;
  assign n12648 = ~pi002 & ~n12647;
  assign n12649 = n3794 & n3897;
  assign n12650 = pi117 & n11630;
  assign n12651 = ~n12649 & ~n12650;
  assign n12652 = ~pi002 & ~n12651;
  assign n12653 = ~pi067 & n3996;
  assign n12654 = ~n3988 & ~n12653;
  assign n12655 = pi117 & ~n12654;
  assign n12656 = ~n4028 & ~n12655;
  assign n12657 = ~n12652 & n12656;
  assign n12658 = ~n12648 & n12657;
  assign n12659 = n12642 & n12658;
  assign n12660 = ~pi036 & ~n12659;
  assign n12661 = n12627 & ~n12660;
  assign n12662 = ~n4161 & n12661;
  assign n12663 = n4161 & ~n12661;
  assign n12664 = ~n12662 & ~n12663;
  assign n12665 = n4267 & ~n8263;
  assign n12666 = ~n4267 & n8263;
  assign n12667 = ~n12665 & ~n12666;
  assign n12668 = ~n12664 & n12667;
  assign n12669 = n12664 & ~n12667;
  assign n12670 = ~n12668 & ~n12669;
  assign n12671 = ~pi281 & ~n3421;
  assign n12672 = pi281 & n3421;
  assign n12673 = ~n12671 & ~n12672;
  assign n12674 = ~n3591 & n11452;
  assign n12675 = n3591 & ~n11452;
  assign n12676 = ~n12674 & ~n12675;
  assign n12677 = ~n12673 & n12676;
  assign n12678 = n12673 & ~n12676;
  assign n12679 = ~n12677 & ~n12678;
  assign n12680 = n12670 & n12679;
  assign n12681 = ~n12670 & ~n12679;
  assign n12682 = ~n12680 & ~n12681;
  assign n12683 = ~pi529 & n12682;
  assign po169 = n12572 | n12683;
  assign n12685 = ~pi172 & pi484;
  assign n12686 = pi172 & ~pi484;
  assign n12687 = ~n12685 & ~n12686;
  assign n12688 = pi529 & ~n12687;
  assign n12689 = ~n3449 & ~n3575;
  assign n12690 = n3436 & ~n12689;
  assign n12691 = pi092 & n12690;
  assign n12692 = ~n11528 & ~n12691;
  assign n12693 = ~pi092 & n3573;
  assign n12694 = n3425 & n3468;
  assign n12695 = ~n3470 & ~n12694;
  assign n12696 = ~pi092 & ~n12695;
  assign n12697 = ~n12693 & ~n12696;
  assign n12698 = ~n3503 & n12697;
  assign n12699 = pi089 & ~n12698;
  assign n12700 = pi028 & n11384;
  assign n12701 = ~n8232 & ~n11420;
  assign n12702 = ~n3552 & n12701;
  assign n12703 = ~pi092 & ~n12702;
  assign n12704 = pi028 & n3530;
  assign n12705 = ~n3494 & ~n12704;
  assign n12706 = ~n8236 & n12705;
  assign n12707 = pi092 & ~n12706;
  assign n12708 = n3449 & n8174;
  assign n12709 = ~n12707 & ~n12708;
  assign n12710 = ~n12703 & n12709;
  assign n12711 = ~n12700 & n12710;
  assign n12712 = ~n8144 & n12711;
  assign n12713 = ~pi089 & ~n12712;
  assign n12714 = ~pi028 & n11438;
  assign n12715 = ~n8161 & ~n12714;
  assign n12716 = n3476 & ~n12715;
  assign n12717 = n3476 & n12219;
  assign n12718 = ~n12716 & ~n12717;
  assign n12719 = ~n12713 & n12718;
  assign n12720 = ~n12699 & n12719;
  assign n12721 = n12692 & n12720;
  assign n12722 = pi085 & n3433;
  assign n12723 = n3467 & n12722;
  assign n12724 = ~n3578 & ~n11489;
  assign n12725 = ~n8180 & n12724;
  assign n12726 = ~pi092 & ~n12725;
  assign n12727 = ~n3566 & ~n12726;
  assign n12728 = ~n3516 & ~n8213;
  assign n12729 = pi092 & ~n12728;
  assign n12730 = n12727 & ~n12729;
  assign n12731 = pi089 & ~n12730;
  assign n12732 = ~n3496 & ~n12271;
  assign n12733 = n3488 & n3555;
  assign n12734 = ~n8236 & ~n12733;
  assign n12735 = ~pi089 & ~n12734;
  assign n12736 = n12732 & ~n12735;
  assign n12737 = ~n12731 & n12736;
  assign n12738 = ~n12723 & n12737;
  assign n12739 = ~pi053 & ~n12738;
  assign n12740 = pi092 & n8212;
  assign n12741 = ~pi028 & pi046;
  assign n12742 = pi085 & n12741;
  assign n12743 = ~n11384 & ~n12742;
  assign n12744 = ~pi092 & ~n12743;
  assign n12745 = ~n12740 & ~n12744;
  assign n12746 = ~n8246 & n12745;
  assign n12747 = pi089 & ~n12746;
  assign n12748 = ~n3440 & ~n3450;
  assign n12749 = ~n3502 & n12748;
  assign n12750 = n3433 & ~n12749;
  assign n12751 = ~n8247 & ~n8252;
  assign n12752 = ~n3509 & n12751;
  assign n12753 = ~n12750 & n12752;
  assign n12754 = pi092 & n11407;
  assign n12755 = ~pi092 & n3438;
  assign n12756 = ~n12225 & ~n12755;
  assign n12757 = ~n11470 & n12756;
  assign n12758 = ~n12754 & n12757;
  assign n12759 = ~n3481 & ~n8172;
  assign n12760 = ~n11519 & n12759;
  assign n12761 = ~n12296 & n12760;
  assign n12762 = n12758 & n12761;
  assign n12763 = ~pi089 & ~n12762;
  assign n12764 = n12753 & ~n12763;
  assign n12765 = ~n12747 & n12764;
  assign n12766 = pi053 & ~n12765;
  assign n12767 = ~n12739 & ~n12766;
  assign n12768 = n12721 & n12767;
  assign n12769 = ~n11452 & n12768;
  assign n12770 = n11452 & ~n12768;
  assign n12771 = ~n12769 & ~n12770;
  assign n12772 = ~n12057 & n12160;
  assign n12773 = n12057 & ~n12160;
  assign n12774 = ~n12772 & ~n12773;
  assign n12775 = ~n12771 & n12774;
  assign n12776 = n12771 & ~n12774;
  assign n12777 = ~n12775 & ~n12776;
  assign n12778 = ~pi075 & pi080;
  assign n12779 = ~pi079 & n12778;
  assign n12780 = ~n3278 & ~n3352;
  assign n12781 = n12779 & ~n12780;
  assign n12782 = ~n11936 & ~n12781;
  assign n12783 = pi079 & n8025;
  assign n12784 = ~n8082 & ~n8130;
  assign n12785 = ~n3338 & n12784;
  assign n12786 = ~pi080 & ~n12785;
  assign n12787 = pi079 & n3385;
  assign n12788 = ~n8109 & ~n12787;
  assign n12789 = ~n3369 & n12788;
  assign n12790 = pi080 & ~n12789;
  assign n12791 = n3278 & n3366;
  assign n12792 = ~n12790 & ~n12791;
  assign n12793 = ~n12786 & n12792;
  assign n12794 = ~n12783 & n12793;
  assign n12795 = ~n11762 & n12794;
  assign n12796 = ~pi073 & ~n12795;
  assign n12797 = ~pi080 & n3358;
  assign n12798 = n3296 & n8061;
  assign n12799 = ~n3262 & ~n12798;
  assign n12800 = ~pi080 & ~n12799;
  assign n12801 = pi080 & n11781;
  assign n12802 = ~n3348 & ~n12801;
  assign n12803 = ~n12800 & n12802;
  assign n12804 = ~n12797 & n12803;
  assign n12805 = pi110 & n3395;
  assign n12806 = ~n3260 & ~n12805;
  assign n12807 = pi080 & ~n12806;
  assign n12808 = n12804 & ~n12807;
  assign n12809 = pi073 & ~n12808;
  assign n12810 = ~n12796 & ~n12809;
  assign n12811 = n12782 & n12810;
  assign n12812 = pi079 & n3350;
  assign n12813 = ~n3355 & ~n12812;
  assign n12814 = ~n11900 & n12813;
  assign n12815 = ~pi080 & ~n12814;
  assign n12816 = ~n3327 & ~n12815;
  assign n12817 = ~n3375 & ~n8026;
  assign n12818 = pi080 & ~n12817;
  assign n12819 = n12816 & ~n12818;
  assign n12820 = pi073 & ~n12819;
  assign n12821 = n3283 & n3339;
  assign n12822 = ~n8109 & ~n12821;
  assign n12823 = ~pi073 & ~n12822;
  assign n12824 = pi075 & n3288;
  assign n12825 = n3259 & n12824;
  assign n12826 = ~n12823 & ~n12825;
  assign n12827 = ~n12820 & n12826;
  assign n12828 = ~pi080 & n11801;
  assign n12829 = ~n3365 & ~n12828;
  assign n12830 = ~pi015 & n12829;
  assign n12831 = n12827 & n12830;
  assign n12832 = n3297 & n3395;
  assign n12833 = ~n3402 & ~n12832;
  assign n12834 = pi015 & n12833;
  assign n12835 = pi080 & n3291;
  assign n12836 = pi042 & n8061;
  assign n12837 = ~n8025 & ~n12836;
  assign n12838 = ~pi080 & ~n12837;
  assign n12839 = ~n12835 & ~n12838;
  assign n12840 = ~pi080 & n11863;
  assign n12841 = n12839 & ~n12840;
  assign n12842 = pi073 & ~n12841;
  assign n12843 = ~n3307 & ~n3394;
  assign n12844 = ~n3293 & n12843;
  assign n12845 = n3288 & ~n12844;
  assign n12846 = ~n11752 & ~n12845;
  assign n12847 = ~pi080 & n3292;
  assign n12848 = pi080 & n8038;
  assign n12849 = ~n11767 & ~n12848;
  assign n12850 = ~n11804 & n12849;
  assign n12851 = ~pi080 & n3260;
  assign n12852 = ~n11818 & ~n12851;
  assign n12853 = n12850 & n12852;
  assign n12854 = ~n12847 & n12853;
  assign n12855 = ~n3279 & ~n8079;
  assign n12856 = n12854 & n12855;
  assign n12857 = ~pi073 & ~n12856;
  assign n12858 = n12846 & ~n12857;
  assign n12859 = ~n12842 & n12858;
  assign n12860 = n12834 & n12859;
  assign n12861 = ~n12831 & ~n12860;
  assign n12862 = n12811 & ~n12861;
  assign n12863 = ~n8140 & n12862;
  assign n12864 = n8140 & ~n12862;
  assign n12865 = ~n12863 & ~n12864;
  assign n12866 = ~pi172 & n11953;
  assign n12867 = pi172 & ~n11953;
  assign n12868 = ~n12866 & ~n12867;
  assign n12869 = ~n12865 & n12868;
  assign n12870 = n12865 & ~n12868;
  assign n12871 = ~n12869 & ~n12870;
  assign n12872 = ~n12777 & n12871;
  assign n12873 = n12777 & ~n12871;
  assign n12874 = ~n12872 & ~n12873;
  assign n12875 = ~pi529 & n12874;
  assign po170 = n12688 | n12875;
  assign n12877 = pi162 & pi485;
  assign n12878 = ~pi162 & ~pi485;
  assign n12879 = ~n12877 & ~n12878;
  assign n12880 = pi529 & n12879;
  assign n12881 = ~n8034 & ~n11752;
  assign n12882 = ~pi079 & n3310;
  assign n12883 = n12881 & ~n12882;
  assign n12884 = ~pi080 & ~n12883;
  assign n12885 = ~n3415 & ~n12840;
  assign n12886 = ~n11884 & ~n12832;
  assign n12887 = pi080 & ~n12886;
  assign n12888 = n12885 & ~n12887;
  assign n12889 = ~n12884 & n12888;
  assign n12890 = ~pi073 & ~n12889;
  assign n12891 = ~pi079 & n3312;
  assign n12892 = ~n3326 & ~n12891;
  assign n12893 = n3290 & ~n12892;
  assign n12894 = ~pi079 & ~n8113;
  assign n12895 = ~n11814 & ~n12894;
  assign n12896 = ~pi073 & ~n12895;
  assign n12897 = ~n3278 & ~n3350;
  assign n12898 = n12778 & ~n12897;
  assign n12899 = pi079 & n12898;
  assign n12900 = n3385 & n3395;
  assign n12901 = ~n11858 & ~n12900;
  assign n12902 = ~pi080 & ~n12901;
  assign n12903 = ~n12899 & ~n12902;
  assign n12904 = ~n3367 & n12903;
  assign n12905 = n3352 & n3366;
  assign n12906 = n3258 & n3302;
  assign n12907 = pi080 & n3372;
  assign n12908 = ~n12906 & ~n12907;
  assign n12909 = ~n12905 & n12908;
  assign n12910 = ~n3291 & ~n8026;
  assign n12911 = n12909 & n12910;
  assign n12912 = pi073 & ~n12911;
  assign n12913 = n12904 & ~n12912;
  assign n12914 = ~n12896 & n12913;
  assign n12915 = ~n12893 & n12914;
  assign n12916 = ~pi015 & ~n12915;
  assign n12917 = ~pi110 & n11826;
  assign n12918 = ~n12812 & ~n12917;
  assign n12919 = ~pi080 & ~n12918;
  assign n12920 = ~n3325 & ~n12919;
  assign n12921 = ~pi080 & n3263;
  assign n12922 = ~n11868 & ~n12921;
  assign n12923 = ~n3394 & n12922;
  assign n12924 = pi073 & ~n12923;
  assign n12925 = n3366 & n8132;
  assign n12926 = ~n3260 & ~n8051;
  assign n12927 = ~n3411 & n12926;
  assign n12928 = pi080 & ~n12927;
  assign n12929 = ~n12925 & ~n12928;
  assign n12930 = pi079 & n11803;
  assign n12931 = ~pi071 & n11826;
  assign n12932 = ~n8079 & ~n12931;
  assign n12933 = ~n12930 & n12932;
  assign n12934 = n12929 & n12933;
  assign n12935 = ~pi073 & ~n12934;
  assign n12936 = ~n3308 & ~n3314;
  assign n12937 = ~n11859 & n12936;
  assign n12938 = pi080 & ~n11762;
  assign n12939 = n12937 & n12938;
  assign n12940 = ~n3294 & ~n8062;
  assign n12941 = ~pi080 & n12940;
  assign n12942 = ~n12939 & ~n12941;
  assign n12943 = ~n12935 & ~n12942;
  assign n12944 = ~n12924 & n12943;
  assign n12945 = n12920 & n12944;
  assign n12946 = ~n11792 & n12945;
  assign n12947 = pi015 & ~n12946;
  assign n12948 = pi080 & n3263;
  assign n12949 = ~pi110 & n12948;
  assign n12950 = n3395 & n12949;
  assign n12951 = ~pi080 & n8109;
  assign n12952 = ~pi079 & n3394;
  assign n12953 = pi080 & n12952;
  assign n12954 = ~n11801 & ~n11879;
  assign n12955 = ~n12953 & n12954;
  assign n12956 = ~n12951 & n12955;
  assign n12957 = ~n11785 & n12956;
  assign n12958 = pi073 & ~n12957;
  assign n12959 = ~pi080 & n12906;
  assign n12960 = ~n12958 & ~n12959;
  assign n12961 = ~n12950 & n12960;
  assign n12962 = ~n12947 & n12961;
  assign n12963 = ~n12916 & n12962;
  assign n12964 = ~n12890 & n12963;
  assign n12965 = ~pi162 & ~n12964;
  assign n12966 = pi162 & n12964;
  assign n12967 = ~n12965 & ~n12966;
  assign n12968 = n3926 & n4267;
  assign n12969 = ~n3926 & ~n4267;
  assign n12970 = ~n12968 & ~n12969;
  assign n12971 = ~n8266 & ~n12970;
  assign n12972 = ~n8264 & n12970;
  assign n12973 = ~n8265 & n12972;
  assign n12974 = ~n12971 & ~n12973;
  assign n12975 = n12967 & n12974;
  assign n12976 = ~n12967 & ~n12974;
  assign n12977 = ~n12975 & ~n12976;
  assign n12978 = ~pi529 & n12977;
  assign po171 = n12880 | n12978;
  assign n12980 = ~pi226 & pi445;
  assign n12981 = pi226 & ~pi445;
  assign n12982 = ~n12980 & ~n12981;
  assign n12983 = pi529 & n12982;
  assign n12984 = n3257 & n11901;
  assign n12985 = ~n3415 & ~n12984;
  assign n12986 = ~pi080 & n3365;
  assign n12987 = pi079 & n3271;
  assign n12988 = ~n12986 & ~n12987;
  assign n12989 = pi073 & ~n12988;
  assign n12990 = ~n12828 & ~n12989;
  assign n12991 = n12985 & n12990;
  assign n12992 = ~n11883 & n12991;
  assign n12993 = ~pi079 & n3313;
  assign n12994 = ~n8082 & ~n12993;
  assign n12995 = ~n3260 & n12994;
  assign n12996 = ~pi080 & ~n12995;
  assign n12997 = n8061 & ~n11891;
  assign n12998 = ~n3295 & ~n12997;
  assign n12999 = pi080 & ~n12998;
  assign n13000 = n3288 & n8054;
  assign n13001 = ~n12999 & ~n13000;
  assign n13002 = ~n3292 & n13001;
  assign n13003 = ~n12996 & n13002;
  assign n13004 = ~pi073 & ~n13003;
  assign n13005 = n12992 & ~n13004;
  assign n13006 = pi075 & n11899;
  assign n13007 = pi071 & n11826;
  assign n13008 = ~n13006 & ~n13007;
  assign n13009 = ~n3386 & n13008;
  assign n13010 = n8117 & ~n13009;
  assign n13011 = ~n3317 & ~n11859;
  assign n13012 = ~n3308 & ~n12930;
  assign n13013 = n13011 & n13012;
  assign n13014 = pi073 & ~n13013;
  assign n13015 = pi080 & n3295;
  assign n13016 = ~n3372 & ~n3375;
  assign n13017 = ~n8078 & n13016;
  assign n13018 = ~pi080 & ~n13017;
  assign n13019 = ~n13015 & ~n13018;
  assign n13020 = ~n11863 & n13019;
  assign n13021 = ~n12851 & n13020;
  assign n13022 = ~n13014 & n13021;
  assign n13023 = ~n13010 & n13022;
  assign n13024 = ~n3295 & ~n3372;
  assign n13025 = ~n8059 & ~n11813;
  assign n13026 = pi080 & ~n13025;
  assign n13027 = ~pi080 & n11828;
  assign n13028 = ~n8037 & ~n13027;
  assign n13029 = ~n13026 & n13028;
  assign n13030 = n13024 & n13029;
  assign n13031 = ~pi073 & ~n13030;
  assign n13032 = ~n11948 & ~n13031;
  assign n13033 = n13023 & n13032;
  assign n13034 = pi015 & ~n13033;
  assign n13035 = pi079 & n3378;
  assign n13036 = ~n3291 & ~n13035;
  assign n13037 = pi079 & n11900;
  assign n13038 = n13036 & ~n13037;
  assign n13039 = ~n12952 & n13038;
  assign n13040 = pi080 & ~n13039;
  assign n13041 = n3270 & n3401;
  assign n13042 = ~n11788 & ~n13041;
  assign n13043 = ~pi079 & n8132;
  assign n13044 = n3288 & n3386;
  assign n13045 = ~n13043 & ~n13044;
  assign n13046 = n13042 & n13045;
  assign n13047 = ~pi073 & ~n13046;
  assign n13048 = ~n8051 & ~n11815;
  assign n13049 = pi080 & ~n13048;
  assign n13050 = ~n3335 & ~n8055;
  assign n13051 = ~pi079 & n3374;
  assign n13052 = n13050 & ~n13051;
  assign n13053 = ~pi080 & ~n13052;
  assign n13054 = ~n3373 & ~n8121;
  assign n13055 = ~n3333 & n13054;
  assign n13056 = ~n3348 & ~n13035;
  assign n13057 = n13055 & n13056;
  assign n13058 = ~n13053 & n13057;
  assign n13059 = ~n13049 & n13058;
  assign n13060 = pi073 & ~n13059;
  assign n13061 = ~n13047 & ~n13060;
  assign n13062 = ~n13040 & n13061;
  assign n13063 = ~pi071 & n8086;
  assign n13064 = n3258 & n13063;
  assign n13065 = n3283 & n13006;
  assign n13066 = ~n12986 & ~n13065;
  assign n13067 = ~n3271 & n13066;
  assign n13068 = ~n13064 & n13067;
  assign n13069 = n13062 & n13068;
  assign n13070 = ~pi015 & ~n13069;
  assign n13071 = ~n13034 & ~n13070;
  assign n13072 = n13005 & n13071;
  assign n13073 = pi226 & ~n13072;
  assign n13074 = ~pi226 & n13072;
  assign n13075 = ~n13073 & ~n13074;
  assign n13076 = ~n11853 & n13075;
  assign n13077 = n11853 & ~n13075;
  assign n13078 = ~n13076 & ~n13077;
  assign n13079 = ~n12252 & n12560;
  assign n13080 = n12252 & ~n12560;
  assign n13081 = ~n13079 & ~n13080;
  assign n13082 = n13078 & n13081;
  assign n13083 = ~n13078 & ~n13081;
  assign n13084 = ~n13082 & ~n13083;
  assign n13085 = ~pi529 & n13084;
  assign po172 = n12983 | n13085;
  assign n13087 = ~pi192 & pi453;
  assign n13088 = pi192 & ~pi453;
  assign n13089 = ~n13087 & ~n13088;
  assign n13090 = pi529 & n13089;
  assign n13091 = pi192 & ~n12964;
  assign n13092 = ~pi192 & n12964;
  assign n13093 = ~n13091 & ~n13092;
  assign n13094 = ~n4042 & n4267;
  assign n13095 = n4042 & ~n4267;
  assign n13096 = ~n13094 & ~n13095;
  assign n13097 = n8263 & ~n11452;
  assign n13098 = ~n8263 & n11452;
  assign n13099 = ~n13097 & ~n13098;
  assign n13100 = n13096 & ~n13099;
  assign n13101 = ~n13096 & n13099;
  assign n13102 = ~n13100 & ~n13101;
  assign n13103 = n13093 & n13102;
  assign n13104 = ~n13093 & ~n13102;
  assign n13105 = ~n13103 & ~n13104;
  assign n13106 = ~pi529 & n13105;
  assign po173 = n13090 | n13106;
  assign n13108 = pi278 & pi513;
  assign n13109 = ~pi278 & ~pi513;
  assign n13110 = ~n13108 & ~n13109;
  assign n13111 = pi529 & n13110;
  assign n13112 = pi074 & n4831;
  assign n13113 = ~n8952 & ~n13112;
  assign n13114 = ~n4919 & n13113;
  assign n13115 = n4882 & ~n13114;
  assign n13116 = ~n5009 & ~n9012;
  assign n13117 = ~pi003 & ~n13116;
  assign n13118 = ~n4925 & ~n8946;
  assign n13119 = ~n4944 & n13118;
  assign n13120 = n9035 & ~n13119;
  assign n13121 = ~n4918 & ~n8951;
  assign n13122 = ~pi074 & n4877;
  assign n13123 = ~pi074 & n4802;
  assign n13124 = ~n4854 & ~n4917;
  assign n13125 = ~n13123 & n13124;
  assign n13126 = ~n13122 & n13125;
  assign n13127 = pi003 & ~pi120;
  assign n13128 = ~n13126 & n13127;
  assign n13129 = n13121 & ~n13128;
  assign n13130 = ~n13120 & n13129;
  assign n13131 = ~pi074 & n4806;
  assign n13132 = ~n9019 & ~n13131;
  assign n13133 = ~n8961 & n13132;
  assign n13134 = n4835 & ~n13133;
  assign n13135 = pi003 & n4828;
  assign n13136 = n8967 & n13135;
  assign n13137 = ~n13134 & ~n13136;
  assign n13138 = n13130 & n13137;
  assign n13139 = ~n13117 & n13138;
  assign n13140 = ~n13115 & n13139;
  assign n13141 = ~n4847 & ~n4929;
  assign n13142 = ~n4985 & n13141;
  assign n13143 = n4882 & ~n13142;
  assign n13144 = ~n4798 & ~n8989;
  assign n13145 = pi003 & ~n13144;
  assign n13146 = ~n4919 & ~n13145;
  assign n13147 = ~n13143 & n13146;
  assign n13148 = ~pi074 & n4913;
  assign n13149 = ~n4921 & ~n4997;
  assign n13150 = ~n4815 & ~n4913;
  assign n13151 = n13149 & n13150;
  assign n13152 = ~pi120 & ~n13151;
  assign n13153 = ~n13148 & ~n13152;
  assign n13154 = n13147 & n13153;
  assign n13155 = ~pi120 & n9029;
  assign n13156 = ~pi074 & n8983;
  assign n13157 = ~n13155 & ~n13156;
  assign n13158 = n4837 & n5007;
  assign n13159 = n13157 & ~n13158;
  assign n13160 = ~n4815 & ~n9030;
  assign n13161 = n13159 & n13160;
  assign n13162 = ~pi003 & ~n13161;
  assign n13163 = pi120 & n9013;
  assign n13164 = ~n13162 & ~n13163;
  assign n13165 = n13154 & n13164;
  assign n13166 = pi044 & ~n13165;
  assign n13167 = n13140 & ~n13166;
  assign n13168 = pi074 & n4817;
  assign n13169 = ~n4976 & ~n13168;
  assign n13170 = ~pi120 & ~n13169;
  assign n13171 = ~n9019 & ~n13170;
  assign n13172 = ~pi074 & ~n4805;
  assign n13173 = pi074 & ~n4929;
  assign n13174 = ~n13172 & ~n13173;
  assign n13175 = ~n4972 & ~n13174;
  assign n13176 = ~pi120 & ~n13175;
  assign n13177 = pi074 & n9042;
  assign n13178 = ~n4795 & ~n13177;
  assign n13179 = ~n13176 & n13178;
  assign n13180 = ~n4829 & n13179;
  assign n13181 = pi003 & ~n13180;
  assign n13182 = ~n4840 & ~n4844;
  assign n13183 = n4882 & ~n13182;
  assign n13184 = ~n13181 & ~n13183;
  assign n13185 = n13171 & n13184;
  assign n13186 = ~pi016 & n9013;
  assign n13187 = ~n5002 & ~n13186;
  assign n13188 = ~pi120 & ~n13187;
  assign n13189 = ~n8955 & ~n13188;
  assign n13190 = ~n13168 & n13189;
  assign n13191 = ~pi003 & ~n13190;
  assign n13192 = n4794 & n4928;
  assign n13193 = pi120 & n8999;
  assign n13194 = ~n13192 & ~n13193;
  assign n13195 = ~pi003 & ~n13194;
  assign n13196 = ~pi074 & n5028;
  assign n13197 = ~n5014 & ~n13196;
  assign n13198 = pi120 & ~n13197;
  assign n13199 = ~n5064 & ~n13198;
  assign n13200 = ~n13195 & n13199;
  assign n13201 = ~n13191 & n13200;
  assign n13202 = n13185 & n13201;
  assign n13203 = ~pi044 & ~n13202;
  assign n13204 = n13167 & ~n13203;
  assign n13205 = ~n5192 & n13204;
  assign n13206 = n5192 & ~n13204;
  assign n13207 = ~n13205 & ~n13206;
  assign n13208 = ~n5298 & n9162;
  assign n13209 = n5298 & ~n9162;
  assign n13210 = ~n13208 & ~n13209;
  assign n13211 = ~n13207 & n13210;
  assign n13212 = n13207 & ~n13210;
  assign n13213 = ~n13211 & ~n13212;
  assign n13214 = ~pi278 & ~n4451;
  assign n13215 = pi278 & n4451;
  assign n13216 = ~n13214 & ~n13215;
  assign n13217 = ~n4620 & n8748;
  assign n13218 = n4620 & ~n8748;
  assign n13219 = ~n13217 & ~n13218;
  assign n13220 = n13216 & n13219;
  assign n13221 = ~n13216 & ~n13219;
  assign n13222 = ~n13220 & ~n13221;
  assign n13223 = ~n13213 & n13222;
  assign n13224 = n13213 & ~n13222;
  assign n13225 = ~n13223 & ~n13224;
  assign n13226 = ~pi529 & n13225;
  assign po174 = n13111 | n13226;
  assign n13228 = pi280 & pi470;
  assign n13229 = ~pi280 & ~pi470;
  assign n13230 = ~n13228 & ~n13229;
  assign n13231 = pi529 & n13230;
  assign n13232 = ~n8423 & n9554;
  assign n13233 = n8423 & ~n9554;
  assign n13234 = ~n13232 & ~n13233;
  assign n13235 = ~pi280 & ~n4451;
  assign n13236 = pi280 & n4451;
  assign n13237 = ~n13235 & ~n13236;
  assign n13238 = n13234 & ~n13237;
  assign n13239 = ~n13234 & n13237;
  assign n13240 = ~n13238 & ~n13239;
  assign n13241 = n4786 & n13204;
  assign n13242 = ~n4786 & ~n13204;
  assign n13243 = ~n13241 & ~n13242;
  assign n13244 = ~n9560 & ~n13243;
  assign n13245 = n4786 & ~n13204;
  assign n13246 = ~n4786 & n13204;
  assign n13247 = ~n13245 & ~n13246;
  assign n13248 = n9560 & ~n13247;
  assign n13249 = ~n13244 & ~n13248;
  assign n13250 = n13240 & n13249;
  assign n13251 = ~n13240 & ~n13249;
  assign n13252 = ~n13250 & ~n13251;
  assign n13253 = ~pi529 & n13252;
  assign po175 = n13231 | n13253;
  assign n13255 = ~pi141 & pi488;
  assign n13256 = pi141 & ~pi488;
  assign n13257 = ~n13255 & ~n13256;
  assign n13258 = pi529 & ~n13257;
  assign n13259 = ~pi120 & n4815;
  assign n13260 = pi120 & n4831;
  assign n13261 = ~n13259 & ~n13260;
  assign n13262 = pi074 & ~n13261;
  assign n13263 = pi120 & n5018;
  assign n13264 = ~n4807 & ~n9042;
  assign n13265 = ~pi120 & ~n13264;
  assign n13266 = ~n5045 & ~n13265;
  assign n13267 = ~n13263 & n13266;
  assign n13268 = ~n8946 & n13267;
  assign n13269 = pi003 & ~n13268;
  assign n13270 = ~n5053 & ~n13177;
  assign n13271 = ~n8999 & n13270;
  assign n13272 = ~pi120 & ~n13271;
  assign n13273 = ~pi045 & ~pi074;
  assign n13274 = pi016 & n13273;
  assign n13275 = ~n4817 & ~n13274;
  assign n13276 = ~pi016 & n4923;
  assign n13277 = ~n5043 & ~n13276;
  assign n13278 = n13275 & n13277;
  assign n13279 = pi120 & ~n13278;
  assign n13280 = ~n13272 & ~n13279;
  assign n13281 = ~pi120 & n4943;
  assign n13282 = pi074 & n4843;
  assign n13283 = ~n4961 & ~n13282;
  assign n13284 = ~n9036 & n13283;
  assign n13285 = ~n13281 & n13284;
  assign n13286 = ~n9039 & n13285;
  assign n13287 = ~pi003 & ~n13286;
  assign n13288 = n13280 & ~n13287;
  assign n13289 = ~n13269 & n13288;
  assign n13290 = pi044 & ~n13289;
  assign n13291 = ~n13262 & ~n13290;
  assign n13292 = n4801 & n4980;
  assign n13293 = ~n4996 & ~n13292;
  assign n13294 = ~n4827 & n13293;
  assign n13295 = pi120 & n4862;
  assign n13296 = n13294 & ~n13295;
  assign n13297 = ~n4846 & ~n4903;
  assign n13298 = pi074 & ~n13297;
  assign n13299 = ~n8981 & ~n13298;
  assign n13300 = ~n5053 & n13299;
  assign n13301 = ~pi120 & ~n13300;
  assign n13302 = n13296 & ~n13301;
  assign n13303 = pi003 & ~n13302;
  assign n13304 = ~n5065 & ~n9012;
  assign n13305 = ~n4878 & ~n13123;
  assign n13306 = ~n4795 & n13305;
  assign n13307 = n13304 & n13306;
  assign n13308 = pi120 & ~n13307;
  assign n13309 = ~pi074 & n4929;
  assign n13310 = ~n13168 & ~n13309;
  assign n13311 = ~n9013 & n13310;
  assign n13312 = ~pi120 & ~n13311;
  assign n13313 = ~n4934 & ~n13312;
  assign n13314 = ~n13308 & n13313;
  assign n13315 = ~n5058 & n13314;
  assign n13316 = ~pi003 & ~n13315;
  assign n13317 = ~n13303 & ~n13316;
  assign n13318 = n4928 & n4947;
  assign n13319 = ~n9010 & ~n13318;
  assign n13320 = pi003 & ~n13319;
  assign n13321 = pi074 & n4983;
  assign n13322 = n4794 & n4890;
  assign n13323 = ~n13321 & ~n13322;
  assign n13324 = ~pi003 & ~n13323;
  assign n13325 = ~n13320 & ~n13324;
  assign n13326 = ~pi074 & n4904;
  assign n13327 = ~n4857 & ~n13326;
  assign n13328 = pi120 & ~n13327;
  assign n13329 = pi003 & n8962;
  assign n13330 = ~n5058 & ~n13329;
  assign n13331 = ~n4949 & ~n13260;
  assign n13332 = ~pi003 & ~n13331;
  assign n13333 = ~pi120 & n4919;
  assign n13334 = ~n13332 & ~n13333;
  assign n13335 = n13330 & n13334;
  assign n13336 = ~pi074 & n4920;
  assign n13337 = ~n4995 & ~n13336;
  assign n13338 = ~n4975 & n13337;
  assign n13339 = n13127 & ~n13338;
  assign n13340 = n13335 & ~n13339;
  assign n13341 = ~n13328 & n13340;
  assign n13342 = n13325 & n13341;
  assign n13343 = ~pi044 & ~n13342;
  assign n13344 = n13317 & ~n13343;
  assign n13345 = n13291 & n13344;
  assign n13346 = n9366 & n13345;
  assign n13347 = ~n9366 & ~n13345;
  assign n13348 = ~n13346 & ~n13347;
  assign n13349 = ~pi118 & n5164;
  assign n13350 = ~pi118 & n4657;
  assign n13351 = ~n13349 & ~n13350;
  assign n13352 = n4642 & n5249;
  assign n13353 = ~n8885 & ~n13352;
  assign n13354 = ~pi066 & n4647;
  assign n13355 = n4733 & n4753;
  assign n13356 = ~n13354 & ~n13355;
  assign n13357 = n13353 & n13356;
  assign n13358 = ~pi034 & ~n13357;
  assign n13359 = ~pi118 & n4706;
  assign n13360 = ~pi118 & n4686;
  assign n13361 = ~n13359 & ~n13360;
  assign n13362 = pi103 & n4748;
  assign n13363 = n8896 & n13362;
  assign n13364 = ~n4759 & ~n13363;
  assign n13365 = n13361 & n13364;
  assign n13366 = pi066 & n4736;
  assign n13367 = ~n4623 & ~n13366;
  assign n13368 = pi066 & n8888;
  assign n13369 = n4636 & n5129;
  assign n13370 = ~n13368 & ~n13369;
  assign n13371 = n13367 & n13370;
  assign n13372 = pi118 & ~n13371;
  assign n13373 = ~n4657 & ~n13366;
  assign n13374 = ~n4663 & ~n5262;
  assign n13375 = ~pi066 & n4723;
  assign n13376 = n13374 & ~n13375;
  assign n13377 = ~pi118 & ~n13376;
  assign n13378 = ~n5147 & ~n9340;
  assign n13379 = pi118 & ~n13378;
  assign n13380 = ~n13377 & ~n13379;
  assign n13381 = n13373 & n13380;
  assign n13382 = ~n4661 & ~n4727;
  assign n13383 = ~n5086 & n13382;
  assign n13384 = n13381 & n13383;
  assign n13385 = pi034 & ~n13384;
  assign n13386 = ~n13372 & ~n13385;
  assign n13387 = n13365 & n13386;
  assign n13388 = ~n13358 & n13387;
  assign n13389 = ~pi038 & ~n13388;
  assign n13390 = ~n4644 & ~n4707;
  assign n13391 = ~n4651 & ~n5141;
  assign n13392 = n13390 & n13391;
  assign n13393 = pi034 & ~n13392;
  assign n13394 = n4726 & ~n5143;
  assign n13395 = ~pi118 & ~n13394;
  assign n13396 = ~n5184 & ~n13395;
  assign n13397 = ~pi118 & n4684;
  assign n13398 = pi118 & n4628;
  assign n13399 = ~n13397 & ~n13398;
  assign n13400 = n13396 & n13399;
  assign n13401 = ~n4628 & ~n4725;
  assign n13402 = ~n5110 & ~n5256;
  assign n13403 = pi118 & ~n13402;
  assign n13404 = ~pi118 & n5169;
  assign n13405 = ~n5271 & ~n13404;
  assign n13406 = ~n13403 & n13405;
  assign n13407 = n13401 & n13406;
  assign n13408 = ~pi034 & ~n13407;
  assign n13409 = ~n8919 & ~n13408;
  assign n13410 = pi066 & pi101;
  assign n13411 = ~pi103 & n13410;
  assign n13412 = ~n13362 & ~n13411;
  assign n13413 = ~n4733 & n13412;
  assign n13414 = ~pi118 & ~n13413;
  assign n13415 = pi034 & n13414;
  assign n13416 = n13409 & ~n13415;
  assign n13417 = n13400 & n13416;
  assign n13418 = ~n13393 & n13417;
  assign n13419 = pi038 & ~n13418;
  assign n13420 = ~pi066 & n4639;
  assign n13421 = ~n4684 & ~n13420;
  assign n13422 = ~n5240 & n13421;
  assign n13423 = n8936 & ~n13422;
  assign n13424 = n5129 & ~n8863;
  assign n13425 = ~n4628 & ~n13424;
  assign n13426 = pi118 & ~n13425;
  assign n13427 = n4753 & n5193;
  assign n13428 = ~n4624 & ~n13427;
  assign n13429 = ~n13426 & n13428;
  assign n13430 = ~pi034 & ~n13429;
  assign n13431 = ~n13423 & ~n13430;
  assign n13432 = pi066 & n4759;
  assign n13433 = ~n13359 & ~n13432;
  assign n13434 = pi034 & ~n13433;
  assign n13435 = n4762 & n8887;
  assign n13436 = ~n4754 & ~n13435;
  assign n13437 = ~n13434 & n13436;
  assign n13438 = n13431 & n13437;
  assign n13439 = ~n13419 & n13438;
  assign n13440 = ~n13389 & n13439;
  assign n13441 = n13351 & n13440;
  assign n13442 = n4490 & n8749;
  assign n13443 = n4550 & ~n8658;
  assign n13444 = ~pi116 & ~n13443;
  assign n13445 = pi116 & n4519;
  assign n13446 = ~n13444 & ~n13445;
  assign n13447 = ~n13442 & n13446;
  assign n13448 = ~n8778 & n13447;
  assign n13449 = pi000 & n8790;
  assign n13450 = pi011 & pi022;
  assign n13451 = ~pi000 & n13450;
  assign n13452 = ~n4562 & ~n13451;
  assign n13453 = ~n13449 & n13452;
  assign n13454 = pi058 & ~n13453;
  assign n13455 = ~pi116 & n13454;
  assign n13456 = ~n4473 & ~n4529;
  assign n13457 = ~n4458 & ~n9113;
  assign n13458 = n13456 & n13457;
  assign n13459 = pi058 & ~n13458;
  assign n13460 = ~n13455 & ~n13459;
  assign n13461 = n13448 & n13460;
  assign n13462 = n4540 & n4582;
  assign n13463 = ~n4519 & ~n4549;
  assign n13464 = ~pi116 & n9149;
  assign n13465 = pi011 & n9069;
  assign n13466 = ~n8670 & ~n13465;
  assign n13467 = pi116 & ~n13466;
  assign n13468 = ~n13464 & ~n13467;
  assign n13469 = n13463 & n13468;
  assign n13470 = ~n8688 & n13469;
  assign n13471 = ~pi058 & ~n13470;
  assign n13472 = ~n13462 & ~n13471;
  assign n13473 = n13461 & n13472;
  assign n13474 = pi060 & ~n13473;
  assign n13475 = pi011 & n8791;
  assign n13476 = pi011 & n4553;
  assign n13477 = ~n8753 & ~n13476;
  assign n13478 = ~n9147 & n13477;
  assign n13479 = ~n13475 & n13478;
  assign n13480 = pi116 & ~n13479;
  assign n13481 = n4471 & n4540;
  assign n13482 = ~n9370 & ~n13481;
  assign n13483 = ~pi011 & n4461;
  assign n13484 = n4481 & n4562;
  assign n13485 = ~n13483 & ~n13484;
  assign n13486 = n13482 & n13485;
  assign n13487 = ~pi058 & ~n13486;
  assign n13488 = ~n4580 & ~n8673;
  assign n13489 = ~pi011 & n4547;
  assign n13490 = n13488 & ~n13489;
  assign n13491 = ~pi116 & ~n13490;
  assign n13492 = ~n4535 & ~n13476;
  assign n13493 = ~n8675 & ~n9388;
  assign n13494 = pi116 & ~n13493;
  assign n13495 = n13492 & ~n13494;
  assign n13496 = ~n13491 & n13495;
  assign n13497 = ~n4551 & ~n4588;
  assign n13498 = ~n8648 & n13497;
  assign n13499 = n13496 & n13498;
  assign n13500 = pi058 & ~n13499;
  assign n13501 = n4484 & n13449;
  assign n13502 = ~pi116 & n4528;
  assign n13503 = ~pi116 & n4502;
  assign n13504 = ~n13502 & ~n13503;
  assign n13505 = ~n4480 & n13504;
  assign n13506 = ~n13501 & n13505;
  assign n13507 = ~n13500 & n13506;
  assign n13508 = ~n13487 & n13507;
  assign n13509 = ~n13480 & n13508;
  assign n13510 = ~pi060 & ~n13509;
  assign n13511 = ~n13474 & ~n13510;
  assign n13512 = pi011 & n4480;
  assign n13513 = ~n13502 & ~n13512;
  assign n13514 = pi058 & ~n13513;
  assign n13515 = ~pi011 & n8675;
  assign n13516 = n4508 & n13515;
  assign n13517 = ~n13514 & ~n13516;
  assign n13518 = ~pi058 & ~pi116;
  assign n13519 = ~pi011 & n4468;
  assign n13520 = ~n8716 & ~n13519;
  assign n13521 = ~n8652 & n13520;
  assign n13522 = n13518 & ~n13521;
  assign n13523 = ~pi116 & n4535;
  assign n13524 = ~n8802 & ~n13523;
  assign n13525 = n4481 & n8638;
  assign n13526 = ~n4460 & ~n4465;
  assign n13527 = n4500 & ~n13526;
  assign n13528 = ~n4519 & ~n13527;
  assign n13529 = pi116 & ~n13528;
  assign n13530 = ~n13525 & ~n13529;
  assign n13531 = ~n4514 & n13530;
  assign n13532 = ~pi058 & ~n13531;
  assign n13533 = ~n4576 & ~n13532;
  assign n13534 = n13524 & n13533;
  assign n13535 = ~n13522 & n13534;
  assign n13536 = n13517 & n13535;
  assign n13537 = n13511 & n13536;
  assign n13538 = ~n13441 & n13537;
  assign n13539 = n13441 & ~n13537;
  assign n13540 = ~n13538 & ~n13539;
  assign n13541 = n4319 & n8598;
  assign n13542 = ~n4381 & ~n8487;
  assign n13543 = ~n13541 & n13542;
  assign n13544 = ~n8565 & n13543;
  assign n13545 = pi019 & n4337;
  assign n13546 = ~n4361 & ~n13545;
  assign n13547 = pi088 & ~n13546;
  assign n13548 = n13544 & ~n13547;
  assign n13549 = ~n8314 & ~n9253;
  assign n13550 = pi090 & ~n13549;
  assign n13551 = ~pi090 & n8602;
  assign n13552 = ~n8323 & ~n13551;
  assign n13553 = ~n13550 & n13552;
  assign n13554 = ~n4349 & ~n4392;
  assign n13555 = n13553 & n13554;
  assign n13556 = ~pi088 & ~n13555;
  assign n13557 = pi090 & n4349;
  assign n13558 = n4395 & ~n8372;
  assign n13559 = ~pi090 & ~n13558;
  assign n13560 = ~n13557 & ~n13559;
  assign n13561 = ~n8453 & n13560;
  assign n13562 = ~n13556 & n13561;
  assign n13563 = ~n8547 & n13562;
  assign n13564 = ~n4289 & ~n9514;
  assign n13565 = ~n4299 & ~n8576;
  assign n13566 = n13564 & n13565;
  assign n13567 = pi088 & ~n13566;
  assign n13568 = pi049 & ~pi086;
  assign n13569 = ~pi051 & n13568;
  assign n13570 = pi019 & pi086;
  assign n13571 = ~pi049 & n13570;
  assign n13572 = ~n13569 & ~n13571;
  assign n13573 = ~n4388 & n13572;
  assign n13574 = n8387 & ~n13573;
  assign n13575 = ~n13567 & ~n13574;
  assign n13576 = ~n8525 & n13575;
  assign n13577 = n13563 & n13576;
  assign n13578 = pi006 & ~n13577;
  assign n13579 = pi019 & n4398;
  assign n13580 = pi019 & n8492;
  assign n13581 = ~n13579 & ~n13580;
  assign n13582 = ~n9472 & n13581;
  assign n13583 = ~n4344 & n13582;
  assign n13584 = pi090 & ~n13583;
  assign n13585 = n4322 & n4388;
  assign n13586 = n4297 & n8324;
  assign n13587 = ~n8603 & ~n13586;
  assign n13588 = ~pi019 & n8355;
  assign n13589 = n13587 & ~n13588;
  assign n13590 = ~n13585 & n13589;
  assign n13591 = ~pi088 & ~n13590;
  assign n13592 = ~n8306 & ~n9250;
  assign n13593 = pi090 & ~n13592;
  assign n13594 = ~n4434 & ~n8310;
  assign n13595 = ~pi019 & n4393;
  assign n13596 = n13594 & ~n13595;
  assign n13597 = ~pi090 & ~n13596;
  assign n13598 = ~n4365 & ~n4436;
  assign n13599 = ~n4391 & n13598;
  assign n13600 = ~n8364 & ~n13579;
  assign n13601 = n13599 & n13600;
  assign n13602 = ~n13597 & n13601;
  assign n13603 = ~n13593 & n13602;
  assign n13604 = pi088 & ~n13603;
  assign n13605 = ~n13591 & ~n13604;
  assign n13606 = ~n13584 & n13605;
  assign n13607 = ~pi090 & n4313;
  assign n13608 = n4328 & n13569;
  assign n13609 = ~n4337 & ~n13608;
  assign n13610 = ~n4361 & n13609;
  assign n13611 = ~n13607 & n13610;
  assign n13612 = n13606 & n13611;
  assign n13613 = ~pi006 & ~n13612;
  assign n13614 = ~pi019 & n4302;
  assign n13615 = ~n8412 & ~n13614;
  assign n13616 = ~n4311 & n13615;
  assign n13617 = ~pi090 & ~n13616;
  assign n13618 = n8304 & ~n8582;
  assign n13619 = ~n4349 & ~n13618;
  assign n13620 = pi090 & ~n13619;
  assign n13621 = n4322 & n8309;
  assign n13622 = ~n13620 & ~n13621;
  assign n13623 = ~n4345 & n13622;
  assign n13624 = ~n13617 & n13623;
  assign n13625 = ~pi088 & ~n13624;
  assign n13626 = ~n13613 & ~n13625;
  assign n13627 = ~n13578 & n13626;
  assign n13628 = n13548 & n13627;
  assign n13629 = ~pi141 & ~n13628;
  assign n13630 = pi141 & n13628;
  assign n13631 = ~n13629 & ~n13630;
  assign n13632 = ~n13540 & n13631;
  assign n13633 = n13540 & ~n13631;
  assign n13634 = ~n13632 & ~n13633;
  assign n13635 = ~n13348 & n13634;
  assign n13636 = n9366 & ~n13345;
  assign n13637 = ~n9366 & n13345;
  assign n13638 = ~n13636 & ~n13637;
  assign n13639 = ~n13634 & ~n13638;
  assign n13640 = ~n13635 & ~n13639;
  assign n13641 = ~pi529 & n13640;
  assign po176 = n13258 | n13641;
  assign n13643 = pi034 & n13349;
  assign n13644 = ~n5165 & ~n13352;
  assign n13645 = ~n8897 & n13644;
  assign n13646 = ~n13643 & n13645;
  assign n13647 = pi066 & n4661;
  assign n13648 = ~n4624 & ~n13647;
  assign n13649 = ~n4643 & n13648;
  assign n13650 = n4762 & ~n13649;
  assign n13651 = pi118 & n9312;
  assign n13652 = ~n4677 & ~n4706;
  assign n13653 = ~n4710 & n13652;
  assign n13654 = ~pi118 & ~n13653;
  assign n13655 = ~n5081 & ~n8913;
  assign n13656 = ~n4666 & n13655;
  assign n13657 = ~n13654 & n13656;
  assign n13658 = ~n13651 & n13657;
  assign n13659 = ~pi034 & ~n13658;
  assign n13660 = pi118 & n4714;
  assign n13661 = ~n13659 & ~n13660;
  assign n13662 = ~pi066 & n8888;
  assign n13663 = ~n5171 & ~n13662;
  assign n13664 = pi118 & ~n13663;
  assign n13665 = ~pi118 & n4759;
  assign n13666 = ~n5240 & ~n13665;
  assign n13667 = ~n13664 & n13666;
  assign n13668 = pi034 & ~n13667;
  assign n13669 = ~n5218 & ~n9326;
  assign n13670 = pi066 & pi119;
  assign n13671 = pi103 & n13670;
  assign n13672 = ~pi118 & n13671;
  assign n13673 = ~pi066 & n5140;
  assign n13674 = ~n13672 & ~n13673;
  assign n13675 = ~n4685 & n13674;
  assign n13676 = ~n4774 & n13675;
  assign n13677 = n13669 & n13676;
  assign n13678 = ~pi034 & ~n13677;
  assign n13679 = ~n13668 & ~n13678;
  assign n13680 = ~n4685 & ~n5114;
  assign n13681 = pi118 & ~n13680;
  assign n13682 = ~pi066 & n5267;
  assign n13683 = pi103 & n4676;
  assign n13684 = ~n13682 & ~n13683;
  assign n13685 = n5103 & ~n9278;
  assign n13686 = ~n4715 & ~n13685;
  assign n13687 = n13684 & n13686;
  assign n13688 = ~pi118 & ~n13687;
  assign n13689 = ~n13681 & ~n13688;
  assign n13690 = n13679 & n13689;
  assign n13691 = ~pi038 & ~n13690;
  assign n13692 = n13661 & ~n13691;
  assign n13693 = ~pi101 & pi103;
  assign n13694 = ~n4732 & ~n13693;
  assign n13695 = n5090 & ~n13694;
  assign n13696 = ~n4651 & ~n13695;
  assign n13697 = ~n4640 & n13696;
  assign n13698 = ~n4661 & ~n5180;
  assign n13699 = ~n4711 & n13698;
  assign n13700 = pi118 & ~n13699;
  assign n13701 = n13697 & ~n13700;
  assign n13702 = pi034 & ~n13701;
  assign n13703 = ~n4636 & ~n13671;
  assign n13704 = pi118 & ~n13703;
  assign n13705 = n4649 & n5090;
  assign n13706 = ~n4706 & ~n13705;
  assign n13707 = ~n13360 & n13706;
  assign n13708 = ~n13363 & n13707;
  assign n13709 = ~n13704 & n13708;
  assign n13710 = ~pi034 & ~n13709;
  assign n13711 = ~n13702 & ~n13710;
  assign n13712 = ~n4774 & ~n5262;
  assign n13713 = ~pi118 & ~n13712;
  assign n13714 = ~n4628 & ~n5169;
  assign n13715 = ~n4759 & n13714;
  assign n13716 = ~n8909 & n13715;
  assign n13717 = pi118 & ~n13716;
  assign n13718 = ~n13713 & ~n13717;
  assign n13719 = n13711 & n13718;
  assign n13720 = pi038 & ~n13719;
  assign n13721 = n13692 & ~n13720;
  assign n13722 = ~n13650 & n13721;
  assign n13723 = n13646 & n13722;
  assign n13724 = n4828 & n4928;
  assign n13725 = ~n5053 & ~n13724;
  assign n13726 = ~n8968 & n13725;
  assign n13727 = pi074 & n8983;
  assign n13728 = ~n9019 & ~n13727;
  assign n13729 = ~n4856 & n13728;
  assign n13730 = n4882 & ~n13729;
  assign n13731 = n13726 & ~n13730;
  assign n13732 = pi120 & n13321;
  assign n13733 = ~n4921 & ~n4975;
  assign n13734 = ~n5002 & n13733;
  assign n13735 = ~pi120 & ~n13734;
  assign n13736 = ~n5066 & ~n8977;
  assign n13737 = ~n9030 & n13736;
  assign n13738 = ~n13735 & n13737;
  assign n13739 = ~n13732 & n13738;
  assign n13740 = ~pi003 & ~n13739;
  assign n13741 = pi120 & n8955;
  assign n13742 = ~n13740 & ~n13741;
  assign n13743 = ~n4854 & ~n4896;
  assign n13744 = ~pi120 & ~n13743;
  assign n13745 = ~pi120 & n13123;
  assign n13746 = ~n4975 & ~n13745;
  assign n13747 = ~pi120 & n4798;
  assign n13748 = pi016 & n8958;
  assign n13749 = n8967 & n13748;
  assign n13750 = ~n13747 & ~n13749;
  assign n13751 = n13746 & n13750;
  assign n13752 = ~pi003 & ~n13751;
  assign n13753 = pi045 & pi074;
  assign n13754 = pi016 & n13753;
  assign n13755 = ~n4814 & ~n13754;
  assign n13756 = n4835 & ~n13755;
  assign n13757 = ~n13752 & ~n13756;
  assign n13758 = ~n4944 & ~n5009;
  assign n13759 = pi003 & ~n13758;
  assign n13760 = ~n4861 & ~n8983;
  assign n13761 = ~n13186 & n13760;
  assign n13762 = n4882 & ~n13761;
  assign n13763 = ~n13759 & ~n13762;
  assign n13764 = ~n4917 & ~n8962;
  assign n13765 = ~n8961 & n13764;
  assign n13766 = pi120 & ~n13765;
  assign n13767 = pi003 & n4890;
  assign n13768 = pi016 & ~pi041;
  assign n13769 = ~n4864 & ~n13768;
  assign n13770 = n13767 & ~n13769;
  assign n13771 = ~n13766 & ~n13770;
  assign n13772 = n13763 & n13771;
  assign n13773 = ~n5044 & n13772;
  assign n13774 = n13757 & n13773;
  assign n13775 = ~n13744 & n13774;
  assign n13776 = pi044 & ~n13775;
  assign n13777 = ~pi120 & n5045;
  assign n13778 = pi003 & n13777;
  assign n13779 = ~n4919 & ~n4973;
  assign n13780 = pi120 & ~n13779;
  assign n13781 = ~pi074 & n4865;
  assign n13782 = pi016 & n4997;
  assign n13783 = ~n13781 & ~n13782;
  assign n13784 = n4969 & ~n13297;
  assign n13785 = ~n8999 & ~n13784;
  assign n13786 = n13783 & n13785;
  assign n13787 = ~pi120 & ~n13786;
  assign n13788 = ~n13780 & ~n13787;
  assign n13789 = ~pi074 & n8959;
  assign n13790 = ~n4845 & ~n13789;
  assign n13791 = pi120 & ~n13790;
  assign n13792 = ~pi120 & n4917;
  assign n13793 = ~n4934 & ~n13792;
  assign n13794 = ~n13791 & n13793;
  assign n13795 = pi003 & ~n13794;
  assign n13796 = ~n4848 & ~n13292;
  assign n13797 = ~pi120 & n13754;
  assign n13798 = ~pi074 & n5018;
  assign n13799 = ~n13797 & ~n13798;
  assign n13800 = ~n4919 & n13799;
  assign n13801 = ~n4854 & n13800;
  assign n13802 = n13796 & n13801;
  assign n13803 = ~pi003 & ~n13802;
  assign n13804 = ~n13795 & ~n13803;
  assign n13805 = n13788 & n13804;
  assign n13806 = ~pi044 & ~n13805;
  assign n13807 = ~n13778 & ~n13806;
  assign n13808 = ~n13776 & n13807;
  assign n13809 = n13742 & n13808;
  assign n13810 = n13731 & n13809;
  assign n13811 = ~n13723 & n13810;
  assign n13812 = n13723 & ~n13810;
  assign n13813 = ~n13811 & ~n13812;
  assign n13814 = ~pi120 & n4975;
  assign n13815 = pi003 & n13814;
  assign n13816 = pi074 & n4917;
  assign n13817 = n4898 & n4928;
  assign n13818 = ~n13816 & ~n13817;
  assign n13819 = pi003 & ~n13818;
  assign n13820 = ~n13815 & ~n13819;
  assign n13821 = ~n4896 & ~n9029;
  assign n13822 = ~pi074 & n9042;
  assign n13823 = n13821 & ~n13822;
  assign n13824 = ~pi120 & ~n13823;
  assign n13825 = pi074 & n4844;
  assign n13826 = ~n9013 & ~n13825;
  assign n13827 = ~n4898 & ~n13282;
  assign n13828 = pi120 & ~n13827;
  assign n13829 = n13826 & ~n13828;
  assign n13830 = ~n13824 & n13829;
  assign n13831 = ~n4829 & ~n8983;
  assign n13832 = ~n4855 & n13831;
  assign n13833 = n13830 & n13832;
  assign n13834 = pi003 & ~n13833;
  assign n13835 = n4806 & n4901;
  assign n13836 = ~n8981 & ~n13835;
  assign n13837 = ~pi003 & ~n13836;
  assign n13838 = ~n4983 & ~n5046;
  assign n13839 = pi120 & ~n13838;
  assign n13840 = pi074 & n8959;
  assign n13841 = ~n13825 & ~n13840;
  assign n13842 = pi120 & ~n13841;
  assign n13843 = ~n13839 & ~n13842;
  assign n13844 = ~n4917 & ~n13749;
  assign n13845 = ~n13814 & n13844;
  assign n13846 = ~n13747 & n13845;
  assign n13847 = n13843 & n13846;
  assign n13848 = n4905 & n4972;
  assign n13849 = ~n13724 & ~n13848;
  assign n13850 = ~pi003 & ~n13849;
  assign n13851 = n13847 & ~n13850;
  assign n13852 = ~n13837 & n13851;
  assign n13853 = ~n13834 & n13852;
  assign n13854 = ~pi044 & ~n13853;
  assign n13855 = n4813 & n4905;
  assign n13856 = ~pi074 & n4943;
  assign n13857 = ~n4934 & ~n13856;
  assign n13858 = ~n4826 & n13857;
  assign n13859 = ~pi120 & ~n13858;
  assign n13860 = ~n13855 & ~n13859;
  assign n13861 = ~n9019 & n13860;
  assign n13862 = n4901 & ~n9027;
  assign n13863 = ~n8961 & ~n13862;
  assign n13864 = pi120 & ~n13863;
  assign n13865 = n13861 & ~n13864;
  assign n13866 = ~pi003 & ~n13865;
  assign n13867 = ~n13854 & ~n13866;
  assign n13868 = n13820 & n13867;
  assign n13869 = pi041 & pi074;
  assign n13870 = ~pi016 & n13869;
  assign n13871 = ~n13748 & ~n13870;
  assign n13872 = ~n4972 & n13871;
  assign n13873 = n13127 & ~n13872;
  assign n13874 = ~n8948 & ~n13873;
  assign n13875 = ~pi120 & n4826;
  assign n13876 = ~n4838 & n13178;
  assign n13877 = ~pi120 & ~n13876;
  assign n13878 = pi120 & n8961;
  assign n13879 = ~n13877 & ~n13878;
  assign n13880 = ~n9023 & n13879;
  assign n13881 = ~n13875 & n13880;
  assign n13882 = ~n4976 & ~n8946;
  assign n13883 = ~n5009 & ~n5019;
  assign n13884 = n13882 & n13883;
  assign n13885 = pi003 & ~n13884;
  assign n13886 = ~n4904 & ~n4960;
  assign n13887 = pi120 & ~n13886;
  assign n13888 = ~pi120 & n5043;
  assign n13889 = ~n13887 & ~n13888;
  assign n13890 = ~n4795 & ~n8961;
  assign n13891 = ~n4869 & n13890;
  assign n13892 = n13889 & n13891;
  assign n13893 = ~pi003 & ~n13892;
  assign n13894 = ~n13885 & ~n13893;
  assign n13895 = n13881 & n13894;
  assign n13896 = n13874 & n13895;
  assign n13897 = pi044 & ~n13896;
  assign n13898 = n13868 & ~n13897;
  assign n13899 = ~pi120 & n9013;
  assign n13900 = ~n5064 & ~n13899;
  assign n13901 = ~n13777 & n13900;
  assign n13902 = n13898 & n13901;
  assign n13903 = ~n13813 & n13902;
  assign n13904 = n13813 & ~n13902;
  assign n13905 = ~n13903 & ~n13904;
  assign n13906 = n4484 & n4528;
  assign n13907 = ~n9154 & ~n13906;
  assign n13908 = pi058 & n8802;
  assign n13909 = n13907 & ~n13908;
  assign n13910 = pi011 & n4588;
  assign n13911 = ~n4514 & ~n13910;
  assign n13912 = ~n4472 & n13911;
  assign n13913 = n4508 & ~n13912;
  assign n13914 = n13909 & ~n13913;
  assign n13915 = ~n4458 & ~n4469;
  assign n13916 = ~n4588 & ~n8681;
  assign n13917 = ~n4536 & n13916;
  assign n13918 = pi116 & ~n13917;
  assign n13919 = pi000 & ~pi022;
  assign n13920 = ~n4478 & ~n13919;
  assign n13921 = n8707 & ~n13920;
  assign n13922 = ~n13918 & ~n13921;
  assign n13923 = n13915 & n13922;
  assign n13924 = pi058 & ~n13923;
  assign n13925 = pi011 & pi097;
  assign n13926 = pi000 & n13925;
  assign n13927 = ~n4465 & ~n13926;
  assign n13928 = pi116 & ~n13927;
  assign n13929 = ~n4528 & ~n8840;
  assign n13930 = ~n13928 & n13929;
  assign n13931 = ~n13501 & n13930;
  assign n13932 = ~n13503 & n13931;
  assign n13933 = ~pi058 & ~n13932;
  assign n13934 = ~n13924 & ~n13933;
  assign n13935 = ~n4480 & ~n9432;
  assign n13936 = ~n4519 & n13935;
  assign n13937 = ~n9149 & n13936;
  assign n13938 = pi116 & ~n13937;
  assign n13939 = ~n4491 & ~n8673;
  assign n13940 = ~pi116 & ~n13939;
  assign n13941 = ~n13938 & ~n13940;
  assign n13942 = n13934 & n13941;
  assign n13943 = pi060 & ~n13942;
  assign n13944 = pi116 & n9438;
  assign n13945 = ~n4528 & ~n4595;
  assign n13946 = ~n4534 & n13945;
  assign n13947 = ~pi116 & ~n13946;
  assign n13948 = pi116 & n4525;
  assign n13949 = ~n9098 & ~n13948;
  assign n13950 = ~n4581 & n13949;
  assign n13951 = ~n13947 & n13950;
  assign n13952 = ~n13944 & n13951;
  assign n13953 = ~pi058 & ~n13952;
  assign n13954 = pi116 & n4542;
  assign n13955 = ~n13953 & ~n13954;
  assign n13956 = ~n13481 & n13955;
  assign n13957 = ~n13943 & n13956;
  assign n13958 = ~pi011 & n8791;
  assign n13959 = ~n8662 & ~n13958;
  assign n13960 = pi116 & ~n13959;
  assign n13961 = ~pi116 & n4480;
  assign n13962 = ~n13960 & ~n13961;
  assign n13963 = ~n8716 & n13962;
  assign n13964 = pi058 & ~n13963;
  assign n13965 = ~n4491 & ~n4501;
  assign n13966 = ~pi011 & n8773;
  assign n13967 = ~pi116 & n13926;
  assign n13968 = ~n13966 & ~n13967;
  assign n13969 = n13965 & n13968;
  assign n13970 = ~n9374 & n13969;
  assign n13971 = ~n8663 & n13970;
  assign n13972 = ~pi058 & ~n13971;
  assign n13973 = ~n13964 & ~n13972;
  assign n13974 = ~pi011 & n8684;
  assign n13975 = pi000 & n4594;
  assign n13976 = n8749 & ~n9368;
  assign n13977 = ~n13975 & ~n13976;
  assign n13978 = ~n4532 & n13977;
  assign n13979 = ~n13974 & n13978;
  assign n13980 = ~pi116 & ~n13979;
  assign n13981 = ~n4501 & ~n9081;
  assign n13982 = pi116 & ~n13981;
  assign n13983 = ~n13980 & ~n13982;
  assign n13984 = n13973 & n13983;
  assign n13985 = ~pi060 & ~n13984;
  assign n13986 = n13957 & ~n13985;
  assign n13987 = n13914 & n13986;
  assign n13988 = n13628 & ~n13987;
  assign n13989 = ~n13628 & n13987;
  assign n13990 = ~n13988 & ~n13989;
  assign n13991 = pi272 & n13990;
  assign n13992 = ~pi272 & ~n13990;
  assign n13993 = ~n13991 & ~n13992;
  assign n13994 = ~n13905 & n13993;
  assign n13995 = n13905 & ~n13993;
  assign n13996 = ~n13994 & ~n13995;
  assign n13997 = ~pi529 & ~n13996;
  assign n13998 = pi272 & pi511;
  assign n13999 = ~pi272 & ~pi511;
  assign n14000 = ~n13998 & ~n13999;
  assign n14001 = pi529 & n14000;
  assign po177 = n13997 | n14001;
  assign n14003 = ~pi130 & pi506;
  assign n14004 = pi130 & ~pi506;
  assign n14005 = ~n14003 & ~n14004;
  assign n14006 = pi529 & ~n14005;
  assign n14007 = ~pi066 & n5234;
  assign n14008 = ~n4684 & ~n14007;
  assign n14009 = n4762 & ~n14008;
  assign n14010 = pi118 & n4667;
  assign n14011 = n4770 & n14010;
  assign n14012 = ~n14009 & ~n14011;
  assign n14013 = ~pi118 & n4695;
  assign n14014 = n4629 & n5129;
  assign n14015 = ~n4686 & ~n14014;
  assign n14016 = ~pi118 & ~n14015;
  assign n14017 = ~n14013 & ~n14016;
  assign n14018 = ~n4657 & n14017;
  assign n14019 = pi034 & ~n14018;
  assign n14020 = ~n4649 & ~n4689;
  assign n14021 = n5078 & ~n14020;
  assign n14022 = pi118 & n14021;
  assign n14023 = ~n8928 & ~n14022;
  assign n14024 = ~n14019 & n14023;
  assign n14025 = pi103 & n4753;
  assign n14026 = n4656 & n14025;
  assign n14027 = ~n4692 & ~n8888;
  assign n14028 = ~n5134 & n14027;
  assign n14029 = ~pi118 & ~n14028;
  assign n14030 = ~n4677 & ~n14029;
  assign n14031 = ~n4724 & ~n5095;
  assign n14032 = pi118 & ~n14031;
  assign n14033 = n14030 & ~n14032;
  assign n14034 = pi034 & ~n14033;
  assign n14035 = ~n4706 & ~n13349;
  assign n14036 = n4669 & n8896;
  assign n14037 = ~n5171 & ~n14036;
  assign n14038 = ~pi034 & ~n14037;
  assign n14039 = n14035 & ~n14038;
  assign n14040 = ~n14034 & n14039;
  assign n14041 = ~n14026 & n14040;
  assign n14042 = ~pi038 & ~n14041;
  assign n14043 = n14024 & ~n14042;
  assign n14044 = pi118 & ~n4623;
  assign n14045 = pi062 & n5129;
  assign n14046 = ~n5267 & ~n14045;
  assign n14047 = ~pi118 & n14046;
  assign n14048 = ~n14044 & ~n14047;
  assign n14049 = ~n5185 & ~n14048;
  assign n14050 = pi034 & ~n14049;
  assign n14051 = pi118 & n5274;
  assign n14052 = ~pi118 & n4624;
  assign n14053 = ~n9346 & ~n14052;
  assign n14054 = ~n8855 & n14053;
  assign n14055 = ~n14051 & n14054;
  assign n14056 = ~n4773 & ~n5144;
  assign n14057 = ~n8935 & n14056;
  assign n14058 = ~n13397 & n14057;
  assign n14059 = n14055 & n14058;
  assign n14060 = ~pi034 & ~n14059;
  assign n14061 = ~n5178 & ~n14060;
  assign n14062 = ~n14050 & n14061;
  assign n14063 = ~n4720 & ~n5080;
  assign n14064 = ~n4650 & ~n4710;
  assign n14065 = ~n4626 & n14064;
  assign n14066 = n4753 & ~n14065;
  assign n14067 = n14063 & ~n14066;
  assign n14068 = n14062 & n14067;
  assign n14069 = pi038 & ~n14068;
  assign n14070 = pi066 & n4732;
  assign n14071 = ~n4705 & ~n14070;
  assign n14072 = ~n5171 & n14071;
  assign n14073 = pi118 & ~n14072;
  assign n14074 = ~n5163 & ~n5240;
  assign n14075 = ~n4666 & n14074;
  assign n14076 = ~pi118 & ~n14075;
  assign n14077 = pi066 & n5267;
  assign n14078 = ~n13705 & ~n14077;
  assign n14079 = ~n14076 & n14078;
  assign n14080 = ~n14073 & n14079;
  assign n14081 = ~n5122 & n14080;
  assign n14082 = ~pi034 & ~n14081;
  assign n14083 = ~n14069 & ~n14082;
  assign n14084 = n14043 & n14083;
  assign n14085 = n14012 & n14084;
  assign n14086 = n9054 & ~n14085;
  assign n14087 = ~n9054 & n14085;
  assign n14088 = ~n14086 & ~n14087;
  assign n14089 = ~n5298 & n8848;
  assign n14090 = n5298 & ~n8848;
  assign n14091 = ~n14089 & ~n14090;
  assign n14092 = n14088 & n14091;
  assign n14093 = ~n14088 & ~n14091;
  assign n14094 = ~n14092 & ~n14093;
  assign n14095 = ~pi130 & ~n8623;
  assign n14096 = pi130 & n8623;
  assign n14097 = ~n14095 & ~n14096;
  assign n14098 = pi000 & ~n13526;
  assign n14099 = ~n4581 & ~n14098;
  assign n14100 = pi116 & ~n14099;
  assign n14101 = ~n8689 & n9083;
  assign n14102 = ~pi116 & ~n14101;
  assign n14103 = ~pi011 & n4486;
  assign n14104 = ~n4527 & ~n14103;
  assign n14105 = ~n8738 & n14104;
  assign n14106 = pi116 & ~n14105;
  assign n14107 = ~n4532 & ~n14106;
  assign n14108 = ~n9138 & n14107;
  assign n14109 = ~n4528 & n14108;
  assign n14110 = ~n8662 & ~n8692;
  assign n14111 = n14109 & n14110;
  assign n14112 = pi058 & ~n14111;
  assign n14113 = ~n13442 & ~n14112;
  assign n14114 = ~n14102 & n14113;
  assign n14115 = ~n14100 & n14114;
  assign n14116 = ~n4514 & ~n9098;
  assign n14117 = ~n4466 & ~n4535;
  assign n14118 = ~pi116 & ~n14117;
  assign n14119 = pi116 & n8658;
  assign n14120 = ~n8771 & ~n14119;
  assign n14121 = ~n9150 & n14120;
  assign n14122 = ~n14118 & n14121;
  assign n14123 = n14116 & n14122;
  assign n14124 = ~n4462 & n14123;
  assign n14125 = ~pi058 & ~n14124;
  assign n14126 = n14115 & ~n14125;
  assign n14127 = pi060 & ~n14126;
  assign n14128 = n4481 & n8791;
  assign n14129 = ~n4519 & ~n9432;
  assign n14130 = ~pi116 & ~n14129;
  assign n14131 = ~pi011 & n4582;
  assign n14132 = ~n14130 & ~n14131;
  assign n14133 = ~n4472 & ~n8689;
  assign n14134 = pi116 & n9069;
  assign n14135 = ~n4467 & ~n4498;
  assign n14136 = n4540 & ~n14135;
  assign n14137 = ~n14134 & ~n14136;
  assign n14138 = n14133 & n14137;
  assign n14139 = ~n13906 & n14138;
  assign n14140 = ~pi058 & ~n14139;
  assign n14141 = ~n13948 & ~n14140;
  assign n14142 = n14132 & n14141;
  assign n14143 = ~n14128 & n14142;
  assign n14144 = ~pi116 & n4588;
  assign n14145 = ~n8791 & ~n13515;
  assign n14146 = pi116 & ~n14145;
  assign n14147 = ~n9149 & ~n9370;
  assign n14148 = ~n4608 & n14147;
  assign n14149 = ~n14146 & n14148;
  assign n14150 = ~n14144 & n14149;
  assign n14151 = pi058 & ~n14150;
  assign n14152 = n14143 & ~n14151;
  assign n14153 = ~pi060 & ~n14152;
  assign n14154 = pi116 & n4473;
  assign n14155 = ~n13462 & ~n14154;
  assign n14156 = ~pi058 & ~n14155;
  assign n14157 = n4481 & n4502;
  assign n14158 = ~n4483 & ~n14157;
  assign n14159 = ~n14156 & n14158;
  assign n14160 = ~n4542 & n14159;
  assign n14161 = n4503 & n8749;
  assign n14162 = ~n4532 & ~n14161;
  assign n14163 = pi116 & ~n14162;
  assign n14164 = ~n8825 & ~n9387;
  assign n14165 = ~n4547 & ~n4588;
  assign n14166 = ~n8684 & n14165;
  assign n14167 = n8707 & ~n14166;
  assign n14168 = n14164 & ~n14167;
  assign n14169 = ~n14163 & n14168;
  assign n14170 = pi058 & ~n14169;
  assign n14171 = n8780 & n13518;
  assign n14172 = ~n14170 & ~n14171;
  assign n14173 = n14160 & n14172;
  assign n14174 = ~n14153 & n14173;
  assign n14175 = ~n14127 & n14174;
  assign n14176 = ~n8748 & n14175;
  assign n14177 = n8748 & ~n14175;
  assign n14178 = ~n14176 & ~n14177;
  assign n14179 = n14097 & ~n14178;
  assign n14180 = ~n14097 & n14178;
  assign n14181 = ~n14179 & ~n14180;
  assign n14182 = ~n14094 & n14181;
  assign n14183 = n14094 & ~n14181;
  assign n14184 = ~n14182 & ~n14183;
  assign n14185 = ~pi529 & n14184;
  assign po178 = n14006 | n14185;
  assign n14187 = pi160 & pi472;
  assign n14188 = ~pi160 & ~pi472;
  assign n14189 = ~n14187 & ~n14188;
  assign n14190 = pi529 & n14189;
  assign n14191 = ~pi160 & ~n9554;
  assign n14192 = pi160 & n9554;
  assign n14193 = ~n14191 & ~n14192;
  assign n14194 = ~n4957 & n5298;
  assign n14195 = n4957 & ~n5298;
  assign n14196 = ~n14194 & ~n14195;
  assign n14197 = ~n9165 & n14196;
  assign n14198 = ~n9163 & ~n14196;
  assign n14199 = ~n9164 & n14198;
  assign n14200 = ~n14197 & ~n14199;
  assign n14201 = n14193 & n14200;
  assign n14202 = ~n14193 & ~n14200;
  assign n14203 = ~n14201 & ~n14202;
  assign n14204 = ~pi529 & n14203;
  assign po179 = n14190 | n14204;
  assign n14206 = n5298 & ~n8748;
  assign n14207 = ~n5298 & n8748;
  assign n14208 = ~n14206 & ~n14207;
  assign n14209 = ~pi161 & ~n8423;
  assign n14210 = pi161 & n8423;
  assign n14211 = ~n14209 & ~n14210;
  assign n14212 = ~n14208 & n14211;
  assign n14213 = n14208 & ~n14211;
  assign n14214 = ~n14212 & ~n14213;
  assign n14215 = n13813 & ~n14214;
  assign n14216 = ~n13813 & n14214;
  assign n14217 = ~n14215 & ~n14216;
  assign n14218 = ~pi529 & ~n14217;
  assign n14219 = ~pi161 & pi409;
  assign n14220 = pi161 & ~pi409;
  assign n14221 = ~n14219 & ~n14220;
  assign n14222 = pi529 & ~n14221;
  assign po180 = n14218 | n14222;
  assign n14224 = ~pi106 & n6175;
  assign n14225 = pi035 & n9852;
  assign n14226 = ~n14224 & ~n14225;
  assign n14227 = pi065 & ~n14226;
  assign n14228 = n6608 & n9872;
  assign n14229 = ~pi106 & n6311;
  assign n14230 = ~n14228 & ~n14229;
  assign n14231 = ~n14227 & n14230;
  assign n14232 = ~n7097 & n14231;
  assign n14233 = ~n11156 & n14232;
  assign n14234 = ~pi035 & n6252;
  assign n14235 = ~n6308 & ~n14234;
  assign n14236 = ~n6220 & n14235;
  assign n14237 = n6654 & ~n14236;
  assign n14238 = n6320 & n9807;
  assign n14239 = n6164 & ~n6595;
  assign n14240 = ~n6630 & ~n14239;
  assign n14241 = pi106 & ~n14240;
  assign n14242 = ~n14238 & ~n14241;
  assign n14243 = ~n6566 & n14242;
  assign n14244 = ~pi065 & ~n14243;
  assign n14245 = ~n14237 & ~n14244;
  assign n14246 = n14233 & n14245;
  assign n14247 = ~n6571 & n10711;
  assign n14248 = ~pi106 & ~n14247;
  assign n14249 = pi106 & n6630;
  assign n14250 = ~n6553 & ~n14249;
  assign n14251 = ~n11131 & n14250;
  assign n14252 = ~n14248 & n14251;
  assign n14253 = pi037 & n6268;
  assign n14254 = pi031 & n6609;
  assign n14255 = ~n14253 & ~n14254;
  assign n14256 = ~n7005 & n14255;
  assign n14257 = pi065 & ~n14256;
  assign n14258 = ~pi106 & n14257;
  assign n14259 = ~n6556 & ~n7053;
  assign n14260 = ~n6261 & ~n7040;
  assign n14261 = n14259 & n14260;
  assign n14262 = pi065 & ~n14261;
  assign n14263 = ~n14258 & ~n14262;
  assign n14264 = n14252 & n14263;
  assign n14265 = ~n6301 & ~n6630;
  assign n14266 = n6191 & n6246;
  assign n14267 = ~n6210 & ~n14266;
  assign n14268 = pi106 & ~n14267;
  assign n14269 = ~pi106 & n6279;
  assign n14270 = ~n14268 & ~n14269;
  assign n14271 = n14265 & n14270;
  assign n14272 = ~n9885 & n14271;
  assign n14273 = ~pi065 & ~n14272;
  assign n14274 = ~n6547 & ~n14273;
  assign n14275 = n14264 & n14274;
  assign n14276 = pi068 & ~n14275;
  assign n14277 = n6617 & n14254;
  assign n14278 = ~pi031 & ~pi106;
  assign n14279 = ~pi037 & n14278;
  assign n14280 = n6165 & n14279;
  assign n14281 = ~n14224 & ~n14280;
  assign n14282 = ~n9852 & n14281;
  assign n14283 = ~n14277 & n14282;
  assign n14284 = n6184 & n6197;
  assign n14285 = ~n6228 & ~n14284;
  assign n14286 = ~pi035 & n6263;
  assign n14287 = n6320 & n7005;
  assign n14288 = ~n14286 & ~n14287;
  assign n14289 = n14285 & n14288;
  assign n14290 = ~pi065 & ~n14289;
  assign n14291 = ~n6245 & ~n6307;
  assign n14292 = pi106 & ~n14291;
  assign n14293 = ~n6597 & ~n9861;
  assign n14294 = ~pi035 & n6262;
  assign n14295 = n14293 & ~n14294;
  assign n14296 = ~pi106 & ~n14295;
  assign n14297 = ~n6311 & ~n6603;
  assign n14298 = ~n9824 & n14297;
  assign n14299 = pi035 & n6584;
  assign n14300 = ~n7075 & ~n14299;
  assign n14301 = n14298 & n14300;
  assign n14302 = ~n14296 & n14301;
  assign n14303 = ~n14292 & n14302;
  assign n14304 = pi065 & ~n14303;
  assign n14305 = ~n6195 & ~n7079;
  assign n14306 = pi035 & n6610;
  assign n14307 = ~n14299 & ~n14306;
  assign n14308 = n14305 & n14307;
  assign n14309 = pi106 & ~n14308;
  assign n14310 = ~n14304 & ~n14309;
  assign n14311 = ~n14290 & n14310;
  assign n14312 = n14283 & n14311;
  assign n14313 = ~pi068 & ~n14312;
  assign n14314 = ~n14276 & ~n14313;
  assign n14315 = n14246 & n14314;
  assign n14316 = ~pi122 & n5384;
  assign n14317 = ~pi043 & n5383;
  assign n14318 = ~n5337 & ~n14317;
  assign n14319 = pi122 & ~n14318;
  assign n14320 = ~n14316 & ~n14319;
  assign n14321 = ~n5377 & n14320;
  assign n14322 = pi039 & ~n14321;
  assign n14323 = ~n5340 & ~n6065;
  assign n14324 = ~pi043 & n6142;
  assign n14325 = pi043 & pi109;
  assign n14326 = pi076 & n14325;
  assign n14327 = ~pi122 & n14326;
  assign n14328 = ~n5358 & ~n5491;
  assign n14329 = ~n14327 & n14328;
  assign n14330 = ~n14324 & n14329;
  assign n14331 = n14323 & n14330;
  assign n14332 = ~pi039 & ~n14331;
  assign n14333 = ~n14322 & ~n14332;
  assign n14334 = ~n5358 & ~n7128;
  assign n14335 = pi122 & ~n14334;
  assign n14336 = ~pi043 & n5413;
  assign n14337 = pi076 & n6100;
  assign n14338 = ~n14336 & ~n14337;
  assign n14339 = n5596 & ~n6113;
  assign n14340 = ~n5493 & ~n14339;
  assign n14341 = n14338 & n14340;
  assign n14342 = ~pi122 & ~n14341;
  assign n14343 = ~n14335 & ~n14342;
  assign n14344 = n14333 & n14343;
  assign n14345 = ~pi017 & ~n14344;
  assign n14346 = pi043 & n5556;
  assign n14347 = ~n5513 & ~n14346;
  assign n14348 = ~n5323 & n14347;
  assign n14349 = n5456 & ~n14348;
  assign n14350 = ~n5409 & ~n5556;
  assign n14351 = ~n10614 & n14350;
  assign n14352 = pi122 & ~n14351;
  assign n14353 = ~pi070 & pi076;
  assign n14354 = ~n5412 & ~n14353;
  assign n14355 = n5444 & ~n14354;
  assign n14356 = ~n14352 & ~n14355;
  assign n14357 = n7136 & n14356;
  assign n14358 = pi039 & ~n14357;
  assign n14359 = ~n5368 & ~n14326;
  assign n14360 = pi122 & ~n14359;
  assign n14361 = pi076 & n5382;
  assign n14362 = n5538 & n14361;
  assign n14363 = ~pi122 & n5464;
  assign n14364 = ~n5486 & ~n6423;
  assign n14365 = ~n14363 & n14364;
  assign n14366 = ~n14362 & n14365;
  assign n14367 = ~n14360 & n14366;
  assign n14368 = ~pi039 & ~n14367;
  assign n14369 = ~n14358 & ~n14368;
  assign n14370 = ~n5384 & ~n5535;
  assign n14371 = ~n5534 & n14370;
  assign n14372 = ~n5517 & n14371;
  assign n14373 = pi122 & ~n14372;
  assign n14374 = ~n5432 & ~n5491;
  assign n14375 = ~pi122 & ~n14374;
  assign n14376 = ~n14373 & ~n14375;
  assign n14377 = n14369 & n14376;
  assign n14378 = pi017 & ~n14377;
  assign n14379 = n5322 & n5362;
  assign n14380 = pi039 & n6140;
  assign n14381 = ~pi122 & n14380;
  assign n14382 = ~n5539 & ~n14381;
  assign n14383 = ~n6116 & n14382;
  assign n14384 = ~n14379 & n14383;
  assign n14385 = pi122 & n5570;
  assign n14386 = pi122 & n6097;
  assign n14387 = ~n5360 & ~n5486;
  assign n14388 = ~n6407 & n14387;
  assign n14389 = ~pi122 & ~n14388;
  assign n14390 = ~n5511 & ~n5551;
  assign n14391 = ~n5527 & n14390;
  assign n14392 = ~n14389 & n14391;
  assign n14393 = ~n14386 & n14392;
  assign n14394 = ~pi039 & ~n14393;
  assign n14395 = ~n14385 & ~n14394;
  assign n14396 = n14384 & n14395;
  assign n14397 = ~n14378 & n14396;
  assign n14398 = ~n14349 & n14397;
  assign n14399 = ~n14345 & n14398;
  assign n14400 = pi005 & n5850;
  assign n14401 = ~n5806 & ~n14400;
  assign n14402 = ~n5624 & n14401;
  assign n14403 = n5697 & ~n14402;
  assign n14404 = pi024 & n6522;
  assign n14405 = ~n5742 & ~n10476;
  assign n14406 = ~pi004 & n5621;
  assign n14407 = ~pi005 & n6493;
  assign n14408 = pi094 & n5796;
  assign n14409 = ~pi091 & n14408;
  assign n14410 = ~n14407 & ~n14409;
  assign n14411 = ~n5652 & n14410;
  assign n14412 = ~n14406 & n14411;
  assign n14413 = n14405 & n14412;
  assign n14414 = ~pi024 & ~n14413;
  assign n14415 = ~n5652 & ~n6923;
  assign n14416 = pi091 & ~n14415;
  assign n14417 = pi004 & n6965;
  assign n14418 = ~pi005 & n5676;
  assign n14419 = n5811 & ~n10478;
  assign n14420 = ~n14418 & ~n14419;
  assign n14421 = ~n14417 & n14420;
  assign n14422 = ~n5774 & n14421;
  assign n14423 = ~pi091 & ~n14422;
  assign n14424 = ~n14416 & ~n14423;
  assign n14425 = ~pi091 & n5610;
  assign n14426 = ~pi005 & n5831;
  assign n14427 = ~n5746 & ~n14426;
  assign n14428 = pi091 & ~n14427;
  assign n14429 = ~n14425 & ~n14428;
  assign n14430 = ~n5623 & n14429;
  assign n14431 = pi024 & ~n14430;
  assign n14432 = n14424 & ~n14431;
  assign n14433 = ~n14414 & n14432;
  assign n14434 = ~pi018 & ~n14433;
  assign n14435 = ~n14404 & ~n14434;
  assign n14436 = ~n5715 & ~n14406;
  assign n14437 = ~pi091 & ~n14436;
  assign n14438 = ~n5659 & ~n14408;
  assign n14439 = n5736 & ~n14438;
  assign n14440 = pi004 & n5830;
  assign n14441 = n5836 & n14440;
  assign n14442 = ~n5773 & ~n6464;
  assign n14443 = ~pi091 & n5752;
  assign n14444 = n14442 & ~n14443;
  assign n14445 = ~n14441 & n14444;
  assign n14446 = ~pi024 & ~n14445;
  assign n14447 = ~n14439 & ~n14446;
  assign n14448 = ~n5632 & ~n6957;
  assign n14449 = pi024 & ~n14448;
  assign n14450 = ~n5673 & ~n5850;
  assign n14451 = ~pi004 & n5798;
  assign n14452 = n14450 & ~n14451;
  assign n14453 = n5697 & ~n14452;
  assign n14454 = ~n14449 & ~n14453;
  assign n14455 = ~n5610 & ~n5826;
  assign n14456 = ~n5825 & n14455;
  assign n14457 = pi091 & ~n14456;
  assign n14458 = pi024 & n5705;
  assign n14459 = pi004 & ~pi084;
  assign n14460 = ~n5608 & ~n14459;
  assign n14461 = n14458 & ~n14460;
  assign n14462 = ~n14457 & ~n14461;
  assign n14463 = n14454 & n14462;
  assign n14464 = ~n5795 & n14463;
  assign n14465 = n14447 & n14464;
  assign n14466 = ~n14437 & n14465;
  assign n14467 = pi018 & ~n14466;
  assign n14468 = ~n5807 & ~n5819;
  assign n14469 = ~n5655 & ~n5773;
  assign n14470 = ~n6475 & n14469;
  assign n14471 = ~pi091 & ~n14470;
  assign n14472 = pi091 & n10537;
  assign n14473 = ~n5829 & ~n14472;
  assign n14474 = ~n14471 & n14473;
  assign n14475 = n14468 & n14474;
  assign n14476 = ~pi024 & ~n14475;
  assign n14477 = pi091 & n5891;
  assign n14478 = ~n14476 & ~n14477;
  assign n14479 = n5609 & n5663;
  assign n14480 = n14478 & ~n14479;
  assign n14481 = ~n14467 & n14480;
  assign n14482 = n14435 & n14481;
  assign n14483 = ~n14403 & n14482;
  assign n14484 = ~n5837 & ~n6980;
  assign n14485 = n14483 & n14484;
  assign n14486 = n14399 & n14485;
  assign n14487 = ~n14399 & ~n14485;
  assign n14488 = ~n14486 & ~n14487;
  assign n14489 = ~n14315 & ~n14488;
  assign n14490 = ~n14399 & n14485;
  assign n14491 = n14399 & ~n14485;
  assign n14492 = ~n14490 & ~n14491;
  assign n14493 = n14315 & ~n14492;
  assign n14494 = ~n14489 & ~n14493;
  assign n14495 = ~pi009 & n6013;
  assign n14496 = ~n6047 & ~n14495;
  assign n14497 = ~n5925 & n14496;
  assign n14498 = ~pi113 & ~n14497;
  assign n14499 = n5994 & ~n6675;
  assign n14500 = ~n6723 & ~n14499;
  assign n14501 = pi113 & ~n14500;
  assign n14502 = n5938 & n6855;
  assign n14503 = ~n14501 & ~n14502;
  assign n14504 = ~n6691 & n14503;
  assign n14505 = ~n14498 & n14504;
  assign n14506 = ~pi096 & ~n14505;
  assign n14507 = n6734 & n6842;
  assign n14508 = ~n9701 & ~n14507;
  assign n14509 = ~n9622 & n14508;
  assign n14510 = ~n6694 & n14509;
  assign n14511 = ~pi113 & n5951;
  assign n14512 = pi009 & n10808;
  assign n14513 = ~n14511 & ~n14512;
  assign n14514 = pi096 & ~n14513;
  assign n14515 = n14510 & ~n14514;
  assign n14516 = pi009 & n6708;
  assign n14517 = ~n5969 & ~n14516;
  assign n14518 = pi009 & n6718;
  assign n14519 = n14517 & ~n14518;
  assign n14520 = ~n9631 & n14519;
  assign n14521 = pi113 & ~n14520;
  assign n14522 = n5916 & n5958;
  assign n14523 = ~n5913 & ~n14522;
  assign n14524 = ~pi009 & n6004;
  assign n14525 = n5938 & n10837;
  assign n14526 = ~n14524 & ~n14525;
  assign n14527 = n14523 & n14526;
  assign n14528 = ~pi096 & ~n14527;
  assign n14529 = ~n6019 & ~n6046;
  assign n14530 = pi113 & ~n14529;
  assign n14531 = ~n6673 & ~n6870;
  assign n14532 = ~pi009 & n6003;
  assign n14533 = n14531 & ~n14532;
  assign n14534 = ~pi113 & ~n14533;
  assign n14535 = ~n6844 & ~n6848;
  assign n14536 = ~n6730 & n14535;
  assign n14537 = ~n6053 & ~n14516;
  assign n14538 = n14536 & n14537;
  assign n14539 = ~n14534 & n14538;
  assign n14540 = ~n14530 & n14539;
  assign n14541 = pi096 & ~n14540;
  assign n14542 = ~n14528 & ~n14541;
  assign n14543 = ~n14521 & n14542;
  assign n14544 = ~pi025 & n6809;
  assign n14545 = n5910 & n14544;
  assign n14546 = pi125 & n6717;
  assign n14547 = n6685 & n14546;
  assign n14548 = ~n14511 & ~n14547;
  assign n14549 = ~n10808 & n14548;
  assign n14550 = ~n14545 & n14549;
  assign n14551 = n14543 & n14550;
  assign n14552 = pi010 & ~n14551;
  assign n14553 = pi025 & n5989;
  assign n14554 = ~n14546 & ~n14553;
  assign n14555 = ~n10837 & n14554;
  assign n14556 = n6854 & ~n14555;
  assign n14557 = pi113 & n6723;
  assign n14558 = ~n6682 & n10830;
  assign n14559 = ~pi113 & ~n14558;
  assign n14560 = ~n14557 & ~n14559;
  assign n14561 = ~n6672 & n14560;
  assign n14562 = ~n6000 & ~n6666;
  assign n14563 = ~n9576 & ~n9587;
  assign n14564 = n14562 & n14563;
  assign n14565 = pi096 & ~n14564;
  assign n14566 = ~n5946 & ~n14565;
  assign n14567 = n14561 & n14566;
  assign n14568 = ~n14556 & n14567;
  assign n14569 = ~n6041 & ~n6723;
  assign n14570 = ~n5980 & ~n6017;
  assign n14571 = pi113 & ~n14570;
  assign n14572 = ~pi113 & n5991;
  assign n14573 = ~n6881 & ~n14572;
  assign n14574 = ~n14571 & n14573;
  assign n14575 = n14569 & n14574;
  assign n14576 = ~pi096 & ~n14575;
  assign n14577 = ~n6778 & ~n14576;
  assign n14578 = n14568 & n14577;
  assign n14579 = ~pi010 & ~n14578;
  assign n14580 = ~n14552 & ~n14579;
  assign n14581 = n14515 & n14580;
  assign n14582 = ~n14506 & n14581;
  assign n14583 = pi096 & n9701;
  assign n14584 = ~n5918 & ~n14583;
  assign n14585 = ~n14522 & n14584;
  assign n14586 = ~n6740 & n14585;
  assign n14587 = pi009 & n6730;
  assign n14588 = ~n6691 & ~n14587;
  assign n14589 = ~n5999 & n14588;
  assign n14590 = n6842 & ~n14589;
  assign n14591 = ~n5903 & ~n6730;
  assign n14592 = ~n10822 & n14591;
  assign n14593 = pi113 & ~n14592;
  assign n14594 = ~pi025 & pi125;
  assign n14595 = ~n6756 & ~n14594;
  assign n14596 = n5966 & ~n14595;
  assign n14597 = ~n14593 & ~n14596;
  assign n14598 = n9577 & n14597;
  assign n14599 = pi096 & ~n14598;
  assign n14600 = pi124 & n5978;
  assign n14601 = ~n5940 & ~n14600;
  assign n14602 = pi113 & ~n14601;
  assign n14603 = ~n9751 & ~n14547;
  assign n14604 = ~n14602 & n14603;
  assign n14605 = ~n14545 & n14604;
  assign n14606 = ~n5951 & n14605;
  assign n14607 = ~pi096 & ~n14606;
  assign n14608 = ~n14599 & ~n14607;
  assign n14609 = ~n6671 & ~n6870;
  assign n14610 = ~pi113 & ~n14609;
  assign n14611 = ~n5956 & ~n10808;
  assign n14612 = ~n6723 & n14611;
  assign n14613 = ~n5991 & n14612;
  assign n14614 = pi113 & ~n14613;
  assign n14615 = ~n14610 & ~n14614;
  assign n14616 = n14608 & n14615;
  assign n14617 = ~pi010 & ~n14616;
  assign n14618 = ~pi113 & n10808;
  assign n14619 = ~pi009 & n6718;
  assign n14620 = ~n6709 & ~n14619;
  assign n14621 = pi113 & ~n14620;
  assign n14622 = ~n14618 & ~n14621;
  assign n14623 = ~n6047 & n14622;
  assign n14624 = pi096 & ~n14623;
  assign n14625 = ~n5923 & ~n6861;
  assign n14626 = ~pi009 & n6007;
  assign n14627 = ~pi113 & n14600;
  assign n14628 = ~n14626 & ~n14627;
  assign n14629 = ~n6671 & n14628;
  assign n14630 = ~n6830 & n14629;
  assign n14631 = n14625 & n14630;
  assign n14632 = ~pi096 & ~n14631;
  assign n14633 = ~n14624 & ~n14632;
  assign n14634 = ~pi009 & n6757;
  assign n14635 = pi125 & n9593;
  assign n14636 = ~n5908 & n5989;
  assign n14637 = ~n6027 & ~n14636;
  assign n14638 = ~n14635 & n14637;
  assign n14639 = ~n14634 & n14638;
  assign n14640 = ~pi113 & ~n14639;
  assign n14641 = ~n6830 & ~n9649;
  assign n14642 = pi113 & ~n14641;
  assign n14643 = ~n14640 & ~n14642;
  assign n14644 = n14633 & n14643;
  assign n14645 = pi010 & ~n14644;
  assign n14646 = pi113 & n5970;
  assign n14647 = ~n5951 & ~n6825;
  assign n14648 = ~n6770 & n14647;
  assign n14649 = ~pi113 & ~n14648;
  assign n14650 = ~n6692 & ~n6720;
  assign n14651 = ~n6674 & n14650;
  assign n14652 = ~n14649 & n14651;
  assign n14653 = ~n14646 & n14652;
  assign n14654 = ~pi096 & ~n14653;
  assign n14655 = pi113 & n6771;
  assign n14656 = ~n14654 & ~n14655;
  assign n14657 = ~n14645 & n14656;
  assign n14658 = ~n14617 & n14657;
  assign n14659 = ~n14590 & n14658;
  assign n14660 = n14586 & n14659;
  assign n14661 = ~pi215 & ~n14660;
  assign n14662 = pi215 & n14660;
  assign n14663 = ~n14661 & ~n14662;
  assign n14664 = n14582 & n14663;
  assign n14665 = ~n14582 & ~n14663;
  assign n14666 = ~n14664 & ~n14665;
  assign n14667 = ~n14494 & ~n14666;
  assign n14668 = n14494 & n14666;
  assign n14669 = ~n14667 & ~n14668;
  assign n14670 = ~pi529 & ~n14669;
  assign n14671 = ~pi215 & pi401;
  assign n14672 = pi215 & ~pi401;
  assign n14673 = ~n14671 & ~n14672;
  assign n14674 = pi529 & ~n14673;
  assign po181 = n14670 | n14674;
  assign n14676 = ~pi122 & n5507;
  assign n14677 = ~n6356 & ~n7185;
  assign n14678 = ~n5463 & ~n5534;
  assign n14679 = ~n5440 & ~n6131;
  assign n14680 = pi122 & ~n14679;
  assign n14681 = ~pi122 & n5517;
  assign n14682 = ~n14680 & ~n14681;
  assign n14683 = n14678 & n14682;
  assign n14684 = ~n5417 & n14683;
  assign n14685 = ~pi039 & ~n14684;
  assign n14686 = ~n5573 & ~n14685;
  assign n14687 = ~n5328 & n10631;
  assign n14688 = ~pi122 & ~n14687;
  assign n14689 = pi122 & n5534;
  assign n14690 = ~n6390 & ~n14689;
  assign n14691 = ~n5492 & n14690;
  assign n14692 = ~n14688 & n14691;
  assign n14693 = pi043 & pi070;
  assign n14694 = ~pi076 & n14693;
  assign n14695 = ~n7127 & ~n14694;
  assign n14696 = ~n14361 & n14695;
  assign n14697 = pi039 & ~n14696;
  assign n14698 = ~pi122 & n14697;
  assign n14699 = ~n7135 & ~n7147;
  assign n14700 = ~n5487 & ~n5571;
  assign n14701 = n14699 & n14700;
  assign n14702 = pi039 & ~n14701;
  assign n14703 = ~n14698 & ~n14702;
  assign n14704 = n14692 & n14703;
  assign n14705 = n14686 & n14704;
  assign n14706 = pi017 & ~n14705;
  assign n14707 = ~n5560 & ~n14379;
  assign n14708 = ~pi043 & n5466;
  assign n14709 = n5381 & n7127;
  assign n14710 = ~n14708 & ~n14709;
  assign n14711 = n14707 & n14710;
  assign n14712 = ~pi039 & ~n14711;
  assign n14713 = ~pi122 & n5486;
  assign n14714 = ~n14363 & ~n14713;
  assign n14715 = ~n5384 & n14714;
  assign n14716 = ~n14362 & n14715;
  assign n14717 = ~n5432 & ~n5526;
  assign n14718 = ~pi043 & n5582;
  assign n14719 = n14717 & ~n14718;
  assign n14720 = ~pi122 & ~n14719;
  assign n14721 = pi043 & n5336;
  assign n14722 = ~n5507 & ~n14721;
  assign n14723 = ~n5376 & ~n6133;
  assign n14724 = pi122 & ~n14723;
  assign n14725 = n14722 & ~n14724;
  assign n14726 = ~n14720 & n14725;
  assign n14727 = ~n5348 & ~n5556;
  assign n14728 = ~n5320 & n14727;
  assign n14729 = n14726 & n14728;
  assign n14730 = pi039 & ~n14729;
  assign n14731 = ~n5512 & ~n14721;
  assign n14732 = pi043 & n5383;
  assign n14733 = n5368 & n5438;
  assign n14734 = ~n14732 & ~n14733;
  assign n14735 = n14731 & n14734;
  assign n14736 = pi122 & ~n14735;
  assign n14737 = ~n14730 & ~n14736;
  assign n14738 = n14716 & n14737;
  assign n14739 = ~n14712 & n14738;
  assign n14740 = ~pi017 & ~n14739;
  assign n14741 = ~n14706 & ~n14740;
  assign n14742 = ~pi043 & n5400;
  assign n14743 = ~n5346 & ~n14742;
  assign n14744 = ~n5377 & n14743;
  assign n14745 = n5593 & ~n14744;
  assign n14746 = n5381 & n5431;
  assign n14747 = n5438 & ~n5528;
  assign n14748 = ~n5534 & ~n14747;
  assign n14749 = pi122 & ~n14748;
  assign n14750 = ~n14746 & ~n14749;
  assign n14751 = ~n5513 & n14750;
  assign n14752 = ~pi039 & ~n14751;
  assign n14753 = pi043 & n5384;
  assign n14754 = ~n14713 & ~n14753;
  assign n14755 = pi039 & ~n14754;
  assign n14756 = n5456 & n5562;
  assign n14757 = ~n14755 & ~n14756;
  assign n14758 = ~n14752 & n14757;
  assign n14759 = ~n14745 & n14758;
  assign n14760 = n14741 & n14759;
  assign n14761 = n14677 & n14760;
  assign n14762 = ~n14676 & n14761;
  assign n14763 = ~n14485 & n14762;
  assign n14764 = n14485 & ~n14762;
  assign n14765 = ~n14763 & ~n14764;
  assign n14766 = n14315 & n14765;
  assign n14767 = ~n14315 & ~n14765;
  assign n14768 = ~n14766 & ~n14767;
  assign n14769 = ~n6232 & ~n6618;
  assign n14770 = pi065 & n11156;
  assign n14771 = n14769 & ~n14770;
  assign n14772 = pi035 & n6603;
  assign n14773 = ~n6212 & ~n14772;
  assign n14774 = ~n6566 & n14773;
  assign n14775 = n9872 & ~n14774;
  assign n14776 = n14771 & ~n14775;
  assign n14777 = pi106 & n6196;
  assign n14778 = ~n6565 & ~n6598;
  assign n14779 = ~n6175 & ~n9817;
  assign n14780 = ~n6540 & n14779;
  assign n14781 = ~pi106 & ~n14780;
  assign n14782 = ~n6633 & ~n14781;
  assign n14783 = n14778 & n14782;
  assign n14784 = ~n14777 & n14783;
  assign n14785 = ~pi065 & ~n14784;
  assign n14786 = pi106 & n6541;
  assign n14787 = ~n14785 & ~n14786;
  assign n14788 = ~n14284 & n14787;
  assign n14789 = pi031 & ~pi037;
  assign n14790 = ~n6647 & ~n14789;
  assign n14791 = n6645 & ~n14790;
  assign n14792 = n7042 & ~n14791;
  assign n14793 = ~n6603 & ~n10718;
  assign n14794 = ~n6181 & n14793;
  assign n14795 = pi106 & ~n14794;
  assign n14796 = n14792 & ~n14795;
  assign n14797 = pi065 & ~n14796;
  assign n14798 = ~n6175 & ~n14277;
  assign n14799 = pi128 & n6246;
  assign n14800 = ~n6322 & ~n14799;
  assign n14801 = pi106 & ~n14800;
  assign n14802 = n14798 & ~n14801;
  assign n14803 = ~n14280 & n14802;
  assign n14804 = ~n11122 & n14803;
  assign n14805 = ~pi065 & ~n14804;
  assign n14806 = ~n14797 & ~n14805;
  assign n14807 = ~n6182 & ~n6279;
  assign n14808 = ~n6630 & n14807;
  assign n14809 = ~n9852 & n14808;
  assign n14810 = pi106 & ~n14809;
  assign n14811 = ~n6552 & ~n9861;
  assign n14812 = ~pi106 & ~n14811;
  assign n14813 = ~n14810 & ~n14812;
  assign n14814 = n14806 & n14813;
  assign n14815 = pi068 & ~n14814;
  assign n14816 = n14788 & ~n14815;
  assign n14817 = ~pi106 & n9852;
  assign n14818 = ~pi035 & n6610;
  assign n14819 = ~n6585 & ~n14818;
  assign n14820 = pi106 & ~n14819;
  assign n14821 = ~n14817 & ~n14820;
  assign n14822 = ~n6308 & n14821;
  assign n14823 = pi065 & ~n14822;
  assign n14824 = ~n6167 & ~n6552;
  assign n14825 = ~pi035 & n6259;
  assign n14826 = ~pi106 & n14799;
  assign n14827 = ~n14825 & ~n14826;
  assign n14828 = n14824 & n14827;
  assign n14829 = ~n6238 & n14828;
  assign n14830 = ~n9833 & n14829;
  assign n14831 = ~pi065 & ~n14830;
  assign n14832 = ~n14823 & ~n14831;
  assign n14833 = pi031 & n6200;
  assign n14834 = ~pi035 & n6648;
  assign n14835 = ~n6224 & n6268;
  assign n14836 = ~n6284 & ~n14835;
  assign n14837 = ~n14834 & n14836;
  assign n14838 = ~n14833 & n14837;
  assign n14839 = ~pi106 & ~n14838;
  assign n14840 = ~n6167 & ~n7006;
  assign n14841 = pi106 & ~n14840;
  assign n14842 = ~n14839 & ~n14841;
  assign n14843 = n14832 & n14842;
  assign n14844 = ~pi068 & ~n14843;
  assign n14845 = n14816 & ~n14844;
  assign n14846 = n14776 & n14845;
  assign n14847 = ~pi275 & ~n14660;
  assign n14848 = pi275 & n14660;
  assign n14849 = ~n14847 & ~n14848;
  assign n14850 = ~n14846 & n14849;
  assign n14851 = n14846 & ~n14849;
  assign n14852 = ~n14850 & ~n14851;
  assign n14853 = ~n14768 & ~n14852;
  assign n14854 = n14768 & n14852;
  assign n14855 = ~n14853 & ~n14854;
  assign n14856 = ~pi529 & ~n14855;
  assign n14857 = ~pi275 & pi523;
  assign n14858 = pi275 & ~pi523;
  assign n14859 = ~n14857 & ~n14858;
  assign n14860 = pi529 & ~n14859;
  assign po182 = n14856 | n14860;
  assign n14862 = pi284 & pi414;
  assign n14863 = ~pi284 & ~pi414;
  assign n14864 = ~n14862 & ~n14863;
  assign n14865 = pi529 & n14864;
  assign n14866 = ~n5610 & ~n14406;
  assign n14867 = ~pi005 & n5692;
  assign n14868 = ~n6463 & ~n14867;
  assign n14869 = n14866 & n14868;
  assign n14870 = n10546 & ~n14869;
  assign n14871 = ~n5660 & ~n5882;
  assign n14872 = ~n5632 & n14871;
  assign n14873 = n5863 & ~n14872;
  assign n14874 = ~n5797 & ~n6957;
  assign n14875 = ~pi024 & ~n14874;
  assign n14876 = ~n14873 & ~n14875;
  assign n14877 = pi005 & n5678;
  assign n14878 = ~n5888 & ~n14877;
  assign n14879 = ~n5652 & n14878;
  assign n14880 = n5697 & ~n14879;
  assign n14881 = ~pi005 & n5706;
  assign n14882 = ~n5806 & ~n14881;
  assign n14883 = ~n5825 & n14882;
  assign n14884 = n5736 & ~n14883;
  assign n14885 = ~n14880 & ~n14884;
  assign n14886 = n14876 & n14885;
  assign n14887 = pi024 & n5609;
  assign n14888 = n5836 & n14887;
  assign n14889 = ~n5611 & ~n14888;
  assign n14890 = ~n5887 & n14889;
  assign n14891 = n14886 & n14890;
  assign n14892 = ~n14870 & n14891;
  assign n14893 = pi091 & n5798;
  assign n14894 = ~pi005 & n5637;
  assign n14895 = ~n5655 & ~n6965;
  assign n14896 = ~n5637 & ~n5761;
  assign n14897 = n14895 & n14896;
  assign n14898 = ~pi091 & ~n14897;
  assign n14899 = ~n5665 & ~n6510;
  assign n14900 = ~n5683 & n14899;
  assign n14901 = n5697 & ~n14900;
  assign n14902 = ~n5752 & ~n5856;
  assign n14903 = pi024 & ~n14902;
  assign n14904 = ~n14901 & ~n14903;
  assign n14905 = ~n5652 & n14904;
  assign n14906 = ~n14898 & n14905;
  assign n14907 = ~n14894 & n14906;
  assign n14908 = ~n14893 & n14907;
  assign n14909 = ~pi091 & n5818;
  assign n14910 = n5612 & n5796;
  assign n14911 = ~pi005 & n5850;
  assign n14912 = ~n14910 & ~n14911;
  assign n14913 = ~n14909 & n14912;
  assign n14914 = ~n5761 & ~n5819;
  assign n14915 = n14913 & n14914;
  assign n14916 = ~pi024 & ~n14915;
  assign n14917 = n14908 & ~n14916;
  assign n14918 = pi018 & ~n14917;
  assign n14919 = n14892 & ~n14918;
  assign n14920 = ~pi005 & ~n5653;
  assign n14921 = pi005 & ~n5665;
  assign n14922 = ~n14920 & ~n14921;
  assign n14923 = ~n6922 & ~n14922;
  assign n14924 = ~pi091 & ~n14923;
  assign n14925 = ~n5751 & ~n6516;
  assign n14926 = ~n14924 & n14925;
  assign n14927 = ~n5739 & n14926;
  assign n14928 = pi024 & ~n14927;
  assign n14929 = ~n5617 & ~n5745;
  assign n14930 = n5697 & ~n14929;
  assign n14931 = ~n5806 & ~n14930;
  assign n14932 = ~n6989 & n14931;
  assign n14933 = ~n14928 & n14932;
  assign n14934 = pi091 & n5774;
  assign n14935 = ~n6473 & ~n14934;
  assign n14936 = ~pi024 & ~n14935;
  assign n14937 = n14933 & ~n14936;
  assign n14938 = ~n5786 & ~n6458;
  assign n14939 = ~pi091 & ~n14938;
  assign n14940 = ~pi005 & n6939;
  assign n14941 = ~n6949 & ~n14940;
  assign n14942 = pi091 & ~n14941;
  assign n14943 = ~n14939 & ~n14942;
  assign n14944 = ~n6475 & ~n14451;
  assign n14945 = ~pi091 & ~n14944;
  assign n14946 = ~n6458 & ~n14945;
  assign n14947 = ~n5891 & n14946;
  assign n14948 = ~pi024 & ~n14947;
  assign n14949 = n14943 & ~n14948;
  assign n14950 = n14937 & n14949;
  assign n14951 = ~pi018 & ~n14950;
  assign n14952 = n14919 & ~n14951;
  assign n14953 = ~n7192 & n14952;
  assign n14954 = n7192 & ~n14952;
  assign n14955 = ~n14953 & ~n14954;
  assign n14956 = n5484 & ~n7102;
  assign n14957 = ~n5484 & n7102;
  assign n14958 = ~n14956 & ~n14957;
  assign n14959 = ~n14955 & n14958;
  assign n14960 = n14955 & ~n14958;
  assign n14961 = ~n14959 & ~n14960;
  assign n14962 = n9897 & ~n10760;
  assign n14963 = ~n9897 & n10760;
  assign n14964 = ~n14962 & ~n14963;
  assign n14965 = ~pi284 & ~n10853;
  assign n14966 = pi284 & n10853;
  assign n14967 = ~n14965 & ~n14966;
  assign n14968 = n14964 & n14967;
  assign n14969 = ~n14964 & ~n14967;
  assign n14970 = ~n14968 & ~n14969;
  assign n14971 = ~n14961 & n14970;
  assign n14972 = n14961 & ~n14970;
  assign n14973 = ~n14971 & ~n14972;
  assign n14974 = ~pi529 & n14973;
  assign po183 = n14865 | n14974;
  assign n14976 = ~pi321 & pi494;
  assign n14977 = pi321 & ~pi494;
  assign n14978 = ~n14976 & ~n14977;
  assign n14979 = pi529 & ~n14978;
  assign n14980 = n6163 & ~n10561;
  assign n14981 = ~n6163 & n10561;
  assign n14982 = ~n14980 & ~n14981;
  assign n14983 = n5898 & ~n14982;
  assign n14984 = ~n5898 & n14982;
  assign n14985 = ~n14983 & ~n14984;
  assign n14986 = pi321 & n6906;
  assign n14987 = ~pi321 & ~n6906;
  assign n14988 = ~n14986 & ~n14987;
  assign n14989 = n6328 & ~n6783;
  assign n14990 = ~n6328 & n6783;
  assign n14991 = ~n14989 & ~n14990;
  assign n14992 = n14988 & n14991;
  assign n14993 = ~n14988 & ~n14991;
  assign n14994 = ~n14992 & ~n14993;
  assign n14995 = ~n14985 & n14994;
  assign n14996 = n14985 & ~n14994;
  assign n14997 = ~n14995 & ~n14996;
  assign n14998 = ~pi529 & n14997;
  assign po184 = n14979 | n14998;
  assign n15000 = n9674 & ~n14846;
  assign n15001 = ~n9674 & n14846;
  assign n15002 = ~n15000 & ~n15001;
  assign n15003 = ~pi233 & ~n6906;
  assign n15004 = pi233 & n6906;
  assign n15005 = ~n15003 & ~n15004;
  assign n15006 = n14660 & n15005;
  assign n15007 = ~n14660 & ~n15005;
  assign n15008 = ~n15006 & ~n15007;
  assign n15009 = ~n15002 & ~n15008;
  assign n15010 = n15002 & n15008;
  assign n15011 = ~n15009 & ~n15010;
  assign n15012 = ~pi529 & ~n15011;
  assign n15013 = ~pi233 & pi477;
  assign n15014 = pi233 & ~pi477;
  assign n15015 = ~n15013 & ~n15014;
  assign n15016 = pi529 & ~n15015;
  assign po185 = n15012 | n15016;
  assign n15018 = n9674 & ~n14485;
  assign n15019 = ~n9674 & n14485;
  assign n15020 = ~n15018 & ~n15019;
  assign n15021 = n9897 & ~n14660;
  assign n15022 = ~n9897 & n14660;
  assign n15023 = ~n15021 & ~n15022;
  assign n15024 = ~pi342 & n15023;
  assign n15025 = pi342 & ~n15023;
  assign n15026 = ~n15024 & ~n15025;
  assign n15027 = ~n15020 & ~n15026;
  assign n15028 = n15020 & n15026;
  assign n15029 = ~n15027 & ~n15028;
  assign n15030 = ~pi529 & ~n15029;
  assign n15031 = ~pi342 & pi467;
  assign n15032 = pi342 & ~pi467;
  assign n15033 = ~n15031 & ~n15032;
  assign n15034 = pi529 & ~n15033;
  assign po186 = n15030 | n15034;
  assign n15036 = ~pi147 & pi463;
  assign n15037 = pi147 & ~pi463;
  assign n15038 = ~n15036 & ~n15037;
  assign n15039 = pi529 & ~n15038;
  assign n15040 = ~pi147 & ~n14660;
  assign n15041 = pi147 & n14660;
  assign n15042 = ~n15040 & ~n15041;
  assign n15043 = ~n14399 & n14846;
  assign n15044 = n14399 & ~n14846;
  assign n15045 = ~n15043 & ~n15044;
  assign n15046 = ~n15042 & n15045;
  assign n15047 = n15042 & ~n15045;
  assign n15048 = ~n15046 & ~n15047;
  assign n15049 = ~n5613 & n14925;
  assign n15050 = ~pi091 & ~n15049;
  assign n15051 = pi091 & n5825;
  assign n15052 = ~n6498 & ~n15051;
  assign n15053 = ~n5812 & n15052;
  assign n15054 = ~n15050 & n15053;
  assign n15055 = ~n5751 & ~n5825;
  assign n15056 = ~pi091 & n5794;
  assign n15057 = ~n5721 & ~n6911;
  assign n15058 = pi091 & ~n15057;
  assign n15059 = ~n15056 & ~n15058;
  assign n15060 = n15055 & n15059;
  assign n15061 = ~n5682 & n15060;
  assign n15062 = ~pi024 & ~n15061;
  assign n15063 = n15054 & ~n15062;
  assign n15064 = ~n5786 & ~n5882;
  assign n15065 = ~n6957 & n15064;
  assign n15066 = ~n6943 & n15065;
  assign n15067 = pi024 & ~n15066;
  assign n15068 = pi005 & pi084;
  assign n15069 = ~pi004 & n15068;
  assign n15070 = ~n14440 & ~n15069;
  assign n15071 = ~n6922 & n15070;
  assign n15072 = n10546 & ~n15071;
  assign n15073 = ~n5884 & ~n15072;
  assign n15074 = ~n15067 & n15073;
  assign n15075 = n15063 & n15074;
  assign n15076 = pi018 & ~n15075;
  assign n15077 = ~pi091 & n5773;
  assign n15078 = pi005 & n5610;
  assign n15079 = n5622 & n5663;
  assign n15080 = ~n15078 & ~n15079;
  assign n15081 = ~n15077 & n15080;
  assign n15082 = pi024 & ~n15081;
  assign n15083 = ~n5715 & ~n5818;
  assign n15084 = ~pi005 & n5872;
  assign n15085 = n15083 & ~n15084;
  assign n15086 = ~pi091 & ~n15085;
  assign n15087 = pi005 & n5745;
  assign n15088 = ~n5798 & ~n15087;
  assign n15089 = ~n5622 & ~n10519;
  assign n15090 = pi091 & ~n15089;
  assign n15091 = n15088 & ~n15090;
  assign n15092 = ~n15086 & n15091;
  assign n15093 = ~n5739 & ~n5850;
  assign n15094 = ~n5732 & n15093;
  assign n15095 = n15092 & n15094;
  assign n15096 = pi024 & ~n15095;
  assign n15097 = n5607 & n6922;
  assign n15098 = ~n14479 & ~n15097;
  assign n15099 = ~pi024 & ~n15098;
  assign n15100 = n5706 & n5719;
  assign n15101 = ~n5848 & ~n15100;
  assign n15102 = ~pi024 & ~n15101;
  assign n15103 = ~n15099 & ~n15102;
  assign n15104 = ~n6485 & ~n6976;
  assign n15105 = pi091 & ~n15104;
  assign n15106 = pi005 & n5831;
  assign n15107 = ~n15087 & ~n15106;
  assign n15108 = pi091 & ~n15107;
  assign n15109 = ~n15105 & ~n15108;
  assign n15110 = ~n5610 & ~n14441;
  assign n15111 = ~n15077 & n15110;
  assign n15112 = ~n14443 & n15111;
  assign n15113 = n15109 & n15112;
  assign n15114 = n15103 & n15113;
  assign n15115 = ~n15096 & n15114;
  assign n15116 = ~pi018 & ~n15115;
  assign n15117 = n5607 & n5714;
  assign n15118 = ~pi005 & n5631;
  assign n15119 = ~n5623 & ~n15118;
  assign n15120 = ~n5651 & n15119;
  assign n15121 = ~pi091 & ~n15120;
  assign n15122 = ~n15117 & ~n15121;
  assign n15123 = ~n5806 & n15122;
  assign n15124 = n5719 & ~n5816;
  assign n15125 = ~n5825 & ~n15124;
  assign n15126 = pi091 & ~n15125;
  assign n15127 = n15123 & ~n15126;
  assign n15128 = ~pi024 & ~n15127;
  assign n15129 = ~n15116 & ~n15128;
  assign n15130 = ~n15082 & n15129;
  assign n15131 = ~n15076 & n15130;
  assign n15132 = ~pi091 & n5798;
  assign n15133 = ~n6989 & ~n15132;
  assign n15134 = ~n6522 & n15133;
  assign n15135 = n15131 & n15134;
  assign n15136 = n14762 & n15135;
  assign n15137 = ~n14762 & ~n15135;
  assign n15138 = ~n15136 & ~n15137;
  assign n15139 = ~n15048 & ~n15138;
  assign n15140 = n15048 & n15138;
  assign n15141 = ~n15139 & ~n15140;
  assign n15142 = ~pi529 & ~n15141;
  assign po187 = n15039 | n15142;
  assign n15144 = ~pi234 & pi428;
  assign n15145 = pi234 & ~pi428;
  assign n15146 = ~n15144 & ~n15145;
  assign n15147 = pi529 & ~n15146;
  assign n15148 = ~pi234 & ~n9668;
  assign n15149 = pi234 & n9668;
  assign n15150 = ~n15148 & ~n15149;
  assign n15151 = ~n6906 & n9897;
  assign n15152 = n6906 & ~n9897;
  assign n15153 = ~n15151 & ~n15152;
  assign n15154 = n7001 & n7192;
  assign n15155 = ~n7001 & ~n7192;
  assign n15156 = ~n15154 & ~n15155;
  assign n15157 = n15153 & n15156;
  assign n15158 = ~n15153 & ~n15156;
  assign n15159 = ~n15157 & ~n15158;
  assign n15160 = n15150 & n15159;
  assign n15161 = ~n15150 & ~n15159;
  assign n15162 = ~n15160 & ~n15161;
  assign n15163 = ~pi529 & n15162;
  assign po188 = n15147 | n15163;
  assign n15165 = pi140 & pi423;
  assign n15166 = ~pi140 & ~pi423;
  assign n15167 = ~n15165 & ~n15166;
  assign n15168 = pi529 & ~n15167;
  assign n15169 = ~n10001 & n10961;
  assign n15170 = n10001 & ~n10961;
  assign n15171 = ~n15169 & ~n15170;
  assign n15172 = pi140 & ~n10453;
  assign n15173 = ~pi140 & n10453;
  assign n15174 = ~n15172 & ~n15173;
  assign n15175 = ~n15171 & n15174;
  assign n15176 = n15171 & ~n15174;
  assign n15177 = ~n15175 & ~n15176;
  assign n15178 = n2081 & n15177;
  assign n15179 = ~n2081 & ~n15177;
  assign n15180 = ~n15178 & ~n15179;
  assign n15181 = ~pi529 & n15180;
  assign po189 = n15168 | n15181;
  assign n15183 = ~n10213 & n10247;
  assign n15184 = n10261 & n15183;
  assign n15185 = ~n10217 & n15184;
  assign n15186 = pi001 & n7848;
  assign n15187 = ~n7373 & ~n15186;
  assign n15188 = ~pi013 & n7383;
  assign n15189 = ~n2911 & ~n15188;
  assign n15190 = pi114 & ~n15189;
  assign n15191 = ~pi007 & ~pi114;
  assign n15192 = ~pi054 & n15191;
  assign n15193 = n1764 & n15192;
  assign n15194 = ~n1848 & ~n15193;
  assign n15195 = ~n15190 & n15194;
  assign n15196 = pi001 & ~n15195;
  assign n15197 = ~n1818 & ~n2907;
  assign n15198 = pi013 & pi098;
  assign n15199 = pi007 & n15198;
  assign n15200 = ~pi114 & n15199;
  assign n15201 = ~pi013 & n1867;
  assign n15202 = ~n15200 & ~n15201;
  assign n15203 = ~n1759 & n15202;
  assign n15204 = ~n10989 & n15203;
  assign n15205 = n15197 & n15204;
  assign n15206 = ~pi001 & ~n15205;
  assign n15207 = ~n15196 & ~n15206;
  assign n15208 = ~n1759 & ~n2959;
  assign n15209 = pi114 & ~n15208;
  assign n15210 = ~pi013 & n2870;
  assign n15211 = pi007 & n2969;
  assign n15212 = ~n15210 & ~n15211;
  assign n15213 = ~n1821 & n2945;
  assign n15214 = ~n1890 & ~n15213;
  assign n15215 = n15212 & n15214;
  assign n15216 = ~pi114 & ~n15215;
  assign n15217 = ~n15209 & ~n15216;
  assign n15218 = n15207 & n15217;
  assign n15219 = ~pi029 & ~n15218;
  assign n15220 = n15187 & ~n15219;
  assign n15221 = ~n2861 & ~n10989;
  assign n15222 = ~pi114 & ~n15221;
  assign n15223 = ~n1778 & ~n7832;
  assign n15224 = ~n10055 & ~n10056;
  assign n15225 = n15223 & n15224;
  assign n15226 = ~pi001 & ~n15225;
  assign n15227 = ~n1862 & ~n15199;
  assign n15228 = n2914 & ~n15227;
  assign n15229 = ~n15226 & ~n15228;
  assign n15230 = ~n2837 & ~n2974;
  assign n15231 = pi001 & ~n15230;
  assign n15232 = ~n1771 & ~n7344;
  assign n15233 = ~n11037 & n15232;
  assign n15234 = n2886 & ~n15233;
  assign n15235 = ~n15231 & ~n15234;
  assign n15236 = ~n1772 & ~n2828;
  assign n15237 = ~n7378 & n15236;
  assign n15238 = pi114 & ~n15237;
  assign n15239 = pi001 & n1791;
  assign n15240 = pi007 & ~pi054;
  assign n15241 = ~n2869 & ~n15240;
  assign n15242 = n15239 & ~n15241;
  assign n15243 = ~n15238 & ~n15242;
  assign n15244 = n15235 & n15243;
  assign n15245 = ~n3013 & n15244;
  assign n15246 = n15229 & n15245;
  assign n15247 = ~n15222 & n15246;
  assign n15248 = pi029 & ~n15247;
  assign n15249 = pi114 & n1795;
  assign n15250 = ~n1778 & ~n2845;
  assign n15251 = ~n2980 & n15250;
  assign n15252 = ~pi114 & ~n15251;
  assign n15253 = ~n3032 & ~n7381;
  assign n15254 = ~n7317 & n15253;
  assign n15255 = ~n15252 & n15254;
  assign n15256 = ~n15249 & n15255;
  assign n15257 = ~pi001 & ~n15256;
  assign n15258 = pi114 & n7362;
  assign n15259 = ~n15257 & ~n15258;
  assign n15260 = ~n1827 & ~n10079;
  assign n15261 = pi013 & n7344;
  assign n15262 = ~n7332 & ~n15261;
  assign n15263 = ~n1766 & n15262;
  assign n15264 = n2886 & ~n15263;
  assign n15265 = n15260 & ~n15264;
  assign n15266 = n15259 & n15265;
  assign n15267 = ~n15248 & n15266;
  assign n15268 = n15220 & n15267;
  assign n15269 = ~n15185 & n15268;
  assign n15270 = n15185 & ~n15268;
  assign n15271 = ~n15269 & ~n15270;
  assign n15272 = n10094 & ~n15271;
  assign n15273 = ~n10094 & n15271;
  assign n15274 = ~n15272 & ~n15273;
  assign n15275 = ~n10348 & n10453;
  assign n15276 = n10348 & ~n10453;
  assign n15277 = ~n15275 & ~n15276;
  assign n15278 = pi169 & n15277;
  assign n15279 = ~pi169 & ~n15277;
  assign n15280 = ~n15278 & ~n15279;
  assign n15281 = ~n15274 & n15280;
  assign n15282 = n15274 & ~n15280;
  assign n15283 = ~n15281 & ~n15282;
  assign n15284 = ~pi529 & ~n15283;
  assign n15285 = pi169 & pi525;
  assign n15286 = ~pi169 & ~pi525;
  assign n15287 = ~n15285 & ~n15286;
  assign n15288 = pi529 & n15287;
  assign po190 = n15284 | n15288;
  assign n15290 = ~pi168 & pi411;
  assign n15291 = pi168 & ~pi411;
  assign n15292 = ~n15290 & ~n15291;
  assign n15293 = pi529 & ~n15292;
  assign n15294 = ~pi168 & ~n10182;
  assign n15295 = pi168 & n10182;
  assign n15296 = ~n15294 & ~n15295;
  assign n15297 = ~n10348 & n15296;
  assign n15298 = n10348 & ~n15296;
  assign n15299 = ~n15297 & ~n15298;
  assign n15300 = n10001 & ~n15268;
  assign n15301 = ~n10001 & n15268;
  assign n15302 = ~n15300 & ~n15301;
  assign n15303 = n10961 & n15302;
  assign n15304 = ~n10961 & ~n15302;
  assign n15305 = ~n15303 & ~n15304;
  assign n15306 = ~n15299 & ~n15305;
  assign n15307 = n15299 & n15305;
  assign n15308 = ~n15306 & ~n15307;
  assign n15309 = ~pi529 & ~n15308;
  assign po191 = n15293 | n15309;
  assign n15311 = ~pi152 & pi421;
  assign n15312 = pi152 & ~pi421;
  assign n15313 = ~n15311 & ~n15312;
  assign n15314 = pi529 & ~n15313;
  assign n15315 = ~n10961 & n15271;
  assign n15316 = n10961 & ~n15271;
  assign n15317 = ~n15315 & ~n15316;
  assign n15318 = ~pi152 & ~n10182;
  assign n15319 = pi152 & n10182;
  assign n15320 = ~n15318 & ~n15319;
  assign n15321 = ~n10453 & ~n15320;
  assign n15322 = n10453 & n15320;
  assign n15323 = ~n15321 & ~n15322;
  assign n15324 = ~n15317 & ~n15323;
  assign n15325 = n15317 & n15323;
  assign n15326 = ~n15324 & ~n15325;
  assign n15327 = ~pi529 & ~n15326;
  assign po192 = n15314 | n15327;
  assign n15329 = pi174 & pi479;
  assign n15330 = ~pi174 & ~pi479;
  assign n15331 = ~n15329 & ~n15330;
  assign n15332 = pi529 & n15331;
  assign n15333 = ~n2365 & n11307;
  assign n15334 = n2365 & ~n11307;
  assign n15335 = ~n15333 & ~n15334;
  assign n15336 = ~pi174 & ~n2586;
  assign n15337 = pi174 & n2586;
  assign n15338 = ~n15336 & ~n15337;
  assign n15339 = n15335 & ~n15338;
  assign n15340 = ~n15335 & n15338;
  assign n15341 = ~n15339 & ~n15340;
  assign n15342 = n2811 & n11067;
  assign n15343 = ~n2811 & ~n11067;
  assign n15344 = ~n15342 & ~n15343;
  assign n15345 = n11332 & ~n15344;
  assign n15346 = n2811 & ~n11067;
  assign n15347 = ~n2811 & n11067;
  assign n15348 = ~n15346 & ~n15347;
  assign n15349 = ~n11332 & ~n15348;
  assign n15350 = ~n15345 & ~n15349;
  assign n15351 = ~n15341 & n15350;
  assign n15352 = n15341 & ~n15350;
  assign n15353 = ~n15351 & ~n15352;
  assign n15354 = ~pi529 & n15353;
  assign po193 = n15332 | n15354;
  assign n15356 = ~pi220 & pi458;
  assign n15357 = pi220 & ~pi458;
  assign n15358 = ~n15356 & ~n15357;
  assign n15359 = pi529 & ~n15358;
  assign n15360 = n1752 & ~n3238;
  assign n15361 = ~n1752 & n3238;
  assign n15362 = ~n15360 & ~n15361;
  assign n15363 = n1915 & n7299;
  assign n15364 = ~n1915 & ~n7299;
  assign n15365 = ~n15363 & ~n15364;
  assign n15366 = n15362 & n15365;
  assign n15367 = ~n15362 & ~n15365;
  assign n15368 = ~n15366 & ~n15367;
  assign n15369 = n1627 & n7504;
  assign n15370 = ~n1627 & ~n7504;
  assign n15371 = ~n15369 & ~n15370;
  assign n15372 = ~pi220 & ~n2243;
  assign n15373 = pi220 & n2243;
  assign n15374 = ~n15372 & ~n15373;
  assign n15375 = n15371 & n15374;
  assign n15376 = ~n15371 & ~n15374;
  assign n15377 = ~n15375 & ~n15376;
  assign n15378 = n15368 & n15377;
  assign n15379 = ~n15368 & ~n15377;
  assign n15380 = ~n15378 & ~n15379;
  assign n15381 = ~pi529 & n15380;
  assign po194 = n15359 | n15381;
  assign n15383 = ~pi155 & pi476;
  assign n15384 = pi155 & ~pi476;
  assign n15385 = ~n15383 & ~n15384;
  assign n15386 = pi529 & ~n15385;
  assign n15387 = ~pi155 & ~n11307;
  assign n15388 = pi155 & n11307;
  assign n15389 = ~n15387 & ~n15388;
  assign n15390 = n1627 & ~n2365;
  assign n15391 = ~n1627 & n2365;
  assign n15392 = ~n15390 & ~n15391;
  assign n15393 = n3040 & n3141;
  assign n15394 = ~n3040 & ~n3141;
  assign n15395 = ~n15393 & ~n15394;
  assign n15396 = n15392 & n15395;
  assign n15397 = ~n15392 & ~n15395;
  assign n15398 = ~n15396 & ~n15397;
  assign n15399 = n15389 & n15398;
  assign n15400 = ~n15389 & ~n15398;
  assign n15401 = ~n15399 & ~n15400;
  assign n15402 = ~pi529 & n15401;
  assign po195 = n15386 | n15402;
  assign n15404 = ~n4154 & ~n12018;
  assign n15405 = pi059 & ~pi095;
  assign n15406 = ~n3610 & ~n15405;
  assign n15407 = n4049 & ~n15406;
  assign n15408 = ~n3740 & ~n15407;
  assign n15409 = ~n3744 & n15408;
  assign n15410 = ~n3633 & ~n4134;
  assign n15411 = ~n3668 & n15410;
  assign n15412 = pi115 & ~n15411;
  assign n15413 = n15409 & ~n15412;
  assign n15414 = pi026 & ~n15413;
  assign n15415 = pi008 & pi099;
  assign n15416 = pi059 & n15415;
  assign n15417 = ~n3625 & ~n15416;
  assign n15418 = pi115 & ~n15417;
  assign n15419 = n3616 & n4049;
  assign n15420 = ~n3703 & ~n15419;
  assign n15421 = ~n12402 & n15420;
  assign n15422 = ~n12404 & n15421;
  assign n15423 = ~n15418 & n15422;
  assign n15424 = ~pi026 & ~n15423;
  assign n15425 = ~n15414 & ~n15424;
  assign n15426 = ~n3722 & ~n4215;
  assign n15427 = ~pi115 & ~n15426;
  assign n15428 = ~n3603 & ~n4145;
  assign n15429 = ~n3612 & n15428;
  assign n15430 = ~n11677 & n15429;
  assign n15431 = pi115 & ~n15430;
  assign n15432 = ~n15427 & ~n15431;
  assign n15433 = n15425 & n15432;
  assign n15434 = pi030 & ~n15433;
  assign n15435 = pi008 & n3633;
  assign n15436 = ~n3595 & ~n15435;
  assign n15437 = ~n3746 & n15436;
  assign n15438 = n3728 & ~n15437;
  assign n15439 = pi026 & n12446;
  assign n15440 = ~pi008 & n12006;
  assign n15441 = ~n4190 & ~n15440;
  assign n15442 = pi115 & ~n15441;
  assign n15443 = ~pi115 & n3612;
  assign n15444 = ~n4249 & ~n15443;
  assign n15445 = ~n15442 & n15444;
  assign n15446 = pi026 & ~n15445;
  assign n15447 = ~n4187 & ~n11652;
  assign n15448 = ~pi115 & n15416;
  assign n15449 = ~pi008 & n4097;
  assign n15450 = ~n15448 & ~n15449;
  assign n15451 = ~n3632 & n15450;
  assign n15452 = ~n3722 & n15451;
  assign n15453 = n15447 & n15452;
  assign n15454 = ~pi026 & ~n15453;
  assign n15455 = ~n15446 & ~n15454;
  assign n15456 = ~n3632 & ~n4065;
  assign n15457 = pi115 & ~n15456;
  assign n15458 = ~pi008 & n4196;
  assign n15459 = pi059 & n3621;
  assign n15460 = ~n15458 & ~n15459;
  assign n15461 = n4060 & ~n11655;
  assign n15462 = ~n3674 & ~n15461;
  assign n15463 = n15460 & n15462;
  assign n15464 = ~pi115 & ~n15463;
  assign n15465 = ~n15457 & ~n15464;
  assign n15466 = n15455 & n15465;
  assign n15467 = ~pi030 & ~n15466;
  assign n15468 = ~n15439 & ~n15467;
  assign n15469 = ~n15438 & n15468;
  assign n15470 = pi115 & n11689;
  assign n15471 = ~n4122 & ~n12027;
  assign n15472 = ~n3623 & ~n3703;
  assign n15473 = ~n3667 & n15472;
  assign n15474 = ~pi115 & ~n15473;
  assign n15475 = ~n3638 & ~n15474;
  assign n15476 = n15471 & n15475;
  assign n15477 = ~n15470 & n15476;
  assign n15478 = ~pi026 & ~n15477;
  assign n15479 = pi115 & n3673;
  assign n15480 = ~n15478 & ~n15479;
  assign n15481 = ~n12407 & n15480;
  assign n15482 = n15469 & n15481;
  assign n15483 = ~n15434 & n15482;
  assign n15484 = n15404 & n15483;
  assign n15485 = ~n8241 & ~n11507;
  assign n15486 = pi089 & n12271;
  assign n15487 = n15485 & ~n15486;
  assign n15488 = pi028 & n3559;
  assign n15489 = ~n3438 & ~n15488;
  assign n15490 = ~n3460 & n15489;
  assign n15491 = n3476 & ~n15490;
  assign n15492 = n15487 & ~n15491;
  assign n15493 = pi092 & n12189;
  assign n15494 = ~n3496 & ~n3566;
  assign n15495 = ~n3502 & n15494;
  assign n15496 = ~pi092 & ~n15495;
  assign n15497 = ~n8248 & ~n11498;
  assign n15498 = ~n3552 & n15497;
  assign n15499 = ~n15496 & n15498;
  assign n15500 = ~n15493 & n15499;
  assign n15501 = ~pi089 & ~n15500;
  assign n15502 = pi092 & n3510;
  assign n15503 = ~n15501 & ~n15502;
  assign n15504 = ~n12326 & n15503;
  assign n15505 = pi085 & ~pi087;
  assign n15506 = ~n3530 & ~n15505;
  assign n15507 = n8174 & ~n15506;
  assign n15508 = ~n3451 & ~n3458;
  assign n15509 = ~n15507 & n15508;
  assign n15510 = ~n3559 & ~n8254;
  assign n15511 = ~n3504 & n15510;
  assign n15512 = pi092 & ~n15511;
  assign n15513 = n15509 & ~n15512;
  assign n15514 = pi089 & ~n15513;
  assign n15515 = pi028 & pi050;
  assign n15516 = pi085 & n15515;
  assign n15517 = ~n3454 & ~n15516;
  assign n15518 = pi092 & ~n15517;
  assign n15519 = ~n3496 & ~n12708;
  assign n15520 = ~n15518 & n15519;
  assign n15521 = ~n12352 & n15520;
  assign n15522 = ~n12353 & n15521;
  assign n15523 = ~pi089 & ~n15522;
  assign n15524 = ~n15514 & ~n15523;
  assign n15525 = ~n3432 & ~n11500;
  assign n15526 = ~n3442 & n15525;
  assign n15527 = ~n8230 & n15526;
  assign n15528 = pi092 & ~n15527;
  assign n15529 = ~n3483 & ~n11395;
  assign n15530 = ~pi092 & ~n15529;
  assign n15531 = ~n15528 & ~n15530;
  assign n15532 = n15524 & n15531;
  assign n15533 = pi053 & ~n15532;
  assign n15534 = n15504 & ~n15533;
  assign n15535 = ~pi028 & n11489;
  assign n15536 = ~n8236 & ~n15535;
  assign n15537 = pi092 & ~n15536;
  assign n15538 = ~pi092 & n3432;
  assign n15539 = ~n15537 & ~n15538;
  assign n15540 = ~n11420 & n15539;
  assign n15541 = pi089 & ~n15540;
  assign n15542 = ~n3469 & ~n3483;
  assign n15543 = ~pi028 & n8168;
  assign n15544 = ~pi092 & n15516;
  assign n15545 = ~n15543 & ~n15544;
  assign n15546 = n15542 & n15545;
  assign n15547 = ~n12173 & n15546;
  assign n15548 = ~n11370 & n15547;
  assign n15549 = ~pi089 & ~n15548;
  assign n15550 = ~n15541 & ~n15549;
  assign n15551 = pi085 & n3565;
  assign n15552 = ~pi028 & n11384;
  assign n15553 = n8199 & ~n12168;
  assign n15554 = ~n15552 & ~n15553;
  assign n15555 = ~n15551 & n15554;
  assign n15556 = ~n3500 & n15555;
  assign n15557 = ~pi092 & ~n15556;
  assign n15558 = ~n3469 & ~n8204;
  assign n15559 = pi092 & ~n15558;
  assign n15560 = ~n15557 & ~n15559;
  assign n15561 = n15550 & n15560;
  assign n15562 = ~pi053 & ~n15561;
  assign n15563 = n15534 & ~n15562;
  assign n15564 = n15492 & n15563;
  assign n15565 = ~n15484 & n15564;
  assign n15566 = n15484 & ~n15564;
  assign n15567 = ~n15565 & ~n15566;
  assign n15568 = ~pi071 & pi075;
  assign n15569 = ~n3385 & ~n15568;
  assign n15570 = n3366 & ~n15569;
  assign n15571 = ~n3308 & ~n15570;
  assign n15572 = ~n3314 & n15571;
  assign n15573 = ~n3333 & ~n8033;
  assign n15574 = ~n3397 & n15573;
  assign n15575 = pi080 & ~n15574;
  assign n15576 = n15572 & ~n15575;
  assign n15577 = pi073 & ~n15576;
  assign n15578 = pi110 & n3302;
  assign n15579 = ~n3310 & ~n15578;
  assign n15580 = pi080 & ~n15579;
  assign n15581 = ~n12791 & ~n13065;
  assign n15582 = ~n3365 & n15581;
  assign n15583 = ~n13064 & n15582;
  assign n15584 = ~n15580 & n15583;
  assign n15585 = ~pi073 & ~n15584;
  assign n15586 = ~n15577 & ~n15585;
  assign n15587 = ~n3273 & ~n8055;
  assign n15588 = ~pi080 & ~n15587;
  assign n15589 = ~n3295 & ~n11828;
  assign n15590 = ~n3271 & ~n11768;
  assign n15591 = n15589 & n15590;
  assign n15592 = pi080 & ~n15591;
  assign n15593 = ~n15588 & ~n15592;
  assign n15594 = n15586 & n15593;
  assign n15595 = pi015 & ~n15594;
  assign n15596 = ~pi080 & n3271;
  assign n15597 = ~pi079 & n11900;
  assign n15598 = ~n8109 & ~n15597;
  assign n15599 = pi080 & ~n15598;
  assign n15600 = ~n15596 & ~n15599;
  assign n15601 = ~n8082 & n15600;
  assign n15602 = pi073 & ~n15601;
  assign n15603 = ~pi080 & n15578;
  assign n15604 = ~pi079 & n11803;
  assign n15605 = ~n15603 & ~n15604;
  assign n15606 = ~n8106 & ~n11796;
  assign n15607 = ~n3261 & ~n3273;
  assign n15608 = n15606 & n15607;
  assign n15609 = n15605 & n15608;
  assign n15610 = ~pi073 & ~n15609;
  assign n15611 = ~n15602 & ~n15610;
  assign n15612 = ~n3261 & ~n12900;
  assign n15613 = pi080 & ~n15612;
  assign n15614 = ~pi079 & n8025;
  assign n15615 = pi075 & n3325;
  assign n15616 = ~n11786 & n11826;
  assign n15617 = ~n15615 & ~n15616;
  assign n15618 = ~n3392 & n15617;
  assign n15619 = ~n15614 & n15618;
  assign n15620 = ~pi080 & ~n15619;
  assign n15621 = ~n15613 & ~n15620;
  assign n15622 = n15611 & n15621;
  assign n15623 = ~pi015 & ~n15622;
  assign n15624 = pi079 & n3333;
  assign n15625 = ~n3292 & ~n15624;
  assign n15626 = ~n3316 & n15625;
  assign n15627 = n3257 & ~n15626;
  assign n15628 = ~n11785 & ~n13041;
  assign n15629 = ~n11908 & n15628;
  assign n15630 = pi073 & n12828;
  assign n15631 = n15629 & ~n15630;
  assign n15632 = ~n15627 & n15631;
  assign n15633 = pi080 & n11755;
  assign n15634 = ~n3327 & ~n3365;
  assign n15635 = ~n3394 & n15634;
  assign n15636 = ~pi080 & ~n15635;
  assign n15637 = ~n11884 & ~n11920;
  assign n15638 = ~n3338 & n15637;
  assign n15639 = ~n15636 & n15638;
  assign n15640 = ~n15633 & n15639;
  assign n15641 = ~pi073 & ~n15640;
  assign n15642 = pi080 & n3403;
  assign n15643 = ~n15641 & ~n15642;
  assign n15644 = n15632 & n15643;
  assign n15645 = ~n15623 & n15644;
  assign n15646 = ~n15595 & n15645;
  assign n15647 = pi146 & ~n15646;
  assign n15648 = ~pi146 & n15646;
  assign n15649 = ~n15647 & ~n15648;
  assign n15650 = ~n15567 & n15649;
  assign n15651 = n15567 & ~n15649;
  assign n15652 = ~n15650 & ~n15651;
  assign n15653 = n12560 & ~n15652;
  assign n15654 = ~n12560 & n15652;
  assign n15655 = ~n15653 & ~n15654;
  assign n15656 = ~pi529 & ~n15655;
  assign n15657 = pi146 & pi514;
  assign n15658 = ~pi146 & ~pi514;
  assign n15659 = ~n15657 & ~n15658;
  assign n15660 = pi529 & ~n15659;
  assign po196 = n15656 | n15660;
  assign n15662 = ~pi273 & ~n15646;
  assign n15663 = pi273 & n15646;
  assign n15664 = ~n15662 & ~n15663;
  assign n15665 = ~n15564 & n15664;
  assign n15666 = n15564 & ~n15664;
  assign n15667 = ~n15665 & ~n15666;
  assign n15668 = ~n12131 & ~n12507;
  assign n15669 = ~n4018 & n15668;
  assign n15670 = pi067 & n12102;
  assign n15671 = ~n12090 & ~n15670;
  assign n15672 = ~n3797 & n15671;
  assign n15673 = n3865 & ~n15672;
  assign n15674 = n15669 & ~n15673;
  assign n15675 = pi117 & n11573;
  assign n15676 = ~n3890 & ~n3929;
  assign n15677 = ~n3970 & n15676;
  assign n15678 = ~pi117 & ~n15677;
  assign n15679 = ~n4030 & ~n12139;
  assign n15680 = ~n12078 & n15679;
  assign n15681 = ~n15678 & n15680;
  assign n15682 = ~n15675 & n15681;
  assign n15683 = ~pi002 & ~n15682;
  assign n15684 = pi117 & n12117;
  assign n15685 = ~n15683 & ~n15684;
  assign n15686 = pi002 & n12555;
  assign n15687 = ~pi067 & n12141;
  assign n15688 = ~n3777 & ~n15687;
  assign n15689 = pi117 & ~n15688;
  assign n15690 = ~pi117 & n3886;
  assign n15691 = ~n3903 & ~n15690;
  assign n15692 = ~n15689 & n15691;
  assign n15693 = pi002 & ~n15692;
  assign n15694 = ~n3772 & ~n11580;
  assign n15695 = pi067 & pi105;
  assign n15696 = pi032 & n15695;
  assign n15697 = ~pi117 & n15696;
  assign n15698 = ~pi067 & n3982;
  assign n15699 = ~n15697 & ~n15698;
  assign n15700 = ~n3888 & n15699;
  assign n15701 = ~n12581 & n15700;
  assign n15702 = n15694 & n15701;
  assign n15703 = ~pi002 & ~n15702;
  assign n15704 = ~n15693 & ~n15703;
  assign n15705 = ~n3888 & ~n3928;
  assign n15706 = pi117 & ~n15705;
  assign n15707 = ~pi067 & n3834;
  assign n15708 = pi032 & n3795;
  assign n15709 = ~n15707 & ~n15708;
  assign n15710 = n3935 & ~n11582;
  assign n15711 = ~n11630 & ~n15710;
  assign n15712 = n15709 & n15711;
  assign n15713 = ~pi117 & ~n15712;
  assign n15714 = ~n15706 & ~n15713;
  assign n15715 = n15704 & n15714;
  assign n15716 = ~pi036 & ~n15715;
  assign n15717 = ~n15686 & ~n15716;
  assign n15718 = ~n3852 & ~n12581;
  assign n15719 = ~pi117 & ~n15718;
  assign n15720 = ~n12482 & ~n12484;
  assign n15721 = ~pi117 & n11594;
  assign n15722 = ~n3929 & ~n15721;
  assign n15723 = n15720 & n15722;
  assign n15724 = ~pi002 & ~n15723;
  assign n15725 = ~n3805 & ~n15696;
  assign n15726 = n3780 & ~n15725;
  assign n15727 = ~n15724 & ~n15726;
  assign n15728 = ~n3913 & ~n3977;
  assign n15729 = pi002 & ~n15728;
  assign n15730 = ~n3830 & ~n12102;
  assign n15731 = ~n12643 & n15730;
  assign n15732 = n3865 & ~n15731;
  assign n15733 = ~n15729 & ~n15732;
  assign n15734 = ~n3886 & ~n11555;
  assign n15735 = ~n12136 & n15734;
  assign n15736 = pi117 & ~n15735;
  assign n15737 = pi002 & n3873;
  assign n15738 = pi032 & ~pi064;
  assign n15739 = ~n3833 & ~n15738;
  assign n15740 = n15737 & ~n15739;
  assign n15741 = ~n15736 & ~n15740;
  assign n15742 = n15733 & n15741;
  assign n15743 = ~n4009 & n15742;
  assign n15744 = n15727 & n15743;
  assign n15745 = ~n15719 & n15744;
  assign n15746 = pi036 & ~n15745;
  assign n15747 = n15717 & ~n15746;
  assign n15748 = n15685 & n15747;
  assign n15749 = n15674 & n15748;
  assign n15750 = n12462 & ~n15749;
  assign n15751 = ~n12462 & n15749;
  assign n15752 = ~n15750 & ~n15751;
  assign n15753 = n12363 & n15752;
  assign n15754 = ~n12363 & ~n15752;
  assign n15755 = ~n15753 & ~n15754;
  assign n15756 = ~n15667 & ~n15755;
  assign n15757 = n15667 & n15755;
  assign n15758 = ~n15756 & ~n15757;
  assign n15759 = ~pi529 & ~n15758;
  assign n15760 = ~pi273 & pi427;
  assign n15761 = pi273 & ~pi427;
  assign n15762 = ~n15760 & ~n15761;
  assign n15763 = pi529 & ~n15762;
  assign po197 = n15759 | n15763;
  assign n15765 = ~n15484 & n15749;
  assign n15766 = n15484 & ~n15749;
  assign n15767 = ~n15765 & ~n15766;
  assign n15768 = n12557 & ~n15767;
  assign n15769 = ~n12557 & n15767;
  assign n15770 = ~n15768 & ~n15769;
  assign n15771 = n13072 & ~n15564;
  assign n15772 = ~n13072 & n15564;
  assign n15773 = ~n15771 & ~n15772;
  assign n15774 = pi274 & n15773;
  assign n15775 = ~pi274 & ~n15773;
  assign n15776 = ~n15774 & ~n15775;
  assign n15777 = ~n15770 & n15776;
  assign n15778 = n15770 & ~n15776;
  assign n15779 = ~n15777 & ~n15778;
  assign n15780 = ~pi529 & ~n15779;
  assign n15781 = pi274 & pi440;
  assign n15782 = ~pi274 & ~pi440;
  assign n15783 = ~n15781 & ~n15782;
  assign n15784 = pi529 & n15783;
  assign po198 = n15780 | n15784;
  assign n15786 = ~pi144 & pi497;
  assign n15787 = pi144 & ~pi497;
  assign n15788 = ~n15786 & ~n15787;
  assign n15789 = pi529 & ~n15788;
  assign n15790 = n12363 & ~n12462;
  assign n15791 = ~n12363 & n12462;
  assign n15792 = ~n15790 & ~n15791;
  assign n15793 = ~pi144 & ~n13072;
  assign n15794 = pi144 & n13072;
  assign n15795 = ~n15793 & ~n15794;
  assign n15796 = ~n15792 & n15795;
  assign n15797 = n15792 & ~n15795;
  assign n15798 = ~n15796 & ~n15797;
  assign n15799 = n11747 & n15798;
  assign n15800 = ~n11747 & ~n15798;
  assign n15801 = ~n15799 & ~n15800;
  assign n15802 = ~pi529 & n15801;
  assign po199 = n15789 | n15802;
  assign n15804 = pi283 & pi498;
  assign n15805 = ~pi283 & ~pi498;
  assign n15806 = ~n15804 & ~n15805;
  assign n15807 = pi529 & n15806;
  assign n15808 = n3755 & n12661;
  assign n15809 = ~n3755 & ~n12661;
  assign n15810 = ~n15808 & ~n15809;
  assign n15811 = n13099 & ~n15810;
  assign n15812 = n3755 & ~n12661;
  assign n15813 = ~n3755 & n12661;
  assign n15814 = ~n15812 & ~n15813;
  assign n15815 = ~n13099 & ~n15814;
  assign n15816 = ~n15811 & ~n15815;
  assign n15817 = ~pi283 & ~n3421;
  assign n15818 = pi283 & n3421;
  assign n15819 = ~n15817 & ~n15818;
  assign n15820 = ~n8140 & n12964;
  assign n15821 = n8140 & ~n12964;
  assign n15822 = ~n15820 & ~n15821;
  assign n15823 = ~n15819 & n15822;
  assign n15824 = n15819 & ~n15822;
  assign n15825 = ~n15823 & ~n15824;
  assign n15826 = n15816 & n15825;
  assign n15827 = ~pi529 & n15826;
  assign n15828 = ~n15816 & ~n15825;
  assign n15829 = ~pi529 & n15828;
  assign n15830 = ~n15827 & ~n15829;
  assign po200 = n15807 | ~n15830;
  assign n15832 = pi131 & pi524;
  assign n15833 = ~pi131 & ~pi524;
  assign n15834 = ~n15832 & ~n15833;
  assign n15835 = pi529 & ~n15834;
  assign n15836 = n4267 & ~n12768;
  assign n15837 = ~n4267 & n12768;
  assign n15838 = ~n15836 & ~n15837;
  assign n15839 = pi008 & n4196;
  assign n15840 = pi008 & n3610;
  assign n15841 = ~n3672 & ~n15840;
  assign n15842 = ~n4190 & n15841;
  assign n15843 = pi115 & ~n15842;
  assign n15844 = ~n4151 & ~n4249;
  assign n15845 = ~n3638 & n15844;
  assign n15846 = ~pi115 & ~n15845;
  assign n15847 = ~n15419 & ~n15846;
  assign n15848 = ~n15843 & n15847;
  assign n15849 = ~n15839 & n15848;
  assign n15850 = ~n4079 & n15849;
  assign n15851 = ~pi026 & ~n15850;
  assign n15852 = pi115 & n4203;
  assign n15853 = ~pi115 & n3595;
  assign n15854 = ~n11678 & ~n11725;
  assign n15855 = ~n15853 & n15854;
  assign n15856 = ~n15852 & n15855;
  assign n15857 = ~n3721 & ~n4101;
  assign n15858 = ~n11718 & n15857;
  assign n15859 = ~n12372 & n15858;
  assign n15860 = n15856 & n15859;
  assign n15861 = ~pi026 & ~n15860;
  assign n15862 = pi115 & n3594;
  assign n15863 = pi056 & n4086;
  assign n15864 = ~n4196 & ~n15863;
  assign n15865 = ~pi115 & ~n15864;
  assign n15866 = ~n15862 & ~n15865;
  assign n15867 = ~n4139 & n15866;
  assign n15868 = pi026 & ~n15867;
  assign n15869 = ~n15861 & ~n15868;
  assign n15870 = ~n3617 & ~n3667;
  assign n15871 = ~n3601 & n15870;
  assign n15872 = n3609 & ~n15871;
  assign n15873 = ~n3679 & ~n4120;
  assign n15874 = ~n15872 & n15873;
  assign n15875 = ~n4132 & n15874;
  assign n15876 = n15869 & n15875;
  assign n15877 = pi030 & ~n15876;
  assign n15878 = ~pi008 & n4244;
  assign n15879 = ~n3631 & ~n15878;
  assign n15880 = n3728 & ~n15879;
  assign n15881 = ~n3616 & ~n3656;
  assign n15882 = n4121 & ~n15881;
  assign n15883 = pi115 & n15882;
  assign n15884 = ~n12043 & ~n15883;
  assign n15885 = ~pi115 & n3652;
  assign n15886 = n3596 & n4086;
  assign n15887 = ~n3651 & ~n15886;
  assign n15888 = ~pi115 & ~n15887;
  assign n15889 = ~n15885 & ~n15888;
  assign n15890 = ~n3649 & n15889;
  assign n15891 = pi026 & ~n15890;
  assign n15892 = pi115 & n3626;
  assign n15893 = n3735 & n15892;
  assign n15894 = ~n15891 & ~n15893;
  assign n15895 = n15884 & n15894;
  assign n15896 = ~n15880 & n15895;
  assign n15897 = pi059 & n3609;
  assign n15898 = n3630 & n15897;
  assign n15899 = ~n3659 & ~n12006;
  assign n15900 = ~n4091 & n15899;
  assign n15901 = ~pi115 & ~n15900;
  assign n15902 = ~n3623 & ~n15901;
  assign n15903 = ~n3683 & ~n4055;
  assign n15904 = pi115 & ~n15903;
  assign n15905 = n15902 & ~n15904;
  assign n15906 = pi026 & ~n15905;
  assign n15907 = ~n3703 & ~n12446;
  assign n15908 = n3640 & n11709;
  assign n15909 = ~n4190 & ~n15908;
  assign n15910 = ~pi026 & ~n15909;
  assign n15911 = n15907 & ~n15910;
  assign n15912 = ~n15906 & n15911;
  assign n15913 = ~n15898 & n15912;
  assign n15914 = ~pi030 & ~n15913;
  assign n15915 = n15896 & ~n15914;
  assign n15916 = ~n15877 & n15915;
  assign n15917 = ~n15851 & n15916;
  assign n15918 = n12160 & ~n15917;
  assign n15919 = ~n12160 & n15917;
  assign n15920 = ~n15918 & ~n15919;
  assign n15921 = ~n15838 & n15920;
  assign n15922 = n15838 & ~n15920;
  assign n15923 = ~n15921 & ~n15922;
  assign n15924 = pi131 & n11953;
  assign n15925 = ~pi131 & ~n11953;
  assign n15926 = ~n15924 & ~n15925;
  assign n15927 = ~n11548 & n15926;
  assign n15928 = n11548 & ~n15926;
  assign n15929 = ~n15927 & ~n15928;
  assign n15930 = ~n15923 & n15929;
  assign n15931 = n15923 & ~n15929;
  assign n15932 = ~n15930 & ~n15931;
  assign n15933 = ~pi529 & n15932;
  assign po201 = n15835 | n15933;
  assign n15935 = pi135 & pi430;
  assign n15936 = ~pi135 & ~pi430;
  assign n15937 = ~n15935 & ~n15936;
  assign n15938 = pi529 & ~n15937;
  assign n15939 = n4267 & n15917;
  assign n15940 = ~n4267 & ~n15917;
  assign n15941 = ~n15939 & ~n15940;
  assign n15942 = ~pi067 & n3910;
  assign n15943 = ~n3785 & ~n15942;
  assign n15944 = n3865 & ~n15943;
  assign n15945 = n3806 & n3861;
  assign n15946 = pi002 & n15945;
  assign n15947 = ~n15944 & ~n15946;
  assign n15948 = ~pi117 & n12152;
  assign n15949 = n3821 & n3857;
  assign n15950 = ~n3816 & ~n15949;
  assign n15951 = ~pi117 & ~n15950;
  assign n15952 = ~n15948 & ~n15951;
  assign n15953 = ~n11602 & n15952;
  assign n15954 = pi002 & ~n15953;
  assign n15955 = ~n3770 & ~n3811;
  assign n15956 = n4017 & ~n15955;
  assign n15957 = pi117 & n15956;
  assign n15958 = ~n12100 & ~n15957;
  assign n15959 = ~n15954 & n15958;
  assign n15960 = n15947 & n15959;
  assign n15961 = pi067 & n3834;
  assign n15962 = ~n3819 & ~n3903;
  assign n15963 = ~n12078 & n15962;
  assign n15964 = ~pi117 & ~n15963;
  assign n15965 = pi067 & n3833;
  assign n15966 = ~n11600 & ~n15965;
  assign n15967 = ~n3777 & n15966;
  assign n15968 = pi117 & ~n15967;
  assign n15969 = ~n15721 & ~n15968;
  assign n15970 = ~n15964 & n15969;
  assign n15971 = ~n15961 & n15970;
  assign n15972 = ~n3964 & n15971;
  assign n15973 = ~pi002 & ~n15972;
  assign n15974 = ~n4022 & ~n4029;
  assign n15975 = ~n3766 & ~n3882;
  assign n15976 = ~n3970 & n15975;
  assign n15977 = n3861 & ~n15976;
  assign n15978 = n15974 & ~n15977;
  assign n15979 = ~n12649 & n15978;
  assign n15980 = pi117 & n3952;
  assign n15981 = pi061 & ~pi067;
  assign n15982 = pi032 & n15981;
  assign n15983 = ~n3834 & ~n15982;
  assign n15984 = ~pi117 & ~n15983;
  assign n15985 = ~n15980 & ~n15984;
  assign n15986 = ~n4027 & n15985;
  assign n15987 = pi002 & ~n15986;
  assign n15988 = n15979 & ~n15987;
  assign n15989 = pi117 & n3841;
  assign n15990 = ~pi117 & n12090;
  assign n15991 = ~n11614 & ~n15990;
  assign n15992 = ~n11560 & n15991;
  assign n15993 = ~n15989 & n15992;
  assign n15994 = ~n3764 & ~n11594;
  assign n15995 = ~n11637 & n15994;
  assign n15996 = ~n12541 & n15995;
  assign n15997 = n15993 & n15996;
  assign n15998 = ~pi002 & ~n15997;
  assign n15999 = n15988 & ~n15998;
  assign n16000 = pi036 & ~n15999;
  assign n16001 = n3762 & n12130;
  assign n16002 = ~n3777 & ~n16001;
  assign n16003 = ~pi002 & ~n16002;
  assign n16004 = pi032 & n3861;
  assign n16005 = n3784 & n16004;
  assign n16006 = ~n3929 & ~n12555;
  assign n16007 = ~n3954 & ~n12141;
  assign n16008 = ~n3998 & n16007;
  assign n16009 = ~pi117 & ~n16008;
  assign n16010 = ~n3890 & ~n16009;
  assign n16011 = ~n3866 & ~n11631;
  assign n16012 = pi117 & ~n16011;
  assign n16013 = n16010 & ~n16012;
  assign n16014 = pi002 & ~n16013;
  assign n16015 = n16006 & ~n16014;
  assign n16016 = ~n16005 & n16015;
  assign n16017 = ~n16003 & n16016;
  assign n16018 = ~pi036 & ~n16017;
  assign n16019 = ~n16000 & ~n16018;
  assign n16020 = ~n15973 & n16019;
  assign n16021 = n15960 & n16020;
  assign n16022 = ~n3926 & n16021;
  assign n16023 = n3926 & ~n16021;
  assign n16024 = ~n16022 & ~n16023;
  assign n16025 = n15941 & n16024;
  assign n16026 = ~n15941 & ~n16024;
  assign n16027 = ~n16025 & ~n16026;
  assign n16028 = n11545 & ~n12057;
  assign n16029 = ~n11545 & n12057;
  assign n16030 = ~n16028 & ~n16029;
  assign n16031 = pi135 & ~n11953;
  assign n16032 = ~pi135 & n11953;
  assign n16033 = ~n16031 & ~n16032;
  assign n16034 = n16030 & n16033;
  assign n16035 = ~n16030 & ~n16033;
  assign n16036 = ~n16034 & ~n16035;
  assign n16037 = ~n16027 & n16036;
  assign n16038 = n16027 & ~n16036;
  assign n16039 = ~n16037 & ~n16038;
  assign n16040 = ~pi529 & n16039;
  assign po202 = n15938 | n16040;
  assign n16042 = ~pi230 & pi491;
  assign n16043 = pi230 & ~pi491;
  assign n16044 = ~n16042 & ~n16043;
  assign n16045 = pi529 & ~n16044;
  assign n16046 = ~pi230 & ~n12964;
  assign n16047 = pi230 & n12964;
  assign n16048 = ~n16046 & ~n16047;
  assign n16049 = ~n8140 & n11452;
  assign n16050 = n8140 & ~n11452;
  assign n16051 = ~n16049 & ~n16050;
  assign n16052 = n4042 & n4161;
  assign n16053 = ~n4042 & ~n4161;
  assign n16054 = ~n16052 & ~n16053;
  assign n16055 = n16051 & n16054;
  assign n16056 = ~n16051 & ~n16054;
  assign n16057 = ~n16055 & ~n16056;
  assign n16058 = n16048 & n16057;
  assign n16059 = ~n16048 & ~n16057;
  assign n16060 = ~n16058 & ~n16059;
  assign n16061 = ~pi529 & n16060;
  assign po203 = n16045 | n16061;
  assign n16063 = ~pi180 & pi402;
  assign n16064 = pi180 & ~pi402;
  assign n16065 = ~n16063 & ~n16064;
  assign n16066 = pi529 & ~n16065;
  assign n16067 = ~pi180 & ~n8140;
  assign n16068 = pi180 & n8140;
  assign n16069 = ~n16067 & ~n16068;
  assign n16070 = ~n11545 & n12862;
  assign n16071 = n11545 & ~n12862;
  assign n16072 = ~n16070 & ~n16071;
  assign n16073 = ~n16069 & n16072;
  assign n16074 = n16069 & ~n16072;
  assign n16075 = ~n16073 & ~n16074;
  assign n16076 = n12774 & n16024;
  assign n16077 = ~n12774 & ~n16024;
  assign n16078 = ~n16076 & ~n16077;
  assign n16079 = ~n16075 & n16078;
  assign n16080 = n16075 & ~n16078;
  assign n16081 = ~n16079 & ~n16080;
  assign n16082 = ~pi529 & n16081;
  assign po204 = n16066 | n16082;
  assign n16084 = ~pi148 & pi519;
  assign n16085 = pi148 & ~pi519;
  assign n16086 = ~n16084 & ~n16085;
  assign n16087 = pi529 & ~n16086;
  assign n16088 = n9366 & n13902;
  assign n16089 = ~n9366 & ~n13902;
  assign n16090 = ~n16088 & ~n16089;
  assign n16091 = n9455 & n16090;
  assign n16092 = ~n9455 & ~n16090;
  assign n16093 = ~n16091 & ~n16092;
  assign n16094 = ~pi148 & ~n13628;
  assign n16095 = pi148 & n13628;
  assign n16096 = ~n16094 & ~n16095;
  assign n16097 = n13537 & n16096;
  assign n16098 = ~n13537 & ~n16096;
  assign n16099 = ~n16097 & ~n16098;
  assign n16100 = ~n16093 & n16099;
  assign n16101 = n16093 & ~n16099;
  assign n16102 = ~n16100 & ~n16101;
  assign n16103 = ~pi529 & n16102;
  assign po205 = n16087 | n16103;
  assign n16105 = pi167 & pi492;
  assign n16106 = ~pi167 & ~pi492;
  assign n16107 = ~n16105 & ~n16106;
  assign n16108 = pi529 & n16107;
  assign n16109 = n9274 & n13537;
  assign n16110 = ~n9274 & ~n13537;
  assign n16111 = ~n16109 & ~n16110;
  assign n16112 = pi167 & n16111;
  assign n16113 = ~pi167 & ~n16111;
  assign n16114 = ~n16112 & ~n16113;
  assign n16115 = ~n13441 & n13902;
  assign n16116 = n13441 & ~n13902;
  assign n16117 = ~n16115 & ~n16116;
  assign n16118 = n13345 & ~n16117;
  assign n16119 = n13441 & n13902;
  assign n16120 = ~n13441 & ~n13902;
  assign n16121 = ~n16119 & ~n16120;
  assign n16122 = ~n13345 & ~n16121;
  assign n16123 = ~n16118 & ~n16122;
  assign n16124 = ~n16114 & n16123;
  assign n16125 = n16114 & ~n16123;
  assign n16126 = ~n16124 & ~n16125;
  assign n16127 = ~pi529 & n16126;
  assign po206 = n16108 | n16127;
  assign n16129 = pi223 & pi518;
  assign n16130 = ~pi223 & ~pi518;
  assign n16131 = ~n16129 & ~n16130;
  assign n16132 = pi529 & n16131;
  assign n16133 = ~pi223 & ~n13628;
  assign n16134 = pi223 & n13628;
  assign n16135 = ~n16133 & ~n16134;
  assign n16136 = ~n9274 & n16135;
  assign n16137 = n9274 & ~n16135;
  assign n16138 = ~n16136 & ~n16137;
  assign n16139 = ~n9455 & ~n16121;
  assign n16140 = n9455 & ~n16117;
  assign n16141 = ~n16139 & ~n16140;
  assign n16142 = n16138 & n16141;
  assign n16143 = ~n16138 & ~n16141;
  assign n16144 = ~n16142 & ~n16143;
  assign n16145 = ~pi529 & n16144;
  assign po207 = n16132 | n16145;
  assign n16147 = pi376 & pi459;
  assign n16148 = ~pi376 & ~pi459;
  assign n16149 = ~n16147 & ~n16148;
  assign n16150 = pi529 & n16149;
  assign n16151 = pi376 & n8423;
  assign n16152 = ~pi376 & ~n8423;
  assign n16153 = ~n16151 & ~n16152;
  assign n16154 = ~n4620 & n9554;
  assign n16155 = n4620 & ~n9554;
  assign n16156 = ~n16154 & ~n16155;
  assign n16157 = ~n16153 & n16156;
  assign n16158 = n16153 & ~n16156;
  assign n16159 = ~n16157 & ~n16158;
  assign n16160 = ~n5077 & ~n13243;
  assign n16161 = ~n5305 & ~n13247;
  assign n16162 = ~n16160 & ~n16161;
  assign n16163 = n16159 & n16162;
  assign n16164 = ~n16159 & ~n16162;
  assign n16165 = ~n16163 & ~n16164;
  assign n16166 = ~pi529 & n16165;
  assign po208 = n16150 | n16166;
  assign n16168 = ~pi134 & pi417;
  assign n16169 = pi134 & ~pi417;
  assign n16170 = ~n16168 & ~n16169;
  assign n16171 = pi529 & ~n16170;
  assign n16172 = n8945 & n14175;
  assign n16173 = ~n8945 & ~n14175;
  assign n16174 = ~n16172 & ~n16173;
  assign n16175 = ~pi134 & ~n8623;
  assign n16176 = pi134 & n8623;
  assign n16177 = ~n16175 & ~n16176;
  assign n16178 = ~n16174 & n16177;
  assign n16179 = n16174 & ~n16177;
  assign n16180 = ~n16178 & ~n16179;
  assign n16181 = ~n5298 & n14085;
  assign n16182 = n5298 & ~n14085;
  assign n16183 = ~n16181 & ~n16182;
  assign n16184 = ~n5058 & ~n5065;
  assign n16185 = pi120 & n4983;
  assign n16186 = ~pi074 & pi081;
  assign n16187 = pi016 & n16186;
  assign n16188 = ~n4865 & ~n16187;
  assign n16189 = ~pi120 & ~n16188;
  assign n16190 = ~n16185 & ~n16189;
  assign n16191 = ~n5063 & n16190;
  assign n16192 = pi003 & ~n16191;
  assign n16193 = pi120 & n4872;
  assign n16194 = ~pi120 & n9019;
  assign n16195 = ~n13263 & ~n16194;
  assign n16196 = ~n9010 & n16195;
  assign n16197 = ~n16193 & n16196;
  assign n16198 = ~n4839 & ~n13123;
  assign n16199 = ~n9036 & n16198;
  assign n16200 = ~n13875 & n16199;
  assign n16201 = n16197 & n16200;
  assign n16202 = ~pi003 & ~n16201;
  assign n16203 = ~n4816 & ~n4913;
  assign n16204 = ~n5002 & n16203;
  assign n16205 = n4905 & ~n16204;
  assign n16206 = ~n13192 & ~n16205;
  assign n16207 = ~n16202 & n16206;
  assign n16208 = ~n16192 & n16207;
  assign n16209 = n16184 & n16208;
  assign n16210 = pi044 & ~n16209;
  assign n16211 = pi074 & n4865;
  assign n16212 = ~n4803 & ~n4934;
  assign n16213 = ~n9030 & n16212;
  assign n16214 = ~pi120 & ~n16213;
  assign n16215 = pi074 & n4864;
  assign n16216 = ~n13168 & ~n16215;
  assign n16217 = ~n4845 & n16216;
  assign n16218 = pi120 & ~n16217;
  assign n16219 = ~n13745 & ~n16218;
  assign n16220 = ~n16214 & n16219;
  assign n16221 = ~n16211 & n16220;
  assign n16222 = ~n4995 & n16221;
  assign n16223 = ~pi003 & ~n16222;
  assign n16224 = ~n16210 & ~n16223;
  assign n16225 = ~pi074 & n4941;
  assign n16226 = ~n4826 & ~n16225;
  assign n16227 = n4882 & ~n16226;
  assign n16228 = ~n4802 & ~n4846;
  assign n16229 = n5052 & ~n16228;
  assign n16230 = pi120 & n16229;
  assign n16231 = ~n9038 & ~n16230;
  assign n16232 = ~pi120 & n8989;
  assign n16233 = n4805 & n4901;
  assign n16234 = ~n4798 & ~n16233;
  assign n16235 = ~pi120 & ~n16234;
  assign n16236 = ~n16232 & ~n16235;
  assign n16237 = ~n9013 & n16236;
  assign n16238 = pi003 & ~n16237;
  assign n16239 = n4815 & n4905;
  assign n16240 = pi003 & n16239;
  assign n16241 = ~n16238 & ~n16240;
  assign n16242 = n16231 & n16241;
  assign n16243 = ~n16227 & n16242;
  assign n16244 = pi016 & n4905;
  assign n16245 = n4797 & n16244;
  assign n16246 = ~n4985 & ~n8959;
  assign n16247 = ~n5030 & n16246;
  assign n16248 = ~pi120 & ~n16247;
  assign n16249 = ~n4921 & ~n16248;
  assign n16250 = ~n4883 & ~n13177;
  assign n16251 = pi120 & ~n16250;
  assign n16252 = n16249 & ~n16251;
  assign n16253 = pi003 & ~n16252;
  assign n16254 = ~n4975 & ~n13777;
  assign n16255 = n4837 & n8967;
  assign n16256 = ~n4845 & ~n16255;
  assign n16257 = ~pi003 & ~n16256;
  assign n16258 = n16254 & ~n16257;
  assign n16259 = ~n16253 & n16258;
  assign n16260 = ~n16245 & n16259;
  assign n16261 = ~pi044 & ~n16260;
  assign n16262 = n16243 & ~n16261;
  assign n16263 = n16224 & n16262;
  assign n16264 = ~n4957 & n16263;
  assign n16265 = n4957 & ~n16263;
  assign n16266 = ~n16264 & ~n16265;
  assign n16267 = ~n16183 & n16266;
  assign n16268 = n16183 & ~n16266;
  assign n16269 = ~n16267 & ~n16268;
  assign n16270 = ~n16180 & n16269;
  assign n16271 = n16180 & ~n16269;
  assign n16272 = ~n16270 & ~n16271;
  assign n16273 = ~pi529 & n16272;
  assign po209 = n16171 | n16273;
  assign n16275 = ~pi319 & pi500;
  assign n16276 = pi319 & ~pi500;
  assign n16277 = ~n16275 & ~n16276;
  assign n16278 = pi529 & ~n16277;
  assign n16279 = pi319 & n8423;
  assign n16280 = ~pi319 & ~n8423;
  assign n16281 = ~n16279 & ~n16280;
  assign n16282 = n8623 & n9455;
  assign n16283 = ~n8623 & ~n9455;
  assign n16284 = ~n16282 & ~n16283;
  assign n16285 = n16281 & n16284;
  assign n16286 = ~n16281 & ~n16284;
  assign n16287 = ~n16285 & ~n16286;
  assign n16288 = n9181 & ~n13348;
  assign n16289 = ~n9181 & ~n13638;
  assign n16290 = ~n16288 & ~n16289;
  assign n16291 = ~n16287 & n16290;
  assign n16292 = n16287 & ~n16290;
  assign n16293 = ~n16291 & ~n16292;
  assign n16294 = ~pi529 & n16293;
  assign po210 = n16278 | n16294;
  assign n16296 = ~pi356 & pi398;
  assign n16297 = pi356 & ~pi398;
  assign n16298 = ~n16296 & ~n16297;
  assign n16299 = pi529 & ~n16298;
  assign n16300 = ~n5298 & n14175;
  assign n16301 = n5298 & ~n14175;
  assign n16302 = ~n16300 & ~n16301;
  assign n16303 = n8945 & n13345;
  assign n16304 = ~n8945 & ~n13345;
  assign n16305 = ~n16303 & ~n16304;
  assign n16306 = n16302 & n16305;
  assign n16307 = ~n16302 & ~n16305;
  assign n16308 = ~n16306 & ~n16307;
  assign n16309 = n8748 & n9455;
  assign n16310 = ~n8748 & ~n9455;
  assign n16311 = ~n16309 & ~n16310;
  assign n16312 = ~pi356 & ~n9274;
  assign n16313 = pi356 & n9274;
  assign n16314 = ~n16312 & ~n16313;
  assign n16315 = n16311 & n16314;
  assign n16316 = ~n16311 & ~n16314;
  assign n16317 = ~n16315 & ~n16316;
  assign n16318 = n16308 & n16317;
  assign n16319 = ~n16308 & ~n16317;
  assign n16320 = ~n16318 & ~n16319;
  assign n16321 = ~pi529 & n16320;
  assign po211 = n16299 | n16321;
  assign n16323 = pi019 & n4436;
  assign n16324 = ~n4298 & ~n16323;
  assign n16325 = ~n4345 & n16324;
  assign n16326 = n4319 & ~n16325;
  assign n16327 = pi090 & n4290;
  assign n16328 = n4295 & n16327;
  assign n16329 = ~n13586 & ~n16328;
  assign n16330 = ~n8588 & n16329;
  assign n16331 = pi088 & n8487;
  assign n16332 = ~n9216 & ~n16331;
  assign n16333 = n16330 & n16332;
  assign n16334 = ~n16326 & n16333;
  assign n16335 = ~n4337 & ~n4349;
  assign n16336 = ~n8602 & ~n8611;
  assign n16337 = n16335 & n16336;
  assign n16338 = pi090 & ~n16337;
  assign n16339 = ~n4332 & ~n8310;
  assign n16340 = ~pi090 & ~n16339;
  assign n16341 = ~n16338 & ~n16340;
  assign n16342 = pi019 & n9525;
  assign n16343 = ~n4295 & ~n16342;
  assign n16344 = pi090 & ~n16343;
  assign n16345 = ~n4360 & ~n8511;
  assign n16346 = ~n16344 & n16345;
  assign n16347 = ~n13608 & n16346;
  assign n16348 = ~n13607 & n16347;
  assign n16349 = ~pi088 & ~n16348;
  assign n16350 = ~n4436 & ~n8319;
  assign n16351 = ~n4366 & n16350;
  assign n16352 = pi090 & ~n16351;
  assign n16353 = n9499 & ~n16352;
  assign n16354 = ~n4387 & ~n13568;
  assign n16355 = n8345 & ~n16354;
  assign n16356 = n16353 & ~n16355;
  assign n16357 = pi088 & ~n16356;
  assign n16358 = ~n16349 & ~n16357;
  assign n16359 = n16341 & n16358;
  assign n16360 = pi006 & ~n16359;
  assign n16361 = ~pi090 & n4337;
  assign n16362 = ~pi019 & n8492;
  assign n16363 = ~n8379 & ~n16362;
  assign n16364 = pi090 & ~n16363;
  assign n16365 = ~n16361 & ~n16364;
  assign n16366 = ~n8412 & n16365;
  assign n16367 = pi088 & ~n16366;
  assign n16368 = ~n4312 & ~n4332;
  assign n16369 = ~pi019 & n8448;
  assign n16370 = ~pi090 & n16342;
  assign n16371 = ~n16369 & ~n16370;
  assign n16372 = ~n8376 & ~n9214;
  assign n16373 = n16371 & n16372;
  assign n16374 = n16368 & n16373;
  assign n16375 = ~pi088 & ~n16374;
  assign n16376 = ~n16367 & ~n16375;
  assign n16377 = ~n4312 & ~n9534;
  assign n16378 = pi090 & ~n16377;
  assign n16379 = ~pi019 & n8318;
  assign n16380 = pi049 & n4376;
  assign n16381 = n8461 & ~n9217;
  assign n16382 = ~n4371 & ~n16381;
  assign n16383 = ~n16380 & n16382;
  assign n16384 = ~n16379 & n16383;
  assign n16385 = ~pi090 & ~n16384;
  assign n16386 = ~n16378 & ~n16385;
  assign n16387 = n16376 & n16386;
  assign n16388 = ~pi006 & ~n16387;
  assign n16389 = ~n4442 & ~n8569;
  assign n16390 = ~n4360 & ~n4367;
  assign n16391 = ~n4414 & n16390;
  assign n16392 = ~pi090 & ~n16391;
  assign n16393 = pi090 & n9199;
  assign n16394 = ~n8614 & ~n16393;
  assign n16395 = ~n16392 & n16394;
  assign n16396 = n16389 & n16395;
  assign n16397 = ~pi088 & ~n16396;
  assign n16398 = ~n16388 & ~n16397;
  assign n16399 = ~n16360 & n16398;
  assign n16400 = n16334 & n16399;
  assign n16401 = ~pi271 & ~n16400;
  assign n16402 = pi271 & n16400;
  assign n16403 = ~n16401 & ~n16402;
  assign n16404 = ~n13987 & n16403;
  assign n16405 = n13987 & ~n16403;
  assign n16406 = ~n16404 & ~n16405;
  assign n16407 = n13441 & ~n13810;
  assign n16408 = ~n13441 & n13810;
  assign n16409 = ~n16407 & ~n16408;
  assign n16410 = n13537 & n16409;
  assign n16411 = ~n13537 & ~n16409;
  assign n16412 = ~n16410 & ~n16411;
  assign n16413 = ~n16406 & ~n16412;
  assign n16414 = n16406 & n16412;
  assign n16415 = ~n16413 & ~n16414;
  assign n16416 = ~pi529 & ~n16415;
  assign n16417 = ~pi271 & pi437;
  assign n16418 = pi271 & ~pi437;
  assign n16419 = ~n16417 & ~n16418;
  assign n16420 = pi529 & ~n16419;
  assign po212 = n16416 | n16420;
  assign n16422 = ~pi225 & pi464;
  assign n16423 = pi225 & ~pi464;
  assign n16424 = ~n16422 & ~n16423;
  assign n16425 = pi529 & ~n16424;
  assign n16426 = ~pi225 & ~n9554;
  assign n16427 = pi225 & n9554;
  assign n16428 = ~n16426 & ~n16427;
  assign n16429 = n8423 & ~n8748;
  assign n16430 = ~n8423 & n8748;
  assign n16431 = ~n16429 & ~n16430;
  assign n16432 = n5074 & n5192;
  assign n16433 = ~n5074 & ~n5192;
  assign n16434 = ~n16432 & ~n16433;
  assign n16435 = n16431 & n16434;
  assign n16436 = ~n16431 & ~n16434;
  assign n16437 = ~n16435 & ~n16436;
  assign n16438 = n16428 & n16437;
  assign n16439 = ~n16428 & ~n16437;
  assign n16440 = ~n16438 & ~n16439;
  assign n16441 = ~pi529 & n16440;
  assign po213 = n16425 | n16441;
  assign n16443 = ~pi181 & pi429;
  assign n16444 = pi181 & ~pi429;
  assign n16445 = ~n16443 & ~n16444;
  assign n16446 = pi529 & ~n16445;
  assign n16447 = ~pi181 & ~n8423;
  assign n16448 = pi181 & n8423;
  assign n16449 = ~n16447 & ~n16448;
  assign n16450 = n8521 & ~n14175;
  assign n16451 = ~n8521 & n14175;
  assign n16452 = ~n16450 & ~n16451;
  assign n16453 = ~n16449 & n16452;
  assign n16454 = n16449 & ~n16452;
  assign n16455 = ~n16453 & ~n16454;
  assign n16456 = n9057 & n16266;
  assign n16457 = ~n9057 & ~n16266;
  assign n16458 = ~n16456 & ~n16457;
  assign n16459 = ~n16455 & n16458;
  assign n16460 = n16455 & ~n16458;
  assign n16461 = ~n16459 & ~n16460;
  assign n16462 = ~pi529 & n16461;
  assign po214 = n16446 | n16462;
  assign n16464 = ~pi349 & pi507;
  assign n16465 = pi349 & ~pi507;
  assign n16466 = ~n16464 & ~n16465;
  assign n16467 = pi529 & ~n16466;
  assign n16468 = ~n14085 & n16263;
  assign n16469 = n14085 & ~n16263;
  assign n16470 = ~n16468 & ~n16469;
  assign n16471 = n13204 & ~n16470;
  assign n16472 = ~n13204 & ~n16468;
  assign n16473 = ~n16469 & n16472;
  assign n16474 = ~n16471 & ~n16473;
  assign n16475 = ~n4451 & n8848;
  assign n16476 = n4451 & ~n8848;
  assign n16477 = ~n16475 & ~n16476;
  assign n16478 = pi349 & n16477;
  assign n16479 = ~pi349 & ~n16477;
  assign n16480 = ~n16478 & ~n16479;
  assign n16481 = n16474 & n16480;
  assign n16482 = ~n16474 & ~n16480;
  assign n16483 = ~n16481 & ~n16482;
  assign n16484 = ~pi529 & n16483;
  assign po215 = n16467 | n16484;
  assign n16486 = ~pi145 & pi469;
  assign n16487 = pi145 & ~pi469;
  assign n16488 = ~n16486 & ~n16487;
  assign n16489 = pi529 & ~n16488;
  assign n16490 = ~n13723 & n13987;
  assign n16491 = n13723 & ~n13987;
  assign n16492 = ~n16490 & ~n16491;
  assign n16493 = ~pi145 & ~n16400;
  assign n16494 = pi145 & n16400;
  assign n16495 = ~n16493 & ~n16494;
  assign n16496 = ~n16492 & n16495;
  assign n16497 = n16492 & ~n16495;
  assign n16498 = ~n16496 & ~n16497;
  assign n16499 = ~n16117 & n16498;
  assign n16500 = ~n16121 & ~n16498;
  assign n16501 = ~n16499 & ~n16500;
  assign n16502 = ~pi529 & ~n16501;
  assign po216 = n16489 | n16502;
  assign n16504 = ~pi256 & pi462;
  assign n16505 = pi256 & ~pi462;
  assign n16506 = ~n16504 & ~n16505;
  assign n16507 = pi529 & ~n16506;
  assign n16508 = ~pi256 & ~n16400;
  assign n16509 = pi256 & n16400;
  assign n16510 = ~n16508 & ~n16509;
  assign n16511 = n13628 & n16510;
  assign n16512 = ~n13628 & ~n16510;
  assign n16513 = ~n16511 & ~n16512;
  assign n16514 = ~n13537 & n13813;
  assign n16515 = n13537 & ~n13813;
  assign n16516 = ~n16514 & ~n16515;
  assign n16517 = ~n16513 & ~n16516;
  assign n16518 = n16513 & n16516;
  assign n16519 = ~n16517 & ~n16518;
  assign n16520 = ~pi529 & ~n16519;
  assign po217 = n16507 | n16520;
  assign n16522 = ~pi222 & pi493;
  assign n16523 = pi222 & ~pi493;
  assign n16524 = ~n16522 & ~n16523;
  assign n16525 = pi529 & ~n16524;
  assign n16526 = ~pi222 & ~n8521;
  assign n16527 = pi222 & n8521;
  assign n16528 = ~n16526 & ~n16527;
  assign n16529 = ~n4451 & n16528;
  assign n16530 = n4451 & ~n16528;
  assign n16531 = ~n16529 & ~n16530;
  assign n16532 = ~n4620 & n16470;
  assign n16533 = n4620 & ~n16470;
  assign n16534 = ~n16532 & ~n16533;
  assign n16535 = n16531 & n16534;
  assign n16536 = ~n16531 & ~n16534;
  assign n16537 = ~n16535 & ~n16536;
  assign n16538 = ~pi529 & n16537;
  assign po218 = n16525 | n16538;
  assign n16540 = pi129 & pi420;
  assign n16541 = ~pi129 & ~pi420;
  assign n16542 = ~n16540 & ~n16541;
  assign n16543 = pi529 & n16542;
  assign n16544 = n14315 & ~n14762;
  assign n16545 = ~n14315 & n14762;
  assign n16546 = ~n16544 & ~n16545;
  assign n16547 = ~pi129 & ~n14582;
  assign n16548 = pi129 & n14582;
  assign n16549 = ~n16547 & ~n16548;
  assign n16550 = ~n16546 & n16549;
  assign n16551 = n16546 & ~n16549;
  assign n16552 = ~n16550 & ~n16551;
  assign n16553 = n14982 & n16552;
  assign n16554 = ~n14982 & ~n16552;
  assign n16555 = ~n16553 & ~n16554;
  assign n16556 = ~pi529 & n16555;
  assign po219 = n16543 | n16556;
  assign n16558 = ~pi270 & pi451;
  assign n16559 = pi270 & ~pi451;
  assign n16560 = ~n16558 & ~n16559;
  assign n16561 = pi529 & ~n16560;
  assign n16562 = ~n11187 & n14982;
  assign n16563 = n11187 & ~n14982;
  assign n16564 = ~n16562 & ~n16563;
  assign n16565 = ~pi270 & ~n6060;
  assign n16566 = pi270 & n6060;
  assign n16567 = ~n16565 & ~n16566;
  assign n16568 = n6783 & ~n6906;
  assign n16569 = ~n6783 & n6906;
  assign n16570 = ~n16568 & ~n16569;
  assign n16571 = ~n16567 & n16570;
  assign n16572 = n16567 & ~n16570;
  assign n16573 = ~n16571 & ~n16572;
  assign n16574 = n16564 & n16573;
  assign n16575 = ~n16564 & ~n16573;
  assign n16576 = ~n16574 & ~n16575;
  assign n16577 = ~pi529 & n16576;
  assign po220 = n16561 | n16577;
  assign n16579 = pi170 & pi522;
  assign n16580 = ~pi170 & ~pi522;
  assign n16581 = ~n16579 & ~n16580;
  assign n16582 = pi529 & n16581;
  assign n16583 = n6060 & ~n14315;
  assign n16584 = ~n6060 & n14315;
  assign n16585 = ~n16583 & ~n16584;
  assign n16586 = ~pi170 & n16585;
  assign n16587 = pi170 & ~n16585;
  assign n16588 = ~n16586 & ~n16587;
  assign n16589 = n10561 & n15138;
  assign n16590 = ~n10561 & ~n15138;
  assign n16591 = ~n16589 & ~n16590;
  assign n16592 = ~n16588 & n16591;
  assign n16593 = n16588 & ~n16591;
  assign n16594 = ~n16592 & ~n16593;
  assign n16595 = ~pi529 & n16594;
  assign po221 = n16582 | n16595;
  assign n16597 = pi232 & pi471;
  assign n16598 = ~pi232 & ~pi471;
  assign n16599 = ~n16597 & ~n16598;
  assign n16600 = pi529 & n16599;
  assign n16601 = ~pi232 & ~n14582;
  assign n16602 = pi232 & n14582;
  assign n16603 = ~n16601 & ~n16602;
  assign n16604 = ~n6060 & n16603;
  assign n16605 = n6060 & ~n16603;
  assign n16606 = ~n16604 & ~n16605;
  assign n16607 = n6328 & n15138;
  assign n16608 = ~n6328 & ~n15138;
  assign n16609 = ~n16607 & ~n16608;
  assign n16610 = n16606 & n16609;
  assign n16611 = ~n16606 & ~n16609;
  assign n16612 = ~n16610 & ~n16611;
  assign n16613 = ~pi529 & n16612;
  assign po222 = n16600 | n16613;
  assign n16615 = pi372 & pi446;
  assign n16616 = ~pi372 & ~pi446;
  assign n16617 = ~n16615 & ~n16616;
  assign n16618 = pi529 & n16617;
  assign n16619 = ~pi372 & ~n6906;
  assign n16620 = pi372 & n6906;
  assign n16621 = ~n16619 & ~n16620;
  assign n16622 = n9668 & ~n10760;
  assign n16623 = ~n9668 & n10760;
  assign n16624 = ~n16622 & ~n16623;
  assign n16625 = ~n16621 & n16624;
  assign n16626 = n16621 & ~n16624;
  assign n16627 = ~n16625 & ~n16626;
  assign n16628 = n10672 & n14952;
  assign n16629 = ~n10672 & ~n14952;
  assign n16630 = ~n16628 & ~n16629;
  assign n16631 = ~n7004 & ~n16630;
  assign n16632 = ~n7199 & n16630;
  assign n16633 = ~n16631 & ~n16632;
  assign n16634 = n16627 & n16633;
  assign n16635 = ~n16627 & ~n16633;
  assign n16636 = ~n16634 & ~n16635;
  assign n16637 = ~pi529 & n16636;
  assign po223 = n16618 | n16637;
  assign n16639 = pi285 & pi455;
  assign n16640 = ~pi285 & ~pi455;
  assign n16641 = ~n16639 & ~n16640;
  assign n16642 = pi529 & n16641;
  assign n16643 = ~n9900 & ~n16630;
  assign n16644 = n9900 & n16630;
  assign n16645 = ~n16643 & ~n16644;
  assign n16646 = ~pi285 & ~n10853;
  assign n16647 = pi285 & n10853;
  assign n16648 = ~n16646 & ~n16647;
  assign n16649 = ~n6906 & n9668;
  assign n16650 = n6906 & ~n9668;
  assign n16651 = ~n16649 & ~n16650;
  assign n16652 = ~n16648 & n16651;
  assign n16653 = n16648 & ~n16651;
  assign n16654 = ~n16652 & ~n16653;
  assign n16655 = n16645 & n16654;
  assign n16656 = ~n16645 & ~n16654;
  assign n16657 = ~n16655 & ~n16656;
  assign n16658 = ~pi529 & n16657;
  assign po224 = n16642 | n16658;
  assign n16660 = pi352 & pi489;
  assign n16661 = ~pi352 & ~pi489;
  assign n16662 = ~n16660 & ~n16661;
  assign n16663 = pi529 & n16662;
  assign n16664 = ~n6431 & n6533;
  assign n16665 = n6431 & ~n6533;
  assign n16666 = ~n16664 & ~n16665;
  assign n16667 = n14952 & ~n16666;
  assign n16668 = ~n14952 & ~n16664;
  assign n16669 = ~n16665 & n16668;
  assign n16670 = ~n16667 & ~n16669;
  assign n16671 = ~n10853 & n11175;
  assign n16672 = n10853 & ~n11175;
  assign n16673 = ~n16671 & ~n16672;
  assign n16674 = pi352 & n16673;
  assign n16675 = ~pi352 & ~n16673;
  assign n16676 = ~n16674 & ~n16675;
  assign n16677 = n16670 & n16676;
  assign n16678 = ~n16670 & ~n16676;
  assign n16679 = ~n16677 & ~n16678;
  assign n16680 = ~pi529 & n16679;
  assign po225 = n16663 | n16680;
  assign n16682 = ~pi207 & pi419;
  assign n16683 = pi207 & ~pi419;
  assign n16684 = ~n16682 & ~n16683;
  assign n16685 = pi529 & ~n16684;
  assign n16686 = n6431 & ~n11175;
  assign n16687 = ~n6431 & n11175;
  assign n16688 = ~n16686 & ~n16687;
  assign n16689 = ~pi207 & ~n9771;
  assign n16690 = pi207 & n9771;
  assign n16691 = ~n16689 & ~n16690;
  assign n16692 = ~n16688 & n16691;
  assign n16693 = n16688 & ~n16691;
  assign n16694 = ~n16692 & ~n16693;
  assign n16695 = ~n16630 & n16694;
  assign n16696 = n16630 & ~n16694;
  assign n16697 = ~n16695 & ~n16696;
  assign n16698 = ~pi529 & n16697;
  assign po226 = n16685 | n16698;
  assign n16700 = ~pi231 & pi460;
  assign n16701 = pi231 & ~pi460;
  assign n16702 = ~n16700 & ~n16701;
  assign n16703 = pi529 & ~n16702;
  assign n16704 = ~pi231 & ~n9771;
  assign n16705 = pi231 & n9771;
  assign n16706 = ~n16704 & ~n16705;
  assign n16707 = ~n10853 & n16706;
  assign n16708 = n10853 & ~n16706;
  assign n16709 = ~n16707 & ~n16708;
  assign n16710 = ~n10760 & n16666;
  assign n16711 = n10760 & ~n16666;
  assign n16712 = ~n16710 & ~n16711;
  assign n16713 = n16709 & n16712;
  assign n16714 = ~n16709 & ~n16712;
  assign n16715 = ~n16713 & ~n16714;
  assign n16716 = ~pi529 & n16715;
  assign po227 = n16703 | n16716;
  assign n16718 = ~pi354 & ~n6906;
  assign n16719 = pi354 & n6906;
  assign n16720 = ~n16718 & ~n16719;
  assign n16721 = ~n9897 & n16720;
  assign n16722 = n9897 & ~n16720;
  assign n16723 = ~n16721 & ~n16722;
  assign n16724 = ~n5772 & n14399;
  assign n16725 = n5772 & ~n14399;
  assign n16726 = ~n16724 & ~n16725;
  assign n16727 = n14846 & n16726;
  assign n16728 = ~n14846 & ~n16726;
  assign n16729 = ~n16727 & ~n16728;
  assign n16730 = ~n16723 & ~n16729;
  assign n16731 = n16723 & n16729;
  assign n16732 = ~n16730 & ~n16731;
  assign n16733 = ~pi529 & ~n16732;
  assign n16734 = ~pi354 & pi434;
  assign n16735 = pi354 & ~pi434;
  assign n16736 = ~n16734 & ~n16735;
  assign n16737 = pi529 & ~n16736;
  assign po228 = n16733 | n16737;
  assign n16739 = ~n5484 & n9897;
  assign n16740 = n5484 & ~n9897;
  assign n16741 = ~n16739 & ~n16740;
  assign n16742 = ~pi166 & ~n6906;
  assign n16743 = pi166 & n6906;
  assign n16744 = ~n16742 & ~n16743;
  assign n16745 = n16741 & n16744;
  assign n16746 = ~n16741 & ~n16744;
  assign n16747 = ~n16745 & ~n16746;
  assign n16748 = ~n14488 & n16747;
  assign n16749 = ~n14492 & ~n16747;
  assign n16750 = ~n16748 & ~n16749;
  assign n16751 = ~pi529 & ~n16750;
  assign n16752 = ~pi166 & pi508;
  assign n16753 = pi166 & ~pi508;
  assign n16754 = ~n16752 & ~n16753;
  assign n16755 = pi529 & ~n16754;
  assign po229 = n16751 | n16755;
  assign n16757 = ~pi133 & pi456;
  assign n16758 = pi133 & ~pi456;
  assign n16759 = ~n16757 & ~n16758;
  assign n16760 = pi529 & ~n16759;
  assign n16761 = n2078 & n10094;
  assign n16762 = ~n2078 & ~n10094;
  assign n16763 = ~n16761 & ~n16762;
  assign n16764 = n7504 & n16763;
  assign n16765 = ~n7504 & ~n16763;
  assign n16766 = ~n16764 & ~n16765;
  assign n16767 = ~pi133 & ~n10453;
  assign n16768 = pi133 & n10453;
  assign n16769 = ~n16767 & ~n16768;
  assign n16770 = n10961 & n16769;
  assign n16771 = ~n10961 & ~n16769;
  assign n16772 = ~n16770 & ~n16771;
  assign n16773 = ~n16766 & n16772;
  assign n16774 = n16766 & ~n16772;
  assign n16775 = ~n16773 & ~n16774;
  assign n16776 = ~pi529 & n16775;
  assign po230 = n16760 | n16776;
  assign n16778 = pi257 & pi486;
  assign n16779 = ~pi257 & ~pi486;
  assign n16780 = ~n16778 & ~n16779;
  assign n16781 = pi529 & n16780;
  assign n16782 = ~pi257 & ~n2365;
  assign n16783 = pi257 & n2365;
  assign n16784 = ~n16782 & ~n16783;
  assign n16785 = ~n2689 & n11307;
  assign n16786 = n2689 & ~n11307;
  assign n16787 = ~n16785 & ~n16786;
  assign n16788 = ~n16784 & n16787;
  assign n16789 = n16784 & ~n16787;
  assign n16790 = ~n16788 & ~n16789;
  assign n16791 = ~n3043 & ~n15344;
  assign n16792 = ~n3245 & ~n15348;
  assign n16793 = ~n16791 & ~n16792;
  assign n16794 = n16790 & n16793;
  assign n16795 = ~n16790 & ~n16793;
  assign n16796 = ~n16794 & ~n16795;
  assign n16797 = ~pi529 & n16796;
  assign po231 = n16781 | n16797;
  assign n16799 = ~pi156 & pi403;
  assign n16800 = pi156 & ~pi403;
  assign n16801 = ~n16799 & ~n16800;
  assign n16802 = pi529 & ~n16801;
  assign n16803 = ~n10348 & n11313;
  assign n16804 = n10348 & ~n11313;
  assign n16805 = ~n16803 & ~n16804;
  assign n16806 = ~pi156 & ~n2365;
  assign n16807 = pi156 & n2365;
  assign n16808 = ~n16806 & ~n16807;
  assign n16809 = n10182 & n16808;
  assign n16810 = ~n10182 & ~n16808;
  assign n16811 = ~n16809 & ~n16810;
  assign n16812 = ~n16805 & ~n16811;
  assign n16813 = n16805 & n16811;
  assign n16814 = ~n16812 & ~n16813;
  assign n16815 = ~pi529 & ~n16814;
  assign po232 = n16802 | n16815;
  assign n16817 = ~pi165 & pi424;
  assign n16818 = pi165 & ~pi424;
  assign n16819 = ~n16817 & ~n16818;
  assign n16820 = pi529 & ~n16819;
  assign n16821 = ~pi165 & ~n2365;
  assign n16822 = pi165 & n2365;
  assign n16823 = ~n16821 & ~n16822;
  assign n16824 = ~n1627 & n3238;
  assign n16825 = n1627 & ~n3238;
  assign n16826 = ~n16824 & ~n16825;
  assign n16827 = ~n16823 & n16826;
  assign n16828 = n16823 & ~n16826;
  assign n16829 = ~n16827 & ~n16828;
  assign n16830 = n15271 & ~n16829;
  assign n16831 = ~n15271 & n16829;
  assign n16832 = ~n16830 & ~n16831;
  assign n16833 = ~pi529 & ~n16832;
  assign po233 = n16820 | n16833;
  assign n16835 = ~pi219 & ~n2365;
  assign n16836 = pi219 & n2365;
  assign n16837 = ~n16835 & ~n16836;
  assign n16838 = n1627 & n16837;
  assign n16839 = ~n1627 & ~n16837;
  assign n16840 = ~n16838 & ~n16839;
  assign n16841 = ~n2937 & n10264;
  assign n16842 = n2937 & ~n10264;
  assign n16843 = ~n16841 & ~n16842;
  assign n16844 = ~n10348 & n16843;
  assign n16845 = n10348 & ~n16843;
  assign n16846 = ~n16844 & ~n16845;
  assign n16847 = ~n16840 & ~n16846;
  assign n16848 = n16840 & n16846;
  assign n16849 = ~n16847 & ~n16848;
  assign n16850 = ~pi529 & ~n16849;
  assign n16851 = ~pi219 & pi422;
  assign n16852 = pi219 & ~pi422;
  assign n16853 = ~n16851 & ~n16852;
  assign n16854 = pi529 & ~n16853;
  assign po234 = n16850 | n16854;
  assign n16856 = ~n12363 & n15767;
  assign n16857 = n12363 & ~n15767;
  assign n16858 = ~n16856 & ~n16857;
  assign n16859 = ~pi227 & ~n15646;
  assign n16860 = pi227 & n15646;
  assign n16861 = ~n16859 & ~n16860;
  assign n16862 = n13072 & n16861;
  assign n16863 = ~n13072 & ~n16861;
  assign n16864 = ~n16862 & ~n16863;
  assign n16865 = ~n16858 & ~n16864;
  assign n16866 = n16858 & n16864;
  assign n16867 = ~n16865 & ~n16866;
  assign n16868 = ~pi529 & ~n16867;
  assign n16869 = ~pi227 & pi425;
  assign n16870 = pi227 & ~pi425;
  assign n16871 = ~n16869 & ~n16870;
  assign n16872 = pi529 & ~n16871;
  assign po235 = n16868 | n16872;
  assign n16874 = pi149 & pi452;
  assign n16875 = ~pi149 & ~pi452;
  assign n16876 = ~n16874 & ~n16875;
  assign n16877 = pi529 & ~n16876;
  assign n16878 = n11744 & n12557;
  assign n16879 = ~n11744 & ~n12557;
  assign n16880 = ~n16878 & ~n16879;
  assign n16881 = n12252 & n16880;
  assign n16882 = ~n12252 & ~n16880;
  assign n16883 = ~n16881 & ~n16882;
  assign n16884 = pi149 & ~n13072;
  assign n16885 = ~pi149 & n13072;
  assign n16886 = ~n16884 & ~n16885;
  assign n16887 = n12363 & n16886;
  assign n16888 = ~n12363 & ~n16886;
  assign n16889 = ~n16887 & ~n16888;
  assign n16890 = ~n16883 & n16889;
  assign n16891 = n16883 & ~n16889;
  assign n16892 = ~n16890 & ~n16891;
  assign n16893 = ~pi529 & n16892;
  assign po236 = n16877 | n16893;
  assign n16895 = pi373 & pi465;
  assign n16896 = ~pi373 & ~pi465;
  assign n16897 = ~n16895 & ~n16896;
  assign n16898 = pi529 & n16897;
  assign n16899 = ~pi373 & ~n8140;
  assign n16900 = pi373 & n8140;
  assign n16901 = ~n16899 & ~n16900;
  assign n16902 = ~n3591 & n12964;
  assign n16903 = n3591 & ~n12964;
  assign n16904 = ~n16902 & ~n16903;
  assign n16905 = ~n16901 & n16904;
  assign n16906 = n16901 & ~n16904;
  assign n16907 = ~n16905 & ~n16906;
  assign n16908 = ~n4045 & ~n15810;
  assign n16909 = ~n4274 & ~n15814;
  assign n16910 = ~n16908 & ~n16909;
  assign n16911 = n16907 & n16910;
  assign n16912 = ~n16907 & ~n16910;
  assign n16913 = ~n16911 & ~n16912;
  assign n16914 = ~pi529 & n16913;
  assign po237 = n16898 | n16914;
  assign n16916 = ~pi357 & pi473;
  assign n16917 = pi357 & ~pi473;
  assign n16918 = ~n16916 & ~n16917;
  assign n16919 = pi529 & ~n16918;
  assign n16920 = ~n4267 & n11545;
  assign n16921 = n4267 & ~n11545;
  assign n16922 = ~n16920 & ~n16921;
  assign n16923 = n11649 & n12057;
  assign n16924 = ~n11649 & ~n12057;
  assign n16925 = ~n16923 & ~n16924;
  assign n16926 = n16922 & n16925;
  assign n16927 = ~n16922 & ~n16925;
  assign n16928 = ~n16926 & ~n16927;
  assign n16929 = n11452 & n12252;
  assign n16930 = ~n11452 & ~n12252;
  assign n16931 = ~n16929 & ~n16930;
  assign n16932 = ~pi357 & ~n11853;
  assign n16933 = pi357 & n11853;
  assign n16934 = ~n16932 & ~n16933;
  assign n16935 = n16931 & n16934;
  assign n16936 = ~n16931 & ~n16934;
  assign n16937 = ~n16935 & ~n16936;
  assign n16938 = n16928 & n16937;
  assign n16939 = ~n16928 & ~n16937;
  assign n16940 = ~n16938 & ~n16939;
  assign n16941 = ~pi529 & n16940;
  assign po238 = n16919 | n16941;
  assign n16943 = pi350 & pi454;
  assign n16944 = ~pi350 & ~pi454;
  assign n16945 = ~n16943 & ~n16944;
  assign n16946 = pi529 & n16945;
  assign n16947 = ~n15917 & n16021;
  assign n16948 = n15917 & ~n16021;
  assign n16949 = ~n16947 & ~n16948;
  assign n16950 = n12661 & ~n16949;
  assign n16951 = ~n12661 & ~n16947;
  assign n16952 = ~n16948 & n16951;
  assign n16953 = ~n16950 & ~n16952;
  assign n16954 = ~n3421 & n12768;
  assign n16955 = n3421 & ~n12768;
  assign n16956 = ~n16954 & ~n16955;
  assign n16957 = pi350 & n16956;
  assign n16958 = ~pi350 & ~n16956;
  assign n16959 = ~n16957 & ~n16958;
  assign n16960 = n16953 & n16959;
  assign n16961 = ~n16953 & ~n16959;
  assign n16962 = ~n16960 & ~n16961;
  assign n16963 = ~pi529 & n16962;
  assign po239 = n16946 | n16963;
  assign n16965 = pi163 & ~n8140;
  assign n16966 = ~pi163 & n8140;
  assign n16967 = ~n16965 & ~n16966;
  assign n16968 = n4267 & ~n11452;
  assign n16969 = ~n4267 & n11452;
  assign n16970 = ~n16968 & ~n16969;
  assign n16971 = n16967 & n16970;
  assign n16972 = ~n16967 & ~n16970;
  assign n16973 = ~n16971 & ~n16972;
  assign n16974 = n15767 & n16973;
  assign n16975 = ~n15767 & ~n16973;
  assign n16976 = ~n16974 & ~n16975;
  assign n16977 = ~pi529 & ~n16976;
  assign n16978 = pi163 & pi504;
  assign n16979 = ~pi163 & ~pi504;
  assign n16980 = ~n16978 & ~n16979;
  assign n16981 = pi529 & ~n16980;
  assign po240 = n16977 | n16981;
  assign n16983 = ~pi229 & pi474;
  assign n16984 = pi229 & ~pi474;
  assign n16985 = ~n16983 & ~n16984;
  assign n16986 = pi529 & ~n16985;
  assign n16987 = ~pi229 & ~n12862;
  assign n16988 = pi229 & n12862;
  assign n16989 = ~n16987 & ~n16988;
  assign n16990 = n3421 & n16989;
  assign n16991 = ~n3421 & ~n16989;
  assign n16992 = ~n16990 & ~n16991;
  assign n16993 = ~n3591 & n16949;
  assign n16994 = n3591 & ~n16949;
  assign n16995 = ~n16993 & ~n16994;
  assign n16996 = ~n16992 & n16995;
  assign n16997 = n16992 & ~n16995;
  assign n16998 = ~n16996 & ~n16997;
  assign n16999 = ~pi529 & n16998;
  assign po241 = n16986 | n16999;
  assign n17001 = ~pi269 & pi415;
  assign n17002 = pi269 & ~pi415;
  assign n17003 = ~n17001 & ~n17002;
  assign n17004 = pi529 & ~n17003;
  assign n17005 = n8423 & ~n8623;
  assign n17006 = ~n8423 & n8623;
  assign n17007 = ~n17005 & ~n17006;
  assign n17008 = ~pi269 & ~n9274;
  assign n17009 = pi269 & n9274;
  assign n17010 = ~n17008 & ~n17009;
  assign n17011 = ~n17007 & n17010;
  assign n17012 = n17007 & ~n17010;
  assign n17013 = ~n17011 & ~n17012;
  assign n17014 = ~n13348 & n14178;
  assign n17015 = ~n13638 & ~n14178;
  assign n17016 = ~n17014 & ~n17015;
  assign n17017 = ~n17013 & n17016;
  assign n17018 = n17013 & ~n17016;
  assign n17019 = ~n17017 & ~n17018;
  assign n17020 = ~pi529 & n17019;
  assign po242 = n17004 | n17020;
  assign n17022 = ~n13987 & n14196;
  assign n17023 = n13987 & ~n14196;
  assign n17024 = ~n17022 & ~n17023;
  assign n17025 = ~pi224 & ~n8423;
  assign n17026 = pi224 & n8423;
  assign n17027 = ~n17025 & ~n17026;
  assign n17028 = ~n16400 & ~n17027;
  assign n17029 = n16400 & n17027;
  assign n17030 = ~n17028 & ~n17029;
  assign n17031 = ~n17024 & ~n17030;
  assign n17032 = n17024 & n17030;
  assign n17033 = ~n17031 & ~n17032;
  assign n17034 = ~pi529 & ~n17033;
  assign n17035 = ~pi224 & pi399;
  assign n17036 = pi224 & ~pi399;
  assign n17037 = ~n17035 & ~n17036;
  assign n17038 = pi529 & ~n17037;
  assign po243 = n17034 | n17038;
  assign n17040 = ~pi353 & ~n8423;
  assign n17041 = pi353 & n8423;
  assign n17042 = ~n17040 & ~n17041;
  assign n17043 = n8748 & n17042;
  assign n17044 = ~n8748 & ~n17042;
  assign n17045 = ~n17043 & ~n17044;
  assign n17046 = ~n4957 & n13723;
  assign n17047 = n4957 & ~n13723;
  assign n17048 = ~n17046 & ~n17047;
  assign n17049 = ~n13987 & n17048;
  assign n17050 = n13987 & ~n17048;
  assign n17051 = ~n17049 & ~n17050;
  assign n17052 = ~n17045 & ~n17051;
  assign n17053 = n17045 & n17051;
  assign n17054 = ~n17052 & ~n17053;
  assign n17055 = ~pi529 & ~n17054;
  assign n17056 = ~pi353 & pi510;
  assign n17057 = pi353 & ~pi510;
  assign n17058 = ~n17056 & ~n17057;
  assign n17059 = pi529 & ~n17058;
  assign po244 = n17055 | n17059;
  assign n17061 = ~pi370 & pi433;
  assign n17062 = pi370 & ~pi433;
  assign n17063 = ~n17061 & ~n17062;
  assign n17064 = pi529 & ~n17063;
  assign n17065 = ~n13810 & n14196;
  assign n17066 = n13810 & ~n14196;
  assign n17067 = ~n17065 & ~n17066;
  assign n17068 = n8748 & ~n16400;
  assign n17069 = ~n8748 & n16400;
  assign n17070 = ~n17068 & ~n17069;
  assign n17071 = ~pi370 & n17070;
  assign n17072 = pi370 & ~n17070;
  assign n17073 = ~n17071 & ~n17072;
  assign n17074 = ~n17067 & n17073;
  assign n17075 = n17067 & ~n17073;
  assign n17076 = ~n17074 & ~n17075;
  assign n17077 = ~pi529 & n17076;
  assign po245 = n17064 | n17077;
  assign n17079 = ~pi157 & pi521;
  assign n17080 = pi157 & ~pi521;
  assign n17081 = ~n17079 & ~n17080;
  assign n17082 = pi529 & ~n17081;
  assign n17083 = n6163 & n15135;
  assign n17084 = ~n6163 & ~n15135;
  assign n17085 = ~n17083 & ~n17084;
  assign n17086 = n6328 & n17085;
  assign n17087 = ~n6328 & ~n17085;
  assign n17088 = ~n17086 & ~n17087;
  assign n17089 = ~pi157 & ~n14582;
  assign n17090 = pi157 & n14582;
  assign n17091 = ~n17089 & ~n17090;
  assign n17092 = n14315 & n17091;
  assign n17093 = ~n14315 & ~n17091;
  assign n17094 = ~n17092 & ~n17093;
  assign n17095 = ~n17088 & n17094;
  assign n17096 = n17088 & ~n17094;
  assign n17097 = ~n17095 & ~n17096;
  assign n17098 = ~pi529 & n17097;
  assign po246 = n17082 | n17098;
  assign n17100 = ~pi276 & pi413;
  assign n17101 = pi276 & ~pi413;
  assign n17102 = ~n17100 & ~n17101;
  assign n17103 = pi529 & ~n17102;
  assign n17104 = ~n14492 & n15135;
  assign n17105 = ~n14488 & ~n15135;
  assign n17106 = ~n17104 & ~n17105;
  assign n17107 = n14582 & ~n14846;
  assign n17108 = ~n14582 & n14846;
  assign n17109 = ~n17107 & ~n17108;
  assign n17110 = pi276 & n17109;
  assign n17111 = ~pi276 & ~n17109;
  assign n17112 = ~n17110 & ~n17111;
  assign n17113 = n17106 & n17112;
  assign n17114 = ~n17106 & ~n17112;
  assign n17115 = ~n17113 & ~n17114;
  assign n17116 = ~pi529 & n17115;
  assign po247 = n17103 | n17116;
  assign n17118 = pi218 & pi461;
  assign n17119 = ~pi218 & ~pi461;
  assign n17120 = ~n17118 & ~n17119;
  assign n17121 = pi529 & n17120;
  assign n17122 = ~n7691 & n7888;
  assign n17123 = n7691 & ~n7888;
  assign n17124 = ~n17122 & ~n17123;
  assign n17125 = n11067 & ~n17124;
  assign n17126 = ~n11067 & ~n17122;
  assign n17127 = ~n17123 & n17126;
  assign n17128 = ~n17125 & ~n17127;
  assign n17129 = ~n2586 & n7605;
  assign n17130 = n2586 & ~n7605;
  assign n17131 = ~n17129 & ~n17130;
  assign n17132 = pi218 & n17131;
  assign n17133 = ~pi218 & ~n17131;
  assign n17134 = ~n17132 & ~n17133;
  assign n17135 = n17128 & n17134;
  assign n17136 = ~n17128 & ~n17134;
  assign n17137 = ~n17135 & ~n17136;
  assign n17138 = ~pi529 & n17137;
  assign po248 = n17121 | n17138;
  assign n17140 = ~pi209 & pi435;
  assign n17141 = pi209 & ~pi435;
  assign n17142 = ~n17140 & ~n17141;
  assign n17143 = pi529 & ~n17142;
  assign n17144 = ~pi209 & ~n7798;
  assign n17145 = pi209 & n7798;
  assign n17146 = ~n17144 & ~n17145;
  assign n17147 = ~n7605 & n7691;
  assign n17148 = n7605 & ~n7691;
  assign n17149 = ~n17147 & ~n17148;
  assign n17150 = n17146 & ~n17149;
  assign n17151 = ~n17146 & n17149;
  assign n17152 = ~n17150 & ~n17151;
  assign n17153 = ~n15344 & n17152;
  assign n17154 = ~n15348 & ~n17152;
  assign n17155 = ~n17153 & ~n17154;
  assign n17156 = ~pi529 & n17155;
  assign po249 = n17143 | n17156;
  assign n17158 = ~pi217 & pi499;
  assign n17159 = pi217 & ~pi499;
  assign n17160 = ~n17158 & ~n17159;
  assign n17161 = pi529 & ~n17160;
  assign n17162 = n2811 & n7888;
  assign n17163 = ~n2811 & ~n7888;
  assign n17164 = ~n17162 & ~n17163;
  assign n17165 = n2689 & n17164;
  assign n17166 = ~n2689 & ~n17164;
  assign n17167 = ~n17165 & ~n17166;
  assign n17168 = ~pi217 & ~n7798;
  assign n17169 = pi217 & n7798;
  assign n17170 = ~n17168 & ~n17169;
  assign n17171 = ~n7605 & n17170;
  assign n17172 = n7605 & ~n17170;
  assign n17173 = ~n17171 & ~n17172;
  assign n17174 = n17167 & n17173;
  assign n17175 = ~n17167 & ~n17173;
  assign n17176 = ~n17174 & ~n17175;
  assign n17177 = ~pi529 & n17176;
  assign po250 = n17161 | n17177;
  assign n17179 = ~pi151 & pi408;
  assign n17180 = pi151 & ~pi408;
  assign n17181 = ~n17179 & ~n17180;
  assign n17182 = pi529 & ~n17181;
  assign n17183 = ~pi151 & ~n7798;
  assign n17184 = pi151 & n7798;
  assign n17185 = ~n17183 & ~n17184;
  assign n17186 = n2586 & n17185;
  assign n17187 = ~n2586 & ~n17185;
  assign n17188 = ~n17186 & ~n17187;
  assign n17189 = ~n2689 & n17124;
  assign n17190 = n2689 & ~n17124;
  assign n17191 = ~n17189 & ~n17190;
  assign n17192 = ~n17188 & n17191;
  assign n17193 = n17188 & ~n17191;
  assign n17194 = ~n17192 & ~n17193;
  assign n17195 = ~pi529 & n17194;
  assign po251 = n17182 | n17195;
  assign n17197 = pi208 & pi449;
  assign n17198 = ~pi208 & ~pi449;
  assign n17199 = ~n17197 & ~n17198;
  assign n17200 = pi529 & ~n17199;
  assign n17201 = pi208 & ~n12862;
  assign n17202 = ~pi208 & n12862;
  assign n17203 = ~n17201 & ~n17202;
  assign n17204 = ~n12768 & n15917;
  assign n17205 = n12768 & ~n15917;
  assign n17206 = ~n17204 & ~n17205;
  assign n17207 = n17203 & ~n17206;
  assign n17208 = ~n17203 & n17206;
  assign n17209 = ~n17207 & ~n17208;
  assign n17210 = ~n15810 & n17209;
  assign n17211 = ~n15814 & ~n17209;
  assign n17212 = ~n17210 & ~n17211;
  assign n17213 = ~pi529 & n17212;
  assign po252 = n17200 | n17213;
  assign n17215 = ~pi346 & pi468;
  assign n17216 = pi346 & ~pi468;
  assign n17217 = ~n17215 & ~n17216;
  assign n17218 = pi529 & ~n17217;
  assign n17219 = n3755 & n16021;
  assign n17220 = ~n3755 & ~n16021;
  assign n17221 = ~n17219 & ~n17220;
  assign n17222 = n3591 & n17221;
  assign n17223 = ~n3591 & ~n17221;
  assign n17224 = ~n17222 & ~n17223;
  assign n17225 = ~pi346 & ~n12862;
  assign n17226 = pi346 & n12862;
  assign n17227 = ~n17225 & ~n17226;
  assign n17228 = ~n12768 & n17227;
  assign n17229 = n12768 & ~n17227;
  assign n17230 = ~n17228 & ~n17229;
  assign n17231 = n17224 & n17230;
  assign n17232 = ~n17224 & ~n17230;
  assign n17233 = ~n17231 & ~n17232;
  assign n17234 = ~pi529 & n17233;
  assign po253 = n17218 | n17234;
  assign n17236 = ~pi375 & ~n8140;
  assign n17237 = pi375 & n8140;
  assign n17238 = ~n17236 & ~n17237;
  assign n17239 = n11452 & n17238;
  assign n17240 = ~n11452 & ~n17238;
  assign n17241 = ~n17239 & ~n17240;
  assign n17242 = ~n3926 & n15484;
  assign n17243 = n3926 & ~n15484;
  assign n17244 = ~n17242 & ~n17243;
  assign n17245 = ~n15564 & n17244;
  assign n17246 = n15564 & ~n17244;
  assign n17247 = ~n17245 & ~n17246;
  assign n17248 = ~n17241 & ~n17247;
  assign n17249 = n17241 & n17247;
  assign n17250 = ~n17248 & ~n17249;
  assign n17251 = ~pi529 & ~n17250;
  assign n17252 = ~pi375 & pi528;
  assign n17253 = pi375 & ~pi528;
  assign n17254 = ~n17252 & ~n17253;
  assign n17255 = pi529 & ~n17254;
  assign po254 = n17251 | n17255;
  assign n17257 = ~pi210 & pi509;
  assign n17258 = pi210 & ~pi509;
  assign n17259 = ~n17257 & ~n17258;
  assign n17260 = pi529 & ~n17259;
  assign n17261 = ~pi210 & ~n8521;
  assign n17262 = pi210 & n8521;
  assign n17263 = ~n17261 & ~n17262;
  assign n17264 = n8848 & ~n14085;
  assign n17265 = ~n8848 & n14085;
  assign n17266 = ~n17264 & ~n17265;
  assign n17267 = ~n17263 & n17266;
  assign n17268 = n17263 & ~n17266;
  assign n17269 = ~n17267 & ~n17268;
  assign n17270 = ~n13243 & n17269;
  assign n17271 = ~n13247 & ~n17269;
  assign n17272 = ~n17270 & ~n17271;
  assign n17273 = ~pi529 & n17272;
  assign po255 = n17260 | n17273;
  assign n17275 = ~pi121 & pi130;
  assign n17276 = pi121 & ~pi130;
  assign n17277 = ~n17275 & ~n17276;
  assign n17278 = ~pi215 & pi233;
  assign n17279 = pi232 & n17278;
  assign n17280 = pi270 & n17279;
  assign n17281 = pi231 & n17280;
  assign n17282 = ~pi270 & n17279;
  assign n17283 = ~pi215 & ~pi232;
  assign n17284 = pi270 & n17283;
  assign n17285 = ~n17282 & ~n17284;
  assign n17286 = pi215 & ~pi233;
  assign n17287 = ~pi270 & n17286;
  assign n17288 = n17285 & ~n17287;
  assign n17289 = ~pi175 & ~pi231;
  assign n17290 = ~n17288 & n17289;
  assign n17291 = ~n17281 & ~n17290;
  assign n17292 = ~pi232 & n17278;
  assign n17293 = ~pi270 & n17292;
  assign n17294 = pi175 & n17293;
  assign n17295 = ~pi231 & n17294;
  assign n17296 = pi175 & pi231;
  assign n17297 = pi215 & pi232;
  assign n17298 = n17296 & n17297;
  assign n17299 = ~pi270 & n17298;
  assign n17300 = pi215 & pi233;
  assign n17301 = ~pi232 & n17300;
  assign n17302 = pi175 & n17301;
  assign n17303 = pi231 & n17302;
  assign n17304 = ~n17299 & ~n17303;
  assign n17305 = ~n17295 & n17304;
  assign n17306 = n17291 & n17305;
  assign n17307 = pi285 & ~n17306;
  assign n17308 = ~pi270 & n17300;
  assign n17309 = pi175 & n17308;
  assign n17310 = ~pi231 & ~pi285;
  assign n17311 = n17309 & n17310;
  assign n17312 = ~n17307 & ~n17311;
  assign n17313 = ~pi215 & ~pi233;
  assign n17314 = ~pi232 & n17313;
  assign n17315 = pi270 & n17314;
  assign n17316 = ~pi175 & n17315;
  assign n17317 = pi231 & n17316;
  assign n17318 = ~pi232 & n17286;
  assign n17319 = ~pi270 & n17318;
  assign n17320 = ~pi175 & pi231;
  assign n17321 = n17319 & n17320;
  assign n17322 = ~n17317 & ~n17321;
  assign n17323 = ~pi285 & ~n17322;
  assign n17324 = ~pi270 & n17301;
  assign n17325 = pi175 & n17324;
  assign n17326 = pi231 & n17325;
  assign n17327 = ~pi233 & ~pi270;
  assign n17328 = ~pi232 & n17327;
  assign n17329 = pi175 & n17328;
  assign n17330 = pi231 & n17329;
  assign n17331 = ~pi232 & pi233;
  assign n17332 = ~pi270 & n17331;
  assign n17333 = ~pi175 & n17332;
  assign n17334 = pi270 & n17313;
  assign n17335 = pi231 & n17334;
  assign n17336 = pi232 & pi233;
  assign n17337 = ~n17300 & ~n17336;
  assign n17338 = n17320 & ~n17337;
  assign n17339 = ~n17335 & ~n17338;
  assign n17340 = ~pi231 & n17280;
  assign n17341 = pi175 & n17340;
  assign n17342 = n17339 & ~n17341;
  assign n17343 = ~n17315 & n17342;
  assign n17344 = ~n17333 & n17343;
  assign n17345 = ~pi285 & ~n17344;
  assign n17346 = pi232 & n17300;
  assign n17347 = ~pi270 & n17346;
  assign n17348 = pi231 & n17347;
  assign n17349 = ~pi231 & n17282;
  assign n17350 = pi232 & n17286;
  assign n17351 = ~pi175 & pi270;
  assign n17352 = n17350 & n17351;
  assign n17353 = ~n17328 & ~n17352;
  assign n17354 = pi231 & ~n17353;
  assign n17355 = pi175 & n17292;
  assign n17356 = pi270 & n17346;
  assign n17357 = pi175 & n17356;
  assign n17358 = ~n17355 & ~n17357;
  assign n17359 = ~pi175 & n17347;
  assign n17360 = n17358 & ~n17359;
  assign n17361 = ~n17354 & n17360;
  assign n17362 = ~n17349 & n17361;
  assign n17363 = pi285 & ~n17362;
  assign n17364 = ~n17348 & ~n17363;
  assign n17365 = ~pi175 & n17356;
  assign n17366 = pi270 & n17286;
  assign n17367 = pi175 & n17366;
  assign n17368 = ~n17365 & ~n17367;
  assign n17369 = ~pi231 & ~n17368;
  assign n17370 = ~pi175 & n17319;
  assign n17371 = ~n17369 & ~n17370;
  assign n17372 = n17364 & n17371;
  assign n17373 = ~n17345 & n17372;
  assign n17374 = ~n17330 & n17373;
  assign n17375 = ~pi234 & ~n17374;
  assign n17376 = ~pi175 & n17280;
  assign n17377 = ~pi231 & n17376;
  assign n17378 = pi175 & n17346;
  assign n17379 = ~n17333 & ~n17378;
  assign n17380 = ~pi231 & ~n17379;
  assign n17381 = ~n17377 & ~n17380;
  assign n17382 = pi175 & ~pi270;
  assign n17383 = n17350 & n17382;
  assign n17384 = ~pi215 & pi232;
  assign n17385 = ~pi175 & n17384;
  assign n17386 = ~n17279 & ~n17385;
  assign n17387 = pi270 & n17331;
  assign n17388 = n17386 & ~n17387;
  assign n17389 = pi231 & ~n17388;
  assign n17390 = ~pi231 & n17314;
  assign n17391 = ~n17280 & ~n17302;
  assign n17392 = ~n17390 & n17391;
  assign n17393 = ~n17389 & n17392;
  assign n17394 = ~pi175 & n17286;
  assign n17395 = ~pi231 & n17394;
  assign n17396 = pi270 & n17336;
  assign n17397 = ~pi175 & n17396;
  assign n17398 = ~n17395 & ~n17397;
  assign n17399 = n17393 & n17398;
  assign n17400 = pi285 & ~n17399;
  assign n17401 = ~n17383 & ~n17400;
  assign n17402 = n17381 & n17401;
  assign n17403 = pi270 & n17292;
  assign n17404 = pi175 & n17403;
  assign n17405 = ~pi175 & ~pi270;
  assign n17406 = ~pi233 & n17405;
  assign n17407 = ~pi215 & n17406;
  assign n17408 = pi232 & ~pi233;
  assign n17409 = ~pi270 & n17408;
  assign n17410 = pi231 & n17409;
  assign n17411 = pi231 & n17350;
  assign n17412 = pi175 & ~pi231;
  assign n17413 = n17318 & n17412;
  assign n17414 = n17292 & n17296;
  assign n17415 = ~n17413 & ~n17414;
  assign n17416 = ~n17411 & n17415;
  assign n17417 = ~n17410 & n17416;
  assign n17418 = ~pi175 & n17301;
  assign n17419 = ~pi231 & n17418;
  assign n17420 = n17417 & ~n17419;
  assign n17421 = ~pi270 & n17297;
  assign n17422 = ~pi175 & n17421;
  assign n17423 = n17420 & ~n17422;
  assign n17424 = ~n17407 & n17423;
  assign n17425 = ~n17404 & n17424;
  assign n17426 = ~pi285 & ~n17425;
  assign n17427 = n17402 & ~n17426;
  assign n17428 = pi175 & n17278;
  assign n17429 = pi270 & n17428;
  assign n17430 = pi270 & n17318;
  assign n17431 = ~n17429 & ~n17430;
  assign n17432 = ~n17403 & n17431;
  assign n17433 = pi231 & ~n17432;
  assign n17434 = n17427 & ~n17433;
  assign n17435 = pi234 & ~n17434;
  assign n17436 = ~n17375 & ~n17435;
  assign n17437 = ~n17326 & n17436;
  assign n17438 = pi231 & n17404;
  assign n17439 = pi175 & n17430;
  assign n17440 = ~n17438 & ~n17439;
  assign n17441 = n17437 & n17440;
  assign n17442 = ~n17323 & n17441;
  assign n17443 = n17312 & n17442;
  assign n17444 = ~pi131 & n17443;
  assign n17445 = pi131 & ~n17443;
  assign n17446 = ~n17444 & ~n17445;
  assign n17447 = ~n17277 & n17446;
  assign n17448 = n17277 & ~n17446;
  assign n17449 = ~n17447 & ~n17448;
  assign n17450 = ~pi532 & ~n17449;
  assign n17451 = pi532 & pi584;
  assign po256 = n17450 | n17451;
  assign n17453 = ~pi371 & pi501;
  assign n17454 = pi371 & ~pi501;
  assign n17455 = ~n17453 & ~n17454;
  assign n17456 = pi529 & ~n17455;
  assign n17457 = n4786 & n16263;
  assign n17458 = ~n4786 & ~n16263;
  assign n17459 = ~n17457 & ~n17458;
  assign n17460 = n4620 & n17459;
  assign n17461 = ~n4620 & ~n17459;
  assign n17462 = ~n17460 & ~n17461;
  assign n17463 = pi371 & n8521;
  assign n17464 = ~pi371 & ~n8521;
  assign n17465 = ~n17463 & ~n17464;
  assign n17466 = ~n8848 & n17465;
  assign n17467 = n8848 & ~n17465;
  assign n17468 = ~n17466 & ~n17467;
  assign n17469 = n17462 & n17468;
  assign n17470 = ~n17462 & ~n17468;
  assign n17471 = ~n17469 & ~n17470;
  assign n17472 = ~pi529 & n17471;
  assign po257 = n17456 | n17472;
  assign n17474 = ~pi351 & pi404;
  assign n17475 = pi351 & ~pi404;
  assign n17476 = ~n17474 & ~n17475;
  assign n17477 = pi529 & ~n17476;
  assign n17478 = n6533 & n10672;
  assign n17479 = ~n6533 & ~n10672;
  assign n17480 = ~n17478 & ~n17479;
  assign n17481 = n10760 & n17480;
  assign n17482 = ~n10760 & ~n17480;
  assign n17483 = ~n17481 & ~n17482;
  assign n17484 = ~pi351 & ~n9771;
  assign n17485 = pi351 & n9771;
  assign n17486 = ~n17484 & ~n17485;
  assign n17487 = n11175 & n17486;
  assign n17488 = ~n11175 & ~n17486;
  assign n17489 = ~n17487 & ~n17488;
  assign n17490 = ~n17483 & n17489;
  assign n17491 = n17483 & ~n17489;
  assign n17492 = ~n17490 & ~n17491;
  assign n17493 = ~pi529 & n17492;
  assign po258 = n17477 | n17493;
  assign n17495 = ~pi258 & pi431;
  assign n17496 = pi258 & ~pi431;
  assign n17497 = ~n17495 & ~n17496;
  assign n17498 = pi529 & ~n17497;
  assign n17499 = n11313 & n15268;
  assign n17500 = ~n11313 & ~n15268;
  assign n17501 = ~n17499 & ~n17500;
  assign n17502 = n1627 & ~n10182;
  assign n17503 = ~n1627 & n10182;
  assign n17504 = ~n17502 & ~n17503;
  assign n17505 = pi258 & n17504;
  assign n17506 = ~pi258 & ~n17504;
  assign n17507 = ~n17505 & ~n17506;
  assign n17508 = ~n17501 & n17507;
  assign n17509 = n17501 & ~n17507;
  assign n17510 = ~n17508 & ~n17509;
  assign n17511 = ~pi529 & n17510;
  assign po259 = n17498 | n17511;
  assign n17513 = ~pi183 & pi480;
  assign n17514 = pi183 & ~pi480;
  assign n17515 = ~n17513 & ~n17514;
  assign n17516 = pi529 & ~n17515;
  assign n17517 = ~n2081 & n7405;
  assign n17518 = n2081 & ~n7405;
  assign n17519 = ~n17517 & ~n17518;
  assign n17520 = ~pi183 & ~n2365;
  assign n17521 = pi183 & n2365;
  assign n17522 = ~n17520 & ~n17521;
  assign n17523 = n2474 & n7504;
  assign n17524 = ~n2474 & ~n7504;
  assign n17525 = ~n17523 & ~n17524;
  assign n17526 = ~n17522 & n17525;
  assign n17527 = n17522 & ~n17525;
  assign n17528 = ~n17526 & ~n17527;
  assign n17529 = ~n17519 & n17528;
  assign n17530 = n17519 & ~n17528;
  assign n17531 = ~n17529 & ~n17530;
  assign n17532 = ~pi529 & n17531;
  assign po260 = n17516 | n17532;
  assign n17534 = ~pi348 & pi526;
  assign n17535 = pi348 & ~pi526;
  assign n17536 = ~n17534 & ~n17535;
  assign n17537 = pi529 & ~n17536;
  assign n17538 = ~n12970 & n15749;
  assign n17539 = n12970 & ~n15749;
  assign n17540 = ~n17538 & ~n17539;
  assign n17541 = n11452 & ~n15646;
  assign n17542 = ~n11452 & n15646;
  assign n17543 = ~n17541 & ~n17542;
  assign n17544 = pi348 & n17543;
  assign n17545 = ~pi348 & ~n17543;
  assign n17546 = ~n17544 & ~n17545;
  assign n17547 = ~n17540 & n17546;
  assign n17548 = n17540 & ~n17546;
  assign n17549 = ~n17547 & ~n17548;
  assign n17550 = ~pi529 & n17549;
  assign po261 = n17537 | n17550;
  assign n17552 = ~pi320 & pi406;
  assign n17553 = pi320 & ~pi406;
  assign n17554 = ~n17552 & ~n17553;
  assign n17555 = pi529 & ~n17554;
  assign n17556 = ~n11747 & n12163;
  assign n17557 = n11747 & ~n12163;
  assign n17558 = ~n17556 & ~n17557;
  assign n17559 = ~pi320 & ~n8140;
  assign n17560 = pi320 & n8140;
  assign n17561 = ~n17559 & ~n17560;
  assign n17562 = n11953 & n12252;
  assign n17563 = ~n11953 & ~n12252;
  assign n17564 = ~n17562 & ~n17563;
  assign n17565 = ~n17561 & n17564;
  assign n17566 = n17561 & ~n17564;
  assign n17567 = ~n17565 & ~n17566;
  assign n17568 = ~n17558 & n17567;
  assign n17569 = n17558 & ~n17567;
  assign n17570 = ~n17568 & ~n17569;
  assign n17571 = ~pi529 & n17570;
  assign po262 = n17555 | n17571;
  assign n17573 = ~pi228 & pi466;
  assign n17574 = pi228 & ~pi466;
  assign n17575 = ~n17573 & ~n17574;
  assign n17576 = pi529 & ~n17575;
  assign n17577 = ~pi228 & ~n8140;
  assign n17578 = pi228 & n8140;
  assign n17579 = ~n17577 & ~n17578;
  assign n17580 = n15646 & n17579;
  assign n17581 = ~n15646 & ~n17579;
  assign n17582 = ~n17580 & ~n17581;
  assign n17583 = ~n12970 & ~n15564;
  assign n17584 = n12970 & n15564;
  assign n17585 = ~n17583 & ~n17584;
  assign n17586 = ~n17582 & n17585;
  assign n17587 = n17582 & ~n17585;
  assign n17588 = ~n17586 & ~n17587;
  assign n17589 = ~pi529 & n17588;
  assign po263 = n17576 | n17589;
  assign n17591 = pi532 & pi562;
  assign n17592 = pi157 & pi354;
  assign n17593 = pi358 & n17592;
  assign n17594 = pi132 & n17593;
  assign n17595 = ~pi275 & ~pi354;
  assign n17596 = ~pi358 & n17595;
  assign n17597 = pi275 & ~pi354;
  assign n17598 = ~pi157 & n17597;
  assign n17599 = pi358 & n17598;
  assign n17600 = ~pi132 & n17599;
  assign n17601 = ~pi354 & ~pi358;
  assign n17602 = ~pi157 & n17601;
  assign n17603 = pi132 & n17602;
  assign n17604 = ~n17600 & ~n17603;
  assign n17605 = ~n17596 & n17604;
  assign n17606 = ~n17594 & n17605;
  assign n17607 = pi351 & ~n17606;
  assign n17608 = pi132 & pi351;
  assign n17609 = n17592 & n17608;
  assign n17610 = ~pi275 & pi354;
  assign n17611 = pi132 & n17610;
  assign n17612 = pi157 & ~pi275;
  assign n17613 = pi358 & n17612;
  assign n17614 = ~pi132 & n17613;
  assign n17615 = ~n17611 & ~n17614;
  assign n17616 = ~pi358 & n17597;
  assign n17617 = ~pi132 & n17616;
  assign n17618 = n17615 & ~n17617;
  assign n17619 = ~pi351 & ~n17618;
  assign n17620 = pi275 & pi354;
  assign n17621 = ~pi157 & n17620;
  assign n17622 = ~pi132 & n17621;
  assign n17623 = ~n17594 & ~n17622;
  assign n17624 = pi157 & n17597;
  assign n17625 = pi358 & n17624;
  assign n17626 = pi351 & n17625;
  assign n17627 = n17623 & ~n17626;
  assign n17628 = ~n17619 & n17627;
  assign n17629 = ~n17609 & n17628;
  assign n17630 = ~pi358 & n17624;
  assign n17631 = ~pi132 & n17630;
  assign n17632 = pi157 & n17610;
  assign n17633 = ~pi358 & n17632;
  assign n17634 = ~pi157 & n17595;
  assign n17635 = pi132 & n17634;
  assign n17636 = ~n17633 & ~n17635;
  assign n17637 = ~n17631 & n17636;
  assign n17638 = n17629 & n17637;
  assign n17639 = pi284 & ~n17638;
  assign n17640 = ~pi358 & n17621;
  assign n17641 = ~pi351 & n17640;
  assign n17642 = ~pi358 & n17634;
  assign n17643 = pi358 & n17632;
  assign n17644 = ~pi351 & n17643;
  assign n17645 = pi132 & ~pi351;
  assign n17646 = ~pi354 & pi358;
  assign n17647 = ~pi157 & n17646;
  assign n17648 = n17645 & n17647;
  assign n17649 = ~n17644 & ~n17648;
  assign n17650 = ~n17642 & n17649;
  assign n17651 = ~n17641 & n17650;
  assign n17652 = pi157 & n17620;
  assign n17653 = ~pi358 & n17652;
  assign n17654 = ~pi132 & n17653;
  assign n17655 = ~pi132 & n17634;
  assign n17656 = pi351 & n17655;
  assign n17657 = ~n17654 & ~n17656;
  assign n17658 = ~pi157 & ~pi275;
  assign n17659 = ~pi358 & n17658;
  assign n17660 = n17608 & n17659;
  assign n17661 = ~pi157 & n17610;
  assign n17662 = pi358 & n17661;
  assign n17663 = ~pi132 & n17662;
  assign n17664 = ~n17660 & ~n17663;
  assign n17665 = n17657 & n17664;
  assign n17666 = ~pi284 & ~n17665;
  assign n17667 = n17651 & ~n17666;
  assign n17668 = ~n17639 & n17667;
  assign n17669 = ~n17607 & n17668;
  assign n17670 = ~pi193 & ~n17669;
  assign n17671 = pi132 & n17624;
  assign n17672 = pi132 & n17616;
  assign n17673 = ~n17671 & ~n17672;
  assign n17674 = pi157 & ~pi354;
  assign n17675 = ~pi358 & n17674;
  assign n17676 = n17673 & ~n17675;
  assign n17677 = ~pi351 & ~n17676;
  assign n17678 = pi358 & n17652;
  assign n17679 = ~pi132 & n17678;
  assign n17680 = pi351 & n17679;
  assign n17681 = pi284 & ~pi351;
  assign n17682 = ~n17647 & ~n17659;
  assign n17683 = n17681 & ~n17682;
  assign n17684 = pi157 & pi284;
  assign n17685 = n17645 & n17684;
  assign n17686 = ~pi358 & n17685;
  assign n17687 = ~pi358 & n17610;
  assign n17688 = pi132 & n17687;
  assign n17689 = ~pi132 & n17643;
  assign n17690 = ~n17688 & ~n17689;
  assign n17691 = pi157 & n17595;
  assign n17692 = pi358 & n17691;
  assign n17693 = pi132 & n17692;
  assign n17694 = pi358 & n17634;
  assign n17695 = ~pi132 & n17694;
  assign n17696 = ~n17693 & ~n17695;
  assign n17697 = n17690 & n17696;
  assign n17698 = pi284 & ~n17697;
  assign n17699 = ~n17686 & ~n17698;
  assign n17700 = ~n17683 & n17699;
  assign n17701 = ~n17680 & n17700;
  assign n17702 = ~pi132 & pi351;
  assign n17703 = ~pi358 & n17598;
  assign n17704 = n17702 & n17703;
  assign n17705 = pi132 & pi358;
  assign n17706 = n17595 & n17705;
  assign n17707 = ~pi157 & pi275;
  assign n17708 = ~pi358 & n17707;
  assign n17709 = ~n17706 & ~n17708;
  assign n17710 = pi351 & n17709;
  assign n17711 = pi132 & n17661;
  assign n17712 = ~pi351 & ~n17711;
  assign n17713 = ~n17710 & ~n17712;
  assign n17714 = ~pi351 & n17624;
  assign n17715 = ~n17671 & ~n17679;
  assign n17716 = ~n17714 & n17715;
  assign n17717 = ~n17713 & n17716;
  assign n17718 = ~pi284 & ~n17717;
  assign n17719 = ~n17704 & ~n17718;
  assign n17720 = pi358 & n17621;
  assign n17721 = ~pi351 & n17720;
  assign n17722 = pi132 & ~pi358;
  assign n17723 = n17624 & n17722;
  assign n17724 = ~n17721 & ~n17723;
  assign n17725 = n17719 & n17724;
  assign n17726 = n17701 & n17725;
  assign n17727 = ~n17677 & n17726;
  assign n17728 = pi193 & ~n17727;
  assign n17729 = ~n17670 & ~n17728;
  assign n17730 = pi132 & n17642;
  assign n17731 = ~n17644 & ~n17730;
  assign n17732 = pi284 & ~n17731;
  assign n17733 = ~pi132 & ~pi351;
  assign n17734 = ~pi358 & n17592;
  assign n17735 = n17733 & n17734;
  assign n17736 = ~n17721 & ~n17735;
  assign n17737 = pi132 & n17625;
  assign n17738 = ~pi351 & n17737;
  assign n17739 = n17736 & ~n17738;
  assign n17740 = ~pi284 & ~n17739;
  assign n17741 = ~pi132 & ~pi358;
  assign n17742 = ~pi354 & n17741;
  assign n17743 = ~pi275 & n17742;
  assign n17744 = pi132 & n17613;
  assign n17745 = ~pi132 & pi358;
  assign n17746 = ~n17598 & ~n17661;
  assign n17747 = n17745 & ~n17746;
  assign n17748 = ~n17744 & ~n17747;
  assign n17749 = ~n17679 & n17748;
  assign n17750 = pi351 & ~n17749;
  assign n17751 = ~n17743 & ~n17750;
  assign n17752 = ~pi284 & ~n17751;
  assign n17753 = ~n17740 & ~n17752;
  assign n17754 = n17625 & n17702;
  assign n17755 = pi284 & n17754;
  assign n17756 = n17753 & ~n17755;
  assign n17757 = ~n17732 & n17756;
  assign n17758 = ~pi358 & n17691;
  assign n17759 = pi132 & n17758;
  assign n17760 = ~pi351 & n17759;
  assign n17761 = pi351 & n17693;
  assign n17762 = ~n17760 & ~n17761;
  assign n17763 = ~pi351 & n17622;
  assign n17764 = n17762 & ~n17763;
  assign n17765 = n17757 & n17764;
  assign n17766 = n17729 & n17765;
  assign n17767 = pi388 & n17766;
  assign n17768 = ~pi388 & ~n17766;
  assign n17769 = ~n17767 & ~n17768;
  assign n17770 = pi140 & pi144;
  assign n17771 = ~pi140 & ~pi144;
  assign n17772 = ~n17770 & ~n17771;
  assign n17773 = pi129 & ~pi141;
  assign n17774 = ~pi129 & pi141;
  assign n17775 = ~n17773 & ~n17774;
  assign n17776 = ~n17772 & n17775;
  assign n17777 = n17772 & ~n17775;
  assign n17778 = ~n17776 & ~n17777;
  assign n17779 = ~n17769 & n17778;
  assign n17780 = ~pi388 & n17766;
  assign n17781 = pi388 & ~n17766;
  assign n17782 = ~n17780 & ~n17781;
  assign n17783 = ~n17778 & ~n17782;
  assign n17784 = ~n17779 & ~n17783;
  assign n17785 = ~pi532 & ~n17784;
  assign po264 = n17591 | n17785;
  assign n17787 = pi532 & pi648;
  assign n17788 = pi130 & n17443;
  assign n17789 = ~pi130 & ~n17443;
  assign n17790 = ~n17788 & ~n17789;
  assign n17791 = ~pi532 & ~n17790;
  assign po265 = n17787 | n17791;
  assign n17793 = pi532 & pi616;
  assign n17794 = ~pi130 & ~pi131;
  assign n17795 = pi130 & pi131;
  assign n17796 = ~n17794 & ~n17795;
  assign n17797 = n17443 & ~n17796;
  assign n17798 = ~n17443 & n17796;
  assign n17799 = ~n17797 & ~n17798;
  assign n17800 = ~pi532 & ~n17799;
  assign po266 = n17793 | n17800;
  assign n17802 = pi532 & pi552;
  assign n17803 = ~pi121 & ~pi131;
  assign n17804 = pi121 & pi131;
  assign n17805 = ~n17803 & ~n17804;
  assign n17806 = ~pi130 & pi132;
  assign n17807 = pi130 & ~pi132;
  assign n17808 = ~n17806 & ~n17807;
  assign n17809 = ~n17805 & n17808;
  assign n17810 = n17805 & ~n17808;
  assign n17811 = ~n17809 & ~n17810;
  assign n17812 = n17443 & ~n17811;
  assign n17813 = ~n17443 & n17811;
  assign n17814 = ~n17812 & ~n17813;
  assign n17815 = ~pi532 & ~n17814;
  assign po267 = n17802 | n17815;
  assign n17817 = ~pi133 & pi148;
  assign n17818 = pi133 & ~pi148;
  assign n17819 = ~n17817 & ~n17818;
  assign n17820 = pi175 & n17350;
  assign n17821 = pi175 & n17287;
  assign n17822 = ~n17820 & ~n17821;
  assign n17823 = ~n17409 & n17822;
  assign n17824 = ~pi231 & ~n17823;
  assign n17825 = pi231 & n17365;
  assign n17826 = ~pi231 & pi285;
  assign n17827 = ~pi270 & n17283;
  assign n17828 = ~pi233 & pi270;
  assign n17829 = ~pi232 & n17828;
  assign n17830 = ~n17827 & ~n17829;
  assign n17831 = n17826 & ~n17830;
  assign n17832 = pi175 & pi232;
  assign n17833 = n17826 & n17832;
  assign n17834 = ~pi270 & n17833;
  assign n17835 = pi232 & n17313;
  assign n17836 = pi270 & n17835;
  assign n17837 = pi175 & n17836;
  assign n17838 = ~pi270 & n17278;
  assign n17839 = pi175 & n17838;
  assign n17840 = ~n17376 & ~n17839;
  assign n17841 = ~n17837 & n17840;
  assign n17842 = ~n17316 & n17841;
  assign n17843 = pi285 & ~n17842;
  assign n17844 = ~n17834 & ~n17843;
  assign n17845 = ~n17831 & n17844;
  assign n17846 = ~n17825 & n17845;
  assign n17847 = pi175 & pi270;
  assign n17848 = n17313 & n17847;
  assign n17849 = pi215 & ~pi232;
  assign n17850 = ~pi270 & n17849;
  assign n17851 = ~n17848 & ~n17850;
  assign n17852 = pi231 & n17851;
  assign n17853 = ~pi231 & ~n17355;
  assign n17854 = ~n17852 & ~n17853;
  assign n17855 = ~pi231 & n17350;
  assign n17856 = ~n17365 & ~n17820;
  assign n17857 = ~n17855 & n17856;
  assign n17858 = ~n17854 & n17857;
  assign n17859 = ~pi285 & ~n17858;
  assign n17860 = ~n17321 & ~n17859;
  assign n17861 = pi270 & n17301;
  assign n17862 = ~pi231 & n17861;
  assign n17863 = ~n17383 & ~n17862;
  assign n17864 = n17860 & n17863;
  assign n17865 = n17846 & n17864;
  assign n17866 = ~n17824 & n17865;
  assign n17867 = pi234 & ~n17866;
  assign n17868 = ~pi175 & n17314;
  assign n17869 = pi231 & n17868;
  assign n17870 = ~n17359 & ~n17869;
  assign n17871 = n17296 & n17827;
  assign n17872 = ~pi175 & n17403;
  assign n17873 = ~n17871 & ~n17872;
  assign n17874 = n17870 & n17873;
  assign n17875 = ~pi285 & ~n17874;
  assign n17876 = pi270 & n17384;
  assign n17877 = ~pi175 & n17876;
  assign n17878 = ~pi175 & n17287;
  assign n17879 = ~n17428 & ~n17878;
  assign n17880 = ~n17877 & n17879;
  assign n17881 = ~pi231 & ~n17880;
  assign n17882 = n17296 & n17336;
  assign n17883 = ~n17881 & ~n17882;
  assign n17884 = pi270 & n17350;
  assign n17885 = pi231 & n17884;
  assign n17886 = pi175 & n17314;
  assign n17887 = ~pi270 & n17350;
  assign n17888 = ~pi175 & n17887;
  assign n17889 = ~n17886 & ~n17888;
  assign n17890 = ~n17282 & n17889;
  assign n17891 = pi175 & n17396;
  assign n17892 = ~n17418 & ~n17891;
  assign n17893 = n17890 & n17892;
  assign n17894 = ~n17885 & n17893;
  assign n17895 = n17883 & n17894;
  assign n17896 = pi285 & ~n17895;
  assign n17897 = ~pi270 & n17313;
  assign n17898 = ~pi175 & n17430;
  assign n17899 = ~n17329 & ~n17898;
  assign n17900 = ~n17897 & n17899;
  assign n17901 = ~n17891 & n17900;
  assign n17902 = pi231 & ~n17901;
  assign n17903 = ~n17896 & ~n17902;
  assign n17904 = ~n17875 & n17903;
  assign n17905 = ~pi231 & n17324;
  assign n17906 = ~pi270 & n17314;
  assign n17907 = n17412 & n17829;
  assign n17908 = ~n17340 & ~n17907;
  assign n17909 = ~n17906 & n17908;
  assign n17910 = ~n17905 & n17909;
  assign n17911 = n17904 & n17910;
  assign n17912 = ~pi234 & ~n17911;
  assign n17913 = ~n17867 & ~n17912;
  assign n17914 = ~pi270 & n17336;
  assign n17915 = n17289 & n17914;
  assign n17916 = ~n17862 & ~n17915;
  assign n17917 = pi232 & n17847;
  assign n17918 = n17286 & n17917;
  assign n17919 = ~pi231 & n17918;
  assign n17920 = n17916 & ~n17919;
  assign n17921 = pi175 & n17876;
  assign n17922 = ~n17292 & ~n17318;
  assign n17923 = n17351 & ~n17922;
  assign n17924 = ~n17921 & ~n17923;
  assign n17925 = ~n17365 & n17924;
  assign n17926 = pi231 & ~n17925;
  assign n17927 = ~n17407 & ~n17926;
  assign n17928 = n17920 & n17927;
  assign n17929 = ~pi285 & ~n17928;
  assign n17930 = pi231 & pi285;
  assign n17931 = n17352 & n17930;
  assign n17932 = ~n17929 & ~n17931;
  assign n17933 = pi175 & n17906;
  assign n17934 = ~n17340 & ~n17933;
  assign n17935 = pi285 & ~n17934;
  assign n17936 = n17932 & ~n17935;
  assign n17937 = ~pi270 & n17835;
  assign n17938 = pi175 & n17937;
  assign n17939 = ~pi231 & n17938;
  assign n17940 = pi231 & n17837;
  assign n17941 = ~n17939 & ~n17940;
  assign n17942 = ~n17419 & n17941;
  assign n17943 = n17936 & n17942;
  assign n17944 = n17913 & n17943;
  assign n17945 = ~pi149 & n17944;
  assign n17946 = pi149 & ~n17944;
  assign n17947 = ~n17945 & ~n17946;
  assign n17948 = ~n17819 & n17947;
  assign n17949 = n17819 & ~n17947;
  assign n17950 = ~n17948 & ~n17949;
  assign n17951 = ~pi532 & ~n17950;
  assign n17952 = pi532 & pi586;
  assign po268 = n17951 | n17952;
  assign n17954 = pi351 & n17603;
  assign n17955 = pi358 & n17595;
  assign n17956 = pi351 & n17955;
  assign n17957 = ~n17592 & ~n17620;
  assign n17958 = n17702 & ~n17957;
  assign n17959 = ~n17956 & ~n17958;
  assign n17960 = pi132 & n17644;
  assign n17961 = n17959 & ~n17960;
  assign n17962 = ~pi157 & pi354;
  assign n17963 = ~pi358 & n17962;
  assign n17964 = ~pi132 & n17963;
  assign n17965 = ~n17694 & ~n17964;
  assign n17966 = n17961 & n17965;
  assign n17967 = ~pi284 & ~n17966;
  assign n17968 = pi351 & n17653;
  assign n17969 = ~pi351 & n17633;
  assign n17970 = n17624 & n17745;
  assign n17971 = ~n17602 & ~n17970;
  assign n17972 = pi351 & ~n17971;
  assign n17973 = pi132 & n17678;
  assign n17974 = ~n17711 & ~n17973;
  assign n17975 = ~n17654 & n17974;
  assign n17976 = ~n17972 & n17975;
  assign n17977 = ~n17969 & n17976;
  assign n17978 = pi284 & ~n17977;
  assign n17979 = ~n17968 & ~n17978;
  assign n17980 = pi358 & n17597;
  assign n17981 = pi132 & n17980;
  assign n17982 = ~n17679 & ~n17981;
  assign n17983 = ~pi351 & ~n17982;
  assign n17984 = ~pi132 & n17703;
  assign n17985 = ~n17983 & ~n17984;
  assign n17986 = n17979 & n17985;
  assign n17987 = ~n17967 & n17986;
  assign n17988 = ~n17954 & n17987;
  assign n17989 = ~pi193 & ~n17988;
  assign n17990 = pi351 & n17695;
  assign n17991 = ~n17704 & ~n17990;
  assign n17992 = ~pi284 & ~n17991;
  assign n17993 = ~pi132 & n17612;
  assign n17994 = ~n17632 & ~n17993;
  assign n17995 = pi358 & n17962;
  assign n17996 = n17994 & ~n17995;
  assign n17997 = pi351 & ~n17996;
  assign n17998 = ~pi351 & n17634;
  assign n17999 = pi132 & n17621;
  assign n18000 = ~n17643 & ~n17999;
  assign n18001 = ~n17998 & n18000;
  assign n18002 = ~n17997 & n18001;
  assign n18003 = ~pi132 & n17597;
  assign n18004 = ~pi351 & n18003;
  assign n18005 = ~pi132 & n17593;
  assign n18006 = ~n18004 & ~n18005;
  assign n18007 = n18002 & n18006;
  assign n18008 = pi284 & ~n18007;
  assign n18009 = ~pi351 & n17689;
  assign n18010 = pi132 & n17652;
  assign n18011 = ~n17964 & ~n18010;
  assign n18012 = ~pi351 & ~n18011;
  assign n18013 = ~n18009 & ~n18012;
  assign n18014 = pi132 & n17662;
  assign n18015 = pi351 & n17675;
  assign n18016 = pi351 & n17624;
  assign n18017 = n17598 & n17645;
  assign n18018 = n17608 & n17661;
  assign n18019 = ~n18017 & ~n18018;
  assign n18020 = ~n18016 & n18019;
  assign n18021 = ~n18015 & n18020;
  assign n18022 = ~n17763 & n18021;
  assign n18023 = pi157 & pi275;
  assign n18024 = ~pi358 & n18023;
  assign n18025 = ~pi132 & n18024;
  assign n18026 = n18022 & ~n18025;
  assign n18027 = ~n17743 & n18026;
  assign n18028 = ~n18014 & n18027;
  assign n18029 = ~pi284 & ~n18028;
  assign n18030 = ~n17723 & ~n18029;
  assign n18031 = n18013 & n18030;
  assign n18032 = ~n18008 & n18031;
  assign n18033 = ~n17599 & ~n17662;
  assign n18034 = pi358 & n17611;
  assign n18035 = n18033 & ~n18034;
  assign n18036 = pi351 & ~n18035;
  assign n18037 = n18032 & ~n18036;
  assign n18038 = pi193 & ~n18037;
  assign n18039 = ~n17992 & ~n18038;
  assign n18040 = ~n17989 & n18039;
  assign n18041 = pi132 & n17640;
  assign n18042 = pi351 & n18041;
  assign n18043 = pi351 & n18014;
  assign n18044 = pi351 & n17643;
  assign n18045 = pi358 & n17658;
  assign n18046 = ~n17616 & ~n17633;
  assign n18047 = ~n18045 & n18046;
  assign n18048 = n17733 & ~n18047;
  assign n18049 = ~n18044 & ~n18048;
  assign n18050 = ~pi358 & n17661;
  assign n18051 = pi132 & n18050;
  assign n18052 = ~pi351 & n18051;
  assign n18053 = n17608 & n18023;
  assign n18054 = ~pi358 & n18053;
  assign n18055 = pi351 & n17999;
  assign n18056 = ~n18054 & ~n18055;
  assign n18057 = ~n18052 & n18056;
  assign n18058 = n18049 & n18057;
  assign n18059 = pi284 & ~n18058;
  assign n18060 = ~pi284 & ~pi351;
  assign n18061 = ~pi358 & n17620;
  assign n18062 = pi132 & n18061;
  assign n18063 = n18060 & n18062;
  assign n18064 = ~n18059 & ~n18063;
  assign n18065 = pi132 & n17599;
  assign n18066 = n18064 & ~n18065;
  assign n18067 = ~n18043 & n18066;
  assign n18068 = ~n18042 & n18067;
  assign n18069 = n18040 & n18068;
  assign n18070 = pi134 & n18069;
  assign n18071 = ~pi134 & ~n18069;
  assign n18072 = ~n18070 & ~n18071;
  assign n18073 = pi386 & n18072;
  assign n18074 = ~pi386 & ~n18072;
  assign n18075 = ~n18073 & ~n18074;
  assign n18076 = ~pi532 & ~n18075;
  assign n18077 = pi532 & pi656;
  assign po269 = n18076 | n18077;
  assign n18079 = ~pi134 & ~pi135;
  assign n18080 = pi134 & pi135;
  assign n18081 = ~n18079 & ~n18080;
  assign n18082 = pi386 & n18069;
  assign n18083 = ~pi386 & ~n18069;
  assign n18084 = ~n18082 & ~n18083;
  assign n18085 = ~n18081 & n18084;
  assign n18086 = n18081 & ~n18084;
  assign n18087 = ~n18085 & ~n18086;
  assign n18088 = ~pi532 & ~n18087;
  assign n18089 = pi532 & pi624;
  assign po270 = n18088 | n18089;
  assign n18091 = ~pi134 & pi136;
  assign n18092 = pi134 & ~pi136;
  assign n18093 = ~n18091 & ~n18092;
  assign n18094 = pi386 & n18093;
  assign n18095 = ~pi386 & ~n18093;
  assign n18096 = ~n18094 & ~n18095;
  assign n18097 = ~pi135 & n18069;
  assign n18098 = pi135 & ~n18069;
  assign n18099 = ~n18097 & ~n18098;
  assign n18100 = ~n18096 & n18099;
  assign n18101 = n18096 & ~n18099;
  assign n18102 = ~n18100 & ~n18101;
  assign n18103 = ~pi532 & ~n18102;
  assign n18104 = pi532 & pi592;
  assign po271 = n18103 | n18104;
  assign n18106 = ~pi137 & pi171;
  assign n18107 = pi137 & ~pi171;
  assign n18108 = ~n18106 & ~n18107;
  assign n18109 = ~pi170 & ~pi342;
  assign n18110 = ~pi321 & n18109;
  assign n18111 = pi182 & n18110;
  assign n18112 = pi352 & n18111;
  assign n18113 = ~pi170 & pi342;
  assign n18114 = ~pi321 & n18113;
  assign n18115 = ~pi182 & n18114;
  assign n18116 = ~pi276 & ~pi342;
  assign n18117 = ~pi170 & n18116;
  assign n18118 = pi321 & n18117;
  assign n18119 = ~pi182 & pi352;
  assign n18120 = pi276 & pi342;
  assign n18121 = pi170 & pi342;
  assign n18122 = ~n18120 & ~n18121;
  assign n18123 = n18119 & ~n18122;
  assign n18124 = pi321 & pi352;
  assign n18125 = n18116 & n18124;
  assign n18126 = ~n18123 & ~n18125;
  assign n18127 = ~pi276 & pi342;
  assign n18128 = pi170 & n18127;
  assign n18129 = pi321 & n18128;
  assign n18130 = ~pi352 & n18129;
  assign n18131 = pi182 & n18130;
  assign n18132 = n18126 & ~n18131;
  assign n18133 = ~n18118 & n18132;
  assign n18134 = ~n18115 & n18133;
  assign n18135 = ~pi372 & ~n18134;
  assign n18136 = ~pi170 & pi276;
  assign n18137 = ~pi342 & n18136;
  assign n18138 = ~pi321 & n18137;
  assign n18139 = ~pi182 & n18138;
  assign n18140 = pi276 & ~pi342;
  assign n18141 = pi321 & n18140;
  assign n18142 = pi182 & n18141;
  assign n18143 = pi170 & n18120;
  assign n18144 = pi321 & n18143;
  assign n18145 = ~pi182 & n18144;
  assign n18146 = ~n18142 & ~n18145;
  assign n18147 = ~pi352 & ~n18146;
  assign n18148 = ~n18139 & ~n18147;
  assign n18149 = ~pi321 & n18143;
  assign n18150 = pi352 & n18149;
  assign n18151 = n18148 & ~n18150;
  assign n18152 = pi170 & n18140;
  assign n18153 = ~pi182 & pi321;
  assign n18154 = n18152 & n18153;
  assign n18155 = ~n18110 & ~n18154;
  assign n18156 = pi352 & n18155;
  assign n18157 = ~pi321 & n18128;
  assign n18158 = ~pi352 & ~n18157;
  assign n18159 = ~n18156 & ~n18158;
  assign n18160 = ~pi182 & n18149;
  assign n18161 = ~pi170 & n18127;
  assign n18162 = pi182 & n18161;
  assign n18163 = pi182 & n18144;
  assign n18164 = ~n18162 & ~n18163;
  assign n18165 = ~n18160 & n18164;
  assign n18166 = ~n18159 & n18165;
  assign n18167 = pi372 & ~n18166;
  assign n18168 = n18151 & ~n18167;
  assign n18169 = ~n18135 & n18168;
  assign n18170 = ~n18112 & n18169;
  assign n18171 = ~pi191 & ~n18170;
  assign n18172 = pi321 & n18113;
  assign n18173 = pi170 & ~pi276;
  assign n18174 = ~pi182 & n18173;
  assign n18175 = ~n18172 & ~n18174;
  assign n18176 = ~n18128 & n18175;
  assign n18177 = pi352 & ~n18176;
  assign n18178 = ~pi182 & n18140;
  assign n18179 = ~pi352 & n18178;
  assign n18180 = ~n18177 & ~n18179;
  assign n18181 = pi321 & n18121;
  assign n18182 = ~pi182 & n18181;
  assign n18183 = ~pi352 & n18117;
  assign n18184 = ~n18129 & ~n18183;
  assign n18185 = ~pi170 & n18120;
  assign n18186 = pi182 & n18185;
  assign n18187 = n18184 & ~n18186;
  assign n18188 = ~n18182 & n18187;
  assign n18189 = n18180 & n18188;
  assign n18190 = pi372 & ~n18189;
  assign n18191 = ~pi321 & n18152;
  assign n18192 = pi182 & n18191;
  assign n18193 = pi182 & n18143;
  assign n18194 = ~n18115 & ~n18193;
  assign n18195 = ~pi352 & ~n18194;
  assign n18196 = ~n18192 & ~n18195;
  assign n18197 = pi352 & n18152;
  assign n18198 = pi182 & pi352;
  assign n18199 = n18161 & n18198;
  assign n18200 = pi170 & ~pi342;
  assign n18201 = ~pi321 & n18200;
  assign n18202 = pi352 & n18201;
  assign n18203 = ~n18199 & ~n18202;
  assign n18204 = ~n18197 & n18203;
  assign n18205 = pi182 & ~pi352;
  assign n18206 = n18137 & n18205;
  assign n18207 = n18204 & ~n18206;
  assign n18208 = ~pi182 & n18185;
  assign n18209 = ~pi352 & n18208;
  assign n18210 = ~pi321 & n18116;
  assign n18211 = ~pi182 & n18210;
  assign n18212 = pi321 & n18161;
  assign n18213 = pi182 & n18212;
  assign n18214 = ~n18211 & ~n18213;
  assign n18215 = ~pi182 & ~pi321;
  assign n18216 = pi170 & pi276;
  assign n18217 = n18215 & n18216;
  assign n18218 = n18214 & ~n18217;
  assign n18219 = ~n18209 & n18218;
  assign n18220 = n18207 & n18219;
  assign n18221 = ~pi372 & ~n18220;
  assign n18222 = ~pi182 & n18129;
  assign n18223 = ~pi352 & n18222;
  assign n18224 = ~n18221 & ~n18223;
  assign n18225 = n18196 & n18224;
  assign n18226 = ~n18190 & n18225;
  assign n18227 = pi321 & n18137;
  assign n18228 = pi182 & n18127;
  assign n18229 = pi321 & n18228;
  assign n18230 = ~n18227 & ~n18229;
  assign n18231 = ~n18212 & n18230;
  assign n18232 = pi352 & ~n18231;
  assign n18233 = n18226 & ~n18232;
  assign n18234 = pi191 & ~n18233;
  assign n18235 = ~n18171 & ~n18234;
  assign n18236 = pi352 & n18139;
  assign n18237 = ~pi182 & n18118;
  assign n18238 = pi352 & n18237;
  assign n18239 = ~n18236 & ~n18238;
  assign n18240 = ~pi372 & ~n18239;
  assign n18241 = n18235 & ~n18240;
  assign n18242 = ~pi321 & n18185;
  assign n18243 = pi182 & n18242;
  assign n18244 = pi352 & n18243;
  assign n18245 = pi182 & n18227;
  assign n18246 = pi352 & n18129;
  assign n18247 = ~pi170 & ~pi276;
  assign n18248 = pi321 & n18247;
  assign n18249 = ~pi321 & n18140;
  assign n18250 = ~n18248 & ~n18249;
  assign n18251 = ~n18157 & n18250;
  assign n18252 = ~pi182 & ~pi352;
  assign n18253 = ~n18251 & n18252;
  assign n18254 = ~n18246 & ~n18253;
  assign n18255 = ~pi321 & n18161;
  assign n18256 = pi182 & n18255;
  assign n18257 = ~pi352 & n18256;
  assign n18258 = n18198 & n18216;
  assign n18259 = ~pi321 & n18258;
  assign n18260 = pi352 & n18186;
  assign n18261 = ~n18259 & ~n18260;
  assign n18262 = ~n18257 & n18261;
  assign n18263 = n18254 & n18262;
  assign n18264 = pi372 & ~n18263;
  assign n18265 = ~pi352 & ~pi372;
  assign n18266 = ~pi321 & n18120;
  assign n18267 = pi182 & n18266;
  assign n18268 = n18265 & n18267;
  assign n18269 = ~n18264 & ~n18268;
  assign n18270 = pi352 & n18213;
  assign n18271 = n18269 & ~n18270;
  assign n18272 = ~n18245 & n18271;
  assign n18273 = ~n18244 & n18272;
  assign n18274 = n18241 & n18273;
  assign n18275 = pi172 & n18274;
  assign n18276 = ~pi172 & ~n18274;
  assign n18277 = ~n18275 & ~n18276;
  assign n18278 = ~n18108 & n18277;
  assign n18279 = n18108 & ~n18277;
  assign n18280 = ~n18278 & ~n18279;
  assign n18281 = ~pi532 & ~n18280;
  assign n18282 = pi532 & pi576;
  assign po272 = n18281 | n18282;
  assign n18284 = ~pi135 & ~pi136;
  assign n18285 = pi135 & pi136;
  assign n18286 = ~n18284 & ~n18285;
  assign n18287 = ~pi134 & pi138;
  assign n18288 = pi134 & ~pi138;
  assign n18289 = ~n18287 & ~n18288;
  assign n18290 = ~n18286 & n18289;
  assign n18291 = n18286 & ~n18289;
  assign n18292 = ~n18290 & ~n18291;
  assign n18293 = n18084 & ~n18292;
  assign n18294 = ~n18084 & n18292;
  assign n18295 = ~n18293 & ~n18294;
  assign n18296 = ~pi532 & ~n18295;
  assign n18297 = pi532 & pi560;
  assign po273 = n18296 | n18297;
  assign n18299 = pi532 & pi557;
  assign n18300 = ~pi351 & n17706;
  assign n18301 = ~n17653 & ~n17703;
  assign n18302 = ~pi132 & ~n18301;
  assign n18303 = ~n18300 & ~n18302;
  assign n18304 = ~pi284 & ~n18303;
  assign n18305 = ~pi284 & n17592;
  assign n18306 = n17702 & n18305;
  assign n18307 = ~n18304 & ~n18306;
  assign n18308 = ~pi132 & n17595;
  assign n18309 = n17620 & n17705;
  assign n18310 = pi351 & n17671;
  assign n18311 = n17733 & n17962;
  assign n18312 = ~n18310 & ~n18311;
  assign n18313 = ~n18309 & n18312;
  assign n18314 = ~n18308 & n18313;
  assign n18315 = ~n17596 & n18314;
  assign n18316 = pi284 & ~n18315;
  assign n18317 = ~pi284 & pi351;
  assign n18318 = n17632 & n18317;
  assign n18319 = ~n17691 & ~n17707;
  assign n18320 = n17608 & ~n18319;
  assign n18321 = ~pi358 & n18320;
  assign n18322 = ~n18318 & ~n18321;
  assign n18323 = ~n18316 & n18322;
  assign n18324 = n18307 & n18323;
  assign n18325 = ~pi132 & n17659;
  assign n18326 = ~n17689 & ~n18325;
  assign n18327 = ~n18010 & n18326;
  assign n18328 = ~pi351 & ~n18327;
  assign n18329 = n18324 & ~n18328;
  assign n18330 = ~pi193 & ~n18329;
  assign n18331 = pi351 & ~n17631;
  assign n18332 = ~pi351 & ~n18309;
  assign n18333 = ~n18331 & ~n18332;
  assign n18334 = ~n17625 & ~n17655;
  assign n18335 = ~n17720 & n18334;
  assign n18336 = pi351 & ~n18335;
  assign n18337 = n17662 & n17733;
  assign n18338 = ~n18336 & ~n18337;
  assign n18339 = ~pi157 & n17722;
  assign n18340 = ~n17688 & ~n18339;
  assign n18341 = ~pi132 & n17675;
  assign n18342 = n18340 & ~n18341;
  assign n18343 = n18338 & n18342;
  assign n18344 = ~pi284 & ~n18343;
  assign n18345 = pi132 & n17734;
  assign n18346 = ~n17693 & ~n18345;
  assign n18347 = ~n17689 & n18346;
  assign n18348 = ~n18050 & n18347;
  assign n18349 = pi351 & ~n18348;
  assign n18350 = pi132 & ~pi354;
  assign n18351 = ~pi358 & n18350;
  assign n18352 = pi132 & n17707;
  assign n18353 = ~n18351 & ~n18352;
  assign n18354 = ~pi351 & ~n18353;
  assign n18355 = n17674 & n17745;
  assign n18356 = ~n17678 & ~n18355;
  assign n18357 = ~pi351 & ~n18356;
  assign n18358 = ~n18354 & ~n18357;
  assign n18359 = ~n18349 & n18358;
  assign n18360 = ~pi132 & n17624;
  assign n18361 = ~n18051 & ~n18360;
  assign n18362 = ~pi351 & n18023;
  assign n18363 = ~n17998 & ~n18362;
  assign n18364 = ~n17599 & n18363;
  assign n18365 = pi284 & ~n18364;
  assign n18366 = n18361 & ~n18365;
  assign n18367 = n18359 & n18366;
  assign n18368 = ~n18344 & n18367;
  assign n18369 = pi193 & ~n18368;
  assign n18370 = ~pi351 & n17723;
  assign n18371 = ~pi132 & n17758;
  assign n18372 = ~pi132 & n17980;
  assign n18373 = ~pi132 & n17598;
  assign n18374 = ~n18372 & ~n18373;
  assign n18375 = ~n18371 & n18374;
  assign n18376 = ~pi351 & ~n18375;
  assign n18377 = ~n18370 & ~n18376;
  assign n18378 = ~n17761 & n18377;
  assign n18379 = ~pi284 & ~n18378;
  assign n18380 = pi351 & n17600;
  assign n18381 = ~pi351 & n18005;
  assign n18382 = ~n18380 & ~n18381;
  assign n18383 = ~pi157 & n17741;
  assign n18384 = n17595 & n18383;
  assign n18385 = ~n17759 & ~n18384;
  assign n18386 = ~n18018 & n18385;
  assign n18387 = n18382 & n18386;
  assign n18388 = pi284 & ~n18387;
  assign n18389 = ~n18379 & ~n18388;
  assign n18390 = pi351 & n18025;
  assign n18391 = ~pi132 & n18050;
  assign n18392 = pi351 & n18391;
  assign n18393 = ~n18390 & ~n18392;
  assign n18394 = ~pi284 & ~n18393;
  assign n18395 = n18389 & ~n18394;
  assign n18396 = ~n18369 & n18395;
  assign n18397 = ~n18333 & n18396;
  assign n18398 = ~n18330 & n18397;
  assign n18399 = ~pi394 & n18398;
  assign n18400 = pi394 & ~n18398;
  assign n18401 = ~n18399 & ~n18400;
  assign n18402 = pi139 & ~pi160;
  assign n18403 = ~pi139 & pi160;
  assign n18404 = ~n18402 & ~n18403;
  assign n18405 = pi162 & ~pi164;
  assign n18406 = ~pi162 & pi164;
  assign n18407 = ~n18405 & ~n18406;
  assign n18408 = ~n18404 & n18407;
  assign n18409 = n18404 & ~n18407;
  assign n18410 = ~n18408 & ~n18409;
  assign n18411 = n18401 & n18410;
  assign n18412 = ~n18401 & ~n18410;
  assign n18413 = ~n18411 & ~n18412;
  assign n18414 = ~pi532 & ~n18413;
  assign po274 = n18299 | n18414;
  assign n18416 = ~pi140 & ~pi141;
  assign n18417 = pi140 & pi141;
  assign n18418 = ~n18416 & ~n18417;
  assign n18419 = pi388 & n18418;
  assign n18420 = ~pi388 & ~n18418;
  assign n18421 = ~n18419 & ~n18420;
  assign n18422 = pi144 & n17766;
  assign n18423 = ~pi144 & ~n17766;
  assign n18424 = ~n18422 & ~n18423;
  assign n18425 = ~n18421 & n18424;
  assign n18426 = n18421 & ~n18424;
  assign n18427 = ~n18425 & ~n18426;
  assign n18428 = ~pi532 & ~n18427;
  assign n18429 = pi532 & pi594;
  assign po275 = n18428 | n18429;
  assign n18431 = pi141 & n17766;
  assign n18432 = ~pi141 & ~n17766;
  assign n18433 = ~n18431 & ~n18432;
  assign n18434 = pi388 & n18433;
  assign n18435 = ~pi388 & ~n18433;
  assign n18436 = ~n18434 & ~n18435;
  assign n18437 = ~pi532 & ~n18436;
  assign n18438 = pi532 & pi658;
  assign po276 = n18437 | n18438;
  assign n18440 = pi142 & ~pi167;
  assign n18441 = ~pi142 & pi167;
  assign n18442 = ~n18440 & ~n18441;
  assign n18443 = pi147 & ~pi166;
  assign n18444 = pi129 & n18443;
  assign n18445 = pi138 & n18444;
  assign n18446 = ~pi185 & n18443;
  assign n18447 = pi138 & n18446;
  assign n18448 = ~n18445 & ~n18447;
  assign n18449 = pi129 & ~pi166;
  assign n18450 = ~pi185 & n18449;
  assign n18451 = n18448 & ~n18450;
  assign n18452 = ~pi207 & ~n18451;
  assign n18453 = pi147 & pi166;
  assign n18454 = pi129 & n18453;
  assign n18455 = pi185 & n18454;
  assign n18456 = ~pi138 & n18455;
  assign n18457 = pi207 & n18456;
  assign n18458 = ~pi207 & pi302;
  assign n18459 = ~pi129 & ~pi147;
  assign n18460 = ~pi185 & n18459;
  assign n18461 = ~pi166 & pi185;
  assign n18462 = ~pi129 & n18461;
  assign n18463 = ~n18460 & ~n18462;
  assign n18464 = n18458 & ~n18463;
  assign n18465 = pi138 & ~pi207;
  assign n18466 = pi129 & pi302;
  assign n18467 = n18465 & n18466;
  assign n18468 = ~pi185 & n18467;
  assign n18469 = ~pi147 & pi166;
  assign n18470 = ~pi185 & n18469;
  assign n18471 = pi138 & n18470;
  assign n18472 = pi129 & n18469;
  assign n18473 = pi185 & n18472;
  assign n18474 = ~pi138 & n18473;
  assign n18475 = ~n18471 & ~n18474;
  assign n18476 = ~pi147 & ~pi166;
  assign n18477 = pi129 & n18476;
  assign n18478 = pi185 & n18477;
  assign n18479 = pi138 & n18478;
  assign n18480 = ~pi129 & n18476;
  assign n18481 = pi185 & n18480;
  assign n18482 = ~pi138 & n18481;
  assign n18483 = ~n18479 & ~n18482;
  assign n18484 = n18475 & n18483;
  assign n18485 = pi302 & ~n18484;
  assign n18486 = ~n18468 & ~n18485;
  assign n18487 = ~n18464 & n18486;
  assign n18488 = ~n18457 & n18487;
  assign n18489 = ~pi138 & pi207;
  assign n18490 = ~pi129 & n18443;
  assign n18491 = ~pi185 & n18490;
  assign n18492 = n18489 & n18491;
  assign n18493 = pi138 & pi185;
  assign n18494 = n18476 & n18493;
  assign n18495 = ~pi129 & pi147;
  assign n18496 = ~pi185 & n18495;
  assign n18497 = ~n18494 & ~n18496;
  assign n18498 = pi207 & ~n18497;
  assign n18499 = ~pi129 & n18469;
  assign n18500 = pi138 & n18499;
  assign n18501 = ~pi207 & n18500;
  assign n18502 = ~n18498 & ~n18501;
  assign n18503 = ~pi207 & n18444;
  assign n18504 = ~n18445 & ~n18456;
  assign n18505 = ~n18503 & n18504;
  assign n18506 = n18502 & n18505;
  assign n18507 = ~pi302 & ~n18506;
  assign n18508 = ~n18492 & ~n18507;
  assign n18509 = ~pi129 & n18453;
  assign n18510 = pi185 & n18509;
  assign n18511 = ~pi207 & n18510;
  assign n18512 = pi138 & ~pi185;
  assign n18513 = n18444 & n18512;
  assign n18514 = ~n18511 & ~n18513;
  assign n18515 = n18508 & n18514;
  assign n18516 = n18488 & n18515;
  assign n18517 = ~n18452 & n18516;
  assign n18518 = pi139 & ~n18517;
  assign n18519 = pi185 & n18444;
  assign n18520 = pi207 & n18519;
  assign n18521 = ~pi138 & n18509;
  assign n18522 = pi129 & pi166;
  assign n18523 = pi185 & n18522;
  assign n18524 = pi138 & n18523;
  assign n18525 = ~n18521 & ~n18524;
  assign n18526 = pi129 & ~pi147;
  assign n18527 = pi185 & n18526;
  assign n18528 = ~pi138 & n18527;
  assign n18529 = ~pi138 & n18446;
  assign n18530 = pi138 & n18469;
  assign n18531 = ~n18529 & ~n18530;
  assign n18532 = ~n18528 & n18531;
  assign n18533 = ~pi207 & ~n18532;
  assign n18534 = pi138 & pi207;
  assign n18535 = n18522 & n18534;
  assign n18536 = ~n18533 & ~n18535;
  assign n18537 = n18525 & n18536;
  assign n18538 = ~n18520 & n18537;
  assign n18539 = ~pi185 & n18444;
  assign n18540 = ~pi138 & n18539;
  assign n18541 = ~pi185 & n18472;
  assign n18542 = pi138 & n18480;
  assign n18543 = ~n18541 & ~n18542;
  assign n18544 = ~n18540 & n18543;
  assign n18545 = n18538 & n18544;
  assign n18546 = pi302 & ~n18545;
  assign n18547 = ~pi138 & ~pi185;
  assign n18548 = n18454 & n18547;
  assign n18549 = ~pi138 & n18480;
  assign n18550 = pi207 & n18549;
  assign n18551 = ~n18548 & ~n18550;
  assign n18552 = n18460 & n18534;
  assign n18553 = pi185 & n18499;
  assign n18554 = ~pi138 & n18553;
  assign n18555 = ~n18552 & ~n18554;
  assign n18556 = n18551 & n18555;
  assign n18557 = ~pi302 & ~n18556;
  assign n18558 = ~pi185 & n18476;
  assign n18559 = pi185 & n18490;
  assign n18560 = ~pi138 & n18559;
  assign n18561 = ~pi166 & ~pi185;
  assign n18562 = ~pi129 & n18561;
  assign n18563 = pi138 & n18562;
  assign n18564 = ~n18560 & ~n18563;
  assign n18565 = ~n18558 & n18564;
  assign n18566 = ~n18524 & n18565;
  assign n18567 = pi207 & ~n18566;
  assign n18568 = ~n18557 & ~n18567;
  assign n18569 = ~n18546 & n18568;
  assign n18570 = ~pi185 & n18453;
  assign n18571 = ~pi129 & n18570;
  assign n18572 = ~pi207 & n18571;
  assign n18573 = ~pi185 & n18480;
  assign n18574 = ~pi207 & n18473;
  assign n18575 = n18462 & n18465;
  assign n18576 = ~n18574 & ~n18575;
  assign n18577 = ~n18573 & n18576;
  assign n18578 = ~n18572 & n18577;
  assign n18579 = n18569 & n18578;
  assign n18580 = ~pi139 & ~n18579;
  assign n18581 = ~n18518 & ~n18580;
  assign n18582 = pi138 & n18573;
  assign n18583 = ~n18574 & ~n18582;
  assign n18584 = pi302 & ~n18583;
  assign n18585 = ~pi138 & ~pi207;
  assign n18586 = ~pi185 & n18522;
  assign n18587 = n18585 & n18586;
  assign n18588 = ~n18511 & ~n18587;
  assign n18589 = pi138 & n18519;
  assign n18590 = ~pi207 & n18589;
  assign n18591 = n18588 & ~n18590;
  assign n18592 = ~pi302 & ~n18591;
  assign n18593 = ~pi166 & n18547;
  assign n18594 = ~pi147 & n18593;
  assign n18595 = pi138 & n18527;
  assign n18596 = ~pi138 & pi185;
  assign n18597 = ~n18490 & ~n18499;
  assign n18598 = n18596 & ~n18597;
  assign n18599 = ~n18595 & ~n18598;
  assign n18600 = ~n18456 & n18599;
  assign n18601 = pi207 & ~n18600;
  assign n18602 = ~n18594 & ~n18601;
  assign n18603 = ~pi302 & ~n18602;
  assign n18604 = ~n18592 & ~n18603;
  assign n18605 = pi302 & n18519;
  assign n18606 = n18489 & n18605;
  assign n18607 = n18604 & ~n18606;
  assign n18608 = ~n18584 & n18607;
  assign n18609 = ~pi185 & n18477;
  assign n18610 = pi138 & n18609;
  assign n18611 = ~pi207 & n18610;
  assign n18612 = pi207 & n18479;
  assign n18613 = ~n18611 & ~n18612;
  assign n18614 = ~pi207 & n18521;
  assign n18615 = n18613 & ~n18614;
  assign n18616 = n18608 & n18615;
  assign n18617 = n18581 & n18616;
  assign n18618 = ~pi178 & n18617;
  assign n18619 = pi178 & ~n18617;
  assign n18620 = ~n18618 & ~n18619;
  assign n18621 = ~n18442 & n18620;
  assign n18622 = n18442 & ~n18620;
  assign n18623 = ~n18621 & ~n18622;
  assign n18624 = ~pi532 & ~n18623;
  assign n18625 = pi532 & pi570;
  assign po277 = n18624 | n18625;
  assign n18627 = ~pi143 & pi181;
  assign n18628 = pi143 & ~pi181;
  assign n18629 = ~n18627 & ~n18628;
  assign n18630 = pi207 & n18563;
  assign n18631 = ~pi129 & pi166;
  assign n18632 = ~pi185 & n18631;
  assign n18633 = ~pi138 & n18632;
  assign n18634 = pi185 & n18476;
  assign n18635 = pi207 & n18634;
  assign n18636 = ~n18453 & ~n18522;
  assign n18637 = n18489 & ~n18636;
  assign n18638 = ~n18635 & ~n18637;
  assign n18639 = pi138 & n18574;
  assign n18640 = n18638 & ~n18639;
  assign n18641 = ~n18481 & n18640;
  assign n18642 = ~n18633 & n18641;
  assign n18643 = ~pi302 & ~n18642;
  assign n18644 = ~pi185 & n18454;
  assign n18645 = pi207 & n18644;
  assign n18646 = pi138 & n18455;
  assign n18647 = ~n18500 & ~n18646;
  assign n18648 = n18444 & n18596;
  assign n18649 = ~n18562 & ~n18648;
  assign n18650 = pi207 & n18649;
  assign n18651 = ~pi207 & ~n18541;
  assign n18652 = ~n18650 & ~n18651;
  assign n18653 = n18647 & ~n18652;
  assign n18654 = ~n18548 & n18653;
  assign n18655 = pi302 & ~n18654;
  assign n18656 = ~n18645 & ~n18655;
  assign n18657 = pi185 & n18443;
  assign n18658 = pi138 & n18657;
  assign n18659 = ~n18456 & ~n18658;
  assign n18660 = ~pi207 & ~n18659;
  assign n18661 = ~pi138 & n18491;
  assign n18662 = ~n18660 & ~n18661;
  assign n18663 = n18656 & n18662;
  assign n18664 = ~n18643 & n18663;
  assign n18665 = ~n18630 & n18664;
  assign n18666 = ~pi139 & ~n18665;
  assign n18667 = ~pi138 & n18526;
  assign n18668 = ~n18472 & ~n18667;
  assign n18669 = pi185 & n18631;
  assign n18670 = n18668 & ~n18669;
  assign n18671 = pi207 & ~n18670;
  assign n18672 = ~pi207 & n18480;
  assign n18673 = pi138 & n18509;
  assign n18674 = ~n18473 & ~n18673;
  assign n18675 = ~n18672 & n18674;
  assign n18676 = ~n18671 & n18675;
  assign n18677 = ~pi138 & n18443;
  assign n18678 = ~pi207 & n18677;
  assign n18679 = ~pi138 & n18523;
  assign n18680 = ~n18678 & ~n18679;
  assign n18681 = n18676 & n18680;
  assign n18682 = pi302 & ~n18681;
  assign n18683 = ~pi207 & n18474;
  assign n18684 = pi138 & n18454;
  assign n18685 = ~n18633 & ~n18684;
  assign n18686 = ~pi207 & ~n18685;
  assign n18687 = ~n18683 & ~n18686;
  assign n18688 = pi138 & n18553;
  assign n18689 = pi207 & n18450;
  assign n18690 = pi207 & n18444;
  assign n18691 = n18465 & n18490;
  assign n18692 = n18499 & n18534;
  assign n18693 = ~n18691 & ~n18692;
  assign n18694 = ~n18690 & n18693;
  assign n18695 = ~n18689 & n18694;
  assign n18696 = ~n18614 & n18695;
  assign n18697 = pi129 & pi147;
  assign n18698 = ~pi185 & n18697;
  assign n18699 = ~pi138 & n18698;
  assign n18700 = n18696 & ~n18699;
  assign n18701 = ~n18594 & n18700;
  assign n18702 = ~n18688 & n18701;
  assign n18703 = ~pi302 & ~n18702;
  assign n18704 = ~n18513 & ~n18703;
  assign n18705 = n18687 & n18704;
  assign n18706 = ~n18682 & n18705;
  assign n18707 = pi185 & n18530;
  assign n18708 = ~n18559 & ~n18707;
  assign n18709 = ~n18553 & n18708;
  assign n18710 = pi207 & ~n18709;
  assign n18711 = n18706 & ~n18710;
  assign n18712 = pi139 & ~n18711;
  assign n18713 = ~n18666 & ~n18712;
  assign n18714 = pi207 & n18482;
  assign n18715 = ~n18492 & ~n18714;
  assign n18716 = ~pi302 & ~n18715;
  assign n18717 = n18713 & ~n18716;
  assign n18718 = pi138 & n18571;
  assign n18719 = pi207 & n18718;
  assign n18720 = pi207 & n18688;
  assign n18721 = pi207 & n18473;
  assign n18722 = pi185 & n18459;
  assign n18723 = ~n18446 & ~n18541;
  assign n18724 = ~n18722 & n18723;
  assign n18725 = n18585 & ~n18724;
  assign n18726 = ~n18721 & ~n18725;
  assign n18727 = ~pi185 & n18499;
  assign n18728 = pi138 & n18727;
  assign n18729 = ~pi207 & n18728;
  assign n18730 = n18534 & n18697;
  assign n18731 = ~pi185 & n18730;
  assign n18732 = pi207 & n18673;
  assign n18733 = ~n18731 & ~n18732;
  assign n18734 = ~n18729 & n18733;
  assign n18735 = n18726 & n18734;
  assign n18736 = pi302 & ~n18735;
  assign n18737 = ~pi207 & ~pi302;
  assign n18738 = pi138 & n18570;
  assign n18739 = n18737 & n18738;
  assign n18740 = ~n18736 & ~n18739;
  assign n18741 = pi138 & n18559;
  assign n18742 = n18740 & ~n18741;
  assign n18743 = ~n18720 & n18742;
  assign n18744 = ~n18719 & n18743;
  assign n18745 = n18717 & n18744;
  assign n18746 = pi180 & n18745;
  assign n18747 = ~pi180 & ~n18745;
  assign n18748 = ~n18746 & ~n18747;
  assign n18749 = ~n18629 & n18748;
  assign n18750 = n18629 & ~n18748;
  assign n18751 = ~n18749 & ~n18750;
  assign n18752 = ~pi532 & ~n18751;
  assign n18753 = pi532 & pi568;
  assign po278 = n18752 | n18753;
  assign n18755 = ~pi141 & pi144;
  assign n18756 = pi141 & ~pi144;
  assign n18757 = ~n18755 & ~n18756;
  assign n18758 = ~n17769 & n18757;
  assign n18759 = ~n17782 & ~n18757;
  assign po279 = n18758 | n18759;
  assign n18761 = ~pi132 & n17691;
  assign n18762 = ~pi351 & n18761;
  assign n18763 = ~n17648 & ~n18762;
  assign n18764 = ~n17641 & n18763;
  assign n18765 = ~n17643 & n18764;
  assign n18766 = pi132 & pi354;
  assign n18767 = pi358 & n18766;
  assign n18768 = ~n17598 & ~n18767;
  assign n18769 = pi351 & ~n18768;
  assign n18770 = n18765 & ~n18769;
  assign n18771 = ~pi284 & ~n18770;
  assign n18772 = ~pi157 & pi358;
  assign n18773 = ~n17658 & ~n18772;
  assign n18774 = n17733 & ~n18773;
  assign n18775 = n18346 & ~n18774;
  assign n18776 = ~n17633 & ~n17980;
  assign n18777 = n17620 & n18383;
  assign n18778 = n18776 & ~n18777;
  assign n18779 = pi351 & ~n18778;
  assign n18780 = n18775 & ~n18779;
  assign n18781 = pi284 & ~n18780;
  assign n18782 = ~n18771 & ~n18781;
  assign n18783 = ~n17679 & ~n17711;
  assign n18784 = ~n17642 & n18783;
  assign n18785 = ~n17981 & n18784;
  assign n18786 = pi351 & ~n18785;
  assign n18787 = ~n17614 & ~n17630;
  assign n18788 = ~pi351 & ~n18787;
  assign n18789 = ~n18786 & ~n18788;
  assign n18790 = n18782 & n18789;
  assign n18791 = pi193 & ~n18790;
  assign n18792 = pi284 & pi351;
  assign n18793 = pi132 & n17633;
  assign n18794 = ~n17743 & ~n18793;
  assign n18795 = ~n17694 & n18794;
  assign n18796 = n18792 & ~n18795;
  assign n18797 = pi284 & n17760;
  assign n18798 = n17621 & n17745;
  assign n18799 = ~n18325 & ~n18798;
  assign n18800 = pi351 & ~n18799;
  assign n18801 = ~pi132 & n18045;
  assign n18802 = pi358 & n18360;
  assign n18803 = ~n17707 & ~n17962;
  assign n18804 = n17722 & ~n18803;
  assign n18805 = ~n17999 & ~n18804;
  assign n18806 = ~n18802 & n18805;
  assign n18807 = ~n18801 & n18806;
  assign n18808 = ~pi351 & ~n18807;
  assign n18809 = ~n18800 & ~n18808;
  assign n18810 = pi132 & n17691;
  assign n18811 = pi351 & n18810;
  assign n18812 = pi132 & n17963;
  assign n18813 = ~n18811 & ~n18812;
  assign n18814 = ~pi132 & n17687;
  assign n18815 = ~pi351 & n18767;
  assign n18816 = ~n17630 & ~n18798;
  assign n18817 = ~n18815 & n18816;
  assign n18818 = ~n18814 & n18817;
  assign n18819 = n18813 & n18818;
  assign n18820 = ~pi284 & ~n18819;
  assign n18821 = n18809 & ~n18820;
  assign n18822 = ~pi351 & n17642;
  assign n18823 = ~n17737 & ~n18822;
  assign n18824 = n17602 & n17702;
  assign n18825 = pi351 & n18005;
  assign n18826 = ~n18824 & ~n18825;
  assign n18827 = n18823 & n18826;
  assign n18828 = pi284 & ~n18827;
  assign n18829 = n18821 & ~n18828;
  assign n18830 = ~pi193 & ~n18829;
  assign n18831 = ~n18797 & ~n18830;
  assign n18832 = ~n18796 & n18831;
  assign n18833 = ~n17960 & ~n18384;
  assign n18834 = pi132 & n17596;
  assign n18835 = pi351 & n18834;
  assign n18836 = pi132 & n17632;
  assign n18837 = ~pi351 & n18836;
  assign n18838 = ~n17644 & ~n18837;
  assign n18839 = ~pi351 & n17599;
  assign n18840 = n18838 & ~n18839;
  assign n18841 = ~n17968 & ~n18025;
  assign n18842 = ~n18034 & n18841;
  assign n18843 = n18840 & n18842;
  assign n18844 = ~n18835 & n18843;
  assign n18845 = ~pi284 & ~n18844;
  assign n18846 = pi351 & n18065;
  assign n18847 = ~n18845 & ~n18846;
  assign n18848 = ~n17656 & n18847;
  assign n18849 = n18833 & n18848;
  assign n18850 = n18832 & n18849;
  assign n18851 = ~n18791 & n18850;
  assign n18852 = pi145 & n18851;
  assign n18853 = ~pi145 & ~n18851;
  assign n18854 = ~n18852 & ~n18853;
  assign n18855 = pi391 & n18854;
  assign n18856 = ~pi391 & ~n18854;
  assign n18857 = ~n18855 & ~n18856;
  assign n18858 = ~pi532 & ~n18857;
  assign n18859 = pi532 & pi659;
  assign po282 = n18858 | n18859;
  assign n18861 = ~pi145 & ~pi146;
  assign n18862 = pi145 & pi146;
  assign n18863 = ~n18861 & ~n18862;
  assign n18864 = pi391 & n18851;
  assign n18865 = ~pi391 & ~n18851;
  assign n18866 = ~n18864 & ~n18865;
  assign n18867 = ~n18863 & n18866;
  assign n18868 = n18863 & ~n18866;
  assign n18869 = ~n18867 & ~n18868;
  assign n18870 = ~pi532 & ~n18869;
  assign n18871 = pi532 & pi627;
  assign po283 = n18870 | n18871;
  assign n18873 = ~pi146 & ~pi153;
  assign n18874 = pi146 & pi153;
  assign n18875 = ~n18873 & ~n18874;
  assign n18876 = ~pi145 & pi147;
  assign n18877 = pi145 & ~pi147;
  assign n18878 = ~n18876 & ~n18877;
  assign n18879 = ~n18875 & n18878;
  assign n18880 = n18875 & ~n18878;
  assign n18881 = ~n18879 & ~n18880;
  assign n18882 = n18866 & ~n18881;
  assign n18883 = ~n18866 & n18881;
  assign n18884 = ~n18882 & ~n18883;
  assign n18885 = ~pi532 & ~n18884;
  assign n18886 = pi532 & pi563;
  assign po284 = n18885 | n18886;
  assign n18888 = pi148 & n17944;
  assign n18889 = ~pi148 & ~n17944;
  assign n18890 = ~n18888 & ~n18889;
  assign n18891 = ~pi532 & ~n18890;
  assign n18892 = pi532 & pi650;
  assign po285 = n18891 | n18892;
  assign n18894 = ~pi148 & ~pi149;
  assign n18895 = pi148 & pi149;
  assign n18896 = ~n18894 & ~n18895;
  assign n18897 = n17944 & ~n18896;
  assign n18898 = ~n17944 & n18896;
  assign n18899 = ~n18897 & ~n18898;
  assign n18900 = ~pi532 & ~n18899;
  assign n18901 = pi532 & pi618;
  assign po286 = n18900 | n18901;
  assign n18903 = pi150 & ~pi187;
  assign n18904 = ~pi150 & pi187;
  assign n18905 = ~n18903 & ~n18904;
  assign n18906 = ~pi207 & n18513;
  assign n18907 = ~pi138 & n18490;
  assign n18908 = ~pi138 & n18609;
  assign n18909 = ~n18907 & ~n18908;
  assign n18910 = ~pi138 & n18657;
  assign n18911 = n18909 & ~n18910;
  assign n18912 = ~pi207 & ~n18911;
  assign n18913 = ~n18906 & ~n18912;
  assign n18914 = ~n18612 & n18913;
  assign n18915 = ~pi302 & ~n18914;
  assign n18916 = pi207 & n18560;
  assign n18917 = ~pi207 & n18679;
  assign n18918 = ~n18916 & ~n18917;
  assign n18919 = ~pi129 & n18547;
  assign n18920 = n18476 & n18919;
  assign n18921 = ~n18610 & ~n18920;
  assign n18922 = ~n18692 & n18921;
  assign n18923 = n18918 & n18922;
  assign n18924 = pi302 & ~n18923;
  assign n18925 = ~n18915 & ~n18924;
  assign n18926 = ~pi138 & n18727;
  assign n18927 = pi207 & n18926;
  assign n18928 = pi207 & n18699;
  assign n18929 = ~n18927 & ~n18928;
  assign n18930 = ~pi302 & ~n18929;
  assign n18931 = pi207 & ~n18540;
  assign n18932 = n18453 & n18493;
  assign n18933 = ~pi207 & ~n18932;
  assign n18934 = ~n18931 & ~n18933;
  assign n18935 = ~n18519 & ~n18549;
  assign n18936 = ~n18510 & n18935;
  assign n18937 = pi207 & ~n18936;
  assign n18938 = n18553 & n18585;
  assign n18939 = ~n18937 & ~n18938;
  assign n18940 = ~pi129 & n18512;
  assign n18941 = ~n18471 & ~n18940;
  assign n18942 = ~pi138 & n18450;
  assign n18943 = n18941 & ~n18942;
  assign n18944 = n18939 & n18943;
  assign n18945 = ~pi302 & ~n18944;
  assign n18946 = pi138 & ~pi166;
  assign n18947 = ~pi185 & n18946;
  assign n18948 = pi138 & n18495;
  assign n18949 = ~n18947 & ~n18948;
  assign n18950 = ~pi207 & ~n18949;
  assign n18951 = n18449 & n18596;
  assign n18952 = ~n18455 & ~n18951;
  assign n18953 = ~pi207 & ~n18952;
  assign n18954 = pi138 & n18586;
  assign n18955 = ~n18479 & ~n18954;
  assign n18956 = ~n18474 & n18955;
  assign n18957 = ~n18727 & n18956;
  assign n18958 = pi207 & ~n18957;
  assign n18959 = ~n18953 & ~n18958;
  assign n18960 = ~n18950 & n18959;
  assign n18961 = ~pi138 & n18444;
  assign n18962 = ~n18728 & ~n18961;
  assign n18963 = ~pi207 & n18697;
  assign n18964 = ~n18672 & ~n18963;
  assign n18965 = ~n18559 & n18964;
  assign n18966 = pi302 & ~n18965;
  assign n18967 = n18962 & ~n18966;
  assign n18968 = n18960 & n18967;
  assign n18969 = ~n18945 & n18968;
  assign n18970 = pi139 & ~n18969;
  assign n18971 = pi207 & ~pi302;
  assign n18972 = n18472 & n18971;
  assign n18973 = ~n18477 & ~n18495;
  assign n18974 = n18534 & ~n18973;
  assign n18975 = ~pi185 & n18974;
  assign n18976 = ~n18972 & ~n18975;
  assign n18977 = ~pi207 & n18494;
  assign n18978 = ~n18491 & ~n18644;
  assign n18979 = ~pi138 & ~n18978;
  assign n18980 = ~n18977 & ~n18979;
  assign n18981 = ~pi302 & ~n18980;
  assign n18982 = ~pi302 & n18522;
  assign n18983 = n18489 & n18982;
  assign n18984 = ~n18981 & ~n18983;
  assign n18985 = ~pi138 & n18460;
  assign n18986 = ~n18474 & ~n18985;
  assign n18987 = ~n18684 & n18986;
  assign n18988 = ~pi207 & ~n18987;
  assign n18989 = ~pi138 & n18476;
  assign n18990 = pi207 & n18445;
  assign n18991 = n18585 & n18631;
  assign n18992 = ~n18990 & ~n18991;
  assign n18993 = ~n18932 & n18992;
  assign n18994 = ~n18989 & n18993;
  assign n18995 = ~n18558 & n18994;
  assign n18996 = pi302 & ~n18995;
  assign n18997 = ~n18988 & ~n18996;
  assign n18998 = n18984 & n18997;
  assign n18999 = n18976 & n18998;
  assign n19000 = ~pi139 & ~n18999;
  assign n19001 = ~n18970 & ~n19000;
  assign n19002 = ~n18934 & n19001;
  assign n19003 = ~n18930 & n19002;
  assign n19004 = n18925 & n19003;
  assign n19005 = ~pi190 & n19004;
  assign n19006 = pi190 & ~n19004;
  assign n19007 = ~n19005 & ~n19006;
  assign n19008 = ~n18905 & n19007;
  assign n19009 = n18905 & ~n19007;
  assign n19010 = ~n19008 & ~n19009;
  assign n19011 = ~pi532 & ~n19010;
  assign n19012 = pi532 & pi565;
  assign po287 = n19011 | n19012;
  assign n19014 = pi151 & ~pi222;
  assign n19015 = ~pi151 & pi222;
  assign n19016 = ~n19014 & ~n19015;
  assign n19017 = pi321 & n18185;
  assign n19018 = pi342 & n18215;
  assign n19019 = ~n19017 & ~n19018;
  assign n19020 = pi352 & pi372;
  assign n19021 = ~n19019 & n19020;
  assign n19022 = ~pi352 & n18163;
  assign n19023 = n18127 & n18153;
  assign n19024 = ~n18242 & ~n19023;
  assign n19025 = ~pi352 & ~n19024;
  assign n19026 = ~n19022 & ~n19025;
  assign n19027 = ~n18208 & n19026;
  assign n19028 = pi372 & ~n19027;
  assign n19029 = pi372 & n18198;
  assign n19030 = n18138 & n19029;
  assign n19031 = ~n19028 & ~n19030;
  assign n19032 = pi170 & n18116;
  assign n19033 = ~n18113 & ~n19032;
  assign n19034 = n18119 & ~n19033;
  assign n19035 = ~pi321 & n19034;
  assign n19036 = ~n18257 & ~n19035;
  assign n19037 = ~pi352 & n18211;
  assign n19038 = pi352 & n18178;
  assign n19039 = ~n18197 & ~n19038;
  assign n19040 = ~pi321 & n18127;
  assign n19041 = pi352 & n19040;
  assign n19042 = n19039 & ~n19041;
  assign n19043 = ~pi352 & n19017;
  assign n19044 = ~n18267 & ~n19043;
  assign n19045 = n19042 & n19044;
  assign n19046 = ~n19037 & n19045;
  assign n19047 = ~pi182 & n19032;
  assign n19048 = ~pi182 & n18201;
  assign n19049 = ~n19047 & ~n19048;
  assign n19050 = n19046 & n19049;
  assign n19051 = ~pi372 & ~n19050;
  assign n19052 = ~pi352 & pi372;
  assign n19053 = pi276 & n18153;
  assign n19054 = ~n18248 & ~n19053;
  assign n19055 = n19052 & ~n19054;
  assign n19056 = n18191 & n18205;
  assign n19057 = pi352 & n18210;
  assign n19058 = ~n19056 & ~n19057;
  assign n19059 = pi372 & ~n19058;
  assign n19060 = ~n19055 & ~n19059;
  assign n19061 = ~n19051 & n19060;
  assign n19062 = ~pi182 & n18152;
  assign n19063 = pi352 & n19062;
  assign n19064 = ~pi321 & n19032;
  assign n19065 = ~pi182 & n19064;
  assign n19066 = pi321 & n19032;
  assign n19067 = ~n18227 & ~n19066;
  assign n19068 = ~n18143 & n19067;
  assign n19069 = n18198 & ~n19068;
  assign n19070 = ~n19065 & ~n19069;
  assign n19071 = ~pi182 & n18255;
  assign n19072 = n19070 & ~n19071;
  assign n19073 = ~n19063 & n19072;
  assign n19074 = n19061 & n19073;
  assign n19075 = pi191 & ~n19074;
  assign n19076 = n18200 & n18205;
  assign n19077 = ~n18182 & ~n19076;
  assign n19078 = ~pi372 & ~n19077;
  assign n19079 = pi182 & n19064;
  assign n19080 = ~pi352 & n19079;
  assign n19081 = ~n18129 & ~n19080;
  assign n19082 = pi182 & n19017;
  assign n19083 = pi352 & n19082;
  assign n19084 = pi182 & n18128;
  assign n19085 = ~pi182 & n18116;
  assign n19086 = pi182 & n18249;
  assign n19087 = ~n19085 & ~n19086;
  assign n19088 = pi352 & ~n19087;
  assign n19089 = pi182 & n18136;
  assign n19090 = pi182 & n18120;
  assign n19091 = ~n19089 & ~n19090;
  assign n19092 = ~n18110 & n19091;
  assign n19093 = ~pi352 & ~n19092;
  assign n19094 = ~n19088 & ~n19093;
  assign n19095 = ~n19084 & n19094;
  assign n19096 = pi372 & ~n19095;
  assign n19097 = ~n19083 & ~n19096;
  assign n19098 = n19081 & n19097;
  assign n19099 = ~n19078 & n19098;
  assign n19100 = ~pi191 & ~n19099;
  assign n19101 = ~n19075 & ~n19100;
  assign n19102 = pi182 & pi321;
  assign n19103 = pi170 & n19102;
  assign n19104 = n18140 & n19103;
  assign n19105 = ~n19064 & ~n19104;
  assign n19106 = ~n18229 & n19105;
  assign n19107 = ~pi352 & ~n19106;
  assign n19108 = pi182 & n18248;
  assign n19109 = ~n19107 & ~n19108;
  assign n19110 = ~pi352 & n19047;
  assign n19111 = pi352 & n18182;
  assign n19112 = ~n18255 & ~n19111;
  assign n19113 = pi182 & n18149;
  assign n19114 = pi182 & n18247;
  assign n19115 = ~n19113 & ~n19114;
  assign n19116 = pi352 & ~n19115;
  assign n19117 = n19112 & ~n19116;
  assign n19118 = ~n19110 & n19117;
  assign n19119 = n19109 & n19118;
  assign n19120 = ~pi372 & ~n19119;
  assign n19121 = n19101 & ~n19120;
  assign n19122 = n19036 & n19121;
  assign n19123 = n19031 & n19122;
  assign n19124 = ~n19021 & n19123;
  assign n19125 = pi229 & n19124;
  assign n19126 = ~pi229 & ~n19124;
  assign n19127 = ~n19125 & ~n19126;
  assign n19128 = ~n19016 & n19127;
  assign n19129 = n19016 & ~n19127;
  assign n19130 = ~n19128 & ~n19129;
  assign n19131 = ~pi532 & ~n19130;
  assign n19132 = pi532 & pi575;
  assign po288 = n19131 | n19132;
  assign n19134 = ~pi152 & pi256;
  assign n19135 = pi152 & ~pi256;
  assign n19136 = ~n19134 & ~n19135;
  assign n19137 = pi182 & n18210;
  assign n19138 = pi352 & n19137;
  assign n19139 = ~pi352 & n18227;
  assign n19140 = ~pi352 & n19084;
  assign n19141 = ~n19139 & ~n19140;
  assign n19142 = ~n18130 & n19141;
  assign n19143 = ~n19138 & n19142;
  assign n19144 = ~n18217 & ~n18229;
  assign n19145 = ~n18150 & n19144;
  assign n19146 = n19143 & n19145;
  assign n19147 = ~pi372 & ~n19146;
  assign n19148 = pi352 & n18245;
  assign n19149 = ~n19147 & ~n19148;
  assign n19150 = ~pi170 & ~pi182;
  assign n19151 = ~pi276 & n19150;
  assign n19152 = ~pi342 & n19151;
  assign n19153 = pi352 & n19152;
  assign n19154 = n19149 & ~n19153;
  assign n19155 = ~pi170 & n18215;
  assign n19156 = n18116 & n19155;
  assign n19157 = ~n18131 & ~n19156;
  assign n19158 = n18153 & n18185;
  assign n19159 = ~pi321 & n18247;
  assign n19160 = ~pi182 & n19159;
  assign n19161 = ~n19158 & ~n19160;
  assign n19162 = pi352 & ~n19161;
  assign n19163 = ~pi182 & n18248;
  assign n19164 = pi321 & n19062;
  assign n19165 = ~n19163 & ~n19164;
  assign n19166 = pi182 & ~pi321;
  assign n19167 = ~n18113 & ~n18136;
  assign n19168 = n19166 & ~n19167;
  assign n19169 = n19165 & ~n19168;
  assign n19170 = ~n18186 & n19169;
  assign n19171 = ~pi352 & ~n19170;
  assign n19172 = ~pi321 & n18117;
  assign n19173 = ~pi352 & n19172;
  assign n19174 = ~n19104 & ~n19173;
  assign n19175 = pi372 & ~n19174;
  assign n19176 = n18110 & n18119;
  assign n19177 = ~n19111 & ~n19176;
  assign n19178 = pi372 & ~n19177;
  assign n19179 = ~n19175 & ~n19178;
  assign n19180 = ~n18191 & ~n19158;
  assign n19181 = pi342 & n19102;
  assign n19182 = ~pi352 & n19181;
  assign n19183 = ~pi182 & n19040;
  assign n19184 = ~n19182 & ~n19183;
  assign n19185 = pi182 & n19032;
  assign n19186 = pi352 & n19185;
  assign n19187 = pi182 & n18114;
  assign n19188 = ~n19186 & ~n19187;
  assign n19189 = n19184 & n19188;
  assign n19190 = n19180 & n19189;
  assign n19191 = ~pi372 & ~n19190;
  assign n19192 = n19179 & ~n19191;
  assign n19193 = ~n19171 & n19192;
  assign n19194 = ~n19162 & n19193;
  assign n19195 = ~pi191 & ~n19194;
  assign n19196 = pi372 & n19080;
  assign n19197 = ~n19195 & ~n19196;
  assign n19198 = pi182 & n18157;
  assign n19199 = ~n18118 & ~n19198;
  assign n19200 = ~n18211 & n19199;
  assign n19201 = n19020 & ~n19200;
  assign n19202 = n19197 & ~n19201;
  assign n19203 = pi182 & n19066;
  assign n19204 = ~pi321 & n18121;
  assign n19205 = pi182 & n19204;
  assign n19206 = ~n19203 & ~n19205;
  assign n19207 = ~pi170 & pi321;
  assign n19208 = ~n18247 & ~n19207;
  assign n19209 = n18252 & ~n19208;
  assign n19210 = n19206 & ~n19209;
  assign n19211 = ~pi182 & n18242;
  assign n19212 = ~n18141 & ~n19211;
  assign n19213 = ~n18157 & n19212;
  assign n19214 = pi352 & ~n19213;
  assign n19215 = n19210 & ~n19214;
  assign n19216 = pi372 & ~n19215;
  assign n19217 = ~n18137 & ~n19181;
  assign n19218 = pi352 & ~n19217;
  assign n19219 = ~pi352 & n18242;
  assign n19220 = pi321 & n18109;
  assign n19221 = n18205 & n19220;
  assign n19222 = ~n19219 & ~n19221;
  assign n19223 = ~n19218 & n19222;
  assign n19224 = ~n18129 & n19223;
  assign n19225 = ~n19110 & n19224;
  assign n19226 = ~pi372 & ~n19225;
  assign n19227 = ~n19216 & ~n19226;
  assign n19228 = ~n18142 & ~n18162;
  assign n19229 = ~n19172 & n19228;
  assign n19230 = ~n18145 & n19229;
  assign n19231 = pi352 & ~n19230;
  assign n19232 = pi321 & n18173;
  assign n19233 = ~pi182 & n19232;
  assign n19234 = ~n18191 & ~n19233;
  assign n19235 = ~pi352 & ~n19234;
  assign n19236 = ~n19231 & ~n19235;
  assign n19237 = n19227 & n19236;
  assign n19238 = pi191 & ~n19237;
  assign n19239 = n19202 & ~n19238;
  assign n19240 = n19157 & n19239;
  assign n19241 = n19154 & n19240;
  assign n19242 = pi227 & n19241;
  assign n19243 = ~pi227 & ~n19241;
  assign n19244 = ~n19242 & ~n19243;
  assign n19245 = ~n19136 & n19244;
  assign n19246 = n19136 & ~n19244;
  assign n19247 = ~n19245 & ~n19246;
  assign n19248 = ~pi532 & ~n19247;
  assign n19249 = pi532 & pi579;
  assign po289 = n19248 | n19249;
  assign n19251 = ~pi145 & pi153;
  assign n19252 = pi145 & ~pi153;
  assign n19253 = ~n19251 & ~n19252;
  assign n19254 = pi391 & n19253;
  assign n19255 = ~pi391 & ~n19253;
  assign n19256 = ~n19254 & ~n19255;
  assign n19257 = ~pi146 & n18851;
  assign n19258 = pi146 & ~n18851;
  assign n19259 = ~n19257 & ~n19258;
  assign n19260 = ~n19256 & n19259;
  assign n19261 = n19256 & ~n19259;
  assign n19262 = ~n19260 & ~n19261;
  assign n19263 = ~pi532 & ~n19262;
  assign n19264 = pi532 & pi595;
  assign po290 = n19263 | n19264;
  assign n19266 = pi154 & ~pi189;
  assign n19267 = ~pi154 & pi189;
  assign n19268 = ~n19266 & ~n19267;
  assign n19269 = ~pi231 & n17383;
  assign n19270 = ~pi175 & n17937;
  assign n19271 = ~pi175 & n17366;
  assign n19272 = ~pi175 & n17318;
  assign n19273 = ~n19271 & ~n19272;
  assign n19274 = ~n19270 & n19273;
  assign n19275 = ~pi231 & ~n19274;
  assign n19276 = ~n19269 & ~n19275;
  assign n19277 = ~n17940 & n19276;
  assign n19278 = ~pi285 & ~n19277;
  assign n19279 = pi231 & n17898;
  assign n19280 = ~pi231 & n17397;
  assign n19281 = ~n19279 & ~n19280;
  assign n19282 = ~pi232 & n17405;
  assign n19283 = n17313 & n19282;
  assign n19284 = ~n17938 & ~n19283;
  assign n19285 = ~n17414 & n19284;
  assign n19286 = n19281 & n19285;
  assign n19287 = pi285 & ~n19286;
  assign n19288 = ~n19278 & ~n19287;
  assign n19289 = ~pi175 & n17293;
  assign n19290 = pi231 & n19289;
  assign n19291 = pi231 & n17422;
  assign n19292 = ~n19290 & ~n19291;
  assign n19293 = ~pi285 & ~n19292;
  assign n19294 = n19288 & ~n19293;
  assign n19295 = pi231 & ~n17888;
  assign n19296 = n17300 & n17847;
  assign n19297 = ~pi231 & ~n19296;
  assign n19298 = ~n19295 & ~n19297;
  assign n19299 = ~n17868 & ~n17884;
  assign n19300 = ~n17861 & n19299;
  assign n19301 = pi231 & ~n19300;
  assign n19302 = n17289 & n17403;
  assign n19303 = ~n19301 & ~n19302;
  assign n19304 = ~pi232 & n17382;
  assign n19305 = ~n17839 & ~n19304;
  assign n19306 = ~pi175 & n17409;
  assign n19307 = n19305 & ~n19306;
  assign n19308 = n19303 & n19307;
  assign n19309 = ~pi285 & ~n19308;
  assign n19310 = n17351 & n17408;
  assign n19311 = ~n17356 & ~n19310;
  assign n19312 = ~pi231 & ~n19311;
  assign n19313 = pi175 & n17914;
  assign n19314 = ~n17837 & ~n19313;
  assign n19315 = ~n17376 & n19314;
  assign n19316 = ~n17293 & n19315;
  assign n19317 = pi231 & ~n19316;
  assign n19318 = ~n19312 & ~n19317;
  assign n19319 = pi175 & ~pi233;
  assign n19320 = ~pi270 & n19319;
  assign n19321 = pi175 & n17849;
  assign n19322 = ~n19320 & ~n19321;
  assign n19323 = ~pi231 & ~n19322;
  assign n19324 = n19318 & ~n19323;
  assign n19325 = ~pi175 & n17350;
  assign n19326 = ~n17294 & ~n19325;
  assign n19327 = ~pi231 & n17297;
  assign n19328 = ~n17390 & ~n19327;
  assign n19329 = ~n17430 & n19328;
  assign n19330 = pi285 & ~n19329;
  assign n19331 = n19326 & ~n19330;
  assign n19332 = n19324 & n19331;
  assign n19333 = ~n19309 & n19332;
  assign n19334 = pi234 & ~n19333;
  assign n19335 = pi231 & ~pi285;
  assign n19336 = n17279 & n19335;
  assign n19337 = ~n17835 & ~n17849;
  assign n19338 = n17296 & ~n19337;
  assign n19339 = ~pi270 & n19338;
  assign n19340 = ~n19336 & ~n19339;
  assign n19341 = ~pi231 & n17848;
  assign n19342 = ~n17319 & ~n17347;
  assign n19343 = ~pi175 & ~n19342;
  assign n19344 = ~n19341 & ~n19343;
  assign n19345 = ~pi285 & ~n19344;
  assign n19346 = ~pi175 & n19335;
  assign n19347 = n17336 & n19346;
  assign n19348 = ~n19345 & ~n19347;
  assign n19349 = ~pi175 & n17827;
  assign n19350 = ~n17376 & ~n19349;
  assign n19351 = ~n17378 & n19350;
  assign n19352 = ~pi231 & ~n19351;
  assign n19353 = ~pi175 & n17313;
  assign n19354 = pi231 & n17820;
  assign n19355 = n17289 & n17331;
  assign n19356 = ~n19354 & ~n19355;
  assign n19357 = ~n19296 & n19356;
  assign n19358 = ~n19353 & n19357;
  assign n19359 = ~n17897 & n19358;
  assign n19360 = pi285 & ~n19359;
  assign n19361 = ~n19352 & ~n19360;
  assign n19362 = n19348 & n19361;
  assign n19363 = n19340 & n19362;
  assign n19364 = ~pi234 & ~n19363;
  assign n19365 = ~n19334 & ~n19364;
  assign n19366 = ~n19298 & n19365;
  assign n19367 = n19294 & n19366;
  assign n19368 = ~pi192 & n19367;
  assign n19369 = pi192 & ~n19367;
  assign n19370 = ~n19368 & ~n19369;
  assign n19371 = ~n19268 & n19370;
  assign n19372 = n19268 & ~n19370;
  assign n19373 = ~n19371 & ~n19372;
  assign n19374 = ~pi532 & ~n19373;
  assign n19375 = pi532 & pi581;
  assign po291 = n19374 | n19375;
  assign n19377 = ~pi155 & pi225;
  assign n19378 = pi155 & ~pi225;
  assign n19379 = ~n19377 & ~n19378;
  assign n19380 = pi352 & ~pi372;
  assign n19381 = n18128 & n19380;
  assign n19382 = ~n18138 & ~n18149;
  assign n19383 = ~pi182 & ~n19382;
  assign n19384 = n18116 & n19102;
  assign n19385 = ~pi352 & n19384;
  assign n19386 = ~n19383 & ~n19385;
  assign n19387 = ~pi372 & ~n19386;
  assign n19388 = ~pi372 & n18121;
  assign n19389 = n18119 & n19388;
  assign n19390 = ~n19387 & ~n19389;
  assign n19391 = pi321 & n19090;
  assign n19392 = pi182 & n18152;
  assign n19393 = pi352 & n19392;
  assign n19394 = n18113 & n18252;
  assign n19395 = ~n19393 & ~n19394;
  assign n19396 = ~n19085 & n19395;
  assign n19397 = ~n18210 & n19396;
  assign n19398 = ~n19391 & n19397;
  assign n19399 = pi372 & ~n19398;
  assign n19400 = ~n18136 & ~n19032;
  assign n19401 = n18198 & ~n19400;
  assign n19402 = ~pi321 & n19401;
  assign n19403 = ~n19399 & ~n19402;
  assign n19404 = n19390 & n19403;
  assign n19405 = ~n19381 & n19404;
  assign n19406 = ~n18193 & ~n18222;
  assign n19407 = ~n19160 & n19406;
  assign n19408 = ~pi352 & ~n19407;
  assign n19409 = n19405 & ~n19408;
  assign n19410 = ~pi191 & ~n19409;
  assign n19411 = ~pi182 & n18191;
  assign n19412 = pi352 & ~n19411;
  assign n19413 = ~pi352 & ~n19391;
  assign n19414 = ~n19412 & ~n19413;
  assign n19415 = ~pi170 & n19166;
  assign n19416 = pi182 & n19040;
  assign n19417 = ~n19415 & ~n19416;
  assign n19418 = ~n19048 & n19417;
  assign n19419 = n18212 & n18252;
  assign n19420 = ~n19017 & ~n19152;
  assign n19421 = pi321 & n18152;
  assign n19422 = n19420 & ~n19421;
  assign n19423 = pi352 & ~n19422;
  assign n19424 = ~n19419 & ~n19423;
  assign n19425 = n19418 & n19424;
  assign n19426 = ~pi372 & ~n19425;
  assign n19427 = ~pi342 & n19166;
  assign n19428 = ~n19089 & ~n19427;
  assign n19429 = ~pi352 & ~n19428;
  assign n19430 = ~n19426 & ~n19429;
  assign n19431 = n18153 & n18200;
  assign n19432 = ~n18144 & ~n19431;
  assign n19433 = ~pi352 & ~n19432;
  assign n19434 = ~n18255 & n19206;
  assign n19435 = ~n18222 & n19434;
  assign n19436 = pi352 & ~n19435;
  assign n19437 = ~n19433 & ~n19436;
  assign n19438 = ~n18256 & ~n19062;
  assign n19439 = ~pi352 & n18216;
  assign n19440 = ~n18227 & ~n19439;
  assign n19441 = ~n18183 & n19440;
  assign n19442 = pi372 & ~n19441;
  assign n19443 = n19438 & ~n19442;
  assign n19444 = n19437 & n19443;
  assign n19445 = n19430 & n19444;
  assign n19446 = pi191 & ~n19445;
  assign n19447 = ~pi182 & n18137;
  assign n19448 = ~pi182 & n18141;
  assign n19449 = ~n19447 & ~n19448;
  assign n19450 = ~n19065 & n19449;
  assign n19451 = ~pi352 & ~n19450;
  assign n19452 = ~n19056 & ~n19451;
  assign n19453 = pi352 & n19203;
  assign n19454 = n19452 & ~n19453;
  assign n19455 = ~pi372 & ~n19454;
  assign n19456 = ~pi182 & n18227;
  assign n19457 = pi352 & ~n19456;
  assign n19458 = ~pi352 & ~n18182;
  assign n19459 = ~n19457 & ~n19458;
  assign n19460 = ~n19079 & ~n19156;
  assign n19461 = ~n18199 & n19460;
  assign n19462 = ~n19459 & n19461;
  assign n19463 = pi372 & ~n19462;
  assign n19464 = ~n19455 & ~n19463;
  assign n19465 = pi352 & n18217;
  assign n19466 = pi352 & n19071;
  assign n19467 = ~n19465 & ~n19466;
  assign n19468 = ~pi372 & ~n19467;
  assign n19469 = n19464 & ~n19468;
  assign n19470 = ~n19446 & n19469;
  assign n19471 = ~n19414 & n19470;
  assign n19472 = ~n19410 & n19471;
  assign n19473 = pi230 & n19472;
  assign n19474 = ~pi230 & ~n19472;
  assign n19475 = ~n19473 & ~n19474;
  assign n19476 = ~n19379 & n19475;
  assign n19477 = n19379 & ~n19475;
  assign n19478 = ~n19476 & ~n19477;
  assign n19479 = ~pi532 & ~n19478;
  assign n19480 = pi532 & pi573;
  assign po292 = n19479 | n19480;
  assign n19482 = ~pi156 & pi224;
  assign n19483 = pi156 & ~pi224;
  assign n19484 = ~n19482 & ~n19483;
  assign n19485 = ~n18248 & ~n19085;
  assign n19486 = pi182 & n18140;
  assign n19487 = pi276 & ~pi321;
  assign n19488 = ~n19486 & ~n19487;
  assign n19489 = n19485 & n19488;
  assign n19490 = n19020 & ~n19489;
  assign n19491 = n18161 & n18252;
  assign n19492 = ~n19082 & ~n19491;
  assign n19493 = pi372 & ~n19492;
  assign n19494 = ~n19490 & ~n19493;
  assign n19495 = ~pi352 & n18152;
  assign n19496 = pi321 & n18216;
  assign n19497 = ~n18141 & ~n18248;
  assign n19498 = ~n19496 & n19497;
  assign n19499 = ~pi352 & ~n19498;
  assign n19500 = ~n19495 & ~n19499;
  assign n19501 = ~pi321 & n18173;
  assign n19502 = pi182 & n19501;
  assign n19503 = ~n19448 & ~n19502;
  assign n19504 = pi352 & n18115;
  assign n19505 = n19503 & ~n19504;
  assign n19506 = ~n18179 & n19505;
  assign n19507 = n19500 & n19506;
  assign n19508 = ~pi372 & ~n19507;
  assign n19509 = ~pi352 & n19448;
  assign n19510 = ~n19508 & ~n19509;
  assign n19511 = ~pi182 & n18266;
  assign n19512 = ~n19233 & ~n19511;
  assign n19513 = pi352 & ~n19512;
  assign n19514 = ~pi321 & n18136;
  assign n19515 = n18198 & n19514;
  assign n19516 = ~n19513 & ~n19515;
  assign n19517 = pi352 & n19421;
  assign n19518 = n19516 & ~n19517;
  assign n19519 = ~n19431 & n19518;
  assign n19520 = n19510 & n19519;
  assign n19521 = n19494 & n19520;
  assign n19522 = pi191 & n19521;
  assign n19523 = ~pi182 & n18143;
  assign n19524 = ~n19048 & ~n19523;
  assign n19525 = ~pi352 & ~n19524;
  assign n19526 = ~pi321 & pi342;
  assign n19527 = n18265 & n19526;
  assign n19528 = ~n19525 & ~n19527;
  assign n19529 = pi352 & n18163;
  assign n19530 = ~pi372 & n19205;
  assign n19531 = n18198 & n19172;
  assign n19532 = ~n19530 & ~n19531;
  assign n19533 = ~n19453 & n19532;
  assign n19534 = ~n19529 & n19533;
  assign n19535 = n18172 & n18198;
  assign n19536 = pi352 & n18117;
  assign n19537 = ~n19535 & ~n19536;
  assign n19538 = ~pi372 & ~n19537;
  assign n19539 = n19534 & ~n19538;
  assign n19540 = ~pi352 & n19104;
  assign n19541 = ~pi352 & n18118;
  assign n19542 = ~n19540 & ~n19541;
  assign n19543 = pi182 & n18137;
  assign n19544 = pi182 & ~pi276;
  assign n19545 = pi321 & n19544;
  assign n19546 = ~n19543 & ~n19545;
  assign n19547 = ~pi352 & ~n19546;
  assign n19548 = pi321 & n18136;
  assign n19549 = n18119 & n19548;
  assign n19550 = ~n19547 & ~n19549;
  assign n19551 = ~n19158 & n19550;
  assign n19552 = ~n19084 & n19551;
  assign n19553 = pi372 & ~n19552;
  assign n19554 = n19542 & ~n19553;
  assign n19555 = n19539 & n19554;
  assign n19556 = n19528 & n19555;
  assign n19557 = ~pi191 & n19556;
  assign n19558 = ~n19522 & ~n19557;
  assign n19559 = pi182 & n18117;
  assign n19560 = ~n19082 & ~n19559;
  assign n19561 = n19380 & ~n19560;
  assign n19562 = ~pi182 & ~pi372;
  assign n19563 = pi352 & n19496;
  assign n19564 = n19562 & n19563;
  assign n19565 = ~n19561 & ~n19564;
  assign n19566 = ~pi352 & n19187;
  assign n19567 = ~n19525 & ~n19566;
  assign n19568 = ~n18182 & n19567;
  assign n19569 = ~pi372 & ~n19568;
  assign n19570 = n19565 & ~n19569;
  assign n19571 = ~pi352 & n19411;
  assign n19572 = pi182 & n19541;
  assign n19573 = ~n19571 & ~n19572;
  assign n19574 = ~n18242 & ~n19392;
  assign n19575 = ~n18212 & ~n19064;
  assign n19576 = ~n18266 & n19575;
  assign n19577 = ~pi182 & ~n19576;
  assign n19578 = n19574 & ~n19577;
  assign n19579 = pi352 & ~n19578;
  assign n19580 = pi182 & ~n19382;
  assign n19581 = ~n19185 & ~n19580;
  assign n19582 = pi182 & n19232;
  assign n19583 = n19581 & ~n19582;
  assign n19584 = ~pi352 & ~n19583;
  assign n19585 = ~n19579 & ~n19584;
  assign n19586 = pi372 & ~n19585;
  assign n19587 = n19573 & ~n19586;
  assign n19588 = n19570 & n19587;
  assign n19589 = ~n19558 & n19588;
  assign n19590 = pi228 & n19589;
  assign n19591 = ~pi228 & ~n19589;
  assign n19592 = ~n19590 & ~n19591;
  assign n19593 = ~n19484 & n19592;
  assign n19594 = n19484 & ~n19592;
  assign n19595 = ~n19593 & ~n19594;
  assign n19596 = ~pi532 & ~n19595;
  assign n19597 = pi532 & pi580;
  assign po293 = n19596 | n19597;
  assign n19599 = ~pi133 & ~pi149;
  assign n19600 = pi133 & pi149;
  assign n19601 = ~n19599 & ~n19600;
  assign n19602 = ~pi148 & pi157;
  assign n19603 = pi148 & ~pi157;
  assign n19604 = ~n19602 & ~n19603;
  assign n19605 = ~n19601 & n19604;
  assign n19606 = n19601 & ~n19604;
  assign n19607 = ~n19605 & ~n19606;
  assign n19608 = n17944 & ~n19607;
  assign n19609 = ~n17944 & n19607;
  assign n19610 = ~n19608 & ~n19609;
  assign n19611 = ~pi532 & ~n19610;
  assign n19612 = pi532 & pi554;
  assign po294 = n19611 | n19612;
  assign n19614 = pi270 & n6328;
  assign n19615 = ~pi270 & ~n6328;
  assign po295 = n19614 | n19615;
  assign n19617 = ~pi159 & pi269;
  assign n19618 = pi159 & ~pi269;
  assign n19619 = ~n19617 & ~n19618;
  assign n19620 = pi352 & n19448;
  assign n19621 = ~n18160 & ~n19156;
  assign n19622 = ~pi352 & ~n19621;
  assign n19623 = n18205 & ~n19167;
  assign n19624 = ~n19622 & ~n19623;
  assign n19625 = ~n18256 & ~n19082;
  assign n19626 = ~n19186 & n19625;
  assign n19627 = n19624 & n19626;
  assign n19628 = ~n19620 & n19627;
  assign n19629 = pi372 & ~n19628;
  assign n19630 = ~pi352 & n19062;
  assign n19631 = ~n19137 & ~n19630;
  assign n19632 = ~n19563 & n19631;
  assign n19633 = ~n19536 & n19632;
  assign n19634 = ~pi372 & ~n19633;
  assign n19635 = ~pi182 & n19514;
  assign n19636 = pi182 & n18118;
  assign n19637 = ~n19635 & ~n19636;
  assign n19638 = pi352 & ~n19637;
  assign n19639 = ~pi352 & n19158;
  assign n19640 = ~n19638 & ~n19639;
  assign n19641 = ~n18142 & ~n18197;
  assign n19642 = ~pi182 & n18128;
  assign n19643 = ~n18129 & ~n19642;
  assign n19644 = ~n18255 & n19643;
  assign n19645 = ~pi352 & ~n19644;
  assign n19646 = n18119 & n18172;
  assign n19647 = ~n19645 & ~n19646;
  assign n19648 = n19641 & n19647;
  assign n19649 = pi372 & ~n19648;
  assign n19650 = ~n19065 & ~n19649;
  assign n19651 = n19640 & n19650;
  assign n19652 = ~n19634 & n19651;
  assign n19653 = ~pi191 & ~n19652;
  assign n19654 = ~n19629 & ~n19653;
  assign n19655 = n18252 & n19548;
  assign n19656 = ~n18209 & ~n19655;
  assign n19657 = ~pi352 & n19113;
  assign n19658 = ~n19392 & ~n19502;
  assign n19659 = ~n18213 & n19658;
  assign n19660 = pi352 & ~n19659;
  assign n19661 = pi352 & n19047;
  assign n19662 = ~n19660 & ~n19661;
  assign n19663 = ~n19466 & n19662;
  assign n19664 = ~n19657 & n19663;
  assign n19665 = n19656 & n19664;
  assign n19666 = ~n19065 & ~n19104;
  assign n19667 = n19665 & n19666;
  assign n19668 = ~pi372 & ~n19667;
  assign n19669 = n19654 & ~n19668;
  assign n19670 = ~pi321 & pi352;
  assign n19671 = n19544 & n19670;
  assign n19672 = ~pi182 & ~pi342;
  assign n19673 = n18124 & n19672;
  assign n19674 = ~n19671 & ~n19673;
  assign n19675 = n18129 & n19380;
  assign n19676 = ~pi352 & n19204;
  assign n19677 = ~n19385 & ~n19676;
  assign n19678 = ~pi372 & ~n19677;
  assign n19679 = ~n19675 & ~n19678;
  assign n19680 = pi182 & n18121;
  assign n19681 = ~n18267 & ~n19680;
  assign n19682 = ~pi372 & ~n19681;
  assign n19683 = n19679 & ~n19682;
  assign n19684 = ~n18150 & n19683;
  assign n19685 = ~n18212 & ~n18249;
  assign n19686 = ~pi352 & ~n19685;
  assign n19687 = ~n18237 & ~n19079;
  assign n19688 = ~n19041 & n19687;
  assign n19689 = ~n19686 & n19688;
  assign n19690 = pi372 & ~n19689;
  assign n19691 = ~n19086 & ~n19156;
  assign n19692 = ~n18186 & n19691;
  assign n19693 = ~pi352 & ~n19692;
  assign n19694 = ~n19690 & ~n19693;
  assign n19695 = n19684 & n19694;
  assign n19696 = ~n18199 & n19695;
  assign n19697 = n19674 & n19696;
  assign n19698 = pi191 & ~n19697;
  assign n19699 = n19669 & ~n19698;
  assign n19700 = ~pi352 & n18138;
  assign n19701 = ~n19563 & ~n19700;
  assign n19702 = pi182 & ~n19701;
  assign n19703 = n19699 & ~n19702;
  assign n19704 = pi301 & n19703;
  assign n19705 = ~pi301 & ~n19703;
  assign n19706 = ~n19704 & ~n19705;
  assign n19707 = ~n19619 & n19706;
  assign n19708 = n19619 & ~n19706;
  assign n19709 = ~n19707 & ~n19708;
  assign n19710 = ~pi532 & ~n19709;
  assign n19711 = pi532 & pi577;
  assign po296 = n19710 | n19711;
  assign n19713 = pi160 & n18398;
  assign n19714 = ~pi160 & ~n18398;
  assign n19715 = ~n19713 & ~n19714;
  assign n19716 = pi394 & n19715;
  assign n19717 = ~pi394 & ~n19715;
  assign n19718 = ~n19716 & ~n19717;
  assign n19719 = ~pi532 & ~n19718;
  assign n19720 = pi532 & pi653;
  assign po297 = n19719 | n19720;
  assign n19722 = pi132 & n17720;
  assign n19723 = n17661 & n17733;
  assign n19724 = ~n19722 & ~n19723;
  assign n19725 = pi284 & ~n19724;
  assign n19726 = pi132 & n17597;
  assign n19727 = pi275 & ~pi358;
  assign n19728 = ~n19726 & ~n19727;
  assign n19729 = ~n18045 & n19728;
  assign n19730 = ~n18308 & n19729;
  assign n19731 = n18792 & ~n19730;
  assign n19732 = ~n19725 & ~n19731;
  assign n19733 = pi358 & n18023;
  assign n19734 = ~n18045 & ~n19733;
  assign n19735 = ~n17980 & n19734;
  assign n19736 = ~pi351 & ~n19735;
  assign n19737 = ~n18004 & ~n19736;
  assign n19738 = ~n17714 & n19737;
  assign n19739 = n17702 & n17963;
  assign n19740 = n19738 & ~n19739;
  assign n19741 = ~pi358 & n17612;
  assign n19742 = pi132 & n19741;
  assign n19743 = ~n18372 & ~n19742;
  assign n19744 = n19740 & n19743;
  assign n19745 = ~pi284 & ~n19744;
  assign n19746 = ~pi351 & n18372;
  assign n19747 = ~n19745 & ~n19746;
  assign n19748 = ~pi132 & n18061;
  assign n19749 = ~n17614 & ~n19748;
  assign n19750 = pi351 & ~n19749;
  assign n19751 = n17608 & n17708;
  assign n19752 = ~n19750 & ~n19751;
  assign n19753 = ~n17626 & n19752;
  assign n19754 = ~n18355 & n19753;
  assign n19755 = n19747 & n19754;
  assign n19756 = n19732 & n19755;
  assign n19757 = pi193 & ~n19756;
  assign n19758 = ~pi132 & n17652;
  assign n19759 = ~n18341 & ~n19758;
  assign n19760 = ~pi351 & ~n19759;
  assign n19761 = ~pi351 & n17694;
  assign n19762 = ~n19760 & ~n19761;
  assign n19763 = ~n17738 & n19762;
  assign n19764 = pi351 & n17634;
  assign n19765 = n17608 & n17995;
  assign n19766 = ~n19764 & ~n19765;
  assign n19767 = ~n18345 & n19766;
  assign n19768 = ~pi284 & ~n19767;
  assign n19769 = ~pi351 & ~pi358;
  assign n19770 = ~pi284 & pi354;
  assign n19771 = n19769 & n19770;
  assign n19772 = ~n19768 & ~n19771;
  assign n19773 = pi132 & ~pi275;
  assign n19774 = pi358 & n19773;
  assign n19775 = pi132 & n17598;
  assign n19776 = ~n19774 & ~n19775;
  assign n19777 = ~pi351 & ~n19776;
  assign n19778 = pi358 & n17707;
  assign n19779 = n17702 & n19778;
  assign n19780 = ~n19777 & ~n19779;
  assign n19781 = ~n18798 & n19780;
  assign n19782 = ~n18836 & n19781;
  assign n19783 = pi284 & ~n19782;
  assign n19784 = pi351 & n17973;
  assign n19785 = ~n17761 & ~n19784;
  assign n19786 = n17608 & n17642;
  assign n19787 = n19785 & ~n19786;
  assign n19788 = ~n19783 & n19787;
  assign n19789 = n19772 & n19788;
  assign n19790 = n19763 & n19789;
  assign n19791 = ~pi193 & ~n19790;
  assign n19792 = ~n19757 & ~n19791;
  assign n19793 = ~n17635 & ~n19722;
  assign n19794 = n18317 & ~n19793;
  assign n19795 = ~pi132 & ~pi284;
  assign n19796 = pi351 & n19733;
  assign n19797 = n19795 & n19796;
  assign n19798 = ~n19794 & ~n19797;
  assign n19799 = ~pi351 & n18812;
  assign n19800 = ~n19760 & ~n19799;
  assign n19801 = ~n18005 & n19800;
  assign n19802 = ~pi284 & ~n19801;
  assign n19803 = n19798 & ~n19802;
  assign n19804 = pi132 & n17694;
  assign n19805 = ~n17631 & ~n19804;
  assign n19806 = ~pi351 & ~n19805;
  assign n19807 = n19803 & ~n19806;
  assign n19808 = pi132 & ~n18301;
  assign n19809 = ~n18810 & ~n19808;
  assign n19810 = ~n17744 & n19809;
  assign n19811 = ~pi351 & ~n19810;
  assign n19812 = ~n17640 & ~n17671;
  assign n19813 = ~n17662 & ~n17758;
  assign n19814 = ~n18061 & n19813;
  assign n19815 = ~pi132 & ~n19814;
  assign n19816 = n19812 & ~n19815;
  assign n19817 = pi351 & ~n19816;
  assign n19818 = ~n19811 & ~n19817;
  assign n19819 = pi284 & ~n19818;
  assign n19820 = n19807 & ~n19819;
  assign n19821 = n19792 & n19820;
  assign n19822 = pi161 & n19821;
  assign n19823 = ~pi161 & ~n19821;
  assign n19824 = ~n19822 & ~n19823;
  assign n19825 = pi392 & n19824;
  assign n19826 = ~pi392 & ~n19824;
  assign n19827 = ~n19825 & ~n19826;
  assign n19828 = ~pi532 & ~n19827;
  assign n19829 = pi532 & pi660;
  assign po298 = n19828 | n19829;
  assign n19831 = ~pi160 & pi162;
  assign n19832 = pi160 & ~pi162;
  assign n19833 = ~n19831 & ~n19832;
  assign n19834 = ~n18401 & ~n19833;
  assign n19835 = n18401 & n19833;
  assign po299 = n19834 | n19835;
  assign n19837 = ~pi161 & ~pi163;
  assign n19838 = pi161 & pi163;
  assign n19839 = ~n19837 & ~n19838;
  assign n19840 = pi392 & n19821;
  assign n19841 = ~pi392 & ~n19821;
  assign n19842 = ~n19840 & ~n19841;
  assign n19843 = ~n19839 & n19842;
  assign n19844 = n19839 & ~n19842;
  assign n19845 = ~n19843 & ~n19844;
  assign n19846 = ~pi532 & ~n19845;
  assign n19847 = pi532 & pi628;
  assign po301 = n19846 | n19847;
  assign n19849 = ~pi160 & pi164;
  assign n19850 = pi160 & ~pi164;
  assign n19851 = ~n19849 & ~n19850;
  assign n19852 = pi394 & n19851;
  assign n19853 = ~pi394 & ~n19851;
  assign n19854 = ~n19852 & ~n19853;
  assign n19855 = pi162 & n18398;
  assign n19856 = ~pi162 & ~n18398;
  assign n19857 = ~n19855 & ~n19856;
  assign n19858 = ~n19854 & n19857;
  assign n19859 = n19854 & ~n19857;
  assign n19860 = ~n19858 & ~n19859;
  assign n19861 = ~pi532 & ~n19860;
  assign n19862 = pi532 & pi589;
  assign po302 = n19861 | n19862;
  assign n19864 = ~pi161 & pi165;
  assign n19865 = pi161 & ~pi165;
  assign n19866 = ~n19864 & ~n19865;
  assign n19867 = pi392 & n19866;
  assign n19868 = ~pi392 & ~n19866;
  assign n19869 = ~n19867 & ~n19868;
  assign n19870 = ~pi163 & n19821;
  assign n19871 = pi163 & ~n19821;
  assign n19872 = ~n19870 & ~n19871;
  assign n19873 = ~n19869 & n19872;
  assign n19874 = n19869 & ~n19872;
  assign n19875 = ~n19873 & ~n19874;
  assign n19876 = ~pi532 & ~n19875;
  assign n19877 = pi532 & pi596;
  assign po303 = n19876 | n19877;
  assign n19879 = ~pi163 & ~pi165;
  assign n19880 = pi163 & pi165;
  assign n19881 = ~n19879 & ~n19880;
  assign n19882 = ~pi161 & pi166;
  assign n19883 = pi161 & ~pi166;
  assign n19884 = ~n19882 & ~n19883;
  assign n19885 = ~n19881 & n19884;
  assign n19886 = n19881 & ~n19884;
  assign n19887 = ~n19885 & ~n19886;
  assign n19888 = n19842 & ~n19887;
  assign n19889 = ~n19842 & n19887;
  assign n19890 = ~n19888 & ~n19889;
  assign n19891 = ~pi532 & ~n19890;
  assign n19892 = pi532 & pi564;
  assign po304 = n19891 | n19892;
  assign n19894 = pi167 & n18617;
  assign n19895 = ~pi167 & ~n18617;
  assign n19896 = ~n19894 & ~n19895;
  assign n19897 = ~pi532 & ~n19896;
  assign n19898 = pi532 & pi634;
  assign po305 = n19897 | n19898;
  assign n19900 = ~pi168 & pi271;
  assign n19901 = pi168 & ~pi271;
  assign n19902 = ~n19900 & ~n19901;
  assign n19903 = ~pi231 & n17430;
  assign n19904 = pi175 & n17279;
  assign n19905 = ~pi231 & n19904;
  assign n19906 = ~n19903 & ~n19905;
  assign n19907 = ~n17340 & n19906;
  assign n19908 = pi175 & n17897;
  assign n19909 = pi231 & n19908;
  assign n19910 = n19907 & ~n19909;
  assign n19911 = ~n17348 & ~n17422;
  assign n19912 = ~n17429 & n19911;
  assign n19913 = n19910 & n19912;
  assign n19914 = ~pi285 & ~n19913;
  assign n19915 = pi231 & n17439;
  assign n19916 = ~n19914 & ~n19915;
  assign n19917 = ~n17869 & n19916;
  assign n19918 = ~n17341 & ~n19283;
  assign n19919 = n17301 & n17351;
  assign n19920 = ~n19349 & ~n19919;
  assign n19921 = pi231 & ~n19920;
  assign n19922 = ~pi175 & n17284;
  assign n19923 = pi270 & n19325;
  assign n19924 = ~n17331 & ~n17849;
  assign n19925 = n17382 & ~n19924;
  assign n19926 = ~n17302 & ~n19925;
  assign n19927 = ~n19923 & n19926;
  assign n19928 = ~n19922 & n19927;
  assign n19929 = ~pi231 & ~n19928;
  assign n19930 = n17320 & n17328;
  assign n19931 = pi231 & n17397;
  assign n19932 = ~n19930 & ~n19931;
  assign n19933 = pi285 & ~n19932;
  assign n19934 = ~pi231 & n17906;
  assign n19935 = ~n17918 & ~n19934;
  assign n19936 = pi285 & ~n19935;
  assign n19937 = ~n19933 & ~n19936;
  assign n19938 = ~n17887 & ~n19919;
  assign n19939 = pi175 & pi233;
  assign n19940 = pi270 & n19939;
  assign n19941 = ~pi231 & n19940;
  assign n19942 = ~pi175 & n17838;
  assign n19943 = ~n19941 & ~n19942;
  assign n19944 = pi175 & n17835;
  assign n19945 = pi231 & n19944;
  assign n19946 = pi175 & n17332;
  assign n19947 = ~n19945 & ~n19946;
  assign n19948 = n19943 & n19947;
  assign n19949 = n19938 & n19948;
  assign n19950 = ~pi285 & ~n19949;
  assign n19951 = n19937 & ~n19950;
  assign n19952 = ~n19929 & n19951;
  assign n19953 = ~n19921 & n19952;
  assign n19954 = ~pi234 & ~n19953;
  assign n19955 = pi285 & n17939;
  assign n19956 = ~n19954 & ~n19955;
  assign n19957 = pi175 & n17282;
  assign n19958 = ~n17407 & ~n19957;
  assign n19959 = ~n17315 & n19958;
  assign n19960 = n17930 & ~n19959;
  assign n19961 = n19956 & ~n19960;
  assign n19962 = ~pi232 & pi270;
  assign n19963 = ~n17283 & ~n19962;
  assign n19964 = n17289 & ~n19963;
  assign n19965 = n19314 & ~n19964;
  assign n19966 = ~n17282 & ~n17366;
  assign n19967 = ~pi175 & n17324;
  assign n19968 = n19966 & ~n19967;
  assign n19969 = pi231 & ~n19968;
  assign n19970 = n19965 & ~n19969;
  assign n19971 = pi285 & n19970;
  assign n19972 = ~pi175 & n17835;
  assign n19973 = ~pi231 & n19972;
  assign n19974 = ~n17907 & ~n19973;
  assign n19975 = ~n17905 & n19974;
  assign n19976 = ~n17280 & n19975;
  assign n19977 = ~n17318 & ~n19940;
  assign n19978 = pi231 & ~n19977;
  assign n19979 = n19976 & ~n19978;
  assign n19980 = ~pi285 & n19979;
  assign n19981 = ~n19971 & ~n19980;
  assign n19982 = ~n17355 & ~n17365;
  assign n19983 = ~n17906 & n19982;
  assign n19984 = ~n17367 & n19983;
  assign n19985 = pi231 & ~n19984;
  assign n19986 = ~n17877 & ~n17887;
  assign n19987 = ~pi231 & ~n19986;
  assign n19988 = ~n19985 & ~n19987;
  assign n19989 = ~n19981 & n19988;
  assign n19990 = pi234 & ~n19989;
  assign n19991 = n19961 & ~n19990;
  assign n19992 = n19918 & n19991;
  assign n19993 = n19917 & n19992;
  assign n19994 = pi273 & n19993;
  assign n19995 = ~pi273 & ~n19993;
  assign n19996 = ~n19994 & ~n19995;
  assign n19997 = ~n19902 & n19996;
  assign n19998 = n19902 & ~n19996;
  assign n19999 = ~n19997 & ~n19998;
  assign n20000 = ~pi532 & ~n19999;
  assign n20001 = pi532 & pi587;
  assign po306 = n20000 | n20001;
  assign n20003 = pi169 & ~pi272;
  assign n20004 = ~pi169 & pi272;
  assign n20005 = ~n20003 & ~n20004;
  assign n20006 = pi138 & n18558;
  assign n20007 = pi207 & n20006;
  assign n20008 = ~pi207 & n18559;
  assign n20009 = pi138 & n18472;
  assign n20010 = ~pi207 & n20009;
  assign n20011 = ~n20008 & ~n20010;
  assign n20012 = ~n18574 & n20011;
  assign n20013 = ~n20007 & n20012;
  assign n20014 = ~n18645 & ~n18699;
  assign n20015 = ~n18707 & n20014;
  assign n20016 = n20013 & n20015;
  assign n20017 = ~pi302 & ~n20016;
  assign n20018 = pi207 & n18741;
  assign n20019 = ~n20017 & ~n20018;
  assign n20020 = ~n18550 & n20019;
  assign n20021 = n18509 & n18596;
  assign n20022 = ~n18985 & ~n20021;
  assign n20023 = pi207 & ~n20022;
  assign n20024 = ~pi138 & n18722;
  assign n20025 = pi185 & n18961;
  assign n20026 = ~n18495 & ~n18631;
  assign n20027 = n18512 & ~n20026;
  assign n20028 = ~n18673 & ~n20027;
  assign n20029 = ~n20025 & n20028;
  assign n20030 = ~n20024 & n20029;
  assign n20031 = ~pi207 & ~n20030;
  assign n20032 = n18489 & n18562;
  assign n20033 = pi207 & n18679;
  assign n20034 = ~n20032 & ~n20033;
  assign n20035 = pi302 & ~n20034;
  assign n20036 = ~pi207 & n18573;
  assign n20037 = ~n18589 & ~n20036;
  assign n20038 = pi302 & ~n20037;
  assign n20039 = ~n20035 & ~n20038;
  assign n20040 = ~n18539 & ~n20021;
  assign n20041 = pi138 & pi166;
  assign n20042 = pi185 & n20041;
  assign n20043 = ~pi207 & n20042;
  assign n20044 = ~pi138 & n18470;
  assign n20045 = ~n20043 & ~n20044;
  assign n20046 = pi138 & n18477;
  assign n20047 = pi207 & n20046;
  assign n20048 = pi138 & n18632;
  assign n20049 = ~n20047 & ~n20048;
  assign n20050 = n20045 & n20049;
  assign n20051 = n20040 & n20050;
  assign n20052 = ~pi302 & ~n20051;
  assign n20053 = n20039 & ~n20052;
  assign n20054 = ~n20031 & n20053;
  assign n20055 = ~n20023 & n20054;
  assign n20056 = ~pi139 & ~n20055;
  assign n20057 = pi302 & n18611;
  assign n20058 = ~n20056 & ~n20057;
  assign n20059 = pi138 & n18541;
  assign n20060 = ~n18594 & ~n20059;
  assign n20061 = ~n18481 & n20060;
  assign n20062 = pi207 & pi302;
  assign n20063 = ~n20061 & n20062;
  assign n20064 = n20058 & ~n20063;
  assign n20065 = ~pi129 & pi185;
  assign n20066 = ~n18459 & ~n20065;
  assign n20067 = n18585 & ~n20066;
  assign n20068 = n18955 & ~n20067;
  assign n20069 = ~pi138 & n18571;
  assign n20070 = ~n18541 & ~n20069;
  assign n20071 = ~n18657 & n20070;
  assign n20072 = pi207 & ~n20071;
  assign n20073 = n20068 & ~n20072;
  assign n20074 = pi302 & n20073;
  assign n20075 = ~pi138 & n18477;
  assign n20076 = ~pi207 & n20075;
  assign n20077 = ~n18575 & ~n20076;
  assign n20078 = ~n18572 & n20077;
  assign n20079 = ~n18473 & n20078;
  assign n20080 = ~n18490 & ~n20042;
  assign n20081 = pi207 & ~n20080;
  assign n20082 = n20079 & ~n20081;
  assign n20083 = ~pi302 & n20082;
  assign n20084 = ~n20074 & ~n20083;
  assign n20085 = ~n18456 & ~n18500;
  assign n20086 = ~n18573 & n20085;
  assign n20087 = ~n18658 & n20086;
  assign n20088 = pi207 & ~n20087;
  assign n20089 = ~n18528 & ~n18539;
  assign n20090 = ~pi207 & ~n20089;
  assign n20091 = ~n20088 & ~n20090;
  assign n20092 = ~n20084 & n20091;
  assign n20093 = pi139 & ~n20092;
  assign n20094 = n20064 & ~n20093;
  assign n20095 = ~n18639 & ~n18920;
  assign n20096 = n20094 & n20095;
  assign n20097 = n20020 & n20096;
  assign n20098 = pi274 & n20097;
  assign n20099 = ~pi274 & ~n20097;
  assign n20100 = ~n20098 & ~n20099;
  assign n20101 = ~n20005 & n20100;
  assign n20102 = n20005 & ~n20100;
  assign n20103 = ~n20101 & ~n20102;
  assign n20104 = ~pi532 & ~n20103;
  assign n20105 = pi532 & pi571;
  assign po307 = n20104 | n20105;
  assign n20107 = ~pi142 & ~pi178;
  assign n20108 = pi142 & pi178;
  assign n20109 = ~n20107 & ~n20108;
  assign n20110 = ~pi167 & pi170;
  assign n20111 = pi167 & ~pi170;
  assign n20112 = ~n20110 & ~n20111;
  assign n20113 = ~n20109 & n20112;
  assign n20114 = n20109 & ~n20112;
  assign n20115 = ~n20113 & ~n20114;
  assign n20116 = n18617 & ~n20115;
  assign n20117 = ~n18617 & n20115;
  assign n20118 = ~n20116 & ~n20117;
  assign n20119 = ~pi532 & ~n20118;
  assign n20120 = pi532 & pi538;
  assign po308 = n20119 | n20120;
  assign n20122 = pi532 & pi640;
  assign n20123 = pi171 & n18274;
  assign n20124 = ~pi171 & ~n18274;
  assign n20125 = ~n20123 & ~n20124;
  assign n20126 = ~pi532 & ~n20125;
  assign po309 = n20122 | n20126;
  assign n20128 = pi532 & pi608;
  assign n20129 = ~pi171 & pi172;
  assign n20130 = pi171 & ~pi172;
  assign n20131 = ~n20129 & ~n20130;
  assign n20132 = n18274 & ~n20131;
  assign n20133 = ~n18274 & n20131;
  assign n20134 = ~n20132 & ~n20133;
  assign n20135 = ~pi532 & ~n20134;
  assign po310 = n20128 | n20135;
  assign n20137 = ~pi173 & pi278;
  assign n20138 = pi173 & ~pi278;
  assign n20139 = ~n20137 & ~n20138;
  assign n20140 = pi270 & n17297;
  assign n20141 = pi175 & n20140;
  assign n20142 = ~n17325 & ~n20141;
  assign n20143 = ~n19919 & n20142;
  assign n20144 = n17930 & ~n20143;
  assign n20145 = ~pi175 & n17292;
  assign n20146 = ~n17407 & ~n20145;
  assign n20147 = ~n17365 & n20146;
  assign n20148 = n19335 & ~n20147;
  assign n20149 = ~n17404 & ~n17837;
  assign n20150 = pi175 & n17318;
  assign n20151 = ~n17316 & ~n20150;
  assign n20152 = ~n19313 & n20151;
  assign n20153 = ~pi231 & ~n20152;
  assign n20154 = n20149 & ~n20153;
  assign n20155 = ~pi285 & ~n20154;
  assign n20156 = ~n20148 & ~n20155;
  assign n20157 = ~n20144 & n20156;
  assign n20158 = pi175 & n17390;
  assign n20159 = ~n17887 & ~n17906;
  assign n20160 = ~pi231 & ~n20159;
  assign n20161 = ~pi270 & n17384;
  assign n20162 = n17289 & n20161;
  assign n20163 = ~n20160 & ~n20162;
  assign n20164 = ~n20158 & n20163;
  assign n20165 = ~n19973 & n20164;
  assign n20166 = pi285 & ~n20165;
  assign n20167 = n20157 & ~n20166;
  assign n20168 = ~pi175 & n17282;
  assign n20169 = ~pi231 & n17428;
  assign n20170 = ~n20168 & ~n20169;
  assign n20171 = n17408 & n17847;
  assign n20172 = ~n17429 & ~n20171;
  assign n20173 = ~n17319 & n20172;
  assign n20174 = n20170 & n20173;
  assign n20175 = ~pi285 & ~n20174;
  assign n20176 = ~n17836 & ~n19325;
  assign n20177 = ~n17319 & n20176;
  assign n20178 = ~n19904 & n20177;
  assign n20179 = ~pi231 & ~n20178;
  assign n20180 = ~pi175 & n17836;
  assign n20181 = ~n20179 & ~n20180;
  assign n20182 = ~n20175 & n20181;
  assign n20183 = ~n19919 & n20182;
  assign n20184 = pi231 & n17418;
  assign n20185 = n20183 & ~n20184;
  assign n20186 = pi270 & n17849;
  assign n20187 = pi175 & n17300;
  assign n20188 = ~n20186 & ~n20187;
  assign n20189 = ~n17332 & n20188;
  assign n20190 = pi231 & ~n20189;
  assign n20191 = ~n17357 & ~n20190;
  assign n20192 = ~n17324 & n20191;
  assign n20193 = pi285 & ~n20192;
  assign n20194 = n20185 & ~n20193;
  assign n20195 = pi234 & ~n20194;
  assign n20196 = ~pi175 & n17346;
  assign n20197 = ~n17396 & ~n20196;
  assign n20198 = pi231 & ~n20197;
  assign n20199 = pi175 & ~n20186;
  assign n20200 = ~pi175 & ~n17278;
  assign n20201 = ~n20199 & ~n20200;
  assign n20202 = ~n17827 & ~n20201;
  assign n20203 = ~pi231 & ~n20202;
  assign n20204 = ~n20198 & ~n20203;
  assign n20205 = n17822 & n20204;
  assign n20206 = ~n17886 & n20205;
  assign n20207 = pi285 & ~n20206;
  assign n20208 = pi231 & n19325;
  assign n20209 = ~n17303 & ~n20208;
  assign n20210 = pi175 & n17347;
  assign n20211 = ~n17439 & ~n19903;
  assign n20212 = ~pi231 & n19967;
  assign n20213 = n20211 & ~n20212;
  assign n20214 = ~n20210 & n20213;
  assign n20215 = n20209 & n20214;
  assign n20216 = ~pi285 & ~n20215;
  assign n20217 = ~n20207 & ~n20216;
  assign n20218 = n17320 & n17327;
  assign n20219 = ~n17869 & ~n20218;
  assign n20220 = ~n17940 & n20219;
  assign n20221 = ~pi231 & n20210;
  assign n20222 = ~n17407 & ~n20221;
  assign n20223 = ~n17377 & n20222;
  assign n20224 = n20220 & n20223;
  assign n20225 = n20217 & n20224;
  assign n20226 = ~pi234 & ~n20225;
  assign n20227 = ~n20195 & ~n20226;
  assign n20228 = n17296 & n17906;
  assign n20229 = ~n17438 & ~n20228;
  assign n20230 = n20227 & n20229;
  assign n20231 = n20167 & n20230;
  assign n20232 = pi281 & n20231;
  assign n20233 = ~pi281 & ~n20231;
  assign n20234 = ~n20232 & ~n20233;
  assign n20235 = ~n20139 & n20234;
  assign n20236 = n20139 & ~n20234;
  assign n20237 = ~n20235 & ~n20236;
  assign n20238 = ~pi532 & ~n20237;
  assign n20239 = pi532 & pi582;
  assign po311 = n20238 | n20239;
  assign n20241 = ~pi174 & pi280;
  assign n20242 = pi174 & ~pi280;
  assign n20243 = ~n20241 & ~n20242;
  assign n20244 = n19670 & n19672;
  assign n20245 = ~n19153 & ~n20244;
  assign n20246 = ~pi352 & n19211;
  assign n20247 = ~n18260 & ~n19063;
  assign n20248 = ~n19113 & ~n19139;
  assign n20249 = n20247 & n20248;
  assign n20250 = ~n18245 & n20249;
  assign n20251 = ~n20246 & n20250;
  assign n20252 = ~pi372 & ~n20251;
  assign n20253 = ~n18181 & ~n19523;
  assign n20254 = pi352 & ~n20253;
  assign n20255 = ~pi182 & ~n18127;
  assign n20256 = pi182 & ~n19548;
  assign n20257 = ~n20255 & ~n20256;
  assign n20258 = ~n19159 & ~n20257;
  assign n20259 = ~pi352 & ~n20258;
  assign n20260 = ~n19086 & ~n19392;
  assign n20261 = ~n19559 & n20260;
  assign n20262 = ~n20259 & n20261;
  assign n20263 = ~n20254 & n20262;
  assign n20264 = pi372 & ~n20263;
  assign n20265 = ~n20252 & ~n20264;
  assign n20266 = ~n18223 & n20265;
  assign n20267 = ~n19453 & n20266;
  assign n20268 = n20245 & n20267;
  assign n20269 = ~n18211 & ~n19657;
  assign n20270 = n20268 & n20269;
  assign n20271 = ~pi191 & ~n20270;
  assign n20272 = ~pi182 & n18157;
  assign n20273 = n18200 & n19102;
  assign n20274 = ~n18229 & ~n20273;
  assign n20275 = ~n18138 & n20274;
  assign n20276 = ~pi352 & n18228;
  assign n20277 = n20275 & ~n20276;
  assign n20278 = ~n20272 & n20277;
  assign n20279 = ~pi372 & ~n20278;
  assign n20280 = ~n19158 & ~n20279;
  assign n20281 = ~n19062 & ~n19084;
  assign n20282 = ~n19066 & n20281;
  assign n20283 = ~n18138 & n20282;
  assign n20284 = ~pi352 & ~n20283;
  assign n20285 = ~pi182 & n19066;
  assign n20286 = ~n20284 & ~n20285;
  assign n20287 = ~n19090 & ~n19548;
  assign n20288 = ~n18114 & n20287;
  assign n20289 = pi352 & ~n20288;
  assign n20290 = ~n18163 & ~n20289;
  assign n20291 = ~n18242 & n20290;
  assign n20292 = pi372 & ~n20291;
  assign n20293 = pi352 & n18208;
  assign n20294 = ~n20292 & ~n20293;
  assign n20295 = n20286 & n20294;
  assign n20296 = n20280 & n20295;
  assign n20297 = pi191 & ~n20296;
  assign n20298 = ~n20271 & ~n20297;
  assign n20299 = pi182 & n19496;
  assign n20300 = ~n19158 & ~n20299;
  assign n20301 = ~n18243 & n20300;
  assign n20302 = n19020 & ~n20301;
  assign n20303 = ~pi182 & n18161;
  assign n20304 = ~n18211 & ~n20303;
  assign n20305 = ~n18145 & n20304;
  assign n20306 = n19380 & ~n20305;
  assign n20307 = ~n18213 & ~n19203;
  assign n20308 = ~n18237 & ~n19205;
  assign n20309 = ~n19543 & n20308;
  assign n20310 = ~pi352 & ~n20309;
  assign n20311 = n20307 & ~n20310;
  assign n20312 = ~pi372 & ~n20311;
  assign n20313 = ~n20306 & ~n20312;
  assign n20314 = ~n20302 & n20313;
  assign n20315 = pi182 & n18183;
  assign n20316 = ~n18191 & ~n19172;
  assign n20317 = ~pi352 & ~n20316;
  assign n20318 = n18252 & n19501;
  assign n20319 = ~n20317 & ~n20318;
  assign n20320 = ~n20315 & n20319;
  assign n20321 = ~n19110 & n20320;
  assign n20322 = pi372 & ~n20321;
  assign n20323 = ~n18270 & ~n19531;
  assign n20324 = ~n20322 & n20323;
  assign n20325 = n20314 & n20324;
  assign n20326 = n20298 & n20325;
  assign n20327 = pi283 & n20326;
  assign n20328 = ~pi283 & ~n20326;
  assign n20329 = ~n20327 & ~n20328;
  assign n20330 = ~n20243 & n20329;
  assign n20331 = n20243 & ~n20329;
  assign n20332 = ~n20330 & ~n20331;
  assign n20333 = ~pi532 & ~n20332;
  assign n20334 = pi532 & pi574;
  assign po312 = n20333 | n20334;
  assign n20336 = pi532 & pi544;
  assign n20337 = pi137 & ~pi172;
  assign n20338 = ~pi137 & pi172;
  assign n20339 = ~n20337 & ~n20338;
  assign n20340 = ~pi171 & pi175;
  assign n20341 = pi171 & ~pi175;
  assign n20342 = ~n20340 & ~n20341;
  assign n20343 = ~n20339 & n20342;
  assign n20344 = n20339 & ~n20342;
  assign n20345 = ~n20343 & ~n20344;
  assign n20346 = n18274 & ~n20345;
  assign n20347 = ~n18274 & n20345;
  assign n20348 = ~n20346 & ~n20347;
  assign n20349 = ~pi532 & ~n20348;
  assign po313 = n20336 | n20349;
  assign n20351 = pi141 & n13902;
  assign n20352 = ~pi141 & ~n13902;
  assign po314 = n20351 | n20352;
  assign n20354 = pi159 & n7504;
  assign n20355 = ~pi159 & ~n7504;
  assign po315 = n20354 | n20355;
  assign n20357 = ~pi167 & ~pi178;
  assign n20358 = pi167 & pi178;
  assign n20359 = ~n20357 & ~n20358;
  assign n20360 = n18617 & ~n20359;
  assign n20361 = ~n18617 & n20359;
  assign n20362 = ~n20360 & ~n20361;
  assign n20363 = ~pi532 & ~n20362;
  assign n20364 = pi532 & pi602;
  assign po316 = n20363 | n20364;
  assign n20366 = ~pi179 & pi223;
  assign n20367 = pi179 & ~pi223;
  assign n20368 = ~n20366 & ~n20367;
  assign n20369 = n18252 & n19204;
  assign n20370 = ~n19043 & ~n20369;
  assign n20371 = ~n19540 & n20370;
  assign n20372 = ~n18137 & ~n18161;
  assign n20373 = n18153 & ~n20372;
  assign n20374 = ~n19582 & ~n20373;
  assign n20375 = ~n18145 & n20374;
  assign n20376 = pi352 & ~n20375;
  assign n20377 = ~n18211 & ~n20376;
  assign n20378 = n20371 & n20377;
  assign n20379 = ~pi372 & ~n20378;
  assign n20380 = pi372 & n18119;
  assign n20381 = n19421 & n20380;
  assign n20382 = pi182 & n19172;
  assign n20383 = ~n18130 & ~n20382;
  assign n20384 = pi372 & ~n20383;
  assign n20385 = ~n20381 & ~n20384;
  assign n20386 = ~n20379 & n20385;
  assign n20387 = ~n19384 & ~n19514;
  assign n20388 = pi352 & n20387;
  assign n20389 = ~pi352 & ~n18162;
  assign n20390 = ~n20388 & ~n20389;
  assign n20391 = ~n18145 & ~n19392;
  assign n20392 = ~n19495 & n20391;
  assign n20393 = ~n20390 & n20392;
  assign n20394 = ~pi372 & ~n20393;
  assign n20395 = ~n18236 & ~n20394;
  assign n20396 = pi352 & n18145;
  assign n20397 = ~n19159 & ~n19220;
  assign n20398 = pi170 & n19166;
  assign n20399 = n20397 & ~n20398;
  assign n20400 = n19052 & ~n20399;
  assign n20401 = ~n18222 & ~n19416;
  assign n20402 = ~n18237 & n20401;
  assign n20403 = ~n19203 & n20402;
  assign n20404 = pi372 & ~n20403;
  assign n20405 = ~n20400 & ~n20404;
  assign n20406 = ~n18192 & ~n19043;
  assign n20407 = ~n18201 & n20260;
  assign n20408 = ~pi352 & ~n20407;
  assign n20409 = n20406 & ~n20408;
  assign n20410 = n20405 & n20409;
  assign n20411 = ~n20396 & n20410;
  assign n20412 = n20395 & n20411;
  assign n20413 = pi191 & ~n20412;
  assign n20414 = n20386 & ~n20413;
  assign n20415 = n18121 & n18198;
  assign n20416 = ~n18228 & ~n19233;
  assign n20417 = ~pi182 & n18249;
  assign n20418 = n20416 & ~n20417;
  assign n20419 = ~pi352 & ~n20418;
  assign n20420 = pi182 & n18181;
  assign n20421 = ~n19411 & ~n20420;
  assign n20422 = ~n19517 & n20421;
  assign n20423 = ~n20419 & n20422;
  assign n20424 = ~n20415 & n20423;
  assign n20425 = ~n18157 & ~n19559;
  assign n20426 = ~n18208 & n20425;
  assign n20427 = n20424 & n20426;
  assign n20428 = pi372 & ~n20427;
  assign n20429 = ~n18111 & ~n20420;
  assign n20430 = ~n18210 & n20429;
  assign n20431 = ~n19456 & n20430;
  assign n20432 = pi352 & ~n20431;
  assign n20433 = ~n20428 & ~n20432;
  assign n20434 = ~pi182 & n18212;
  assign n20435 = n18198 & n19159;
  assign n20436 = ~n20434 & ~n20435;
  assign n20437 = ~n18160 & n20436;
  assign n20438 = ~n19153 & n20437;
  assign n20439 = ~pi372 & ~n20438;
  assign n20440 = n19222 & ~n20439;
  assign n20441 = n20433 & n20440;
  assign n20442 = ~n19172 & n20441;
  assign n20443 = ~n18130 & n20442;
  assign n20444 = ~pi191 & ~n20443;
  assign n20445 = n20414 & ~n20444;
  assign n20446 = ~n18209 & n20445;
  assign n20447 = ~n19453 & n20446;
  assign n20448 = ~n19080 & n20447;
  assign n20449 = ~pi226 & n20448;
  assign n20450 = pi226 & ~n20448;
  assign n20451 = ~n20449 & ~n20450;
  assign n20452 = ~n20368 & n20451;
  assign n20453 = n20368 & ~n20451;
  assign n20454 = ~n20452 & ~n20453;
  assign n20455 = ~pi532 & ~n20454;
  assign n20456 = pi532 & pi578;
  assign po317 = n20455 | n20456;
  assign n20458 = pi532 & pi600;
  assign n20459 = pi180 & ~pi181;
  assign n20460 = ~pi180 & pi181;
  assign n20461 = ~n20459 & ~n20460;
  assign n20462 = n18745 & ~n20461;
  assign n20463 = ~n18745 & n20461;
  assign n20464 = ~n20462 & ~n20463;
  assign n20465 = ~pi532 & ~n20464;
  assign po318 = n20458 | n20465;
  assign n20467 = pi532 & pi632;
  assign n20468 = pi181 & n18745;
  assign n20469 = ~pi181 & ~n18745;
  assign n20470 = ~n20468 & ~n20469;
  assign n20471 = ~pi532 & ~n20470;
  assign po319 = n20467 | n20471;
  assign n20473 = pi532 & pi536;
  assign n20474 = pi143 & ~pi180;
  assign n20475 = ~pi143 & pi180;
  assign n20476 = ~n20474 & ~n20475;
  assign n20477 = ~pi181 & pi182;
  assign n20478 = pi181 & ~pi182;
  assign n20479 = ~n20477 & ~n20478;
  assign n20480 = ~n20476 & n20479;
  assign n20481 = n20476 & ~n20479;
  assign n20482 = ~n20480 & ~n20481;
  assign n20483 = n18745 & ~n20482;
  assign n20484 = ~n18745 & n20482;
  assign n20485 = ~n20483 & ~n20484;
  assign n20486 = ~pi532 & ~n20485;
  assign po320 = n20473 | n20486;
  assign n20488 = ~pi183 & pi319;
  assign n20489 = pi183 & ~pi319;
  assign n20490 = ~n20488 & ~n20489;
  assign n20491 = ~pi207 & n20021;
  assign n20492 = pi207 & n18480;
  assign n20493 = pi185 & n18697;
  assign n20494 = pi207 & n20493;
  assign n20495 = ~pi207 & n18961;
  assign n20496 = ~n20006 & ~n20495;
  assign n20497 = ~n20494 & n20496;
  assign n20498 = ~n20492 & n20497;
  assign n20499 = ~pi302 & ~n20498;
  assign n20500 = ~n20491 & ~n20499;
  assign n20501 = ~pi138 & n18496;
  assign n20502 = pi138 & n18481;
  assign n20503 = ~n20501 & ~n20502;
  assign n20504 = pi207 & ~n20503;
  assign n20505 = ~pi138 & n18472;
  assign n20506 = ~n18473 & ~n20505;
  assign n20507 = ~n18727 & n20506;
  assign n20508 = ~pi207 & ~n20507;
  assign n20509 = n18489 & n18669;
  assign n20510 = ~n20508 & ~n20509;
  assign n20511 = ~n18690 & n20510;
  assign n20512 = ~n18658 & n20511;
  assign n20513 = pi302 & ~n20512;
  assign n20514 = ~n18908 & ~n20513;
  assign n20515 = ~n20504 & n20514;
  assign n20516 = n20500 & n20515;
  assign n20517 = ~pi139 & ~n20516;
  assign n20518 = pi185 & n18495;
  assign n20519 = n18585 & n20518;
  assign n20520 = pi138 & n18644;
  assign n20521 = ~pi207 & n20520;
  assign n20522 = ~n20519 & ~n20521;
  assign n20523 = ~n18614 & n20522;
  assign n20524 = pi207 & n20075;
  assign n20525 = ~pi185 & n18526;
  assign n20526 = pi138 & n20525;
  assign n20527 = ~n18688 & ~n20526;
  assign n20528 = ~n18445 & n20527;
  assign n20529 = pi207 & ~n20528;
  assign n20530 = ~n20524 & ~n20529;
  assign n20531 = n20523 & n20530;
  assign n20532 = ~n18927 & n20531;
  assign n20533 = ~n18589 & ~n18908;
  assign n20534 = n20532 & n20533;
  assign n20535 = ~pi302 & ~n20534;
  assign n20536 = pi207 & n18910;
  assign n20537 = ~n18548 & ~n18920;
  assign n20538 = ~pi207 & ~n20537;
  assign n20539 = n18465 & ~n20026;
  assign n20540 = ~n20538 & ~n20539;
  assign n20541 = pi138 & n18510;
  assign n20542 = ~n20047 & ~n20541;
  assign n20543 = ~n18728 & n20542;
  assign n20544 = n20540 & n20543;
  assign n20545 = ~n20536 & n20544;
  assign n20546 = pi302 & ~n20545;
  assign n20547 = ~n20535 & ~n20546;
  assign n20548 = ~pi207 & n18491;
  assign n20549 = ~n20494 & ~n20548;
  assign n20550 = pi138 & ~n20549;
  assign n20551 = ~pi147 & ~pi185;
  assign n20552 = n18534 & n20551;
  assign n20553 = ~n18692 & ~n20552;
  assign n20554 = n18461 & n18489;
  assign n20555 = n20553 & ~n20554;
  assign n20556 = n18473 & n18971;
  assign n20557 = ~pi207 & n18586;
  assign n20558 = ~n18977 & ~n20557;
  assign n20559 = ~pi302 & ~n20558;
  assign n20560 = ~n20556 & ~n20559;
  assign n20561 = pi138 & n18522;
  assign n20562 = ~n18738 & ~n20561;
  assign n20563 = ~pi302 & ~n20562;
  assign n20564 = n20560 & ~n20563;
  assign n20565 = ~n18447 & ~n18673;
  assign n20566 = ~n18920 & n20565;
  assign n20567 = ~pi207 & ~n20566;
  assign n20568 = n20564 & ~n20567;
  assign n20569 = ~n18446 & ~n18553;
  assign n20570 = ~pi207 & ~n20569;
  assign n20571 = pi207 & n18470;
  assign n20572 = ~n18482 & ~n18610;
  assign n20573 = ~n20571 & n20572;
  assign n20574 = ~n20570 & n20573;
  assign n20575 = pi302 & ~n20574;
  assign n20576 = n20568 & ~n20575;
  assign n20577 = ~n18645 & n20576;
  assign n20578 = n20555 & n20577;
  assign n20579 = pi139 & ~n20578;
  assign n20580 = ~n20550 & ~n20579;
  assign n20581 = n20547 & n20580;
  assign n20582 = ~n20517 & n20581;
  assign n20583 = pi320 & n20582;
  assign n20584 = ~pi320 & ~n20582;
  assign n20585 = ~n20583 & ~n20584;
  assign n20586 = ~n20490 & n20585;
  assign n20587 = n20490 & ~n20585;
  assign n20588 = ~n20586 & ~n20587;
  assign n20589 = ~pi532 & ~n20588;
  assign n20590 = pi532 & pi569;
  assign po321 = n20589 | n20590;
  assign n20592 = pi532 & pi625;
  assign n20593 = ~pi184 & ~pi255;
  assign n20594 = pi184 & pi255;
  assign n20595 = ~n20593 & ~n20594;
  assign n20596 = ~pi351 & n18798;
  assign n20597 = ~pi351 & n18360;
  assign n20598 = ~n18834 & ~n20597;
  assign n20599 = ~n19796 & n20598;
  assign n20600 = ~n19764 & n20599;
  assign n20601 = ~pi284 & ~n20600;
  assign n20602 = ~n20596 & ~n20601;
  assign n20603 = ~pi132 & n17708;
  assign n20604 = ~n19804 & ~n20603;
  assign n20605 = pi351 & ~n20604;
  assign n20606 = ~pi132 & n17632;
  assign n20607 = ~n17643 & ~n20606;
  assign n20608 = ~n18050 & n20607;
  assign n20609 = ~pi351 & ~n20608;
  assign n20610 = n17702 & n17995;
  assign n20611 = ~n20609 & ~n20610;
  assign n20612 = ~n18016 & n20611;
  assign n20613 = ~n17981 & n20612;
  assign n20614 = pi284 & ~n20613;
  assign n20615 = ~n18371 & ~n20614;
  assign n20616 = ~n20605 & n20615;
  assign n20617 = n20602 & n20616;
  assign n20618 = ~pi193 & ~n20617;
  assign n20619 = pi351 & n18761;
  assign n20620 = ~n17671 & ~n19742;
  assign n20621 = ~n18014 & n20620;
  assign n20622 = pi351 & ~n20621;
  assign n20623 = ~n20619 & ~n20622;
  assign n20624 = ~n18392 & n20623;
  assign n20625 = pi132 & n17653;
  assign n20626 = ~pi351 & n20625;
  assign n20627 = n17733 & n19778;
  assign n20628 = ~n17763 & ~n20627;
  assign n20629 = ~n20626 & n20628;
  assign n20630 = n20624 & n20629;
  assign n20631 = ~n17737 & ~n18371;
  assign n20632 = n20630 & n20631;
  assign n20633 = ~pi284 & ~n20632;
  assign n20634 = pi351 & n18372;
  assign n20635 = ~n17654 & ~n18384;
  assign n20636 = ~pi351 & ~n20635;
  assign n20637 = n17645 & ~n18803;
  assign n20638 = ~n20636 & ~n20637;
  assign n20639 = ~n18811 & ~n19722;
  assign n20640 = ~n18051 & n20639;
  assign n20641 = n20638 & n20640;
  assign n20642 = ~n20634 & n20641;
  assign n20643 = pi284 & ~n20642;
  assign n20644 = ~n20633 & ~n20643;
  assign n20645 = ~pi351 & n17703;
  assign n20646 = ~n19796 & ~n20645;
  assign n20647 = pi132 & ~n20646;
  assign n20648 = ~pi275 & ~pi358;
  assign n20649 = n17608 & n20648;
  assign n20650 = ~n18018 & ~n20649;
  assign n20651 = n17646 & n17702;
  assign n20652 = n20650 & ~n20651;
  assign n20653 = n17643 & n18317;
  assign n20654 = ~pi351 & n17734;
  assign n20655 = ~n18300 & ~n20654;
  assign n20656 = ~pi284 & ~n20655;
  assign n20657 = ~n20653 & ~n20656;
  assign n20658 = pi132 & n17592;
  assign n20659 = ~n18062 & ~n20658;
  assign n20660 = ~pi284 & ~n20659;
  assign n20661 = n20657 & ~n20660;
  assign n20662 = ~n17672 & ~n17999;
  assign n20663 = ~n18384 & n20662;
  assign n20664 = ~pi351 & ~n20663;
  assign n20665 = n20661 & ~n20664;
  assign n20666 = ~n17616 & ~n17662;
  assign n20667 = ~pi351 & ~n20666;
  assign n20668 = pi351 & n17687;
  assign n20669 = ~n17695 & ~n17759;
  assign n20670 = ~n20668 & n20669;
  assign n20671 = ~n20667 & n20670;
  assign n20672 = pi284 & ~n20671;
  assign n20673 = n20665 & ~n20672;
  assign n20674 = ~n17968 & n20673;
  assign n20675 = n20652 & n20674;
  assign n20676 = pi193 & ~n20675;
  assign n20677 = ~n20647 & ~n20676;
  assign n20678 = n20644 & n20677;
  assign n20679 = ~n20618 & n20678;
  assign n20680 = pi384 & ~n20679;
  assign n20681 = ~pi384 & n20679;
  assign n20682 = ~n20680 & ~n20681;
  assign n20683 = ~n20595 & n20682;
  assign n20684 = n20595 & ~n20682;
  assign n20685 = ~n20683 & ~n20684;
  assign n20686 = ~pi532 & ~n20685;
  assign po322 = n20592 | n20686;
  assign n20688 = pi532 & pi561;
  assign n20689 = ~pi184 & ~pi221;
  assign n20690 = pi184 & pi221;
  assign n20691 = ~n20689 & ~n20690;
  assign n20692 = pi185 & ~pi255;
  assign n20693 = ~pi185 & pi255;
  assign n20694 = ~n20692 & ~n20693;
  assign n20695 = ~n20691 & n20694;
  assign n20696 = n20691 & ~n20694;
  assign n20697 = ~n20695 & ~n20696;
  assign n20698 = n20682 & ~n20697;
  assign n20699 = ~n20682 & n20697;
  assign n20700 = ~n20698 & ~n20699;
  assign n20701 = ~pi532 & ~n20700;
  assign po323 = n20688 | n20701;
  assign n20703 = pi144 & n12557;
  assign n20704 = ~pi144 & ~n12557;
  assign po324 = n20703 | n20704;
  assign n20706 = pi532 & pi629;
  assign n20707 = pi187 & n19004;
  assign n20708 = ~pi187 & ~n19004;
  assign n20709 = ~n20707 & ~n20708;
  assign n20710 = ~pi532 & ~n20709;
  assign po325 = n20706 | n20710;
  assign n20712 = ~pi140 & n10094;
  assign n20713 = pi140 & ~n10094;
  assign po326 = n20712 | n20713;
  assign n20715 = pi532 & pi645;
  assign n20716 = pi189 & n19367;
  assign n20717 = ~pi189 & ~n19367;
  assign n20718 = ~n20716 & ~n20717;
  assign n20719 = ~pi532 & ~n20718;
  assign po327 = n20715 | n20719;
  assign n20721 = pi532 & pi597;
  assign n20722 = pi187 & pi190;
  assign n20723 = ~pi187 & ~pi190;
  assign n20724 = ~n20722 & ~n20723;
  assign n20725 = n19004 & ~n20724;
  assign n20726 = ~n19004 & n20724;
  assign n20727 = ~n20725 & ~n20726;
  assign n20728 = ~pi532 & ~n20727;
  assign po328 = n20721 | n20728;
  assign n20730 = pi532 & pi533;
  assign n20731 = pi150 & pi190;
  assign n20732 = ~pi150 & ~pi190;
  assign n20733 = ~n20731 & ~n20732;
  assign n20734 = pi187 & ~pi191;
  assign n20735 = ~pi187 & pi191;
  assign n20736 = ~n20734 & ~n20735;
  assign n20737 = ~n20733 & n20736;
  assign n20738 = n20733 & ~n20736;
  assign n20739 = ~n20737 & ~n20738;
  assign n20740 = n19004 & ~n20739;
  assign n20741 = ~n19004 & n20739;
  assign n20742 = ~n20740 & ~n20741;
  assign n20743 = ~pi532 & ~n20742;
  assign po329 = n20730 | n20743;
  assign n20745 = pi532 & pi613;
  assign n20746 = ~pi189 & ~pi192;
  assign n20747 = pi189 & pi192;
  assign n20748 = ~n20746 & ~n20747;
  assign n20749 = n19367 & ~n20748;
  assign n20750 = ~n19367 & n20748;
  assign n20751 = ~n20749 & ~n20750;
  assign n20752 = ~pi532 & ~n20751;
  assign po330 = n20745 | n20752;
  assign n20754 = pi532 & pi549;
  assign n20755 = ~pi154 & ~pi192;
  assign n20756 = pi154 & pi192;
  assign n20757 = ~n20755 & ~n20756;
  assign n20758 = ~pi189 & pi193;
  assign n20759 = pi189 & ~pi193;
  assign n20760 = ~n20758 & ~n20759;
  assign n20761 = ~n20757 & n20760;
  assign n20762 = n20757 & ~n20760;
  assign n20763 = ~n20761 & ~n20762;
  assign n20764 = n19367 & ~n20763;
  assign n20765 = ~n19367 & n20763;
  assign n20766 = ~n20764 & ~n20765;
  assign n20767 = ~pi532 & ~n20766;
  assign po331 = n20754 | n20767;
  assign n20769 = pi167 & n13628;
  assign n20770 = ~pi167 & ~n13628;
  assign po332 = n20769 | n20770;
  assign n20772 = pi269 & n9455;
  assign n20773 = ~pi269 & ~n9455;
  assign po333 = n20772 | n20773;
  assign n20775 = pi137 & n1752;
  assign n20776 = ~pi137 & ~n1752;
  assign po334 = n20775 | n20776;
  assign n20778 = pi223 & n13537;
  assign n20779 = ~pi223 & ~n13537;
  assign po335 = n20778 | n20779;
  assign n20781 = pi148 & n13441;
  assign n20782 = ~pi148 & ~n13441;
  assign po336 = n20781 | n20782;
  assign n20784 = pi301 & n12252;
  assign n20785 = ~pi301 & ~n12252;
  assign po337 = n20784 | n20785;
  assign n20787 = pi224 & n8748;
  assign n20788 = ~pi224 & ~n8748;
  assign po338 = n20787 | n20788;
  assign n20790 = pi154 & n3141;
  assign n20791 = ~pi154 & ~n3141;
  assign po339 = n20790 | n20791;
  assign n20793 = ~pi192 & n4161;
  assign n20794 = pi192 & ~n4161;
  assign po340 = n20793 | n20794;
  assign n20796 = pi189 & n5192;
  assign n20797 = ~pi189 & ~n5192;
  assign po341 = n20796 | n20797;
  assign n20799 = pi152 & n10348;
  assign n20800 = ~pi152 & ~n10348;
  assign po342 = n20799 | n20800;
  assign n20802 = pi145 & n13810;
  assign n20803 = ~pi145 & ~n13810;
  assign po343 = n20802 | n20803;
  assign n20805 = ~pi231 & ~n11175;
  assign n20806 = pi231 & n11175;
  assign po344 = n20805 | n20806;
  assign n20808 = ~pi208 & ~pi209;
  assign n20809 = pi208 & pi209;
  assign n20810 = ~n20808 & ~n20809;
  assign n20811 = pi207 & ~pi210;
  assign n20812 = ~pi207 & pi210;
  assign n20813 = ~n20811 & ~n20812;
  assign n20814 = ~n20810 & n20813;
  assign n20815 = n20810 & ~n20813;
  assign n20816 = ~n20814 & ~n20815;
  assign n20817 = ~n17737 & ~n18034;
  assign n20818 = ~n17758 & n20817;
  assign n20819 = ~pi351 & ~n20818;
  assign n20820 = pi132 & n18045;
  assign n20821 = ~n20819 & ~n20820;
  assign n20822 = ~n18762 & n20821;
  assign n20823 = pi132 & n17658;
  assign n20824 = ~n20625 & ~n20823;
  assign n20825 = pi351 & ~n20824;
  assign n20826 = n20822 & ~n20825;
  assign n20827 = ~n18050 & ~n18825;
  assign n20828 = n20826 & n20827;
  assign n20829 = ~pi284 & ~n20828;
  assign n20830 = pi275 & pi358;
  assign n20831 = ~pi132 & n20830;
  assign n20832 = ~n18045 & ~n20831;
  assign n20833 = n17681 & ~n20832;
  assign n20834 = pi351 & n17596;
  assign n20835 = ~n18370 & ~n20834;
  assign n20836 = pi284 & ~n20835;
  assign n20837 = ~n20833 & ~n20836;
  assign n20838 = pi351 & n18003;
  assign n20839 = ~pi351 & n17743;
  assign n20840 = ~n20668 & ~n20839;
  assign n20841 = ~n18016 & n20840;
  assign n20842 = ~n20838 & n20841;
  assign n20843 = ~n17721 & n20842;
  assign n20844 = ~n18062 & n20843;
  assign n20845 = ~n18341 & n20844;
  assign n20846 = ~n18761 & n20845;
  assign n20847 = ~pi284 & ~n20846;
  assign n20848 = n20837 & ~n20847;
  assign n20849 = pi351 & n18360;
  assign n20850 = ~n17599 & ~n17692;
  assign n20851 = ~n17652 & n20850;
  assign n20852 = n17608 & ~n20851;
  assign n20853 = ~n20849 & ~n20852;
  assign n20854 = ~n18371 & ~n18391;
  assign n20855 = n20853 & n20854;
  assign n20856 = n20848 & n20855;
  assign n20857 = pi193 & ~n20856;
  assign n20858 = ~n17672 & ~n18308;
  assign n20859 = pi351 & ~n20858;
  assign n20860 = pi132 & n17620;
  assign n20861 = ~n18352 & ~n20860;
  assign n20862 = ~n17602 & n20861;
  assign n20863 = ~pi351 & ~n20862;
  assign n20864 = ~n20859 & ~n20863;
  assign n20865 = ~n18836 & n20864;
  assign n20866 = pi284 & ~n20865;
  assign n20867 = pi351 & n19722;
  assign n20868 = ~n20866 & ~n20867;
  assign n20869 = n17645 & n17674;
  assign n20870 = ~n18005 & ~n20869;
  assign n20871 = ~pi284 & ~n20870;
  assign n20872 = ~n17643 & ~n17760;
  assign n20873 = ~n20871 & n20872;
  assign n20874 = n20868 & n20873;
  assign n20875 = ~pi193 & ~n20874;
  assign n20876 = ~n20857 & ~n20875;
  assign n20877 = ~n17691 & ~n17962;
  assign n20878 = n17702 & ~n20877;
  assign n20879 = ~pi358 & n20878;
  assign n20880 = ~n18052 & ~n20879;
  assign n20881 = n17608 & n17703;
  assign n20882 = pi284 & n20881;
  assign n20883 = n17610 & n17745;
  assign n20884 = ~n17640 & ~n20883;
  assign n20885 = ~pi351 & ~n20884;
  assign n20886 = ~n17622 & ~n20885;
  assign n20887 = ~pi351 & n17973;
  assign n20888 = n20886 & ~n20887;
  assign n20889 = pi284 & ~n20888;
  assign n20890 = ~n20882 & ~n20889;
  assign n20891 = pi354 & ~pi358;
  assign n20892 = ~pi132 & n20891;
  assign n20893 = ~n17720 & ~n20892;
  assign n20894 = n18792 & ~n20893;
  assign n20895 = n20890 & ~n20894;
  assign n20896 = n20880 & n20895;
  assign n20897 = n20876 & n20896;
  assign n20898 = ~n20829 & n20897;
  assign n20899 = pi385 & n20898;
  assign n20900 = ~pi385 & ~n20898;
  assign n20901 = ~n20899 & ~n20900;
  assign n20902 = ~n20816 & n20901;
  assign n20903 = n20816 & ~n20901;
  assign n20904 = ~n20902 & ~n20903;
  assign n20905 = ~pi532 & ~n20904;
  assign n20906 = pi532 & pi559;
  assign po345 = n20905 | n20906;
  assign n20908 = ~pi208 & ~pi210;
  assign n20909 = pi208 & pi210;
  assign n20910 = ~n20908 & ~n20909;
  assign n20911 = n20901 & ~n20910;
  assign n20912 = ~n20901 & n20910;
  assign n20913 = ~n20911 & ~n20912;
  assign n20914 = ~pi532 & ~n20913;
  assign n20915 = pi532 & pi623;
  assign po346 = n20914 | n20915;
  assign n20917 = pi209 & ~pi210;
  assign n20918 = ~pi209 & pi210;
  assign n20919 = ~n20917 & ~n20918;
  assign n20920 = pi385 & n20919;
  assign n20921 = ~pi385 & ~n20919;
  assign n20922 = ~n20920 & ~n20921;
  assign n20923 = ~pi208 & n20898;
  assign n20924 = pi208 & ~n20898;
  assign n20925 = ~n20923 & ~n20924;
  assign n20926 = ~n20922 & n20925;
  assign n20927 = n20922 & ~n20925;
  assign n20928 = ~n20926 & ~n20927;
  assign n20929 = ~pi532 & ~n20928;
  assign n20930 = pi532 & pi591;
  assign po347 = n20929 | n20930;
  assign n20932 = pi210 & n20898;
  assign n20933 = ~pi210 & ~n20898;
  assign n20934 = ~n20932 & ~n20933;
  assign n20935 = pi385 & n20934;
  assign n20936 = ~pi385 & ~n20934;
  assign n20937 = ~n20935 & ~n20936;
  assign n20938 = ~pi532 & ~n20937;
  assign n20939 = pi532 & pi655;
  assign po348 = n20938 | n20939;
  assign n20941 = pi191 & n9668;
  assign n20942 = ~pi191 & ~n9668;
  assign po349 = n20941 | n20942;
  assign n20944 = pi321 & n6060;
  assign n20945 = ~pi321 & ~n6060;
  assign po350 = n20944 | n20945;
  assign n20947 = pi276 & n14660;
  assign n20948 = ~pi276 & ~n14660;
  assign po351 = n20947 | n20948;
  assign n20950 = pi150 & n11307;
  assign n20951 = ~pi150 & ~n11307;
  assign po352 = n20950 | n20951;
  assign n20953 = pi532 & pi547;
  assign n20954 = pi152 & ~pi227;
  assign n20955 = ~pi152 & pi227;
  assign n20956 = ~n20954 & ~n20955;
  assign n20957 = pi215 & ~pi256;
  assign n20958 = ~pi215 & pi256;
  assign n20959 = ~n20957 & ~n20958;
  assign n20960 = ~n20956 & n20959;
  assign n20961 = n20956 & ~n20959;
  assign n20962 = ~n20960 & ~n20961;
  assign n20963 = n19241 & ~n20962;
  assign n20964 = ~n19241 & n20962;
  assign n20965 = ~n20963 & ~n20964;
  assign n20966 = ~pi532 & ~n20965;
  assign po353 = n20953 | n20966;
  assign n20968 = ~pi190 & n12964;
  assign n20969 = pi190 & ~n12964;
  assign po354 = n20968 | n20969;
  assign n20971 = ~pi217 & pi371;
  assign n20972 = pi217 & ~pi371;
  assign n20973 = ~n20971 & ~n20972;
  assign n20974 = ~n17429 & ~n17918;
  assign n20975 = ~n17937 & n20974;
  assign n20976 = ~pi231 & ~n20975;
  assign n20977 = pi175 & n17284;
  assign n20978 = ~n20976 & ~n20977;
  assign n20979 = ~n19973 & n20978;
  assign n20980 = pi175 & n17283;
  assign n20981 = ~n20210 & ~n20980;
  assign n20982 = pi231 & ~n20981;
  assign n20983 = n20979 & ~n20982;
  assign n20984 = ~n17293 & ~n19931;
  assign n20985 = n20983 & n20984;
  assign n20986 = ~pi285 & ~n20985;
  assign n20987 = pi215 & pi270;
  assign n20988 = ~pi175 & n20987;
  assign n20989 = ~n17284 & ~n20988;
  assign n20990 = n17826 & ~n20989;
  assign n20991 = pi231 & n17897;
  assign n20992 = ~n19269 & ~n20991;
  assign n20993 = pi285 & ~n20992;
  assign n20994 = ~n20990 & ~n20993;
  assign n20995 = pi231 & n17394;
  assign n20996 = ~pi231 & n17407;
  assign n20997 = pi231 & n17838;
  assign n20998 = ~n20996 & ~n20997;
  assign n20999 = ~n17411 & n20998;
  assign n21000 = ~n20995 & n20999;
  assign n21001 = ~n19306 & ~n19972;
  assign n21002 = ~n17309 & n21001;
  assign n21003 = ~n17862 & n21002;
  assign n21004 = n21000 & n21003;
  assign n21005 = ~pi285 & ~n21004;
  assign n21006 = n20994 & ~n21005;
  assign n21007 = ~n17430 & ~n17836;
  assign n21008 = ~n17346 & n21007;
  assign n21009 = n17296 & ~n21008;
  assign n21010 = ~n20208 & ~n21009;
  assign n21011 = ~n19270 & ~n19289;
  assign n21012 = n21010 & n21011;
  assign n21013 = n21006 & n21012;
  assign n21014 = pi234 & ~n21013;
  assign n21015 = n17408 & n17412;
  assign n21016 = ~n17397 & ~n21015;
  assign n21017 = ~pi285 & ~n21016;
  assign n21018 = ~n17280 & ~n17939;
  assign n21019 = ~n19321 & ~n20187;
  assign n21020 = ~n17328 & n21019;
  assign n21021 = ~pi231 & ~n21020;
  assign n21022 = ~n19904 & ~n21021;
  assign n21023 = ~n17821 & ~n19353;
  assign n21024 = pi231 & ~n21023;
  assign n21025 = n21022 & ~n21024;
  assign n21026 = pi285 & ~n21025;
  assign n21027 = pi175 & n17861;
  assign n21028 = pi231 & n21027;
  assign n21029 = ~n21026 & ~n21028;
  assign n21030 = n21018 & n21029;
  assign n21031 = ~n21017 & n21030;
  assign n21032 = ~pi234 & ~n21031;
  assign n21033 = ~n21014 & ~n21032;
  assign n21034 = ~n17331 & ~n17835;
  assign n21035 = n17320 & ~n21034;
  assign n21036 = ~pi270 & n21035;
  assign n21037 = ~n17295 & ~n21036;
  assign n21038 = pi175 & n17319;
  assign n21039 = n17930 & n21038;
  assign n21040 = n17278 & n17351;
  assign n21041 = ~n17324 & ~n21040;
  assign n21042 = ~pi231 & ~n21041;
  assign n21043 = ~n17418 & ~n21042;
  assign n21044 = ~pi231 & n17357;
  assign n21045 = n21043 & ~n21044;
  assign n21046 = pi285 & ~n21045;
  assign n21047 = ~n21039 & ~n21046;
  assign n21048 = pi233 & ~pi270;
  assign n21049 = ~pi175 & n21048;
  assign n21050 = ~n17861 & ~n21049;
  assign n21051 = n17930 & ~n21050;
  assign n21052 = n21047 & ~n21051;
  assign n21053 = n21037 & n21052;
  assign n21054 = n21033 & n21053;
  assign n21055 = ~n20986 & n21054;
  assign n21056 = pi346 & n21055;
  assign n21057 = ~pi346 & ~n21055;
  assign n21058 = ~n21056 & ~n21057;
  assign n21059 = ~n20973 & n21058;
  assign n21060 = n20973 & ~n21058;
  assign n21061 = ~n21059 & ~n21060;
  assign n21062 = ~pi532 & ~n21061;
  assign n21063 = pi532 & pi583;
  assign po355 = n21062 | n21063;
  assign n21065 = pi218 & ~pi349;
  assign n21066 = ~pi218 & pi349;
  assign n21067 = ~n21065 & ~n21066;
  assign n21068 = ~n18589 & ~n18707;
  assign n21069 = ~n18609 & n21068;
  assign n21070 = ~pi207 & ~n21069;
  assign n21071 = pi138 & n18722;
  assign n21072 = ~n21070 & ~n21071;
  assign n21073 = ~n20076 & n21072;
  assign n21074 = pi138 & n18459;
  assign n21075 = ~n20520 & ~n21074;
  assign n21076 = pi207 & ~n21075;
  assign n21077 = n21073 & ~n21076;
  assign n21078 = ~n18727 & ~n20033;
  assign n21079 = n21077 & n21078;
  assign n21080 = ~pi302 & ~n21079;
  assign n21081 = pi147 & pi185;
  assign n21082 = ~pi138 & n21081;
  assign n21083 = ~n18722 & ~n21082;
  assign n21084 = n18458 & ~n21083;
  assign n21085 = pi207 & n18558;
  assign n21086 = ~n18906 & ~n21085;
  assign n21087 = pi302 & ~n21086;
  assign n21088 = ~n21084 & ~n21087;
  assign n21089 = pi207 & n18677;
  assign n21090 = ~pi207 & n18594;
  assign n21091 = ~n20571 & ~n21090;
  assign n21092 = ~n18690 & n21091;
  assign n21093 = ~n21089 & n21092;
  assign n21094 = ~n18511 & n21093;
  assign n21095 = ~n18738 & n21094;
  assign n21096 = ~n18942 & n21095;
  assign n21097 = ~n20075 & n21096;
  assign n21098 = ~pi302 & ~n21097;
  assign n21099 = n21088 & ~n21098;
  assign n21100 = pi207 & n18961;
  assign n21101 = ~n18478 & ~n18559;
  assign n21102 = ~n18454 & n21101;
  assign n21103 = n18534 & ~n21102;
  assign n21104 = ~n21100 & ~n21103;
  assign n21105 = ~n18908 & ~n18926;
  assign n21106 = n21104 & n21105;
  assign n21107 = n21099 & n21106;
  assign n21108 = pi139 & ~n21107;
  assign n21109 = n18449 & n18465;
  assign n21110 = ~n18679 & ~n21109;
  assign n21111 = ~pi302 & ~n21110;
  assign n21112 = ~n18473 & ~n18611;
  assign n21113 = ~n18447 & ~n18989;
  assign n21114 = pi207 & ~n21113;
  assign n21115 = pi138 & n18453;
  assign n21116 = ~n18948 & ~n21115;
  assign n21117 = ~n18562 & n21116;
  assign n21118 = ~pi207 & ~n21117;
  assign n21119 = ~n21114 & ~n21118;
  assign n21120 = ~n20009 & n21119;
  assign n21121 = pi302 & ~n21120;
  assign n21122 = pi207 & n20541;
  assign n21123 = ~n21121 & ~n21122;
  assign n21124 = n21112 & n21123;
  assign n21125 = ~n21111 & n21124;
  assign n21126 = ~pi139 & ~n21125;
  assign n21127 = ~n21108 & ~n21126;
  assign n21128 = ~n18477 & ~n18631;
  assign n21129 = n18489 & ~n21128;
  assign n21130 = ~pi185 & n21129;
  assign n21131 = ~n18729 & ~n21130;
  assign n21132 = pi166 & ~pi185;
  assign n21133 = ~pi138 & n21132;
  assign n21134 = ~n18510 & ~n21133;
  assign n21135 = n20062 & ~n21134;
  assign n21136 = n18491 & n18534;
  assign n21137 = pi302 & n21136;
  assign n21138 = n18469 & n18596;
  assign n21139 = ~n18571 & ~n21138;
  assign n21140 = ~pi207 & ~n21139;
  assign n21141 = ~n18521 & ~n21140;
  assign n21142 = ~pi207 & n18646;
  assign n21143 = n21141 & ~n21142;
  assign n21144 = pi302 & ~n21143;
  assign n21145 = ~n21137 & ~n21144;
  assign n21146 = ~n21135 & n21145;
  assign n21147 = n21131 & n21146;
  assign n21148 = n21127 & n21147;
  assign n21149 = ~n21080 & n21148;
  assign n21150 = pi350 & n21149;
  assign n21151 = ~pi350 & ~n21149;
  assign n21152 = ~n21150 & ~n21151;
  assign n21153 = ~n21067 & n21152;
  assign n21154 = n21067 & ~n21152;
  assign n21155 = ~n21153 & ~n21154;
  assign n21156 = ~pi532 & ~n21155;
  assign n21157 = pi532 & pi567;
  assign po356 = n21156 | n21157;
  assign n21159 = ~pi219 & pi353;
  assign n21160 = pi219 & ~pi353;
  assign n21161 = ~n21159 & ~n21160;
  assign n21162 = ~n17886 & ~n21027;
  assign n21163 = n19335 & ~n21162;
  assign n21164 = ~pi175 & ~pi285;
  assign n21165 = pi231 & n20140;
  assign n21166 = n21164 & n21165;
  assign n21167 = ~n21163 & ~n21166;
  assign n21168 = ~n19306 & ~n20196;
  assign n21169 = ~pi231 & ~n21168;
  assign n21170 = ~pi231 & n19946;
  assign n21171 = ~n21169 & ~n21170;
  assign n21172 = ~n17397 & n21171;
  assign n21173 = ~pi285 & ~n21172;
  assign n21174 = n21167 & ~n21173;
  assign n21175 = pi175 & n17315;
  assign n21176 = ~n17888 & ~n21175;
  assign n21177 = ~pi231 & ~n21176;
  assign n21178 = n21174 & ~n21177;
  assign n21179 = ~pi231 & n17315;
  assign n21180 = ~n21169 & ~n21179;
  assign n21181 = pi231 & n17314;
  assign n21182 = n17296 & n17387;
  assign n21183 = ~n21181 & ~n21182;
  assign n21184 = ~pi285 & ~n21183;
  assign n21185 = n17310 & n21048;
  assign n21186 = ~n21184 & ~n21185;
  assign n21187 = ~pi285 & n19313;
  assign n21188 = n21186 & ~n21187;
  assign n21189 = ~n17919 & n21188;
  assign n21190 = n21180 & n21189;
  assign n21191 = pi231 & n17357;
  assign n21192 = ~n20228 & ~n21191;
  assign n21193 = ~n17940 & n21192;
  assign n21194 = n21190 & n21193;
  assign n21195 = pi175 & ~pi215;
  assign n21196 = pi270 & n21195;
  assign n21197 = ~n20150 & ~n21196;
  assign n21198 = ~pi231 & ~n21197;
  assign n21199 = n17320 & n20186;
  assign n21200 = ~n21198 & ~n21199;
  assign n21201 = ~n19919 & n21200;
  assign n21202 = ~n19904 & n21201;
  assign n21203 = pi285 & ~n21202;
  assign n21204 = n21194 & ~n21203;
  assign n21205 = ~pi234 & ~n21204;
  assign n21206 = n17289 & n17292;
  assign n21207 = ~n21027 & ~n21206;
  assign n21208 = pi285 & ~n21207;
  assign n21209 = pi175 & n17286;
  assign n21210 = pi215 & ~pi270;
  assign n21211 = ~n21209 & ~n21210;
  assign n21212 = ~n17284 & n21211;
  assign n21213 = ~n19353 & n21212;
  assign n21214 = n17930 & ~n21213;
  assign n21215 = ~n21208 & ~n21214;
  assign n21216 = ~n17284 & ~n17366;
  assign n21217 = ~n20140 & n21216;
  assign n21218 = ~pi231 & ~n21217;
  assign n21219 = ~n17855 & ~n21218;
  assign n21220 = pi175 & n20161;
  assign n21221 = ~n19271 & ~n21220;
  assign n21222 = pi231 & n17333;
  assign n21223 = n21221 & ~n21222;
  assign n21224 = ~n17395 & n21223;
  assign n21225 = n21219 & n21224;
  assign n21226 = ~pi285 & ~n21225;
  assign n21227 = ~pi231 & n19271;
  assign n21228 = ~n21226 & ~n21227;
  assign n21229 = ~pi175 & n17308;
  assign n21230 = ~n17877 & ~n21229;
  assign n21231 = pi231 & ~n21230;
  assign n21232 = n17296 & n17850;
  assign n21233 = ~n21231 & ~n21232;
  assign n21234 = ~n17885 & n21233;
  assign n21235 = ~n19310 & n21234;
  assign n21236 = n21228 & n21235;
  assign n21237 = n21215 & n21236;
  assign n21238 = pi234 & ~n21237;
  assign n21239 = ~n21205 & ~n21238;
  assign n21240 = pi175 & ~n19342;
  assign n21241 = ~n19944 & ~n21240;
  assign n21242 = ~n17921 & n21241;
  assign n21243 = ~pi231 & ~n21242;
  assign n21244 = ~n17324 & ~n17820;
  assign n21245 = ~n17403 & ~n17937;
  assign n21246 = ~n17308 & n21245;
  assign n21247 = ~pi175 & ~n21246;
  assign n21248 = n21244 & ~n21247;
  assign n21249 = pi231 & ~n21248;
  assign n21250 = ~n21243 & ~n21249;
  assign n21251 = pi285 & ~n21250;
  assign n21252 = n21239 & ~n21251;
  assign n21253 = n21178 & n21252;
  assign n21254 = pi375 & n21253;
  assign n21255 = ~pi375 & ~n21253;
  assign n21256 = ~n21254 & ~n21255;
  assign n21257 = ~n21161 & n21256;
  assign n21258 = n21161 & ~n21256;
  assign n21259 = ~n21257 & ~n21258;
  assign n21260 = ~pi532 & ~n21259;
  assign n21261 = pi532 & pi588;
  assign po357 = n21260 | n21261;
  assign n21263 = ~pi220 & pi356;
  assign n21264 = pi220 & ~pi356;
  assign n21265 = ~n21263 & ~n21264;
  assign n21266 = ~pi231 & n19919;
  assign n21267 = ~pi231 & n19325;
  assign n21268 = ~n19908 & ~n21267;
  assign n21269 = ~n21165 & n21268;
  assign n21270 = ~n21181 & n21269;
  assign n21271 = ~pi285 & ~n21270;
  assign n21272 = ~n21266 & ~n21271;
  assign n21273 = ~pi175 & n17850;
  assign n21274 = ~n21175 & ~n21273;
  assign n21275 = pi231 & ~n21274;
  assign n21276 = ~pi175 & n17279;
  assign n21277 = ~n17280 & ~n21276;
  assign n21278 = ~n17293 & n21277;
  assign n21279 = ~pi231 & ~n21278;
  assign n21280 = n17320 & n17387;
  assign n21281 = ~n21279 & ~n21280;
  assign n21282 = ~n17411 & n21281;
  assign n21283 = ~n17367 & n21282;
  assign n21284 = pi285 & ~n21283;
  assign n21285 = ~n19270 & ~n21284;
  assign n21286 = ~n21275 & n21285;
  assign n21287 = n21272 & n21286;
  assign n21288 = ~pi234 & ~n21287;
  assign n21289 = n17289 & n20186;
  assign n21290 = ~n20221 & ~n21289;
  assign n21291 = pi231 & n19972;
  assign n21292 = ~n17404 & ~n21220;
  assign n21293 = ~n17820 & n21292;
  assign n21294 = pi231 & ~n21293;
  assign n21295 = ~n21291 & ~n21294;
  assign n21296 = ~n19290 & n21295;
  assign n21297 = ~n17419 & n21296;
  assign n21298 = n21290 & n21297;
  assign n21299 = ~n17918 & ~n19270;
  assign n21300 = n21298 & n21299;
  assign n21301 = ~pi285 & ~n21300;
  assign n21302 = pi231 & n19271;
  assign n21303 = ~n17359 & ~n19283;
  assign n21304 = ~pi231 & ~n21303;
  assign n21305 = n17412 & ~n19924;
  assign n21306 = ~n21304 & ~n21305;
  assign n21307 = ~n19945 & ~n21027;
  assign n21308 = ~n17294 & n21307;
  assign n21309 = n21306 & n21308;
  assign n21310 = ~n21302 & n21309;
  assign n21311 = pi285 & ~n21310;
  assign n21312 = ~n21301 & ~n21311;
  assign n21313 = ~pi231 & n17319;
  assign n21314 = ~n21165 & ~n21313;
  assign n21315 = pi175 & ~n21314;
  assign n21316 = ~pi215 & ~pi270;
  assign n21317 = n17296 & n21316;
  assign n21318 = ~n17414 & ~n21317;
  assign n21319 = n17320 & n17828;
  assign n21320 = n21318 & ~n21319;
  assign n21321 = n17280 & n19335;
  assign n21322 = ~pi231 & n17914;
  assign n21323 = ~n19341 & ~n21322;
  assign n21324 = ~pi285 & ~n21323;
  assign n21325 = ~n21321 & ~n21324;
  assign n21326 = pi175 & n17336;
  assign n21327 = ~n17309 & ~n21326;
  assign n21328 = ~pi285 & ~n21327;
  assign n21329 = n21325 & ~n21328;
  assign n21330 = ~n17302 & ~n17821;
  assign n21331 = ~n19283 & n21330;
  assign n21332 = ~pi231 & ~n21331;
  assign n21333 = n21329 & ~n21332;
  assign n21334 = ~n17287 & ~n17403;
  assign n21335 = ~pi231 & ~n21334;
  assign n21336 = ~n17316 & ~n17938;
  assign n21337 = ~n20997 & n21336;
  assign n21338 = ~n21335 & n21337;
  assign n21339 = pi285 & ~n21338;
  assign n21340 = n21333 & ~n21339;
  assign n21341 = ~n17348 & n21340;
  assign n21342 = n21320 & n21341;
  assign n21343 = pi234 & ~n21342;
  assign n21344 = ~n21315 & ~n21343;
  assign n21345 = n21312 & n21344;
  assign n21346 = ~n21288 & n21345;
  assign n21347 = pi357 & n21346;
  assign n21348 = ~pi357 & ~n21346;
  assign n21349 = ~n21347 & ~n21348;
  assign n21350 = ~n21265 & n21349;
  assign n21351 = n21265 & ~n21349;
  assign n21352 = ~n21350 & ~n21351;
  assign n21353 = ~pi532 & ~n21352;
  assign n21354 = pi532 & pi585;
  assign po358 = n21353 | n21354;
  assign n21356 = pi221 & ~pi255;
  assign n21357 = ~pi221 & pi255;
  assign n21358 = ~n21356 & ~n21357;
  assign n21359 = pi384 & n21358;
  assign n21360 = ~pi384 & ~n21358;
  assign n21361 = ~n21359 & ~n21360;
  assign n21362 = pi184 & n20679;
  assign n21363 = ~pi184 & ~n20679;
  assign n21364 = ~n21362 & ~n21363;
  assign n21365 = ~n21361 & n21364;
  assign n21366 = n21361 & ~n21364;
  assign n21367 = ~n21365 & ~n21366;
  assign n21368 = ~pi532 & ~n21367;
  assign n21369 = pi532 & pi593;
  assign po359 = n21368 | n21369;
  assign n21371 = pi532 & pi639;
  assign n21372 = pi222 & n19124;
  assign n21373 = ~pi222 & ~n19124;
  assign n21374 = ~n21372 & ~n21373;
  assign n21375 = ~pi532 & ~n21374;
  assign po360 = n21371 | n21375;
  assign n21377 = pi532 & pi642;
  assign n21378 = pi223 & n20448;
  assign n21379 = ~pi223 & ~n20448;
  assign n21380 = ~n21378 & ~n21379;
  assign n21381 = ~pi532 & ~n21380;
  assign po361 = n21377 | n21381;
  assign n21383 = pi532 & pi644;
  assign n21384 = pi224 & n19589;
  assign n21385 = ~pi224 & ~n19589;
  assign n21386 = ~n21384 & ~n21385;
  assign n21387 = ~pi532 & ~n21386;
  assign po362 = n21383 | n21387;
  assign n21389 = pi532 & pi637;
  assign n21390 = pi225 & n19472;
  assign n21391 = ~pi225 & ~n19472;
  assign n21392 = ~n21390 & ~n21391;
  assign n21393 = ~pi532 & ~n21392;
  assign po363 = n21389 | n21393;
  assign n21395 = pi532 & pi610;
  assign n21396 = ~pi223 & ~pi226;
  assign n21397 = pi223 & pi226;
  assign n21398 = ~n21396 & ~n21397;
  assign n21399 = n20448 & ~n21398;
  assign n21400 = ~n20448 & n21398;
  assign n21401 = ~n21399 & ~n21400;
  assign n21402 = ~pi532 & ~n21401;
  assign po364 = n21395 | n21402;
  assign n21404 = pi532 & pi611;
  assign n21405 = pi227 & ~pi256;
  assign n21406 = ~pi227 & pi256;
  assign n21407 = ~n21405 & ~n21406;
  assign n21408 = n19241 & ~n21407;
  assign n21409 = ~n19241 & n21407;
  assign n21410 = ~n21408 & ~n21409;
  assign n21411 = ~pi532 & ~n21410;
  assign po365 = n21404 | n21411;
  assign n21413 = pi532 & pi612;
  assign n21414 = pi224 & ~pi228;
  assign n21415 = ~pi224 & pi228;
  assign n21416 = ~n21414 & ~n21415;
  assign n21417 = n19589 & ~n21416;
  assign n21418 = ~n19589 & n21416;
  assign n21419 = ~n21417 & ~n21418;
  assign n21420 = ~pi532 & ~n21419;
  assign po366 = n21413 | n21420;
  assign n21422 = pi532 & pi607;
  assign n21423 = ~pi222 & pi229;
  assign n21424 = pi222 & ~pi229;
  assign n21425 = ~n21423 & ~n21424;
  assign n21426 = n19124 & ~n21425;
  assign n21427 = ~n19124 & n21425;
  assign n21428 = ~n21426 & ~n21427;
  assign n21429 = ~pi532 & ~n21428;
  assign po367 = n21422 | n21429;
  assign n21431 = pi532 & pi605;
  assign n21432 = ~pi225 & pi230;
  assign n21433 = pi225 & ~pi230;
  assign n21434 = ~n21432 & ~n21433;
  assign n21435 = n19472 & ~n21434;
  assign n21436 = ~n19472 & n21434;
  assign n21437 = ~n21435 & ~n21436;
  assign n21438 = ~pi532 & ~n21437;
  assign po368 = n21431 | n21438;
  assign n21440 = pi532 & pi543;
  assign n21441 = pi151 & ~pi229;
  assign n21442 = ~pi151 & pi229;
  assign n21443 = ~n21441 & ~n21442;
  assign n21444 = ~pi222 & pi231;
  assign n21445 = pi222 & ~pi231;
  assign n21446 = ~n21444 & ~n21445;
  assign n21447 = ~n21443 & n21446;
  assign n21448 = n21443 & ~n21446;
  assign n21449 = ~n21447 & ~n21448;
  assign n21450 = n19124 & ~n21449;
  assign n21451 = ~n19124 & n21449;
  assign n21452 = ~n21450 & ~n21451;
  assign n21453 = ~pi532 & ~n21452;
  assign po369 = n21440 | n21453;
  assign n21455 = pi532 & pi546;
  assign n21456 = ~pi179 & ~pi226;
  assign n21457 = pi179 & pi226;
  assign n21458 = ~n21456 & ~n21457;
  assign n21459 = ~pi223 & pi232;
  assign n21460 = pi223 & ~pi232;
  assign n21461 = ~n21459 & ~n21460;
  assign n21462 = ~n21458 & n21461;
  assign n21463 = n21458 & ~n21461;
  assign n21464 = ~n21462 & ~n21463;
  assign n21465 = n20448 & ~n21464;
  assign n21466 = ~n20448 & n21464;
  assign n21467 = ~n21465 & ~n21466;
  assign n21468 = ~pi532 & ~n21467;
  assign po370 = n21455 | n21468;
  assign n21470 = pi532 & pi548;
  assign n21471 = ~pi156 & pi228;
  assign n21472 = pi156 & ~pi228;
  assign n21473 = ~n21471 & ~n21472;
  assign n21474 = ~pi224 & pi233;
  assign n21475 = pi224 & ~pi233;
  assign n21476 = ~n21474 & ~n21475;
  assign n21477 = ~n21473 & n21476;
  assign n21478 = n21473 & ~n21476;
  assign n21479 = ~n21477 & ~n21478;
  assign n21480 = n19589 & ~n21479;
  assign n21481 = ~n19589 & n21479;
  assign n21482 = ~n21480 & ~n21481;
  assign n21483 = ~pi532 & ~n21482;
  assign po371 = n21470 | n21483;
  assign n21485 = pi532 & pi541;
  assign n21486 = pi155 & ~pi230;
  assign n21487 = ~pi155 & pi230;
  assign n21488 = ~n21486 & ~n21487;
  assign n21489 = ~pi225 & pi234;
  assign n21490 = pi225 & ~pi234;
  assign n21491 = ~n21489 & ~n21490;
  assign n21492 = ~n21488 & n21491;
  assign n21493 = n21488 & ~n21491;
  assign n21494 = ~n21492 & ~n21493;
  assign n21495 = n19472 & ~n21494;
  assign n21496 = ~n19472 & n21494;
  assign n21497 = ~n21495 & ~n21496;
  assign n21498 = ~pi532 & ~n21497;
  assign po372 = n21485 | n21498;
  assign n21500 = pi129 & n15135;
  assign n21501 = ~pi129 & ~n15135;
  assign po373 = n21500 | n21501;
  assign n21503 = pi121 & n7299;
  assign n21504 = ~pi121 & ~n7299;
  assign po374 = n21503 | n21504;
  assign n21506 = pi179 & n10961;
  assign n21507 = ~pi179 & ~n10961;
  assign po375 = n21506 | n21507;
  assign n21509 = pi280 & n4620;
  assign n21510 = ~pi280 & ~n4620;
  assign po376 = n21509 | n21510;
  assign n21512 = pi225 & n9162;
  assign n21513 = ~pi225 & ~n9162;
  assign po377 = n21512 | n21513;
  assign n21515 = ~pi226 & n12363;
  assign n21516 = pi226 & ~n12363;
  assign po378 = n21515 | n21516;
  assign n21518 = pi232 & n14315;
  assign n21519 = ~pi232 & ~n14315;
  assign po379 = n21518 | n21519;
  assign n21521 = pi130 & n8945;
  assign n21522 = ~pi130 & ~n8945;
  assign po380 = n21521 | n21522;
  assign n21524 = pi132 & n5603;
  assign n21525 = ~pi132 & ~n5603;
  assign po381 = n21524 | n21525;
  assign n21527 = pi156 & n1627;
  assign n21528 = ~pi156 & ~n1627;
  assign po382 = n21527 | n21528;
  assign n21530 = ~pi151 & ~n7605;
  assign n21531 = pi151 & n7605;
  assign po383 = n21530 | n21531;
  assign n21533 = pi228 & n11452;
  assign n21534 = ~pi228 & ~n11452;
  assign po384 = n21533 | n21534;
  assign n21536 = ~pi229 & ~n12768;
  assign n21537 = pi229 & n12768;
  assign po385 = n21536 | n21537;
  assign n21539 = pi319 & n9274;
  assign n21540 = ~pi319 & ~n9274;
  assign po386 = n21539 | n21540;
  assign n21542 = pi153 & n15268;
  assign n21543 = ~pi153 & ~n15268;
  assign po387 = n21542 | n21543;
  assign n21545 = ~pi146 & n15749;
  assign n21546 = pi146 & ~n15749;
  assign po388 = n21545 | n21546;
  assign n21548 = pi256 & n13987;
  assign n21549 = ~pi256 & ~n13987;
  assign po389 = n21548 | n21549;
  assign n21551 = pi227 & n15564;
  assign n21552 = ~pi227 & ~n15564;
  assign po390 = n21551 | n21552;
  assign n21554 = pi303 & n13204;
  assign n21555 = ~pi303 & ~n13204;
  assign po391 = n21554 | n21555;
  assign n21557 = pi255 & n13345;
  assign n21558 = ~pi255 & ~n13345;
  assign po392 = n21557 | n21558;
  assign n21560 = ~pi255 & n20679;
  assign n21561 = pi255 & ~n20679;
  assign n21562 = ~n21560 & ~n21561;
  assign n21563 = pi384 & n21562;
  assign n21564 = ~pi384 & ~n21562;
  assign n21565 = ~n21563 & ~n21564;
  assign n21566 = ~pi532 & ~n21565;
  assign n21567 = pi532 & pi657;
  assign po393 = n21566 | n21567;
  assign n21569 = pi532 & pi643;
  assign n21570 = pi256 & n19241;
  assign n21571 = ~pi256 & ~n19241;
  assign n21572 = ~n21570 & ~n21571;
  assign n21573 = ~pi532 & ~n21572;
  assign po394 = n21569 | n21573;
  assign n21575 = ~pi257 & pi376;
  assign n21576 = pi257 & ~pi376;
  assign n21577 = ~n21575 & ~n21576;
  assign n21578 = n18534 & n18573;
  assign n21579 = ~n18720 & ~n21578;
  assign n21580 = pi138 & n20493;
  assign n21581 = ~n18718 & ~n21580;
  assign n21582 = ~n20021 & n21581;
  assign n21583 = n20062 & ~n21582;
  assign n21584 = ~pi138 & n18499;
  assign n21585 = ~n18594 & ~n21584;
  assign n21586 = ~n18456 & n21585;
  assign n21587 = n18971 & ~n21586;
  assign n21588 = ~n18479 & ~n18688;
  assign n21589 = pi138 & n18490;
  assign n21590 = ~n18482 & ~n21589;
  assign n21591 = ~n18954 & n21590;
  assign n21592 = ~pi207 & ~n21591;
  assign n21593 = n21588 & ~n21592;
  assign n21594 = ~pi302 & ~n21593;
  assign n21595 = ~n21587 & ~n21594;
  assign n21596 = ~n21583 & n21595;
  assign n21597 = pi138 & n18672;
  assign n21598 = ~n18539 & ~n18573;
  assign n21599 = ~pi207 & ~n21598;
  assign n21600 = n18585 & n20525;
  assign n21601 = ~n21599 & ~n21600;
  assign n21602 = ~n21597 & n21601;
  assign n21603 = ~n20076 & n21602;
  assign n21604 = pi302 & ~n21603;
  assign n21605 = n21596 & ~n21604;
  assign n21606 = n18489 & n18561;
  assign n21607 = ~n18550 & ~n21606;
  assign n21608 = ~pi207 & n20069;
  assign n21609 = ~n18732 & ~n21100;
  assign n21610 = ~n18741 & ~n20008;
  assign n21611 = n21609 & n21610;
  assign n21612 = ~n20520 & n21611;
  assign n21613 = ~n21608 & n21612;
  assign n21614 = ~pi302 & ~n21613;
  assign n21615 = ~pi138 & n18454;
  assign n21616 = ~n18523 & ~n21615;
  assign n21617 = pi207 & ~n21616;
  assign n21618 = ~pi138 & ~n18469;
  assign n21619 = pi138 & ~n20518;
  assign n21620 = ~n21618 & ~n21619;
  assign n21621 = ~n18460 & ~n21620;
  assign n21622 = ~pi207 & ~n21621;
  assign n21623 = n18448 & ~n18542;
  assign n21624 = ~n21622 & n21623;
  assign n21625 = ~n21617 & n21624;
  assign n21626 = pi302 & ~n21625;
  assign n21627 = ~n21614 & ~n21626;
  assign n21628 = ~n18683 & n21627;
  assign n21629 = ~n18612 & n21628;
  assign n21630 = n21607 & n21629;
  assign n21631 = ~n18594 & ~n20521;
  assign n21632 = n21630 & n21631;
  assign n21633 = ~pi139 & ~n21632;
  assign n21634 = ~n18478 & ~n18961;
  assign n21635 = ~n18491 & n21634;
  assign n21636 = ~n20009 & n21635;
  assign n21637 = ~pi207 & ~n21636;
  assign n21638 = ~pi138 & n18478;
  assign n21639 = ~n21637 & ~n21638;
  assign n21640 = pi207 & n18521;
  assign n21641 = ~pi207 & n18530;
  assign n21642 = ~pi138 & n18541;
  assign n21643 = ~n21641 & ~n21642;
  assign n21644 = n18449 & n18493;
  assign n21645 = ~n18707 & ~n21644;
  assign n21646 = ~n18491 & n21645;
  assign n21647 = n21643 & n21646;
  assign n21648 = ~pi302 & ~n21647;
  assign n21649 = ~n21640 & ~n21648;
  assign n21650 = ~n20021 & n21649;
  assign n21651 = n21639 & n21650;
  assign n21652 = ~n18571 & ~n18646;
  assign n21653 = ~n20518 & ~n21115;
  assign n21654 = ~n18632 & n21653;
  assign n21655 = pi207 & ~n21654;
  assign n21656 = n21652 & ~n21655;
  assign n21657 = pi302 & ~n21656;
  assign n21658 = n21651 & ~n21657;
  assign n21659 = pi139 & ~n21658;
  assign n21660 = ~n21633 & ~n21659;
  assign n21661 = n21605 & n21660;
  assign n21662 = n21579 & n21661;
  assign n21663 = pi373 & n21662;
  assign n21664 = ~pi373 & ~n21662;
  assign n21665 = ~n21663 & ~n21664;
  assign n21666 = ~n21577 & n21665;
  assign n21667 = n21577 & ~n21665;
  assign n21668 = ~n21666 & ~n21667;
  assign n21669 = ~pi532 & ~n21668;
  assign n21670 = pi532 & pi566;
  assign po395 = n21669 | n21670;
  assign n21672 = pi258 & ~pi370;
  assign n21673 = ~pi258 & pi370;
  assign n21674 = ~n21672 & ~n21673;
  assign n21675 = ~n18722 & ~n18989;
  assign n21676 = pi138 & n18443;
  assign n21677 = pi147 & ~pi185;
  assign n21678 = ~n21676 & ~n21677;
  assign n21679 = n21675 & n21678;
  assign n21680 = n20062 & ~n21679;
  assign n21681 = n18499 & n18585;
  assign n21682 = ~n20541 & ~n21681;
  assign n21683 = pi302 & ~n21682;
  assign n21684 = ~n21680 & ~n21683;
  assign n21685 = ~n18657 & ~n18722;
  assign n21686 = ~n20493 & n21685;
  assign n21687 = ~pi207 & ~n21686;
  assign n21688 = ~n18503 & ~n21687;
  assign n21689 = ~n18910 & ~n20526;
  assign n21690 = pi207 & n18633;
  assign n21691 = n21689 & ~n21690;
  assign n21692 = ~n18678 & n21691;
  assign n21693 = n21688 & n21692;
  assign n21694 = ~pi302 & ~n21693;
  assign n21695 = ~pi207 & n18910;
  assign n21696 = ~n21694 & ~n21695;
  assign n21697 = ~pi138 & n18570;
  assign n21698 = ~n18528 & ~n21697;
  assign n21699 = pi207 & ~n21698;
  assign n21700 = n18496 & n18534;
  assign n21701 = ~n21699 & ~n21700;
  assign n21702 = ~n18520 & n21701;
  assign n21703 = ~n18951 & n21702;
  assign n21704 = n21696 & n21703;
  assign n21705 = n21684 & n21704;
  assign n21706 = pi139 & ~n21705;
  assign n21707 = n18534 & n18669;
  assign n21708 = ~n20492 & ~n21707;
  assign n21709 = ~n18954 & n21708;
  assign n21710 = ~pi302 & ~n21709;
  assign n21711 = ~pi185 & ~pi207;
  assign n21712 = pi166 & ~pi302;
  assign n21713 = n21711 & n21712;
  assign n21714 = ~n21710 & ~n21713;
  assign n21715 = pi207 & n18646;
  assign n21716 = ~n21578 & ~n21715;
  assign n21717 = ~n18612 & n21716;
  assign n21718 = n18489 & n20518;
  assign n21719 = pi138 & ~pi147;
  assign n21720 = pi185 & n21719;
  assign n21721 = ~n21589 & ~n21720;
  assign n21722 = ~pi207 & ~n21721;
  assign n21723 = ~n20009 & ~n20021;
  assign n21724 = ~n21722 & n21723;
  assign n21725 = ~n21718 & n21724;
  assign n21726 = pi302 & ~n21725;
  assign n21727 = n21717 & ~n21726;
  assign n21728 = ~n18942 & ~n21615;
  assign n21729 = ~pi207 & ~n21728;
  assign n21730 = ~pi207 & n18481;
  assign n21731 = ~n21729 & ~n21730;
  assign n21732 = ~n18590 & n21731;
  assign n21733 = n21727 & n21732;
  assign n21734 = n21714 & n21733;
  assign n21735 = ~pi139 & ~n21734;
  assign n21736 = ~n21706 & ~n21735;
  assign n21737 = ~n18542 & ~n20541;
  assign n21738 = n18971 & ~n21737;
  assign n21739 = ~pi138 & ~pi302;
  assign n21740 = n20494 & n21739;
  assign n21741 = ~n21738 & ~n21740;
  assign n21742 = ~pi207 & n20048;
  assign n21743 = ~n21729 & ~n21742;
  assign n21744 = ~n18679 & n21743;
  assign n21745 = ~pi302 & ~n21744;
  assign n21746 = n21741 & ~n21745;
  assign n21747 = ~n18540 & ~n20502;
  assign n21748 = ~pi207 & ~n21747;
  assign n21749 = n21746 & ~n21748;
  assign n21750 = pi138 & ~n18978;
  assign n21751 = ~n20046 & ~n21750;
  assign n21752 = ~n18595 & n21751;
  assign n21753 = ~pi207 & ~n21752;
  assign n21754 = ~n18445 & ~n18571;
  assign n21755 = ~n18553 & ~n18609;
  assign n21756 = ~n18570 & n21755;
  assign n21757 = ~pi138 & ~n21756;
  assign n21758 = n21754 & ~n21757;
  assign n21759 = pi207 & ~n21758;
  assign n21760 = ~n21753 & ~n21759;
  assign n21761 = pi302 & ~n21760;
  assign n21762 = n21749 & ~n21761;
  assign n21763 = n21736 & n21762;
  assign n21764 = pi348 & n21763;
  assign n21765 = ~pi348 & ~n21763;
  assign n21766 = ~n21764 & ~n21765;
  assign n21767 = ~n21674 & n21766;
  assign n21768 = n21674 & ~n21766;
  assign n21769 = ~n21767 & ~n21768;
  assign n21770 = ~pi532 & ~n21769;
  assign n21771 = pi532 & pi572;
  assign po396 = n21770 | n21771;
  assign n21773 = pi157 & n14762;
  assign n21774 = ~pi157 & ~n14762;
  assign po397 = n21773 | n21774;
  assign n21776 = pi160 & n5074;
  assign n21777 = ~pi160 & ~n5074;
  assign po398 = n21776 | n21777;
  assign n21779 = pi193 & n7192;
  assign n21780 = ~pi193 & ~n7192;
  assign po399 = n21779 | n21780;
  assign n21782 = ~pi170 & ~n14582;
  assign n21783 = pi170 & n14582;
  assign po400 = n21782 | n21783;
  assign n21785 = ~pi142 & ~n10453;
  assign n21786 = pi142 & n10453;
  assign po401 = n21785 | n21786;
  assign n21788 = pi143 & n2474;
  assign n21789 = ~pi143 & ~n2474;
  assign po402 = n21788 | n21789;
  assign n21791 = pi178 & ~n13072;
  assign n21792 = ~pi178 & n13072;
  assign po403 = n21791 | n21792;
  assign n21794 = pi180 & n11953;
  assign n21795 = ~pi180 & ~n11953;
  assign po404 = n21794 | n21795;
  assign n21797 = pi267 & ~pi303;
  assign n21798 = ~pi267 & pi303;
  assign n21799 = ~n21797 & ~n21798;
  assign n21800 = pi389 & n21799;
  assign n21801 = ~pi389 & ~n21799;
  assign n21802 = ~n21800 & ~n21801;
  assign n21803 = ~n18043 & ~n19786;
  assign n21804 = pi132 & n19733;
  assign n21805 = ~n18041 & ~n21804;
  assign n21806 = ~n18798 & n21805;
  assign n21807 = n18792 & ~n21806;
  assign n21808 = ~pi132 & n17661;
  assign n21809 = ~n17743 & ~n21808;
  assign n21810 = ~n17679 & n21809;
  assign n21811 = n18317 & ~n21810;
  assign n21812 = ~n17693 & ~n18014;
  assign n21813 = ~n17695 & ~n19775;
  assign n21814 = ~n18345 & n21813;
  assign n21815 = ~pi351 & ~n21814;
  assign n21816 = n21812 & ~n21815;
  assign n21817 = ~pi284 & ~n21816;
  assign n21818 = ~n21811 & ~n21817;
  assign n21819 = ~n21807 & n21818;
  assign n21820 = pi132 & n17998;
  assign n21821 = ~n17630 & ~n17642;
  assign n21822 = ~pi351 & ~n21821;
  assign n21823 = n17733 & n19741;
  assign n21824 = ~n21822 & ~n21823;
  assign n21825 = ~n21820 & n21824;
  assign n21826 = ~n18762 & n21825;
  assign n21827 = pi284 & ~n21826;
  assign n21828 = n21819 & ~n21827;
  assign n21829 = n17601 & n17702;
  assign n21830 = ~n17656 & ~n21829;
  assign n21831 = ~pi351 & n18777;
  assign n21832 = ~n18055 & ~n20849;
  assign n21833 = ~n18065 & ~n18839;
  assign n21834 = n21832 & n21833;
  assign n21835 = ~n20625 & n21834;
  assign n21836 = ~n21831 & n21835;
  assign n21837 = ~pi284 & ~n21836;
  assign n21838 = ~n17593 & ~n19758;
  assign n21839 = pi351 & ~n21838;
  assign n21840 = ~pi132 & ~n17610;
  assign n21841 = pi132 & ~n19778;
  assign n21842 = ~n21840 & ~n21841;
  assign n21843 = ~n17659 & ~n21842;
  assign n21844 = ~pi351 & ~n21843;
  assign n21845 = ~n17635 & n17673;
  assign n21846 = ~n21844 & n21845;
  assign n21847 = ~n21839 & n21846;
  assign n21848 = pi284 & ~n21847;
  assign n21849 = ~n21837 & ~n21848;
  assign n21850 = ~n18009 & n21849;
  assign n21851 = ~n17761 & n21850;
  assign n21852 = n21830 & n21851;
  assign n21853 = ~n17743 & ~n20626;
  assign n21854 = n21852 & n21853;
  assign n21855 = ~pi193 & ~n21854;
  assign n21856 = ~n17692 & ~n18360;
  assign n21857 = ~n18836 & n21856;
  assign n21858 = ~n17703 & n21857;
  assign n21859 = ~pi351 & ~n21858;
  assign n21860 = ~pi132 & n17692;
  assign n21861 = ~n21859 & ~n21860;
  assign n21862 = pi351 & n17622;
  assign n21863 = ~pi351 & n17611;
  assign n21864 = ~pi132 & n17633;
  assign n21865 = ~n21863 & ~n21864;
  assign n21866 = n17674 & n17705;
  assign n21867 = ~n18034 & ~n21866;
  assign n21868 = ~n17703 & n21867;
  assign n21869 = n21865 & n21868;
  assign n21870 = ~pi284 & ~n21869;
  assign n21871 = ~n21862 & ~n21870;
  assign n21872 = ~n18798 & n21871;
  assign n21873 = n21861 & n21872;
  assign n21874 = ~n17640 & ~n17973;
  assign n21875 = ~n17963 & ~n19778;
  assign n21876 = ~n20860 & n21875;
  assign n21877 = pi351 & ~n21876;
  assign n21878 = n21874 & ~n21877;
  assign n21879 = pi284 & ~n21878;
  assign n21880 = n21873 & ~n21879;
  assign n21881 = pi193 & ~n21880;
  assign n21882 = ~n21855 & ~n21881;
  assign n21883 = n21828 & n21882;
  assign n21884 = n21803 & n21883;
  assign n21885 = ~pi268 & n21884;
  assign n21886 = pi268 & ~n21884;
  assign n21887 = ~n21885 & ~n21886;
  assign n21888 = ~n21802 & n21887;
  assign n21889 = n21802 & ~n21887;
  assign n21890 = ~n21888 & ~n21889;
  assign n21891 = ~pi532 & ~n21890;
  assign n21892 = pi532 & pi590;
  assign po405 = n21891 | n21892;
  assign n21894 = pi532 & pi622;
  assign n21895 = ~pi268 & ~pi303;
  assign n21896 = pi268 & pi303;
  assign n21897 = ~n21895 & ~n21896;
  assign n21898 = pi389 & n21884;
  assign n21899 = ~pi389 & ~n21884;
  assign n21900 = ~n21898 & ~n21899;
  assign n21901 = ~n21897 & n21900;
  assign n21902 = n21897 & ~n21900;
  assign n21903 = ~n21901 & ~n21902;
  assign n21904 = ~pi532 & ~n21903;
  assign po406 = n21894 | n21904;
  assign n21906 = pi269 & n19703;
  assign n21907 = ~pi269 & ~n19703;
  assign n21908 = ~n21906 & ~n21907;
  assign n21909 = ~pi532 & ~n21908;
  assign n21910 = pi532 & pi641;
  assign po407 = n21909 | n21910;
  assign n21912 = pi159 & ~pi301;
  assign n21913 = ~pi159 & pi301;
  assign n21914 = ~n21912 & ~n21913;
  assign n21915 = ~pi269 & pi270;
  assign n21916 = pi269 & ~pi270;
  assign n21917 = ~n21915 & ~n21916;
  assign n21918 = ~n21914 & n21917;
  assign n21919 = n21914 & ~n21917;
  assign n21920 = ~n21918 & ~n21919;
  assign n21921 = n19703 & ~n21920;
  assign n21922 = ~n19703 & n21920;
  assign n21923 = ~n21921 & ~n21922;
  assign n21924 = ~pi532 & ~n21923;
  assign n21925 = pi532 & pi545;
  assign po408 = n21924 | n21925;
  assign n21927 = pi271 & n19993;
  assign n21928 = ~pi271 & ~n19993;
  assign n21929 = ~n21927 & ~n21928;
  assign n21930 = ~pi532 & ~n21929;
  assign n21931 = pi532 & pi651;
  assign po409 = n21930 | n21931;
  assign n21933 = pi532 & pi635;
  assign n21934 = pi272 & n20097;
  assign n21935 = ~pi272 & ~n20097;
  assign n21936 = ~n21934 & ~n21935;
  assign n21937 = ~pi532 & ~n21936;
  assign po410 = n21933 | n21937;
  assign n21939 = pi532 & pi619;
  assign n21940 = ~pi271 & pi273;
  assign n21941 = pi271 & ~pi273;
  assign n21942 = ~n21940 & ~n21941;
  assign n21943 = n19993 & ~n21942;
  assign n21944 = ~n19993 & n21942;
  assign n21945 = ~n21943 & ~n21944;
  assign n21946 = ~pi532 & ~n21945;
  assign po411 = n21939 | n21946;
  assign n21948 = pi532 & pi603;
  assign n21949 = ~pi272 & pi274;
  assign n21950 = pi272 & ~pi274;
  assign n21951 = ~n21949 & ~n21950;
  assign n21952 = n20097 & ~n21951;
  assign n21953 = ~n20097 & n21951;
  assign n21954 = ~n21952 & ~n21953;
  assign n21955 = ~pi532 & ~n21954;
  assign po412 = n21948 | n21955;
  assign n21957 = pi532 & pi555;
  assign n21958 = pi168 & ~pi273;
  assign n21959 = ~pi168 & pi273;
  assign n21960 = ~n21958 & ~n21959;
  assign n21961 = ~pi271 & pi275;
  assign n21962 = pi271 & ~pi275;
  assign n21963 = ~n21961 & ~n21962;
  assign n21964 = ~n21960 & n21963;
  assign n21965 = n21960 & ~n21963;
  assign n21966 = ~n21964 & ~n21965;
  assign n21967 = n19993 & ~n21966;
  assign n21968 = ~n19993 & n21966;
  assign n21969 = ~n21967 & ~n21968;
  assign n21970 = ~pi532 & ~n21969;
  assign po413 = n21957 | n21970;
  assign n21972 = pi532 & pi539;
  assign n21973 = pi169 & ~pi274;
  assign n21974 = ~pi169 & pi274;
  assign n21975 = ~n21973 & ~n21974;
  assign n21976 = ~pi272 & pi276;
  assign n21977 = pi272 & ~pi276;
  assign n21978 = ~n21976 & ~n21977;
  assign n21979 = ~n21975 & n21978;
  assign n21980 = n21975 & ~n21978;
  assign n21981 = ~n21979 & ~n21980;
  assign n21982 = n20097 & ~n21981;
  assign n21983 = ~n20097 & n21981;
  assign n21984 = ~n21982 & ~n21983;
  assign n21985 = ~pi532 & ~n21984;
  assign po414 = n21972 | n21985;
  assign n21987 = pi164 & n3040;
  assign n21988 = ~pi164 & ~n3040;
  assign po415 = n21987 | n21988;
  assign n21990 = pi278 & n20231;
  assign n21991 = ~pi278 & ~n20231;
  assign n21992 = ~n21990 & ~n21991;
  assign n21993 = ~pi532 & ~n21992;
  assign n21994 = pi532 & pi646;
  assign po416 = n21993 | n21994;
  assign n21996 = pi162 & n4042;
  assign n21997 = ~pi162 & ~n4042;
  assign po417 = n21996 | n21997;
  assign n21999 = pi532 & pi638;
  assign n22000 = pi280 & n20326;
  assign n22001 = ~pi280 & ~n20326;
  assign n22002 = ~n22000 & ~n22001;
  assign n22003 = ~pi532 & ~n22002;
  assign po418 = n21999 | n22003;
  assign n22005 = ~pi278 & pi281;
  assign n22006 = pi278 & ~pi281;
  assign n22007 = ~n22005 & ~n22006;
  assign n22008 = n20231 & ~n22007;
  assign n22009 = ~n20231 & n22007;
  assign n22010 = ~n22008 & ~n22009;
  assign n22011 = ~pi532 & ~n22010;
  assign n22012 = pi532 & pi614;
  assign po419 = n22011 | n22012;
  assign n22014 = pi133 & n10001;
  assign n22015 = ~pi133 & ~n10001;
  assign po420 = n22014 | n22015;
  assign n22017 = pi532 & pi606;
  assign n22018 = ~pi280 & pi283;
  assign n22019 = pi280 & ~pi283;
  assign n22020 = ~n22018 & ~n22019;
  assign n22021 = n20326 & ~n22020;
  assign n22022 = ~n20326 & n22020;
  assign n22023 = ~n22021 & ~n22022;
  assign n22024 = ~pi532 & ~n22023;
  assign po421 = n22017 | n22024;
  assign n22026 = pi173 & ~pi281;
  assign n22027 = ~pi173 & pi281;
  assign n22028 = ~n22026 & ~n22027;
  assign n22029 = ~pi278 & pi284;
  assign n22030 = pi278 & ~pi284;
  assign n22031 = ~n22029 & ~n22030;
  assign n22032 = ~n22028 & n22031;
  assign n22033 = n22028 & ~n22031;
  assign n22034 = ~n22032 & ~n22033;
  assign n22035 = n20231 & ~n22034;
  assign n22036 = ~n20231 & n22034;
  assign n22037 = ~n22035 & ~n22036;
  assign n22038 = ~pi532 & ~n22037;
  assign n22039 = pi532 & pi550;
  assign po422 = n22038 | n22039;
  assign n22041 = pi532 & pi542;
  assign n22042 = pi174 & ~pi283;
  assign n22043 = ~pi174 & pi283;
  assign n22044 = ~n22042 & ~n22043;
  assign n22045 = ~pi280 & pi285;
  assign n22046 = pi280 & ~pi285;
  assign n22047 = ~n22045 & ~n22046;
  assign n22048 = ~n22044 & n22047;
  assign n22049 = n22044 & ~n22047;
  assign n22050 = ~n22048 & ~n22049;
  assign n22051 = n20326 & ~n22050;
  assign n22052 = ~n20326 & n22050;
  assign n22053 = ~n22051 & ~n22052;
  assign n22054 = ~pi532 & ~n22053;
  assign po423 = n22041 | n22054;
  assign n22056 = ~pi149 & n12462;
  assign n22057 = pi149 & ~n12462;
  assign po424 = n22056 | n22057;
  assign n22059 = ~pi131 & n12057;
  assign n22060 = pi131 & ~n12057;
  assign po425 = n22059 | n22060;
  assign n22062 = pi139 & n7001;
  assign n22063 = ~pi139 & ~n7001;
  assign po426 = n22062 | n22063;
  assign n22065 = pi172 & n11545;
  assign n22066 = ~pi172 & ~n11545;
  assign po427 = n22065 | n22066;
  assign n22068 = pi134 & n9054;
  assign n22069 = ~pi134 & ~n9054;
  assign po428 = n22068 | n22069;
  assign n22071 = pi283 & n3591;
  assign n22072 = ~pi283 & ~n3591;
  assign po429 = n22071 | n22072;
  assign n22074 = pi222 & n8848;
  assign n22075 = ~pi222 & ~n8848;
  assign po430 = n22074 | n22075;
  assign n22077 = pi346 & n15917;
  assign n22078 = ~pi346 & ~n15917;
  assign po431 = n22077 | n22078;
  assign n22080 = pi147 & n14485;
  assign n22081 = ~pi147 & ~n14485;
  assign po432 = n22080 | n22081;
  assign n22083 = pi354 & n5484;
  assign n22084 = ~pi354 & ~n5484;
  assign po433 = n22083 | n22084;
  assign n22086 = pi351 & n6431;
  assign n22087 = ~pi351 & ~n6431;
  assign po434 = n22086 | n22087;
  assign n22089 = pi371 & n14085;
  assign n22090 = ~pi371 & ~n14085;
  assign po435 = n22089 | n22090;
  assign n22092 = pi267 & n11067;
  assign n22093 = ~pi267 & ~n11067;
  assign po436 = n22092 | n22093;
  assign n22095 = ~pi268 & n12661;
  assign n22096 = pi268 & ~n12661;
  assign po437 = n22095 | n22096;
  assign n22098 = pi221 & n1915;
  assign n22099 = ~pi221 & ~n1915;
  assign po438 = n22098 | n22099;
  assign n22101 = ~pi269 & pi301;
  assign n22102 = pi269 & ~pi301;
  assign n22103 = ~n22101 & ~n22102;
  assign n22104 = n19703 & ~n22103;
  assign n22105 = ~n19703 & n22103;
  assign n22106 = ~n22104 & ~n22105;
  assign n22107 = ~pi532 & ~n22106;
  assign n22108 = pi532 & pi609;
  assign po439 = n22107 | n22108;
  assign n22110 = pi532 & pi558;
  assign n22111 = ~pi267 & ~pi268;
  assign n22112 = pi267 & pi268;
  assign n22113 = ~n22111 & ~n22112;
  assign n22114 = pi302 & ~pi303;
  assign n22115 = ~pi302 & pi303;
  assign n22116 = ~n22114 & ~n22115;
  assign n22117 = ~n22113 & n22116;
  assign n22118 = n22113 & ~n22116;
  assign n22119 = ~n22117 & ~n22118;
  assign n22120 = n21900 & ~n22119;
  assign n22121 = ~n21900 & n22119;
  assign n22122 = ~n22120 & ~n22121;
  assign n22123 = ~pi532 & ~n22122;
  assign po440 = n22110 | n22123;
  assign n22125 = pi303 & n21884;
  assign n22126 = ~pi303 & ~n21884;
  assign n22127 = ~n22125 & ~n22126;
  assign n22128 = pi389 & n22127;
  assign n22129 = ~pi389 & ~n22127;
  assign n22130 = ~n22128 & ~n22129;
  assign n22131 = ~pi532 & ~n22130;
  assign n22132 = pi532 & pi654;
  assign po441 = n22131 | n22132;
  assign n22134 = pi174 & n2689;
  assign n22135 = ~pi174 & ~n2689;
  assign po442 = n22134 | n22135;
  assign n22137 = pi372 & n10853;
  assign n22138 = ~pi372 & ~n10853;
  assign po443 = n22137 | n22138;
  assign n22140 = ~pi342 & ~n6906;
  assign n22141 = pi342 & n6906;
  assign po444 = n22140 | n22141;
  assign n22143 = pi169 & n10182;
  assign n22144 = ~pi169 & ~n10182;
  assign po445 = n22143 | n22144;
  assign n22146 = pi183 & n2243;
  assign n22147 = ~pi183 & ~n2243;
  assign po446 = n22146 | n22147;
  assign n22149 = pi257 & n2586;
  assign n22150 = ~pi257 & ~n2586;
  assign po447 = n22149 | n22150;
  assign n22152 = ~pi258 & ~n2365;
  assign n22153 = pi258 & n2365;
  assign po448 = n22152 | n22153;
  assign n22155 = pi320 & n11853;
  assign n22156 = ~pi320 & ~n11853;
  assign po449 = n22155 | n22156;
  assign n22158 = pi274 & n15646;
  assign n22159 = ~pi274 & ~n15646;
  assign po450 = n22158 | n22159;
  assign n22161 = ~pi348 & ~n8140;
  assign n22162 = pi348 & n8140;
  assign po451 = n22161 | n22162;
  assign n22164 = pi217 & n7691;
  assign n22165 = ~pi217 & ~n7691;
  assign po452 = n22164 | n22165;
  assign n22167 = pi136 & n7402;
  assign n22168 = ~pi136 & ~n7402;
  assign po453 = n22167 | n22168;
  assign n22170 = ~pi135 & n12160;
  assign n22171 = pi135 & ~n12160;
  assign po454 = n22170 | n22171;
  assign n22173 = pi155 & n7988;
  assign n22174 = ~pi155 & ~n7988;
  assign po455 = n22173 | n22174;
  assign n22176 = pi230 & n8263;
  assign n22177 = ~pi230 & ~n8263;
  assign po456 = n22176 | n22177;
  assign n22179 = pi319 & n20582;
  assign n22180 = ~pi319 & ~n20582;
  assign n22181 = ~n22179 & ~n22180;
  assign n22182 = ~pi532 & ~n22181;
  assign n22183 = pi532 & pi633;
  assign po457 = n22182 | n22183;
  assign n22185 = pi319 & ~pi320;
  assign n22186 = ~pi319 & pi320;
  assign n22187 = ~n22185 & ~n22186;
  assign n22188 = n20582 & ~n22187;
  assign n22189 = ~n20582 & n22187;
  assign n22190 = ~n22188 & ~n22189;
  assign n22191 = ~pi532 & ~n22190;
  assign n22192 = pi532 & pi601;
  assign po458 = n22191 | n22192;
  assign n22194 = pi183 & ~pi320;
  assign n22195 = ~pi183 & pi320;
  assign n22196 = ~n22194 & ~n22195;
  assign n22197 = ~pi319 & pi321;
  assign n22198 = pi319 & ~pi321;
  assign n22199 = ~n22197 & ~n22198;
  assign n22200 = ~n22196 & n22199;
  assign n22201 = n22196 & ~n22199;
  assign n22202 = ~n22200 & ~n22201;
  assign n22203 = n20582 & ~n22202;
  assign n22204 = ~n20582 & n22202;
  assign n22205 = ~n22203 & ~n22204;
  assign n22206 = ~pi532 & ~n22205;
  assign n22207 = pi532 & pi537;
  assign po459 = n22206 | n22207;
  assign n22209 = pi285 & n10760;
  assign n22210 = ~pi285 & ~n10760;
  assign po460 = n22209 | n22210;
  assign n22212 = pi166 & n5772;
  assign n22213 = ~pi166 & ~n5772;
  assign po461 = n22212 | n22213;
  assign n22215 = ~pi272 & ~n16400;
  assign n22216 = pi272 & n16400;
  assign po462 = n22215 | n22216;
  assign n22218 = pi219 & n3238;
  assign n22219 = ~pi219 & ~n3238;
  assign po463 = n22218 | n22219;
  assign n22221 = pi168 & n10264;
  assign n22222 = ~pi168 & ~n10264;
  assign po464 = n22221 | n22222;
  assign n22224 = ~pi208 & n16021;
  assign n22225 = pi208 & ~n16021;
  assign po465 = n22224 | n22225;
  assign n22227 = pi353 & n5298;
  assign n22228 = ~pi353 & ~n5298;
  assign po466 = n22227 | n22228;
  assign n22230 = pi275 & n14399;
  assign n22231 = ~pi275 & ~n14399;
  assign po467 = n22230 | n22231;
  assign n22233 = ~pi370 & ~n8423;
  assign n22234 = pi370 & n8423;
  assign po468 = n22233 | n22234;
  assign n22236 = pi233 & n9897;
  assign n22237 = ~pi233 & ~n9897;
  assign po469 = n22236 | n22237;
  assign n22239 = pi215 & n14846;
  assign n22240 = ~pi215 & ~n14846;
  assign po470 = n22239 | n22240;
  assign n22242 = ~pi184 & n11649;
  assign n22243 = pi184 & ~n11649;
  assign po471 = n22242 | n22243;
  assign n22245 = pi356 & n9366;
  assign n22246 = ~pi356 & ~n9366;
  assign po472 = n22245 | n22246;
  assign n22248 = pi350 & n12862;
  assign n22249 = ~pi350 & ~n12862;
  assign po473 = n22248 | n22249;
  assign n22251 = pi175 & n6659;
  assign n22252 = ~pi175 & ~n6659;
  assign po474 = n22251 | n22252;
  assign n22254 = pi218 & n7798;
  assign n22255 = ~pi218 & ~n7798;
  assign po475 = n22254 | n22255;
  assign n22257 = pi138 & n9779;
  assign n22258 = ~pi138 & ~n9779;
  assign po476 = n22257 | n22258;
  assign n22260 = pi352 & n9771;
  assign n22261 = ~pi352 & ~n9771;
  assign po477 = n22260 | n22261;
  assign n22263 = pi185 & n10561;
  assign n22264 = ~pi185 & ~n10561;
  assign po478 = n22263 | n22264;
  assign n22266 = pi302 & n14952;
  assign n22267 = ~pi302 & ~n14952;
  assign po479 = n22266 | n22267;
  assign n22269 = pi532 & pi540;
  assign n22270 = pi258 & ~pi348;
  assign n22271 = ~pi258 & pi348;
  assign n22272 = ~n22270 & ~n22271;
  assign n22273 = pi342 & ~pi370;
  assign n22274 = ~pi342 & pi370;
  assign n22275 = ~n22273 & ~n22274;
  assign n22276 = ~n22272 & n22275;
  assign n22277 = n22272 & ~n22275;
  assign n22278 = ~n22276 & ~n22277;
  assign n22279 = n21763 & ~n22278;
  assign n22280 = ~n21763 & n22278;
  assign n22281 = ~n22279 & ~n22280;
  assign n22282 = ~pi532 & ~n22281;
  assign po480 = n22269 | n22282;
  assign n22284 = pi209 & n7888;
  assign n22285 = ~pi209 & ~n7888;
  assign po481 = n22284 | n22285;
  assign n22287 = pi210 & n16263;
  assign n22288 = ~pi210 & ~n16263;
  assign po482 = n22287 | n22288;
  assign n22290 = pi182 & n6783;
  assign n22291 = ~pi182 & ~n6783;
  assign po483 = n22290 | n22291;
  assign n22293 = pi532 & pi615;
  assign n22294 = ~pi346 & pi371;
  assign n22295 = pi346 & ~pi371;
  assign n22296 = ~n22294 & ~n22295;
  assign n22297 = n21055 & ~n22296;
  assign n22298 = ~n21055 & n22296;
  assign n22299 = ~n22297 & ~n22298;
  assign n22300 = ~pi532 & ~n22299;
  assign po484 = n22293 | n22300;
  assign n22302 = pi373 & n3421;
  assign n22303 = ~pi373 & ~n3421;
  assign po485 = n22302 | n22303;
  assign n22305 = pi532 & pi604;
  assign n22306 = pi348 & ~pi370;
  assign n22307 = ~pi348 & pi370;
  assign n22308 = ~n22306 & ~n22307;
  assign n22309 = n21763 & ~n22308;
  assign n22310 = ~n21763 & n22308;
  assign n22311 = ~n22309 & ~n22310;
  assign n22312 = ~pi532 & ~n22311;
  assign po486 = n22305 | n22312;
  assign n22314 = pi532 & pi631;
  assign n22315 = pi349 & n21149;
  assign n22316 = ~pi349 & ~n21149;
  assign n22317 = ~n22315 & ~n22316;
  assign n22318 = ~pi532 & ~n22317;
  assign po487 = n22314 | n22318;
  assign n22320 = pi532 & pi599;
  assign n22321 = ~pi349 & pi350;
  assign n22322 = pi349 & ~pi350;
  assign n22323 = ~n22321 & ~n22322;
  assign n22324 = n21149 & ~n22323;
  assign n22325 = ~n21149 & n22323;
  assign n22326 = ~n22324 & ~n22325;
  assign n22327 = ~pi532 & ~n22326;
  assign po488 = n22320 | n22327;
  assign n22329 = pi532 & pi551;
  assign n22330 = pi217 & ~pi346;
  assign n22331 = ~pi217 & pi346;
  assign n22332 = ~n22330 & ~n22331;
  assign n22333 = pi351 & ~pi371;
  assign n22334 = ~pi351 & pi371;
  assign n22335 = ~n22333 & ~n22334;
  assign n22336 = ~n22332 & n22335;
  assign n22337 = n22332 & ~n22335;
  assign n22338 = ~n22336 & ~n22337;
  assign n22339 = n21055 & ~n22338;
  assign n22340 = ~n21055 & n22338;
  assign n22341 = ~n22339 & ~n22340;
  assign n22342 = ~pi532 & ~n22341;
  assign po489 = n22329 | n22342;
  assign n22344 = pi532 & pi535;
  assign n22345 = pi218 & ~pi350;
  assign n22346 = ~pi218 & pi350;
  assign n22347 = ~n22345 & ~n22346;
  assign n22348 = ~pi349 & pi352;
  assign n22349 = pi349 & ~pi352;
  assign n22350 = ~n22348 & ~n22349;
  assign n22351 = ~n22347 & n22350;
  assign n22352 = n22347 & ~n22350;
  assign n22353 = ~n22351 & ~n22352;
  assign n22354 = n21149 & ~n22353;
  assign n22355 = ~n21149 & n22353;
  assign n22356 = ~n22354 & ~n22355;
  assign n22357 = ~pi532 & ~n22356;
  assign po490 = n22344 | n22357;
  assign n22359 = pi532 & pi652;
  assign n22360 = pi353 & n21253;
  assign n22361 = ~pi353 & ~n21253;
  assign n22362 = ~n22360 & ~n22361;
  assign n22363 = ~pi532 & ~n22362;
  assign po491 = n22359 | n22363;
  assign n22365 = pi532 & pi556;
  assign n22366 = ~pi219 & pi375;
  assign n22367 = pi219 & ~pi375;
  assign n22368 = ~n22366 & ~n22367;
  assign n22369 = ~pi353 & pi354;
  assign n22370 = pi353 & ~pi354;
  assign n22371 = ~n22369 & ~n22370;
  assign n22372 = ~n22368 & n22371;
  assign n22373 = n22368 & ~n22371;
  assign n22374 = ~n22372 & ~n22373;
  assign n22375 = n21253 & ~n22374;
  assign n22376 = ~n21253 & n22374;
  assign n22377 = ~n22375 & ~n22376;
  assign n22378 = ~pi532 & ~n22377;
  assign po492 = n22365 | n22378;
  assign n22380 = pi171 & n14175;
  assign n22381 = ~pi171 & ~n14175;
  assign po493 = n22380 | n22381;
  assign n22383 = pi532 & pi649;
  assign n22384 = pi356 & n21346;
  assign n22385 = ~pi356 & ~n21346;
  assign n22386 = ~n22384 & ~n22385;
  assign n22387 = ~pi532 & ~n22386;
  assign po494 = n22383 | n22387;
  assign n22389 = pi532 & pi617;
  assign n22390 = ~pi356 & pi357;
  assign n22391 = pi356 & ~pi357;
  assign n22392 = ~n22390 & ~n22391;
  assign n22393 = n21346 & ~n22392;
  assign n22394 = ~n21346 & n22392;
  assign n22395 = ~n22393 & ~n22394;
  assign n22396 = ~pi532 & ~n22395;
  assign po495 = n22389 | n22396;
  assign n22398 = pi532 & pi553;
  assign n22399 = pi220 & ~pi357;
  assign n22400 = ~pi220 & pi357;
  assign n22401 = ~n22399 & ~n22400;
  assign n22402 = ~pi356 & pi358;
  assign n22403 = pi356 & ~pi358;
  assign n22404 = ~n22402 & ~n22403;
  assign n22405 = ~n22401 & n22404;
  assign n22406 = n22401 & ~n22404;
  assign n22407 = ~n22405 & ~n22406;
  assign n22408 = n21346 & ~n22407;
  assign n22409 = ~n21346 & n22407;
  assign n22410 = ~n22408 & ~n22409;
  assign n22411 = ~pi532 & ~n22410;
  assign po496 = n22398 | n22411;
  assign n22413 = pi376 & n4451;
  assign n22414 = ~pi376 & ~n4451;
  assign po497 = n22413 | n22414;
  assign n22416 = pi165 & n2937;
  assign n22417 = ~pi165 & ~n2937;
  assign po498 = n22416 | n22417;
  assign n22419 = pi187 & n9554;
  assign n22420 = ~pi187 & ~n9554;
  assign po499 = n22419 | n22420;
  assign n22422 = pi278 & n4786;
  assign n22423 = ~pi278 & ~n4786;
  assign po500 = n22422 | n22423;
  assign n22425 = pi161 & n4957;
  assign n22426 = ~pi161 & ~n4957;
  assign po501 = n22425 | n22426;
  assign n22428 = pi271 & n13723;
  assign n22429 = ~pi271 & ~n13723;
  assign po502 = n22428 | n22429;
  assign n22431 = pi207 & n6533;
  assign n22432 = ~pi207 & ~n6533;
  assign po503 = n22431 | n22432;
  assign n22434 = ~pi349 & ~n8521;
  assign n22435 = pi349 & n8521;
  assign po504 = n22434 | n22435;
  assign n22437 = pi220 & n2078;
  assign n22438 = ~pi220 & ~n2078;
  assign po505 = n22437 | n22438;
  assign n22440 = pi357 & n11744;
  assign n22441 = ~pi357 & ~n11744;
  assign po506 = n22440 | n22441;
  assign n22443 = ~pi163 & n3926;
  assign n22444 = pi163 & ~n3926;
  assign po507 = n22443 | n22444;
  assign n22446 = pi532 & pi636;
  assign n22447 = pi370 & n21763;
  assign n22448 = ~pi370 & ~n21763;
  assign n22449 = ~n22447 & ~n22448;
  assign n22450 = ~pi532 & ~n22449;
  assign po508 = n22446 | n22450;
  assign n22452 = pi532 & pi647;
  assign n22453 = pi371 & n21055;
  assign n22454 = ~pi371 & ~n21055;
  assign n22455 = ~n22453 & ~n22454;
  assign n22456 = ~pi532 & ~n22455;
  assign po509 = n22452 | n22456;
  assign n22458 = pi257 & ~pi373;
  assign n22459 = ~pi257 & pi373;
  assign n22460 = ~n22458 & ~n22459;
  assign n22461 = pi372 & ~pi376;
  assign n22462 = ~pi372 & pi376;
  assign n22463 = ~n22461 & ~n22462;
  assign n22464 = ~n22460 & n22463;
  assign n22465 = n22460 & ~n22463;
  assign n22466 = ~n22464 & ~n22465;
  assign n22467 = n21662 & ~n22466;
  assign n22468 = ~n21662 & n22466;
  assign n22469 = ~n22467 & ~n22468;
  assign n22470 = ~pi532 & ~n22469;
  assign n22471 = pi532 & pi534;
  assign po510 = n22470 | n22471;
  assign n22473 = pi373 & ~pi376;
  assign n22474 = ~pi373 & pi376;
  assign n22475 = ~n22473 & ~n22474;
  assign n22476 = n21662 & ~n22475;
  assign n22477 = ~n21662 & n22475;
  assign n22478 = ~n22476 & ~n22477;
  assign n22479 = ~pi532 & ~n22478;
  assign n22480 = pi532 & pi598;
  assign po511 = n22479 | n22480;
  assign n22482 = pi358 & n6163;
  assign n22483 = ~pi358 & ~n6163;
  assign po512 = n22482 | n22483;
  assign n22485 = pi532 & pi620;
  assign n22486 = pi353 & ~pi375;
  assign n22487 = ~pi353 & pi375;
  assign n22488 = ~n22486 & ~n22487;
  assign n22489 = n21253 & ~n22488;
  assign n22490 = ~n21253 & n22488;
  assign n22491 = ~n22489 & ~n22490;
  assign n22492 = ~pi532 & ~n22491;
  assign po513 = n22485 | n22492;
  assign n22494 = pi376 & n21662;
  assign n22495 = ~pi376 & ~n21662;
  assign n22496 = ~n22494 & ~n22495;
  assign n22497 = ~pi532 & ~n22496;
  assign n22498 = pi532 & pi630;
  assign po514 = n22497 | n22498;
  assign n22500 = pi273 & n15484;
  assign n22501 = ~pi273 & ~n15484;
  assign po515 = n22500 | n22501;
  assign n22503 = pi281 & n3755;
  assign n22504 = ~pi281 & ~n3755;
  assign po516 = n22503 | n22504;
  assign n22506 = pi181 & n8623;
  assign n22507 = ~pi181 & ~n8623;
  assign po517 = n22506 | n22507;
  assign n22509 = pi375 & n4267;
  assign n22510 = ~pi375 & ~n4267;
  assign po518 = n22509 | n22510;
  assign n22512 = pi284 & n10672;
  assign n22513 = ~pi284 & ~n10672;
  assign po519 = n22512 | n22513;
  assign n22515 = pi173 & n2811;
  assign n22516 = ~pi173 & ~n2811;
  assign po520 = n22515 | n22516;
  assign n22518 = pi234 & n7102;
  assign n22519 = ~pi234 & ~n7102;
  assign po521 = n22518 | n22519;
  assign n22521 = pi487 & pi520;
  assign n22522 = ~pi487 & ~pi520;
  assign n22523 = ~n22521 & ~n22522;
  assign n22524 = pi482 & n22521;
  assign n22525 = pi396 & ~n22524;
  assign n22526 = ~pi396 & n22524;
  assign n22527 = ~n22525 & ~n22526;
  assign n22528 = ~pi482 & ~n22521;
  assign n22529 = ~n22524 & ~n22528;
  assign n22530 = n22527 & n22529;
  assign n22531 = ~n22523 & n22530;
  assign n22532 = pi520 & n22531;
  assign n22533 = ~n22527 & ~n22529;
  assign n22534 = ~n22523 & n22533;
  assign n22535 = ~n22532 & ~n22534;
  assign po522 = ~pi532 & ~n22535;
  assign n22537 = ~pi520 & ~n22534;
  assign n22538 = n22527 & ~n22529;
  assign n22539 = n22523 & n22538;
  assign n22540 = pi520 & ~n22539;
  assign n22541 = ~n22537 & ~n22540;
  assign po523 = ~pi532 & n22541;
  assign n22543 = ~pi520 & ~n22539;
  assign n22544 = pi520 & ~n22534;
  assign n22545 = ~n22543 & ~n22544;
  assign po524 = ~pi532 & n22545;
  assign n22547 = pi531 & pi532;
  assign n22548 = ~pi393 & ~pi395;
  assign n22549 = ~pi387 & ~pi390;
  assign n22550 = n22548 & n22549;
  assign n22551 = ~pi390 & n22548;
  assign n22552 = pi387 & ~n22551;
  assign n22553 = ~n22550 & ~n22552;
  assign n22554 = ~n22550 & ~n22553;
  assign n22555 = pi387 & n22550;
  assign n22556 = ~n22554 & ~n22555;
  assign n22557 = pi531 & ~n22556;
  assign po525 = n22547 | n22557;
  assign po658 = ~pi520 & ~pi532;
  assign n22560 = ~n22531 & ~n22534;
  assign po526 = po658 & ~n22560;
  assign n22562 = ~pi520 & ~n22523;
  assign n22563 = ~n22529 & n22562;
  assign n22564 = ~n22534 & ~n22563;
  assign po527 = ~pi532 & ~n22564;
  assign n22566 = n22548 & ~n22550;
  assign n22567 = pi390 & ~n22566;
  assign n22568 = ~n22550 & n22551;
  assign n22569 = ~n22567 & ~n22568;
  assign n22570 = pi531 & ~n22569;
  assign po528 = ~pi532 & n22570;
  assign po625 = ~pi532 & n22523;
  assign n22573 = pi520 & po625;
  assign po529 = n22530 & n22573;
  assign n22575 = ~pi520 & po625;
  assign po530 = n22530 & n22575;
  assign n22577 = pi393 & pi395;
  assign n22578 = ~n22548 & ~n22577;
  assign n22579 = ~n22550 & ~n22578;
  assign n22580 = pi393 & n22550;
  assign n22581 = ~n22579 & ~n22580;
  assign n22582 = pi531 & ~n22581;
  assign po531 = n22547 | n22582;
  assign n22584 = pi520 & ~n22523;
  assign n22585 = ~n22529 & n22584;
  assign po532 = pi532 | n22585;
  assign n22587 = pi395 & ~n22550;
  assign n22588 = ~pi395 & n22550;
  assign n22589 = ~n22587 & ~n22588;
  assign n22590 = pi531 & n22589;
  assign po533 = n22547 | n22590;
  assign po534 = ~pi532 & ~n22527;
  assign n22593 = pi395 & n22549;
  assign n22594 = ~pi532 & n22593;
  assign po535 = ~pi393 & n22594;
  assign n22596 = pi398 & ~pi532;
  assign n22597 = pi532 & pi777;
  assign po536 = n22596 | n22597;
  assign n22599 = pi399 & ~pi532;
  assign n22600 = pi532 & pi772;
  assign po537 = n22599 | n22600;
  assign n22602 = pi400 & ~pi532;
  assign n22603 = pi532 & pi698;
  assign po538 = n22602 | n22603;
  assign n22605 = pi401 & ~pi532;
  assign n22606 = pi532 & pi675;
  assign po539 = n22605 | n22606;
  assign n22608 = pi402 & ~pi532;
  assign n22609 = pi532 & pi728;
  assign po540 = n22608 | n22609;
  assign n22611 = pi403 & ~pi532;
  assign n22612 = pi532 & pi708;
  assign po541 = n22611 | n22612;
  assign n22614 = pi404 & ~pi532;
  assign n22615 = pi532 & pi679;
  assign po542 = n22614 | n22615;
  assign n22617 = pi405 & ~pi532;
  assign n22618 = pi532 & pi661;
  assign po543 = n22617 | n22618;
  assign n22620 = pi406 & ~pi532;
  assign n22621 = pi532 & pi729;
  assign po544 = n22620 | n22621;
  assign n22623 = pi407 & ~pi532;
  assign n22624 = pi532 & pi710;
  assign po545 = n22623 | n22624;
  assign n22626 = pi408 & ~pi532;
  assign n22627 = pi532 & pi703;
  assign po546 = n22626 | n22627;
  assign n22629 = pi409 & ~pi532;
  assign n22630 = pi532 & pi788;
  assign po547 = n22629 | n22630;
  assign n22632 = pi410 & ~pi532;
  assign n22633 = pi532 & pi725;
  assign po548 = n22632 | n22633;
  assign n22635 = pi411 & ~pi532;
  assign n22636 = pi532 & pi715;
  assign po549 = n22635 | n22636;
  assign n22638 = pi412 & ~pi532;
  assign n22639 = pi532 & pi696;
  assign po550 = n22638 | n22639;
  assign n22641 = pi413 & ~pi532;
  assign n22642 = pi532 & pi667;
  assign po551 = n22641 | n22642;
  assign n22644 = pi414 & ~pi532;
  assign n22645 = pi532 & pi678;
  assign po552 = n22644 | n22645;
  assign n22647 = pi415 & ~pi532;
  assign n22648 = pi532 & pi769;
  assign po553 = n22647 | n22648;
  assign n22650 = pi416 & ~pi532;
  assign n22651 = pi532 & pi672;
  assign po554 = n22650 | n22651;
  assign n22653 = pi417 & ~pi532;
  assign n22654 = pi532 & pi784;
  assign po555 = n22653 | n22654;
  assign n22656 = pi418 & ~pi532;
  assign n22657 = pi532 & pi685;
  assign po556 = n22656 | n22657;
  assign n22659 = pi419 & ~pi532;
  assign n22660 = pi532 & pi687;
  assign po557 = n22659 | n22660;
  assign n22662 = pi420 & ~pi532;
  assign n22663 = pi532 & pi690;
  assign po558 = n22662 | n22663;
  assign n22665 = pi421 & ~pi532;
  assign n22666 = pi532 & pi707;
  assign po559 = n22665 | n22666;
  assign n22668 = pi422 & ~pi532;
  assign n22669 = pi532 & pi716;
  assign po560 = n22668 | n22669;
  assign n22671 = pi423 & ~pi532;
  assign n22672 = pi532 & pi722;
  assign po561 = n22671 | n22672;
  assign n22674 = pi424 & ~pi532;
  assign n22675 = pi532 & pi724;
  assign po562 = n22674 | n22675;
  assign n22677 = pi425 & ~pi532;
  assign n22678 = pi532 & pi739;
  assign po563 = n22677 | n22678;
  assign n22680 = pi426 & ~pi532;
  assign n22681 = pi532 & pi742;
  assign po564 = n22680 | n22681;
  assign n22683 = pi427 & ~pi532;
  assign n22684 = pi532 & pi747;
  assign po565 = n22683 | n22684;
  assign n22686 = pi428 & ~pi532;
  assign n22687 = pi532 & pi669;
  assign po566 = n22686 | n22687;
  assign n22689 = pi429 & ~pi532;
  assign n22690 = pi532 & pi760;
  assign po567 = n22689 | n22690;
  assign n22692 = pi430 & ~pi532;
  assign n22693 = pi532 & pi752;
  assign po568 = n22692 | n22693;
  assign n22695 = pi431 & ~pi532;
  assign n22696 = pi532 & pi700;
  assign po569 = n22695 | n22696;
  assign n22698 = pi432 & ~pi532;
  assign n22699 = pi532 & pi721;
  assign po570 = n22698 | n22699;
  assign n22701 = pi433 & ~pi532;
  assign n22702 = pi532 & pi764;
  assign po571 = n22701 | n22702;
  assign n22704 = pi434 & ~pi532;
  assign n22705 = pi532 & pi684;
  assign po572 = n22704 | n22705;
  assign n22707 = pi435 & ~pi532;
  assign n22708 = pi532 & pi719;
  assign po573 = n22707 | n22708;
  assign n22710 = pi436 & ~pi532;
  assign n22711 = pi532 & pi664;
  assign po574 = n22710 | n22711;
  assign n22713 = pi437 & ~pi532;
  assign n22714 = pi532 & pi779;
  assign po575 = n22713 | n22714;
  assign n22716 = pi438 & ~pi532;
  assign n22717 = pi532 & pi720;
  assign po576 = n22716 | n22717;
  assign n22719 = pi439 & ~pi532;
  assign n22720 = pi532 & pi757;
  assign po577 = n22719 | n22720;
  assign n22722 = pi440 & ~pi532;
  assign n22723 = pi532 & pi731;
  assign po578 = n22722 | n22723;
  assign n22725 = pi441 & ~pi532;
  assign n22726 = pi532 & pi712;
  assign po579 = n22725 | n22726;
  assign n22728 = pi442 & ~pi532;
  assign n22729 = pi532 & pi753;
  assign po580 = n22728 | n22729;
  assign n22731 = pi443 & ~pi532;
  assign n22732 = pi532 & pi768;
  assign po581 = n22731 | n22732;
  assign n22734 = pi444 & ~pi532;
  assign n22735 = pi532 & pi689;
  assign po582 = n22734 | n22735;
  assign n22737 = pi445 & ~pi532;
  assign n22738 = pi532 & pi738;
  assign po583 = n22737 | n22738;
  assign n22740 = pi446 & ~pi532;
  assign n22741 = pi532 & pi662;
  assign po584 = n22740 | n22741;
  assign n22743 = pi447 & ~pi532;
  assign n22744 = pi532 & pi680;
  assign po585 = n22743 | n22744;
  assign n22746 = pi448 & ~pi532;
  assign n22747 = pi532 & pi717;
  assign po586 = n22746 | n22747;
  assign n22749 = pi449 & ~pi532;
  assign n22750 = pi532 & pi751;
  assign po587 = n22749 | n22750;
  assign n22752 = pi450 & ~pi532;
  assign n22753 = pi532 & pi730;
  assign po588 = n22752 | n22753;
  assign n22755 = pi451 & ~pi532;
  assign n22756 = pi532 & pi673;
  assign po589 = n22755 | n22756;
  assign n22758 = pi452 & ~pi532;
  assign n22759 = pi532 & pi746;
  assign po590 = n22758 | n22759;
  assign n22761 = pi453 & ~pi532;
  assign n22762 = pi532 & pi741;
  assign po591 = n22761 | n22762;
  assign n22764 = pi454 & ~pi532;
  assign n22765 = pi532 & pi727;
  assign po592 = n22764 | n22765;
  assign n22767 = pi455 & ~pi532;
  assign n22768 = pi532 & pi670;
  assign po593 = n22767 | n22768;
  assign n22770 = pi456 & ~pi532;
  assign n22771 = pi532 & pi714;
  assign po594 = n22770 | n22771;
  assign n22773 = pi457 & ~pi532;
  assign n22774 = pi532 & pi706;
  assign po595 = n22773 | n22774;
  assign n22776 = pi458 & ~pi532;
  assign n22777 = pi532 & pi713;
  assign po596 = n22776 | n22777;
  assign n22779 = pi459 & ~pi532;
  assign n22780 = pi532 & pi758;
  assign po597 = n22779 | n22780;
  assign n22782 = pi460 & ~pi532;
  assign n22783 = pi532 & pi671;
  assign po598 = n22782 | n22783;
  assign n22785 = pi461 & ~pi532;
  assign n22786 = pi532 & pi695;
  assign po599 = n22785 | n22786;
  assign n22788 = pi462 & ~pi532;
  assign n22789 = pi532 & pi771;
  assign po600 = n22788 | n22789;
  assign n22791 = pi463 & ~pi532;
  assign n22792 = pi532 & pi691;
  assign po601 = n22791 | n22792;
  assign n22794 = pi464 & ~pi532;
  assign n22795 = pi532 & pi765;
  assign po602 = n22794 | n22795;
  assign n22797 = pi465 & ~pi532;
  assign n22798 = pi532 & pi726;
  assign po603 = n22797 | n22798;
  assign n22800 = pi466 & ~pi532;
  assign n22801 = pi532 & pi740;
  assign po604 = n22800 | n22801;
  assign n22803 = pi467 & ~pi532;
  assign n22804 = pi532 & pi668;
  assign po605 = n22803 | n22804;
  assign n22806 = pi468 & ~pi532;
  assign n22807 = pi532 & pi743;
  assign po606 = n22806 | n22807;
  assign n22809 = pi469 & ~pi532;
  assign n22810 = pi532 & pi787;
  assign po607 = n22809 | n22810;
  assign n22812 = pi470 & ~pi532;
  assign n22813 = pi532 & pi766;
  assign po608 = n22812 | n22813;
  assign n22815 = pi471 & ~pi532;
  assign n22816 = pi532 & pi674;
  assign po609 = n22815 | n22816;
  assign n22818 = pi472 & ~pi532;
  assign n22819 = pi532 & pi781;
  assign po610 = n22818 | n22819;
  assign n22821 = pi473 & ~pi532;
  assign n22822 = pi532 & pi745;
  assign po611 = n22821 | n22822;
  assign n22824 = pi474 & ~pi532;
  assign n22825 = pi532 & pi735;
  assign po612 = n22824 | n22825;
  assign n22827 = pi475 & ~pi532;
  assign n22828 = pi532 & pi677;
  assign po613 = n22827 | n22828;
  assign n22830 = pi476 & ~pi532;
  assign n22831 = pi532 & pi701;
  assign po614 = n22830 | n22831;
  assign n22833 = pi477 & ~pi532;
  assign n22834 = pi532 & pi676;
  assign po615 = n22833 | n22834;
  assign n22836 = pi478 & ~pi532;
  assign n22837 = pi532 & pi782;
  assign po616 = n22836 | n22837;
  assign n22839 = pi479 & ~pi532;
  assign n22840 = pi532 & pi702;
  assign po617 = n22839 | n22840;
  assign n22842 = pi480 & ~pi532;
  assign n22843 = pi532 & pi697;
  assign po618 = n22842 | n22843;
  assign n22845 = pi481 & ~pi532;
  assign n22846 = pi532 & pi681;
  assign po619 = n22845 | n22846;
  assign po620 = ~pi532 & n22529;
  assign n22849 = pi483 & ~pi532;
  assign n22850 = pi532 & pi693;
  assign po621 = n22849 | n22850;
  assign n22852 = pi484 & ~pi532;
  assign n22853 = pi532 & pi736;
  assign po622 = n22852 | n22853;
  assign n22855 = pi485 & ~pi532;
  assign n22856 = pi532 & pi749;
  assign po623 = n22855 | n22856;
  assign n22858 = pi486 & ~pi532;
  assign n22859 = pi532 & pi694;
  assign po624 = n22858 | n22859;
  assign n22861 = pi488 & ~pi532;
  assign n22862 = pi532 & pi786;
  assign po626 = n22861 | n22862;
  assign n22864 = pi489 & ~pi532;
  assign n22865 = pi532 & pi663;
  assign po627 = n22864 | n22865;
  assign n22867 = pi490 & ~pi532;
  assign n22868 = pi532 & pi705;
  assign po628 = n22867 | n22868;
  assign n22870 = pi491 & ~pi532;
  assign n22871 = pi532 & pi733;
  assign po629 = n22870 | n22871;
  assign n22873 = pi492 & ~pi532;
  assign n22874 = pi532 & pi762;
  assign po630 = n22873 | n22874;
  assign n22876 = pi493 & ~pi532;
  assign n22877 = pi532 & pi767;
  assign po631 = n22876 | n22877;
  assign n22879 = pi494 & ~pi532;
  assign n22880 = pi532 & pi665;
  assign po632 = n22879 | n22880;
  assign n22882 = pi495 & ~pi532;
  assign n22883 = pi532 & pi704;
  assign po633 = n22882 | n22883;
  assign n22885 = pi496 & ~pi532;
  assign n22886 = pi532 & pi773;
  assign po634 = n22885 | n22886;
  assign n22888 = pi497 & ~pi532;
  assign n22889 = pi532 & pi754;
  assign po635 = n22888 | n22889;
  assign n22891 = pi498 & ~pi532;
  assign n22892 = pi532 & pi734;
  assign po636 = n22891 | n22892;
  assign n22894 = pi499 & ~pi532;
  assign n22895 = pi532 & pi711;
  assign po637 = n22894 | n22895;
  assign n22897 = pi500 & ~pi532;
  assign n22898 = pi532 & pi761;
  assign po638 = n22897 | n22898;
  assign n22900 = pi501 & ~pi532;
  assign n22901 = pi532 & pi775;
  assign po639 = n22900 | n22901;
  assign n22903 = pi502 & ~pi532;
  assign n22904 = pi532 & pi686;
  assign po640 = n22903 | n22904;
  assign n22906 = pi503 & ~pi532;
  assign n22907 = pi532 & pi718;
  assign po641 = n22906 | n22907;
  assign n22909 = pi504 & ~pi532;
  assign n22910 = pi532 & pi756;
  assign po642 = n22909 | n22910;
  assign n22912 = pi505 & ~pi532;
  assign n22913 = pi532 & pi785;
  assign po643 = n22912 | n22913;
  assign n22915 = pi506 & ~pi532;
  assign n22916 = pi532 & pi776;
  assign po644 = n22915 | n22916;
  assign n22918 = pi507 & ~pi532;
  assign n22919 = pi532 & pi759;
  assign po645 = n22918 | n22919;
  assign n22921 = pi508 & ~pi532;
  assign n22922 = pi532 & pi692;
  assign po646 = n22921 | n22922;
  assign n22924 = pi509 & ~pi532;
  assign n22925 = pi532 & pi783;
  assign po647 = n22924 | n22925;
  assign n22927 = pi510 & ~pi532;
  assign n22928 = pi532 & pi780;
  assign po648 = n22927 | n22928;
  assign n22930 = pi511 & ~pi532;
  assign n22931 = pi532 & pi763;
  assign po649 = n22930 | n22931;
  assign n22933 = pi512 & ~pi532;
  assign n22934 = pi532 & pi737;
  assign po650 = n22933 | n22934;
  assign n22936 = pi513 & ~pi532;
  assign n22937 = pi532 & pi774;
  assign po651 = n22936 | n22937;
  assign n22939 = pi514 & ~pi532;
  assign n22940 = pi532 & pi755;
  assign po652 = n22939 | n22940;
  assign n22942 = pi515 & ~pi532;
  assign n22943 = pi532 & pi723;
  assign po653 = n22942 | n22943;
  assign n22945 = pi516 & ~pi532;
  assign n22946 = pi532 & pi709;
  assign po654 = n22945 | n22946;
  assign n22948 = pi517 & ~pi532;
  assign n22949 = pi532 & pi688;
  assign po655 = n22948 | n22949;
  assign n22951 = pi518 & ~pi532;
  assign n22952 = pi532 & pi770;
  assign po656 = n22951 | n22952;
  assign n22954 = pi519 & ~pi532;
  assign n22955 = pi532 & pi778;
  assign po657 = n22954 | n22955;
  assign n22957 = pi521 & ~pi532;
  assign n22958 = pi532 & pi682;
  assign po659 = n22957 | n22958;
  assign n22960 = pi522 & ~pi532;
  assign n22961 = pi532 & pi666;
  assign po660 = n22960 | n22961;
  assign n22963 = pi523 & ~pi532;
  assign n22964 = pi532 & pi683;
  assign po661 = n22963 | n22964;
  assign n22966 = pi524 & ~pi532;
  assign n22967 = pi532 & pi744;
  assign po662 = n22966 | n22967;
  assign n22969 = pi525 & ~pi532;
  assign n22970 = pi532 & pi699;
  assign po663 = n22969 | n22970;
  assign n22972 = pi526 & ~pi532;
  assign n22973 = pi532 & pi732;
  assign po664 = n22972 | n22973;
  assign n22975 = pi527 & ~pi532;
  assign n22976 = pi532 & pi750;
  assign po665 = n22975 | n22976;
  assign n22978 = pi528 & ~pi532;
  assign n22979 = pi532 & pi748;
  assign po666 = n22978 | n22979;
  assign po140 = 1'b1;
  assign po000 = pi397;
  assign po001 = pi211;
  assign po002 = pi305;
  assign po003 = pi339;
  assign po004 = pi345;
  assign po005 = pi212;
  assign po006 = pi262;
  assign po007 = pi213;
  assign po008 = pi306;
  assign po009 = pi383;
  assign po010 = pi322;
  assign po011 = pi206;
  assign po012 = pi336;
  assign po013 = pi158;
  assign po014 = pi241;
  assign po015 = pi332;
  assign po016 = pi331;
  assign po017 = pi261;
  assign po018 = pi381;
  assign po019 = pi296;
  assign po020 = pi243;
  assign po021 = pi374;
  assign po022 = pi259;
  assign po023 = pi329;
  assign po024 = pi295;
  assign po025 = pi288;
  assign po026 = pi341;
  assign po027 = pi365;
  assign po028 = pi338;
  assign po029 = pi340;
  assign po030 = pi235;
  assign po031 = pi294;
  assign po032 = pi323;
  assign po033 = pi214;
  assign po034 = pi309;
  assign po035 = pi337;
  assign po036 = pi264;
  assign po037 = pi308;
  assign po038 = pi263;
  assign po039 = pi307;
  assign po040 = pi310;
  assign po041 = pi317;
  assign po042 = pi304;
  assign po043 = pi245;
  assign po044 = pi196;
  assign po045 = pi177;
  assign po046 = pi237;
  assign po047 = pi204;
  assign po048 = pi244;
  assign po049 = pi201;
  assign po050 = pi382;
  assign po051 = pi314;
  assign po052 = pi236;
  assign po053 = pi367;
  assign po054 = pi282;
  assign po055 = pi326;
  assign po056 = pi325;
  assign po057 = pi277;
  assign po058 = pi298;
  assign po059 = pi343;
  assign po060 = pi315;
  assign po061 = pi300;
  assign po062 = pi188;
  assign po063 = pi249;
  assign po064 = pi360;
  assign po065 = pi216;
  assign po066 = pi347;
  assign po067 = pi335;
  assign po068 = pi266;
  assign po069 = pi311;
  assign po070 = pi265;
  assign po071 = pi312;
  assign po072 = pi313;
  assign po073 = pi318;
  assign po074 = pi291;
  assign po075 = pi247;
  assign po076 = pi289;
  assign po077 = pi199;
  assign po078 = pi240;
  assign po079 = pi252;
  assign po080 = pi246;
  assign po081 = pi202;
  assign po082 = pi378;
  assign po083 = pi293;
  assign po084 = pi287;
  assign po085 = pi368;
  assign po086 = pi286;
  assign po087 = pi377;
  assign po088 = pi380;
  assign po089 = pi279;
  assign po090 = pi299;
  assign po091 = pi327;
  assign po092 = pi316;
  assign po093 = pi333;
  assign po094 = pi186;
  assign po095 = pi250;
  assign po096 = pi369;
  assign po097 = pi361;
  assign po098 = pi359;
  assign po099 = pi366;
  assign po100 = pi379;
  assign po101 = pi248;
  assign po102 = pi194;
  assign po103 = pi324;
  assign po104 = pi330;
  assign po105 = pi239;
  assign po106 = pi238;
  assign po107 = pi292;
  assign po108 = pi355;
  assign po109 = pi195;
  assign po110 = pi197;
  assign po111 = pi251;
  assign po112 = pi200;
  assign po113 = pi203;
  assign po114 = pi362;
  assign po115 = pi297;
  assign po116 = pi242;
  assign po117 = pi334;
  assign po118 = pi198;
  assign po119 = pi364;
  assign po120 = pi328;
  assign po121 = pi260;
  assign po122 = pi253;
  assign po123 = pi344;
  assign po124 = pi290;
  assign po125 = pi254;
  assign po126 = pi176;
  assign po127 = pi205;
  assign po128 = pi363;
  assign po129 = pi530;
  assign po142 = pi529;
  assign po280 = pi532;
  assign po281 = pi626;
  assign po300 = pi621;
  assign po667 = pi532;
endmodule


