// Benchmark "usb_phy" written by ABC on Wed Apr 29 13:55:16 2015

module usb_phy ( 
    pi000, pi001, pi002, pi003, pi004, pi005, pi006, pi007, pi008, pi009,
    pi010, pi011, pi012, pi013, pi014, pi015, pi016, pi017, pi018, pi019,
    pi020, pi021, pi022, pi023, pi024, pi025, pi026, pi027, pi028, pi029,
    pi030, pi031, pi032, pi033, pi034, pi035, pi036, pi037, pi038, pi039,
    pi040, pi041, pi042, pi043, pi044, pi045, pi046, pi047, pi048, pi049,
    pi050, pi051, pi052, pi053, pi054, pi055, pi056, pi057, pi058, pi059,
    pi060, pi061, pi062, pi063, pi064, pi065, pi066, pi067, pi068, pi069,
    pi070, pi071, pi072, pi073, pi074, pi075, pi076, pi077, pi078, pi079,
    pi080, pi081, pi082, pi083, pi084, pi085, pi086, pi087, pi088, pi089,
    pi090, pi091, pi092, pi093, pi094, pi095, pi096, pi097, pi098, pi099,
    pi100, pi101, pi102, pi103, pi104, pi105, pi106, pi107, pi108, pi109,
    pi110, pi111, pi112,
    po000, po001, po002, po003, po004, po005, po006, po007, po008, po009,
    po010, po011, po012, po013, po014, po015, po016, po017, po018, po019,
    po020, po021, po022, po023, po024, po025, po026, po027, po028, po029,
    po030, po031, po032, po033, po034, po035, po036, po037, po038, po039,
    po040, po041, po042, po043, po044, po045, po046, po047, po048, po049,
    po050, po051, po052, po053, po054, po055, po056, po057, po058, po059,
    po060, po061, po062, po063, po064, po065, po066, po067, po068, po069,
    po070, po071, po072, po073, po074, po075, po076, po077, po078, po079,
    po080, po081, po082, po083, po084, po085, po086, po087, po088, po089,
    po090, po091, po092, po093, po094, po095, po096, po097, po098, po099,
    po100, po101, po102, po103, po104, po105, po106, po107, po108, po109,
    po110  );
  input  pi000, pi001, pi002, pi003, pi004, pi005, pi006, pi007, pi008,
    pi009, pi010, pi011, pi012, pi013, pi014, pi015, pi016, pi017, pi018,
    pi019, pi020, pi021, pi022, pi023, pi024, pi025, pi026, pi027, pi028,
    pi029, pi030, pi031, pi032, pi033, pi034, pi035, pi036, pi037, pi038,
    pi039, pi040, pi041, pi042, pi043, pi044, pi045, pi046, pi047, pi048,
    pi049, pi050, pi051, pi052, pi053, pi054, pi055, pi056, pi057, pi058,
    pi059, pi060, pi061, pi062, pi063, pi064, pi065, pi066, pi067, pi068,
    pi069, pi070, pi071, pi072, pi073, pi074, pi075, pi076, pi077, pi078,
    pi079, pi080, pi081, pi082, pi083, pi084, pi085, pi086, pi087, pi088,
    pi089, pi090, pi091, pi092, pi093, pi094, pi095, pi096, pi097, pi098,
    pi099, pi100, pi101, pi102, pi103, pi104, pi105, pi106, pi107, pi108,
    pi109, pi110, pi111, pi112;
  output po000, po001, po002, po003, po004, po005, po006, po007, po008, po009,
    po010, po011, po012, po013, po014, po015, po016, po017, po018, po019,
    po020, po021, po022, po023, po024, po025, po026, po027, po028, po029,
    po030, po031, po032, po033, po034, po035, po036, po037, po038, po039,
    po040, po041, po042, po043, po044, po045, po046, po047, po048, po049,
    po050, po051, po052, po053, po054, po055, po056, po057, po058, po059,
    po060, po061, po062, po063, po064, po065, po066, po067, po068, po069,
    po070, po071, po072, po073, po074, po075, po076, po077, po078, po079,
    po080, po081, po082, po083, po084, po085, po086, po087, po088, po089,
    po090, po091, po092, po093, po094, po095, po096, po097, po098, po099,
    po100, po101, po102, po103, po104, po105, po106, po107, po108, po109,
    po110;
  wire n226, n228, n230, n231, n232, n233, n234, n235, n236, n237, n238,
    n239, n240, n241, n242, n243, n244, n245, n246, n247, n248, n250, n251,
    n252, n253, n254, n255, n256, n257, n258, n259, n260, n261, n262, n263,
    n264, n265, n266, n268, n269, n270, n271, n272, n273, n275, n276, n277,
    n278, n279, n280, n281, n282, n283, n284, n285, n286, n287, n288, n290,
    n291, n292, n293, n294, n295, n296, n297, n299, n300, n301, n302, n303,
    n304, n305, n307, n308, n309, n311, n312, n313, n314, n315, n316, n318,
    n319, n320, n321, n322, n324, n325, n326, n328, n329, n330, n332, n333,
    n334, n336, n337, n338, n340, n341, n342, n344, n345, n346, n348, n349,
    n350, n352, n353, n355, n356, n357, n358, n359, n360, n361, n362, n363,
    n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
    n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n387, n388,
    n389, n390, n392, n393, n394, n395, n396, n397, n398, n400, n401, n402,
    n403, n404, n405, n407, n408, n409, n410, n411, n412, n413, n415, n417,
    n419, n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n431,
    n432, n433, n435, n436, n437, n438, n440, n441, n442, n443, n444, n445,
    n447, n448, n449, n450, n451, n452, n453, n454, n456, n457, n458, n459,
    n460, n461, n462, n463, n464, n465, n467, n468, n469, n470, n471, n472,
    n474, n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
    n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497,
    n498, n500, n501, n502, n503, n504, n505, n507, n508, n509, n510, n511,
    n512, n513, n514, n515, n517, n518, n520, n521, n522, n523, n525, n526,
    n527, n529, n530, n531, n532, n533, n534, n536, n537, n538, n539, n540,
    n542, n543, n544, n545, n546, n547, n548, n549, n551, n552, n553, n554,
    n555, n556, n557, n559, n560, n561, n562, n563, n564, n565, n566, n568,
    n569, n570, n572, n573, n574, n575, n577, n578, n579, n580, n584, n585,
    n587, n588, n589, n590, n591, n592, n594, n595, n596, n597, n598, n599,
    n600, n602, n603, n604, n605, n606, n607, n608, n610, n611, n612, n613,
    n615, n616, n617, n619, n620, n621, n622, n623, n624, n626, n627, n628,
    n629, n630, n632, n633, n634, n635, n641, n642, n644, n645, n646, n648,
    n649, n650, n652, n653, n654, n656, n657, n658, n660, n661, n662, n664,
    n665, n666, n667, n668, n669, n670, n671, n673, n674, n675, n677, n678,
    n679, n681, n682, n684;
  assign n226 = pi003 & pi006;
  assign po007 = ~pi008 | ~n226;
  assign n228 = ~pi002 & pi073;
  assign po043 = ~pi062 & ~pi063;
  assign n230 = n228 & ~po043;
  assign n231 = ~pi016 & n230;
  assign n232 = pi062 & ~pi063;
  assign n233 = pi095 & n232;
  assign n234 = pi063 & pi095;
  assign n235 = ~pi062 & n234;
  assign n236 = n233 & ~n235;
  assign n237 = pi001 & pi005;
  assign n238 = pi004 & n237;
  assign n239 = ~pi004 & n237;
  assign n240 = ~n238 & n239;
  assign n241 = n236 & n240;
  assign n242 = n232 & ~n239;
  assign n243 = n238 & n242;
  assign n244 = ~n241 & ~n243;
  assign n245 = n231 & ~n244;
  assign n246 = ~pi002 & ~n245;
  assign n247 = pi073 & ~n246;
  assign n248 = pi000 & ~pi073;
  assign po020 = n247 | n248;
  assign n250 = ~pi001 & pi005;
  assign n251 = pi004 & n250;
  assign n252 = n233 & n251;
  assign n253 = ~pi004 & n250;
  assign n254 = n233 & n253;
  assign n255 = ~n252 & ~n254;
  assign n256 = ~pi001 & ~pi005;
  assign n257 = pi004 & n256;
  assign n258 = n233 & n257;
  assign n259 = ~pi001 & ~n233;
  assign n260 = ~pi004 & ~n259;
  assign n261 = n256 & n260;
  assign n262 = ~n258 & ~n261;
  assign n263 = n231 & n262;
  assign n264 = n255 & n263;
  assign n265 = ~pi001 & ~n231;
  assign n266 = ~n264 & ~n265;
  assign po021 = pi099 & n266;
  assign n268 = pi095 & pi099;
  assign n269 = n231 & n268;
  assign n270 = ~n244 & n269;
  assign n271 = pi022 & po043;
  assign n272 = pi002 & ~n271;
  assign n273 = pi099 & n272;
  assign po022 = n270 | n273;
  assign n275 = pi001 & ~pi005;
  assign n276 = pi004 & n275;
  assign n277 = ~n235 & n276;
  assign n278 = ~n233 & n257;
  assign n279 = ~n277 & ~n278;
  assign n280 = ~pi004 & n275;
  assign n281 = ~n235 & n280;
  assign n282 = n279 & ~n281;
  assign n283 = ~n235 & n239;
  assign n284 = ~n253 & ~n283;
  assign n285 = ~n251 & n284;
  assign n286 = ~n233 & ~n285;
  assign n287 = n282 & ~n286;
  assign n288 = ~pi002 & n231;
  assign po023 = ~n287 & n288;
  assign n290 = pi004 & ~n231;
  assign n291 = n235 & n280;
  assign n292 = n235 & n239;
  assign n293 = ~n258 & ~n292;
  assign n294 = ~n252 & n293;
  assign n295 = ~n291 & n294;
  assign n296 = n231 & ~n295;
  assign n297 = ~n290 & ~n296;
  assign po024 = pi099 & ~n297;
  assign n299 = n235 & n276;
  assign n300 = ~n252 & ~n299;
  assign n301 = ~n254 & ~n292;
  assign n302 = n300 & n301;
  assign n303 = n231 & ~n302;
  assign n304 = pi005 & ~n231;
  assign n305 = ~n303 & ~n304;
  assign po025 = pi099 & ~n305;
  assign n307 = ~pi031 & ~pi036;
  assign n308 = pi023 & ~n307;
  assign n309 = pi002 & po043;
  assign po026 = n308 & n309;
  assign n311 = pi007 & pi037;
  assign n312 = ~pi019 & ~pi027;
  assign n313 = ~pi017 & n312;
  assign n314 = pi104 & n313;
  assign n315 = ~pi037 & pi112;
  assign n316 = ~n314 & ~n315;
  assign po027 = n311 | ~n316;
  assign n318 = pi028 & pi029;
  assign n319 = ~pi034 & n318;
  assign n320 = pi002 & pi073;
  assign n321 = n319 & n320;
  assign n322 = ~po043 & n321;
  assign po028 = pi056 & n322;
  assign n324 = ~pi037 & pi105;
  assign n325 = pi009 & pi037;
  assign n326 = ~n324 & ~n325;
  assign po029 = ~n314 & ~n326;
  assign n328 = ~pi037 & pi106;
  assign n329 = pi010 & pi037;
  assign n330 = ~n328 & ~n329;
  assign po030 = ~n314 & ~n330;
  assign n332 = ~pi037 & pi107;
  assign n333 = pi011 & pi037;
  assign n334 = ~n332 & ~n333;
  assign po031 = ~n314 & ~n334;
  assign n336 = ~pi037 & pi108;
  assign n337 = pi012 & pi037;
  assign n338 = ~n336 & ~n337;
  assign po032 = ~n314 & ~n338;
  assign n340 = ~pi037 & pi109;
  assign n341 = pi013 & pi037;
  assign n342 = ~n340 & ~n341;
  assign po033 = ~n314 & ~n342;
  assign n344 = ~pi037 & pi110;
  assign n345 = pi014 & pi037;
  assign n346 = ~n344 & ~n345;
  assign po034 = ~n314 & ~n346;
  assign n348 = ~pi037 & pi111;
  assign n349 = pi015 & pi037;
  assign n350 = ~n348 & ~n349;
  assign po035 = ~n314 & ~n350;
  assign n352 = pi073 & po043;
  assign n353 = pi016 & ~pi073;
  assign po036 = n352 | n353;
  assign n355 = pi064 & ~pi091;
  assign n356 = ~pi019 & n355;
  assign n357 = ~pi017 & ~pi077;
  assign n358 = pi027 & n357;
  assign n359 = n356 & n358;
  assign n360 = pi019 & ~pi027;
  assign n361 = ~pi017 & n360;
  assign n362 = ~n313 & ~n361;
  assign n363 = pi017 & ~n362;
  assign n364 = ~pi060 & pi073;
  assign n365 = n361 & n364;
  assign n366 = ~n314 & ~n365;
  assign n367 = ~pi017 & ~pi019;
  assign n368 = pi027 & n367;
  assign n369 = pi017 & n368;
  assign n370 = n366 & ~n369;
  assign n371 = ~n363 & n370;
  assign n372 = ~n359 & n371;
  assign n373 = ~pi019 & pi027;
  assign n374 = pi017 & n373;
  assign n375 = pi017 & ~pi060;
  assign n376 = n374 & n375;
  assign n377 = ~pi027 & ~pi073;
  assign n378 = pi019 & n377;
  assign n379 = pi017 & n378;
  assign n380 = pi017 & n312;
  assign n381 = ~n355 & n380;
  assign n382 = ~n379 & ~n381;
  assign n383 = pi017 & ~n382;
  assign n384 = ~n376 & ~n383;
  assign n385 = n372 & n384;
  assign po037 = pi099 & ~n385;
  assign n387 = pi074 & pi081;
  assign n388 = ~pi074 & ~pi081;
  assign n389 = ~n387 & ~n388;
  assign n390 = pi095 & n389;
  assign po094 = pi018 & ~pi021;
  assign n392 = n390 & po094;
  assign n393 = ~pi018 & ~pi021;
  assign n394 = ~n390 & n393;
  assign n395 = ~n392 & ~n394;
  assign n396 = pi021 & ~n390;
  assign n397 = ~pi018 & n396;
  assign n398 = n395 & ~n397;
  assign po038 = ~pi099 | ~n398;
  assign n400 = ~n361 & ~n379;
  assign n401 = pi019 & ~n400;
  assign n402 = ~n365 & ~n401;
  assign n403 = ~pi019 & ~pi060;
  assign n404 = n374 & ~n403;
  assign n405 = n402 & ~n404;
  assign po039 = pi099 & ~n405;
  assign n407 = pi073 & ~n319;
  assign n408 = pi020 & ~n407;
  assign n409 = pi099 & n408;
  assign n410 = pi035 & pi036;
  assign n411 = pi031 & n407;
  assign n412 = pi099 & n411;
  assign n413 = n410 & n412;
  assign po040 = n409 | n413;
  assign n415 = ~po094 & ~n397;
  assign po041 = pi099 & ~n415;
  assign n417 = pi022 & ~pi073;
  assign po042 = pi044 | n417;
  assign n419 = ~pi070 & pi073;
  assign n420 = pi054 & pi058;
  assign n421 = pi026 & n420;
  assign n422 = pi024 & ~n421;
  assign n423 = ~pi024 & n421;
  assign n424 = ~n422 & ~n423;
  assign n425 = n419 & ~n424;
  assign n426 = pi024 & ~n419;
  assign n427 = ~n425 & ~n426;
  assign n428 = ~pi082 & ~pi084;
  assign n429 = pi099 & n428;
  assign po044 = ~n427 & n429;
  assign n431 = pi025 & ~n419;
  assign n432 = pi024 & pi026;
  assign n433 = n420 & n432;
  assign po084 = pi025 & n433;
  assign n435 = ~pi025 & ~n433;
  assign n436 = ~po084 & ~n435;
  assign n437 = n419 & n436;
  assign n438 = ~n431 & ~n437;
  assign po045 = n429 & ~n438;
  assign n440 = ~pi026 & n420;
  assign n441 = pi026 & ~n420;
  assign n442 = ~n440 & ~n441;
  assign n443 = n419 & ~n442;
  assign n444 = pi026 & ~n419;
  assign n445 = ~n443 & ~n444;
  assign po046 = n429 & ~n445;
  assign n447 = pi027 & n368;
  assign n448 = pi027 & ~pi060;
  assign n449 = n374 & n448;
  assign n450 = ~pi027 & ~n355;
  assign n451 = n380 & ~n450;
  assign n452 = ~n449 & ~n451;
  assign n453 = ~n447 & n452;
  assign n454 = ~n359 & n453;
  assign po047 = pi099 & ~n454;
  assign n456 = pi000 & pi099;
  assign n457 = pi029 & pi034;
  assign n458 = pi028 & ~n457;
  assign n459 = ~pi028 & n457;
  assign n460 = ~n458 & ~n459;
  assign n461 = pi056 & ~n319;
  assign n462 = pi073 & n461;
  assign n463 = ~n460 & n462;
  assign n464 = pi028 & ~pi073;
  assign n465 = ~n463 & ~n464;
  assign po048 = n456 & ~n465;
  assign n467 = pi029 & ~pi073;
  assign n468 = pi029 & ~pi034;
  assign n469 = ~pi029 & pi034;
  assign n470 = ~n468 & ~n469;
  assign n471 = n462 & ~n470;
  assign n472 = ~n467 & ~n471;
  assign po049 = n456 & ~n472;
  assign n474 = pi041 & pi042;
  assign n475 = pi096 & n474;
  assign n476 = pi032 & n475;
  assign n477 = ~pi032 & n474;
  assign n478 = ~pi088 & n477;
  assign n479 = ~n476 & ~n478;
  assign n480 = pi041 & ~pi042;
  assign n481 = ~pi085 & n480;
  assign n482 = ~pi041 & ~pi042;
  assign n483 = pi092 & n482;
  assign n484 = ~n481 & ~n483;
  assign n485 = ~pi032 & ~n484;
  assign n486 = n479 & ~n485;
  assign n487 = pi097 & n482;
  assign n488 = pi032 & n487;
  assign n489 = ~pi041 & pi042;
  assign n490 = ~pi032 & pi094;
  assign n491 = n489 & n490;
  assign n492 = ~n488 & ~n491;
  assign n493 = ~pi090 & n489;
  assign n494 = ~pi086 & n480;
  assign n495 = ~n493 & ~n494;
  assign n496 = pi032 & ~n495;
  assign n497 = n492 & ~n496;
  assign n498 = n486 & n497;
  assign po050 = pi065 & ~n498;
  assign n500 = pi031 & ~n407;
  assign n501 = pi031 & ~n410;
  assign n502 = ~pi031 & n410;
  assign n503 = ~n501 & ~n502;
  assign n504 = n407 & ~n503;
  assign n505 = ~n500 & ~n504;
  assign po051 = n456 & ~n505;
  assign n507 = pi038 & pi039;
  assign n508 = ~pi043 & n507;
  assign n509 = pi073 & ~n508;
  assign n510 = pi032 & ~n474;
  assign n511 = ~n477 & ~n510;
  assign n512 = n509 & ~n511;
  assign n513 = pi032 & ~n509;
  assign n514 = ~n512 & ~n513;
  assign n515 = pi065 & pi099;
  assign po052 = ~n514 & n515;
  assign n517 = pi033 & ~pi068;
  assign n518 = ~n359 & ~n517;
  assign po053 = pi099 & ~n518;
  assign n520 = pi034 & ~pi073;
  assign n521 = ~pi034 & n461;
  assign n522 = pi073 & n521;
  assign n523 = ~n520 & ~n522;
  assign po054 = n456 & ~n523;
  assign n525 = pi035 & ~n407;
  assign n526 = ~pi035 & n407;
  assign n527 = ~n525 & ~n526;
  assign po055 = n456 & ~n527;
  assign n529 = pi036 & ~n407;
  assign n530 = ~pi035 & pi036;
  assign n531 = pi035 & ~pi036;
  assign n532 = ~n530 & ~n531;
  assign n533 = n407 & ~n532;
  assign n534 = ~n529 & ~n533;
  assign po056 = n456 & ~n534;
  assign n536 = pi077 & n355;
  assign n537 = n368 & n536;
  assign n538 = ~n380 & n537;
  assign n539 = n355 & n380;
  assign n540 = ~n368 & n539;
  assign po057 = n538 | n540;
  assign n542 = pi038 & ~pi073;
  assign n543 = pi038 & ~pi043;
  assign n544 = ~pi038 & pi043;
  assign n545 = ~n543 & ~n544;
  assign n546 = pi030 & ~n508;
  assign n547 = pi073 & n546;
  assign n548 = ~n545 & n547;
  assign n549 = ~n542 & ~n548;
  assign po058 = n515 & ~n549;
  assign n551 = pi039 & ~pi073;
  assign n552 = pi038 & pi043;
  assign n553 = pi039 & ~n552;
  assign n554 = ~pi039 & n552;
  assign n555 = ~n553 & ~n554;
  assign n556 = n547 & ~n555;
  assign n557 = ~n551 & ~n556;
  assign po059 = n515 & ~n557;
  assign n559 = pi099 & pi104;
  assign n560 = ~pi017 & pi027;
  assign n561 = n559 & ~n560;
  assign n562 = n539 & n561;
  assign n563 = ~pi017 & ~n380;
  assign n564 = n536 & n563;
  assign n565 = pi027 & n564;
  assign n566 = n559 & n565;
  assign po060 = n562 | n566;
  assign n568 = pi041 & ~n509;
  assign n569 = ~pi041 & n509;
  assign n570 = ~n568 & ~n569;
  assign po061 = n515 & ~n570;
  assign n572 = pi042 & ~n509;
  assign n573 = ~n480 & ~n489;
  assign n574 = n509 & ~n573;
  assign n575 = ~n572 & ~n574;
  assign po062 = n515 & ~n575;
  assign n577 = pi043 & ~pi073;
  assign n578 = ~pi043 & n546;
  assign n579 = pi073 & n578;
  assign n580 = ~n577 & ~n579;
  assign po063 = n515 & ~n580;
  assign po064 = pi020 & n407;
  assign po065 = ~pi000 | ~n407;
  assign n584 = pi053 & ~pi060;
  assign n585 = ~n314 & ~n584;
  assign po067 = pi099 & ~n585;
  assign n587 = pi054 & ~n419;
  assign n588 = pi054 & ~pi058;
  assign n589 = ~pi054 & pi058;
  assign n590 = ~n588 & ~n589;
  assign n591 = n419 & ~n590;
  assign n592 = ~n587 & ~n591;
  assign po068 = n429 & ~n592;
  assign n594 = pi073 & ~pi100;
  assign n595 = pi073 & pi100;
  assign n596 = ~pi060 & n595;
  assign n597 = ~n594 & ~n596;
  assign n598 = pi071 & ~n597;
  assign n599 = pi055 & ~pi073;
  assign n600 = ~n598 & ~n599;
  assign po069 = ~pi099 | ~n600;
  assign n602 = pi074 & pi075;
  assign n603 = ~pi074 & ~pi075;
  assign n604 = ~n602 & ~n603;
  assign n605 = n320 & ~n604;
  assign n606 = pi056 & ~n320;
  assign n607 = ~n605 & ~n606;
  assign n608 = pi002 & n607;
  assign po070 = pi099 & ~n608;
  assign n610 = ~pi073 & pi099;
  assign n611 = pi057 & n610;
  assign n612 = pi030 & n509;
  assign n613 = n515 & n612;
  assign po071 = n611 | n613;
  assign n615 = ~pi058 & n419;
  assign n616 = pi058 & ~n419;
  assign n617 = ~n615 & ~n616;
  assign po072 = n429 & ~n617;
  assign n619 = pi059 & ~pi073;
  assign n620 = pi060 & ~n594;
  assign n621 = ~pi071 & n595;
  assign n622 = ~pi060 & ~n621;
  assign n623 = ~n620 & ~n622;
  assign n624 = ~n619 & ~n623;
  assign po073 = pi099 & ~n624;
  assign n626 = pi060 & n610;
  assign n627 = pi060 & ~pi072;
  assign n628 = ~pi068 & ~n627;
  assign n629 = pi073 & ~n628;
  assign n630 = pi099 & n629;
  assign po074 = n626 | n630;
  assign n632 = ~pi066 & ~pi069;
  assign n633 = pi073 & n632;
  assign n634 = pi061 & ~pi073;
  assign n635 = ~n633 & ~n634;
  assign po075 = ~pi099 | ~n635;
  assign po092 = pi082 & pi089;
  assign po076 = ~pi078 | po092;
  assign po093 = pi084 & pi093;
  assign po077 = ~pi079 | po093;
  assign n641 = pi042 & ~n508;
  assign n642 = pi032 & n641;
  assign po078 = pi041 & n642;
  assign n644 = pi053 & pi073;
  assign n645 = pi065 & ~pi073;
  assign n646 = ~n644 & ~n645;
  assign po079 = pi099 & ~n646;
  assign n648 = pi065 & pi073;
  assign n649 = pi066 & ~pi073;
  assign n650 = ~n648 & ~n649;
  assign po080 = pi099 & ~n650;
  assign n652 = pi033 & pi073;
  assign n653 = pi067 & ~pi073;
  assign n654 = ~n652 & ~n653;
  assign po081 = pi099 & ~n654;
  assign n656 = pi067 & pi073;
  assign n657 = pi068 & ~pi073;
  assign n658 = ~n656 & ~n657;
  assign po082 = pi099 & ~n658;
  assign n660 = pi069 & ~pi073;
  assign n661 = pi066 & pi073;
  assign n662 = ~n660 & ~n661;
  assign po083 = pi099 & ~n662;
  assign n664 = pi057 & pi071;
  assign n665 = ~pi057 & ~pi071;
  assign n666 = ~n664 & ~n665;
  assign n667 = pi073 & ~n666;
  assign n668 = pi071 & ~pi073;
  assign n669 = ~n667 & ~n668;
  assign n670 = pi065 & n669;
  assign n671 = pi099 & n670;
  assign po085 = ~pi066 | ~n671;
  assign n673 = pi072 & ~pi073;
  assign n674 = pi060 & pi073;
  assign n675 = ~n673 & ~n674;
  assign po086 = pi099 & ~n675;
  assign n677 = pi074 & pi087;
  assign n678 = ~pi074 & ~pi087;
  assign n679 = ~pi083 & ~n678;
  assign po088 = n677 | n679;
  assign n681 = pi073 & pi074;
  assign n682 = ~pi073 & pi075;
  assign po089 = n681 | n682;
  assign n684 = pi053 & ~pi077;
  assign po091 = n559 & ~n684;
  assign po018 = 1'b1;
  assign po000 = pi070;
  assign po001 = pi055;
  assign po002 = pi059;
  assign po003 = pi061;
  assign po004 = pi040;
  assign po005 = pi044;
  assign po006 = pi002;
  assign po008 = pi047;
  assign po009 = pi048;
  assign po010 = pi049;
  assign po011 = pi050;
  assign po012 = pi046;
  assign po013 = pi051;
  assign po014 = pi045;
  assign po015 = pi052;
  assign po016 = pi084;
  assign po017 = pi082;
  assign po019 = pi098;
  assign po066 = pi056;
  assign po087 = pi076;
  assign po090 = pi080;
  assign po095 = pi074;
  assign po096 = pi089;
  assign po097 = pi087;
  assign po098 = pi093;
  assign po099 = pi010;
  assign po100 = pi014;
  assign po101 = pi101;
  assign po102 = pi012;
  assign po103 = pi103;
  assign po104 = pi015;
  assign po105 = pi064;
  assign po106 = pi009;
  assign po107 = pi102;
  assign po108 = pi011;
  assign po109 = pi007;
  assign po110 = pi013;
endmodule


