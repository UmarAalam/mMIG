//Written by the Majority Logic Package Wed Apr 29 21:27:03 2015
module top (
            pi000, pi001, pi002, pi003, pi004, pi005, pi006, pi007, pi008, pi009, pi010, pi011, pi012, pi013, pi014, pi015, pi016, pi017, pi018, pi019, pi020, pi021, pi022, pi023, pi024, pi025, pi026, pi027, pi028, pi029, pi030, pi031, pi032, pi033, pi034, pi035, pi036, pi037, pi038, pi039, pi040, pi041, pi042, pi043, pi044, pi045, pi046, pi047, pi048, pi049, pi050, pi051, pi052, pi053, pi054, pi055, pi056, pi057, pi058, pi059, pi060, pi061, pi062, pi063, pi064, pi065, pi066, pi067, pi068, pi069, pi070, pi071, pi072, pi073, pi074, pi075, pi076, pi077, pi078, pi079, pi080, pi081, pi082, pi083, pi084, pi085, pi086, pi087, pi088, pi089, pi090, pi091, pi092, pi093, pi094, pi095, pi096, pi097, pi098, pi099, pi100, pi101, pi102, pi103, pi104, pi105, pi106, pi107, pi108, pi109, pi110, pi111, pi112, pi113, pi114, pi115, pi116, pi117, pi118, pi119, pi120, pi121, pi122, pi123, pi124, pi125, pi126, pi127, pi128, pi129, pi130, pi131, pi132, pi133, pi134, pi135, pi136, pi137, pi138, pi139, pi140, pi141, pi142, pi143, pi144, pi145, pi146, pi147, pi148, pi149, pi150, pi151, pi152, pi153, pi154, pi155, pi156, pi157, pi158, pi159, pi160, pi161, pi162, pi163, pi164, pi165, pi166, pi167, pi168, pi169, pi170, pi171, pi172, pi173, pi174, pi175, pi176, pi177, pi178, pi179, pi180, pi181, pi182, pi183, pi184, pi185, pi186, pi187, pi188, pi189, pi190, pi191, pi192, pi193, pi194, pi195, pi196, pi197, pi198, pi199, pi200, pi201, pi202, pi203, pi204, pi205, pi206, pi207, pi208, pi209, pi210, pi211, pi212, pi213, pi214, pi215, pi216, pi217, pi218, pi219, pi220, pi221, pi222, pi223, pi224, pi225, pi226, pi227, pi228, pi229, pi230, pi231, pi232, pi233, pi234, pi235, pi236, pi237, pi238, pi239, pi240, pi241, pi242, pi243, pi244, pi245, pi246, pi247, pi248, pi249, pi250, pi251, pi252, pi253, pi254, pi255, pi256, pi257, pi258, pi259, pi260, pi261, pi262, pi263, pi264, pi265, pi266, pi267, pi268, pi269, pi270, pi271, pi272, pi273, pi274, pi275, pi276, pi277, pi278, pi279, pi280, pi281, pi282, pi283, pi284, pi285, pi286, pi287, pi288, pi289, pi290, pi291, pi292, pi293, pi294, pi295, pi296, pi297, pi298, pi299, pi300, pi301, pi302, pi303, pi304, pi305, pi306, pi307, pi308, pi309, pi310, pi311, pi312, pi313, pi314, pi315, pi316, pi317, pi318, pi319, pi320, pi321, pi322, pi323, pi324, pi325, pi326, pi327, pi328, pi329, pi330, pi331, pi332, pi333, pi334, pi335, pi336, pi337, pi338, pi339, pi340, pi341, pi342, pi343, pi344, pi345, pi346, pi347, pi348, pi349, pi350, pi351, pi352, pi353, pi354, pi355, pi356, pi357, pi358, pi359, pi360, pi361, pi362, pi363, pi364, pi365, pi366, pi367, 
            po00, po01, po02, po03, po04, po05, po06, po07, po08, po09, po10, po11, po12, po13, po14, po15, po16, po17, po18, po19, po20, po21, po22, po23, po24, po25, po26, po27, po28, po29, po30, po31, po32, po33, po34, po35, po36, po37, po38, po39, po40, po41, po42, po43, po44, po45, po46, po47, po48, po49, po50, po51, po52, po53, po54, po55, po56, po57, po58, po59, po60, po61, po62, po63, po64, po65, po66, po67, po68, po69, po70, po71);
input pi000, pi001, pi002, pi003, pi004, pi005, pi006, pi007, pi008, pi009, pi010, pi011, pi012, pi013, pi014, pi015, pi016, pi017, pi018, pi019, pi020, pi021, pi022, pi023, pi024, pi025, pi026, pi027, pi028, pi029, pi030, pi031, pi032, pi033, pi034, pi035, pi036, pi037, pi038, pi039, pi040, pi041, pi042, pi043, pi044, pi045, pi046, pi047, pi048, pi049, pi050, pi051, pi052, pi053, pi054, pi055, pi056, pi057, pi058, pi059, pi060, pi061, pi062, pi063, pi064, pi065, pi066, pi067, pi068, pi069, pi070, pi071, pi072, pi073, pi074, pi075, pi076, pi077, pi078, pi079, pi080, pi081, pi082, pi083, pi084, pi085, pi086, pi087, pi088, pi089, pi090, pi091, pi092, pi093, pi094, pi095, pi096, pi097, pi098, pi099, pi100, pi101, pi102, pi103, pi104, pi105, pi106, pi107, pi108, pi109, pi110, pi111, pi112, pi113, pi114, pi115, pi116, pi117, pi118, pi119, pi120, pi121, pi122, pi123, pi124, pi125, pi126, pi127, pi128, pi129, pi130, pi131, pi132, pi133, pi134, pi135, pi136, pi137, pi138, pi139, pi140, pi141, pi142, pi143, pi144, pi145, pi146, pi147, pi148, pi149, pi150, pi151, pi152, pi153, pi154, pi155, pi156, pi157, pi158, pi159, pi160, pi161, pi162, pi163, pi164, pi165, pi166, pi167, pi168, pi169, pi170, pi171, pi172, pi173, pi174, pi175, pi176, pi177, pi178, pi179, pi180, pi181, pi182, pi183, pi184, pi185, pi186, pi187, pi188, pi189, pi190, pi191, pi192, pi193, pi194, pi195, pi196, pi197, pi198, pi199, pi200, pi201, pi202, pi203, pi204, pi205, pi206, pi207, pi208, pi209, pi210, pi211, pi212, pi213, pi214, pi215, pi216, pi217, pi218, pi219, pi220, pi221, pi222, pi223, pi224, pi225, pi226, pi227, pi228, pi229, pi230, pi231, pi232, pi233, pi234, pi235, pi236, pi237, pi238, pi239, pi240, pi241, pi242, pi243, pi244, pi245, pi246, pi247, pi248, pi249, pi250, pi251, pi252, pi253, pi254, pi255, pi256, pi257, pi258, pi259, pi260, pi261, pi262, pi263, pi264, pi265, pi266, pi267, pi268, pi269, pi270, pi271, pi272, pi273, pi274, pi275, pi276, pi277, pi278, pi279, pi280, pi281, pi282, pi283, pi284, pi285, pi286, pi287, pi288, pi289, pi290, pi291, pi292, pi293, pi294, pi295, pi296, pi297, pi298, pi299, pi300, pi301, pi302, pi303, pi304, pi305, pi306, pi307, pi308, pi309, pi310, pi311, pi312, pi313, pi314, pi315, pi316, pi317, pi318, pi319, pi320, pi321, pi322, pi323, pi324, pi325, pi326, pi327, pi328, pi329, pi330, pi331, pi332, pi333, pi334, pi335, pi336, pi337, pi338, pi339, pi340, pi341, pi342, pi343, pi344, pi345, pi346, pi347, pi348, pi349, pi350, pi351, pi352, pi353, pi354, pi355, pi356, pi357, pi358, pi359, pi360, pi361, pi362, pi363, pi364, pi365, pi366, pi367;
output po00, po01, po02, po03, po04, po05, po06, po07, po08, po09, po10, po11, po12, po13, po14, po15, po16, po17, po18, po19, po20, po21, po22, po23, po24, po25, po26, po27, po28, po29, po30, po31, po32, po33, po34, po35, po36, po37, po38, po39, po40, po41, po42, po43, po44, po45, po46, po47, po48, po49, po50, po51, po52, po53, po54, po55, po56, po57, po58, po59, po60, po61, po62, po63, po64, po65, po66, po67, po68, po69, po70, po71;
wire one,v0, v1, v2, v3, v4, v5, v6, v7, v8, v9, v10, v11, v12, v13, v14, v15, v16, v17, v18, v19, v20, v21, v22, v23, v24, v25, v26, v27, v28, v29, v30, v31, v32, v33, v34, v35, v36, v37, v38, v39, v40, v41, v42, v43, v44, v45, v46, v47, v48, v49, v50, v51, v52, v53, v54, v55, v56, v57, v58, v59, v60, v61, v62, v63, v64, v65, v66, v67, v68, v69, v70, v71, v72, v73, v74, v75, v76, v77, v78, v79, v80, v81, v82, v83, v84, v85, v86, v87, v88, v89, v90, v91, v92, v93, v94, v95, v96, v97, v98, v99, v100, v101, v102, v103, v104, v105, v106, v107, v108, v109, v110, v111, v112, v113, v114, v115, v116, v117, v118, v119, v120, v121, v122, v123, v124, v125, v126, v127, v128, v129, v130, v131, v132, v133, v134, v135, v136, v137, v138, v139, v140, v141, v142, v143, v144, v145, v146, v147, v148, v149, v150, v151, v152, v153, v154, v155, v156, v157, v158, v159, v160, v161, v162, v163, v164, v165, v166, v167, v168, v169, v170, v171, v172, v173, v174, v175, v176, v177, v178, v179, v180, v181, v182, v183, v184, v185, v186, v187, v188, v189, v190, v191, v192, v193, v194, v195, v196, v197, v198, v199, v200, v201, v202, v203, v204, v205, v206, v207, v208, v209, v210, v211, v212, v213, v214, v215, v216, v217, v218, v219, v220, v221, v222, v223, v224, v225, v226, v227, v228, v229, v230, v231, v232, v233, v234, v235, v236, v237, v238, v239, v240, v241, v242, v243, v244, v245, v246, v247, v248, v249, v250, v251, v252, v253, v254, v255, v256, v257, v258, v259, v260, v261, v262, v263, v264, v265, v266, v267, v268, v269, v270, v271, v272, v273, v274, v275, v276, v277, v278, v279, v280, v281, v282, v283, v284, v285, v286, v287, v288, v289, v290, v291, v292, v293, v294, v295, v296, v297, v298, v299, v300, v301, v302, v303, v304, v305, v306, v307, v308, v309, v310, v311, v312, v313, v314, v315, v316, v317, v318, v319, v320, v321, v322, v323, v324, v325, v326, v327, v328, v329, v330, v331, v332, v333, v334, v335, v336, v337, v338, v339, v340, v341, v342, v343, v344, v345, v346, v347, v348, v349, v350, v351, v352, v353, v354, v355, v356, v357, v358, v359, v360, v361, v362, v363, v364, v365, v366, v367, v368, v369, v370, v371, v372, v373, v374, v375, v376, v377, v378, v379, v380, v381, v382, v383, v384, v385, v386, v387, v388, v389, v390, v391, v392, v393, v394, v395, v396, v397, v398, v399, v400, v401, v402, v403, v404, v405, v406, v407, v408, v409, v410, v411, v412, v413, v414, v415, v416, v417, v418, v419, v420, v421, v422, v423, v424, v425, v426, v427, v428, v429, v430, v431, v432, v433, v434, v435, v436, v437, v438, v439, v440, v441, v442, v443, v444, v445, v446, v447, v448, v449, v450, v451, v452, v453, v454, v455, v456, v457, v458, v459, v460, v461, v462, v463, v464, v465, v466, v467, v468, v469, v470, v471, v472, v473, v474, v475, v476, v477, v478, v479, v480, v481, v482, v483, v484, v485, v486, v487, v488, v489, v490, v491, v492, v493, v494, v495, v496, v497, v498, v499, v500, v501, v502, v503, v504, v505, v506, v507, v508, v509, v510, v511, v512, v513, v514, v515, v516, v517, v518, v519, v520, v521, v522, v523, v524, v525, v526, v527, v528, v529, v530, v531, v532, v533, v534, v535, v536, v537, v538, v539, v540, v541, v542, v543, v544, v545, v546, v547, v548, v549, v550, v551, v552, v553, v554, v555, v556, v557, v558, v559, v560, v561, v562, v563, v564, v565, v566, v567, v568, v569, v570, v571, v572, v573, v574, v575, v576, v577, v578, v579, v580, v581, v582, v583, v584, v585, v586, v587, v588, v589, v590, v591, v592, v593, v594, v595, v596, v597, v598, v599, v600, v601, v602, v603, v604, v605, v606, v607, v608, v609, v610, v611, v612, v613, v614, v615, v616, v617, v618, v619, v620, v621, v622, v623, v624, v625, v626, v627, v628, v629, v630, v631, v632, v633, v634, v635, v636, v637, v638, v639, v640, v641, v642, v643, v644, v645, v646, v647, v648, v649, v650, v651, v652, v653, v654, v655, v656, v657, v658, v659, v660, v661, v662, v663, v664, v665, v666, v667, v668, v669, v670, v671, v672, v673, v674, v675, v676, v677, v678, v679, v680, v681, v682, v683, v684, v685, v686, v687, v688, v689, v690, v691, v692, v693, v694, v695, v696, v697, v698, v699, v700, v701, v702, v703, v704, v705, v706, v707, v708, v709, v710, v711, v712, v713, v714, v715, v716, v717, v718, v719, v720, v721, v722, v723, v724, v725, v726, v727, v728, v729, v730, v731, v732, v733, v734, v735, v736, v737, v738, v739, v740, v741, v742, v743, v744, v745, v746, v747, v748, v749, v750, v751, v752, v753, v754, v755, v756, v757, v758, v759, v760, v761, v762, v763, v764, v765, v766, v767, v768, v769, v770, v771, v772, v773, v774, v775, v776, v777, v778, v779, v780, v781, v782, v783, v784, v785, v786, v787, v788, v789, v790, v791, v792, v793, v794, v795, v796, v797, v798, v799, v800, v801, v802, v803, v804, v805, v806, v807, v808, v809, v810, v811, v812, v813, v814, v815, v816, v817, v818, v819, v820, v821, v822, v823, v824, v825, v826, v827, v828, v829, v830, v831, v832, v833, v834, v835, v836, v837, v838, v839, v840, v841, v842, v843, v844, v845, v846, v847, v848, v849, v850, v851, v852, v853, v854, v855, v856, v857, v858, v859, v860, v861, v862, v863, v864, v865, v866, v867, v868, v869, v870, v871, v872, v873, v874, v875, v876, v877, v878, v879, v880, v881, v882, v883, v884, v885, v886, v887, v888, v889, v890, v891, v892, v893, v894, v895, v896, v897, v898, v899, v900, v901, v902, v903, v904, v905, v906, v907, v908, v909, v910, v911, v912, v913, v914, v915, v916, v917, v918, v919, v920, v921, v922, v923, v924, v925, v926, v927, v928, v929, v930, v931, v932, v933, v934, v935, v936, v937, v938, v939, v940, v941, v942, v943, v944, v945, v946, v947, v948, v949, v950, v951, v952, v953, v954, v955, v956, v957, v958, v959, v960, v961, v962, v963, v964, v965, v966, v967, v968, v969, v970, v971, v972, v973, v974, v975, v976, v977, v978, v979, v980, v981, v982, v983, v984, v985, v986, v987, v988, v989, v990, v991, v992, v993, v994, v995, v996, v997, v998, v999, v1000, v1001, v1002, v1003, v1004, v1005, v1006, v1007, v1008, v1009, v1010, v1011, v1012, v1013, v1014, v1015, v1016, v1017, v1018, v1019, v1020, v1021, v1022, v1023, v1024, v1025, v1026, v1027, v1028, v1029, v1030, v1031, v1032, v1033, v1034, v1035, v1036, v1037, v1038, v1039, v1040, v1041, v1042, v1043, v1044, v1045, v1046, v1047, v1048, v1049, v1050, v1051, v1052, v1053, v1054, v1055, v1056, v1057, v1058, v1059, v1060, v1061, v1062, v1063, v1064, v1065, v1066, v1067, v1068, v1069, v1070, v1071, v1072, v1073, v1074, v1075, v1076, v1077, v1078, v1079, v1080, v1081, v1082, v1083, v1084, v1085, v1086, v1087, v1088, v1089, v1090, v1091, v1092, v1093, v1094, v1095, v1096, v1097, v1098, v1099, v1100, v1101, v1102, v1103, v1104, v1105, v1106, v1107, v1108, v1109, v1110, v1111, v1112, v1113, v1114, v1115, v1116, v1117, v1118, v1119, v1120, v1121, v1122, v1123, v1124, v1125, v1126, v1127, v1128, v1129, v1130, v1131, v1132, v1133, v1134, v1135, v1136, v1137, v1138, v1139, v1140, v1141, v1142, v1143, v1144, v1145, v1146, v1147, v1148, v1149, v1150, v1151, v1152, v1153, v1154, v1155, v1156, v1157, v1158, v1159, v1160, v1161, v1162, v1163, v1164, v1165, v1166, v1167, v1168, v1169, v1170, v1171, v1172, v1173, v1174, v1175, v1176, v1177, v1178, v1179, v1180, v1181, v1182, v1183, v1184, v1185, v1186, v1187, v1188, v1189, v1190, v1191, v1192, v1193, v1194, v1195, v1196, v1197, v1198, v1199, v1200, v1201, v1202, v1203, v1204, v1205, v1206, v1207, v1208, v1209, v1210, v1211, v1212, v1213, v1214, v1215, v1216, v1217, v1218, v1219, v1220, v1221, v1222, v1223, v1224, v1225, v1226, v1227, v1228, v1229, v1230, v1231, v1232, v1233, v1234, v1235, v1236, v1237, v1238, v1239, v1240, v1241, v1242, v1243, v1244, v1245, v1246, v1247, v1248, v1249, v1250, v1251, v1252, v1253, v1254, v1255, v1256, v1257, v1258, v1259, v1260, v1261, v1262, v1263, v1264, v1265, v1266, v1267, v1268, v1269, v1270, v1271, v1272, v1273, v1274, v1275, v1276, v1277, v1278, v1279, v1280, v1281, v1282, v1283, v1284, v1285, v1286, v1287, v1288, v1289, v1290, v1291, v1292, v1293, v1294, v1295, v1296, v1297, v1298, v1299, v1300, v1301, v1302, v1303, v1304, v1305, v1306, v1307, v1308, v1309, v1310, v1311, v1312, v1313, v1314, v1315, v1316, v1317, v1318, v1319, v1320, v1321, v1322, v1323, v1324, v1325, v1326, v1327, v1328, v1329, v1330, v1331, v1332, v1333, v1334, v1335, v1336, v1337, v1338, v1339, v1340, v1341, v1342, v1343, v1344, v1345, v1346, v1347, v1348, v1349, v1350, v1351, v1352, v1353, v1354, v1355, v1356, v1357, v1358, v1359, v1360, v1361, v1362, v1363, v1364, v1365, v1366, v1367, v1368, v1369, v1370, v1371, v1372, v1373, v1374, v1375, v1376, v1377, v1378, v1379, v1380, v1381, v1382, v1383, v1384, v1385, v1386, v1387, v1388, v1389, v1390, v1391, v1392, v1393, v1394, v1395, v1396, v1397, v1398, v1399, v1400, v1401, v1402, v1403, v1404, v1405, v1406, v1407, v1408, v1409, v1410, v1411, v1412, v1413, v1414, v1415, v1416, v1417, v1418, v1419, v1420, v1421, v1422, v1423, v1424, v1425, v1426, v1427, v1428, v1429, v1430, v1431, v1432, v1433, v1434, v1435, v1436, v1437, v1438, v1439, v1440, v1441, v1442, v1443, v1444, v1445, v1446, v1447, v1448, v1449, v1450, v1451, v1452, v1453, v1454, v1455, v1456, v1457, v1458, v1459, v1460, v1461, v1462, v1463, v1464, v1465, v1466, v1467, v1468, v1469, v1470, v1471, v1472, v1473, v1474, v1475, v1476, v1477, v1478, v1479, v1480, v1481, v1482, v1483, v1484, v1485, v1486, v1487, v1488, v1489, v1490, v1491, v1492, v1493, v1494, v1495, v1496, v1497, v1498, v1499, v1500, v1501, v1502, v1503, v1504, v1505,
w0, w1, w2, w3, w4, w5, w6, w7, w8, w9, w10, w11, w12, w13, w14, w15, w16, w17, w18, w19, w20, w21, w22, w23, w24, w25, w26, w27, w28, w29, w30, w31, w32, w33, w34, w35, w36, w37, w38, w39, w40, w41, w42, w43, w44, w45, w46, w47, w48, w49, w50, w51, w52, w53, w54, w55, w56, w57, w58, w59, w60, w61, w62, w63, w64, w65, w66, w67, w68, w69, w70, w71, w72, w73, w74, w75, w76, w77, w78, w79, w80, w81, w82, w83, w84, w85, w86, w87, w88, w89, w90, w91, w92, w93, w94, w95, w96, w97, w98, w99, w100, w101, w102, w103, w104, w105, w106, w107, w108, w109, w110, w111, w112, w113, w114, w115, w116, w117, w118, w119, w120, w121, w122, w123, w124, w125, w126, w127, w128, w129, w130, w131, w132, w133, w134, w135, w136, w137, w138, w139, w140, w141, w142, w143, w144, w145, w146, w147, w148, w149, w150, w151, w152, w153, w154, w155, w156, w157, w158, w159, w160, w161, w162, w163, w164, w165, w166, w167, w168, w169, w170, w171, w172, w173, w174, w175, w176, w177, w178, w179, w180, w181, w182, w183, w184, w185, w186, w187, w188, w189, w190, w191, w192, w193, w194, w195, w196, w197, w198, w199, w200, w201, w202, w203, w204, w205, w206, w207, w208, w209, w210, w211, w212, w213, w214, w215, w216, w217, w218, w219, w220, w221, w222, w223, w224, w225, w226, w227, w228, w229, w230, w231, w232, w233, w234, w235, w236, w237, w238, w239, w240, w241, w242, w243, w244, w245, w246, w247, w248, w249, w250, w251, w252, w253, w254, w255, w256, w257, w258, w259, w260, w261, w262, w263, w264, w265, w266, w267, w268, w269, w270, w271, w272, w273, w274, w275, w276, w277, w278, w279, w280, w281, w282, w283, w284, w285, w286, w287, w288, w289, w290, w291, w292, w293, w294, w295, w296, w297, w298, w299, w300, w301, w302, w303, w304, w305, w306, w307, w308, w309, w310, w311, w312, w313, w314, w315, w316, w317, w318, w319, w320, w321, w322, w323, w324, w325, w326, w327, w328, w329, w330, w331, w332, w333, w334, w335, w336, w337, w338, w339, w340, w341, w342, w343, w344, w345, w346, w347, w348, w349, w350, w351, w352, w353, w354, w355, w356, w357, w358, w359, w360, w361, w362, w363, w364, w365, w366, w367, w368, w369, w370, w371, w372, w373, w374, w375, w376, w377, w378, w379, w380, w381, w382, w383, w384, w385, w386, w387, w388, w389, w390, w391, w392, w393, w394, w395, w396, w397, w398, w399, w400, w401, w402, w403, w404, w405, w406, w407, w408, w409, w410, w411, w412, w413, w414, w415, w416, w417, w418, w419, w420, w421, w422, w423, w424, w425, w426, w427, w428, w429, w430, w431, w432, w433, w434, w435, w436, w437, w438, w439, w440, w441, w442, w443, w444, w445, w446, w447, w448, w449, w450, w451, w452, w453, w454, w455, w456, w457, w458, w459, w460, w461, w462, w463, w464, w465, w466, w467, w468, w469, w470, w471, w472, w473, w474, w475, w476, w477, w478, w479, w480, w481, w482, w483, w484, w485, w486, w487, w488, w489, w490, w491, w492, w493, w494, w495, w496, w497, w498, w499, w500, w501, w502, w503, w504, w505, w506, w507, w508, w509, w510, w511, w512, w513, w514, w515, w516, w517, w518, w519, w520, w521, w522, w523, w524, w525, w526, w527, w528, w529, w530, w531, w532, w533, w534, w535, w536, w537, w538, w539, w540, w541, w542, w543, w544, w545, w546, w547, w548, w549, w550, w551, w552, w553, w554, w555, w556, w557, w558, w559, w560, w561, w562, w563, w564, w565, w566, w567, w568, w569, w570, w571, w572, w573, w574, w575, w576, w577, w578, w579, w580, w581, w582, w583, w584, w585, w586, w587, w588, w589, w590, w591, w592, w593, w594, w595, w596, w597, w598, w599, w600, w601, w602, w603, w604, w605, w606, w607, w608, w609, w610, w611, w612, w613, w614, w615, w616, w617, w618, w619, w620, w621, w622, w623, w624, w625, w626, w627, w628, w629, w630, w631, w632, w633, w634, w635, w636, w637, w638, w639, w640, w641, w642, w643, w644, w645, w646, w647, w648, w649, w650, w651, w652, w653, w654, w655, w656, w657, w658, w659, w660, w661, w662, w663, w664, w665, w666, w667, w668, w669, w670, w671, w672, w673, w674, w675, w676, w677, w678, w679, w680, w681, w682, w683, w684, w685, w686, w687, w688, w689, w690, w691, w692, w693, w694, w695, w696, w697, w698, w699, w700, w701, w702, w703, w704, w705, w706, w707, w708, w709, w710, w711, w712, w713, w714, w715, w716, w717, w718, w719, w720, w721, w722, w723, w724, w725, w726, w727, w728, w729, w730, w731, w732, w733, w734, w735, w736, w737, w738, w739, w740, w741, w742, w743, w744, w745, w746, w747, w748, w749, w750, w751, w752, w753, w754, w755, w756, w757, w758, w759, w760, w761, w762, w763, w764, w765, w766, w767, w768, w769, w770, w771, w772, w773, w774, w775, w776, w777, w778, w779, w780, w781, w782, w783, w784, w785, w786, w787, w788, w789, w790, w791, w792, w793, w794, w795, w796, w797, w798, w799, w800, w801, w802, w803, w804, w805, w806, w807, w808, w809, w810, w811, w812, w813, w814, w815, w816, w817, w818, w819, w820, w821, w822, w823, w824, w825, w826, w827, w828, w829, w830, w831, w832, w833, w834, w835, w836, w837, w838, w839, w840, w841, w842, w843, w844, w845, w846, w847, w848, w849, w850, w851, w852, w853, w854, w855, w856, w857, w858, w859, w860, w861, w862, w863, w864, w865, w866, w867, w868, w869, w870, w871, w872, w873, w874, w875, w876, w877, w878, w879, w880, w881, w882, w883, w884, w885, w886, w887, w888, w889, w890, w891, w892, w893, w894, w895, w896, w897, w898, w899, w900, w901, w902, w903, w904, w905, w906, w907, w908, w909, w910, w911, w912, w913, w914, w915, w916, w917, w918, w919, w920, w921, w922, w923, w924, w925, w926, w927, w928, w929, w930, w931, w932, w933, w934, w935, w936, w937, w938, w939, w940, w941, w942, w943, w944, w945, w946, w947, w948, w949, w950, w951, w952, w953, w954, w955, w956, w957, w958, w959, w960, w961, w962, w963, w964, w965, w966, w967, w968, w969, w970, w971, w972, w973, w974, w975, w976, w977, w978, w979, w980, w981, w982, w983, w984, w985, w986, w987, w988, w989, w990, w991, w992, w993, w994, w995, w996, w997, w998, w999, w1000, w1001, w1002, w1003, w1004, w1005, w1006, w1007, w1008, w1009, w1010, w1011, w1012, w1013, w1014, w1015, w1016, w1017, w1018, w1019, w1020, w1021, w1022, w1023, w1024, w1025, w1026, w1027, w1028, w1029, w1030, w1031, w1032, w1033, w1034, w1035, w1036, w1037, w1038, w1039, w1040, w1041, w1042, w1043, w1044, w1045, w1046, w1047, w1048, w1049, w1050, w1051, w1052, w1053, w1054, w1055, w1056, w1057, w1058, w1059, w1060, w1061, w1062, w1063, w1064, w1065, w1066, w1067, w1068, w1069, w1070, w1071, w1072, w1073, w1074, w1075, w1076, w1077, w1078, w1079, w1080, w1081, w1082, w1083, w1084, w1085, w1086, w1087, w1088, w1089, w1090, w1091, w1092, w1093, w1094, w1095, w1096, w1097, w1098, w1099, w1100, w1101, w1102, w1103, w1104, w1105, w1106, w1107, w1108, w1109, w1110, w1111, w1112, w1113, w1114, w1115, w1116, w1117, w1118, w1119, w1120, w1121, w1122, w1123, w1124, w1125, w1126, w1127, w1128, w1129, w1130, w1131, w1132, w1133, w1134, w1135, w1136, w1137, w1138, w1139, w1140, w1141, w1142, w1143, w1144, w1145, w1146, w1147, w1148, w1149, w1150, w1151, w1152, w1153, w1154, w1155, w1156, w1157, w1158, w1159, w1160, w1161, w1162, w1163, w1164, w1165, w1166, w1167, w1168, w1169, w1170, w1171, w1172, w1173, w1174, w1175, w1176, w1177, w1178, w1179, w1180, w1181, w1182, w1183, w1184, w1185, w1186, w1187, w1188, w1189, w1190, w1191, w1192, w1193, w1194, w1195, w1196, w1197, w1198, w1199, w1200, w1201, w1202, w1203, w1204, w1205, w1206, w1207, w1208, w1209, w1210, w1211, w1212, w1213, w1214, w1215, w1216, w1217, w1218, w1219, w1220, w1221, w1222, w1223, w1224, w1225, w1226, w1227, w1228, w1229, w1230, w1231, w1232, w1233, w1234, w1235, w1236, w1237, w1238, w1239, w1240, w1241, w1242, w1243, w1244, w1245, w1246, w1247, w1248, w1249, w1250, w1251, w1252, w1253, w1254, w1255, w1256, w1257, w1258, w1259, w1260, w1261, w1262, w1263, w1264, w1265, w1266, w1267, w1268, w1269, w1270, w1271, w1272, w1273, w1274, w1275, w1276, w1277, w1278, w1279, w1280, w1281, w1282, w1283, w1284, w1285, w1286, w1287, w1288, w1289, w1290, w1291, w1292, w1293, w1294, w1295, w1296, w1297, w1298, w1299, w1300, w1301, w1302, w1303, w1304, w1305, w1306, w1307, w1308, w1309, w1310, w1311, w1312, w1313, w1314, w1315, w1316, w1317, w1318, w1319, w1320, w1321, w1322, w1323, w1324, w1325, w1326, w1327, w1328, w1329, w1330, w1331, w1332, w1333, w1334, w1335, w1336, w1337, w1338, w1339, w1340, w1341, w1342, w1343, w1344, w1345, w1346, w1347, w1348, w1349, w1350, w1351, w1352, w1353, w1354, w1355, w1356, w1357, w1358, w1359, w1360, w1361, w1362, w1363, w1364, w1365, w1366, w1367, w1368, w1369, w1370, w1371, w1372, w1373, w1374, w1375, w1376, w1377, w1378, w1379, w1380, w1381, w1382, w1383, w1384, w1385, w1386, w1387, w1388, w1389, w1390, w1391, w1392, w1393, w1394, w1395, w1396, w1397, w1398, w1399, w1400, w1401, w1402, w1403, w1404, w1405, w1406, w1407, w1408, w1409, w1410, w1411, w1412, w1413, w1414, w1415, w1416, w1417, w1418, w1419, w1420, w1421, w1422, w1423, w1424, w1425, w1426, w1427, w1428, w1429, w1430, w1431, w1432, w1433, w1434, w1435, w1436, w1437, w1438, w1439, w1440, w1441, w1442, w1443, w1444, w1445, w1446, w1447, w1448, w1449, w1450, w1451, w1452, w1453, w1454, w1455, w1456, w1457, w1458, w1459, w1460, w1461, w1462, w1463, w1464, w1465, w1466, w1467, w1468, w1469, w1470, w1471, w1472, w1473, w1474, w1475, w1476, w1477, w1478, w1479, w1480, w1481, w1482, w1483, w1484, w1485, w1486, w1487, w1488, w1489, w1490, w1491, w1492, w1493, w1494, w1495, w1496, w1497, w1498, w1499, w1500, w1501, w1502, w1503, w1504, w1505, w1506, w1507, w1508, w1509, w1510, w1511, w1512, w1513, w1514, w1515, w1516, w1517, w1518, w1519, w1520, w1521, w1522, w1523, w1524, w1525, w1526, w1527, w1528, w1529, w1530, w1531, w1532, w1533, w1534, w1535, w1536, w1537, w1538, w1539, w1540, w1541, w1542, w1543, w1544, w1545, w1546, w1547, w1548, w1549, w1550, w1551, w1552, w1553, w1554, w1555, w1556, w1557, w1558, w1559, w1560, w1561, w1562, w1563, w1564, w1565, w1566, w1567, w1568, w1569, w1570, w1571, w1572, w1573, w1574, w1575, w1576, w1577, w1578, w1579, w1580, w1581, w1582, w1583, w1584, w1585, w1586, w1587, w1588, w1589, w1590, w1591, w1592, w1593, w1594, w1595, w1596, w1597, w1598, w1599, w1600, w1601, w1602, w1603, w1604, w1605, w1606, w1607, w1608, w1609, w1610, w1611, w1612, w1613, w1614, w1615, w1616, w1617, w1618, w1619, w1620, w1621, w1622, w1623, w1624, w1625, w1626, w1627, w1628, w1629, w1630, w1631, w1632, w1633, w1634, w1635, w1636, w1637, w1638, w1639, w1640, w1641, w1642, w1643, w1644, w1645, w1646, w1647, w1648, w1649, w1650, w1651, w1652, w1653, w1654, w1655, w1656, w1657, w1658, w1659, w1660, w1661, w1662, w1663, w1664, w1665, w1666, w1667, w1668, w1669, w1670, w1671, w1672, w1673, w1674, w1675, w1676, w1677, w1678, w1679, w1680, w1681, w1682, w1683, w1684, w1685, w1686, w1687, w1688, w1689, w1690, w1691, w1692, w1693, w1694, w1695, w1696, w1697, w1698, w1699, w1700, w1701, w1702, w1703, w1704, w1705, w1706, w1707, w1708, w1709, w1710, w1711, w1712, w1713, w1714, w1715, w1716, w1717, w1718, w1719, w1720, w1721, w1722, w1723, w1724, w1725, w1726, w1727, w1728, w1729, w1730, w1731, w1732, w1733, w1734, w1735, w1736, w1737, w1738, w1739, w1740, w1741, w1742, w1743, w1744, w1745, w1746, w1747, w1748, w1749, w1750, w1751, w1752, w1753, w1754, w1755, w1756, w1757, w1758, w1759, w1760, w1761, w1762, w1763, w1764, w1765, w1766, w1767, w1768, w1769, w1770, w1771, w1772, w1773, w1774, w1775, w1776, w1777, w1778, w1779, w1780, w1781, w1782, w1783, w1784, w1785, w1786, w1787, w1788, w1789, w1790, w1791, w1792, w1793, w1794, w1795, w1796, w1797, w1798, w1799, w1800, w1801, w1802, w1803, w1804, w1805, w1806, w1807, w1808, w1809, w1810, w1811, w1812, w1813, w1814, w1815, w1816, w1817, w1818, w1819, w1820, w1821, w1822, w1823, w1824, w1825, w1826, w1827, w1828, w1829, w1830, w1831, w1832, w1833, w1834, w1835, w1836, w1837, w1838, w1839, w1840, w1841, w1842, w1843, w1844, w1845, w1846, w1847, w1848, w1849, w1850, w1851, w1852, w1853, w1854, w1855, w1856, w1857, w1858, w1859, w1860, w1861, w1862, w1863, w1864, w1865, w1866, w1867, w1868, w1869, w1870, w1871, w1872, w1873, w1874, w1875, w1876, w1877, w1878, w1879, w1880, w1881, w1882, w1883, w1884, w1885, w1886, w1887, w1888, w1889, w1890, w1891, w1892, w1893, w1894, w1895, w1896, w1897, w1898, w1899, w1900, w1901, w1902, w1903, w1904, w1905, w1906, w1907, w1908, w1909, w1910, w1911, w1912, w1913, w1914, w1915, w1916, w1917, w1918, w1919, w1920, w1921, w1922, w1923, w1924, w1925, w1926, w1927, w1928, w1929, w1930, w1931, w1932, w1933, w1934, w1935, w1936, w1937, w1938, w1939, w1940, w1941, w1942, w1943, w1944, w1945, w1946, w1947, w1948, w1949, w1950, w1951, w1952, w1953, w1954, w1955, w1956, w1957, w1958, w1959, w1960, w1961, w1962, w1963, w1964, w1965, w1966, w1967, w1968, w1969, w1970, w1971, w1972, w1973, w1974, w1975, w1976, w1977, w1978, w1979, w1980, w1981, w1982, w1983, w1984, w1985, w1986, w1987, w1988, w1989, w1990, w1991, w1992, w1993, w1994, w1995, w1996, w1997, w1998, w1999, w2000, w2001, w2002, w2003, w2004, w2005, w2006, w2007, w2008, w2009, w2010, w2011, w2012, w2013, w2014, w2015, w2016, w2017, w2018, w2019, w2020, w2021, w2022, w2023, w2024, w2025, w2026, w2027, w2028, w2029, w2030, w2031, w2032, w2033, w2034, w2035, w2036, w2037, w2038, w2039, w2040, w2041, w2042, w2043, w2044, w2045, w2046, w2047, w2048, w2049, w2050, w2051, w2052, w2053, w2054, w2055, w2056, w2057, w2058, w2059, w2060, w2061, w2062, w2063, w2064, w2065, w2066, w2067, w2068, w2069, w2070, w2071, w2072, w2073, w2074, w2075, w2076, w2077, w2078, w2079, w2080, w2081, w2082, w2083, w2084, w2085, w2086, w2087, w2088, w2089, w2090, w2091, w2092, w2093, w2094, w2095, w2096, w2097, w2098, w2099, w2100, w2101, w2102, w2103, w2104, w2105, w2106, w2107, w2108, w2109, w2110, w2111, w2112, w2113, w2114, w2115, w2116, w2117, w2118, w2119, w2120, w2121, w2122, w2123, w2124, w2125, w2126, w2127, w2128, w2129, w2130, w2131, w2132, w2133, w2134, w2135, w2136, w2137, w2138, w2139, w2140, w2141, w2142, w2143, w2144, w2145, w2146, w2147, w2148, w2149, w2150, w2151, w2152, w2153, w2154, w2155, w2156, w2157, w2158, w2159, w2160, w2161, w2162, w2163, w2164, w2165, w2166, w2167, w2168, w2169, w2170, w2171, w2172, w2173, w2174, w2175, w2176, w2177, w2178, w2179, w2180, w2181, w2182, w2183, w2184, w2185, w2186, w2187, w2188, w2189, w2190, w2191, w2192, w2193, w2194, w2195, w2196, w2197, w2198, w2199, w2200, w2201, w2202, w2203, w2204, w2205, w2206, w2207, w2208, w2209, w2210, w2211, w2212, w2213, w2214, w2215, w2216, w2217, w2218, w2219, w2220, w2221, w2222, w2223, w2224, w2225, w2226, w2227, w2228, w2229, w2230, w2231, w2232, w2233, w2234, w2235, w2236, w2237, w2238, w2239, w2240, w2241, w2242, w2243, w2244, w2245, w2246, w2247, w2248, w2249, w2250, w2251, w2252, w2253, w2254, w2255, w2256, w2257, w2258, w2259, w2260, w2261, w2262, w2263, w2264, w2265, w2266, w2267, w2268, w2269, w2270, w2271, w2272, w2273, w2274, w2275, w2276, w2277, w2278, w2279, w2280, w2281, w2282, w2283, w2284, w2285, w2286, w2287, w2288, w2289, w2290, w2291, w2292, w2293, w2294, w2295, w2296, w2297, w2298, w2299, w2300, w2301, w2302, w2303, w2304, w2305, w2306, w2307, w2308, w2309, w2310, w2311, w2312, w2313, w2314, w2315, w2316, w2317, w2318, w2319, w2320, w2321, w2322, w2323, w2324, w2325, w2326, w2327, w2328, w2329, w2330, w2331, w2332, w2333, w2334, w2335, w2336, w2337, w2338, w2339, w2340, w2341, w2342, w2343, w2344, w2345, w2346, w2347, w2348, w2349, w2350, w2351, w2352, w2353, w2354, w2355, w2356, w2357, w2358, w2359, w2360, w2361, w2362, w2363, w2364, w2365, w2366, w2367, w2368, w2369, w2370, w2371, w2372, w2373, w2374, w2375, w2376, w2377, w2378, w2379, w2380, w2381, w2382, w2383, w2384, w2385, w2386, w2387, w2388, w2389, w2390, w2391, w2392, w2393, w2394, w2395, w2396, w2397, w2398, w2399, w2400, w2401, w2402, w2403, w2404, w2405, w2406, w2407, w2408, w2409, w2410, w2411, w2412, w2413, w2414, w2415, w2416, w2417, w2418, w2419, w2420, w2421, w2422, w2423, w2424, w2425, w2426, w2427, w2428, w2429, w2430, w2431, w2432, w2433, w2434, w2435, w2436, w2437, w2438, w2439, w2440, w2441, w2442, w2443, w2444, w2445, w2446, w2447, w2448, w2449, w2450, w2451, w2452, w2453, w2454, w2455, w2456, w2457, w2458, w2459, w2460, w2461, w2462, w2463, w2464, w2465, w2466, w2467, w2468, w2469, w2470, w2471, w2472, w2473, w2474, w2475, w2476, w2477, w2478, w2479, w2480, w2481, w2482, w2483, w2484, w2485, w2486, w2487, w2488, w2489, w2490, w2491, w2492, w2493, w2494, w2495, w2496, w2497, w2498, w2499, w2500, w2501, w2502, w2503, w2504, w2505, w2506, w2507, w2508, w2509, w2510, w2511, w2512, w2513, w2514, w2515, w2516, w2517, w2518, w2519, w2520, w2521, w2522, w2523, w2524, w2525, w2526, w2527, w2528, w2529, w2530, w2531, w2532, w2533, w2534, w2535, w2536, w2537, w2538, w2539, w2540, w2541, w2542, w2543, w2544, w2545, w2546, w2547, w2548, w2549, w2550, w2551, w2552, w2553, w2554, w2555, w2556, w2557, w2558, w2559, w2560, w2561, w2562, w2563, w2564, w2565, w2566, w2567, w2568, w2569, w2570, w2571, w2572, w2573, w2574, w2575, w2576, w2577, w2578, w2579, w2580, w2581, w2582, w2583, w2584, w2585, w2586, w2587, w2588, w2589, w2590, w2591, w2592, w2593, w2594, w2595, w2596, w2597, w2598, w2599, w2600, w2601, w2602, w2603, w2604, w2605, w2606, w2607, w2608, w2609, w2610, w2611, w2612, w2613, w2614, w2615, w2616, w2617, w2618, w2619, w2620, w2621, w2622, w2623, w2624, w2625, w2626, w2627, w2628, w2629, w2630, w2631, w2632, w2633, w2634, w2635, w2636, w2637, w2638, w2639, w2640, w2641, w2642, w2643, w2644, w2645, w2646, w2647, w2648, w2649, w2650, w2651, w2652, w2653, w2654, w2655, w2656, w2657, w2658, w2659, w2660, w2661, w2662, w2663, w2664, w2665, w2666, w2667, w2668, w2669, w2670, w2671, w2672, w2673, w2674, w2675, w2676, w2677, w2678, w2679, w2680, w2681, w2682, w2683, w2684, w2685, w2686, w2687, w2688, w2689, w2690, w2691, w2692, w2693, w2694, w2695, w2696, w2697, w2698, w2699, w2700, w2701, w2702, w2703, w2704, w2705, w2706, w2707, w2708, w2709, w2710, w2711, w2712, w2713, w2714, w2715, w2716, w2717, w2718, w2719, w2720, w2721, w2722, w2723, w2724, w2725, w2726, w2727, w2728, w2729, w2730, w2731, w2732, w2733, w2734, w2735, w2736, w2737, w2738, w2739, w2740, w2741, w2742, w2743, w2744, w2745, w2746, w2747, w2748, w2749, w2750, w2751, w2752, w2753, w2754, w2755, w2756, w2757, w2758, w2759, w2760, w2761, w2762, w2763, w2764, w2765, w2766, w2767, w2768, w2769, w2770, w2771, w2772, w2773, w2774, w2775, w2776, w2777, w2778, w2779, w2780, w2781, w2782, w2783, w2784, w2785, w2786, w2787, w2788, w2789, w2790, w2791, w2792, w2793, w2794, w2795, w2796, w2797, w2798, w2799, w2800, w2801, w2802, w2803, w2804, w2805, w2806, w2807, w2808, w2809, w2810, w2811, w2812, w2813, w2814, w2815, w2816, w2817, w2818, w2819, w2820, w2821, w2822, w2823, w2824, w2825, w2826, w2827, w2828, w2829, w2830, w2831, w2832, w2833, w2834, w2835, w2836, w2837, w2838, w2839, w2840, w2841, w2842, w2843, w2844, w2845, w2846, w2847, w2848, w2849, w2850, w2851, w2852, w2853, w2854, w2855, w2856, w2857, w2858, w2859, w2860, w2861, w2862, w2863, w2864, w2865, w2866, w2867, w2868, w2869, w2870, w2871, w2872, w2873, w2874, w2875, w2876, w2877, w2878, w2879, w2880, w2881, w2882, w2883, w2884, w2885, w2886, w2887, w2888, w2889, w2890, w2891, w2892, w2893, w2894, w2895, w2896, w2897, w2898, w2899, w2900, w2901, w2902, w2903, w2904, w2905, w2906, w2907, w2908, w2909, w2910, w2911, w2912, w2913, w2914, w2915, w2916, w2917, w2918, w2919, w2920, w2921, w2922, w2923, w2924, w2925, w2926, w2927, w2928, w2929, w2930, w2931, w2932, w2933, w2934, w2935, w2936, w2937, w2938, w2939, w2940, w2941, w2942, w2943, w2944, w2945, w2946, w2947, w2948, w2949, w2950, w2951, w2952, w2953, w2954, w2955, w2956, w2957, w2958, w2959, w2960, w2961, w2962, w2963, w2964, w2965, w2966, w2967, w2968, w2969, w2970, w2971, w2972, w2973, w2974, w2975, w2976, w2977, w2978, w2979, w2980, w2981, w2982, w2983, w2984, w2985, w2986, w2987, w2988, w2989, w2990, w2991, w2992, w2993, w2994, w2995, w2996, w2997, w2998, w2999, w3000, w3001, w3002, w3003, w3004, w3005, w3006, w3007, w3008, w3009, w3010, w3011, w3012, w3013, w3014, w3015, w3016, w3017, w3018, w3019, w3020, w3021, w3022, w3023, w3024, w3025, w3026, w3027, w3028, w3029, w3030, w3031, w3032, w3033, w3034, w3035, w3036, w3037, w3038, w3039, w3040, w3041, w3042, w3043, w3044, w3045, w3046, w3047, w3048, w3049, w3050, w3051, w3052, w3053, w3054, w3055, w3056, w3057, w3058, w3059, w3060, w3061, w3062, w3063, w3064, w3065, w3066, w3067, w3068, w3069, w3070, w3071, w3072, w3073, w3074, w3075, w3076, w3077, w3078, w3079, w3080, w3081, w3082, w3083, w3084, w3085, w3086, w3087, w3088, w3089, w3090, w3091, w3092, w3093, w3094, w3095, w3096, w3097, w3098, w3099, w3100, w3101, w3102, w3103, w3104, w3105, w3106, w3107, w3108, w3109, w3110, w3111, w3112, w3113, w3114, w3115, w3116, w3117, w3118, w3119, w3120, w3121, w3122, w3123, w3124, w3125, w3126, w3127, w3128, w3129, w3130, w3131, w3132, w3133, w3134, w3135, w3136, w3137, w3138, w3139, w3140, w3141, w3142, w3143, w3144, w3145, w3146, w3147, w3148, w3149, w3150, w3151, w3152, w3153, w3154, w3155, w3156, w3157, w3158, w3159, w3160, w3161, w3162, w3163, w3164, w3165, w3166, w3167, w3168, w3169, w3170, w3171, w3172, w3173, w3174, w3175, w3176, w3177, w3178, w3179, w3180, w3181, w3182, w3183, w3184, w3185, w3186, w3187, w3188, w3189, w3190, w3191, w3192, w3193, w3194, w3195, w3196, w3197, w3198, w3199, w3200, w3201, w3202, w3203, w3204, w3205, w3206, w3207, w3208, w3209, w3210, w3211, w3212, w3213, w3214, w3215, w3216, w3217, w3218, w3219, w3220, w3221, w3222, w3223, w3224, w3225, w3226, w3227, w3228, w3229, w3230, w3231, w3232, w3233, w3234, w3235, w3236, w3237, w3238, w3239, w3240, w3241, w3242, w3243, w3244, w3245, w3246, w3247, w3248, w3249, w3250, w3251, w3252, w3253, w3254, w3255, w3256, w3257, w3258, w3259, w3260, w3261, w3262, w3263, w3264, w3265, w3266, w3267, w3268, w3269, w3270, w3271, w3272, w3273, w3274, w3275, w3276, w3277, w3278, w3279, w3280, w3281, w3282, w3283, w3284, w3285, w3286, w3287, w3288, w3289, w3290, w3291, w3292, w3293, w3294, w3295, w3296, w3297, w3298, w3299, w3300, w3301, w3302, w3303, w3304, w3305, w3306, w3307, w3308, w3309, w3310, w3311, w3312, w3313, w3314, w3315, w3316, w3317, w3318, w3319, w3320, w3321, w3322, w3323, w3324, w3325, w3326, w3327, w3328, w3329, w3330, w3331, w3332, w3333, w3334, w3335, w3336, w3337, w3338, w3339, w3340, w3341, w3342, w3343, w3344, w3345, w3346, w3347, w3348, w3349, w3350, w3351, w3352, w3353, w3354, w3355, w3356, w3357, w3358, w3359, w3360, w3361, w3362, w3363, w3364, w3365, w3366, w3367, w3368, w3369, w3370, w3371, w3372, w3373, w3374, w3375, w3376, w3377, w3378, w3379, w3380, w3381, w3382, w3383, w3384, w3385, w3386, w3387, w3388, w3389, w3390, w3391, w3392, w3393, w3394, w3395, w3396, w3397, w3398, w3399, w3400, w3401, w3402, w3403, w3404, w3405, w3406, w3407, w3408, w3409, w3410, w3411, w3412, w3413, w3414, w3415, w3416, w3417, w3418, w3419, w3420, w3421, w3422, w3423, w3424, w3425, w3426, w3427, w3428, w3429, w3430, w3431, w3432, w3433, w3434, w3435, w3436, w3437, w3438, w3439, w3440, w3441, w3442, w3443, w3444, w3445, w3446, w3447, w3448, w3449, w3450, w3451, w3452, w3453, w3454, w3455, w3456, w3457, w3458, w3459, w3460, w3461, w3462, w3463, w3464, w3465, w3466, w3467, w3468, w3469, w3470, w3471, w3472, w3473, w3474, w3475, w3476, w3477, w3478, w3479, w3480, w3481, w3482, w3483, w3484, w3485, w3486, w3487, w3488, w3489, w3490, w3491, w3492, w3493, w3494, w3495, w3496, w3497, w3498, w3499, w3500, w3501, w3502, w3503, w3504, w3505, w3506, w3507, w3508, w3509, w3510, w3511, w3512, w3513, w3514, w3515, w3516, w3517, w3518, w3519, w3520, w3521, w3522, w3523, w3524, w3525, w3526, w3527, w3528, w3529, w3530, w3531, w3532, w3533, w3534, w3535, w3536, w3537, w3538, w3539, w3540, w3541, w3542, w3543, w3544, w3545, w3546, w3547, w3548, w3549, w3550, w3551, w3552, w3553, w3554, w3555, w3556, w3557, w3558, w3559, w3560, w3561, w3562, w3563, w3564, w3565, w3566, w3567, w3568, w3569, w3570, w3571, w3572, w3573, w3574, w3575, w3576, w3577, w3578, w3579, w3580, w3581, w3582, w3583, w3584, w3585, w3586, w3587, w3588, w3589, w3590, w3591, w3592, w3593, w3594, w3595, w3596, w3597, w3598, w3599, w3600, w3601, w3602, w3603, w3604, w3605, w3606, w3607, w3608, w3609, w3610, w3611, w3612, w3613, w3614, w3615, w3616, w3617, w3618, w3619, w3620, w3621, w3622, w3623, w3624, w3625, w3626, w3627, w3628, w3629, w3630, w3631, w3632, w3633, w3634, w3635, w3636, w3637, w3638, w3639, w3640, w3641, w3642, w3643, w3644, w3645, w3646, w3647, w3648, w3649, w3650, w3651, w3652, w3653, w3654, w3655, w3656, w3657, w3658, w3659, w3660, w3661, w3662, w3663, w3664, w3665, w3666, w3667, w3668, w3669, w3670, w3671, w3672, w3673, w3674, w3675, w3676, w3677, w3678, w3679, w3680, w3681, w3682, w3683, w3684, w3685, w3686, w3687, w3688, w3689, w3690, w3691, w3692, w3693, w3694, w3695, w3696, w3697, w3698, w3699, w3700, w3701, w3702, w3703, w3704, w3705, w3706, w3707, w3708, w3709, w3710, w3711, w3712, w3713, w3714, w3715, w3716, w3717, w3718, w3719, w3720, w3721, w3722, w3723, w3724, w3725, w3726, w3727, w3728, w3729, w3730, w3731, w3732, w3733, w3734, w3735, w3736, w3737, w3738, w3739, w3740, w3741, w3742, w3743, w3744, w3745, w3746, w3747, w3748, w3749, w3750, w3751, w3752, w3753, w3754, w3755, w3756, w3757, w3758, w3759, w3760, w3761, w3762, w3763, w3764, w3765, w3766, w3767, w3768, w3769, w3770, w3771, w3772, w3773, w3774, w3775, w3776, w3777, w3778, w3779, w3780, w3781, w3782, w3783, w3784, w3785, w3786, w3787, w3788, w3789, w3790, w3791, w3792, w3793, w3794, w3795, w3796, w3797, w3798, w3799, w3800, w3801, w3802, w3803, w3804, w3805, w3806, w3807, w3808, w3809, w3810, w3811, w3812, w3813, w3814, w3815, w3816, w3817, w3818, w3819, w3820, w3821, w3822, w3823, w3824, w3825, w3826, w3827, w3828, w3829, w3830, w3831, w3832, w3833, w3834, w3835, w3836, w3837, w3838, w3839, w3840, w3841, w3842, w3843, w3844, w3845, w3846, w3847, w3848, w3849, w3850, w3851, w3852, w3853, w3854, w3855, w3856, w3857, w3858, w3859, w3860, w3861, w3862, w3863, w3864, w3865, w3866, w3867, w3868, w3869, w3870, w3871, w3872, w3873, w3874, w3875, w3876, w3877, w3878, w3879, w3880, w3881, w3882, w3883, w3884, w3885, w3886, w3887, w3888, w3889, w3890, w3891, w3892, w3893, w3894, w3895, w3896, w3897, w3898, w3899, w3900, w3901, w3902, w3903, w3904, w3905, w3906, w3907, w3908, w3909, w3910, w3911, w3912, w3913, w3914, w3915, w3916, w3917, w3918, w3919, w3920, w3921, w3922, w3923, w3924, w3925, w3926, w3927, w3928, w3929, w3930, w3931, w3932, w3933, w3934, w3935, w3936, w3937, w3938, w3939, w3940, w3941, w3942, w3943, w3944, w3945, w3946, w3947, w3948, w3949, w3950, w3951, w3952, w3953, w3954, w3955, w3956, w3957, w3958, w3959, w3960, w3961, w3962, w3963, w3964, w3965, w3966, w3967, w3968, w3969, w3970, w3971, w3972, w3973, w3974, w3975, w3976, w3977, w3978, w3979, w3980, w3981, w3982, w3983, w3984, w3985, w3986, w3987, w3988, w3989, w3990, w3991, w3992, w3993, w3994, w3995, w3996, w3997, w3998, w3999, w4000, w4001, w4002, w4003, w4004, w4005, w4006, w4007, w4008, w4009, w4010, w4011, w4012, w4013, w4014, w4015, w4016, w4017, w4018, w4019, w4020, w4021, w4022, w4023, w4024, w4025, w4026, w4027, w4028, w4029, w4030, w4031, w4032, w4033, w4034, w4035, w4036, w4037, w4038, w4039, w4040, w4041, w4042, w4043, w4044, w4045, w4046, w4047, w4048, w4049, w4050, w4051, w4052, w4053, w4054, w4055, w4056, w4057, w4058, w4059, w4060, w4061, w4062, w4063, w4064, w4065, w4066, w4067, w4068, w4069, w4070, w4071, w4072, w4073, w4074, w4075, w4076, w4077, w4078, w4079, w4080, w4081, w4082, w4083, w4084, w4085, w4086, w4087, w4088, w4089, w4090, w4091, w4092, w4093, w4094, w4095, w4096, w4097, w4098, w4099, w4100, w4101, w4102, w4103, w4104, w4105, w4106, w4107, w4108, w4109, w4110, w4111, w4112, w4113, w4114, w4115, w4116, w4117, w4118, w4119, w4120, w4121, w4122, w4123, w4124, w4125, w4126, w4127, w4128, w4129, w4130, w4131, w4132, w4133, w4134, w4135, w4136, w4137, w4138, w4139, w4140, w4141, w4142, w4143, w4144, w4145, w4146, w4147, w4148, w4149, w4150, w4151, w4152, w4153, w4154, w4155, w4156, w4157, w4158, w4159, w4160, w4161, w4162, w4163, w4164, w4165, w4166, w4167, w4168, w4169, w4170, w4171, w4172, w4173, w4174, w4175, w4176, w4177, w4178, w4179, w4180, w4181, w4182, w4183, w4184, w4185;
assign w0 = ~w1386 & w1039;
assign v0 = ~(w497 | w2518);
assign w1 = v0;
assign v1 = ~(w1377 | w3149);
assign w2 = v1;
assign v2 = ~(w1970 | w3722);
assign w3 = v2;
assign w4 = (~w1469 & ~w1099) | (~w1469 & w1690) | (~w1099 & w1690);
assign w5 = w426 & ~w1629;
assign w6 = ~pi366 & pi218;
assign v3 = ~(w744 | w1590);
assign w7 = v3;
assign v4 = ~(w1574 | w3030);
assign w8 = v4;
assign v5 = ~(w2583 | w997);
assign w9 = v5;
assign v6 = ~(w566 | w4007);
assign w10 = v6;
assign v7 = ~(w1324 | w83);
assign w11 = v7;
assign w12 = w2484 & ~w442;
assign v8 = ~(w1801 | w2089);
assign w13 = v8;
assign w14 = pi106 & w570;
assign v9 = ~(w2693 | w763);
assign w15 = v9;
assign w16 = w4005 & w3227;
assign v10 = ~(w4121 | w665);
assign w17 = v10;
assign w18 = w2443 & ~w2285;
assign w19 = ~w1996 & w4012;
assign v11 = ~(w2297 | w628);
assign w20 = v11;
assign w21 = ~w2776 & w1555;
assign w22 = pi267 & w2362;
assign v12 = ~(w2289 | w29);
assign w23 = v12;
assign w24 = w871 & ~w445;
assign w25 = w1005 & ~w1342;
assign w26 = w1995 & w2912;
assign w27 = w2602 & w3807;
assign v13 = ~(w2968 | w1182);
assign w28 = v13;
assign v14 = ~(w179 | w3160);
assign w29 = v14;
assign w30 = (pi069 & ~w1654) | (pi069 & w2920) | (~w1654 & w2920);
assign w31 = w350 & ~w1469;
assign v15 = ~(w165 | w425);
assign w32 = v15;
assign w33 = (w2443 & w3477) | (w2443 & w236) | (w3477 & w236);
assign w34 = pi306 & ~pi366;
assign w35 = ~w1806 & w1175;
assign w36 = pi350 & ~pi366;
assign w37 = (w1698 & w429) | (w1698 & w3306) | (w429 & w3306);
assign v16 = ~(w1654 | w1182);
assign w38 = v16;
assign w39 = w2000 & ~w2436;
assign w40 = w1570 & w2218;
assign v17 = ~(w1754 | w3722);
assign w41 = v17;
assign w42 = (w3380 & ~w3606) | (w3380 & w369) | (~w3606 & w369);
assign w43 = w2717 & ~w3317;
assign v18 = ~(w15 | w2484);
assign w44 = v18;
assign w45 = ~w3094 & w1327;
assign v19 = ~(w1900 | w590);
assign w46 = v19;
assign w47 = w1743 & w2455;
assign w48 = ~w1486 & w2530;
assign w49 = w2324 & w2898;
assign v20 = ~(w2966 | w2331);
assign w50 = v20;
assign v21 = ~(w177 | w3252);
assign w51 = v21;
assign w52 = pi189 & w1570;
assign v22 = ~(w1509 | w3455);
assign w53 = v22;
assign v23 = ~(w2615 | w3844);
assign w54 = v23;
assign v24 = ~(w1661 | w3462);
assign w55 = v24;
assign w56 = w15 & w2484;
assign w57 = w2194 & w342;
assign w58 = ~w2646 & w244;
assign w59 = (w1469 & ~w2613) | (w1469 & w3250) | (~w2613 & w3250);
assign v25 = ~(w994 | w3894);
assign w60 = v25;
assign w61 = w2731 & w2395;
assign v26 = ~(w46 | w1893);
assign w62 = v26;
assign w63 = w2420 & ~w89;
assign w64 = w3048 & w732;
assign v27 = ~(w2396 | w2207);
assign w65 = v27;
assign w66 = ~w2646 & w3180;
assign v28 = ~(w3111 | w662);
assign w67 = v28;
assign w68 = (w3505 & w638) | (w3505 & w2399) | (w638 & w2399);
assign w69 = ~w1135 & w2061;
assign w70 = w656 & ~w1607;
assign w71 = w3024 & w1654;
assign w72 = w253 & w3032;
assign w73 = ~w3094 & w3005;
assign v29 = ~(w1957 | w3892);
assign w74 = v29;
assign w75 = w1199 & ~w1102;
assign w76 = w4037 & w1664;
assign w77 = ~w2606 & w946;
assign w78 = ~w3094 & w2100;
assign w79 = pi273 & w2362;
assign w80 = pi134 & ~pi364;
assign w81 = w656 & ~w1782;
assign w82 = ~w513 & w3706;
assign w83 = (~w1469 & ~w2562) | (~w1469 & w139) | (~w2562 & w139);
assign v30 = ~(w3160 | w3858);
assign w84 = v30;
assign w85 = ~pi366 & pi241;
assign w86 = w378 & ~w2459;
assign w87 = pi340 & ~pi366;
assign w88 = w73 & w1469;
assign w89 = w3262 & ~w1089;
assign w90 = w118 & pi047;
assign w91 = ~w1510 & w3803;
assign v31 = ~(w362 | w3478);
assign w92 = v31;
assign w93 = w47 & w643;
assign w94 = w1689 & w1631;
assign v32 = ~(w3685 | w978);
assign w95 = v32;
assign w96 = w2420 & w559;
assign w97 = ~w1071 & w307;
assign v33 = ~(w2304 | w109);
assign w98 = v33;
assign w99 = pi307 & ~pi366;
assign v34 = ~(w1754 | w3277);
assign w100 = v34;
assign v35 = ~(w1918 | w834);
assign w101 = v35;
assign v36 = ~(w3182 | w2104);
assign w102 = v36;
assign v37 = ~(w954 | w3414);
assign w103 = v37;
assign w104 = w1924 & w2910;
assign w105 = w1662 & ~w2832;
assign v38 = ~(w2667 | w1324);
assign w106 = v38;
assign v39 = ~(w4180 | w3205);
assign w107 = v39;
assign v40 = ~(w981 | w3056);
assign w108 = v40;
assign w109 = ~w1987 & w213;
assign v41 = ~(w1642 | w3563);
assign w110 = v41;
assign w111 = w3928 & ~w1469;
assign w112 = w118 & pi054;
assign w113 = pi358 & ~pi366;
assign w114 = w344 & w2153;
assign v42 = ~(w794 | w3878);
assign w115 = v42;
assign w116 = w2825 & w1469;
assign v43 = ~(w2627 | w1535);
assign w117 = v43;
assign w118 = pi366 & pi367;
assign v44 = ~(w994 | w1810);
assign w119 = v44;
assign w120 = pi308 & ~pi366;
assign w121 = ~w138 & w2605;
assign w122 = w3669 & ~w3425;
assign w123 = w271 & w1182;
assign w124 = w1381 & w2659;
assign v45 = ~(w2475 | w3977);
assign w125 = v45;
assign w126 = ~w4049 & w3322;
assign w127 = w2717 & ~w3277;
assign v46 = ~(w1680 | w1898);
assign w128 = v46;
assign w129 = (pi071 & ~w1654) | (pi071 & w3291) | (~w1654 & w3291);
assign v47 = ~(w2643 | w820);
assign w130 = v47;
assign v48 = ~(w2917 | w2068);
assign w131 = v48;
assign w132 = (~w1886 & ~w2830) | (~w1886 & w2183) | (~w2830 & w2183);
assign w133 = pi297 & w2362;
assign w134 = w2587 & w1654;
assign w135 = (~w1089 & ~w2004) | (~w1089 & w2159) | (~w2004 & w2159);
assign w136 = w1473 & w3854;
assign v49 = ~(w334 | w375);
assign w137 = v49;
assign v50 = ~(w1202 | w3121);
assign w138 = v50;
assign w139 = w3144 & ~w1469;
assign v51 = ~(w2799 | w2123);
assign w140 = v51;
assign v52 = ~(w4116 | w3053);
assign w141 = v52;
assign w142 = ~w3658 & w1314;
assign w143 = w2359 & ~w1469;
assign w144 = w1510 & w2764;
assign w145 = ~w3064 & w1714;
assign w146 = ~pi366 & pi247;
assign w147 = ~w1671 & w2788;
assign w148 = ~w3094 & w3428;
assign w149 = ~w1772 & w1260;
assign w150 = (w227 & w3501) | (w227 & w829) | (w3501 & w829);
assign w151 = w118 & pi072;
assign w152 = ~w2046 & w1499;
assign v53 = ~(w1146 | w1144);
assign w153 = v53;
assign v54 = ~(w4038 | w422);
assign w154 = v54;
assign w155 = w2626 & ~w3677;
assign v55 = ~(w4159 | w1955);
assign w156 = v55;
assign v56 = ~(w244 | w3180);
assign w157 = v56;
assign w158 = pi144 & w1570;
assign w159 = w260 & w374;
assign w160 = (w252 & ~w2918) | (w252 & w474) | (~w2918 & w474);
assign w161 = w1443 & w1469;
assign w162 = w2022 & w3628;
assign w163 = w2397 & ~w2769;
assign w164 = (w1024 & ~w2114) | (w1024 & w2639) | (~w2114 & w2639);
assign w165 = ~w15 & w2484;
assign v57 = ~(w1352 | w2277);
assign w166 = v57;
assign v58 = ~(w2451 | w1507);
assign w167 = v58;
assign w168 = w118 & pi057;
assign v59 = ~(w722 | w3328);
assign w169 = v59;
assign w170 = w3094 & w535;
assign w171 = w2717 & ~w1607;
assign w172 = w361 & ~w3626;
assign w173 = w394 & ~w772;
assign w174 = w1610 & w2015;
assign w175 = w435 & w2373;
assign w176 = (pi013 & ~w1654) | (pi013 & w2939) | (~w1654 & w2939);
assign w177 = w2058 & w1628;
assign w178 = w3094 & w904;
assign w179 = ~w45 & w1916;
assign w180 = w1313 & w1654;
assign w181 = w2484 & ~w1539;
assign v60 = ~(w2475 | w1782);
assign w182 = v60;
assign v61 = ~(w1871 | w2118);
assign w183 = v61;
assign w184 = ~w3094 & w3789;
assign w185 = w705 & w2156;
assign w186 = pi264 & w2362;
assign w187 = w2268 & ~w2324;
assign w188 = w2566 & w2330;
assign w189 = w2373 & w3443;
assign v62 = ~(w3277 | w2475);
assign w190 = v62;
assign w191 = w2471 & w1469;
assign v63 = ~(w2938 | w3717);
assign w192 = v63;
assign v64 = ~(w889 | w661);
assign w193 = v64;
assign v65 = ~(w3284 | w3772);
assign w194 = v65;
assign v66 = ~(w2487 | w1507);
assign w195 = v66;
assign v67 = ~(w779 | w2992);
assign w196 = v67;
assign w197 = w4155 & w2686;
assign v68 = ~(w956 | w55);
assign w198 = v68;
assign v69 = ~(w3312 | w3977);
assign w199 = v69;
assign w200 = w354 & ~w1387;
assign w201 = w460 & w2973;
assign w202 = ~w226 & w183;
assign v70 = ~(w2379 | w2808);
assign w203 = v70;
assign w204 = (w1654 & w1670) | (w1654 & w3617) | (w1670 & w3617);
assign w205 = w1570 & w80;
assign w206 = (w1249 & w3342) | (w1249 & w3453) | (w3342 & w3453);
assign v71 = ~(w2936 | w3068);
assign w207 = v71;
assign v72 = ~(w2335 | w57);
assign w208 = v72;
assign w209 = w3094 & w2943;
assign w210 = w2717 & ~w3131;
assign v73 = ~(w708 | w2180);
assign w211 = v73;
assign w212 = w44 & ~w4130;
assign v74 = ~(w2936 | w2539);
assign w213 = v74;
assign w214 = w672 & ~w3565;
assign v75 = ~(w317 | w3113);
assign w215 = v75;
assign w216 = w92 & ~w2133;
assign w217 = w2646 & w244;
assign w218 = w893 & ~w3794;
assign v76 = ~(w2175 | w357);
assign w219 = v76;
assign v77 = ~(w2536 | w2708);
assign w220 = v77;
assign v78 = ~(w409 | w1967);
assign w221 = v78;
assign w222 = w3144 & w1469;
assign v79 = ~(w4038 | w1592);
assign w223 = v79;
assign w224 = w1057 & w3467;
assign v80 = ~(w882 | w2200);
assign w225 = v80;
assign v81 = ~(w2748 | w3361);
assign w226 = v81;
assign v82 = ~(w2473 | w450);
assign w227 = v82;
assign v83 = ~(w3259 | w398);
assign w228 = v83;
assign w229 = w3769 & w3191;
assign w230 = ~w1145 & w2564;
assign v84 = ~(w2393 | w3008);
assign w231 = v84;
assign w232 = ~w2570 & w3793;
assign v85 = ~(w250 | w2889);
assign w233 = v85;
assign w234 = ~w3041 & w3669;
assign v86 = ~(w371 | w2052);
assign w235 = v86;
assign w236 = w424 & w2443;
assign w237 = w1638 & w3522;
assign v87 = ~(w3312 | w357);
assign w238 = v87;
assign v88 = ~(w4160 | w1842);
assign w239 = v88;
assign w240 = ~pi366 & pi210;
assign w241 = ~w128 & w3159;
assign v89 = ~(w170 | w1986);
assign w242 = v89;
assign w243 = w3883 & w3571;
assign v90 = ~(w82 | w264);
assign w244 = v90;
assign w245 = w2759 & w1469;
assign v91 = ~(w2175 | w3317);
assign w246 = v91;
assign v92 = ~(w2287 | w1095);
assign w247 = v92;
assign w248 = ~w802 & w1304;
assign w249 = w1358 & ~w3729;
assign w250 = ~w871 & w1635;
assign v93 = ~(w3608 | w3257);
assign w251 = v93;
assign w252 = (w2998 & w328) | (w2998 & w977) | (w328 & w977);
assign w253 = w1932 & w3705;
assign w254 = w2646 & ~w244;
assign w255 = w3945 & w1469;
assign w256 = (w1654 & w1029) | (w1654 & w1947) | (w1029 & w1947);
assign v94 = ~(w3506 | w3245);
assign w257 = v94;
assign w258 = w2690 & ~w3026;
assign w259 = (w3838 & ~w3585) | (w3838 & w1064) | (~w3585 & w1064);
assign v95 = ~(w3362 | w2413);
assign w260 = v95;
assign v96 = ~(w2109 | w1965);
assign w261 = v96;
assign v97 = ~(w1754 | w2412);
assign w262 = v97;
assign w263 = w1571 & w1046;
assign w264 = w513 & ~w3706;
assign w265 = (w2764 & ~w3803) | (w2764 & w144) | (~w3803 & w144);
assign w266 = w705 & w2630;
assign w267 = w4120 & w1005;
assign w268 = ~w1992 & w2350;
assign w269 = w1804 & w3244;
assign w270 = w2717 & ~w1633;
assign w271 = (~w1469 & ~w4127) | (~w1469 & w143) | (~w4127 & w143);
assign w272 = pi248 & w2362;
assign w273 = (w324 & ~w1689) | (w324 & w969) | (~w1689 & w969);
assign w274 = ~pi366 & pi197;
assign v98 = ~(w2175 | w3343);
assign w275 = v98;
assign w276 = (w1469 & ~w567) | (w1469 & w1185) | (~w567 & w1185);
assign w277 = w3094 & w461;
assign v99 = ~(w2799 | w2085);
assign w278 = v99;
assign w279 = w3585 & w405;
assign w280 = w45 & w1469;
assign v100 = ~(w2178 | w2082);
assign w281 = v100;
assign w282 = w118 & pi024;
assign v101 = ~(w2799 | w1667);
assign w283 = v101;
assign w284 = w705 & w414;
assign w285 = w2046 & ~w3179;
assign w286 = w3159 & ~w2000;
assign v102 = ~(w1072 | w2169);
assign w287 = v102;
assign v103 = ~(w4038 | w1164);
assign w288 = v103;
assign w289 = w766 & w619;
assign w290 = w194 & w2854;
assign w291 = w1179 & w2188;
assign w292 = (w1318 & w2817) | (w1318 & w1572) | (w2817 & w1572);
assign w293 = w656 & ~w422;
assign w294 = w141 & ~w2315;
assign w295 = w3262 & w1089;
assign v104 = ~(w907 | w270);
assign w296 = v104;
assign w297 = w1716 & w1654;
assign w298 = (w1654 & w2246) | (w1654 & w1228) | (w2246 & w1228);
assign w299 = w1469 & w2690;
assign w300 = w2099 & ~w2642;
assign w301 = (w2989 & ~w653) | (w2989 & w3558) | (~w653 & w3558);
assign w302 = w1182 & ~w3605;
assign w303 = ~w2268 & w2324;
assign w304 = ~w2322 & w1328;
assign v105 = ~(w1140 | w3312);
assign w305 = v105;
assign w306 = w1830 & ~w920;
assign w307 = w771 & w3035;
assign w308 = (w1469 & ~w947) | (w1469 & w2847) | (~w947 & w2847);
assign w309 = w3370 & w3154;
assign w310 = w3069 & w3756;
assign w311 = ~w3022 & w1154;
assign w312 = w3189 & w3972;
assign w313 = (w1654 & w2674) | (w1654 & w2512) | (w2674 & w2512);
assign v106 = ~(w179 | w3312);
assign w314 = v106;
assign w315 = w1774 & w1499;
assign v107 = ~(w1059 | w1733);
assign w316 = v107;
assign v108 = ~(w1754 | w3131);
assign w317 = v108;
assign w318 = (w1853 & ~w3069) | (w1853 & w1236) | (~w3069 & w1236);
assign w319 = w451 & ~w911;
assign w320 = w1028 & w2330;
assign v109 = ~(w1117 | w2326);
assign w321 = v109;
assign w322 = w730 & w1654;
assign w323 = w118 & pi052;
assign w324 = ~w2553 & w2112;
assign v110 = ~(w1502 | w2139);
assign w325 = v110;
assign v111 = ~(w698 | w1758);
assign w326 = v111;
assign w327 = ~w3710 & w3669;
assign w328 = w3068 & ~w3180;
assign w329 = ~w847 & w2378;
assign w330 = w1297 & w1654;
assign w331 = ~w2070 & w2125;
assign w332 = w1830 & ~w557;
assign v112 = ~(w1550 | w2590);
assign w333 = v112;
assign w334 = ~w2542 & w331;
assign w335 = w64 & w2996;
assign w336 = ~w580 & w600;
assign w337 = ~w2373 & w3179;
assign w338 = w950 & ~w867;
assign w339 = w3262 & w2440;
assign w340 = w806 & w846;
assign w341 = ~w173 & w1083;
assign w342 = w4047 & w2502;
assign w343 = w1334 & w511;
assign v113 = ~(w738 | w1765);
assign w344 = v113;
assign w345 = w1272 & w1626;
assign w346 = w1249 & ~w781;
assign v114 = ~(w2475 | w3414);
assign w347 = v114;
assign w348 = ~w1222 & w4091;
assign w349 = w1330 & ~w335;
assign w350 = ~w3094 & w2192;
assign w351 = w1008 & w289;
assign w352 = w595 & w748;
assign w353 = w1654 & w570;
assign v115 = ~(w3436 | w2948);
assign w354 = v115;
assign w355 = w2397 & ~w1541;
assign w356 = pi046 & w353;
assign w357 = ~w3394 & w567;
assign w358 = w705 & w2012;
assign v116 = ~(w954 | w149);
assign w359 = v116;
assign w360 = ~w425 & w2461;
assign v117 = ~(w3137 | w4131);
assign w361 = v117;
assign w362 = (w1654 & w2447) | (w1654 & w3758) | (w2447 & w3758);
assign w363 = ~w2099 & w2642;
assign w364 = (~w1662 & w2892) | (~w1662 & w3413) | (w2892 & w3413);
assign w365 = ~w2140 & w3246;
assign w366 = w991 & ~w1132;
assign w367 = (w2594 & ~w709) | (w2594 & w2903) | (~w709 & w2903);
assign v118 = ~(w4146 | w3860);
assign w368 = v118;
assign w369 = ~w2965 & w3380;
assign w370 = ~w2606 & w4171;
assign v119 = ~(w1970 | w3414);
assign w371 = v119;
assign w372 = ~w1447 & w932;
assign v120 = ~(w785 | w2193);
assign w373 = v120;
assign v121 = ~(w1694 | w2054);
assign w374 = v121;
assign w375 = ~w3551 & w292;
assign w376 = (w1469 & ~w1260) | (w1469 & w1974) | (~w1260 & w1974);
assign w377 = w3714 & w1877;
assign w378 = w4000 & w3547;
assign v122 = ~(w1757 | w4133);
assign w379 = v122;
assign v123 = ~(w1177 | w1529);
assign w380 = v123;
assign v124 = ~(w204 | w1568);
assign w381 = v124;
assign v125 = ~(w603 | w1984);
assign w382 = v125;
assign w383 = ~w775 & w1539;
assign v126 = ~(w3530 | w2384);
assign w384 = v126;
assign v127 = ~(w3264 | w3970);
assign w385 = v127;
assign v128 = ~(w4148 | w3170);
assign w386 = v128;
assign w387 = w2405 & w3689;
assign w388 = ~w3094 & w3519;
assign w389 = w1469 & w2626;
assign v129 = ~(w2876 | w1934);
assign w390 = v129;
assign w391 = w2523 & w1332;
assign v130 = ~(w4038 | w1881);
assign w392 = v130;
assign w393 = w3094 & w3636;
assign v131 = ~(w433 | w2394);
assign w394 = v131;
assign w395 = pi179 & w1570;
assign w396 = ~pi366 & pi237;
assign w397 = ~pi366 & pi228;
assign w398 = ~w2759 & w251;
assign w399 = w571 & w2201;
assign w400 = w3196 & w4014;
assign v132 = ~(w2848 | w1927);
assign w401 = v132;
assign v133 = ~(w2317 | w2536);
assign w402 = v133;
assign w403 = w3216 & ~w1762;
assign w404 = w130 & w3888;
assign w405 = (~w492 & w2223) | (~w492 & w2886) | (w2223 & w2886);
assign w406 = w3064 & ~w1714;
assign w407 = ~w2172 & w3447;
assign v134 = ~(w3792 | w2811);
assign w408 = v134;
assign v135 = ~(w3160 | w3168);
assign w409 = v135;
assign w410 = w891 & w377;
assign w411 = pi184 & w1570;
assign w412 = w2860 & w3207;
assign w413 = ~w2501 & w798;
assign w414 = w1570 & w2585;
assign w415 = ~w834 & w2487;
assign w416 = w2082 & w2706;
assign v136 = ~(w216 | w1402);
assign w417 = v136;
assign w418 = (w1654 & w3502) | (w1654 & w463) | (w3502 & w463);
assign v137 = ~(w868 | w283);
assign w419 = v137;
assign w420 = w1081 & ~w157;
assign w421 = w2244 & ~w1525;
assign w422 = ~w3740 & w242;
assign w423 = w1663 & w325;
assign w424 = (w1469 & ~w709) | (w1469 & w1485) | (~w709 & w1485);
assign w425 = w15 & ~w4074;
assign v138 = ~(w874 | w2747);
assign w426 = v138;
assign w427 = w1762 & w2079;
assign v139 = ~(w4087 | w2475);
assign w428 = v139;
assign w429 = w3068 & ~w2031;
assign w430 = w946 & w303;
assign w431 = pi312 & ~pi366;
assign w432 = w1830 & ~w3848;
assign v140 = ~(w349 | w2614);
assign w433 = v140;
assign w434 = (w1654 & w3631) | (w1654 & w2597) | (w3631 & w2597);
assign v141 = ~(w2923 | w3063);
assign w435 = v141;
assign v142 = ~(w2878 | w1679);
assign w436 = v142;
assign v143 = ~(w2527 | w3115);
assign w437 = v143;
assign w438 = w2690 & ~w3679;
assign w439 = w851 & ~w3764;
assign v144 = ~(w1318 | w304);
assign w440 = v144;
assign w441 = w2743 & w1654;
assign v145 = ~(w3274 | w4081);
assign w442 = v145;
assign w443 = w2831 & w1021;
assign v146 = ~(w3160 | w923);
assign w444 = v146;
assign v147 = ~(w4010 | w162);
assign w445 = v147;
assign w446 = ~w3856 & w1688;
assign v148 = ~(w2175 | w1533);
assign w447 = v148;
assign w448 = ~w3928 & w767;
assign w449 = (~w943 & w3518) | (~w943 & w2032) | (w3518 & w2032);
assign w450 = (pi126 & ~w1654) | (pi126 & w1280) | (~w1654 & w1280);
assign w451 = w2122 & ~w285;
assign v149 = ~(w1673 | w4038);
assign w452 = v149;
assign v150 = ~(w2475 | w149);
assign w453 = v150;
assign w454 = (~w162 & w871) | (~w162 & w1307) | (w871 & w1307);
assign w455 = w466 & w983;
assign w456 = (w943 & w1699) | (w943 & w1162) | (w1699 & w1162);
assign v151 = ~(w3929 | w1970);
assign w457 = v151;
assign w458 = w3408 & w3215;
assign w459 = ~w269 & w2099;
assign w460 = w616 & w2066;
assign w461 = pi334 & ~pi366;
assign v152 = ~(w2000 | w128);
assign w462 = v152;
assign w463 = w4179 & w1654;
assign v153 = ~(w1346 | w1265);
assign w464 = v153;
assign w465 = w1199 & ~w919;
assign w466 = w1385 & w2559;
assign w467 = pi191 & ~pi364;
assign w468 = w705 & w2002;
assign w469 = w1565 & w1851;
assign v154 = ~(w256 | w1730);
assign w470 = v154;
assign v155 = ~(w3216 | w2628);
assign w471 = v155;
assign w472 = w2717 & ~w1104;
assign w473 = w1830 & ~w3943;
assign w474 = w4056 & w252;
assign w475 = w3086 & w3127;
assign v156 = ~(w1970 | w3131);
assign w476 = v156;
assign w477 = pi173 & ~pi364;
assign v157 = ~(w3837 | w3955);
assign w478 = v157;
assign v158 = ~(w1673 | w3878);
assign w479 = v158;
assign w480 = w2484 & ~w2523;
assign w481 = w3042 & w1322;
assign w482 = w2626 & ~w119;
assign w483 = w2268 & w660;
assign w484 = ~w3094 & w85;
assign w485 = w656 & ~w3131;
assign w486 = ~w3067 & w613;
assign w487 = (w1469 & ~w3440) | (w1469 & w3668) | (~w3440 & w3668);
assign v159 = ~(w1318 | w1038);
assign w488 = v159;
assign v160 = ~(w4022 | w453);
assign w489 = v160;
assign w490 = ~w1245 & w3542;
assign v161 = ~(w318 | w310);
assign w491 = v161;
assign w492 = w984 & ~w320;
assign w493 = w118 & pi127;
assign v162 = ~(w4038 | w3977);
assign w494 = v162;
assign w495 = w1920 & ~w1469;
assign v163 = ~(w1139 | w433);
assign w496 = v163;
assign w497 = ~w48 & w2717;
assign w498 = ~w1920 & w108;
assign v164 = ~(w3303 | w230);
assign w499 = v164;
assign v165 = ~(w3159 | w128);
assign w500 = v165;
assign w501 = ~w1607 & w1830;
assign w502 = w9 & w2620;
assign w503 = (w1654 & w4002) | (w1654 & w3374) | (w4002 & w3374);
assign w504 = ~w3094 & w1206;
assign w505 = w2055 & w3305;
assign w506 = pi324 & ~pi366;
assign w507 = pi287 & w2362;
assign w508 = w705 & w4129;
assign v166 = ~(w4159 | w2085);
assign w509 = v166;
assign w510 = (w1469 & ~w4170) | (w1469 & w1350) | (~w4170 & w1350);
assign v167 = ~(w3753 | w3174);
assign w511 = v167;
assign w512 = w1120 & w2777;
assign w513 = w3989 & w1232;
assign w514 = (w2215 & ~w2055) | (w2215 & w1911) | (~w2055 & w1911);
assign v168 = ~(w3312 | w2412);
assign w515 = v168;
assign w516 = (pi087 & ~w1654) | (pi087 & w4026) | (~w1654 & w4026);
assign w517 = w1740 & w3409;
assign v169 = ~(w630 | w2098);
assign w518 = v169;
assign v170 = ~(w2140 | w2022);
assign w519 = v170;
assign w520 = w4150 & w3419;
assign v171 = ~(w3457 | w3973);
assign w521 = v171;
assign v172 = ~(w2833 | w133);
assign w522 = v172;
assign v173 = ~(w3160 | w920);
assign w523 = v173;
assign v174 = ~(w2475 | w1533);
assign w524 = v174;
assign w525 = ~pi366 & pi239;
assign w526 = pi326 & ~pi366;
assign w527 = pi321 & ~pi366;
assign w528 = ~w3094 & w2344;
assign v175 = ~(w1104 | w3905);
assign w529 = v175;
assign w530 = w378 & ~w211;
assign w531 = ~w717 & w1873;
assign w532 = ~pi366 & pi212;
assign v176 = ~(w2175 | w2412);
assign w533 = v176;
assign w534 = w2717 & ~w179;
assign w535 = pi356 & ~pi366;
assign v177 = ~(w1970 | w542);
assign w536 = v177;
assign w537 = w3150 & w3863;
assign w538 = w1473 & w2177;
assign v178 = ~(w3379 | w3760);
assign w539 = v178;
assign v179 = ~(w3160 | w1533);
assign w540 = v179;
assign w541 = w2717 & ~w3385;
assign w542 = ~w2283 & w1217;
assign v180 = ~(w3905 | w3722);
assign w543 = v180;
assign v181 = ~(w2640 | w3894);
assign w544 = v181;
assign v182 = ~(w2244 | w2610);
assign w545 = v182;
assign w546 = ~w3094 & w146;
assign v183 = ~(w1661 | w3426);
assign w547 = v183;
assign w548 = ~pi366 & pi222;
assign w549 = ~w2325 & w3887;
assign w550 = w1830 & ~w1955;
assign w551 = ~w1022 & w1436;
assign v184 = ~(w3149 | w3470);
assign w552 = v184;
assign w553 = w118 & pi067;
assign v185 = ~(w1025 | w2418);
assign w554 = v185;
assign w555 = w2563 & w2306;
assign w556 = pi349 & ~pi366;
assign w557 = ~w2001 & w1268;
assign v186 = ~(w1754 | w794);
assign w558 = v186;
assign w559 = w2315 & w964;
assign v187 = ~(w2740 | w3776);
assign w560 = v187;
assign v188 = ~(pi360 | pi367);
assign w561 = v188;
assign w562 = (~w1469 & ~w117) | (~w1469 & w1713) | (~w117 & w1713);
assign v189 = ~(w4159 | w91);
assign w563 = v189;
assign w564 = w2690 & ~w65;
assign w565 = w3262 & w964;
assign w566 = w1005 & ~w2288;
assign v190 = ~(w1426 | w1106);
assign w567 = v190;
assign w568 = w2207 & w838;
assign v191 = ~(w3842 | w2248);
assign w569 = v191;
assign v192 = ~(w1570 | w118);
assign w570 = v192;
assign w571 = w2321 & w3834;
assign w572 = (~w1469 & ~w2678) | (~w1469 & w3237) | (~w2678 & w3237);
assign v193 = ~(w3160 | w448);
assign w573 = v193;
assign v194 = ~(w1220 | w3840);
assign w574 = v194;
assign v195 = ~(w4052 | w4089);
assign w575 = v195;
assign w576 = w2956 & ~w3665;
assign w577 = w4119 & w389;
assign w578 = w7 & w1490;
assign w579 = (w1469 & ~w478) | (w1469 & w1362) | (~w478 & w1362);
assign w580 = w2717 & ~w1444;
assign v196 = ~(w4016 | w1828);
assign w581 = v196;
assign w582 = ~w4140 & w2692;
assign v197 = ~(w1594 | w3637);
assign w583 = v197;
assign w584 = pi299 & w2362;
assign v198 = ~(w3160 | w1881);
assign w585 = v198;
assign w586 = ~w3279 & w531;
assign w587 = w3094 & w1311;
assign w588 = w118 & pi031;
assign w589 = ~w2774 & w2922;
assign w590 = ~w2968 & w410;
assign w591 = pi259 & w2362;
assign w592 = ~w419 & w3380;
assign v199 = ~(w4159 | w542);
assign w593 = v199;
assign v200 = ~(w4159 | w1592);
assign w594 = v200;
assign w595 = w840 & w1420;
assign v201 = ~(w2328 | w3335);
assign w596 = v201;
assign w597 = (w1626 & w2298) | (w1626 & w345) | (w2298 & w345);
assign v202 = ~(w1324 | w562);
assign w598 = v202;
assign v203 = ~(w3161 | w22);
assign w599 = v203;
assign v204 = ~(w2844 | w4079);
assign w600 = v204;
assign w601 = w3995 & w1086;
assign v205 = ~(w479 | w2008);
assign w602 = v205;
assign w603 = w2717 & ~w3848;
assign v206 = ~(w2475 | w3263);
assign w604 = v206;
assign w605 = w3208 & w606;
assign v207 = ~(w2499 | w3610);
assign w606 = v207;
assign v208 = ~(w359 | w4173);
assign w607 = v208;
assign w608 = w3094 & w2490;
assign w609 = w378 & ~w674;
assign v209 = ~(w3588 | w1635);
assign w610 = v209;
assign v210 = ~(w3696 | w572);
assign w611 = v210;
assign w612 = (~w991 & ~w1250) | (~w991 & w2267) | (~w1250 & w2267);
assign w613 = ~w3159 & w539;
assign w614 = ~pi048 & w353;
assign w615 = ~w391 & w3830;
assign w616 = w3833 & w4118;
assign v211 = ~(w1970 | w4087);
assign w617 = v211;
assign v212 = ~(w846 | w1343);
assign w618 = v212;
assign v213 = ~(w1737 | w678);
assign w619 = v213;
assign w620 = w1976 & w1469;
assign w621 = w2367 & w2507;
assign w622 = (w2993 & ~w4150) | (w2993 & w3429) | (~w4150 & w3429);
assign v214 = ~(w1604 | w3259);
assign w623 = v214;
assign v215 = ~(w754 | w2953);
assign w624 = v215;
assign w625 = ~w4017 & w3773;
assign w626 = ~w1318 & w2108;
assign w627 = w2397 & ~w1991;
assign v216 = ~(w2799 | w1164);
assign w628 = v216;
assign v217 = ~(w3312 | w3131);
assign w629 = v217;
assign v218 = ~(w2799 | w1444);
assign w630 = v218;
assign w631 = w118 & pi043;
assign w632 = (w3318 & ~w478) | (w3318 & w852) | (~w478 & w852);
assign w633 = w1733 & w3669;
assign v219 = ~(w1661 | w3943);
assign w634 = v219;
assign w635 = w571 & w94;
assign w636 = (~w1758 & ~w2367) | (~w1758 & w326) | (~w2367 & w326);
assign v220 = ~(w3180 | w254);
assign w637 = v220;
assign w638 = w846 & w3759;
assign w639 = (pi030 & ~w1654) | (pi030 & w3211) | (~w1654 & w3211);
assign w640 = (~w381 & w263) | (~w381 & w4151) | (w263 & w4151);
assign w641 = ~w3129 & w1471;
assign v221 = ~(w2936 | w3919);
assign w642 = v221;
assign w643 = w839 & ~w3422;
assign v222 = ~(w1300 | w43);
assign w644 = v222;
assign v223 = ~(w2007 | w4167);
assign w645 = v223;
assign w646 = (w1654 & w2778) | (w1654 & w2930) | (w2778 & w2930);
assign w647 = w1834 & w3518;
assign w648 = w15 & w4074;
assign w649 = w677 & ~w311;
assign v224 = ~(w1019 | w2839);
assign w650 = v224;
assign v225 = ~(w1104 | w1661);
assign w651 = v225;
assign w652 = w400 & w2795;
assign w653 = ~w2871 & w2661;
assign w654 = w656 & ~w398;
assign v226 = ~(w1695 | w3792);
assign w655 = v226;
assign v227 = ~(w897 | w1464);
assign w656 = v227;
assign w657 = ~w2632 & w2604;
assign w658 = w2126 & ~w2528;
assign w659 = ~w1469 & w2397;
assign w660 = ~w2893 & w4047;
assign w661 = (w1469 & ~w2562) | (w1469 & w222) | (~w2562 & w222);
assign v228 = ~(w1661 | w1667);
assign w662 = v228;
assign w663 = w838 & ~w3054;
assign w664 = (pi098 & ~w1654) | (pi098 & w2111) | (~w1654 & w2111);
assign w665 = (~w1343 & w4138) | (~w1343 & w618) | (w4138 & w618);
assign v229 = ~(w2123 | w1970);
assign w666 = v229;
assign v230 = ~(w2136 | w550);
assign w667 = v230;
assign w668 = ~w3094 & w3939;
assign w669 = w3158 & w1388;
assign v231 = ~(w3259 | w2209);
assign w670 = v231;
assign v232 = ~(w2799 | w149);
assign w671 = v232;
assign w672 = w2006 & w1273;
assign w673 = ~w1277 & w1973;
assign v233 = ~(w3921 | w562);
assign w674 = v233;
assign v234 = ~(w627 | w3148);
assign w675 = v234;
assign w676 = w2936 & w2082;
assign v235 = ~(w3537 | w2875);
assign w677 = v235;
assign w678 = w1830 & ~w657;
assign w679 = ~w1803 & w1582;
assign w680 = pi076 & w353;
assign v236 = ~(w1546 | w1171);
assign w681 = v236;
assign v237 = ~(w3259 | w1444);
assign w682 = v237;
assign w683 = w856 & w23;
assign w684 = w1139 & ~w3188;
assign v238 = ~(w1844 | w2059);
assign w685 = v238;
assign w686 = w118 & pi110;
assign w687 = w3546 & ~w1287;
assign v239 = ~(w651 | w2934);
assign w688 = v239;
assign w689 = ~pi366 & pi211;
assign w690 = w2086 & ~w2914;
assign w691 = (w3380 & ~w174) | (w3380 & w592) | (~w174 & w592);
assign w692 = w3509 & ~w1469;
assign w693 = w1910 & w2901;
assign v240 = ~(w999 | w3095);
assign w694 = v240;
assign v241 = ~(w48 | w4159);
assign w695 = v241;
assign v242 = ~(w3160 | w4105);
assign w696 = v242;
assign w697 = ~w1709 & w348;
assign w698 = w800 & w3068;
assign w699 = w3094 & w113;
assign w700 = (~w1469 & ~w3803) | (~w1469 & w1797) | (~w3803 & w1797);
assign v243 = ~(w2799 | w557);
assign w701 = v243;
assign w702 = w198 & w2047;
assign w703 = w2964 & w1654;
assign v244 = ~(w452 | w3725);
assign w704 = v244;
assign w705 = ~pi365 & w2357;
assign w706 = w3992 & w3622;
assign v245 = ~(w1657 | w2972);
assign w707 = v245;
assign w708 = (w1469 & ~w3803) | (w1469 & w2115) | (~w3803 & w2115);
assign v246 = ~(w1323 | w79);
assign w709 = v246;
assign v247 = ~(w1721 | w2756);
assign w710 = v247;
assign v248 = ~(w48 | w2175);
assign w711 = v248;
assign w712 = w3094 & w34;
assign v249 = ~(w447 | w1914);
assign w713 = v249;
assign v250 = ~(w3180 | w217);
assign w714 = v250;
assign w715 = w4073 & ~w2626;
assign w716 = ~w538 & w2535;
assign w717 = w1114 & w1705;
assign w718 = ~w800 & w2646;
assign w719 = ~w1492 & w3360;
assign w720 = w3102 & w3987;
assign v251 = ~(w1878 | w2423);
assign w721 = v251;
assign v252 = ~(w1604 | w3312);
assign w722 = v252;
assign w723 = ~w3094 & w3190;
assign w724 = w1531 & w1398;
assign w725 = ~w3094 & w6;
assign w726 = w118 & pi016;
assign v253 = ~(w3312 | w3943);
assign w727 = v253;
assign v254 = ~(w2475 | w1444);
assign w728 = v254;
assign w729 = (w1318 & w1549) | (w1318 & w3220) | (w1549 & w3220);
assign w730 = pi153 & w1570;
assign w731 = ~w2383 & w3913;
assign w732 = w3868 & w1355;
assign w733 = w2247 & ~w1469;
assign w734 = ~w4049 & w3601;
assign w735 = (w1469 & ~w2678) | (w1469 & w620) | (~w2678 & w620);
assign w736 = w4074 & ~w138;
assign w737 = w433 & ~w1113;
assign v255 = ~(w3878 | w1633);
assign w738 = v255;
assign v256 = ~(w1754 | w1782);
assign w739 = v256;
assign w740 = w1631 & ~w2993;
assign w741 = w1486 & w1469;
assign w742 = pi341 & ~pi366;
assign v257 = ~(w1231 | w433);
assign w743 = v257;
assign v258 = ~(w2475 | w398);
assign w744 = v258;
assign w745 = (w1654 & w1423) | (w1654 & w134) | (w1423 & w134);
assign w746 = w3669 & ~w1100;
assign w747 = w2058 & w3145;
assign w748 = w4128 & ~w324;
assign w749 = w1830 & ~w4087;
assign w750 = (w187 & ~w1227) | (w187 & w3935) | (~w1227 & w3935);
assign v259 = ~(w2300 | w1377);
assign w751 = v259;
assign w752 = pi137 & ~pi364;
assign w753 = ~w1447 & w3216;
assign w754 = w3094 & w2561;
assign w755 = (pi005 & ~w1654) | (pi005 & w3465) | (~w1654 & w3465);
assign w756 = (w1005 & w3342) | (w1005 & w267) | (w3342 & w267);
assign w757 = w4070 & w1662;
assign w758 = w354 & ~w183;
assign w759 = (pi023 & ~w1654) | (pi023 & w1052) | (~w1654 & w1052);
assign v260 = ~(w3081 | w1169);
assign w760 = v260;
assign w761 = pi346 & ~pi366;
assign w762 = w1005 & ~w1866;
assign w763 = w1101 & w93;
assign w764 = (w1654 & w1744) | (w1654 & w441) | (w1744 & w441);
assign v261 = ~(w970 | w4103);
assign w765 = v261;
assign v262 = ~(w2522 | w3976);
assign w766 = v262;
assign v263 = ~(w3877 | w2265);
assign w767 = v263;
assign w768 = (w2461 & w1061) | (w2461 & w803) | (w1061 & w803);
assign v264 = ~(w2307 | w2915);
assign w769 = v264;
assign w770 = (pi090 & ~w1654) | (pi090 & w3909) | (~w1654 & w3909);
assign v265 = ~(w4065 | w138);
assign w771 = v265;
assign w772 = w871 & w3483;
assign w773 = ~w1626 & w1779;
assign w774 = w3191 & w3724;
assign w775 = (~w2076 & w2408) | (~w2076 & w3936) | (w2408 & w3936);
assign v266 = ~(w451 | w3827);
assign w776 = v266;
assign w777 = w876 & ~w2398;
assign v267 = ~(w3847 | w1936);
assign w778 = v267;
assign w779 = w2443 & ~w2971;
assign v268 = ~(w1480 | w1854);
assign w780 = v268;
assign v269 = ~(w4120 | w271);
assign w781 = v269;
assign v270 = ~(w4038 | w3385);
assign w782 = v270;
assign w783 = pi020 & w570;
assign v271 = ~(w1715 | w1964);
assign w784 = v271;
assign w785 = (w1654 & w2818) | (w1654 & w3142) | (w2818 & w3142);
assign v272 = ~(w2042 | w609);
assign w786 = v272;
assign w787 = w67 & w3497;
assign w788 = (w1034 & ~w709) | (w1034 & w3829) | (~w709 & w3829);
assign w789 = w3514 & w2658;
assign v273 = ~(w48 | w3905);
assign w790 = v273;
assign v274 = ~(w1754 | w91);
assign w791 = v274;
assign w792 = w1278 & ~w3079;
assign v275 = ~(w1754 | w1604);
assign w793 = v275;
assign w794 = ~w3144 & w2562;
assign w795 = w2315 & ~w89;
assign v276 = ~(w4159 | w557);
assign w796 = v276;
assign w797 = w2717 & ~w3426;
assign v277 = ~(w2461 | w425);
assign w798 = v277;
assign w799 = w656 & ~w2085;
assign v278 = ~(w2545 | w1917);
assign w800 = v278;
assign w801 = w1303 & w2495;
assign w802 = w1616 & w1293;
assign w803 = w425 & w2461;
assign w804 = w656 & ~w4105;
assign w805 = ~w3094 & w396;
assign w806 = w3159 & w539;
assign w807 = (w2484 & ~w3128) | (w2484 & w3607) | (~w3128 & w3607);
assign v279 = ~(w2022 | w4010);
assign w808 = v279;
assign w809 = pi038 & w570;
assign w810 = (w1005 & w3696) | (w1005 & w2338) | (w3696 & w2338);
assign v280 = ~(w271 | w1425);
assign w811 = v280;
assign w812 = w3094 & w2648;
assign v281 = ~(w2812 | w2372);
assign w813 = v281;
assign v282 = ~(w2117 | w1129);
assign w814 = v282;
assign w815 = w1830 & ~w3426;
assign v283 = ~(w3312 | w2085);
assign w816 = v283;
assign v284 = ~(w1741 | w4003);
assign w817 = v284;
assign w818 = pi128 & w1570;
assign w819 = w528 & w1469;
assign w820 = ~w2080 & w3228;
assign w821 = ~w1455 & w3859;
assign v285 = ~(w2191 | w3836);
assign w822 = v285;
assign w823 = w1830 & ~w357;
assign v286 = ~(w1970 | w923);
assign w824 = v286;
assign w825 = ~w4108 & w849;
assign v287 = ~(w1989 | w3534);
assign w826 = v287;
assign v288 = ~(w3216 | w2668);
assign w827 = v288;
assign w828 = (w1654 & w2991) | (w1654 & w3698) | (w2991 & w3698);
assign w829 = w63 & w3157;
assign v289 = ~(w2175 | w498);
assign w830 = v289;
assign v290 = ~(w4025 | w472);
assign w831 = v290;
assign v291 = ~(w3027 | w1978);
assign w832 = v291;
assign w833 = (w324 & ~w595) | (w324 & w1901) | (~w595 & w1901);
assign w834 = ~w4065 & w138;
assign v292 = ~(w59 | w3187);
assign w835 = v292;
assign w836 = ~w76 & w641;
assign v293 = ~(w48 | w1661);
assign w837 = v293;
assign w838 = w4000 & w2006;
assign v294 = ~(w2303 | w3268);
assign w839 = v294;
assign v295 = ~(w1982 | w939);
assign w840 = v295;
assign w841 = w1250 & w850;
assign w842 = ~w2123 & w656;
assign v296 = ~(w3878 | w1881);
assign w843 = v296;
assign v297 = ~(w2088 | w4);
assign w844 = v297;
assign w845 = (~w1469 & ~w2530) | (~w1469 & w975) | (~w2530 & w975);
assign w846 = w2000 & ~w128;
assign w847 = ~w2053 & w1981;
assign v298 = ~(w1794 | w1545);
assign w848 = v298;
assign w849 = ~w768 & w878;
assign w850 = (~w991 & ~w2194) | (~w991 & w3441) | (~w2194 & w3441);
assign w851 = w15 & w4065;
assign w852 = w388 & w3318;
assign w853 = ~w1007 & w3084;
assign v299 = ~(w3469 | w2710);
assign w854 = v299;
assign v300 = ~(w1617 | w3952);
assign w855 = v300;
assign v301 = ~(w1685 | w1094);
assign w856 = v301;
assign v302 = ~(w1970 | w422);
assign w857 = v302;
assign w858 = pi077 & w570;
assign w859 = ~w1469 & w3630;
assign v303 = ~(w3281 | w3292);
assign w860 = v303;
assign w861 = (~w3068 & ~w58) | (~w3068 & w207) | (~w58 & w207);
assign w862 = ~w2995 & w147;
assign w863 = ~w3159 & w128;
assign v304 = ~(w212 | w3752);
assign w864 = v304;
assign w865 = (w2330 & ~w1722) | (w2330 & w188) | (~w1722 & w188);
assign w866 = w3158 & w3206;
assign v305 = ~(w1749 | w1733);
assign w867 = v305;
assign v306 = ~(w1673 | w1661);
assign w868 = v306;
assign w869 = ~w4158 & w3331;
assign v307 = ~(w884 | w2281);
assign w870 = v307;
assign v308 = ~(w519 | w3588);
assign w871 = v308;
assign w872 = w3838 & w2037;
assign w873 = ~w1658 & w237;
assign v309 = ~(w226 | w183);
assign w874 = v309;
assign v310 = ~(w756 | w1538);
assign w875 = v310;
assign v311 = ~(w2609 | w2284);
assign w876 = v311;
assign v312 = ~(w954 | w3131);
assign w877 = v312;
assign w878 = (~w2487 & w2560) | (~w2487 & w1465) | (w2560 & w1465);
assign w879 = ~w3262 & w141;
assign v313 = ~(w3905 | w3168);
assign w880 = v313;
assign w881 = w1009 & w2850;
assign w882 = w1249 & ~w2549;
assign w883 = pi187 & w1570;
assign w884 = w575 & ~w3345;
assign w885 = (pi067 & ~w1654) | (pi067 & w553) | (~w1654 & w553);
assign v314 = ~(w3850 | w4001);
assign w886 = v314;
assign w887 = w2128 & ~w2358;
assign w888 = ~w860 & w3084;
assign w889 = (~w1469 & ~w2613) | (~w1469 & w1309) | (~w2613 & w1309);
assign v315 = ~(w372 | w2469);
assign w890 = v315;
assign w891 = w1215 & w3474;
assign v316 = ~(w1611 | w182);
assign w892 = v316;
assign v317 = ~(w1876 | w1760);
assign w893 = v317;
assign w894 = (pi044 & ~w1654) | (pi044 & w3251) | (~w1654 & w3251);
assign w895 = ~w1631 & w2993;
assign w896 = ~w3262 & w2610;
assign v318 = ~(w1469 | w950);
assign w897 = v318;
assign w898 = ~w162 & w1458;
assign w899 = w672 & ~w3993;
assign w900 = pi171 & w1570;
assign w901 = (~w1469 & ~w2407) | (~w1469 & w1859) | (~w2407 & w1859);
assign v319 = ~(w1104 | w2175);
assign w902 = v319;
assign w903 = (pi072 & ~w1654) | (pi072 & w151) | (~w1654 & w151);
assign w904 = pi338 & ~pi366;
assign v320 = ~(w3878 | w3131);
assign w905 = v320;
assign w906 = ~w871 & w1579;
assign v321 = ~(w48 | w3878);
assign w907 = v321;
assign v322 = ~(w428 | w1542);
assign w908 = v322;
assign w909 = pi166 & w1570;
assign v323 = ~(w1295 | w2497);
assign w910 = v323;
assign w911 = w46 & ~w4099;
assign w912 = (pi001 & ~w1654) | (pi001 & w3550) | (~w1654 & w3550);
assign v324 = ~(w646 | w770);
assign w913 = v324;
assign v325 = ~(w1852 | w857);
assign w914 = v325;
assign v326 = ~(w3475 | w1711);
assign w915 = v326;
assign w916 = w2690 & w3269;
assign v327 = ~(w1970 | w498);
assign w917 = v327;
assign w918 = w4171 & w2267;
assign v328 = ~(w1749 | w1878);
assign w919 = v328;
assign w920 = ~w528 & w1793;
assign v329 = ~(w2623 | w41);
assign w921 = v329;
assign w922 = (w2179 & ~w2349) | (w2179 & w3675) | (~w2349 & w3675);
assign w923 = ~w3775 & w1569;
assign v330 = ~(w59 | w83);
assign w924 = v330;
assign w925 = ~w3850 & w3534;
assign v331 = ~(w3953 | w663);
assign w926 = v331;
assign v332 = ~(w523 | w2456);
assign w927 = v332;
assign w928 = ~w446 & w239;
assign w929 = pi170 & w1570;
assign w930 = pi364 & pi365;
assign v333 = ~(w2799 | w1533);
assign w931 = v333;
assign w932 = w3216 & ~w3179;
assign w933 = w118 & pi017;
assign v334 = ~(w1970 | w3263);
assign w934 = v334;
assign v335 = ~(w954 | w2412);
assign w935 = v335;
assign w936 = w1245 & w226;
assign v336 = ~(w2175 | w3168);
assign w937 = v336;
assign w938 = w2443 & ~w2963;
assign v337 = ~(w3259 | w3385);
assign w939 = v337;
assign w940 = (w1469 & ~w3673) | (w1469 & w4063) | (~w3673 & w4063);
assign w941 = pi280 & w2362;
assign w942 = w2028 & w2258;
assign v338 = ~(w2476 | w2067);
assign w943 = v338;
assign w944 = w321 & w1070;
assign w945 = pi254 & w2362;
assign w946 = w4171 & ~w2129;
assign v339 = ~(w1532 | w1585);
assign w947 = v339;
assign v340 = ~(w3259 | w3105);
assign w948 = v340;
assign w949 = w324 & w4015;
assign w950 = w2006 & w3118;
assign w951 = w834 & w44;
assign w952 = w3620 & w3532;
assign w953 = (w3630 & w3342) | (w3630 & w1925) | (w3342 & w1925);
assign v341 = ~(w859 | w1895);
assign w954 = v341;
assign w955 = w1469 & w1005;
assign v342 = ~(w2475 | w3343);
assign w956 = v342;
assign v343 = ~(w887 | w3072);
assign w957 = v343;
assign v344 = ~(w2305 | w2529);
assign w958 = v344;
assign v345 = ~(w2244 | w1853);
assign w959 = v345;
assign w960 = w2663 & w131;
assign v346 = ~(w3262 | w2315);
assign w961 = v346;
assign w962 = ~w3094 & w240;
assign w963 = (pi064 & ~w1654) | (pi064 & w1013) | (~w1654 & w1013);
assign v347 = ~(w3979 | w3270);
assign w964 = v347;
assign w965 = ~w1707 & w1526;
assign w966 = w1317 & ~w2859;
assign w967 = w3159 & w2000;
assign w968 = ~w56 & w2487;
assign w969 = (w2173 & w949) | (w2173 & w2558) | (w949 & w2558);
assign v348 = ~(w3878 | w91);
assign w970 = v348;
assign w971 = ~w4113 & w1764;
assign w972 = pi150 & w1570;
assign w973 = ~w2779 & w3479;
assign w974 = (w1469 & ~w117) | (w1469 & w4044) | (~w117 & w4044);
assign w975 = w1486 & ~w1469;
assign w976 = pi302 & w2362;
assign w977 = w3068 & ~w2936;
assign v349 = ~(w3905 | w1633);
assign w978 = v349;
assign v350 = ~(w917 | w2237);
assign w979 = v350;
assign w980 = (w1654 & w3219) | (w1654 & w3171) | (w3219 & w3171);
assign w981 = w3094 & w2217;
assign w982 = w725 & ~w1469;
assign w983 = w3548 & w2629;
assign v351 = ~(w3957 | w1576);
assign w984 = v351;
assign v352 = ~(w2324 | w3199);
assign w985 = v352;
assign v353 = ~(w1661 | w4087);
assign w986 = v353;
assign w987 = w101 & w3348;
assign v354 = ~(w2799 | w1607);
assign w988 = v354;
assign w989 = w162 & w2574;
assign w990 = w1188 & w681;
assign v355 = ~(w406 | w145);
assign w991 = v355;
assign v356 = ~(w727 | w782);
assign w992 = v356;
assign w993 = w3334 & ~w1469;
assign w994 = (~w1469 & ~w4139) | (~w1469 & w31) | (~w4139 & w31);
assign w995 = (w2397 & w940) | (w2397 & w3971) | (w940 & w3971);
assign v357 = ~(w954 | w4105);
assign w996 = v357;
assign w997 = (w955 & ~w4139) | (w955 & w2961) | (~w4139 & w2961);
assign w998 = (~w2076 & w3745) | (~w2076 & w3407) | (w3745 & w3407);
assign v358 = ~(w250 | w610);
assign w999 = v358;
assign v359 = ~(w3312 | w422);
assign w1000 = v359;
assign w1001 = w1036 & w704;
assign w1002 = w2087 & w1233;
assign v360 = ~(w954 | w91);
assign w1003 = v360;
assign w1004 = ~w135 & w1161;
assign w1005 = w3547 & w3118;
assign w1006 = ~w3501 & w3463;
assign w1007 = w226 & ~w860;
assign w1008 = w1515 & w257;
assign v361 = ~(w2426 | w1952);
assign w1009 = v361;
assign v362 = ~(w2936 | w3687);
assign w1010 = v362;
assign v363 = ~(w3312 | w149);
assign w1011 = v363;
assign v364 = ~(w2123 | w954);
assign w1012 = v364;
assign w1013 = w118 & pi064;
assign v365 = ~(w2300 | w2767);
assign w1014 = v365;
assign v366 = ~(w3080 | w2485);
assign w1015 = v366;
assign w1016 = w705 & w205;
assign w1017 = (w2993 & ~w1689) | (w2993 & w895) | (~w1689 & w895);
assign w1018 = ~w1469 & w1249;
assign w1019 = w3630 & ~w2467;
assign v367 = ~(w1970 | w794);
assign w1020 = v367;
assign v368 = ~(w2186 | w1321);
assign w1021 = v368;
assign w1022 = w1219 & w426;
assign w1023 = w3780 & w1856;
assign w1024 = ~w1971 & w3674;
assign v369 = ~(w2799 | w2955);
assign w1025 = v369;
assign v370 = ~(w150 | w1006);
assign w1026 = v370;
assign v371 = ~(w4159 | w1782);
assign w1027 = v371;
assign w1028 = w2936 & w718;
assign w1029 = pi119 & w570;
assign w1030 = pi162 & w1570;
assign v372 = ~(w1148 | w501);
assign w1031 = v372;
assign w1032 = ~pi366 & pi199;
assign w1033 = w3838 & w3350;
assign w1034 = ~w1469 & w838;
assign w1035 = ~w346 & w1002;
assign v373 = ~(w996 | w2538);
assign w1036 = v373;
assign w1037 = w158 & w1654;
assign w1038 = w2817 & w462;
assign w1039 = w1105 & ~w597;
assign w1040 = ~w3659 & w281;
assign w1041 = ~w1119 & w3879;
assign w1042 = w3817 & w2690;
assign w1043 = ~pi366 & pi224;
assign v374 = ~(w1354 | w258);
assign w1044 = v374;
assign w1045 = w656 & ~w3848;
assign v375 = ~(w2228 | w2556);
assign w1046 = v375;
assign v376 = ~(w954 | w357);
assign w1047 = v376;
assign w1048 = w3094 & w1632;
assign w1049 = ~w2746 & w2361;
assign w1050 = w1457 & w3283;
assign w1051 = w3427 & ~w1469;
assign w1052 = w118 & pi023;
assign w1053 = w3730 & w1654;
assign w1054 = w2747 & w2466;
assign v377 = ~(w622 | w520);
assign w1055 = v377;
assign w1056 = w2717 & ~w2085;
assign w1057 = w2387 & w808;
assign w1058 = (pi015 & ~w1654) | (pi015 & w1935) | (~w1654 & w1935);
assign w1059 = (w1469 & ~w1099) | (w1469 & w3958) | (~w1099 & w3958);
assign w1060 = pi328 & ~pi366;
assign w1061 = (~w2484 & w138) | (~w2484 & w1891) | (w138 & w1891);
assign w1062 = (w128 & w1318) | (w128 & w4156) | (w1318 & w4156);
assign w1063 = w705 & w1786;
assign w1064 = (w492 & w872) | (w492 & w1033) | (w872 & w1033);
assign v378 = ~(w487 | w2180);
assign w1065 = v378;
assign w1066 = w2411 & ~w555;
assign v379 = ~(w214 | w3326);
assign w1067 = v379;
assign v380 = ~(w3259 | w3943);
assign w1068 = v380;
assign w1069 = w1249 & ~w3489;
assign v381 = ~(w2314 | w1224);
assign w1070 = v381;
assign w1071 = ~w413 & w773;
assign w1072 = w2717 & ~w1604;
assign v382 = ~(w510 | w3817);
assign w1073 = v382;
assign v383 = ~(w2864 | w3470);
assign w1074 = v383;
assign w1075 = w1469 & w838;
assign w1076 = ~w539 & w2000;
assign v384 = ~(w3312 | w657);
assign w1077 = v384;
assign v385 = ~(w2475 | w357);
assign w1078 = v385;
assign v386 = ~(w456 | w1484);
assign w1079 = v386;
assign w1080 = ~w3686 & w3358;
assign w1081 = w3531 & ~w2330;
assign v387 = ~(w434 | w2916);
assign w1082 = v387;
assign v388 = ~(w2695 | w3889);
assign w1083 = v388;
assign w1084 = w838 & ~w2662;
assign w1085 = (~w2324 & ~w1227) | (~w2324 & w2198) | (~w1227 & w2198);
assign w1086 = w786 & w2520;
assign v389 = ~(w179 | w4038);
assign w1087 = v389;
assign v390 = ~(w2048 | w931);
assign w1088 = v390;
assign v391 = ~(w2879 | w2734);
assign w1089 = v391;
assign w1090 = pi167 & ~pi364;
assign v392 = ~(w3312 | w923);
assign w1091 = v392;
assign w1092 = (~w2626 & w2570) | (~w2626 & w715) | (w2570 & w715);
assign v393 = ~(w1534 | w3507);
assign w1093 = v393;
assign w1094 = ~w2874 & w656;
assign w1095 = ~w1629 & w1884;
assign w1096 = w3094 & w1641;
assign v394 = ~(w4120 | w3932);
assign w1097 = v394;
assign v395 = ~(w3878 | w3414);
assign w1098 = v395;
assign v396 = ~(w2346 | w2709);
assign w1099 = v396;
assign v397 = ~(w2941 | w2640);
assign w1100 = v397;
assign w1101 = w1198 & w4183;
assign v398 = ~(w2660 | w2767);
assign w1102 = v398;
assign v399 = ~(w539 | w361);
assign w1103 = v399;
assign w1104 = ~w3945 & w2299;
assign w1105 = (w2487 & ~w951) | (w2487 & w3733) | (~w951 & w3733);
assign w1106 = pi290 & w2362;
assign w1107 = ~w2417 & w2763;
assign w1108 = ~w2268 & w991;
assign v400 = ~(w1673 | w3312);
assign w1109 = v400;
assign w1110 = ~pi366 & pi232;
assign w1111 = pi319 & ~pi366;
assign v401 = ~(w1421 | w711);
assign w1112 = v401;
assign w1113 = w2519 & w3085;
assign v402 = ~(w2893 | w187);
assign w1114 = v402;
assign v403 = ~(w2799 | w3317);
assign w1115 = v403;
assign w1116 = w3732 & w309;
assign v404 = ~(w4087 | w3878);
assign w1117 = v404;
assign w1118 = w135 & ~w2044;
assign w1119 = ~w1390 & w3398;
assign v405 = ~(w1442 | w696);
assign w1120 = v405;
assign v406 = ~(w3908 | w186);
assign w1121 = v406;
assign w1122 = w2471 & ~w1469;
assign v407 = ~(w3806 | w2130);
assign w1123 = v407;
assign w1124 = ~w2846 & w1552;
assign v408 = ~(w1205 | w2184);
assign w1125 = v408;
assign w1126 = w1829 & ~w521;
assign v409 = ~(w827 | w2469);
assign w1127 = v409;
assign w1128 = w2084 & w2786;
assign w1129 = w705 & w4058;
assign w1130 = w2870 & w1138;
assign w1131 = w2463 & w1520;
assign v410 = ~(w2324 | w4047);
assign w1132 = v410;
assign w1133 = pi108 & w353;
assign w1134 = w672 & ~w3193;
assign v411 = ~(w0 | w1353);
assign w1135 = v411;
assign w1136 = (w1333 & ~w4109) | (w1333 & w2264) | (~w4109 & w2264);
assign v412 = ~(w2137 | w4101);
assign w1137 = v412;
assign v413 = ~(w3693 | w3353);
assign w1138 = v413;
assign v414 = ~(w1821 | w2292);
assign w1139 = v414;
assign w1140 = ~w78 & w1356;
assign w1141 = w382 & w3099;
assign w1142 = w4049 & ~w354;
assign v415 = ~(w1373 | w3448);
assign w1143 = v415;
assign v416 = ~(w2123 | w3878);
assign w1144 = v416;
assign v417 = ~(w3594 | w2806);
assign w1145 = v417;
assign v418 = ~(w2799 | w1104);
assign w1146 = v418;
assign w1147 = w656 & ~w4087;
assign v419 = ~(w1140 | w1970);
assign w1148 = v419;
assign w1149 = w1888 & w1869;
assign w1150 = (pi091 & ~w1654) | (pi091 & w3177) | (~w1654 & w3177);
assign w1151 = pi283 & w2362;
assign v420 = ~(w3515 | w2167);
assign w1152 = v420;
assign v421 = ~(w1197 | w515);
assign w1153 = v421;
assign w1154 = ~w3690 & w961;
assign v422 = ~(w1970 | w3168);
assign w1155 = v422;
assign w1156 = w578 & w1818;
assign w1157 = w3588 & ~w1139;
assign v423 = ~(w749 | w3151);
assign w1158 = v423;
assign w1159 = w2373 & ~w1774;
assign v424 = ~(w1661 | w3722);
assign w1160 = v424;
assign w1161 = w2976 & w2489;
assign w1162 = ~w3518 & w3016;
assign v425 = ~(w2689 | w3629);
assign w1163 = v425;
assign w1164 = ~w962 & w1896;
assign w1165 = w221 & w710;
assign w1166 = w3527 & w2142;
assign w1167 = w1320 & w3468;
assign v426 = ~(w3878 | w1899);
assign w1168 = v426;
assign v427 = ~(w3878 | w3385);
assign w1169 = v427;
assign w1170 = w865 & ~w3068;
assign w1171 = w656 & ~w1104;
assign v428 = ~(w734 | w2482);
assign w1172 = v428;
assign v429 = ~(w425 | w834);
assign w1173 = v429;
assign w1174 = w3094 & w3458;
assign v430 = ~(w3974 | w1437);
assign w1175 = v430;
assign w1176 = w656 & ~w3168;
assign w1177 = (w1539 & w2030) | (w1539 & w383) | (w2030 & w383);
assign v431 = ~(w444 | w2716);
assign w1178 = v431;
assign v432 = ~(w2516 | w4154);
assign w1179 = v432;
assign w1180 = w1830 & ~w1592;
assign w1181 = w118 & pi065;
assign w1182 = w930 & w3547;
assign w1183 = (w1654 & w2339) | (w1654 & w297) | (w2339 & w297);
assign w1184 = w2082 & w2126;
assign w1185 = w3394 & w1469;
assign v433 = ~(w2162 | w3357);
assign w1186 = v433;
assign v434 = ~(w3484 | w4085);
assign w1187 = v434;
assign v435 = ~(w3090 | w2796);
assign w1188 = v435;
assign w1189 = w1834 & ~w3315;
assign w1190 = w1727 & w2670;
assign w1191 = w4158 & ~w3331;
assign w1192 = ~w1184 & w3986;
assign w1193 = w118 & pi117;
assign v436 = ~(w4038 | w2085);
assign w1194 = v436;
assign w1195 = (w1075 & ~w2369) | (w1075 & w3618) | (~w2369 & w3618);
assign v437 = ~(w1799 | w3390);
assign w1196 = v437;
assign v438 = ~(w2799 | w3131);
assign w1197 = v438;
assign w1198 = w1165 & w1723;
assign w1199 = w3062 & w3118;
assign v439 = ~(w2175 | w923);
assign w1200 = v439;
assign v440 = ~(w991 | w1441);
assign w1201 = v440;
assign w1202 = (w2179 & ~w2572) | (w2179 & w922) | (~w2572 & w922);
assign w1203 = pi314 & ~pi366;
assign w1204 = (w1654 & w3818) | (w1654 & w330) | (w3818 & w330);
assign v441 = ~(w954 | w4087);
assign w1205 = v441;
assign w1206 = ~pi366 & pi194;
assign w1207 = w3180 & ~w658;
assign w1208 = (~w1469 & ~w1121) | (~w1469 & w2789) | (~w1121 & w2789);
assign w1209 = w3549 & w3846;
assign v442 = ~(w1661 | w3977);
assign w1210 = v442;
assign w1211 = (~w1469 & ~w1838) | (~w1469 & w1122) | (~w1838 & w1122);
assign w1212 = w1570 & w477;
assign w1213 = (w1654 & w2725) | (w1654 & w1053) | (w2725 & w1053);
assign v443 = ~(w1717 | w3400);
assign w1214 = v443;
assign w1215 = w3967 & w1240;
assign w1216 = pi135 & ~pi364;
assign v444 = ~(w1406 | w941);
assign w1217 = v444;
assign w1218 = ~w831 & w2631;
assign w1219 = w860 & ~w3061;
assign v445 = ~(w3878 | w3105);
assign w1220 = v445;
assign v446 = ~(w3878 | w2085);
assign w1221 = v446;
assign w1222 = w3179 & ~w2131;
assign w1223 = w425 & ~w2484;
assign v447 = ~(w2175 | w4105);
assign w1224 = v447;
assign v448 = ~(w3160 | w357);
assign w1225 = v448;
assign v449 = ~(w3312 | w3848);
assign w1226 = v449;
assign v450 = ~(w3294 | w3495);
assign w1227 = v450;
assign w1228 = w2370 & w1654;
assign w1229 = w2244 & w1853;
assign w1230 = w3372 & w384;
assign w1231 = ~w1139 & w162;
assign w1232 = w2039 & w3699;
assign v451 = ~(w1747 | w1945);
assign w1233 = v451;
assign w1234 = w118 & pi096;
assign w1235 = pi352 & ~pi366;
assign w1236 = ~w2896 & w1229;
assign w1237 = ~w439 & w3313;
assign w1238 = w118 & pi116;
assign w1239 = w656 & ~w3462;
assign v452 = ~(w810 | w206);
assign w1240 = v452;
assign v453 = ~(w3507 | w2367);
assign w1241 = v453;
assign w1242 = w3451 & w107;
assign v454 = ~(w294 | w559);
assign w1243 = v454;
assign w1244 = w2325 & ~w3887;
assign w1245 = w860 & ~w183;
assign w1246 = ~w3094 & w3389;
assign w1247 = w2022 & ~w1139;
assign w1248 = (w1080 & ~w3656) | (w1080 & w2276) | (~w3656 & w2276);
assign w1249 = w2357 & w1273;
assign w1250 = w2893 & w4047;
assign v455 = ~(w3929 | w1754);
assign w1251 = v455;
assign w1252 = pi085 & w570;
assign v456 = ~(w2625 | w2040);
assign w1253 = v456;
assign v457 = ~(w1622 | w2146);
assign w1254 = v457;
assign v458 = ~(w4174 | w1756);
assign w1255 = v458;
assign w1256 = pi181 & ~pi364;
assign w1257 = w3222 & w290;
assign w1258 = pi156 & w1570;
assign v459 = ~(w3175 | w1418);
assign w1259 = v459;
assign v460 = ~(w2754 | w3266);
assign w1260 = v460;
assign w1261 = w688 & w385;
assign w1262 = (w3422 & ~w47) | (w3422 & w2798) | (~w47 & w2798);
assign v461 = ~(w954 | w3263);
assign w1263 = v461;
assign w1264 = ~w1389 & w965;
assign w1265 = w1127 & w62;
assign v462 = ~(w790 | w654);
assign w1266 = v462;
assign v463 = ~(w3312 | w3964);
assign w1267 = v463;
assign v464 = ~(w1349 | w2171);
assign w1268 = v464;
assign w1269 = (w3226 & w4083) | (w3226 & w621) | (w4083 & w621);
assign w1270 = ~w3001 & w2166;
assign w1271 = pi004 & w570;
assign w1272 = w138 & w3825;
assign w1273 = pi364 & ~pi365;
assign w1274 = w3159 & ~w361;
assign v465 = ~(w3160 | w3343);
assign w1275 = v465;
assign v466 = ~(w2905 | w487);
assign w1276 = v466;
assign w1277 = w3813 & w2554;
assign v467 = ~(w370 | w985);
assign w1278 = v467;
assign w1279 = ~pi366 & pi198;
assign w1280 = w118 & pi126;
assign v468 = ~(w2475 | w91);
assign w1281 = v468;
assign v469 = ~(w4038 | w657);
assign w1282 = v469;
assign w1283 = (w2631 & ~w578) | (w2631 & w1218) | (~w578 & w1218);
assign v470 = ~(w1754 | w3977);
assign w1284 = v470;
assign v471 = ~(w797 | w1147);
assign w1285 = v471;
assign v472 = ~(w1754 | w557);
assign w1286 = v472;
assign w1287 = ~w1798 & w1784;
assign w1288 = w2626 & ~w1405;
assign v473 = ~(w3628 | w2460);
assign w1289 = v473;
assign v474 = ~(w3878 | w3848);
assign w1290 = v474;
assign v475 = ~(w1157 | w1556);
assign w1291 = v475;
assign w1292 = ~w3094 & w2049;
assign v476 = ~(w1089 | w294);
assign w1293 = v476;
assign w1294 = pi152 & w1570;
assign v477 = ~(w2373 | w3179);
assign w1295 = v477;
assign w1296 = (w1249 & w1603) | (w1249 & w2190) | (w1603 & w2190);
assign w1297 = pi154 & w1570;
assign w1298 = w2004 & ~w964;
assign w1299 = (w1566 & ~w2860) | (w1566 & w3503) | (~w2860 & w3503);
assign v478 = ~(w954 | w923);
assign w1300 = v478;
assign v479 = ~(w4049 | w3084);
assign w1301 = v479;
assign w1302 = w1022 & w2750;
assign v480 = ~(w3779 | w33);
assign w1303 = v480;
assign w1304 = w649 & w142;
assign w1305 = w2022 & w4010;
assign w1306 = w3300 & w1702;
assign v481 = ~(w1579 | w162);
assign w1307 = v481;
assign w1308 = w2813 & w1625;
assign w1309 = w2578 & ~w1469;
assign w1310 = w2058 & ~w3667;
assign w1311 = pi333 & ~pi366;
assign v482 = ~(w1661 | w557);
assign w1312 = v482;
assign w1313 = pi160 & w1570;
assign w1314 = w2244 & ~w4001;
assign w1315 = w1089 & w565;
assign w1316 = (w1653 & ~w1605) | (w1653 & w2308) | (~w1605 & w2308);
assign w1317 = ~w3544 & w1259;
assign v483 = ~(w2651 | w635);
assign w1318 = v483;
assign w1319 = w4074 & ~w4065;
assign w1320 = w554 & w1802;
assign v484 = ~(w3160 | w1140);
assign w1321 = v484;
assign w1322 = w1137 & w3755;
assign w1323 = w3094 & w3336;
assign w1324 = (w1469 & ~w1660) | (w1469 & w2712) | (~w1660 & w2712);
assign v485 = ~(w1977 | w2647);
assign w1325 = v485;
assign w1326 = w3183 & ~w3422;
assign w1327 = ~pi366 & pi221;
assign v486 = ~(w1865 | w4121);
assign w1328 = v486;
assign v487 = ~(w3312 | w1633);
assign w1329 = v487;
assign v488 = ~(w1913 | w3638);
assign w1330 = v488;
assign w1331 = ~w2484 & w442;
assign w1332 = ~w2461 & w2428;
assign w1333 = ~w4135 & w1850;
assign v489 = ~(w547 | w3043);
assign w1334 = v489;
assign w1335 = w118 & pi027;
assign v490 = ~(w3261 | w2510);
assign w1336 = v490;
assign v491 = ~(w2802 | w3355);
assign w1337 = v491;
assign w1338 = w3735 & w3459;
assign w1339 = w705 & w3937;
assign w1340 = pi121 & w353;
assign v492 = ~(w3312 | w1592);
assign w1341 = v492;
assign v493 = ~(w2941 | w2300);
assign w1342 = v493;
assign w1343 = w539 & w361;
assign w1344 = (~w2484 & w121) | (~w2484 & w3903) | (w121 & w3903);
assign w1345 = w3694 & ~w834;
assign w1346 = ~w2942 & w2464;
assign w1347 = pi186 & w1570;
assign w1348 = w141 & w565;
assign w1349 = w3094 & w506;
assign w1350 = w4119 & w1469;
assign w1351 = (w1654 & w1540) | (w1654 & w2404) | (w1540 & w2404);
assign v494 = ~(w4038 | w3343);
assign w1352 = v494;
assign w1353 = w1382 & w864;
assign w1354 = w838 & ~w2881;
assign v495 = ~(w3204 | w1855);
assign w1355 = v495;
assign v496 = ~(w3872 | w3652);
assign w1356 = v496;
assign w1357 = w1376 & w4075;
assign v497 = ~(w2509 | w1366);
assign w1358 = v497;
assign v498 = ~(w4137 | w46);
assign w1359 = v498;
assign v499 = ~(w2525 | w35);
assign w1360 = v499;
assign w1361 = (w838 & w2168) | (w838 & w1460) | (w2168 & w1460);
assign w1362 = w388 & w1469;
assign w1363 = ~w1469 & w4015;
assign w1364 = w1637 & ~w2933;
assign w1365 = w1830 & ~w1604;
assign w1366 = (pi117 & ~w1654) | (pi117 & w1193) | (~w1654 & w1193);
assign w1367 = w16 & w2069;
assign v500 = ~(w2475 | w448);
assign w1368 = v500;
assign v501 = ~(w3153 | w960);
assign w1369 = v501;
assign w1370 = w378 & ~w1501;
assign v502 = ~(w2132 | w468);
assign w1371 = v502;
assign v503 = ~(w3878 | w3343);
assign w1372 = v503;
assign w1373 = ~w807 & w3395;
assign v504 = ~(w3905 | w3848);
assign w1374 = v504;
assign w1375 = w735 & w1654;
assign v505 = ~(w1180 | w2909);
assign w1376 = v505;
assign w1377 = (w1469 & ~w2434) | (w1469 & w1946) | (~w2434 & w1946);
assign v506 = ~(w1673 | w1970);
assign w1378 = v506;
assign w1379 = w4015 & ~w2821;
assign v507 = ~(w4159 | w1667);
assign w1380 = v507;
assign v508 = ~(w2019 | w4050);
assign w1381 = v508;
assign w1382 = w3738 & ~w1778;
assign v509 = ~(w708 | w83);
assign w1383 = v509;
assign w1384 = (pi120 & ~w1654) | (pi120 & w1488) | (~w1654 & w1488);
assign w1385 = w1088 & w1835;
assign v510 = ~(w1996 | w3260);
assign w1386 = v510;
assign w1387 = ~w226 & w860;
assign v511 = ~(w1662 | w49);
assign w1388 = v511;
assign v512 = ~(w2877 | w2479);
assign w1389 = v512;
assign w1390 = (~w1458 & w1291) | (~w1458 & w1687) | (w1291 & w1687);
assign w1391 = ~w2004 & w2315;
assign v513 = ~(w2799 | w3462);
assign w1392 = v513;
assign v514 = ~(w2423 | w901);
assign w1393 = v514;
assign v515 = ~(w2226 | w3404);
assign w1394 = v515;
assign w1395 = pi165 & ~pi364;
assign w1396 = w3094 & w3267;
assign w1397 = w1285 & w914;
assign w1398 = w3378 & w1244;
assign w1399 = w1107 & ~w3323;
assign w1400 = ~w4114 & w152;
assign w1401 = w433 & ~w2807;
assign w1402 = ~w92 & w2133;
assign v516 = ~(w56 | w2461);
assign w1403 = v516;
assign w1404 = (w354 & w2592) | (w354 & w2622) | (w2592 & w2622);
assign v517 = ~(w2074 | w661);
assign w1405 = v517;
assign w1406 = w3094 & w3136;
assign w1407 = w705 & w2744;
assign v518 = ~(w2640 | w2767);
assign w1408 = v518;
assign v519 = ~(w4159 | w657);
assign w1409 = v519;
assign v520 = ~(w465 | w1655);
assign w1410 = v520;
assign v521 = ~(w2227 | w306);
assign w1411 = v521;
assign w1412 = w4049 & w1387;
assign v522 = ~(w2874 | w3312);
assign w1413 = v522;
assign w1414 = w2993 & w729;
assign v523 = ~(w2936 | w217);
assign w1415 = v523;
assign v524 = ~(w2175 | w657);
assign w1416 = v524;
assign v525 = ~(w2377 | w332);
assign w1417 = v525;
assign w1418 = w705 & w4086;
assign v526 = ~(w319 | w776);
assign w1419 = v526;
assign v527 = ~(w2206 | w3643);
assign w1420 = v527;
assign v528 = ~(w954 | w422);
assign w1421 = v528;
assign w1422 = pi252 & w2362;
assign w1423 = pi025 & w570;
assign v529 = ~(w954 | w542);
assign w1424 = v529;
assign w1425 = (w1469 & ~w1838) | (w1469 & w191) | (~w1838 & w191);
assign w1426 = w3094 & w761;
assign w1427 = w1486 & w2094;
assign v530 = ~(w4038 | w3943);
assign w1428 = v530;
assign w1429 = w354 & w3061;
assign w1430 = w2283 & ~w1469;
assign w1431 = pi178 & w1570;
assign v531 = ~(w1089 | w1864);
assign w1432 = v531;
assign w1433 = w2717 & ~w1782;
assign w1434 = w3994 & ~w1630;
assign w1435 = pi292 & w2362;
assign w1436 = ~w853 & w126;
assign w1437 = ~w3352 & w2711;
assign w1438 = ~w1985 & w893;
assign w1439 = w909 & w1654;
assign w1440 = w4092 & w2422;
assign v532 = ~(w3654 | w483);
assign w1441 = v532;
assign v533 = ~(w954 | w398);
assign w1442 = v533;
assign w1443 = ~w3094 & w3642;
assign w1444 = ~w2371 & w2718;
assign v534 = ~(w1598 | w1251);
assign w1445 = v534;
assign w1446 = w2022 & ~w2050;
assign w1447 = ~w2046 & w435;
assign v535 = ~(w3894 | w2864);
assign w1448 = v535;
assign w1449 = pi251 & w2362;
assign v536 = ~(w1661 | w3263);
assign w1450 = v536;
assign v537 = ~(w2898 | w3294);
assign w1451 = v537;
assign w1452 = w778 & ~w784;
assign w1453 = w734 & w2967;
assign v538 = ~(w1979 | w1949);
assign w1454 = v538;
assign w1455 = w433 & ~w2959;
assign v539 = ~(w3761 | w1109);
assign w1456 = v539;
assign w1457 = w1650 & w3376;
assign w1458 = w4010 & ~w1139;
assign w1459 = w2397 & ~w2;
assign w1460 = w1878 & w838;
assign w1461 = w2717 & ~w422;
assign w1462 = ~w2504 & w1318;
assign w1463 = (~w1469 & ~w1950) | (~w1469 & w2809) | (~w1950 & w2809);
assign w1464 = w1469 & ~w3630;
assign v540 = ~(w1883 | w2487);
assign w1465 = v540;
assign w1466 = pi111 & w570;
assign v541 = ~(w800 | w2058);
assign w1467 = v541;
assign w1468 = pi301 & w2362;
assign v542 = ~(w2263 | w4043);
assign w1469 = v542;
assign v543 = ~(w2315 | w1089);
assign w1470 = v543;
assign v544 = ~(w2424 | w1295);
assign w1471 = v544;
assign w1472 = pi036 & w570;
assign v545 = ~(w906 | w3997);
assign w1473 = v545;
assign w1474 = w2568 & w4098;
assign v546 = ~(w791 | w2900);
assign w1475 = v546;
assign v547 = ~(w3810 | w4008);
assign w1476 = v547;
assign w1477 = pi159 & ~pi364;
assign w1478 = ~w778 & w784;
assign w1479 = w1387 & w2477;
assign v548 = ~(w2799 | w3722);
assign w1480 = v548;
assign v549 = ~(w2387 | w2574);
assign w1481 = v549;
assign v550 = ~(w1661 | w1533);
assign w1482 = v550;
assign w1483 = w1249 & ~w2990;
assign w1484 = ~w1699 & w449;
assign w1485 = w1776 & w1469;
assign w1486 = ~w3094 & w1676;
assign v551 = ~(w3920 | w3010);
assign w1487 = v551;
assign w1488 = w118 & pi120;
assign v552 = ~(w3169 | w1312);
assign w1489 = v552;
assign v553 = ~(w3050 | w816);
assign w1490 = v553;
assign w1491 = (~w3323 & w3285) | (~w3323 & w1399) | (w3285 & w1399);
assign v554 = ~(w2373 | w3216);
assign w1492 = v554;
assign w1493 = ~w3031 & w1270;
assign v555 = ~(w894 | w358);
assign w1494 = v555;
assign v556 = ~(w3878 | w557);
assign w1495 = v556;
assign v557 = ~(w954 | w3722);
assign w1496 = v557;
assign w1497 = pi342 & ~pi366;
assign v558 = ~(w3307 | w1718);
assign w1498 = v558;
assign w1499 = w2373 & w3216;
assign w1500 = w950 & ~w402;
assign v559 = ~(w1059 | w1211);
assign w1501 = v559;
assign w1502 = w2717 & ~w923;
assign v560 = ~(w954 | w3385);
assign w1503 = v560;
assign w1504 = w354 & ~w874;
assign v561 = ~(w3259 | w1782);
assign w1505 = v561;
assign w1506 = w1469 & w378;
assign w1507 = w1319 & w56;
assign w1508 = ~w1759 & w647;
assign v562 = ~(w4038 | w3414);
assign w1509 = v562;
assign w1510 = ~w3094 & w2035;
assign w1511 = (pi065 & ~w1654) | (pi065 & w1181) | (~w1654 & w1181);
assign v563 = ~(w995 | w3597);
assign w1512 = v563;
assign v564 = ~(w3297 | w3143);
assign w1513 = v564;
assign w1514 = w4094 & w589;
assign v565 = ~(w2888 | w593);
assign w1515 = v565;
assign w1516 = (w1469 & ~w4127) | (w1469 & w3681) | (~w4127 & w3681);
assign v566 = ~(w324 | w4015);
assign w1517 = v566;
assign w1518 = w73 & ~w1469;
assign w1519 = w2690 & ~w544;
assign w1520 = w2141 & w2781;
assign w1521 = pi018 & w570;
assign w1522 = (~w3226 & w3229) | (~w3226 & w636) | (w3229 & w636);
assign v567 = ~(w1754 | w1104);
assign w1523 = v567;
assign v568 = ~(w301 | w3247);
assign w1524 = v568;
assign w1525 = ~w964 & w961;
assign w1526 = ~w1318 & w361;
assign v569 = ~(w1768 | w2791);
assign w1527 = v569;
assign w1528 = (~w1469 & ~w2299) | (~w1469 & w3564) | (~w2299 & w3564);
assign w1529 = ~w2030 & w998;
assign v570 = ~(w4038 | w1667);
assign w1530 = v570;
assign w1531 = w3347 & w875;
assign w1532 = w3094 & w3580;
assign w1533 = ~w1976 & w2678;
assign w1534 = w2058 & w2213;
assign w1535 = pi284 & w2362;
assign w1536 = w4119 & ~w1469;
assign v571 = ~(w1970 | w1633);
assign w1537 = v571;
assign w1538 = (w1249 & w3696) | (w1249 & w4132) | (w3696 & w4132);
assign w1539 = ~w2576 & w3708;
assign w1540 = pi053 & w570;
assign v572 = ~(w1810 | w2660);
assign w1541 = v572;
assign v573 = ~(w3426 | w3312);
assign w1542 = v573;
assign v574 = ~(w103 | w1739);
assign w1543 = v574;
assign w1544 = pi100 & w570;
assign w1545 = pi276 & w2362;
assign v575 = ~(w2799 | w4105);
assign w1546 = v575;
assign w1547 = ~w3628 & w1458;
assign w1548 = w979 & w2014;
assign w1549 = ~w846 & w486;
assign w1550 = (w3191 & w1022) | (w3191 & w229) | (w1022 & w229);
assign w1551 = pi112 & w353;
assign w1552 = ~w1400 & w2232;
assign v576 = ~(w687 | w2072);
assign w1553 = v576;
assign w1554 = w292 & w39;
assign w1555 = ~w3126 & w2820;
assign w1556 = w2774 & ~w1247;
assign w1557 = w1586 & w2366;
assign v577 = ~(w3160 | w3964);
assign w1558 = v577;
assign w1559 = w656 & ~w3426;
assign w1560 = (w3382 & ~w2433) | (w3382 & w1589) | (~w2433 & w1589);
assign v578 = ~(w728 | w701);
assign w1561 = v578;
assign v579 = ~(w324 | w1425);
assign w1562 = v579;
assign w1563 = w2717 & ~w1955;
assign w1564 = pi133 & ~pi364;
assign v580 = ~(w3832 | w457);
assign w1565 = v580;
assign v581 = ~(w3371 | w2758);
assign w1566 = v581;
assign w1567 = w3094 & w1111;
assign w1568 = (pi068 & ~w1654) | (pi068 & w2843) | (~w1654 & w2843);
assign v582 = ~(w3924 | w591);
assign w1569 = v582;
assign v583 = ~(pi366 | pi367);
assign w1570 = v583;
assign w1571 = ~w2836 & w677;
assign w1572 = ~w361 & w1318;
assign w1573 = w1735 & w2701;
assign w1574 = (pi017 & ~w1654) | (pi017 & w933) | (~w1654 & w933);
assign v584 = ~(w48 | w954);
assign w1575 = v584;
assign w1576 = w2178 & w676;
assign w1577 = ~w1140 & w1830;
assign w1578 = ~w3795 & w789;
assign w1579 = ~w4010 & w3628;
assign w1580 = w2234 & ~w1057;
assign v585 = ~(w712 | w1672);
assign w1581 = v585;
assign w1582 = (w2487 & ~w771) | (w2487 & w968) | (~w771 & w968);
assign w1583 = ~w1071 & w1237;
assign v586 = ~(w2968 | w1425);
assign w1584 = v586;
assign w1585 = pi289 & w2362;
assign v587 = ~(w3324 | w3709);
assign w1586 = v587;
assign w1587 = w433 & ~w1514;
assign w1588 = w569 & ~w1491;
assign w1589 = w3541 & w3382;
assign v588 = ~(w2175 | w3722);
assign w1590 = v588;
assign w1591 = w3341 & w3286;
assign w1592 = ~w4053 & w947;
assign v589 = ~(w935 | w1495);
assign w1593 = v589;
assign w1594 = w656 & ~w3977;
assign v590 = ~(w2123 | w2175);
assign w1595 = v590;
assign w1596 = w1619 & w640;
assign w1597 = ~w2817 & w3573;
assign v591 = ~(w3160 | w1607);
assign w1598 = v591;
assign v592 = ~(w1607 | w4038);
assign w1599 = v592;
assign w1600 = ~w3094 & w397;
assign w1601 = w2965 & ~w3380;
assign v593 = ~(w3160 | w1592);
assign w1602 = v593;
assign w1603 = (w1469 & ~w1217) | (w1469 & w1668) | (~w1217 & w1668);
assign w1604 = ~w1443 & w1121;
assign v594 = ~(w18 | w1483);
assign w1605 = v594;
assign w1606 = pi347 & ~pi366;
assign w1607 = ~w723 & w2251;
assign v595 = ~(w2475 | w557);
assign w1608 = v595;
assign v596 = ~(w2875 | w3713);
assign w1609 = v596;
assign v597 = ~(w4080 | w509);
assign w1610 = v597;
assign v598 = ~(w2123 | w4038);
assign w1611 = v598;
assign w1612 = w2717 & ~w542;
assign v599 = ~(w4038 | w357);
assign w1613 = v599;
assign w1614 = w1475 & w3133;
assign v600 = ~(w2945 | w288);
assign w1615 = v600;
assign v601 = ~(w2440 | w2976);
assign w1616 = v601;
assign w1617 = w913 & ~w3931;
assign v602 = ~(w1754 | w398);
assign w1618 = v602;
assign w1619 = ~w3586 & w2488;
assign v603 = ~(w3061 | w1629);
assign w1620 = v603;
assign w1621 = w626 & w1062;
assign w1622 = w656 & ~w448;
assign w1623 = w1548 & w1261;
assign w1624 = (~w3269 & w3412) | (~w3269 & w2493) | (w3412 & w2493);
assign v604 = ~(w86 | w3743);
assign w1625 = v604;
assign w1626 = w4074 & w138;
assign w1627 = w950 & ~w2946;
assign w1628 = w800 & w2936;
assign v605 = ~(w1007 | w1387);
assign w1629 = v605;
assign w1630 = (w2940 & w1827) | (w2940 & w4024) | (w1827 & w4024);
assign w1631 = (~w2173 & w1517) | (~w2173 & w1562) | (w1517 & w1562);
assign w1632 = pi348 & ~pi366;
assign w1633 = ~w3334 & w3319;
assign w1634 = pi185 & ~pi364;
assign w1635 = w4010 & w3628;
assign v606 = ~(w1882 | w1047);
assign w1636 = v606;
assign v607 = ~(w1204 | w2700);
assign w1637 = v607;
assign w1638 = ~w2726 & w3886;
assign v608 = ~(w1703 | w2093);
assign w1639 = v608;
assign w1640 = (w2993 & ~w571) | (w2993 & w1017) | (~w571 & w1017);
assign w1641 = pi310 & ~pi366;
assign v609 = ~(w3160 | w3105);
assign w1642 = v609;
assign w1643 = w560 & w765;
assign v610 = ~(w2432 | w2259);
assign w1644 = v610;
assign w1645 = ~w132 & w3051;
assign v611 = ~(w1661 | w3414);
assign w1646 = v611;
assign w1647 = w1471 & ~w46;
assign w1648 = w838 & ~w1408;
assign w1649 = ~w2682 & w2182;
assign v612 = ~(w902 | w2448);
assign w1650 = v612;
assign w1651 = w174 & w3975;
assign w1652 = w2213 & w1767;
assign v613 = ~(w2570 | w4073);
assign w1653 = v613;
assign w1654 = w2357 & w4000;
assign w1655 = w838 & ~w1692;
assign w1656 = (w1654 & w2483) | (w1654 & w3567) | (w2483 & w3567);
assign v614 = ~(w2175 | w3977);
assign w1657 = v614;
assign v615 = ~(w825 | w2727);
assign w1658 = v615;
assign v616 = ~(w3108 | w1868);
assign w1659 = v616;
assign v617 = ~(w812 | w3508);
assign w1660 = v617;
assign v618 = ~(w3898 | w3983);
assign w1661 = v618;
assign v619 = ~(w966 | w1845);
assign w1662 = v619;
assign v620 = ~(w2320 | w3851);
assign w1663 = v620;
assign v621 = ~(w315 | w4182);
assign w1664 = v621;
assign w1665 = (pi016 & ~w1654) | (pi016 & w726) | (~w1654 & w726);
assign w1666 = w929 & w1654;
assign w1667 = ~w805 & w1950;
assign w1668 = w2283 & w1469;
assign w1669 = w3094 & w4062;
assign w1670 = pi002 & w570;
assign w1671 = (w361 & ~w2070) | (w361 & w1812) | (~w2070 & w1812);
assign w1672 = pi250 & w2362;
assign w1673 = ~w1246 & w1660;
assign w1674 = w656 & ~w2955;
assign v622 = ~(w2616 | w821);
assign w1675 = v622;
assign w1676 = ~pi366 & pi200;
assign v623 = ~(w880 | w4034);
assign w1677 = v623;
assign w1678 = (~w1139 & w4094) | (~w1139 & w1247) | (w4094 & w1247);
assign w1679 = w838 & ~w1065;
assign w1680 = (w3706 & ~w2540) | (w3706 & w3442) | (~w2540 & w3442);
assign w1681 = w2443 & ~w2617;
assign v624 = ~(w3823 | w1059);
assign w1682 = v624;
assign w1683 = (w3085 & w365) | (w3085 & w2204) | (w365 & w2204);
assign w1684 = ~w2624 & w3002;
assign v625 = ~(w3277 | w954);
assign w1685 = v625;
assign v626 = ~(w4038 | w557);
assign w1686 = v626;
assign w1687 = w496 & ~w1458;
assign w1688 = w3199 & ~w2018;
assign v627 = ~(w438 | w1370);
assign w1689 = v627;
assign w1690 = w1292 & ~w1469;
assign v628 = ~(w3160 | w1444);
assign w1691 = v628;
assign v629 = ~(w1695 | w2088);
assign w1692 = v629;
assign v630 = ~(w2175 | w3263);
assign w1693 = v630;
assign w1694 = w656 & ~w3414;
assign w1695 = (~w1469 & ~w2369) | (~w1469 & w3058) | (~w2369 & w3058);
assign w1696 = w484 & ~w1469;
assign v631 = ~(w3946 | w3657);
assign w1697 = v631;
assign v632 = ~(w1351 | w1511);
assign w1698 = v632;
assign v633 = ~(w2810 | w1419);
assign w1699 = v633;
assign w1700 = ~w1857 & w98;
assign w1701 = w1837 & w801;
assign w1702 = w1985 & ~w893;
assign v634 = ~(w1104 | w3160);
assign w1703 = v634;
assign v635 = ~(w3178 | w3893);
assign w1704 = v635;
assign w1705 = w991 & ~w2280;
assign v636 = ~(w432 | w3146);
assign w1706 = v636;
assign w1707 = w128 & w2479;
assign w1708 = (w3898 & ~w947) | (w3898 & w3103) | (~w947 & w3103);
assign w1709 = ~w910 & w2208;
assign w1710 = (~w3669 & w298) | (~w3669 & w3646) | (w298 & w3646);
assign v637 = ~(w1661 | w1633);
assign w1711 = v637;
assign w1712 = w3061 & ~w874;
assign w1713 = w1600 & ~w1469;
assign w1714 = w1023 & w4031;
assign w1715 = ~w1196 & w2381;
assign w1716 = pi163 & w1570;
assign w1717 = w838 & ~w2636;
assign w1718 = (~w1469 & ~w2434) | (~w1469 & w2982) | (~w2434 & w2982);
assign w1719 = w3420 & ~w3256;
assign w1720 = ~w106 & w2397;
assign v638 = ~(w1661 | w2209);
assign w1721 = v638;
assign v639 = ~(w3531 | w217);
assign w1722 = v639;
assign w1723 = w235 & w1187;
assign w1724 = w2717 & ~w3414;
assign w1725 = (w893 & ~w3300) | (w893 & w1438) | (~w3300 & w1438);
assign w1726 = w3656 & w3218;
assign v640 = ~(w1069 | w530);
assign w1727 = v640;
assign w1728 = w1870 & ~w1469;
assign v641 = ~(w1754 | w3943);
assign w1729 = v641;
assign w1730 = (pi049 & ~w1654) | (pi049 & w2239) | (~w1654 & w2239);
assign w1731 = w118 & pi056;
assign v642 = ~(w954 | w1955);
assign w1732 = v642;
assign w1733 = (~w1469 & ~w1260) | (~w1469 & w3525) | (~w1260 & w3525);
assign w1734 = w3718 & w3393;
assign w1735 = w2185 & w2675;
assign v643 = ~(w3949 | w2638);
assign w1736 = v643;
assign v644 = ~(w2799 | w1592);
assign w1737 = v644;
assign v645 = ~(w3910 | w266);
assign w1738 = v645;
assign v646 = ~(w3905 | w542);
assign w1739 = v646;
assign v647 = ~(w3981 | w1915);
assign w1740 = v647;
assign v648 = ~(w3259 | w91);
assign w1741 = v648;
assign w1742 = w4109 & w2038;
assign v649 = ~(w2654 | w843);
assign w1743 = v649;
assign w1744 = pi103 & w570;
assign w1745 = w3467 & w1289;
assign w1746 = ~w1712 & w3384;
assign v650 = ~(w4159 | w3168);
assign w1747 = v650;
assign v651 = ~(w277 | w2457);
assign w1748 = v651;
assign w1749 = (w1469 & ~w2433) | (w1469 & w3397) | (~w2433 & w3397);
assign w1750 = ~w987 & w615;
assign w1751 = w378 & ~w3298;
assign v652 = ~(w3905 | w2955);
assign w1752 = v652;
assign w1753 = w2814 & w1654;
assign v653 = ~(w2094 | w4149);
assign w1754 = v653;
assign v654 = ~(w2475 | w2209);
assign w1755 = v654;
assign w1756 = w1830 & ~w3105;
assign v655 = ~(w4159 | w3426);
assign w1757 = v655;
assign v656 = ~(w1656 | w1843);
assign w1758 = v656;
assign w1759 = ~w719 & w3258;
assign w1760 = (pi063 & ~w1654) | (pi063 & w1943) | (~w1654 & w1943);
assign v657 = ~(w2683 | w793);
assign w1761 = v657;
assign w1762 = w435 & w3179;
assign w1763 = w118 & pi073;
assign w1764 = ~w3635 & w3496;
assign v658 = ~(w2475 | w1667);
assign w1765 = v658;
assign v659 = ~(w3948 | w3996);
assign w1766 = v659;
assign w1767 = (~w3180 & ~w2082) | (~w3180 & w3575) | (~w2082 & w3575);
assign v660 = ~(w954 | w1782);
assign w1768 = v660;
assign w1769 = w2207 & w3669;
assign w1770 = ~pi366 & pi215;
assign w1771 = ~w1469 & w2690;
assign w1772 = ~w3094 & w3815;
assign v661 = ~(w3823 | w2109);
assign w1773 = v661;
assign v662 = ~(w2046 | w435);
assign w1774 = v662;
assign w1775 = ~w2373 & w1774;
assign w1776 = ~w3094 & w2714;
assign v663 = ~(w276 | w1528);
assign w1777 = v663;
assign w1778 = w851 & w2428;
assign v664 = ~(w2484 | w851);
assign w1779 = v664;
assign w1780 = w2690 & ~w1773;
assign v665 = ~(w3224 | w1596);
assign w1781 = v665;
assign w1782 = ~w73 & w848;
assign w1783 = w876 & ~w2612;
assign w1784 = ~w1404 & w333;
assign v666 = ~(w1754 | w2874);
assign w1785 = v666;
assign w1786 = w1570 & w1216;
assign w1787 = (w718 & w2170) | (w718 & w2621) | (w2170 & w2621);
assign w1788 = (~w1469 & ~w3319) | (~w1469 & w993) | (~w3319 & w993);
assign v667 = ~(w700 | w2708);
assign w1789 = v667;
assign v668 = ~(w1380 | w2895);
assign w1790 = v668;
assign w1791 = w546 & w2594;
assign w1792 = w78 & ~w1469;
assign v669 = ~(w3855 | w3445);
assign w1793 = v669;
assign w1794 = w3094 & w3004;
assign v670 = ~(w1272 | w3645);
assign w1795 = v670;
assign w1796 = w4015 & ~w1014;
assign w1797 = w1510 & ~w1469;
assign w1798 = (~w3191 & ~w247) | (~w3191 & w2555) | (~w247 & w2555);
assign v671 = ~(w4121 | w3209);
assign w1799 = v671;
assign w1800 = ~w1616 & w1432;
assign v672 = ~(w2475 | w3722);
assign w1801 = v672;
assign v673 = ~(w585 | w2772);
assign w1802 = v673;
assign w1803 = w834 & w1223;
assign w1804 = w1839 & w423;
assign w1805 = ~pi366 & pi195;
assign w1806 = ~w356 & w4161;
assign w1807 = w2811 & w838;
assign w1808 = w1830 & ~w1444;
assign v674 = ~(w3259 | w657);
assign w1809 = v674;
assign w1810 = (w1469 & ~w1793) | (w1469 & w819) | (~w1793 & w819);
assign w1811 = w683 & w3013;
assign w1812 = w128 & w361;
assign v675 = ~(w1301 | w3191);
assign w1813 = v675;
assign w1814 = ~w841 & w586;
assign v676 = ~(w2738 | w4078);
assign w1815 = v676;
assign w1816 = ~w1637 & w2933;
assign w1817 = w3825 & w2224;
assign w1818 = w831 & ~w2631;
assign w1819 = (~w1469 & ~w1394) | (~w1469 & w1728) | (~w1394 & w1728);
assign w1820 = w1678 & w1057;
assign w1821 = w2462 & ~w72;
assign w1822 = (~w1653 & w1498) | (~w1653 & w1092) | (w1498 & w1092);
assign w1823 = w2387 & w1305;
assign w1824 = w2397 & ~w2034;
assign w1825 = w175 & w4137;
assign w1826 = ~w3262 & w1089;
assign w1827 = ~w3249 & w2853;
assign v677 = ~(w2175 | w3462);
assign w1828 = v677;
assign w1829 = ~w1278 & w1841;
assign v678 = ~(w2144 | w2211);
assign w1830 = v678;
assign v679 = ~(w2799 | w794);
assign w1831 = v679;
assign w1832 = (w3887 & ~w1531) | (w3887 & w2600) | (~w1531 & w2600);
assign w1833 = pi335 & ~pi366;
assign w1834 = w46 & ~w2057;
assign v680 = ~(w1409 | w392);
assign w1835 = v680;
assign v681 = ~(w3878 | w3858);
assign w1836 = v681;
assign w1837 = w124 & w2309;
assign v682 = ~(w699 | w976);
assign w1838 = v682;
assign w1839 = w1706 & w3330;
assign v683 = ~(w3905 | w3317);
assign w1840 = v683;
assign w1841 = w991 & ~w2898;
assign w1842 = ~w3199 & w1705;
assign w1843 = (pi074 & ~w1654) | (pi074 & w3185) | (~w1654 & w3185);
assign w1844 = w1830 & ~w1899;
assign w1845 = ~w1317 & w2859;
assign v684 = ~(w2908 | w3911);
assign w1846 = v684;
assign v685 = ~(w3747 | w3390);
assign w1847 = v685;
assign w1848 = ~w3900 & w2551;
assign w1849 = (~w1469 & ~w624) | (~w1469 & w2619) | (~w624 & w2619);
assign v686 = ~(w176 | w3210);
assign w1850 = v686;
assign v687 = ~(w1563 | w1413);
assign w1851 = v687;
assign v688 = ~(w1607 | w1661);
assign w1852 = v688;
assign v689 = ~(w418 | w885);
assign w1853 = v689;
assign v690 = ~(w1140 | w3878);
assign w1854 = v690;
assign w1855 = w3630 & ~w60;
assign w1856 = w667 & w1659;
assign w1857 = (~w3068 & ~w1241) | (~w3068 & w1170) | (~w1241 & w1170);
assign w1858 = (w3773 & ~w3189) | (w3773 & w625) | (~w3189 & w625);
assign w1859 = w184 & ~w1469;
assign w1860 = pi355 & ~pi366;
assign w1861 = w3741 & ~w1054;
assign w1862 = w118 & pi097;
assign w1863 = (pi045 & ~w1654) | (pi045 & w4117) | (~w1654 & w4117);
assign w1864 = ~w565 & w2440;
assign w1865 = w2070 & w1671;
assign v691 = ~(w308 | w3932);
assign w1866 = v691;
assign w1867 = ~w1201 & w1388;
assign w1868 = ~w1673 & w2717;
assign w1869 = w4115 & w2230;
assign w1870 = ~w3094 & w3202;
assign w1871 = (w3380 & ~w2241) | (w3380 & w691) | (~w2241 & w691);
assign w1872 = w3094 & w3876;
assign w1873 = ~w918 & w105;
assign w1874 = w3804 & w602;
assign v692 = ~(w3046 | w1239);
assign w1875 = v692;
assign w1876 = (w1654 & w3540) | (w1654 & w3517) | (w3540 & w3517);
assign w1877 = w650 & w3737;
assign w1878 = (~w1469 & ~w947) | (~w1469 & w3968) | (~w947 & w3968);
assign w1879 = w546 & w1892;
assign w1880 = ~w3094 & w3480;
assign w1881 = ~w3509 & w3673;
assign w1882 = w656 & ~w794;
assign w1883 = w4065 & w165;
assign v693 = ~(w3061 | w202);
assign w1884 = v693;
assign v694 = ~(w3874 | w2752);
assign w1885 = v694;
assign w1886 = (~w3180 & ~w2936) | (~w3180 & w2998) | (~w2936 & w2998);
assign v695 = ~(w1450 | w3849);
assign w1887 = v695;
assign w1888 = w3757 & w2222;
assign w1889 = w2573 & w3711;
assign w1890 = w1469 & w2397;
assign v696 = ~(w4065 | w2484);
assign w1891 = v696;
assign w1892 = w1469 & w2443;
assign w1893 = w2668 & ~w471;
assign w1894 = pi339 & ~pi366;
assign w1895 = w1469 & w950;
assign v697 = ~(w1174 | w3584);
assign w1896 = v697;
assign w1897 = (w123 & w2214) | (w123 & w3754) | (w2214 & w3754);
assign w1898 = w2540 & w2911;
assign w1899 = ~w1870 & w1394;
assign w1900 = w2968 & ~w410;
assign w1901 = ~w4128 & w324;
assign v698 = ~(w3240 | w1482);
assign w1902 = v698;
assign w1903 = w368 & w296;
assign v699 = ~(w4038 | w920);
assign w1904 = v699;
assign v700 = ~(w2175 | w1881);
assign w1905 = v700;
assign v701 = ~(w1754 | w1607);
assign w1906 = v701;
assign v702 = ~(w1754 | w3343);
assign w1907 = v702;
assign w1908 = w3248 & w1326;
assign v703 = ~(w762 | w3598);
assign w1909 = v703;
assign v704 = ~(w3087 | w2152);
assign w1910 = v704;
assign w1911 = ~w1697 & w2215;
assign v705 = ~(w2941 | w2536);
assign w1912 = v705;
assign w1913 = (w1654 & w2687) | (w1654 & w322) | (w2687 & w322);
assign w1914 = w2717 & ~w3263;
assign w1915 = w1830 & ~w398;
assign v706 = ~(w587 | w3197);
assign w1916 = v706;
assign w1917 = w455 & ~w1317;
assign w1918 = w4065 & ~w138;
assign w1919 = w2221 & w2160;
assign w1920 = ~w3094 & w1770;
assign v707 = ~(w2475 | w657);
assign w1921 = v707;
assign w1922 = w1605 & w1822;
assign w1923 = w2250 & ~w1333;
assign w1924 = ~w3923 & w2110;
assign w1925 = w735 & w3630;
assign v708 = ~(w2244 | w2044);
assign w1926 = v708;
assign v709 = ~(w954 | w2209);
assign w1927 = v709;
assign w1928 = w1199 & ~w3344;
assign v710 = ~(w877 | w1200);
assign w1929 = v710;
assign w1930 = w2397 & ~w1073;
assign w1931 = ~w3392 & w1186;
assign w1932 = w1445 & w3712;
assign v711 = ~(w226 | w3061);
assign w1933 = v711;
assign v712 = ~(w3152 | w2885);
assign w1934 = v712;
assign w1935 = w118 & pi015;
assign w1936 = (pi070 & ~w1654) | (pi070 & w2680) | (~w1654 & w2680);
assign v713 = ~(w2799 | w448);
assign w1937 = v713;
assign v714 = ~(w3037 | w1530);
assign w1938 = v714;
assign w1939 = w1005 & ~w3843;
assign w1940 = w118 & pi059;
assign w1941 = (~w2469 & w3518) | (~w2469 & w890) | (w3518 & w890);
assign w1942 = w921 & w2785;
assign w1943 = w118 & pi063;
assign v715 = ~(w2819 | w3356);
assign w1944 = v715;
assign v716 = ~(w1970 | w3317);
assign w1945 = v716;
assign w1946 = w2907 & w1469;
assign w1947 = w4020 & w1654;
assign w1948 = w656 & ~w657;
assign w1949 = (w965 & w1597) | (w965 & w1264) | (w1597 & w1264);
assign v717 = ~(w2386 | w2077);
assign w1950 = v717;
assign w1951 = w962 & w1469;
assign v718 = ~(w2799 | w542);
assign w1952 = v718;
assign v719 = ~(w179 | w1661);
assign w1953 = v719;
assign v720 = ~(w3167 | w2537);
assign w1954 = v720;
assign w1955 = ~w2247 & w3440;
assign w1956 = w128 & w2000;
assign w1957 = w3094 & w3777;
assign v721 = ~(w2646 | w3068);
assign w1958 = v721;
assign w1959 = w1969 & w3750;
assign v722 = ~(w2799 | w3385);
assign w1960 = v722;
assign v723 = ~(w1661 | w542);
assign w1961 = v723;
assign v724 = ~(w3719 | w3234);
assign w1962 = v724;
assign w1963 = (w1654 & w3477) | (w1654 & w1375) | (w3477 & w1375);
assign w1964 = ~w17 & w2203;
assign w1965 = (~w1469 & ~w709) | (~w1469 & w2694) | (~w709 & w2694);
assign v725 = ~(w1139 | w1983);
assign w1966 = v725;
assign w1967 = w656 & ~w1164;
assign w1968 = (w3669 & w2168) | (w3669 & w633) | (w2168 & w633);
assign v726 = ~(w3907 | w1078);
assign w1969 = v726;
assign v727 = ~(w1363 | w1506);
assign w1970 = v727;
assign w1971 = pi113 & w353;
assign w1972 = ~w694 & w1966;
assign w1973 = ~w2685 & w2017;
assign w1974 = w1772 & w1469;
assign v728 = ~(w3933 | w122);
assign w1975 = v728;
assign w1976 = ~w3094 & w1110;
assign v729 = ~(w3259 | w1899);
assign w1977 = v729;
assign w1978 = w1525 & w826;
assign w1979 = (w3127 & w1684) | (w3127 & w475) | (w1684 & w475);
assign w1980 = w2897 & w2534;
assign v730 = ~(w1665 | w2913);
assign w1981 = v730;
assign v731 = ~(w2475 | w3943);
assign w1982 = v731;
assign w1983 = (w433 & ~w3085) | (w433 & w3155) | (~w3085 & w3155);
assign v732 = ~(w3312 | w3317);
assign w1984 = v732;
assign w1985 = w3232 & w693;
assign w1986 = pi300 & w2362;
assign w1987 = ~w2528 & w1767;
assign v733 = ~(w1970 | w1667);
assign w1988 = v733;
assign v734 = ~(w1470 | w964);
assign w1989 = v734;
assign w1990 = w1474 & w2671;
assign v735 = ~(w1819 | w1059);
assign w1991 = v735;
assign w1992 = w391 & ~w3401;
assign w1993 = w3669 & ~w3605;
assign w1994 = w404 & w2391;
assign v736 = ~(w293 | w3055);
assign w1995 = v736;
assign w1996 = w32 & w101;
assign v737 = ~(w2475 | w542);
assign w1997 = v737;
assign w1998 = w2579 & w3074;
assign w1999 = (pi127 & ~w1654) | (pi127 & w493) | (~w1654 & w493);
assign v738 = ~(w2575 | w3276);
assign w2000 = v738;
assign w2001 = ~w3094 & w532;
assign w2002 = w1570 & w1256;
assign w2003 = pi129 & w1570;
assign w2004 = w3262 & ~w141;
assign v739 = ~(w524 | w948);
assign w2005 = v739;
assign w2006 = pi362 & ~pi363;
assign w2007 = w4015 & ~w721;
assign v740 = ~(w3277 | w1661);
assign w2008 = v740;
assign v741 = ~(w2667 | w487);
assign w2009 = v741;
assign v742 = ~(w2862 | w1751);
assign w2010 = v742;
assign w2011 = (w1062 & ~w3573) | (w1062 & w1621) | (~w3573 & w1621);
assign w2012 = w1570 & w2828;
assign v743 = ~(w4038 | w149);
assign w2013 = v743;
assign v744 = ~(w3798 | w278);
assign w2014 = v744;
assign v745 = ~(w3299 | w529);
assign w2015 = v745;
assign w2016 = w3094 & w431;
assign w2017 = ~w2020 & w2705;
assign w2018 = ~w2324 & w991;
assign w2019 = w1830 & ~w3168;
assign w2020 = ~w1504 & w1479;
assign v746 = ~(w1504 | w3191);
assign w2021 = v746;
assign v747 = ~(w777 | w2771);
assign w2022 = v747;
assign w2023 = w4093 & w137;
assign w2024 = ~w51 & w3141;
assign w2025 = ~w893 & w3794;
assign v748 = ~(w1928 | w2782);
assign w2026 = v748;
assign v749 = ~(w1275 | w3678);
assign w2027 = v749;
assign v750 = ~(w2446 | w3857);
assign w2028 = v750;
assign w2029 = ~w303 & w1662;
assign v751 = ~(w2515 | w1750);
assign w2030 = v751;
assign w2031 = ~w1010 & w3295;
assign v752 = ~(w372 | w943);
assign w2032 = v752;
assign v753 = ~(w3929 | w3905);
assign w2033 = v753;
assign v754 = ~(w579 | w700);
assign w2034 = v754;
assign w2035 = ~pi366 & pi207;
assign v755 = ~(w3041 | w2837);
assign w2036 = v755;
assign w2037 = w718 & w2161;
assign w2038 = w2834 & ~w1333;
assign w2039 = w3092 & w518;
assign w2040 = w2717 & ~w657;
assign w2041 = w3394 & ~w1469;
assign w2042 = w3630 & ~w2009;
assign v756 = ~(w4087 | w3259);
assign w2043 = v756;
assign w2044 = w3690 & w961;
assign w2045 = ~pi366 & pi206;
assign v757 = ~(w2723 | w3704);
assign w2046 = v757;
assign v758 = ~(w1168 | w3788);
assign w2047 = v758;
assign w2048 = w656 & ~w1899;
assign w2049 = ~pi366 & pi209;
assign v759 = ~(w1458 | w3188);
assign w2050 = v759;
assign v760 = ~(w249 | w2947);
assign w2051 = v760;
assign v761 = ~(w3312 | w1899);
assign w2052 = v761;
assign w2053 = pi123 & w353;
assign v762 = ~(w4159 | w3263);
assign w2054 = v762;
assign w2055 = w3093 & w13;
assign w2056 = w1325 & w644;
assign w2057 = w1447 & w1492;
assign v763 = ~(w58 | w254);
assign w2058 = v763;
assign v764 = ~(w3878 | w2955);
assign w2059 = v764;
assign w2060 = w1570 & w2884;
assign w2061 = (~w973 & w1143) | (~w973 & w3915) | (w1143 & w3915);
assign v765 = ~(w2075 | w2496);
assign w2062 = v765;
assign w2063 = w3928 & w1469;
assign w2064 = ~w2250 & w1333;
assign w2065 = ~w355 & w1337;
assign w2066 = ~w1720 & w1397;
assign w2067 = (pi092 & ~w1654) | (pi092 & w3602) | (~w1654 & w3602);
assign v766 = ~(w3262 | w3022);
assign w2068 = v766;
assign w2069 = w1015 & w4181;
assign w2070 = w539 & w2000;
assign v767 = ~(w3671 | w284);
assign w2071 = v767;
assign w2072 = ~w3546 & w1287;
assign v768 = ~(w1054 | w200);
assign w2073 = v768;
assign w2074 = (~w1469 & ~w1660) | (~w1469 & w3523) | (~w1660 & w3523);
assign v769 = ~(w4038 | w3722);
assign w2075 = v769;
assign w2076 = w3260 & w480;
assign w2077 = pi293 & w2362;
assign w2078 = w847 & ~w2378;
assign w2079 = w2046 & ~w2373;
assign v770 = ~(w1219 | w2466);
assign w2080 = v770;
assign v771 = ~(w1718 | w4059);
assign w2081 = v771;
assign w2082 = w800 & ~w244;
assign w2083 = w3216 & ~w337;
assign v772 = ~(w2919 | w1960);
assign w2084 = v772;
assign w2085 = ~w1600 & w117;
assign v773 = ~(w503 | w4068);
assign w2086 = v773;
assign v774 = ~(w485 | w2013);
assign w2087 = v774;
assign w2088 = (w1469 & ~w1394) | (w1469 & w4107) | (~w1394 & w4107);
assign v775 = ~(w4038 | w4087);
assign w2089 = v775;
assign w2090 = w3912 & w3826;
assign w2091 = w2717 & ~w3105;
assign w2092 = w2732 & ~w1469;
assign v776 = ~(w1754 | w422);
assign w2093 = v776;
assign w2094 = ~w1469 & w1005;
assign v777 = ~(w2874 | w3160);
assign w2095 = v777;
assign v778 = ~(w3101 | w171);
assign w2096 = v778;
assign v779 = ~(w954 | w657);
assign w2097 = v779;
assign w2098 = w656 & ~w2209;
assign w2099 = ~w1133 & w3604;
assign w2100 = ~pi366 & pi235;
assign v780 = ~(w494 | w3186);
assign w2101 = v780;
assign w2102 = ~w1192 & w642;
assign v781 = ~(w3878 | w3943);
assign w2103 = v781;
assign w2104 = w950 & ~w408;
assign w2105 = (w1758 & ~w3950) | (w1758 & w1269) | (~w3950 & w1269);
assign w2106 = w3094 & w4147;
assign v782 = ~(w1604 | w2175);
assign w2107 = v782;
assign w2108 = ~w3159 & w2000;
assign w2109 = (w1469 & ~w3570) | (w1469 & w2481) | (~w3570 & w2481);
assign v783 = ~(w3116 | w3726);
assign w2110 = v783;
assign w2111 = w118 & pi098;
assign v784 = ~(w3421 | w3966);
assign w2112 = v784;
assign v785 = ~(w1263 | w1752);
assign w2113 = v785;
assign w2114 = w2005 & w813;
assign w2115 = w1510 & w1469;
assign w2116 = w4082 & w908;
assign w2117 = (pi027 & ~w1654) | (pi027 & w1335) | (~w1654 & w1335);
assign w2118 = w2241 & w1651;
assign v786 = ~(w2757 | w2271);
assign w2119 = v786;
assign w2120 = w2606 & w4047;
assign w2121 = w2966 & ~w2477;
assign v787 = ~(w189 | w2329);
assign w2122 = v787;
assign w2123 = ~w504 & w1581;
assign w2124 = w89 & ~w559;
assign w2125 = w1318 & w361;
assign w2126 = (~w3068 & ~w2082) | (~w3068 & w1958) | (~w2082 & w1958);
assign w2127 = w2438 & w990;
assign v788 = ~(w2979 | w30);
assign w2128 = v788;
assign w2129 = w2324 & w991;
assign v789 = ~(w1661 | w657);
assign w2130 = v789;
assign v790 = ~(w4182 | w1825);
assign w2131 = v790;
assign w2132 = (pi009 & ~w1654) | (pi009 & w3978) | (~w1654 & w3978);
assign v791 = ~(w697 | w3364);
assign w2133 = v791;
assign w2134 = w546 & w1469;
assign w2135 = w175 & w4066;
assign v792 = ~(w48 | w2475);
assign w2136 = v792;
assign v793 = ~(w422 | w3259);
assign w2137 = v793;
assign w2138 = w1570 & w2242;
assign v794 = ~(w954 | w1592);
assign w2139 = v794;
assign v795 = ~(w1136 | w1742);
assign w2140 = v795;
assign v796 = ~(w3386 | w3700);
assign w2141 = v796;
assign w2142 = w2514 & w1128;
assign w2143 = pi269 & w2362;
assign v797 = ~(w1469 | w378);
assign w2144 = v797;
assign w2145 = w426 & w2466;
assign w2146 = w1830 & ~w3462;
assign v798 = ~(w276 | w1718);
assign w2147 = v798;
assign w2148 = ~w97 & w268;
assign w2149 = w3094 & w1060;
assign v799 = ~(w3307 | w3187);
assign w2150 = v799;
assign w2151 = ~w876 & w2612;
assign w2152 = w1199 & ~w4076;
assign v800 = ~(w543 | w739);
assign w2153 = v800;
assign w2154 = w3740 & ~w1469;
assign w2155 = w705 & w2138;
assign w2156 = w1570 & w3028;
assign v801 = ~(w2364 | w2999);
assign w2157 = v801;
assign v802 = ~(w1661 | w1955);
assign w2158 = v802;
assign w2159 = w2315 & ~w1089;
assign w2160 = w1636 & w3925;
assign w2161 = w2936 & w3068;
assign w2162 = w2747 & w4071;
assign v803 = ~(w2804 | w69);
assign w2163 = v803;
assign v804 = ~(w2175 | w557);
assign w2164 = v804;
assign v805 = ~(w823 | w1160);
assign w2165 = v805;
assign w2166 = w2487 & ~w2501;
assign v806 = ~(w2475 | w3131);
assign w2167 = v806;
assign w2168 = (w1469 & ~w624) | (w1469 & w2421) | (~w624 & w2421);
assign v807 = ~(w2799 | w1633);
assign w2169 = v807;
assign w2170 = ~w3068 & w2646;
assign w2171 = pi268 & w2362;
assign w2172 = w1005 & ~w1074;
assign w2173 = w4 & w4015;
assign v808 = ~(w4037 | w1941);
assign w2174 = v808;
assign v809 = ~(w299 | w1034);
assign w2175 = v809;
assign w2176 = w2876 & w1934;
assign w2177 = w1139 & ~w3467;
assign w2178 = w2646 & w3180;
assign v810 = ~(w298 | w3710);
assign w2179 = v810;
assign w2180 = (~w1469 & ~w242) | (~w1469 & w2154) | (~w242 & w2154);
assign v811 = ~(w1459 | w1681);
assign w2181 = v811;
assign v812 = ~(w366 | w660);
assign w2182 = v812;
assign w2183 = w157 & ~w1886;
assign v813 = ~(w4038 | w1955);
assign w2184 = v813;
assign v814 = ~(w2927 | w1809);
assign w2185 = v814;
assign v815 = ~(w3277 | w4159);
assign w2186 = v815;
assign w2187 = ~pi366 & pi225;
assign v816 = ~(w2256 | w1755);
assign w2188 = v816;
assign w2189 = w950 & ~w2838;
assign w2190 = w1878 & w1249;
assign w2191 = w2717 & ~w2955;
assign w2192 = ~pi366 & pi236;
assign w2193 = (pi054 & ~w1654) | (pi054 & w112) | (~w1654 & w112);
assign v817 = ~(w187 | w303);
assign w2194 = v817;
assign w2195 = w1253 & w2225;
assign w2196 = w3094 & w2458;
assign w2197 = w1654 & ~w2;
assign w2198 = w2502 & w2291;
assign w2199 = (~w46 & ~w3129) | (~w46 & w1647) | (~w3129 & w1647);
assign w2200 = w2690 & ~w2633;
assign w2201 = w1689 & w740;
assign w2202 = w3094 & w36;
assign w2203 = (w1318 & w1847) | (w1318 & w1462) | (w1847 & w1462);
assign w2204 = w1547 & w3085;
assign v818 = ~(w4159 | w1604);
assign w2205 = v818;
assign w2206 = w1830 & ~w923;
assign w2207 = (w1469 & ~w74) | (w1469 & w2567) | (~w74 & w2567);
assign v819 = ~(w3749 | w753);
assign w2208 = v819;
assign w2209 = ~w2359 & w4127;
assign w2210 = (w1654 & w1544) | (w1654 & w2261) | (w1544 & w2261);
assign w2211 = w1469 & ~w4015;
assign w2212 = w926 & w1909;
assign v820 = ~(w2936 | w3799);
assign w2213 = v820;
assign w2214 = w2968 & w1182;
assign v821 = ~(w3321 | w912);
assign w2215 = v821;
assign v822 = ~(w4038 | w1633);
assign w2216 = v822;
assign w2217 = pi327 & ~pi366;
assign w2218 = pi136 & ~pi364;
assign w2219 = ~w2411 & w555;
assign w2220 = pi320 & ~pi366;
assign w2221 = w1456 & w4172;
assign w2222 = w3029 & w3839;
assign v823 = ~(w3838 | w2037);
assign w2223 = v823;
assign w2224 = w15 & w138;
assign v824 = ~(w2618 | w1045);
assign w2225 = v824;
assign w2226 = w3094 & w1203;
assign v825 = ~(w3426 | w2475);
assign w2227 = v825;
assign w2228 = ~w2917 & w2124;
assign w2229 = (w3068 & w2936) | (w3068 & w3410) | (w2936 & w3410);
assign w2230 = w1875 & w1561;
assign v826 = ~(w1970 | w2085);
assign w2231 = v826;
assign v827 = ~(w2135 | w2765);
assign w2232 = v827;
assign w2233 = w2550 & w386;
assign v828 = ~(w2531 | w4123);
assign w2234 = v828;
assign w2235 = w3960 & ~w3781;
assign w2236 = pi354 & ~pi366;
assign v829 = ~(w4159 | w3858);
assign w2237 = v829;
assign v830 = ~(w4159 | w3343);
assign w2238 = v830;
assign w2239 = w118 & pi049;
assign v831 = ~(w3930 | w2737);
assign w2240 = v831;
assign w2241 = w2513 & w3703;
assign w2242 = pi151 & ~pi364;
assign w2243 = pi256 & w2362;
assign v832 = ~(w1783 | w2151);
assign w2244 = v832;
assign w2245 = ~w2244 & w381;
assign w2246 = pi075 & w570;
assign w2247 = ~w3094 & w2045;
assign w2248 = (pi093 & ~w1654) | (pi093 & w2337) | (~w1654 & w2337);
assign w2249 = ~w750 & w582;
assign w2250 = w1623 & w2403;
assign v833 = ~(w2106 | w2143);
assign w2251 = v833;
assign w2252 = w1182 & ~w751;
assign w2253 = w1258 & w1654;
assign v834 = ~(w393 | w507);
assign w2254 = v834;
assign w2255 = ~pi366 & pi244;
assign v835 = ~(w3160 | w1164);
assign w2256 = v835;
assign v836 = ~(w954 | w1881);
assign w2257 = v836;
assign v837 = ~(w695 | w3119);
assign w2258 = v837;
assign w2259 = ~w3810 & w4112;
assign w2260 = (w2646 & w2936) | (w2646 & w718) | (w2936 & w718);
assign w2261 = w900 & w1654;
assign w2262 = (w4015 & w1603) | (w4015 & w2392) | (w1603 & w2392);
assign w2263 = pi360 & ~pi366;
assign w2264 = ~w2834 & w1333;
assign w2265 = pi275 & w2362;
assign v838 = ~(w1953 | w1225);
assign w2266 = v838;
assign v839 = ~(w2268 | w991);
assign w2267 = v839;
assign v840 = ~(w2273 | w201);
assign w2268 = v840;
assign w2269 = w3391 & ~w3841;
assign v841 = ~(w558 | w3082);
assign w2270 = v841;
assign w2271 = w2717 & ~w1881;
assign v842 = ~(w209 | w1468);
assign w2272 = v842;
assign w2273 = (w3269 & ~w460) | (w3269 & w3767) | (~w460 & w3767);
assign w2274 = w2827 & w1654;
assign w2275 = ~w3412 & w916;
assign w2276 = ~w4064 & w1080;
assign v843 = ~(w3878 | w1533);
assign w2277 = v843;
assign w2278 = ~pi366 & pi192;
assign w2279 = pi104 & w353;
assign w2280 = w2324 & ~w4047;
assign w2281 = ~w575 & w3345;
assign w2282 = w2717 & ~w3858;
assign w2283 = ~w3094 & w1043;
assign w2284 = (pi061 & ~w1654) | (pi061 & w2390) | (~w1654 & w2390);
assign v844 = ~(w1463 | w1377);
assign w2285 = v844;
assign w2286 = w2519 & w3332;
assign w2287 = ~w50 & w1429;
assign v845 = ~(w2480 | w1516);
assign w2288 = v845;
assign v846 = ~(w1104 | w4159);
assign w2289 = v846;
assign v847 = ~(w3312 | w542);
assign w2290 = v847;
assign w2291 = w4047 & ~w2324;
assign w2292 = ~w2462 & w72;
assign w2293 = w1662 & ~w342;
assign w2294 = w2626 & ~w3100;
assign v848 = ~(w2606 | w1132);
assign w2295 = v848;
assign v849 = ~(w2469 | w3988);
assign w2296 = v849;
assign v850 = ~(w4038 | w1444);
assign w2297 = v850;
assign w2298 = ~w834 & w1061;
assign v851 = ~(w4177 | w584);
assign w2299 = v851;
assign w2300 = (~w1469 & ~w567) | (~w1469 & w2041) | (~w567 & w2041);
assign w2301 = pi318 & ~pi366;
assign v852 = ~(w3438 | w899);
assign w2302 = v852;
assign v853 = ~(w1754 | w3462);
assign w2303 = v853;
assign w2304 = (~w3180 & w3507) | (~w3180 & w3824) | (w3507 & w3824);
assign w2305 = w656 & ~w3964;
assign w2306 = w2056 & w1130;
assign v854 = ~(w4159 | w3131);
assign w2307 = v854;
assign w2308 = ~w1498 & w232;
assign w2309 = w1230 & w3481;
assign w2310 = ~pi366 & pi238;
assign v855 = ~(w1661 | w4105);
assign w2311 = v855;
assign v856 = ~(w800 | w3068);
assign w2312 = v856;
assign v857 = ~(w2799 | w2412);
assign w2313 = v857;
assign v858 = ~(w4159 | w422);
assign w2314 = v858;
assign v859 = ~(w3524 | w3366);
assign w2315 = v859;
assign w2316 = w2836 & ~w649;
assign w2317 = (w1469 & ~w522) | (w1469 & w2449) | (~w522 & w2449);
assign w2318 = pi109 & w353;
assign w2319 = w1570 & w1395;
assign v860 = ~(w2799 | w2209);
assign w2320 = v860;
assign w2321 = w2719 & w2548;
assign w2322 = (~w3747 & ~w2551) | (~w3747 & w3066) | (~w2551 & w3066);
assign w2323 = w853 & w1504;
assign v861 = ~(w2064 | w1923);
assign w2324 = v861;
assign v862 = ~(w347 | w3896);
assign w2325 = v862;
assign w2326 = ~w3929 & w1830;
assign w2327 = pi323 & ~pi366;
assign w2328 = w1199 & ~w1383;
assign w2329 = w1447 & w3179;
assign w2330 = w244 & w3180;
assign w2331 = w183 & w3021;
assign w2332 = (w2018 & w370) | (w2018 & w2974) | (w370 & w2974);
assign v863 = ~(w3929 | w4159);
assign w2333 = v863;
assign w2334 = (w3380 & ~w3992) | (w3380 & w42) | (~w3992 & w42);
assign w2335 = (w850 & w3223) | (w850 & w3012) | (w3223 & w3012);
assign v864 = ~(w1662 | w3625);
assign w2336 = v864;
assign w2337 = w118 & pi093;
assign w2338 = w1878 & w1005;
assign w2339 = pi101 & w570;
assign w2340 = w1487 & w153;
assign w2341 = ~w3664 & w3649;
assign w2342 = w1759 & w4072;
assign v865 = ~(w3160 | w2412);
assign w2343 = v865;
assign w2344 = ~pi366 & pi242;
assign v866 = ~(w2394 | w989);
assign w2345 = v866;
assign w2346 = w3094 & w527;
assign v867 = ~(w1012 | w228);
assign w2347 = v867;
assign v868 = ~(w3312 | w3722);
assign w2348 = v868;
assign v869 = ~(w3402 | w953);
assign w2349 = v869;
assign v870 = ~(w1803 | w2726);
assign w2350 = v870;
assign w2351 = pi360 & ~w2362;
assign w2352 = (w1654 & w2453) | (w1654 & w3471) | (w2453 & w3471);
assign w2353 = w1654 & ~w1991;
assign w2354 = w376 & w2397;
assign w2355 = (w442 & ~w1638) | (w442 & w243) | (~w1638 & w243);
assign w2356 = (w2750 & ~w3917) | (w2750 & w1302) | (~w3917 & w1302);
assign v871 = ~(pi362 | pi363);
assign w2357 = v871;
assign w2358 = ~w2336 & w3097;
assign w2359 = ~w3094 & w2699;
assign w2360 = w539 & w863;
assign w2361 = ~w1745 & w3377;
assign w2362 = pi366 & ~pi367;
assign v872 = ~(w3312 | w3343);
assign w2363 = v872;
assign v873 = ~(w179 | w3878);
assign w2364 = v873;
assign v874 = ~(w986 | w305);
assign w2365 = v874;
assign v875 = ~(w3106 | w988);
assign w2366 = v875;
assign v876 = ~(w2260 | w2706);
assign w2367 = v876;
assign w2368 = w481 & w2790;
assign v877 = ~(w2202 | w3600);
assign w2369 = v877;
assign w2370 = pi131 & w1570;
assign w2371 = ~w3094 & w3278;
assign v878 = ~(w3160 | w3263);
assign w2372 = v878;
assign v879 = ~(w3235 | w2382);
assign w2373 = v879;
assign v880 = ~(w3822 | w851);
assign w2374 = v880;
assign v881 = ~(w3312 | w920);
assign w2375 = v881;
assign w2376 = w4046 & w605;
assign v882 = ~(w1754 | w3263);
assign w2377 = v882;
assign w2378 = w2409 & w952;
assign w2379 = (pi042 & ~w1654) | (pi042 & w2645) | (~w1654 & w2645);
assign w2380 = w3466 & w4015;
assign w2381 = ~w1889 & w488;
assign w2382 = w2761 & w2824;
assign w2383 = (~w1403 & w2679) | (~w1403 & w1345) | (w2679 & w1345);
assign v883 = ~(w1970 | w3977);
assign w2384 = v883;
assign w2385 = w118 & pi032;
assign w2386 = w3094 & w556;
assign w2387 = w2140 & w3628;
assign w2388 = w2717 & ~w557;
assign w2389 = w5 & w2720;
assign w2390 = w118 & pi061;
assign v884 = ~(w2425 | w1453);
assign w2391 = v884;
assign w2392 = w2480 & w4015;
assign w2393 = w361 & ~w2817;
assign w2394 = w519 & w2460;
assign v885 = ~(w2036 | w3951);
assign w2395 = v885;
assign w2396 = (~w1469 & ~w2433) | (~w1469 & w2454) | (~w2433 & w2454);
assign w2397 = w2357 & w3118;
assign w2398 = w4084 & w1131;
assign w2399 = w3067 & w3505;
assign w2400 = pi311 & ~pi366;
assign v886 = ~(w1754 | w149);
assign w2401 = v886;
assign v887 = ~(w1661 | w3385);
assign w2402 = v887;
assign w2403 = w1942 & w2445;
assign w2404 = w1431 & w1654;
assign v888 = ~(w1719 | w1972);
assign w2405 = v888;
assign w2406 = w3094 & w2301;
assign v889 = ~(w1872 | w2478);
assign w2407 = v889;
assign v890 = ~(w3287 | w480);
assign w2408 = v890;
assign w2409 = w2543 & w2980;
assign w2410 = w118 & pi041;
assign w2411 = ~w1551 & w3415;
assign w2412 = ~w1292 & w1099;
assign v891 = ~(w1661 | w3168);
assign w2413 = v891;
assign w2414 = w3650 & w3862;
assign v892 = ~(w2800 | w905);
assign w2415 = v892;
assign w2416 = ~w3969 & w3543;
assign v893 = ~(w2517 | w1705);
assign w2417 = v893;
assign w2418 = w2717 & ~w3943;
assign w2419 = ~w2624 & w3390;
assign v894 = ~(w2004 | w879);
assign w2420 = v894;
assign w2421 = w3808 & w1469;
assign v895 = ~(w3899 | w3692);
assign w2422 = v895;
assign w2423 = (w1469 & ~w2369) | (w1469 & w4165) | (~w2369 & w4165);
assign w2424 = w2373 & w3179;
assign w2425 = (w1504 & ~w126) | (w1504 & w2323) | (~w126 & w2323);
assign v896 = ~(w1754 | w657);
assign w2426 = v896;
assign w2427 = pi040 & w570;
assign w2428 = w2484 & ~w138;
assign w2429 = w652 & w3512;
assign v897 = ~(w1428 | w2704);
assign w2430 = v897;
assign w2431 = (w838 & w1849) | (w838 & w568) | (w1849 & w568);
assign w2432 = w2420 & ~w3589;
assign v898 = ~(w2869 | w2696);
assign w2433 = v898;
assign v899 = ~(w3399 | w1151);
assign w2434 = v899;
assign w2435 = ~w2123 & w1830;
assign w2436 = (~w361 & ~w2070) | (~w361 & w4156) | (~w2070 & w4156);
assign v900 = ~(w4010 | w1139);
assign w2437 = v900;
assign w2438 = w1790 & w2165;
assign w2439 = w95 & w3941;
assign w2440 = ~w141 & w2315;
assign w2441 = w1301 & ~w2967;
assign w2442 = w3630 & ~w3293;
assign w2443 = w4000 & w3062;
assign w2444 = (w1767 & ~w1310) | (w1767 & w1652) | (~w1310 & w1652);
assign w2445 = w817 & w3670;
assign v901 = ~(w3878 | w920);
assign w2446 = v901;
assign w2447 = pi060 & w570;
assign v902 = ~(w1661 | w357);
assign w2448 = v902;
assign w2449 = w484 & w1469;
assign w2450 = w2987 & w215;
assign v903 = ~(w4074 | w165);
assign w2451 = v903;
assign v904 = ~(w954 | w1604);
assign w2452 = v904;
assign w2453 = pi022 & w570;
assign w2454 = w3541 & ~w1469;
assign v905 = ~(w210 | w2581);
assign w2455 = v905;
assign v906 = ~(w954 | w3858);
assign w2456 = v906;
assign w2457 = pi278 & w2362;
assign w2458 = pi337 & ~pi366;
assign v907 = ~(w59 | w1788);
assign w2459 = v907;
assign w2460 = ~w4010 & w1139;
assign w2461 = ~w4074 & w4065;
assign w2462 = ~w3176 & w1494;
assign w2463 = w1527 & w3513;
assign v908 = ~(w46 | w3179);
assign w2464 = v908;
assign w2465 = pi083 & w570;
assign w2466 = ~w860 & w3061;
assign v909 = ~(w376 | w2396);
assign w2467 = v909;
assign w2468 = w2443 & ~w11;
assign w2469 = ~w2046 & w2424;
assign w2470 = ~w2280 & w1114;
assign w2471 = ~w3094 & w3070;
assign w2472 = w118 & pi019;
assign w2473 = (w1654 & w3641) | (w1654 & w180) | (w3641 & w180);
assign v910 = ~(w4169 | w4166);
assign w2474 = v910;
assign v911 = ~(w1771 | w1075);
assign w2475 = v911;
assign w2476 = (w1654 & w2427) | (w1654 & w703) | (w2427 & w703);
assign v912 = ~(w4071 | w1429);
assign w2477 = v912;
assign w2478 = pi261 & w2362;
assign v913 = ~(w539 | w2000);
assign w2479 = v913;
assign w2480 = (~w1469 & ~w767) | (~w1469 & w111) | (~w767 & w111);
assign w2481 = w3427 & w1469;
assign w2482 = (w226 & w888) | (w226 & w936) | (w888 & w936);
assign w2483 = pi026 & w570;
assign v914 = ~(w3454 | w3723);
assign w2484 = v914;
assign v915 = ~(w3312 | w557);
assign w2485 = v915;
assign w2486 = w806 & w3067;
assign v916 = ~(w1725 | w1306);
assign w2487 = v916;
assign w2488 = ~w2316 & w832;
assign v917 = ~(w294 | w2440);
assign w2489 = v917;
assign w2490 = pi304 & ~pi366;
assign w2491 = w3073 & w2415;
assign w2492 = ~w58 & w2312;
assign v918 = ~(w2690 | w3269);
assign w2493 = v918;
assign v919 = ~(w4059 | w3301);
assign w2494 = v919;
assign w2495 = (~w123 & w28) | (~w123 & w1584) | (w28 & w1584);
assign v920 = ~(w1754 | w920);
assign w2496 = v920;
assign v921 = ~(w1447 | w3443);
assign w2497 = v921;
assign v922 = ~(w1115 | w1602);
assign w2498 = v922;
assign w2499 = w1830 & ~w1533;
assign w2500 = w208 & w2882;
assign w2501 = ~w15 & w1319;
assign w2502 = ~w2893 & w991;
assign w2503 = pi158 & w1570;
assign v923 = ~(w2393 | w2904);
assign w2504 = v923;
assign v924 = ~(w3566 | w1613);
assign w2505 = v924;
assign w2506 = ~w2189 & w114;
assign w2507 = w698 & w1758;
assign w2508 = pi281 & w2362;
assign w2509 = (w1654 & w3529) | (w1654 & w2722) | (w3529 & w2722);
assign w2510 = w4015 & ~w835;
assign w2511 = pi172 & w1570;
assign w2512 = w3801 & w1654;
assign w2513 = w2090 & w458;
assign w2514 = w3254 & w2653;
assign w2515 = ~w19 & w1493;
assign w2516 = w1830 & ~w149;
assign v925 = ~(w3199 | w4185);
assign w2517 = v925;
assign v926 = ~(w2123 | w1754);
assign w2518 = v926;
assign v927 = ~(w2774 | w2387);
assign w2519 = v927;
assign v928 = ~(w3367 | w1939);
assign w2520 = v928;
assign w2521 = w1654 & ~w2769;
assign v929 = ~(w3905 | w557);
assign w2522 = v929;
assign v930 = ~(w1319 | w648);
assign w2523 = v930;
assign w2524 = w962 & ~w1469;
assign w2525 = w1806 & ~w1175;
assign w2526 = w2444 & w3068;
assign w2527 = w378 & ~w3221;
assign w2528 = ~w800 & w58;
assign v931 = ~(w2175 | w149);
assign w2529 = v931;
assign v932 = ~(w2016 | w2243);
assign w2530 = v932;
assign w2531 = ~w2140 & w2437;
assign w2532 = pi141 & ~pi364;
assign w2533 = w521 & w2293;
assign v933 = ~(w837 | w3609);
assign w2534 = v933;
assign w2535 = ~w1820 & w737;
assign w2536 = (~w1469 & ~w3440) | (~w1469 & w733) | (~w3440 & w733);
assign v934 = ~(w1970 | w1444);
assign w2537 = v934;
assign v935 = ~(w3259 | w498);
assign w2538 = v935;
assign w2539 = (w3180 & ~w3799) | (w3180 & w66) | (~w3799 & w66);
assign w2540 = w2672 & w645;
assign w2541 = pi014 & w570;
assign v936 = ~(w846 | w3067);
assign w2542 = v936;
assign w2543 = w2760 & w53;
assign v937 = ~(w1904 | w2311);
assign w2544 = v937;
assign w2545 = ~w455 & w1317;
assign w2546 = w3504 & w1654;
assign v938 = ~(w1213 | w664);
assign w2547 = v938;
assign w2548 = w1489 & w166;
assign v939 = ~(w974 | w1463);
assign w2549 = v939;
assign v940 = ~(w3621 | w1618);
assign w2550 = v940;
assign v941 = ~(w1274 | w340);
assign w2551 = v941;
assign w2552 = ~w879 & w4004;
assign w2553 = pi102 & w353;
assign w2554 = w1504 & ~w1007;
assign v942 = ~(w1931 | w3191);
assign w2555 = v942;
assign w2556 = w1826 & ~w1243;
assign v943 = ~(w2205 | w2216);
assign w2557 = v943;
assign w2558 = w324 & w1425;
assign w2559 = w3728 & w2240;
assign w2560 = w2461 & w3128;
assign w2561 = pi309 & ~pi366;
assign v944 = ~(w3437 | w4162);
assign w2562 = v944;
assign w2563 = w3583 & w159;
assign w2564 = w1041 & ~w3683;
assign v945 = ~(w226 | w860);
assign w2565 = v945;
assign w2566 = w800 & ~w2936;
assign w2567 = w725 & w1469;
assign v946 = ~(w476 | w473);
assign w2568 = v946;
assign w2569 = w1902 & w4100;
assign w2570 = (w1654 & w1466) | (w1654 & w2546) | (w1466 & w2546);
assign v947 = ~(w3878 | w3964);
assign w2571 = v947;
assign w2572 = w1990 & w1578;
assign v948 = ~(w539 | w846);
assign w2573 = v948;
assign w2574 = ~w2140 & w4010;
assign w2575 = (w1080 & ~w2429) | (w1080 & w1248) | (~w2429 & w1248);
assign w2576 = pi055 & w353;
assign w2577 = ~w1673 & w1830;
assign w2578 = ~w3094 & w2278;
assign w2579 = w130 & ~w551;
assign w2580 = w3655 & w1257;
assign v949 = ~(w954 | w2955);
assign w2581 = v949;
assign v950 = ~(w2799 | w422);
assign w2582 = v950;
assign v951 = ~(w1607 | w2475);
assign w2583 = v951;
assign w2584 = (~w1469 & ~w251) | (~w1469 & w3473) | (~w251 & w3473);
assign w2585 = pi138 & ~pi364;
assign w2586 = w787 & w2233;
assign w2587 = pi164 & w1570;
assign v952 = ~(w1267 | w3736);
assign w2588 = v952;
assign v953 = ~(w1933 | w2331);
assign w2589 = v953;
assign w2590 = ~w1301 & w1479;
assign v954 = ~(w1661 | w923);
assign w2591 = v954;
assign w2592 = w1301 & w774;
assign w2593 = (w2765 & w1400) | (w2765 & w2677) | (w1400 & w2677);
assign w2594 = ~w1469 & w2626;
assign w2595 = ~w2125 & w3766;
assign v955 = ~(w1089 | w964);
assign w2596 = v955;
assign w2597 = w411 & w1654;
assign w2598 = pi142 & w1570;
assign v956 = ~(w731 | w1583);
assign w2599 = v956;
assign w2600 = (w3887 & ~w3378) | (w3887 & w549) | (~w3378 & w549);
assign w2601 = w2420 & ~w2315;
assign w2602 = w1944 & w3796;
assign v957 = ~(w682 | w3555);
assign w2603 = v957;
assign v958 = ~(w1096 | w945);
assign w2604 = v958;
assign w2605 = w4074 & w4065;
assign v959 = ~(w2268 | w2324);
assign w2606 = v959;
assign w2607 = w656 & ~w91;
assign v960 = ~(w2751 | w666);
assign w2608 = v960;
assign w2609 = (w1654 & w858) | (w1654 & w3316) | (w858 & w3316);
assign w2610 = w1989 & w3534;
assign w2611 = w169 & w3192;
assign w2612 = w1734 & w3616;
assign v961 = ~(w608 | w272);
assign w2613 = v961;
assign w2614 = ~w1330 & w335;
assign w2615 = w366 & ~w3727;
assign w2616 = (w1082 & w1455) | (w1082 & w2803) | (w1455 & w2803);
assign v962 = ~(w3162 | w3052);
assign w2617 = v962;
assign v963 = ~(w4159 | w3462);
assign w2618 = v963;
assign w2619 = w3808 & ~w1469;
assign v964 = ~(w2805 | w2452);
assign w2620 = v964;
assign w2621 = ~w3068 & w2936;
assign w2622 = w2482 & w354;
assign v965 = ~(w3878 | w357);
assign w2623 = v965;
assign v966 = ~(w967 | w1707);
assign w2624 = v966;
assign v967 = ~(w2475 | w3317);
assign w2625 = v967;
assign w2626 = w930 & w2006;
assign w2627 = w3094 & w87;
assign v968 = ~(w435 | w3179);
assign w2628 = v968;
assign w2629 = w1255 & w1677;
assign w2630 = w1570 & w1090;
assign v969 = ~(w2210 | w1058);
assign w2631 = v969;
assign w2632 = ~w3094 & w1279;
assign v970 = ~(w2667 | w4059);
assign w2633 = v970;
assign w2634 = (~w1469 & ~w1704) | (~w1469 & w3556) | (~w1704 & w3556);
assign w2635 = ~w217 & w3180;
assign v971 = ~(w3644 | w1788);
assign w2636 = v971;
assign w2637 = w3498 & ~w1024;
assign w2638 = ~w1814 & w390;
assign w2639 = ~w3498 & w1024;
assign w2640 = (~w1469 & ~w1748) | (~w1469 & w2866) | (~w1748 & w2866);
assign v972 = ~(w3576 | w3156);
assign w2641 = v972;
assign w2642 = w3203 & w3423;
assign w2643 = w426 & w3406;
assign v973 = ~(w954 | w794);
assign w2644 = v973;
assign w2645 = w118 & pi042;
assign v974 = ~(w459 | w3439);
assign w2646 = v974;
assign v975 = ~(w3312 | w3385);
assign w2647 = v975;
assign w2648 = pi305 & ~pi366;
assign w2649 = w118 & pi066;
assign w2650 = w378 & ~w1276;
assign w2651 = (w324 & ~w571) | (w324 & w273) | (~w571 & w273);
assign v976 = ~(w2475 | w1633);
assign w2652 = v976;
assign v977 = ~(w2238 | w1098);
assign w2653 = v977;
assign v978 = ~(w4038 | w542);
assign w2654 = v978;
assign v979 = ~(w2986 | w1905);
assign w2655 = v979;
assign w2656 = (w1654 & w3895) | (w1654 & w2935) | (w3895 & w2935);
assign v980 = ~(w4038 | w3426);
assign w2657 = v980;
assign v981 = ~(w3424 | w2571);
assign w2658 = v981;
assign w2659 = w574 & w2474;
assign w2660 = (~w1469 & ~w1356) | (~w1469 & w1792) | (~w1356 & w1792);
assign v982 = ~(w2011 | w1554);
assign w2661 = v982;
assign v983 = ~(w2317 | w3149);
assign w2662 = v983;
assign w2663 = (w1089 & ~w2440) | (w1089 & w1826) | (~w2440 & w1826);
assign w2664 = ~pi366 & pi234;
assign w2665 = ~w4041 & w3984;
assign w2666 = w3687 & w3488;
assign w2667 = (~w1469 & ~w522) | (~w1469 & w1696) | (~w522 & w1696);
assign v984 = ~(w3354 | w175);
assign w2668 = v984;
assign w2669 = w1919 & w3038;
assign v985 = ~(w163 | w2197);
assign w2670 = v985;
assign w2671 = w3243 & w2498;
assign w2672 = w2195 & w2450;
assign w2673 = w2062 & w3071;
assign w2674 = ~pi058 & w570;
assign v986 = ~(w2164 | w1937);
assign w2675 = v986;
assign v987 = ~(w764 | w1863);
assign w2676 = v987;
assign w2677 = w2135 & w2765;
assign v988 = ~(w1396 | w3225);
assign w2678 = v988;
assign w2679 = w3694 & w2461;
assign w2680 = w118 & pi070;
assign w2681 = ~w2817 & w1812;
assign v989 = ~(w2898 | w2120);
assign w2682 = v989;
assign v990 = ~(w3312 | w794);
assign w2683 = v990;
assign w2684 = pi257 & w2362;
assign w2685 = ~w1620 & w1746;
assign v991 = ~(w1575 | w2333);
assign w2686 = v991;
assign w2687 = pi081 & w570;
assign v992 = ~(w755 | w185);
assign w2688 = v992;
assign w2689 = w378 & ~w1097;
assign w2690 = w3062 & w930;
assign w2691 = (w442 & w1658) | (w442 & w2355) | (w1658 & w2355);
assign w2692 = (w1662 & ~w946) | (w1662 & w2029) | (~w946 & w2029);
assign w2693 = (w3422 & ~w1101) | (w3422 & w1262) | (~w1101 & w1262);
assign w2694 = w1776 & ~w1469;
assign w2695 = w1139 & w1057;
assign w2696 = pi295 & w2362;
assign w2697 = ~w2668 & w403;
assign v993 = ~(w482 | w1519);
assign w2698 = v993;
assign w2699 = ~pi366 & pi196;
assign w2700 = (pi116 & ~w1654) | (pi116 & w1238) | (~w1654 & w1238);
assign w2701 = w2588 & w3472;
assign w2702 = pi161 & ~pi364;
assign w2703 = ~w1 & w203;
assign v994 = ~(w1970 | w2209);
assign w2704 = v994;
assign w2705 = (~w1054 & ~w490) | (~w1054 & w1861) | (~w490 & w1861);
assign v995 = ~(w2646 | w157);
assign w2706 = v995;
assign w2707 = w1512 & w3351;
assign w2708 = (w1469 & ~w242) | (w1469 & w3853) | (~w242 & w3853);
assign w2709 = pi265 & w2362;
assign w2710 = (w1199 & w2634) | (w1199 & w3748) | (w2634 & w3748);
assign w2711 = w3828 & w1093;
assign w2712 = w1246 & w1469;
assign w2713 = w118 & pi007;
assign w2714 = ~pi366 & pi217;
assign v996 = ~(w2102 | w1645);
assign w2715 = v996;
assign v997 = ~(w1970 | w3385);
assign w2716 = v997;
assign w2717 = w2799 & ~w38;
assign v998 = ~(w178 | w3288);
assign w2718 = v998;
assign v999 = ~(w4096 | w1226);
assign w2719 = v999;
assign w2720 = w2477 & ~w200;
assign v1000 = ~(w3160 | w422);
assign w2721 = v1000;
assign w2722 = w2511 & w1654;
assign w2723 = (w3422 & ~w2414) | (w3422 & w4009) | (~w2414 & w4009);
assign w2724 = ~w3179 & w175;
assign w2725 = pi006 & w570;
assign w2726 = w2428 & w3821;
assign w2727 = ~w1373 & w679;
assign w2728 = w3191 & ~w1412;
assign v1001 = ~(w4038 | w2955);
assign w2729 = v1001;
assign w2730 = w2865 & w3096;
assign w2731 = w2929 & w3867;
assign w2732 = ~w3094 & w2783;
assign v1002 = ~(w954 | w3105);
assign w2733 = v1002;
assign w2734 = ~w373 & w3375;
assign w2735 = w118 & pi034;
assign v1003 = ~(w3878 | w3263);
assign w2736 = v1003;
assign v1004 = ~(w954 | w557);
assign w2737 = v1004;
assign w2738 = w656 & ~w923;
assign v1005 = ~(w3307 | w562);
assign w2739 = v1005;
assign v1006 = ~(w1661 | w422);
assign w2740 = v1006;
assign v1007 = ~(w690 | w3785);
assign w2741 = v1007;
assign w2742 = w3431 & w4102;
assign w2743 = pi175 & w1570;
assign w2744 = w1570 & w3329;
assign v1008 = ~(w1819 | w2423);
assign w2745 = v1008;
assign w2746 = ~w1157 & w1446;
assign w2747 = w226 & w183;
assign w2748 = w2179 & ~w2580;
assign w2749 = ~pi366 & pi223;
assign v1009 = ~(w354 | w1007);
assign w2750 = v1009;
assign v1010 = ~(w179 | w2475);
assign w2751 = v1010;
assign v1011 = ~(w2175 | w1955);
assign w2752 = v1011;
assign v1012 = ~(w4038 | w398);
assign w2753 = v1012;
assign w2754 = w3094 & w3040;
assign w2755 = (pi057 & ~w1654) | (pi057 & w168) | (~w1654 & w168);
assign v1013 = ~(w2799 | w3343);
assign w2756 = v1013;
assign v1014 = ~(w4159 | w1533);
assign w2757 = v1014;
assign w2758 = (pi003 & ~w1654) | (pi003 & w2768) | (~w1654 & w2768);
assign w2759 = ~w3094 & w2749;
assign v1015 = ~(w2925 | w1176);
assign w2760 = v1015;
assign w2761 = w1367 & w675;
assign w2762 = w2244 & ~w1348;
assign w2763 = w364 & ~w2332;
assign w2764 = w1469 & w3669;
assign v1016 = ~(w828 | w3771);
assign w2765 = v1016;
assign v1017 = ~(w3246 | w3332);
assign w2766 = v1017;
assign w2767 = (w1469 & ~w2299) | (w1469 & w255) | (~w2299 & w255);
assign w2768 = w118 & pi003;
assign v1018 = ~(w2941 | w1208);
assign w2769 = v1018;
assign w2770 = (pi007 & ~w1654) | (pi007 & w2713) | (~w1654 & w2713);
assign w2771 = ~w876 & w2398;
assign w2772 = w1830 & ~w1164;
assign w2773 = w2557 & w1885;
assign v1019 = ~(w2140 | w3628);
assign w2774 = v1019;
assign w2775 = w3922 & w3639;
assign w2776 = (~w2373 & w4113) | (~w2373 & w427) | (w4113 & w427);
assign v1020 = ~(w219 | w2231);
assign w2777 = v1020;
assign w2778 = pi000 & w570;
assign w2779 = pi035 & w353;
assign w2780 = (w1654 & w2997) | (w1654 & w3057) | (w2997 & w3057);
assign v1021 = ~(w156 | w3688);
assign w2781 = v1021;
assign w2782 = w950 & ~w1448;
assign w2783 = ~pi366 & pi230;
assign w2784 = w3094 & w99;
assign v1022 = ~(w3746 | w1732);
assign w2785 = v1022;
assign v1023 = ~(w4067 | w223);
assign w2786 = v1023;
assign w2787 = ~w1469 & w2443;
assign w2788 = ~w1318 & w3747;
assign w2789 = w1443 & ~w1469;
assign w2790 = w1614 & w2841;
assign v1024 = ~(w3160 | w498);
assign w2791 = v1024;
assign w2792 = ~w3994 & w1630;
assign v1025 = ~(w1595 | w3325);
assign w2793 = v1025;
assign w2794 = ~w179 & w1830;
assign w2795 = w1593 & w583;
assign v1026 = ~(w3277 | w4038);
assign w2796 = v1026;
assign w2797 = w3904 & w4111;
assign w2798 = ~w839 & w3422;
assign v1027 = ~(w4069 | w3304);
assign w2799 = v1027;
assign v1028 = ~(w954 | w448);
assign w2800 = v1028;
assign w2801 = w2861 & w1513;
assign v1029 = ~(w1673 | w1754);
assign w2802 = v1029;
assign w2803 = ~w2822 & w1082;
assign w2804 = (w973 & w1135) | (w973 & w2857) | (w1135 & w2857);
assign v1030 = ~(w2175 | w3858);
assign w2805 = v1030;
assign w2806 = ~w3812 & w1587;
assign w2807 = w1678 & ~w24;
assign w2808 = (w1654 & w3885) | (w1654 & w71) | (w3885 & w71);
assign w2809 = w805 & ~w1469;
assign w2810 = ~w836 & w2199;
assign w2811 = (~w1469 & ~w3570) | (~w1469 & w1051) | (~w3570 & w1051);
assign w2812 = w1830 & ~w3343;
assign w2813 = w942 & w1001;
assign w2814 = pi140 & w1570;
assign w2815 = (~w2574 & ~w3085) | (~w2574 & w1481) | (~w3085 & w1481);
assign v1031 = ~(w2646 | w800);
assign w2816 = v1031;
assign w2817 = w3159 & ~w539;
assign w2818 = pi078 & w570;
assign v1032 = ~(w2799 | w498);
assign w2819 = v1032;
assign w2820 = w1834 & ~w3988;
assign v1033 = ~(w2584 | w974);
assign w2821 = v1033;
assign w2822 = (w1083 & w3482) | (w1083 & w341) | (w3482 & w341);
assign v1034 = ~(w3878 | w542);
assign w2823 = v1034;
assign w2824 = w2114 & w2637;
assign w2825 = ~w3094 & w548;
assign w2826 = w2365 & w3720;
assign w2827 = pi149 & w1570;
assign w2828 = pi145 & ~pi364;
assign w2829 = w3094 & w120;
assign w2830 = w3531 & w2058;
assign v1035 = ~(w1559 | w3464);
assign w2831 = v1035;
assign w2832 = w2898 & w1132;
assign w2833 = w3094 & w3520;
assign w2834 = w3446 & w3581;
assign w2835 = w350 & w1469;
assign w2836 = ~w1391 & w1989;
assign v1036 = ~(w4069 | w299);
assign w2837 = v1036;
assign v1037 = ~(w2074 | w974);
assign w2838 = v1037;
assign w2839 = (w3669 & w3477) | (w3669 & w1769) | (w3477 & w1769);
assign w2840 = ~w2318 & w2688;
assign w2841 = w192 & w2266;
assign w2842 = w4015 & ~w1912;
assign w2843 = w118 & pi068;
assign v1038 = ~(w1754 | w3848);
assign w2844 = v1038;
assign v1039 = ~(w2993 | w729);
assign w2845 = v1039;
assign v1040 = ~(w3236 | w21);
assign w2846 = v1040;
assign w2847 = w4053 & w1469;
assign v1041 = ~(w1661 | w149);
assign w2848 = v1041;
assign v1042 = ~(w1695 | w308);
assign w2849 = v1042;
assign v1043 = ~(w1195 | w788);
assign w2850 = v1043;
assign w2851 = pi286 & w2362;
assign w2852 = w336 & w2569;
assign w2853 = w2728 & ~w2162;
assign v1044 = ~(w1365 | w3104);
assign w2854 = v1044;
assign v1045 = ~(w1907 | w2313);
assign w2855 = v1045;
assign v1046 = ~(w1970 | w657);
assign w2856 = v1046;
assign w2857 = ~w1143 & w3954;
assign w2858 = (w1388 & w1085) | (w1388 & w669) | (w1085 & w669);
assign w2859 = w2775 & w104;
assign w2860 = w2852 & w2010;
assign v1047 = ~(w3861 | w1729);
assign w2861 = v1047;
assign w2862 = w4015 & ~w316;
assign w2863 = ~w3138 & w3593;
assign w2864 = (~w1469 & ~w1916) | (~w1469 & w2969) | (~w1916 & w2969);
assign w2865 = w291 & w2491;
assign w2866 = w2825 & ~w1469;
assign w2867 = w388 & ~w1469;
assign w2868 = w1040 & w1787;
assign w2869 = w3094 & w4184;
assign v1048 = ~(w1608 | w1691);
assign w2870 = v1048;
assign w2871 = w1318 & ~w3568;
assign w2872 = w2439 & w197;
assign v1049 = ~(w4159 | w3317);
assign w2873 = v1049;
assign w2874 = ~w2825 & w1748;
assign w2875 = w879 & w559;
assign w2876 = w1867 & w3112;
assign w2877 = w2070 & ~w128;
assign w2878 = w2626 & ~w552;
assign w2879 = w373 & ~w3375;
assign v1050 = ~(w4159 | w3964);
assign w2880 = v1050;
assign v1051 = ~(w974 | w700);
assign w2881 = v1051;
assign v1052 = ~(w2533 | w2858);
assign w2882 = v1052;
assign w2883 = ~w2651 & w1640;
assign w2884 = pi143 & ~pi364;
assign w2885 = (pi094 & ~w1654) | (pi094 & w3965) | (~w1654 & w3965);
assign v1053 = ~(w3838 | w3350);
assign w2886 = v1053;
assign v1054 = ~(w3312 | w3168);
assign w2887 = v1054;
assign v1055 = ~(w954 | w3964);
assign w2888 = v1055;
assign w2889 = (w2022 & w3388) | (w2022 & w3676) | (w3388 & w3676);
assign w2890 = w1254 & w3982;
assign w2891 = pi099 & w353;
assign w2892 = (w991 & ~w1250) | (w991 & w1108) | (~w1250 & w1108);
assign v1056 = ~(w3275 | w2928);
assign w2893 = v1056;
assign v1057 = ~(w271 | w3466);
assign w2894 = v1057;
assign v1058 = ~(w3312 | w1955);
assign w2895 = v1058;
assign w2896 = w3591 & w1476;
assign v1059 = ~(w3627 | w2282);
assign w2897 = v1059;
assign w2898 = w2268 & ~w2893;
assign v1060 = ~(w2905 | w3644);
assign w2899 = v1060;
assign v1061 = ~(w1104 | w3878);
assign w2900 = v1061;
assign v1062 = ~(w564 | w3521);
assign w2901 = v1062;
assign v1063 = ~(w1091 | w1921);
assign w2902 = v1063;
assign w2903 = w1776 & w2594;
assign v1064 = ~(w1103 | w3067);
assign w2904 = v1064;
assign w2905 = (~w1469 & ~w108) | (~w1469 & w495) | (~w108 & w495);
assign w2906 = (w1654 & w1252) | (w1654 & w3672) | (w1252 & w3672);
assign w2907 = ~w3094 & w4141;
assign w2908 = (pi034 & ~w1654) | (pi034 & w2735) | (~w1654 & w2735);
assign v1065 = ~(w3160 | w3462);
assign w2909 = v1065;
assign w2910 = w436 & w3320;
assign w2911 = w3239 & w3914;
assign v1066 = ~(w238 | w4145);
assign w2912 = v1066;
assign w2913 = w705 & w1212;
assign w2914 = w3875 & w4055;
assign w2915 = w2717 & ~w3977;
assign w2916 = (pi089 & ~w1654) | (pi089 & w3460) | (~w1654 & w3460);
assign v1067 = ~(w2315 | w964);
assign w2917 = v1067;
assign v1068 = ~(w2816 | w3715);
assign w2918 = v1068;
assign v1069 = ~(w1661 | w3317);
assign w2919 = v1069;
assign w2920 = w118 & pi069;
assign w2921 = pi263 & w2362;
assign w2922 = w2022 & w1139;
assign w2923 = (w324 & ~w720) | (w324 & w833) | (~w720 & w833);
assign w2924 = w2349 & w3802;
assign w2925 = w1830 & ~w3977;
assign w2926 = (pi056 & ~w1654) | (pi056 & w1731) | (~w1654 & w1731);
assign w2927 = (w2594 & ~w1704) | (w2594 & w1791) | (~w1704 & w1791);
assign w2928 = ~w1330 & w2669;
assign w2929 = w2960 & w4018;
assign w2930 = w818 & w1654;
assign w2931 = ~w866 & w3373;
assign w2932 = w1116 & w601;
assign w2933 = ~w2599 & w2148;
assign w2934 = w2717 & ~w1140;
assign w2935 = w2503 & w1654;
assign v1070 = ~(w1858 | w312);
assign w2936 = v1070;
assign w2937 = ~w3094 & w3117;
assign w2938 = w656 & ~w1140;
assign w2939 = w118 & pi013;
assign v1071 = ~(w2121 | w2389);
assign w2940 = v1071;
assign w2941 = (w1469 & ~w108) | (w1469 & w3114) | (~w108 & w3114);
assign w2942 = ~w3749 & w2122;
assign w2943 = pi357 & ~pi366;
assign v1072 = ~(w1970 | w1899);
assign w2944 = v1072;
assign v1073 = ~(w4159 | w3385);
assign w2945 = v1073;
assign v1074 = ~(w1788 | w3162);
assign w2946 = v1074;
assign w2947 = ~w1358 & w3729;
assign w2948 = w61 & w1811;
assign w2949 = w1469 & w1199;
assign w2950 = w3233 & w2376;
assign v1075 = ~(w3878 | w3977);
assign w2951 = v1075;
assign w2952 = w2717 & ~w3168;
assign w2953 = pi253 & w2362;
assign v1076 = ~(w3814 | w1372);
assign w2954 = v1076;
assign w2955 = ~w2937 & w2272;
assign w2956 = ~w3759 & w462;
assign w2957 = pi180 & w1570;
assign w2958 = w2215 & ~w4143;
assign w2959 = ~w3784 & w4122;
assign v1077 = ~(w1000 | w2043);
assign w2960 = v1077;
assign w2961 = w350 & w955;
assign v1078 = ~(w2799 | w179);
assign w2962 = v1078;
assign v1079 = ~(w3076 | w2536);
assign w2963 = v1079;
assign w2964 = pi174 & w1570;
assign v1080 = ~(w534 | w3871);
assign w2965 = v1080;
assign w2966 = ~w183 & w2565;
assign v1081 = ~(w426 | w2466);
assign w2967 = v1081;
assign w2968 = ~w1340 & w1846;
assign w2969 = w45 & ~w1469;
assign w2970 = w705 & w3000;
assign v1082 = ~(w1516 | w1733);
assign w2971 = v1082;
assign v1083 = ~(w2799 | w3964);
assign w2972 = v1083;
assign w2973 = w3290 & w1624;
assign w2974 = w660 & w2018;
assign v1084 = ~(w3312 | w4105);
assign w2975 = v1084;
assign v1085 = ~(w964 | w961);
assign w2976 = v1085;
assign w2977 = w3770 & w343;
assign w2978 = (~w227 & w961) | (~w227 & w4048) | (w961 & w4048);
assign w2979 = (w1654 & w1472) | (w1654 & w1037) | (w1472 & w1037);
assign w2980 = w2855 & w1954;
assign w2981 = w3614 & w3742;
assign w2982 = w2907 & ~w1469;
assign w2983 = ~w1787 & w1028;
assign w2984 = w1929 & w3198;
assign w2985 = ~w3296 & w1207;
assign v1086 = ~(w4038 | w3462);
assign w2986 = v1086;
assign v1087 = ~(w1068 | w2823);
assign w2987 = v1087;
assign w2988 = w1454 & ~w2989;
assign v1088 = ~(w745 | w1150);
assign w2989 = v1088;
assign v1089 = ~(w3076 | w994);
assign w2990 = v1089;
assign w2991 = pi062 & w570;
assign w2992 = (w4015 & w3342) | (w4015 & w2380) | (w3342 & w2380);
assign v1090 = ~(w2352 | w1384);
assign w2993 = v1090;
assign v1091 = ~(w4159 | w1633);
assign w2994 = v1091;
assign w2995 = (~w361 & w2877) | (~w361 & w3485) | (w2877 & w3485);
assign w2996 = w3791 & w3383;
assign w2997 = pi008 & w570;
assign w2998 = w800 & ~w3180;
assign v1092 = ~(w3277 | w1970);
assign w2999 = v1092;
assign w3000 = w1570 & w1564;
assign w3001 = w165 & ~w3800;
assign v1093 = ~(w2070 | w2542);
assign w3002 = v1093;
assign w3003 = ~w3882 & w2194;
assign w3004 = pi332 & ~pi366;
assign w3005 = ~pi366 & pi220;
assign w3006 = w736 & ~w2484;
assign v1094 = ~(w2584 | w1810);
assign w3007 = v1094;
assign w3008 = w1103 & w1956;
assign w3009 = (w838 & w940) | (w838 & w1807) | (w940 & w1807);
assign w3010 = ~w3929 & w656;
assign w3011 = w705 & w40;
assign w3012 = w2194 & w850;
assign w3013 = w1 & ~w203;
assign w3014 = (w2968 & ~w1837) | (w2968 & w3985) | (~w1837 & w3985);
assign w3015 = w3916 & w1761;
assign w3016 = w372 & w943;
assign w3017 = w3628 & w1139;
assign w3018 = w1830 & ~w1667;
assign w3019 = ~w298 & w327;
assign v1095 = ~(w1673 | w954);
assign w3020 = v1095;
assign w3021 = w226 & w3061;
assign v1096 = ~(w141 | w964);
assign w3022 = v1096;
assign v1097 = ~(w1500 | w4124);
assign w3023 = v1097;
assign w3024 = pi147 & w1570;
assign v1098 = ~(w3259 | w2085);
assign w3025 = v1098;
assign v1099 = ~(w562 | w708);
assign w3026 = v1099;
assign w3027 = w4004 & ~w886;
assign w3028 = pi183 & ~pi364;
assign v1100 = ~(w3516 | w246);
assign w3029 = v1100;
assign w3030 = w705 & w2060;
assign w3031 = w736 & ~w2374;
assign w3032 = w2611 & w1980;
assign v1101 = ~(w3259 | w3263);
assign w3033 = v1101;
assign w3034 = pi039 & w570;
assign v1102 = ~(w425 | w2487);
assign w3035 = v1102;
assign w3036 = w1153 & w2101;
assign v1103 = ~(w1607 | w3312);
assign w3037 = v1103;
assign w3038 = w1643 & w3065;
assign w3039 = ~w1391 & w2596;
assign w3040 = pi316 & ~pi366;
assign v1104 = ~(w2317 | w2074);
assign w3041 = v1104;
assign w3042 = w892 & w2096;
assign v1105 = ~(w1140 | w2475);
assign w3043 = v1105;
assign w3044 = (w2547 & ~w2405) | (w2547 & w3634) | (~w2405 & w3634);
assign w3045 = w2717 & ~w3722;
assign v1106 = ~(w4159 | w923);
assign w3046 = v1106;
assign w3047 = w3969 & ~w3543;
assign w3048 = w225 & w3387;
assign v1107 = ~(w3076 | w889);
assign w3049 = v1107;
assign v1108 = ~(w1661 | w1782);
assign w3050 = v1108;
assign w3051 = ~w2646 & w2936;
assign w3052 = (~w1469 & ~w1793) | (~w1469 & w3242) | (~w1793 & w3242);
assign w3053 = w3535 & w505;
assign v1109 = ~(w1749 | w3817);
assign w3054 = v1109;
assign w3055 = w1830 & ~w91;
assign w3056 = pi271 & w2362;
assign w3057 = w2957 & w1654;
assign w3058 = w3417 & ~w1469;
assign w3059 = pi157 & ~pi364;
assign v1110 = ~(w68 | w172);
assign w3060 = v1110;
assign v1111 = ~(w218 | w2025);
assign w3061 = v1111;
assign w3062 = ~pi362 & pi363;
assign w3063 = w720 & w352;
assign v1112 = ~(w2906 | w639);
assign w3064 = v1112;
assign w3065 = w2793 & w287;
assign w3066 = w3900 & ~w3747;
assign w3067 = ~w2000 & w128;
assign v1113 = ~(w1066 | w2219);
assign w3068 = v1113;
assign w3069 = ~w3582 & w3739;
assign w3070 = ~pi366 & pi246;
assign v1114 = ~(w1505 | w1836);
assign w3071 = v1114;
assign w3072 = ~w2128 & w2358;
assign v1115 = ~(w1341 | w2873);
assign w3073 = v1115;
assign w3074 = w3309 & ~w3405;
assign v1116 = ~(w2799 | w398);
assign w3075 = v1116;
assign w3076 = (w1469 & ~w2530) | (w1469 & w741) | (~w2530 & w741);
assign v1117 = ~(w1780 | w1930);
assign w3077 = v1117;
assign w3078 = w308 & w2690;
assign w3079 = ~w3294 & w1841;
assign v1118 = ~(w3878 | w1444);
assign w3080 = v1118;
assign v1119 = ~(w1661 | w3105);
assign w3081 = v1119;
assign v1120 = ~(w3277 | w3160);
assign w3082 = v1120;
assign v1121 = ~(w3595 | w199);
assign w3083 = v1121;
assign w3084 = ~w3061 & w183;
assign v1122 = ~(w1305 | w808);
assign w3085 = v1122;
assign w3086 = w613 & w462;
assign w3087 = w2626 & ~w3869;
assign w3088 = ~pi366 & pi216;
assign w3089 = w1030 & w1654;
assign v1123 = ~(w1673 | w3259);
assign w3090 = v1123;
assign w3091 = ~w3039 & w2762;
assign v1124 = ~(w3452 | w1840);
assign w3092 = v1124;
assign v1125 = ~(w3020 | w70);
assign w3093 = v1125;
assign v1126 = ~(w561 | w3963);
assign w3094 = v1126;
assign w3095 = w519 & w4094;
assign w3096 = w3577 & w2742;
assign w3097 = ~w3363 & w3500;
assign w3098 = (~w3068 & ~w492) | (~w3068 & w2868) | (~w492 & w2868);
assign v1127 = ~(w3751 | w3434);
assign w3099 = v1127;
assign v1128 = ~(w845 | w487);
assign w3100 = v1128;
assign w3101 = ~w3277 & w1830;
assign w3102 = w4175 & w3816;
assign w3103 = w4053 & w3898;
assign v1129 = ~(w954 | w179);
assign w3104 = v1129;
assign w3105 = ~w3808 & w624;
assign v1130 = ~(w1754 | w4105);
assign w3106 = v1130;
assign w3107 = (w1654 & w1271) | (w1654 & w3991) | (w1271 & w3991);
assign v1131 = ~(w3929 | w2799);
assign w3108 = v1131;
assign w3109 = w800 & ~w2646;
assign w3110 = w3396 & w3255;
assign w3111 = w656 & ~w3858;
assign v1132 = ~(w1829 | w4021);
assign w3112 = v1132;
assign v1133 = ~(w3312 | w1164);
assign w3113 = v1133;
assign w3114 = w1920 & w1469;
assign w3115 = w1005 & ~w2739;
assign w3116 = w3630 & ~w3765;
assign w3117 = ~pi366 & pi245;
assign w3118 = ~pi364 & pi365;
assign v1134 = ~(w2799 | w3426);
assign w3119 = v1134;
assign w3120 = w1249 & ~w3783;
assign w3121 = w2572 & w2924;
assign w3122 = ~pi366 & pi219;
assign w3123 = w2932 & ~w1653;
assign w3124 = ~w1041 & w3683;
assign w3125 = pi188 & w1570;
assign w3126 = ~w2083 & w4144;
assign v1135 = ~(w1318 | w361);
assign w3127 = v1135;
assign w3128 = ~w15 & w138;
assign v1136 = ~(w2497 | w753);
assign w3129 = v1136;
assign w3130 = w1570 & w3059;
assign w3131 = ~w546 & w1704;
assign w3132 = ~w4045 & w3569;
assign v1137 = ~(w1378 | w2994);
assign w3133 = v1137;
assign v1138 = ~(w3881 | w2353);
assign w3134 = v1138;
assign v1139 = ~(w3304 | w1034);
assign w3135 = v1139;
assign w3136 = pi336 & ~pi366;
assign w3137 = w2840 & ~w3721;
assign w3138 = w1775 & ~w2697;
assign w3139 = w2505 & w1411;
assign v1140 = ~(w1826 | w565);
assign w3140 = v1140;
assign v1141 = ~(w3068 | w3659);
assign w3141 = v1141;
assign w3142 = w395 & w1654;
assign v1142 = ~(w3878 | w149);
assign w3143 = v1142;
assign w3144 = ~w3094 & w1032;
assign w3145 = w3531 & ~w157;
assign v1143 = ~(w1970 | w3964);
assign w3146 = v1143;
assign w3147 = w2663 & w1609;
assign w3148 = w3669 & ~w844;
assign w3149 = (~w1469 & ~w848) | (~w1469 & w1518) | (~w848 & w1518);
assign v1144 = ~(w1785 | w2962);
assign w3150 = v1144;
assign v1145 = ~(w1607 | w3878);
assign w3151 = v1145;
assign w3152 = (w1654 & w3034) | (w1654 & w3089) | (w3034 & w3089);
assign w3153 = ~w2228 & w925;
assign v1146 = ~(w1379 | w1134);
assign w3154 = v1146;
assign w3155 = ~w2387 & w433;
assign v1147 = ~(w2799 | w91);
assign w3156 = v1147;
assign w3157 = ~w961 & w3403;
assign w3158 = ~w660 & w2129;
assign v1148 = ~(w4125 | w4097);
assign w3159 = v1148;
assign v1149 = ~(w1892 | w2594);
assign w3160 = v1149;
assign w3161 = w3094 & w2327;
assign w3162 = (w1469 & ~w4139) | (w1469 & w2835) | (~w4139 & w2835);
assign w3163 = pi272 & w2362;
assign w3164 = w489 & w2603;
assign w3165 = w705 & w2319;
assign v1150 = ~(w632 | w265);
assign w3166 = v1150;
assign v1151 = ~(w2175 | w1899);
assign w3167 = v1151;
assign w3168 = ~w3265 & w599;
assign v1152 = ~(w3160 | w3943);
assign w3169 = v1152;
assign v1153 = ~(w4159 | w1607);
assign w3170 = v1153;
assign w3171 = w3282 & w1654;
assign v1154 = ~(w3942 | w540);
assign w3172 = v1154;
assign w3173 = w2936 & ~w3180;
assign v1155 = ~(w1970 | w1604);
assign w3174 = v1155;
assign w3175 = (pi052 & ~w1654) | (pi052 & w323) | (~w1654 & w323);
assign w3176 = pi082 & w353;
assign w3177 = w118 & pi091;
assign w3178 = w3094 & w3491;
assign v1156 = ~(w3956 | w4134);
assign w3179 = v1156;
assign v1157 = ~(w1832 | w724);
assign w3180 = v1157;
assign w3181 = pi033 & w570;
assign w3182 = w3630 & ~w3349;
assign v1158 = ~(w2591 | w2091);
assign w3183 = v1158;
assign w3184 = ~w3183 & w3422;
assign w3185 = w118 & pi074;
assign v1159 = ~(w3878 | w657);
assign w3186 = v1159;
assign w3187 = (~w1469 & ~w478) | (~w1469 & w2867) | (~w478 & w2867);
assign v1160 = ~(w4010 | w3628);
assign w3188 = v1160;
assign w3189 = w1167 & w1035;
assign w3190 = ~pi366 & pi213;
assign v1161 = ~(w3902 | w3123);
assign w3191 = v1161;
assign v1162 = ~(w815 | w1194);
assign w3192 = v1162;
assign v1163 = ~(w845 | w59);
assign w3193 = v1163;
assign v1164 = ~(w3696 | w2634);
assign w3194 = v1164;
assign w3195 = w184 & w1469;
assign v1165 = ~(w2952 | w1077);
assign w3196 = v1165;
assign w3197 = pi277 & w2362;
assign v1166 = ~(w1011 | w1290);
assign w3198 = v1166;
assign w3199 = ~w2268 & w2893;
assign w3200 = (w2374 & ~w1539) | (w2374 & w3680) | (~w1539 & w3680);
assign v1167 = ~(w3430 | w3230);
assign w3201 = v1167;
assign w3202 = ~pi366 & pi202;
assign w3203 = w2773 & w1557;
assign w3204 = w2397 & ~w2899;
assign v1168 = ~(w48 | w1970);
assign w3205 = v1168;
assign v1169 = ~(w4171 | w4185);
assign w3206 = v1169;
assign w3207 = w1573 & ~w1566;
assign v1170 = ~(w541 | w1997);
assign w3208 = v1170;
assign w3209 = ~w286 & w2436;
assign w3210 = w705 & w3444;
assign w3211 = w118 & pi030;
assign v1171 = ~(w1537 | w3774);
assign w3212 = v1171;
assign w3213 = ~w2487 & w12;
assign w3214 = w2663 & ~w2601;
assign v1172 = ~(w1329 | w4060);
assign w3215 = v1172;
assign v1173 = ~(w1299 | w412);
assign w3216 = v1173;
assign w3217 = w510 & w1182;
assign w3218 = w4064 & ~w1080;
assign w3219 = pi028 & w570;
assign w3220 = w2681 & w1318;
assign v1174 = ~(w889 | w579);
assign w3221 = v1174;
assign w3222 = w3590 & w3661;
assign w3223 = w2517 & w1441;
assign w3224 = (w381 & ~w1619) | (w381 & w3536) | (~w1619 & w3536);
assign w3225 = pi288 & w2362;
assign w3226 = (~w157 & ~w2918) | (~w157 & w420) | (~w2918 & w420);
assign v1175 = ~(w1674 | w824);
assign w3227 = v1175;
assign w3228 = w758 & ~w1629;
assign v1176 = ~(w1758 | w3068);
assign w3229 = v1176;
assign w3230 = pi285 & w2362;
assign w3231 = (w389 & ~w4170) | (w389 & w577) | (~w4170 & w577);
assign w3232 = w102 & w196;
assign w3233 = w3640 & w2984;
assign v1177 = ~(w1970 | w3105);
assign w3234 = v1177;
assign w3235 = (w1024 & ~w2761) | (w1024 & w164) | (~w2761 & w164);
assign w3236 = ~w971 & w2863;
assign w3237 = w1976 & ~w1469;
assign v1178 = ~(w1132 | w1688);
assign w3238 = v1178;
assign w3239 = w401 & w3662;
assign v1179 = ~(w4038 | w923);
assign w3240 = v1179;
assign v1180 = ~(w2480 | w2423);
assign w3241 = v1180;
assign w3242 = w528 & ~w1469;
assign v1181 = ~(w1416 | w2290);
assign w3243 = v1181;
assign w3244 = w2801 & w1591;
assign v1182 = ~(w1970 | w3848);
assign w3245 = v1182;
assign w3246 = (w1139 & w2460) | (w1139 & w3017) | (w2460 & w3017);
assign w3247 = w653 & w2988;
assign w3248 = w1417 & w4126;
assign w3249 = ~w2073 & w2441;
assign w3250 = w2578 & w1469;
assign w3251 = w118 & pi044;
assign w3252 = w281 & w1415;
assign v1183 = ~(w533 | w3560);
assign w3253 = v1183;
assign v1184 = ~(w2733 | w3884);
assign w3254 = v1184;
assign v1185 = ~(w2944 | w1612);
assign w3255 = v1185;
assign v1186 = ~(w906 | w394);
assign w3256 = v1186;
assign w3257 = pi279 & w2362;
assign w3258 = w1664 & ~w2697;
assign v1187 = ~(w2787 | w389);
assign w3259 = v1187;
assign v1188 = ~(w648 | w771);
assign w3260 = v1188;
assign w3261 = w1654 & ~w2147;
assign v1189 = ~(w2334 | w706);
assign w3262 = v1189;
assign w3263 = ~w2471 & w1838;
assign v1190 = ~(w3312 | w1782);
assign w3264 = v1190;
assign w3265 = ~w3094 & w689;
assign w3266 = pi260 & w2362;
assign w3267 = pi344 & ~pi366;
assign v1191 = ~(w3905 | w448);
assign w3268 = v1191;
assign w3269 = ~w3962 & w3918;
assign w3270 = w1308 & w1156;
assign v1192 = ~(w1661 | w3848);
assign w3271 = v1192;
assign w3272 = (pi011 & ~w1654) | (pi011 & w3651) | (~w1654 & w3651);
assign w3273 = ~w3615 & w1371;
assign w3274 = (w1654 & w809) | (w1654 & w1753) | (w809 & w1753);
assign w3275 = w1330 & ~w2669;
assign w3276 = w2429 & w1726;
assign w3277 = ~w2732 & w4157;
assign w3278 = ~pi366 & pi226;
assign w3279 = w3003 & ~w792;
assign v1193 = ~(w2294 | w746);
assign w3280 = v1193;
assign w3281 = w470 & ~w2368;
assign w3282 = pi190 & w1570;
assign w3283 = w3864 & w3166;
assign v1194 = ~(w3426 | w2175);
assign w3284 = v1194;
assign w3285 = ~w928 & w2249;
assign v1195 = ~(w1948 | w629);
assign w3286 = v1195;
assign w3287 = ~w2374 & w3006;
assign w3288 = pi282 & w2362;
assign v1196 = ~(w1588 | w4029);
assign w3289 = v1196;
assign v1197 = ~(w234 | w1648);
assign w3290 = v1197;
assign w3291 = w118 & pi071;
assign w3292 = ~w470 & w2368;
assign v1198 = ~(w2811 | w424);
assign w3293 = v1198;
assign w3294 = ~w2268 & w4171;
assign w3295 = w984 & ~w747;
assign w3296 = w1722 & w2229;
assign v1199 = ~(w1661 | w2412);
assign w3297 = v1199;
assign v1200 = ~(w4 | w376);
assign w3298 = v1200;
assign v1201 = ~(w3277 | w2175);
assign w3299 = v1201;
assign w3300 = w2212 & w2707;
assign w3301 = (~w1469 & ~w4157) | (~w1469 & w2092) | (~w4157 & w2092);
assign w3302 = (pi043 & ~w1654) | (pi043 & w631) | (~w1654 & w631);
assign w3303 = (w3683 & w1145) | (w3683 & w3124) | (w1145 & w3124);
assign w3304 = w1469 & w1182;
assign w3305 = w1697 & ~w2215;
assign w3306 = ~w1700 & w1698;
assign w3307 = (w1469 & ~w1950) | (w1469 & w3890) | (~w1950 & w3890);
assign w3308 = pi168 & w1570;
assign w3309 = (~w3191 & ~w5) | (~w3191 & w1813) | (~w5 & w1813);
assign w3310 = w950 & ~w261;
assign w3311 = pi331 & ~pi366;
assign v1202 = ~(w3382 | w2949);
assign w3312 = v1202;
assign w3313 = (w2487 & w32) | (w2487 & w415) | (w32 & w415);
assign w3314 = pi315 & ~pi366;
assign w3315 = ~w827 & w2296;
assign w3316 = w883 & w1654;
assign w3317 = ~w184 & w2407;
assign w3318 = ~w1469 & w3669;
assign v1203 = ~(w1669 | w2684);
assign w3319 = v1203;
assign v1204 = ~(w1796 | w3493);
assign w3320 = v1204;
assign w3321 = (w1654 & w14) | (w1654 & w4153) | (w14 & w4153);
assign w3322 = w354 & ~w2466;
assign w3323 = w3079 & w3494;
assign v1205 = ~(w3259 | w3858);
assign w3324 = v1205;
assign v1206 = ~(w3160 | w3722);
assign w3325 = v1206;
assign w3326 = w2690 & ~w220;
assign w3327 = ~w2373 & w3216;
assign v1207 = ~(w4159 | w1140);
assign w3328 = v1207;
assign w3329 = pi132 & ~pi364;
assign v1208 = ~(w1693 | w3797);
assign w3330 = v1208;
assign w3331 = w3553 & w2981;
assign w3332 = ~w519 & w684;
assign v1209 = ~(w1708 | w1560);
assign w3333 = v1209;
assign w3334 = ~w3094 & w3845;
assign w3335 = w672 & ~w3416;
assign w3336 = pi329 & ~pi366;
assign w3337 = pi148 & w1570;
assign w3338 = w2234 & w743;
assign w3339 = pi105 & w353;
assign w3340 = ~w2424 & w1774;
assign v1210 = ~(w1686 | w4023);
assign w3341 = v1210;
assign w3342 = (~w1469 & ~w1896) | (~w1469 & w2524) | (~w1896 & w2524);
assign w3343 = ~w148 & w3611;
assign v1211 = ~(w2941 | w700);
assign w3344 = v1211;
assign v1212 = ~(w136 | w716);
assign w3345 = v1212;
assign w3346 = w2797 & w3139;
assign w3347 = w1357 & w1141;
assign w3348 = w32 & w4065;
assign v1213 = ~(w901 | w2109);
assign w3349 = v1213;
assign w3350 = (w1028 & ~w1040) | (w1028 & w2983) | (~w1040 & w2983);
assign v1214 = ~(w1963 | w1296);
assign w3351 = v1214;
assign w3352 = w1040 & ~w714;
assign v1215 = ~(w1970 | w3343);
assign w3353 = v1215;
assign w3354 = ~w2046 & w3179;
assign v1216 = ~(w3878 | w3722);
assign w3355 = v1216;
assign w3356 = w2717 & ~w2874;
assign w3357 = w3021 & w1245;
assign v1217 = ~(w3490 | w2970);
assign w3358 = v1217;
assign w3359 = w118 & pi088;
assign w3360 = w1447 & ~w3179;
assign w3361 = ~w2179 & w2580;
assign v1218 = ~(w2799 | w657);
assign w3362 = v1218;
assign w3363 = (w1662 & ~w2931) | (w1662 & w757) | (~w2931 & w757);
assign w3364 = ~w3623 & w2342;
assign v1219 = ~(w2175 | w1667);
assign w3365 = v1219;
assign w3366 = w1338 & w1922;
assign w3367 = w3669 & ~w2081;
assign w3368 = w118 & ~pi118;
assign w3369 = w4039 & ~w430;
assign v1220 = ~(w2521 | w302);
assign w3370 = v1220;
assign w3371 = (w1654 & w2465) | (w1654 & w2274) | (w2465 & w2274);
assign v1221 = ~(w3231 | w2363);
assign w3372 = v1221;
assign v1222 = ~(w77 | w2120);
assign w3373 = v1222;
assign w3374 = w3308 & w1654;
assign w3375 = w4033 & w2586;
assign v1223 = ~(w2375 | w127);
assign w3376 = v1223;
assign v1224 = ~(w433 | w1823);
assign w3377 = v1224;
assign w3378 = w958 & w2430;
assign w3379 = w2411 & ~w1149;
assign v1225 = ~(w1183 | w3302);
assign w3380 = v1225;
assign w3381 = (w1469 & ~w1916) | (w1469 & w280) | (~w1916 & w280);
assign w3382 = ~w1469 & w672;
assign w3383 = w1336 & w3280;
assign w3384 = w2750 & ~w3191;
assign w3385 = ~w1776 & w709;
assign v1226 = ~(w1140 | w2175);
assign w3386 = v1226;
assign v1227 = ~(w3613 | w1627);
assign w3387 = v1227;
assign w3388 = w2140 & w2460;
assign w3389 = ~pi366 & pi193;
assign w3390 = ~w286 & w2573;
assign v1228 = ~(w2656 | w3852);
assign w3391 = v1228;
assign w3392 = w3601 & w202;
assign w3393 = w3559 & w2302;
assign w3394 = ~w3094 & w2664;
assign v1229 = ~(w425 | w1061);
assign w3395 = v1229;
assign v1230 = ~(w125 | w670);
assign w3396 = v1230;
assign w3397 = w3541 & w1469;
assign v1231 = ~(w2050 | w898);
assign w3398 = v1231;
assign w3399 = w3094 & w1894;
assign w3400 = w1199 & ~w3049;
assign w3401 = ~w834 & w56;
assign w3402 = w950 & ~w611;
assign w3403 = ~w964 & w227;
assign w3404 = pi258 & w2362;
assign w3405 = (~w354 & w4006) | (~w354 & w3782) | (w4006 & w3782);
assign w3406 = ~w354 & w1219;
assign w3407 = w3200 & ~w1996;
assign v1232 = ~(w1087 | w2607);
assign w3408 = v1232;
assign v1233 = ~(w799 | w1831);
assign w3409 = v1233;
assign w3410 = ~w800 & w3068;
assign w3411 = ~w2215 & w4143;
assign v1234 = ~(w3644 | w1528);
assign w3412 = v1234;
assign v1235 = ~(w3856 | w1662);
assign w3413 = v1235;
assign w3414 = ~w4119 & w4170;
assign v1236 = ~(w3272 | w508);
assign w3415 = v1236;
assign v1237 = ~(w700 | w661);
assign w3416 = v1237;
assign w3417 = ~w3094 & w2310;
assign v1238 = ~(w1754 | w923);
assign w3418 = v1238;
assign w3419 = (~w4035 & w3653) | (~w4035 & w2845) | (w3653 & w2845);
assign v1239 = ~(w999 | w2766);
assign w3420 = v1239;
assign w3421 = (pi032 & ~w1654) | (pi032 & w2385) | (~w1654 & w2385);
assign w3422 = ~w3339 & w3865;
assign w3423 = w2116 & w1242;
assign v1240 = ~(w3905 | w2412);
assign w3424 = v1240;
assign v1241 = ~(w3052 | w4027);
assign w3425 = v1241;
assign w3426 = ~w350 & w4139;
assign w3427 = ~w3094 & w1805;
assign w3428 = ~pi366 & pi240;
assign w3429 = (w4035 & w2883) | (w4035 & w1414) | (w2883 & w1414);
assign w3430 = w3094 & w742;
assign v1242 = ~(w634 | w1392);
assign w3431 = v1242;
assign w3432 = (pi041 & ~w1654) | (pi041 & w2410) | (~w1654 & w2410);
assign v1243 = ~(w1452 | w1478);
assign w3433 = v1243;
assign v1244 = ~(w4159 | w1899);
assign w3434 = v1244;
assign w3435 = w78 & w1469;
assign w3436 = (w203 & ~w61) | (w203 & w3660) | (~w61 & w3660);
assign w3437 = w3094 & w2400;
assign w3438 = w4015 & ~w1789;
assign w3439 = w269 & ~w2099;
assign v1245 = ~(w2406 | w3612);
assign w3440 = v1245;
assign w3441 = w3882 & ~w991;
assign w3442 = (w3706 & ~w3239) | (w3706 & w4110) | (~w3239 & w4110);
assign w3443 = w2046 & ~w435;
assign w3444 = w1570 & w2702;
assign w3445 = pi298 & w2362;
assign v1246 = ~(w4057 | w2842);
assign w3446 = v1246;
assign v1247 = ~(w1993 | w4019);
assign w3447 = v1247;
assign w3448 = (w15 & w2298) | (w15 & w1817) | (w2298 & w1817);
assign w3449 = w3961 & w1125;
assign v1248 = ~(w1084 | w4142);
assign w3450 = v1248;
assign v1249 = ~(w3499 | w1433);
assign w3451 = v1249;
assign v1250 = ~(w954 | w3977);
assign w3452 = v1250;
assign w3453 = w308 & w1249;
assign w3454 = w3273 & ~w1166;
assign v1251 = ~(w3160 | w557);
assign w3455 = v1251;
assign v1252 = ~(w1434 | w2792);
assign w3456 = v1252;
assign v1253 = ~(w2502 | w2295);
assign w3457 = v1253;
assign w3458 = pi322 & ~pi366;
assign w3459 = w517 & w469;
assign w3460 = w118 & pi089;
assign w3461 = w118 & pi095;
assign w3462 = ~w3541 & w2433;
assign w3463 = (~w227 & ~w63) | (~w227 & w2978) | (~w63 & w2978);
assign v1254 = ~(w2874 | w1661);
assign w3464 = v1254;
assign w3465 = w118 & pi005;
assign w3466 = (w1469 & ~w1704) | (w1469 & w2134) | (~w1704 & w2134);
assign w3467 = w2140 & ~w2022;
assign w3468 = w3333 & w1543;
assign w3469 = w672 & ~w2894;
assign w3470 = (w1469 & ~w4157) | (w1469 & w3526) | (~w4157 & w3526);
assign w3471 = w2598 & w1654;
assign v1255 = ~(w3763 | w1424);
assign w3472 = v1255;
assign w3473 = w2759 & ~w1469;
assign w3474 = w3077 & w1163;
assign w3475 = w656 & ~w498;
assign v1256 = ~(w179 | w3905);
assign w3476 = v1256;
assign w3477 = (~w1469 & ~w4170) | (~w1469 & w1536) | (~w4170 & w1536);
assign w3478 = (pi073 & ~w1654) | (pi073 & w1763) | (~w1654 & w1763);
assign v1257 = ~(w3927 | w3011);
assign w3479 = v1257;
assign w3480 = ~pi366 & pi229;
assign w3481 = w3778 & w581;
assign w3482 = w1580 & w233;
assign w3483 = ~w1139 & w3188;
assign w3484 = w1830 & ~w3317;
assign w3485 = w2479 & ~w361;
assign v1258 = ~(w1139 | w24);
assign w3486 = v1258;
assign w3487 = w1182 & ~w844;
assign w3488 = (w3180 & w3531) | (w3180 & w2635) | (w3531 & w2635);
assign v1259 = ~(w3381 | w3301);
assign w3489 = v1259;
assign w3490 = (pi047 & ~w1654) | (pi047 & w90) | (~w1654 & w90);
assign w3491 = pi359 & ~pi366;
assign v1260 = ~(w1364 | w1816);
assign w3492 = v1260;
assign w3493 = w378 & ~w1777;
assign w3494 = w2606 & ~w342;
assign w3495 = w2893 & ~w991;
assign w3496 = w3216 & ~w1774;
assign v1261 = ~(w3025 | w2095);
assign w3497 = v1261;
assign v1262 = ~(w2097 | w1210);
assign w3498 = v1262;
assign v1263 = ~(w3878 | w398);
assign w3499 = v1263;
assign w3500 = (~w430 & ~w1649) | (~w430 & w3369) | (~w1649 & w3369);
assign v1264 = ~(w3648 | w248);
assign w3501 = v1264;
assign w3502 = pi037 & w570;
assign w3503 = ~w1573 & w1566;
assign w3504 = pi155 & w1570;
assign v1265 = ~(w1318 | w3159);
assign w3505 = v1265;
assign v1266 = ~(w1754 | w1533);
assign w3506 = v1266;
assign w3507 = w3531 & w254;
assign w3508 = pi249 & w2362;
assign w3509 = ~w3094 & w3088;
assign w3510 = (w2690 & w1849) | (w2690 & w3078) | (w1849 & w3078);
assign v1267 = ~(w2729 | w934);
assign w3511 = v1267;
assign v1268 = ~(w2431 | w4088);
assign w3512 = v1268;
assign v1269 = ~(w1523 | w3);
assign w3513 = v1269;
assign v1270 = ~(w3271 | w2401);
assign w3514 = v1270;
assign v1271 = ~(w3878 | w2412);
assign w3515 = v1271;
assign w3516 = w2717 & ~w448;
assign w3517 = w52 & w1654;
assign v1272 = ~(w1159 | w1775);
assign w3518 = v1272;
assign w3519 = ~pi366 & pi214;
assign w3520 = pi353 & ~pi366;
assign w3521 = w3669 & ~w1682;
assign w3522 = (~w442 & ~w3883) | (~w442 & w3213) | (~w3883 & w3213);
assign w3523 = w1246 & ~w1469;
assign w3524 = (w1653 & ~w1338) | (w1653 & w1316) | (~w1338 & w1316);
assign w3525 = w1772 & ~w1469;
assign w3526 = w2732 & w1469;
assign w3527 = w2890 & w3110;
assign v1273 = ~(w259 | w279);
assign w3528 = v1273;
assign w3529 = pi021 & w570;
assign v1274 = ~(w1754 | w2955);
assign w3530 = v1274;
assign w3531 = ~w800 & w2936;
assign w3532 = w760 & w2119;
assign w3533 = pi169 & ~pi364;
assign v1275 = ~(w1089 | w3022);
assign w3534 = v1275;
assign w3535 = w27 & w596;
assign w3536 = ~w263 & w2245;
assign w3537 = w2596 & w2440;
assign w3538 = w3591 & w4032;
assign v1276 = ~(w1754 | w3105);
assign w3539 = v1276;
assign w3540 = pi107 & w570;
assign w3541 = ~w3094 & w525;
assign w3542 = w226 & ~w3191;
assign w3543 = ~w614 & w2071;
assign w3544 = pi086 & w353;
assign v1277 = ~(w2799 | w3848);
assign w3545 = v1277;
assign v1278 = ~(w980 | w516);
assign w3546 = v1278;
assign w3547 = pi362 & pi363;
assign w3548 = w2954 & w1178;
assign w3549 = w1815 & w1887;
assign w3550 = w118 & pi001;
assign v1279 = ~(w486 | w2956);
assign w3551 = v1279;
assign w3552 = ~w4138 & w846;
assign w3553 = w443 & w3015;
assign v1280 = ~(w889 | w3894);
assign w3554 = v1280;
assign v1281 = ~(w3160 | w3848);
assign w3555 = v1281;
assign w3556 = w546 & ~w1469;
assign w3557 = w2345 & ~w772;
assign w3558 = ~w1454 & w2989;
assign v1282 = ~(w2468 | w75);
assign w3559 = v1282;
assign v1283 = ~(w4038 | w1533);
assign w3560 = v1283;
assign w3561 = w118 & pi115;
assign w3562 = w1700 & ~w1698;
assign w3563 = w1830 & ~w1881;
assign w3564 = w3945 & ~w1469;
assign v1284 = ~(w2905 | w708);
assign w3565 = v1284;
assign v1285 = ~(w3160 | w398);
assign w3566 = v1285;
assign w3567 = w3624 & w1654;
assign w3568 = ~w2419 & w3835;
assign w3569 = (~w3191 & ~w3813) | (~w3191 & w2021) | (~w3813 & w2021);
assign v1286 = ~(w2784 | w1449);
assign w3570 = v1286;
assign w3571 = (w442 & w2487) | (w442 & w1331) | (w2487 & w1331);
assign w3572 = w1570 & w467;
assign v1287 = ~(w486 | w2486);
assign w3573 = v1287;
assign v1288 = ~(w4104 | w1374);
assign w3574 = v1288;
assign v1289 = ~(w2646 | w3180);
assign w3575 = v1289;
assign w3576 = w2717 & ~w4105;
assign w3577 = w713 & w3574;
assign v1290 = ~(w2799 | w1881);
assign w3578 = v1290;
assign w3579 = w705 & w4061;
assign w3580 = pi345 & ~pi366;
assign v1291 = ~(w2650 | w1824);
assign w3581 = v1291;
assign v1292 = ~(w2244 | w1644);
assign w3582 = v1292;
assign w3583 = w2655 & w4152;
assign w3584 = pi266 & w2362;
assign w3585 = ~w2024 & w3633;
assign w3586 = ~w1369 & w421;
assign w3587 = ~w429 & w3562;
assign w3588 = w2140 & w2022;
assign v1293 = ~(w1470 | w3850);
assign w3589 = v1293;
assign v1294 = ~(w1906 | w563);
assign w3590 = v1294;
assign v1295 = ~(w311 | w1298);
assign w3591 = v1295;
assign v1296 = ~(w4176 | w2657);
assign w3592 = v1296;
assign w3593 = (~w46 & w4114) | (~w46 & w1359) | (w4114 & w1359);
assign w3594 = ~w3647 & w1049;
assign v1297 = ~(w4038 | w2209);
assign w3595 = v1297;
assign w3596 = w3334 & w1469;
assign w3597 = (w1182 & w572) | (w1182 & w3217) | (w572 & w3217);
assign w3598 = w672 & ~w3241;
assign v1298 = ~(w2269 | w3959);
assign w3599 = v1298;
assign w3600 = pi294 & w2362;
assign v1299 = ~(w354 | w1219);
assign w3601 = v1299;
assign w3602 = w118 & pi092;
assign w3603 = (w2765 & w2846) | (w2765 & w2593) | (w2846 & w2593);
assign v1300 = ~(w2926 | w1063);
assign w3604 = v1300;
assign v1301 = ~(w2905 | w3716);
assign w3605 = v1301;
assign w3606 = w927 & w3212;
assign w3607 = ~w2461 & w2484;
assign w3608 = w3094 & w1833;
assign v1302 = ~(w794 | w2475);
assign w3609 = v1302;
assign w3610 = w656 & ~w557;
assign v1303 = ~(w3702 | w3947);
assign w3611 = v1303;
assign w3612 = pi262 & w2362;
assign w3613 = w672 & ~w3007;
assign w3614 = w1112 & w2608;
assign w3615 = pi080 & w353;
assign w3616 = w407 & w1190;
assign w3617 = w3337 & w1654;
assign w3618 = w3417 & w1075;
assign w3619 = w1918 & w2451;
assign w3620 = w2902 & w2113;
assign w3621 = w1830 & ~w4105;
assign w3622 = w3606 & w1601;
assign v1304 = ~(w3216 | w2942);
assign w3623 = v1304;
assign w3624 = pi176 & w1570;
assign w3625 = ~w1126 & w4013;
assign v1305 = ~(w1038 | w2360);
assign w3626 = v1305;
assign v1306 = ~(w2874 | w3878);
assign w3627 = v1306;
assign v1307 = ~(w1191 | w869);
assign w3628 = v1307;
assign w3629 = w2626 & ~w1393;
assign w3630 = w3062 & w1273;
assign w3631 = pi051 & w570;
assign w3632 = w118 & pi122;
assign v1308 = ~(w2985 | w160);
assign w3633 = v1308;
assign w3634 = w3938 & w2547;
assign w3635 = w2046 & w1762;
assign w3636 = pi343 & ~pi366;
assign v1309 = ~(w4159 | w3943);
assign w3637 = v1309;
assign w3638 = (pi024 & ~w1654) | (pi024 & w282) | (~w1654 & w282);
assign w3639 = w2065 & w2026;
assign w3640 = w3684 & w4036;
assign w3641 = pi012 & w570;
assign w3642 = ~pi366 & pi208;
assign w3643 = w656 & ~w3343;
assign w3644 = (w1469 & ~w1748) | (w1469 & w116) | (~w1748 & w116);
assign w3645 = ~w425 & w771;
assign w3646 = w3710 & ~w3669;
assign w3647 = w3486 & ~w454;
assign w3648 = ~w3538 & w3666;
assign w3649 = ~w2356 & w3191;
assign w3650 = w3164 & w3036;
assign w3651 = w118 & pi011;
assign w3652 = pi291 & w2362;
assign w3653 = (~w2993 & w2651) | (~w2993 & w399) | (w2651 & w399);
assign w3654 = ~w2893 & w2280;
assign w3655 = w2340 & w2826;
assign w3656 = w3172 & w3511;
assign v1310 = ~(w2123 | w3259);
assign w3657 = v1310;
assign w3658 = ~w2489 & w1315;
assign w3659 = ~w800 & w244;
assign w3660 = (w203 & ~w683) | (w203 & w2703) | (~w683 & w2703);
assign v1311 = ~(w2721 | w4028);
assign w3661 = v1311;
assign v1312 = ~(w573 | w3578);
assign w3662 = v1312;
assign v1313 = ~(w954 | w2874);
assign w3663 = v1313;
assign w3664 = w4178 & w1172;
assign w3665 = w3159 & w361;
assign w3666 = ~w1800 & w1926;
assign w3667 = w2936 & w3799;
assign w3668 = w2247 & w1469;
assign w3669 = w3547 & w1273;
assign v1314 = ~(w154 | w2577);
assign w3670 = v1314;
assign w3671 = (~pi118 & ~w1654) | (~pi118 & w3368) | (~w1654 & w3368);
assign w3672 = w4164 & w1654;
assign v1315 = ~(w2149 | w3163);
assign w3673 = v1315;
assign v1316 = ~(w3432 | w1339);
assign w3674 = v1316;
assign w3675 = ~w811 & w3019;
assign w3676 = w2774 & w2022;
assign w3677 = pi366 & w561;
assign v1317 = ~(w1754 | w3168);
assign w3678 = v1317;
assign v1318 = ~(w1695 | w424);
assign w3679 = v1318;
assign w3680 = (~w1539 & w181) | (~w1539 & ~w736) | (w181 & ~w736);
assign w3681 = w2359 & w1469;
assign v1319 = ~(w2475 | w3858);
assign w3682 = v1319;
assign v1320 = ~(w4040 | w3820);
assign w3683 = v1320;
assign v1321 = ~(w262 | w3033);
assign w3684 = v1321;
assign v1322 = ~(w2799 | w2874);
assign w3685 = v1322;
assign w3686 = pi125 & w353;
assign v1323 = ~(w1467 | w416);
assign w3687 = v1323;
assign v1324 = ~(w4038 | w794);
assign w3688 = v1324;
assign v1325 = ~(w3938 | w2547);
assign w3689 = v1325;
assign w3690 = w141 & w964;
assign v1326 = ~(w2175 | w1164);
assign w3691 = v1326;
assign w3692 = w2717 & ~w1592;
assign w3693 = w1830 & ~w2955;
assign w3694 = w2484 & w138;
assign v1327 = ~(w3312 | w2955);
assign w3695 = v1327;
assign w3696 = (w1469 & ~w1896) | (w1469 & w1951) | (~w1896 & w1951);
assign v1328 = ~(w1604 | w2475);
assign w3697 = v1328;
assign w3698 = w3125 & w1654;
assign w3699 = w110 & w1615;
assign w3700 = w2717 & ~w2123;
assign v1329 = ~(w3365 | w2582);
assign w3701 = v1329;
assign w3702 = w3094 & w1235;
assign v1330 = ~(w25 | w3120);
assign w3703 = v1330;
assign w3704 = w2414 & w1908;
assign w3705 = w2347 & w3701;
assign w3706 = ~w2279 & w1738;
assign w3707 = (pi097 & ~w1654) | (pi097 & w1862) | (~w1654 & w1862);
assign v1331 = ~(w3707 | w1016);
assign w3708 = v1331;
assign w3709 = w656 & ~w920;
assign w3710 = (pi059 & ~w1654) | (pi059 & w1940) | (~w1654 & w1940);
assign w3711 = ~w286 & w361;
assign v1332 = ~(w617 | w804);
assign w3712 = v1332;
assign w3713 = ~w964 & w294;
assign w3714 = w3134 & w854;
assign w3715 = w2936 & w58;
assign w3716 = (w1469 & ~w1121) | (w1469 & w161) | (~w1121 & w161);
assign v1333 = ~(w954 | w498);
assign w3717 = v1333;
assign w3718 = ~w1288 & w1959;
assign v1334 = ~(w3259 | w1881);
assign w3719 = v1334;
assign v1335 = ~(w190 | w1020);
assign w3720 = v1335;
assign w3721 = w351 & w1209;
assign w3722 = ~w1880 & w3201;
assign w3723 = ~w3273 & w1166;
assign v1336 = ~(w226 | w1219);
assign w3724 = v1336;
assign v1337 = ~(w3160 | w1667);
assign w3725 = v1337;
assign w3726 = w1654 & ~w193;
assign w3727 = ~w2268 & w3856;
assign v1338 = ~(w1284 | w604);
assign w3728 = v1338;
assign v1339 = ~(w1998 | w1994);
assign w3729 = v1339;
assign w3730 = pi182 & w1570;
assign v1340 = ~(w2435 | w1003);
assign w3731 = v1340;
assign w3732 = w1214 & w3023;
assign w3733 = ~w2523 & w2487;
assign w3734 = w3094 & w1497;
assign w3735 = w2544 & w502;
assign v1341 = ~(w4159 | w1164);
assign w3736 = v1341;
assign v1342 = ~(w3009 | w2262);
assign w3737 = v1342;
assign w3738 = (~w2487 & ~w834) | (~w2487 & w3035) | (~w834 & w3035);
assign v1343 = ~(w2316 | w896);
assign w3739 = v1343;
assign w3740 = ~w3094 & w2255;
assign v1344 = ~(w1219 | w758);
assign w3741 = v1344;
assign w3742 = w2641 & w1158;
assign w3743 = w4015 & ~w3554;
assign v1345 = ~(w1516 | w1211);
assign w3744 = v1345;
assign w3745 = w3200 & ~w480;
assign w3746 = ~w3277 & w656;
assign w3747 = (w3159 & ~w1103) | (w3159 & w241) | (~w1103 & w241);
assign w3748 = w1516 & w1199;
assign w3749 = w1295 & w2497;
assign v1346 = ~(w1496 | w842);
assign w3750 = v1346;
assign v1347 = ~(w2799 | w3168);
assign w3751 = v1347;
assign w3752 = (~w1403 & w360) | (~w1403 & w1173) | (w360 & w1173);
assign v1348 = ~(w2123 | w3160);
assign w3753 = v1348;
assign w3754 = w2968 & w1425;
assign v1349 = ~(w2348 | w3944);
assign w3755 = v1349;
assign w3756 = (~w1853 & w2896) | (~w1853 & w959) | (w2896 & w959);
assign w3757 = w3083 & w685;
assign w3758 = w1347 & w1654;
assign v1350 = ~(w3159 | w361);
assign w3759 = v1350;
assign w3760 = ~w2411 & w1149;
assign v1351 = ~(w1104 | w1970);
assign w3761 = v1351;
assign w3762 = w1830 & ~w3722;
assign w3763 = w656 & ~w3263;
assign v1352 = ~(w2428 | w1626);
assign w3764 = v1352;
assign v1353 = ~(w1788 | w3381);
assign w3765 = v1353;
assign w3766 = w1076 & ~w863;
assign w3767 = (w3269 & ~w3290) | (w3269 & w2275) | (~w3290 & w2275);
assign v1354 = ~(w1754 | w3385);
assign w3768 = v1354;
assign w3769 = ~w354 & w2466;
assign w3770 = w1938 & w1266;
assign w3771 = (pi095 & ~w1654) | (pi095 & w3461) | (~w1654 & w3461);
assign v1355 = ~(w2874 | w3905);
assign w3772 = v1355;
assign w3773 = ~w680 & w4077;
assign v1356 = ~(w3878 | w1782);
assign w3774 = v1356;
assign w3775 = ~w3094 & w4054;
assign v1357 = ~(w1140 | w3905);
assign w3776 = v1357;
assign w3777 = pi330 & ~pi366;
assign v1358 = ~(w367 | w796);
assign w3778 = v1358;
assign w3779 = w1654 & ~w3744;
assign w3780 = w379 & w915;
assign v1359 = ~(w3906 | w3214);
assign w3781 = v1359;
assign w3782 = w1629 & w1142;
assign v1360 = ~(w2905 | w276);
assign w3783 = v1360;
assign w3784 = w3486 & ~w2815;
assign w3785 = ~w2086 & w2914;
assign v1361 = ~(w1754 | w3858);
assign w3786 = v1361;
assign v1362 = ~(w3921 | w3052);
assign w3787 = v1362;
assign v1363 = ~(w2175 | w448);
assign w3788 = v1363;
assign w3789 = ~pi366 & pi205;
assign v1364 = ~(w1286 | w2736);
assign w3790 = v1364;
assign w3791 = w437 & w3450;
assign w3792 = (w1469 & ~w2407) | (w1469 & w3195) | (~w2407 & w3195);
assign w3793 = ~w4073 & w2626;
assign w3794 = w3805 & w2977;
assign w3795 = w2397 & ~w3744;
assign v1365 = ~(w1577 | w2107);
assign w3796 = v1365;
assign v1366 = ~(w3160 | w542);
assign w3797 = v1366;
assign v1367 = ~(w3160 | w1633);
assign w3798 = v1367;
assign w3799 = w800 & w244;
assign v1368 = ~(w138 | w2461);
assign w3800 = v1368;
assign w3801 = pi130 & w1570;
assign w3802 = (~w2179 & w811) | (~w2179 & w1710) | (w811 & w1710);
assign v1369 = ~(w1567 | w2921);
assign w3803 = v1369;
assign v1370 = ~(w3476 | w2652);
assign w3804 = v1370;
assign w3805 = w537 & w944;
assign v1371 = ~(w1970 | w3943);
assign w3806 = v1371;
assign w3807 = w2157 & w1639;
assign w3808 = ~w3094 & w274;
assign v1372 = ~(w314 | w623);
assign w3809 = v1372;
assign w3810 = w3140 & w795;
assign w3811 = ~w2351 & w155;
assign w3812 = (w3467 & ~w2234) | (w3467 & w224) | (~w2234 & w224);
assign v1373 = ~(w1219 | w1301);
assign w3813 = v1373;
assign v1374 = ~(w3312 | w1444);
assign w3814 = v1374;
assign w3815 = ~pi366 & pi204;
assign w3816 = w3790 & w822;
assign w3817 = (~w1469 & ~w74) | (~w1469 & w982) | (~w74 & w982);
assign w3818 = pi029 & w570;
assign w3819 = w660 & w187;
assign w3820 = (pi096 & ~w1654) | (pi096 & w1234) | (~w1654 & w1234);
assign w3821 = w851 & ~w4074;
assign v1375 = ~(w15 | w4065);
assign w3822 = v1375;
assign w3823 = (~w1469 & ~w3673) | (~w1469 & w692) | (~w3673 & w692);
assign w3824 = w3109 & w3173;
assign w3825 = w2484 & ~w4065;
assign v1376 = ~(w3897 | w3682);
assign w3826 = v1376;
assign w3827 = w46 & ~w3496;
assign w3828 = ~w1576 & w861;
assign w3829 = w1776 & w1034;
assign w3830 = w3738 & ~w3619;
assign w3831 = w1294 & w1654;
assign v1377 = ~(w2123 | w4159);
assign w3832 = v1377;
assign w3833 = w3731 & w3809;
assign w3834 = w4011 & w881;
assign v1378 = ~(w638 | w576);
assign w3835 = v1378;
assign v1379 = ~(w954 | w3848);
assign w3836 = v1379;
assign w3837 = w3094 & w526;
assign v1380 = ~(w313 | w129);
assign w3838 = v1380;
assign v1381 = ~(w1503 | w1646);
assign w3839 = v1381;
assign v1382 = ~(w2475 | w923);
assign w3840 = v1382;
assign w3841 = (~w3781 & w2665) | (~w3781 & w2235) | (w2665 & w2235);
assign w3842 = (w1654 & w1521) | (w1654 & w1439) | (w1521 & w1439);
assign v1383 = ~(w1463 | w579);
assign w3843 = v1383;
assign w3844 = ~w3654 & w612;
assign w3845 = ~pi366 & pi201;
assign w3846 = w992 & w1152;
assign w3847 = (w1654 & w783) | (w1654 & w3831) | (w783 & w3831);
assign w3848 = ~w725 & w74;
assign w3849 = w2717 & ~w3343;
assign w3850 = w2315 & w3690;
assign v1384 = ~(w4159 | w448);
assign w3851 = v1384;
assign w3852 = (pi122 & ~w1654) | (pi122 & w3632) | (~w1654 & w3632);
assign w3853 = w3740 & w1469;
assign w3854 = ~w3934 & w3338;
assign w3855 = w3094 & w2236;
assign w3856 = w2324 & w4047;
assign w3857 = w656 & ~w357;
assign w3858 = ~w2578 & w2613;
assign w3859 = w2822 & ~w1082;
assign v1385 = ~(w2175 | w920);
assign w3860 = v1385;
assign v1386 = ~(w2475 | w1164);
assign w3861 = v1386;
assign v1387 = ~(w2442 | w3310);
assign w3862 = v1387;
assign v1388 = ~(w2644 | w1056);
assign w3863 = v1388;
assign v1389 = ~(w3075 | w84);
assign w3864 = v1389;
assign v1390 = ~(w759 | w3165);
assign w3865 = v1390;
assign w3866 = (w2397 & w1849) | (w2397 & w2354) | (w1849 & w2354);
assign w3867 = w1031 & w3592;
assign v1391 = ~(w938 | w2252);
assign w3868 = v1391;
assign v1392 = ~(w271 | w376);
assign w3869 = v1392;
assign w3870 = ~w3552 & w2595;
assign v1393 = ~(w1754 | w498);
assign w3871 = v1393;
assign w3872 = w3094 & w1606;
assign w3873 = ~pi366 & pi243;
assign v1394 = ~(w3929 | w3160);
assign w3874 = v1394;
assign w3875 = ~w1189 & w464;
assign w3876 = pi317 & ~pi366;
assign w3877 = w3094 & w3311;
assign v1395 = ~(w955 | w1018);
assign w3878 = v1395;
assign v1396 = ~(w1683 | w2695);
assign w3879 = v1396;
assign v1397 = ~(w3603 | w1124);
assign w3880 = v1397;
assign w3881 = w2443 & ~w655;
assign v1398 = ~(w2893 | w4047);
assign w3882 = v1398;
assign w3883 = ~w2374 & w1626;
assign v1399 = ~(w3160 | w2955);
assign w3884 = v1399;
assign w3885 = pi084 & w570;
assign w3886 = (~w1507 & ~w3645) | (~w1507 & w167) | (~w3645 & w167);
assign w3887 = ~w4051 & w8;
assign w3888 = w2728 & ~w2145;
assign w3889 = w898 & ~w610;
assign w3890 = w805 & w1469;
assign v1400 = ~(w1661 | w1444);
assign w3891 = v1400;
assign w3892 = pi274 & w2362;
assign w3893 = pi303 & w2362;
assign w3894 = (w1469 & ~w3319) | (w1469 & w3596) | (~w3319 & w3596);
assign w3895 = pi010 & w570;
assign v1401 = ~(w3259 | w3131);
assign w3896 = v1401;
assign v1402 = ~(w3160 | w1955);
assign w3897 = v1402;
assign w3898 = w1469 & w672;
assign v1403 = ~(w1754 | w3414);
assign w3899 = v1403;
assign w3900 = ~w2070 & w500;
assign w3901 = ~w3870 & w3060;
assign w3902 = ~w2932 & w1653;
assign w3903 = w3128 & ~w2484;
assign v1404 = ~(w2158 | w3045);
assign w3904 = v1404;
assign v1405 = ~(w2787 | w3811);
assign w3905 = v1405;
assign v1406 = ~(w826 | w96);
assign w3906 = v1406;
assign v1407 = ~(w1607 | w2175);
assign w3907 = v1407;
assign w3908 = w3094 & w2220;
assign w3909 = w118 & pi090;
assign w3910 = (pi019 & ~w1654) | (pi019 & w2472) | (~w1654 & w2472);
assign w3911 = w705 & w3130;
assign v1408 = ~(w1461 | w3762);
assign w3912 = v1408;
assign w3913 = ~w1344 & w195;
assign w3914 = w3253 & ~w3706;
assign w3915 = w4074 & ~w973;
assign v1409 = ~(w2033 | w2753);
assign w3916 = v1409;
assign w3917 = ~w1933 & w50;
assign v1410 = ~(w2755 | w3579);
assign w3918 = v1410;
assign w3919 = ~w2492 & w637;
assign v1411 = ~(w48 | w4038);
assign w3920 = v1411;
assign w3921 = (w1469 & ~w251) | (w1469 & w245) | (~w251 & w245);
assign w3922 = w1067 & w1975;
assign w3923 = w2443 & ~w2494;
assign w3924 = w3094 & w3314;
assign v1412 = ~(w1599 | w100);
assign w3925 = v1412;
assign v1413 = ~(w2105 | w3990);
assign w3926 = v1413;
assign w3927 = (pi088 & ~w1654) | (pi088 & w3359) | (~w1654 & w3359);
assign w3928 = ~w3094 & w3122;
assign w3929 = ~w484 & w522;
assign v1414 = ~(w1661 | w2955);
assign w3930 = v1414;
assign w3931 = ~w2341 & w673;
assign w3932 = (~w1469 & ~w1217) | (~w1469 & w1430) | (~w1217 & w1430);
assign w3933 = w1182 & ~w924;
assign w3934 = w2460 & w3467;
assign w3935 = w342 & w187;
assign v1415 = ~(w3287 | w1996);
assign w3936 = v1415;
assign w3937 = w1570 & w2532;
assign w3938 = ~w3420 & w1401;
assign w3939 = ~pi366 & pi231;
assign w3940 = ~w3199 & w2324;
assign v1416 = ~(w81 | w1221);
assign w3941 = v1416;
assign v1417 = ~(w3905 | w3343);
assign w3942 = v1417;
assign w3943 = ~w3427 & w3570;
assign v1418 = ~(w2799 | w1955);
assign w3944 = v1418;
assign w3945 = ~w3094 & w3873;
assign v1419 = ~(w4159 | w357);
assign w3946 = v1419;
assign w3947 = pi296 & w2362;
assign w3948 = w3998 & ~w2500;
assign w3949 = (w1934 & w1814) | (w1934 & w2176) | (w1814 & w2176);
assign w3950 = ~w3098 & w2715;
assign v1420 = ~(w106 | w3135);
assign w3951 = v1420;
assign w3952 = ~w913 & w3931;
assign w3953 = w378 & ~w3194;
assign w3954 = ~w4074 & w973;
assign w3955 = pi270 & w2362;
assign w3956 = w1080 & ~w2950;
assign w3957 = w3799 & w714;
assign w3958 = w1292 & w1469;
assign w3959 = ~w3391 & w3841;
assign w3960 = ~w1004 & w3091;
assign v1421 = ~(w140 | w3697);
assign w3961 = v1421;
assign w3962 = pi079 & w353;
assign w3963 = pi360 & pi367;
assign w3964 = ~w3417 & w2369;
assign w3965 = w118 & pi094;
assign w3966 = w705 & w3572;
assign v1422 = ~(w338 | w3487);
assign w3967 = v1422;
assign w3968 = w4053 & ~w1469;
assign w3969 = ~w440 & w2023;
assign v1423 = ~(w2475 | w920);
assign w3970 = v1423;
assign w3971 = w4 & w2397;
assign w3972 = w4017 & ~w3773;
assign w3973 = ~w4185 & w3940;
assign w3974 = (w3068 & w2666) | (w3068 & w2526) | (w2666 & w2526);
assign w3975 = w419 & ~w3380;
assign v1424 = ~(w3160 | w149);
assign w3976 = v1424;
assign w3977 = ~w668 & w2254;
assign w3978 = w118 & pi009;
assign w3979 = (w2631 & ~w1308) | (w2631 & w1283) | (~w1308 & w1283);
assign w3980 = w15 & ~w2484;
assign w3981 = (w2094 & ~w2530) | (w2094 & w1427) | (~w2530 & w1427);
assign v1425 = ~(w3691 | w2887);
assign w3982 = v1425;
assign w3983 = ~w1469 & w1199;
assign w3984 = ~w3999 & w545;
assign w3985 = (w2968 & ~w1303) | (w2968 & w1897) | (~w1303 & w1897);
assign w3986 = ~w2528 & w2539;
assign v1426 = ~(w3866 | w1968);
assign w3987 = v1426;
assign w3988 = w2424 & w3443;
assign w3989 = w1440 & w702;
assign w3990 = w3950 & w1522;
assign w3991 = w972 & w1654;
assign w3992 = w2127 & w1044;
assign v1427 = ~(w4027 | w1528);
assign w3993 = v1427;
assign v1428 = ~(w3107 | w903);
assign w3994 = v1428;
assign w3995 = w2181 & w2698;
assign w3996 = ~w3998 & w2500;
assign w3997 = ~w2519 & w3085;
assign v1429 = ~(w2780 | w963);
assign w3998 = v1429;
assign w3999 = w1391 & w3022;
assign v1430 = ~(pi364 | pi365);
assign w4000 = v1430;
assign w4001 = w2917 & w295;
assign w4002 = ~pi050 & w570;
assign v1431 = ~(w179 | w2175);
assign w4003 = v1431;
assign w4004 = w1089 & ~w294;
assign v1432 = ~(w3768 | w1724);
assign w4005 = v1432;
assign v1433 = ~(w2967 | w2589);
assign w4006 = v1433;
assign w4007 = w2690 & ~w2745;
assign w4008 = ~w3140 & w294;
assign w4009 = (w3422 & ~w3248) | (w3422 & w3184) | (~w3248 & w3184);
assign v1434 = ~(w2958 | w3411);
assign w4010 = v1434;
assign w4011 = w769 & w607;
assign w4012 = (w1891 & w3980) | (w1891 & w2224) | (w3980 & w2224);
assign v1435 = ~(w54 | w3819);
assign w4013 = v1435;
assign v1436 = ~(w671 | w2402);
assign w4014 = v1436;
assign w4015 = w2357 & w930;
assign v1437 = ~(w4038 | w3317);
assign w4016 = v1437;
assign w4017 = w1410 & w10;
assign v1438 = ~(w115 | w1281);
assign w4018 = v1438;
assign w4019 = w1182 & ~w2081;
assign w4020 = pi139 & w1570;
assign w4021 = w1451 & ~w3238;
assign v1439 = ~(w1970 | w1533);
assign w4022 = v1439;
assign v1440 = ~(w3259 | w1533);
assign w4023 = v1440;
assign w4024 = w3132 & w2940;
assign v1441 = ~(w1754 | w1955);
assign w4025 = v1441;
assign w4026 = w118 & pi087;
assign w4027 = (w1469 & ~w1356) | (w1469 & w3435) | (~w1356 & w3435);
assign w4028 = w2717 & ~w398;
assign w4029 = ~w569 & w1491;
assign v1442 = ~(w2416 | w3047);
assign w4030 = v1442;
assign w4031 = w2673 & w512;
assign w4032 = ~w339 & w2552;
assign w4033 = w1903 & w3449;
assign w4034 = w2717 & ~w3462;
assign w4035 = ~w1848 & w2995;
assign v1443 = ~(w1558 | w594);
assign w4036 = v1443;
assign w4037 = w2083 & ~w2724;
assign v1444 = ~(w2764 | w659);
assign w4038 = v1444;
assign w4039 = ~w2280 & w4160;
assign w4040 = (w1654 & w2541) | (w1654 & w1666) | (w2541 & w1666);
assign v1445 = ~(w1118 | w3147);
assign w4041 = v1445;
assign v1446 = ~(w37 | w3587);
assign w4042 = v1446;
assign w4043 = ~pi360 & pi366;
assign w4044 = w1600 & w1469;
assign w4045 = ~w3813 & w2073;
assign w4046 = w1123 & w20;
assign v1447 = ~(w300 | w363);
assign w4047 = v1447;
assign w4048 = w964 & ~w227;
assign w4049 = w3061 & ~w183;
assign v1448 = ~(w954 | w1444);
assign w4050 = v1448;
assign w4051 = pi114 & w353;
assign w4052 = (w1654 & w3181) | (w1654 & w2253) | (w3181 & w2253);
assign w4053 = ~w3094 & w4163;
assign w4054 = ~pi366 & pi203;
assign v1449 = ~(w2174 | w1508);
assign w4055 = v1449;
assign w4056 = w2646 & w2082;
assign w4057 = w3630 & ~w598;
assign w4058 = w1570 & w752;
assign w4059 = (w1469 & ~w848) | (w1469 & w88) | (~w848 & w88);
assign v1450 = ~(w1970 | w1782);
assign w4060 = v1450;
assign w4061 = w1570 & w3533;
assign w4062 = pi313 & ~pi366;
assign w4063 = w3509 & w1469;
assign v1451 = ~(w1808 | w3418);
assign w4064 = v1451;
assign v1452 = ~(w3014 | w1701);
assign w4065 = v1452;
assign v1453 = ~(w3179 | w3216);
assign w4066 = v1453;
assign v1454 = ~(w1754 | w1881);
assign w4067 = v1454;
assign w4068 = (pi066 & ~w1654) | (pi066 & w2649) | (~w1654 & w2649);
assign w4069 = w1654 & ~w1469;
assign w4070 = ~w3079 & w2470;
assign v1455 = ~(w354 | w3061);
assign w4071 = v1455;
assign w4072 = (~w46 & w2131) | (~w46 & w2464) | (w2131 & w2464);
assign w4073 = (pi031 & ~w1654) | (pi031 & w588) | (~w1654 & w588);
assign v1456 = ~(w2078 | w329);
assign w4074 = v1456;
assign v1457 = ~(w1961 | w2257);
assign w4075 = v1457;
assign v1458 = ~(w4120 | w1695);
assign w4076 = v1458;
assign v1459 = ~(w2770 | w2155);
assign w4077 = v1459;
assign v1460 = ~(w2175 | w1444);
assign w4078 = v1460;
assign v1461 = ~(w2475 | w1592);
assign w4079 = v1461;
assign v1462 = ~(w954 | w920);
assign w4080 = v1462;
assign w4081 = (pi115 & ~w1654) | (pi115 & w3561) | (~w1654 & w3561);
assign v1463 = ~(w3663 | w3018);
assign w4082 = v1463;
assign w4083 = w1758 & w3068;
assign w4084 = w26 & w1874;
assign v1464 = ~(w4159 | w3977);
assign w4085 = v1464;
assign w4086 = w1570 & w1634;
assign w4087 = ~w2907 & w2434;
assign w4088 = (w2690 & w2168) | (w2690 & w1042) | (w2168 & w1042);
assign w4089 = (pi110 & ~w1654) | (pi110 & w686) | (~w1654 & w686);
assign v1465 = ~(w2343 | w3891);
assign w4090 = v1465;
assign w4091 = w46 & ~w76;
assign v1466 = ~(w1155 | w3695);
assign w4092 = v1466;
assign w4093 = (~w3008 & w2624) | (~w3008 & w231) | (w2624 & w231);
assign v1467 = ~(w1635 | w3188);
assign w4094 = v1467;
assign v1468 = ~(w2691 | w873);
assign w4095 = v1468;
assign v1469 = ~(w3259 | w923);
assign w4096 = v1469;
assign w4097 = ~w2676 & w2730;
assign v1470 = ~(w1368 | w2388);
assign w4098 = v1470;
assign v1471 = ~(w3496 | w3340);
assign w4099 = v1471;
assign v1472 = ~(w2103 | w4168);
assign w4100 = v1472;
assign v1473 = ~(w794 | w2175);
assign w4101 = v1473;
assign v1474 = ~(w536 | w1282);
assign w4102 = v1474;
assign v1475 = ~(w2475 | w498);
assign w4103 = v1475;
assign v1476 = ~(w1754 | w3964);
assign w4104 = v1476;
assign w4105 = ~w388 & w478;
assign v1477 = ~(w3044 | w387);
assign w4106 = v1477;
assign w4107 = w1870 & w1469;
assign v1478 = ~(w480 | w1795);
assign w4108 = v1478;
assign w4109 = w1050 & w2506;
assign w4110 = ~w3253 & w3706;
assign v1479 = ~(w2975 | w3786);
assign w4111 = v1479;
assign w4112 = ~w961 & w4004;
assign v1480 = ~(w3179 | w2497);
assign w4113 = v1480;
assign v1481 = ~(w2628 | w1762);
assign w4114 = v1481;
assign w4115 = w1962 & w2027;
assign w4116 = (w2215 & ~w3535) | (w2215 & w514) | (~w3535 & w514);
assign w4117 = w118 & pi045;
assign w4118 = w2270 & w780;
assign w4119 = ~w3094 & w2187;
assign w4120 = (w1469 & ~w767) | (w1469 & w2063) | (~w767 & w2063);
assign w4121 = w806 & ~w2542;
assign w4122 = ~w2286 & w3557;
assign w4123 = w2140 & w1458;
assign w4124 = w1249 & ~w2150;
assign w4125 = w2676 & ~w2730;
assign v1482 = ~(w275 | w2880);
assign w4126 = v1482;
assign v1483 = ~(w2829 | w1422);
assign w4127 = v1483;
assign v1484 = ~(w2856 | w4136);
assign w4128 = v1484;
assign w4129 = w1570 & w1477;
assign w4130 = ~w1319 & w138;
assign w4131 = ~w2840 & w3721;
assign w4132 = w2480 & w1249;
assign v1485 = ~(w3312 | w1667);
assign w4133 = v1485;
assign w4134 = ~w1080 & w2950;
assign w4135 = pi124 & w353;
assign v1486 = ~(w3312 | w1533);
assign w4136 = v1486;
assign w4137 = w2046 & ~w3216;
assign v1487 = ~(w3159 | w2070);
assign w4138 = v1487;
assign v1488 = ~(w1048 | w1435);
assign w4139 = v1488;
assign w4140 = w2898 & w3856;
assign w4141 = ~pi366 & pi227;
assign w4142 = w1199 & ~w3787;
assign w4143 = w3346 & w2872;
assign w4144 = ~w1492 & w1774;
assign v1489 = ~(w2799 | w920);
assign w4145 = v1489;
assign v1490 = ~(w1970 | w3426);
assign w4146 = v1490;
assign w4147 = pi325 & ~pi366;
assign v1491 = ~(w3929 | w3312);
assign w4148 = v1491;
assign w4149 = w1469 & w1249;
assign w4150 = ~w862 & w3901;
assign w4151 = w2244 & ~w381;
assign v1492 = ~(w2951 | w3539);
assign w4152 = v1492;
assign w4153 = w2003 & w1654;
assign w4154 = w656 & ~w2412;
assign v1493 = ~(w830 | w1988);
assign w4155 = v1493;
assign w4156 = w128 & ~w361;
assign v1494 = ~(w3734 | w2851);
assign w4157 = v1494;
assign w4158 = ~w2891 & w814;
assign v1495 = ~(w3318 | w1890);
assign w4159 = v1495;
assign v1496 = ~(w2606 | w991);
assign w4160 = v1496;
assign v1497 = ~(w1999 | w1407);
assign w4161 = v1497;
assign w4162 = pi255 & w2362;
assign w4163 = ~pi366 & pi233;
assign w4164 = pi177 & w1570;
assign w4165 = w3417 & w1469;
assign v1498 = ~(w1661 | w1899);
assign w4166 = v1498;
assign w4167 = w378 & ~w2849;
assign w4168 = (w1892 & ~w1704) | (w1892 & w1879) | (~w1704 & w1879);
assign w4169 = w656 & ~w1881;
assign v1499 = ~(w2196 | w2508);
assign w4170 = v1499;
assign w4171 = w2893 & ~w4047;
assign v1500 = ~(w2794 | w1027);
assign w4172 = v1500;
assign w4173 = w656 & ~w1444;
assign v1501 = ~(w2175 | w3414);
assign w4174 = v1501;
assign w4175 = w4090 & w707;
assign v1502 = ~(w1661 | w1604);
assign w4176 = v1502;
assign w4177 = w3094 & w1860;
assign w4178 = ~w1022 & w3917;
assign w4179 = pi146 & w1570;
assign v1503 = ~(w1661 | w2085);
assign w4180 = v1503;
assign v1504 = ~(w3545 | w937);
assign w4181 = v1504;
assign w4182 = w3443 & w3327;
assign v1505 = ~(w3510 | w1361);
assign w4183 = v1505;
assign w4184 = pi351 & ~pi366;
assign w4185 = w2268 & w3882;
assign one = 1;
assign po00 = ~w855;// level 22
assign po01 = ~w2215;// level 5
assign po02 = ~w3528;// level 21
assign po03 = ~w2179;// level 5
assign po04 = w1360;// level 21
assign po05 = ~w1080;// level 5
assign po06 = ~w380;// level 21
assign po07 = ~w2099;// level 5
assign po08 = ~w2163;// level 21
assign po09 = ~w4158;// level 5
assign po10 = ~w4030;// level 21
assign po11 = ~w470;// level 5
assign po12 = ~w4095;// level 21
assign po13 = ~w1024;// level 5
assign po14 = ~w1055;// level 21
assign po15 = ~w3887;// level 5
assign po16 = ~w957;// level 22
assign po17 = ~w2462;// level 5
assign po18 = ~w491;// level 21
assign po19 = ~w203;// level 5
assign po20 = w1781;// level 21
assign po21 = ~w1566;// level 5
assign po22 = ~w3456;// level 21
assign po23 = ~w3773;// level 5
assign po24 = w3433;// level 21
assign po25 = ~w1330;// level 5
assign po26 = ~w3492;// level 21
assign po27 = ~w1653;// level 5
assign po28 = w870;// level 21
assign po29 = ~w2968;// level 5
assign po30 = ~w3599;// level 21
assign po31 = ~w2411;// level 5
assign po32 = w1026;// level 21
assign po33 = ~w1333;// level 5
assign po34 = w1736;// level 21
assign po35 = ~w3380;// level 5
assign po36 = w1524;// level 21
assign po37 = ~w3422;// level 5
assign po38 = w3289;// level 21
assign po39 = ~w3706;// level 5
assign po40 = w2741;// level 22
assign po41 = ~w3269;// level 5
assign po42 = ~w499;// level 21
assign po43 = ~w2631;// level 5
assign po44 = w2051;// level 22
assign po45 = ~w847;// level 5
assign po46 = ~w1079;// level 21
assign po47 = ~w2676;// level 5
assign po48 = ~w3926;// level 21
assign po49 = ~w3064;// level 5
assign po50 = w4042;// level 21
assign po51 = ~w373;// level 5
assign po52 = ~w1766;// level 21
assign po53 = ~w3273;// level 5
assign po54 = ~w4106;// level 21
assign po55 = ~w2840;// level 5
assign po56 = ~w1675;// level 21
assign po57 = ~w1317;// level 5
assign po58 = w417;// level 22
assign po59 = ~w876;// level 5
assign po60 = ~w3880;// level 21
assign po61 = ~w893;// level 5
assign po62 = ~w1553;// level 21
assign po63 = ~w324;// level 5
assign po64 = pi361;// level 0
assign po65 = one;// level 0
assign po66 = w1781;// level 21
assign po67 = w1524;// level 21
assign po68 = ~w1553;// level 21
assign po69 = ~w957;// level 22
assign po70 = ~w4030;// level 21
assign po71 = w417;// level 22
endmodule
