// Benchmark "simple_spi" written by ABC on Wed Apr 29 13:50:50 2015

module simple_spi ( 
    pi000, pi001, pi002, pi003, pi004, pi005, pi006, pi007, pi008, pi009,
    pi010, pi011, pi012, pi013, pi014, pi015, pi016, pi017, pi018, pi019,
    pi020, pi021, pi022, pi023, pi024, pi025, pi026, pi027, pi028, pi029,
    pi030, pi031, pi032, pi033, pi034, pi035, pi036, pi037, pi038, pi039,
    pi040, pi041, pi042, pi043, pi044, pi045, pi046, pi047, pi048, pi049,
    pi050, pi051, pi052, pi053, pi054, pi055, pi056, pi057, pi058, pi059,
    pi060, pi061, pi062, pi063, pi064, pi065, pi066, pi067, pi068, pi069,
    pi070, pi071, pi072, pi073, pi074, pi075, pi076, pi077, pi078, pi079,
    pi080, pi081, pi082, pi083, pi084, pi085, pi086, pi087, pi088, pi089,
    pi090, pi091, pi092, pi093, pi094, pi095, pi096, pi097, pi098, pi099,
    pi100, pi101, pi102, pi103, pi104, pi105, pi106, pi107, pi108, pi109,
    pi110, pi111, pi112, pi113, pi114, pi115, pi116, pi117, pi118, pi119,
    pi120, pi121, pi122, pi123, pi124, pi125, pi126, pi127, pi128, pi129,
    pi130, pi131, pi132, pi133, pi134, pi135, pi136, pi137, pi138, pi139,
    pi140, pi141, pi142, pi143, pi144, pi145, pi146, pi147,
    po000, po001, po002, po003, po004, po005, po006, po007, po008, po009,
    po010, po011, po012, po013, po014, po015, po016, po017, po018, po019,
    po020, po021, po022, po023, po024, po025, po026, po027, po028, po029,
    po030, po031, po032, po033, po034, po035, po036, po037, po038, po039,
    po040, po041, po042, po043, po044, po045, po046, po047, po048, po049,
    po050, po051, po052, po053, po054, po055, po056, po057, po058, po059,
    po060, po061, po062, po063, po064, po065, po066, po067, po068, po069,
    po070, po071, po072, po073, po074, po075, po076, po077, po078, po079,
    po080, po081, po082, po083, po084, po085, po086, po087, po088, po089,
    po090, po091, po092, po093, po094, po095, po096, po097, po098, po099,
    po100, po101, po102, po103, po104, po105, po106, po107, po108, po109,
    po110, po111, po112, po113, po114, po115, po116, po117, po118, po119,
    po120, po121, po122, po123, po124, po125, po126, po127, po128, po129,
    po130, po131, po132, po133, po134, po135, po136, po137, po138, po139,
    po140, po141, po142, po143, po144, po145, po146  );
  input  pi000, pi001, pi002, pi003, pi004, pi005, pi006, pi007, pi008,
    pi009, pi010, pi011, pi012, pi013, pi014, pi015, pi016, pi017, pi018,
    pi019, pi020, pi021, pi022, pi023, pi024, pi025, pi026, pi027, pi028,
    pi029, pi030, pi031, pi032, pi033, pi034, pi035, pi036, pi037, pi038,
    pi039, pi040, pi041, pi042, pi043, pi044, pi045, pi046, pi047, pi048,
    pi049, pi050, pi051, pi052, pi053, pi054, pi055, pi056, pi057, pi058,
    pi059, pi060, pi061, pi062, pi063, pi064, pi065, pi066, pi067, pi068,
    pi069, pi070, pi071, pi072, pi073, pi074, pi075, pi076, pi077, pi078,
    pi079, pi080, pi081, pi082, pi083, pi084, pi085, pi086, pi087, pi088,
    pi089, pi090, pi091, pi092, pi093, pi094, pi095, pi096, pi097, pi098,
    pi099, pi100, pi101, pi102, pi103, pi104, pi105, pi106, pi107, pi108,
    pi109, pi110, pi111, pi112, pi113, pi114, pi115, pi116, pi117, pi118,
    pi119, pi120, pi121, pi122, pi123, pi124, pi125, pi126, pi127, pi128,
    pi129, pi130, pi131, pi132, pi133, pi134, pi135, pi136, pi137, pi138,
    pi139, pi140, pi141, pi142, pi143, pi144, pi145, pi146, pi147;
  output po000, po001, po002, po003, po004, po005, po006, po007, po008, po009,
    po010, po011, po012, po013, po014, po015, po016, po017, po018, po019,
    po020, po021, po022, po023, po024, po025, po026, po027, po028, po029,
    po030, po031, po032, po033, po034, po035, po036, po037, po038, po039,
    po040, po041, po042, po043, po044, po045, po046, po047, po048, po049,
    po050, po051, po052, po053, po054, po055, po056, po057, po058, po059,
    po060, po061, po062, po063, po064, po065, po066, po067, po068, po069,
    po070, po071, po072, po073, po074, po075, po076, po077, po078, po079,
    po080, po081, po082, po083, po084, po085, po086, po087, po088, po089,
    po090, po091, po092, po093, po094, po095, po096, po097, po098, po099,
    po100, po101, po102, po103, po104, po105, po106, po107, po108, po109,
    po110, po111, po112, po113, po114, po115, po116, po117, po118, po119,
    po120, po121, po122, po123, po124, po125, po126, po127, po128, po129,
    po130, po131, po132, po133, po134, po135, po136, po137, po138, po139,
    po140, po141, po142, po143, po144, po145, po146;
  wire n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, n307,
    n308, n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
    n321, n322, n323, n324, n325, n326, n327, n328, n330, n331, n332, n333,
    n334, n335, n336, n337, n339, n340, n341, n342, n343, n344, n345, n346,
    n347, n349, n350, n351, n353, n354, n355, n357, n358, n359, n360, n361,
    n363, n364, n365, n366, n367, n369, n370, n371, n372, n373, n375, n376,
    n377, n378, n379, n381, n382, n383, n384, n385, n387, n388, n389, n390,
    n391, n393, n394, n395, n396, n397, n399, n400, n401, n402, n403, n405,
    n406, n407, n408, n409, n411, n412, n413, n414, n415, n417, n418, n419,
    n420, n421, n423, n424, n425, n426, n427, n429, n430, n431, n432, n433,
    n435, n436, n437, n438, n439, n441, n442, n443, n444, n445, n447, n448,
    n449, n450, n451, n453, n454, n455, n456, n457, n458, n460, n461, n462,
    n463, n464, n466, n467, n468, n469, n470, n472, n473, n474, n475, n476,
    n478, n479, n480, n481, n482, n484, n485, n486, n487, n488, n490, n491,
    n492, n493, n494, n496, n497, n498, n499, n500, n502, n503, n504, n505,
    n506, n507, n509, n510, n511, n512, n513, n515, n516, n517, n518, n519,
    n521, n522, n523, n524, n525, n527, n528, n529, n530, n531, n533, n534,
    n535, n536, n537, n539, n540, n541, n542, n543, n545, n546, n547, n548,
    n549, n551, n552, n553, n554, n555, n556, n557, n558, n559, n560, n561,
    n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
    n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585,
    n586, n587, n588, n589, n590, n591, n592, n593, n594, n595, n596, n597,
    n598, n599, n600, n601, n602, n603, n604, n606, n607, n608, n609, n610,
    n611, n612, n613, n614, n615, n616, n618, n619, n620, n621, n622, n623,
    n624, n625, n626, n627, n629, n630, n631, n632, n633, n634, n635, n636,
    n637, n639, n640, n641, n642, n643, n644, n645, n646, n647, n648, n649,
    n650, n651, n652, n654, n655, n656, n657, n658, n659, n660, n661, n662,
    n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, n674, n675,
    n676, n677, n678, n679, n680, n681, n682, n684, n685, n686, n687, n688,
    n689, n690, n691, n692, n693, n694, n695, n696, n697, n698, n700, n701,
    n702, n703, n704, n705, n706, n707, n708, n709, n710, n711, n712, n713,
    n714, n716, n717, n718, n719, n720, n721, n722, n723, n724, n725, n726,
    n727, n728, n729, n730, n732, n733, n734, n735, n736, n737, n738, n739,
    n740, n741, n742, n743, n744, n745, n746, n748, n749, n750, n751, n752,
    n753, n754, n755, n756, n757, n758, n759, n760, n761, n762, n764, n765,
    n766, n767, n768, n769, n770, n771, n772, n773, n774, n775, n776, n777,
    n778, n780, n781, n782, n783, n784, n785, n786, n787, n788, n789, n790,
    n791, n792, n793, n794, n796, n797, n798, n799, n800, n801, n802, n803,
    n804, n805, n806, n808, n809, n810, n811, n812, n813, n814, n816, n817,
    n818, n819, n820, n821, n822, n823, n824, n825, n827, n828, n829, n830,
    n831, n832, n833, n834, n836, n837, n838, n839, n840, n841, n842, n844,
    n845, n846, n847, n848, n849, n850, n851, n852, n853, n854, n856, n857,
    n858, n859, n860, n861, n863, n864, n865, n866, n867, n869, n870, n871,
    n873, n874, n875, n876, n878, n879, n880, n881, n883, n884, n886, n887,
    n888, n889, n890, n891, n892, n893, n895, n896, n897, n898, n899, n900,
    n901, n902, n903, n904, n905, n906, n907, n908, n909, n910, n911, n912,
    n913, n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925,
    n927, n928, n929, n930, n931, n932, n933, n934, n935, n936, n937, n938,
    n939, n940, n942, n943, n944, n945, n946, n947, n948, n949, n950, n951,
    n952, n953, n954, n956, n957, n958, n959, n960, n961, n962, n963, n964,
    n965, n966, n967, n968, n969, n970, n971, n972, n973, n975, n976, n977,
    n978, n979, n980, n981, n982, n983, n984, n985, n987, n988, n989, n990,
    n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1002,
    n1003, n1004, n1005, n1006, n1008, n1009, n1010, n1011, n1012, n1013,
    n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1022, n1023, n1024,
    n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1034, n1035,
    n1036, n1037, n1039, n1040, n1041, n1042, n1044, n1045, n1046, n1048,
    n1049, n1050, n1051, n1052, n1054, n1055, n1056, n1057, n1058, n1060,
    n1061, n1062, n1063, n1064, n1066, n1067, n1068, n1069, n1070, n1072,
    n1073, n1074, n1076, n1077, n1078, n1080, n1081, n1082, n1083, n1084,
    n1086, n1087, n1088, n1089, n1090, n1092, n1093, n1094, n1095, n1096,
    n1098, n1099, n1100, n1101, n1102, n1104, n1105, n1106, n1107, n1108,
    n1110, n1111, n1112, n1113, n1114, n1116, n1117, n1118, n1119, n1120,
    n1122, n1123, n1124, n1125, n1126, n1128, n1129, n1130, n1131, n1132,
    n1134, n1135, n1136, n1137, n1138, n1140, n1141, n1142, n1143, n1144,
    n1146, n1147, n1148, n1149, n1150, n1152, n1153, n1154, n1155, n1156,
    n1157, n1159, n1160, n1161, n1162, n1163, n1164, n1166, n1167, n1168,
    n1169, n1170, n1172, n1173, n1174, n1175, n1176, n1178, n1179, n1180,
    n1181, n1182, n1184, n1185, n1186, n1187, n1188, n1190, n1191, n1192,
    n1193, n1194, n1196, n1197, n1198, n1199, n1200, n1202, n1203, n1204,
    n1205, n1206, n1208, n1209, n1210, n1211, n1212, n1214, n1215, n1216,
    n1217, n1218, n1220, n1221, n1222, n1223, n1224, n1226, n1227, n1228,
    n1229, n1230, n1232, n1233, n1234, n1235, n1236, n1238, n1239, n1240,
    n1241, n1242, n1244, n1245, n1246, n1247, n1248, n1250, n1251, n1252,
    n1253, n1254, n1256, n1258, n1259, n1260, n1261, n1262, n1264, n1265,
    n1266, n1267, n1268, n1270, n1271, n1272, n1273, n1274, n1276, n1277,
    n1278, n1279, n1280, n1282, n1283, n1284, n1285, n1286, n1288, n1289,
    n1290, n1291, n1292, n1294, n1295, n1296, n1297, n1298, n1300, n1301,
    n1302, n1303, n1304, n1306, n1307, n1308, n1309, n1310, n1312, n1313,
    n1314, n1315, n1316, n1318, n1319, n1320, n1321, n1322, n1324, n1326,
    n1327, n1328, n1329, n1330, n1332, n1333, n1334, n1335, n1336, n1338,
    n1339, n1340, n1341, n1342, n1344, n1345, n1346;
  assign n297 = pi000 & pi128;
  assign n298 = pi063 & n297;
  assign n299 = pi120 & ~pi128;
  assign n300 = ~n298 & ~n299;
  assign n301 = ~pi063 & pi120;
  assign n302 = ~pi000 & ~pi002;
  assign n303 = n301 & n302;
  assign n304 = pi000 & ~pi063;
  assign n305 = ~n302 & n304;
  assign n306 = pi002 & n305;
  assign n307 = ~n303 & ~n306;
  assign n308 = pi128 & ~n307;
  assign po014 = ~n300 | n308;
  assign n310 = pi128 & pi133;
  assign n311 = ~pi138 & pi139;
  assign n312 = pi130 & n311;
  assign n313 = pi134 & pi135;
  assign n314 = ~pi136 & n313;
  assign n315 = n312 & n314;
  assign n316 = pi001 & ~n315;
  assign n317 = pi004 & ~pi005;
  assign n318 = ~pi004 & pi005;
  assign n319 = ~n317 & ~n318;
  assign n320 = pi075 & n319;
  assign n321 = ~pi075 & ~n319;
  assign n322 = ~n320 & ~n321;
  assign n323 = ~pi063 & n322;
  assign n324 = ~pi005 & ~pi077;
  assign n325 = pi005 & pi077;
  assign n326 = ~n324 & ~n325;
  assign n327 = n323 & n326;
  assign n328 = ~n316 & ~n327;
  assign po015 = n310 & ~n328;
  assign n330 = pi119 & ~pi128;
  assign n331 = pi002 & pi063;
  assign n332 = ~pi002 & ~n302;
  assign n333 = pi119 & n302;
  assign n334 = ~n332 & ~n333;
  assign n335 = ~pi063 & ~n334;
  assign n336 = ~n331 & ~n335;
  assign n337 = pi128 & ~n336;
  assign po016 = n330 | n337;
  assign n339 = pi003 & pi128;
  assign n340 = pi136 & n313;
  assign n341 = pi138 & ~pi139;
  assign n342 = pi147 & n341;
  assign n343 = n340 & n342;
  assign n344 = n339 & ~n343;
  assign n345 = ~pi063 & pi128;
  assign n346 = ~n343 & n345;
  assign n347 = n302 & n346;
  assign po017 = n344 | n347;
  assign n349 = pi004 & pi063;
  assign n350 = ~pi063 & ~n319;
  assign n351 = ~n349 & ~n350;
  assign po019 = pi128 & ~n351;
  assign n353 = pi005 & pi063;
  assign n354 = ~pi005 & ~pi063;
  assign n355 = ~n353 & ~n354;
  assign po020 = pi128 & ~n355;
  assign n357 = pi046 & n318;
  assign n358 = pi006 & ~n318;
  assign n359 = ~n357 & ~n358;
  assign n360 = ~pi063 & ~n359;
  assign n361 = pi006 & pi063;
  assign po021 = n360 | n361;
  assign n363 = pi047 & n318;
  assign n364 = pi007 & ~n318;
  assign n365 = ~n363 & ~n364;
  assign n366 = ~pi063 & ~n365;
  assign n367 = pi007 & pi063;
  assign po022 = n366 | n367;
  assign n369 = pi048 & n318;
  assign n370 = pi008 & ~n318;
  assign n371 = ~n369 & ~n370;
  assign n372 = ~pi063 & ~n371;
  assign n373 = pi008 & pi063;
  assign po023 = n372 | n373;
  assign n375 = pi049 & n318;
  assign n376 = pi009 & ~n318;
  assign n377 = ~n375 & ~n376;
  assign n378 = ~pi063 & ~n377;
  assign n379 = pi009 & pi063;
  assign po024 = n378 | n379;
  assign n381 = pi043 & n318;
  assign n382 = pi010 & ~n318;
  assign n383 = ~n381 & ~n382;
  assign n384 = ~pi063 & ~n383;
  assign n385 = pi010 & pi063;
  assign po025 = n384 | n385;
  assign n387 = pi050 & n317;
  assign n388 = pi011 & ~n317;
  assign n389 = ~n387 & ~n388;
  assign n390 = ~pi063 & ~n389;
  assign n391 = pi011 & pi063;
  assign po026 = n390 | n391;
  assign n393 = pi051 & n317;
  assign n394 = pi012 & ~n317;
  assign n395 = ~n393 & ~n394;
  assign n396 = ~pi063 & ~n395;
  assign n397 = pi012 & pi063;
  assign po027 = n396 | n397;
  assign n399 = pi045 & n317;
  assign n400 = pi013 & ~n317;
  assign n401 = ~n399 & ~n400;
  assign n402 = ~pi063 & ~n401;
  assign n403 = pi013 & pi063;
  assign po028 = n402 | n403;
  assign n405 = pi046 & n317;
  assign n406 = pi014 & ~n317;
  assign n407 = ~n405 & ~n406;
  assign n408 = ~pi063 & ~n407;
  assign n409 = pi014 & pi063;
  assign po029 = n408 | n409;
  assign n411 = pi047 & n317;
  assign n412 = pi015 & ~n317;
  assign n413 = ~n411 & ~n412;
  assign n414 = ~pi063 & ~n413;
  assign n415 = pi015 & pi063;
  assign po030 = n414 | n415;
  assign n417 = pi048 & n317;
  assign n418 = pi016 & ~n317;
  assign n419 = ~n417 & ~n418;
  assign n420 = ~pi063 & ~n419;
  assign n421 = pi016 & pi063;
  assign po031 = n420 | n421;
  assign n423 = pi049 & n317;
  assign n424 = pi017 & ~n317;
  assign n425 = ~n423 & ~n424;
  assign n426 = ~pi063 & ~n425;
  assign n427 = pi017 & pi063;
  assign po032 = n426 | n427;
  assign n429 = pi043 & n317;
  assign n430 = pi018 & ~n317;
  assign n431 = ~n429 & ~n430;
  assign n432 = ~pi063 & ~n431;
  assign n433 = pi018 & pi063;
  assign po033 = n432 | n433;
  assign n435 = pi050 & n318;
  assign n436 = pi019 & ~n318;
  assign n437 = ~n435 & ~n436;
  assign n438 = ~pi063 & ~n437;
  assign n439 = pi019 & pi063;
  assign po034 = n438 | n439;
  assign n441 = pi051 & n318;
  assign n442 = pi020 & ~n318;
  assign n443 = ~n441 & ~n442;
  assign n444 = ~pi063 & ~n443;
  assign n445 = pi020 & pi063;
  assign po035 = n444 | n445;
  assign n447 = pi045 & n318;
  assign n448 = pi021 & ~n318;
  assign n449 = ~n447 & ~n448;
  assign n450 = ~pi063 & ~n449;
  assign n451 = pi021 & pi063;
  assign po036 = n450 | n451;
  assign n453 = pi004 & pi005;
  assign n454 = pi050 & n453;
  assign n455 = pi022 & ~n453;
  assign n456 = ~n454 & ~n455;
  assign n457 = ~pi063 & ~n456;
  assign n458 = pi022 & pi063;
  assign po037 = n457 | n458;
  assign n460 = pi051 & n453;
  assign n461 = pi023 & ~n453;
  assign n462 = ~n460 & ~n461;
  assign n463 = ~pi063 & ~n462;
  assign n464 = pi023 & pi063;
  assign po038 = n463 | n464;
  assign n466 = pi045 & n453;
  assign n467 = pi024 & ~n453;
  assign n468 = ~n466 & ~n467;
  assign n469 = ~pi063 & ~n468;
  assign n470 = pi024 & pi063;
  assign po039 = n469 | n470;
  assign n472 = pi046 & n453;
  assign n473 = pi025 & ~n453;
  assign n474 = ~n472 & ~n473;
  assign n475 = ~pi063 & ~n474;
  assign n476 = pi025 & pi063;
  assign po040 = n475 | n476;
  assign n478 = pi047 & n453;
  assign n479 = pi026 & ~n453;
  assign n480 = ~n478 & ~n479;
  assign n481 = ~pi063 & ~n480;
  assign n482 = pi026 & pi063;
  assign po041 = n481 | n482;
  assign n484 = pi048 & n453;
  assign n485 = pi027 & ~n453;
  assign n486 = ~n484 & ~n485;
  assign n487 = ~pi063 & ~n486;
  assign n488 = pi027 & pi063;
  assign po042 = n487 | n488;
  assign n490 = pi049 & n453;
  assign n491 = pi028 & ~n453;
  assign n492 = ~n490 & ~n491;
  assign n493 = ~pi063 & ~n492;
  assign n494 = pi028 & pi063;
  assign po043 = n493 | n494;
  assign n496 = pi043 & n453;
  assign n497 = pi029 & ~n453;
  assign n498 = ~n496 & ~n497;
  assign n499 = ~pi063 & ~n498;
  assign n500 = pi029 & pi063;
  assign po044 = n499 | n500;
  assign n502 = ~pi004 & ~pi005;
  assign n503 = pi030 & ~n502;
  assign n504 = pi050 & n502;
  assign n505 = ~n503 & ~n504;
  assign n506 = ~pi063 & ~n505;
  assign n507 = pi030 & pi063;
  assign po045 = n506 | n507;
  assign n509 = pi031 & ~n502;
  assign n510 = pi051 & n502;
  assign n511 = ~n509 & ~n510;
  assign n512 = ~pi063 & ~n511;
  assign n513 = pi031 & pi063;
  assign po046 = n512 | n513;
  assign n515 = pi032 & ~n502;
  assign n516 = pi046 & n502;
  assign n517 = ~n515 & ~n516;
  assign n518 = ~pi063 & ~n517;
  assign n519 = pi032 & pi063;
  assign po047 = n518 | n519;
  assign n521 = pi033 & ~n502;
  assign n522 = pi047 & n502;
  assign n523 = ~n521 & ~n522;
  assign n524 = ~pi063 & ~n523;
  assign n525 = pi033 & pi063;
  assign po048 = n524 | n525;
  assign n527 = pi034 & ~n502;
  assign n528 = pi048 & n502;
  assign n529 = ~n527 & ~n528;
  assign n530 = ~pi063 & ~n529;
  assign n531 = pi034 & pi063;
  assign po049 = n530 | n531;
  assign n533 = pi035 & ~n502;
  assign n534 = pi043 & n502;
  assign n535 = ~n533 & ~n534;
  assign n536 = ~pi063 & ~n535;
  assign n537 = pi035 & pi063;
  assign po050 = n536 | n537;
  assign n539 = pi036 & ~n502;
  assign n540 = pi045 & n502;
  assign n541 = ~n539 & ~n540;
  assign n542 = ~pi063 & ~n541;
  assign n543 = pi036 & pi063;
  assign po051 = n542 | n543;
  assign n545 = pi037 & ~n502;
  assign n546 = pi049 & n502;
  assign n547 = ~n545 & ~n546;
  assign n548 = ~pi063 & ~n547;
  assign n549 = pi037 & pi063;
  assign po052 = n548 | n549;
  assign n551 = pi076 & pi082;
  assign n552 = ~pi076 & ~pi082;
  assign n553 = ~n551 & ~n552;
  assign n554 = ~pi083 & ~pi129;
  assign n555 = pi083 & pi129;
  assign n556 = ~n554 & ~n555;
  assign n557 = ~n553 & ~n556;
  assign n558 = ~pi066 & n557;
  assign n559 = ~pi038 & pi124;
  assign n560 = ~pi124 & pi127;
  assign n561 = ~n559 & ~n560;
  assign n562 = ~n558 & ~n561;
  assign n563 = pi127 & ~n553;
  assign n564 = ~pi066 & n563;
  assign n565 = ~n556 & n564;
  assign n566 = ~n562 & ~n565;
  assign n567 = ~pi039 & ~pi062;
  assign n568 = ~n566 & n567;
  assign n569 = ~pi058 & ~pi060;
  assign n570 = ~pi056 & ~pi061;
  assign n571 = n569 & n570;
  assign n572 = ~pi052 & ~pi064;
  assign n573 = ~pi042 & ~pi057;
  assign n574 = n572 & n573;
  assign n575 = ~pi053 & ~pi054;
  assign n576 = ~pi055 & ~pi059;
  assign n577 = n575 & n576;
  assign n578 = n574 & n577;
  assign n579 = n571 & n578;
  assign n580 = ~pi038 & n579;
  assign n581 = pi038 & ~n579;
  assign n582 = ~n580 & ~n581;
  assign n583 = pi039 & ~pi062;
  assign n584 = ~n582 & n583;
  assign n585 = ~pi039 & pi062;
  assign n586 = pi038 & n585;
  assign n587 = pi039 & pi062;
  assign n588 = ~pi059 & ~pi060;
  assign n589 = ~pi055 & ~pi058;
  assign n590 = n588 & n589;
  assign n591 = ~pi040 & ~pi044;
  assign n592 = ~pi041 & n591;
  assign n593 = pi127 & n592;
  assign n594 = ~pi038 & ~n592;
  assign n595 = ~n593 & ~n594;
  assign n596 = n570 & n575;
  assign n597 = n574 & n596;
  assign n598 = ~n595 & n597;
  assign n599 = n590 & n598;
  assign n600 = ~n581 & ~n599;
  assign n601 = n587 & ~n600;
  assign n602 = ~n586 & ~n601;
  assign n603 = ~n584 & n602;
  assign n604 = ~n568 & n603;
  assign po053 = pi128 & ~n604;
  assign n606 = pi039 & n583;
  assign n607 = n579 & ~n592;
  assign n608 = pi039 & ~n579;
  assign n609 = ~n607 & ~n608;
  assign n610 = n587 & ~n609;
  assign n611 = n579 & n583;
  assign n612 = ~pi039 & n558;
  assign n613 = n567 & ~n612;
  assign n614 = ~n611 & ~n613;
  assign n615 = ~n610 & n614;
  assign n616 = ~n606 & n615;
  assign po054 = pi128 & ~n616;
  assign n618 = ~n583 & ~n585;
  assign n619 = pi040 & ~n618;
  assign n620 = ~n567 & ~n619;
  assign n621 = pi128 & ~n620;
  assign n622 = pi040 & n579;
  assign n623 = ~pi040 & ~n579;
  assign n624 = ~n622 & ~n623;
  assign n625 = pi062 & pi128;
  assign n626 = pi039 & n625;
  assign n627 = n624 & n626;
  assign po055 = n621 | n627;
  assign n629 = pi041 & ~n591;
  assign n630 = ~n592 & ~n629;
  assign n631 = n579 & ~n630;
  assign n632 = pi041 & ~n579;
  assign n633 = ~n631 & ~n632;
  assign n634 = n587 & ~n633;
  assign n635 = pi041 & ~n618;
  assign n636 = ~n634 & ~n635;
  assign n637 = ~n567 & n636;
  assign po056 = pi128 & ~n637;
  assign n639 = pi128 & ~n567;
  assign n640 = ~n579 & n639;
  assign n641 = pi115 & pi123;
  assign n642 = ~n640 & n641;
  assign n643 = ~pi059 & n589;
  assign n644 = ~pi060 & n643;
  assign n645 = n596 & n644;
  assign n646 = ~pi042 & n645;
  assign n647 = pi042 & ~n645;
  assign n648 = ~n646 & ~n647;
  assign n649 = n640 & ~n648;
  assign n650 = ~n642 & ~n649;
  assign n651 = pi115 & pi126;
  assign n652 = ~n640 & n651;
  assign po057 = ~n650 | n652;
  assign n654 = pi049 & n579;
  assign n655 = pi043 & ~n579;
  assign n656 = ~n654 & ~n655;
  assign n657 = n587 & ~n656;
  assign n658 = pi043 & ~n618;
  assign n659 = ~n657 & ~n658;
  assign n660 = pi076 & ~pi129;
  assign n661 = pi095 & n660;
  assign n662 = pi076 & pi129;
  assign n663 = pi111 & n662;
  assign n664 = ~n661 & ~n663;
  assign n665 = ~pi076 & ~pi129;
  assign n666 = pi099 & n665;
  assign n667 = ~pi076 & pi129;
  assign n668 = pi089 & n667;
  assign n669 = ~n666 & ~n668;
  assign n670 = n664 & n669;
  assign n671 = n567 & ~n670;
  assign n672 = n659 & ~n671;
  assign po058 = pi128 & ~n672;
  assign n674 = pi040 & pi044;
  assign n675 = ~n591 & ~n674;
  assign n676 = n579 & ~n675;
  assign n677 = pi044 & ~n579;
  assign n678 = ~n676 & ~n677;
  assign n679 = n587 & ~n678;
  assign n680 = pi044 & ~n618;
  assign n681 = ~n679 & ~n680;
  assign n682 = ~n567 & n681;
  assign po059 = pi128 & ~n682;
  assign n684 = pi107 & n662;
  assign n685 = pi086 & n667;
  assign n686 = ~n684 & ~n685;
  assign n687 = pi102 & n665;
  assign n688 = pi091 & n660;
  assign n689 = ~n687 & ~n688;
  assign n690 = n686 & n689;
  assign n691 = n567 & ~n690;
  assign n692 = pi051 & n579;
  assign n693 = pi045 & ~n579;
  assign n694 = ~n692 & ~n693;
  assign n695 = n587 & ~n694;
  assign n696 = pi045 & ~n618;
  assign n697 = ~n695 & ~n696;
  assign n698 = ~n691 & n697;
  assign po060 = pi128 & ~n698;
  assign n700 = pi092 & n660;
  assign n701 = pi108 & n662;
  assign n702 = ~n700 & ~n701;
  assign n703 = pi103 & n665;
  assign n704 = pi087 & n667;
  assign n705 = ~n703 & ~n704;
  assign n706 = n702 & n705;
  assign n707 = n567 & ~n706;
  assign n708 = pi045 & n579;
  assign n709 = pi046 & ~n579;
  assign n710 = ~n708 & ~n709;
  assign n711 = n587 & ~n710;
  assign n712 = pi046 & ~n618;
  assign n713 = ~n711 & ~n712;
  assign n714 = ~n707 & n713;
  assign po061 = pi128 & ~n714;
  assign n716 = pi078 & n660;
  assign n717 = pi097 & n662;
  assign n718 = ~n716 & ~n717;
  assign n719 = pi096 & n665;
  assign n720 = pi081 & n667;
  assign n721 = ~n719 & ~n720;
  assign n722 = n718 & n721;
  assign n723 = n567 & ~n722;
  assign n724 = pi046 & n579;
  assign n725 = pi047 & ~n579;
  assign n726 = ~n724 & ~n725;
  assign n727 = n587 & ~n726;
  assign n728 = pi047 & ~n618;
  assign n729 = ~n727 & ~n728;
  assign n730 = ~n723 & n729;
  assign po062 = pi128 & ~n730;
  assign n732 = pi093 & n660;
  assign n733 = pi109 & n662;
  assign n734 = ~n732 & ~n733;
  assign n735 = pi105 & n665;
  assign n736 = pi088 & n667;
  assign n737 = ~n735 & ~n736;
  assign n738 = n734 & n737;
  assign n739 = n567 & ~n738;
  assign n740 = pi047 & n579;
  assign n741 = pi048 & ~n579;
  assign n742 = ~n740 & ~n741;
  assign n743 = n587 & ~n742;
  assign n744 = pi048 & ~n618;
  assign n745 = ~n743 & ~n744;
  assign n746 = ~n739 & n745;
  assign po063 = pi128 & ~n746;
  assign n748 = pi094 & n660;
  assign n749 = pi110 & n662;
  assign n750 = ~n748 & ~n749;
  assign n751 = pi104 & n665;
  assign n752 = pi079 & n667;
  assign n753 = ~n751 & ~n752;
  assign n754 = n750 & n753;
  assign n755 = n567 & ~n754;
  assign n756 = pi048 & n579;
  assign n757 = pi049 & ~n579;
  assign n758 = ~n756 & ~n757;
  assign n759 = n587 & ~n758;
  assign n760 = pi049 & ~n618;
  assign n761 = ~n759 & ~n760;
  assign n762 = ~n755 & n761;
  assign po064 = pi128 & ~n762;
  assign n764 = pi098 & n662;
  assign n765 = pi084 & n667;
  assign n766 = ~n764 & ~n765;
  assign n767 = pi100 & n665;
  assign n768 = pi080 & n660;
  assign n769 = ~n767 & ~n768;
  assign n770 = n766 & n769;
  assign n771 = n567 & ~n770;
  assign n772 = pi137 & n579;
  assign n773 = pi050 & ~n579;
  assign n774 = ~n772 & ~n773;
  assign n775 = n587 & ~n774;
  assign n776 = pi050 & ~n618;
  assign n777 = ~n775 & ~n776;
  assign n778 = ~n771 & n777;
  assign po065 = pi128 & ~n778;
  assign n780 = pi090 & n660;
  assign n781 = pi106 & n662;
  assign n782 = ~n780 & ~n781;
  assign n783 = pi101 & n665;
  assign n784 = pi085 & n667;
  assign n785 = ~n783 & ~n784;
  assign n786 = n782 & n785;
  assign n787 = n567 & ~n786;
  assign n788 = pi050 & n579;
  assign n789 = pi051 & ~n579;
  assign n790 = ~n788 & ~n789;
  assign n791 = n587 & ~n790;
  assign n792 = pi051 & ~n618;
  assign n793 = ~n791 & ~n792;
  assign n794 = ~n787 & n793;
  assign po066 = pi128 & ~n794;
  assign n796 = ~pi053 & ~pi056;
  assign n797 = n573 & n796;
  assign n798 = ~pi054 & ~pi061;
  assign n799 = n588 & n798;
  assign n800 = n589 & n799;
  assign n801 = n797 & n800;
  assign n802 = pi052 & ~n801;
  assign n803 = ~pi052 & n801;
  assign n804 = ~n802 & ~n803;
  assign n805 = n640 & ~n804;
  assign n806 = pi123 & n652;
  assign po067 = n805 | n806;
  assign n808 = pi115 & ~n640;
  assign n809 = ~pi056 & n798;
  assign n810 = n644 & n809;
  assign n811 = pi053 & ~n810;
  assign n812 = ~pi053 & n810;
  assign n813 = ~n811 & ~n812;
  assign n814 = n640 & ~n813;
  assign po068 = n808 | n814;
  assign n816 = pi114 & ~pi123;
  assign n817 = ~n640 & ~n816;
  assign n818 = pi054 & n644;
  assign n819 = ~pi054 & ~n644;
  assign n820 = ~n818 & ~n819;
  assign n821 = n640 & ~n820;
  assign n822 = ~n817 & ~n821;
  assign n823 = pi114 & pi126;
  assign n824 = ~pi115 & ~n823;
  assign n825 = ~n640 & ~n824;
  assign po069 = n822 | n825;
  assign n827 = ~pi058 & n588;
  assign n828 = pi055 & ~n827;
  assign n829 = ~n644 & ~n828;
  assign n830 = n640 & ~n829;
  assign n831 = ~pi115 & ~n816;
  assign n832 = pi123 & pi126;
  assign n833 = n831 & ~n832;
  assign n834 = ~n640 & ~n833;
  assign po070 = n830 | n834;
  assign n836 = pi056 & ~n800;
  assign n837 = ~pi056 & n800;
  assign n838 = ~n836 & ~n837;
  assign n839 = n640 & ~n838;
  assign n840 = pi123 & n823;
  assign n841 = ~pi115 & ~n840;
  assign n842 = ~n640 & ~n841;
  assign po071 = n839 | n842;
  assign n844 = ~pi042 & ~pi061;
  assign n845 = ~pi054 & ~pi059;
  assign n846 = ~pi060 & n589;
  assign n847 = n845 & n846;
  assign n848 = ~pi053 & n847;
  assign n849 = ~pi056 & n848;
  assign n850 = n844 & n849;
  assign n851 = pi057 & ~n850;
  assign n852 = ~pi057 & n850;
  assign n853 = ~n851 & ~n852;
  assign n854 = n640 & ~n853;
  assign po072 = n652 | n854;
  assign n856 = pi058 & ~n588;
  assign n857 = ~n827 & ~n856;
  assign n858 = n640 & ~n857;
  assign n859 = ~pi114 & ~pi115;
  assign n860 = ~n832 & n859;
  assign n861 = ~n640 & ~n860;
  assign po073 = n858 | n861;
  assign n863 = ~pi123 & ~n640;
  assign n864 = pi059 & n640;
  assign n865 = ~n863 & ~n864;
  assign n866 = ~pi126 & n859;
  assign n867 = ~n640 & ~n866;
  assign po074 = n865 | n867;
  assign n869 = pi059 & pi060;
  assign n870 = ~n588 & ~n869;
  assign n871 = n640 & ~n870;
  assign po075 = n867 | n871;
  assign n873 = pi061 & ~n847;
  assign n874 = ~pi061 & n847;
  assign n875 = ~n873 & ~n874;
  assign n876 = n640 & ~n875;
  assign po076 = n825 | n876;
  assign n878 = ~n579 & n587;
  assign n879 = pi062 & n878;
  assign n880 = pi128 & n879;
  assign n881 = pi128 & n611;
  assign po077 = n880 | n881;
  assign n883 = n579 & n592;
  assign n884 = pi128 & n883;
  assign po078 = n587 & n884;
  assign n886 = ~pi052 & ~pi053;
  assign n887 = n573 & n886;
  assign n888 = n810 & n887;
  assign n889 = pi064 & ~n888;
  assign n890 = ~pi064 & n886;
  assign n891 = n810 & n890;
  assign n892 = n573 & n891;
  assign n893 = ~n889 & ~n892;
  assign po079 = n640 & ~n893;
  assign n895 = ~pi075 & pi077;
  assign n896 = pi009 & n895;
  assign n897 = pi075 & pi077;
  assign n898 = pi028 & n897;
  assign n899 = ~n896 & ~n898;
  assign n900 = ~pi075 & ~pi077;
  assign n901 = pi037 & n900;
  assign n902 = pi075 & ~pi077;
  assign n903 = pi017 & n902;
  assign n904 = ~n901 & ~n903;
  assign n905 = n899 & n904;
  assign n906 = n311 & ~n905;
  assign n907 = ~pi138 & ~pi139;
  assign n908 = pi128 & n907;
  assign n909 = ~n906 & ~n908;
  assign n910 = pi138 & pi139;
  assign n911 = pi119 & n910;
  assign n912 = ~pi072 & n341;
  assign n913 = ~n911 & ~n912;
  assign po080 = ~n909 | ~n913;
  assign n915 = pi066 & ~pi113;
  assign n916 = n312 & n340;
  assign n917 = pi082 & ~pi083;
  assign n918 = ~pi082 & pi083;
  assign n919 = ~n917 & ~n918;
  assign n920 = pi076 & ~n919;
  assign n921 = ~pi076 & n919;
  assign n922 = ~n920 & ~n921;
  assign n923 = n556 & ~n922;
  assign n924 = n916 & n923;
  assign n925 = ~n915 & ~n924;
  assign po081 = n310 & ~n925;
  assign n927 = pi006 & n895;
  assign n928 = pi014 & n902;
  assign n929 = ~n927 & ~n928;
  assign n930 = pi032 & n900;
  assign n931 = pi025 & n897;
  assign n932 = ~n930 & ~n931;
  assign n933 = n929 & n932;
  assign n934 = n311 & ~n933;
  assign n935 = pi066 & n557;
  assign n936 = n341 & n935;
  assign n937 = ~n934 & ~n936;
  assign n938 = pi127 & n907;
  assign n939 = pi117 & n910;
  assign n940 = ~n938 & ~n939;
  assign po082 = ~n937 | ~n940;
  assign n942 = pi013 & n902;
  assign n943 = pi036 & n900;
  assign n944 = ~n942 & ~n943;
  assign n945 = pi024 & n897;
  assign n946 = pi021 & n895;
  assign n947 = ~n945 & ~n946;
  assign n948 = n944 & n947;
  assign n949 = n311 & ~n948;
  assign n950 = n341 & n558;
  assign n951 = ~n949 & ~n950;
  assign n952 = pi124 & n907;
  assign n953 = pi116 & n910;
  assign n954 = ~n952 & ~n953;
  assign po083 = ~n951 | ~n954;
  assign n956 = pi012 & n902;
  assign n957 = pi023 & n897;
  assign n958 = ~n956 & ~n957;
  assign n959 = pi031 & n900;
  assign n960 = pi020 & n895;
  assign n961 = ~n959 & ~n960;
  assign n962 = n958 & n961;
  assign n963 = n311 & ~n962;
  assign n964 = pi126 & n907;
  assign n965 = pi115 & n910;
  assign n966 = ~n964 & ~n965;
  assign n967 = ~pi004 & pi075;
  assign n968 = pi004 & ~pi075;
  assign n969 = ~n967 & ~n968;
  assign n970 = ~n326 & n969;
  assign n971 = pi001 & n970;
  assign n972 = n341 & n971;
  assign n973 = n966 & ~n972;
  assign po084 = n963 | ~n973;
  assign n975 = pi122 & n907;
  assign n976 = pi112 & n910;
  assign n977 = ~n975 & ~n976;
  assign n978 = pi027 & n897;
  assign n979 = pi008 & n895;
  assign n980 = pi016 & n902;
  assign n981 = ~n979 & ~n980;
  assign n982 = ~n978 & n981;
  assign n983 = pi034 & n900;
  assign n984 = n982 & ~n983;
  assign n985 = n311 & ~n984;
  assign po085 = ~n977 | n985;
  assign n987 = pi123 & n907;
  assign n988 = pi114 & n910;
  assign n989 = ~n987 & ~n988;
  assign n990 = pi022 & n897;
  assign n991 = pi011 & n902;
  assign n992 = ~n990 & ~n991;
  assign n993 = pi030 & n900;
  assign n994 = pi019 & n895;
  assign n995 = ~n993 & ~n994;
  assign n996 = n992 & n995;
  assign n997 = n311 & ~n996;
  assign n998 = ~pi001 & n341;
  assign n999 = n970 & n998;
  assign n1000 = ~n997 & ~n999;
  assign po086 = ~n989 | ~n1000;
  assign n1002 = n916 & n935;
  assign n1003 = pi072 & ~n1002;
  assign n1004 = pi128 & ~n1003;
  assign n1005 = pi146 & n340;
  assign n1006 = n341 & n1005;
  assign po087 = n1004 & ~n1006;
  assign n1008 = pi029 & n897;
  assign n1009 = pi018 & n902;
  assign n1010 = ~n1008 & ~n1009;
  assign n1011 = pi035 & n900;
  assign n1012 = pi010 & n895;
  assign n1013 = ~n1011 & ~n1012;
  assign n1014 = n1010 & n1013;
  assign n1015 = n311 & ~n1014;
  assign n1016 = pi120 & n910;
  assign n1017 = ~n1015 & ~n1016;
  assign n1018 = pi121 & n907;
  assign n1019 = pi003 & n341;
  assign n1020 = ~n1018 & ~n1019;
  assign po088 = ~n1017 | ~n1020;
  assign n1022 = pi125 & n907;
  assign n1023 = pi118 & n910;
  assign n1024 = ~n1022 & ~n1023;
  assign n1025 = pi026 & n897;
  assign n1026 = pi007 & n895;
  assign n1027 = pi015 & n902;
  assign n1028 = ~n1026 & ~n1027;
  assign n1029 = ~n1025 & n1028;
  assign n1030 = pi033 & n900;
  assign n1031 = n1029 & ~n1030;
  assign n1032 = n311 & ~n1031;
  assign po089 = ~n1024 | n1032;
  assign n1034 = ~n895 & ~n902;
  assign n1035 = n315 & ~n1034;
  assign n1036 = pi075 & ~n315;
  assign n1037 = ~n1035 & ~n1036;
  assign po090 = pi128 & ~n1037;
  assign n1039 = ~n660 & ~n667;
  assign n1040 = pi113 & ~n1039;
  assign n1041 = pi076 & ~pi113;
  assign n1042 = ~n1040 & ~n1041;
  assign po091 = pi128 & ~n1042;
  assign n1044 = pi077 & ~n315;
  assign n1045 = ~pi077 & n315;
  assign n1046 = ~n1044 & ~n1045;
  assign po092 = pi128 & ~n1046;
  assign n1048 = pi078 & ~n916;
  assign n1049 = pi144 & n917;
  assign n1050 = pi078 & ~n917;
  assign n1051 = ~n1049 & ~n1050;
  assign n1052 = n916 & ~n1051;
  assign po093 = n1048 | n1052;
  assign n1054 = pi079 & ~n916;
  assign n1055 = pi146 & n918;
  assign n1056 = pi079 & ~n918;
  assign n1057 = ~n1055 & ~n1056;
  assign n1058 = n916 & ~n1057;
  assign po094 = n1054 | n1058;
  assign n1060 = pi080 & ~n916;
  assign n1061 = pi140 & n917;
  assign n1062 = pi080 & ~n917;
  assign n1063 = ~n1061 & ~n1062;
  assign n1064 = n916 & ~n1063;
  assign po095 = n1060 | n1064;
  assign n1066 = pi081 & ~n916;
  assign n1067 = pi144 & n918;
  assign n1068 = pi081 & ~n918;
  assign n1069 = ~n1067 & ~n1068;
  assign n1070 = n916 & ~n1069;
  assign po096 = n1066 | n1070;
  assign n1072 = pi082 & ~n916;
  assign n1073 = n916 & ~n919;
  assign n1074 = ~n1072 & ~n1073;
  assign po097 = pi128 & ~n1074;
  assign n1076 = pi083 & ~n916;
  assign n1077 = ~pi083 & n916;
  assign n1078 = ~n1076 & ~n1077;
  assign po098 = pi128 & ~n1078;
  assign n1080 = pi084 & ~n916;
  assign n1081 = pi140 & n918;
  assign n1082 = pi084 & ~n918;
  assign n1083 = ~n1081 & ~n1082;
  assign n1084 = n916 & ~n1083;
  assign po099 = n1080 | n1084;
  assign n1086 = pi085 & ~n916;
  assign n1087 = pi141 & n918;
  assign n1088 = pi085 & ~n918;
  assign n1089 = ~n1087 & ~n1088;
  assign n1090 = n916 & ~n1089;
  assign po100 = n1086 | n1090;
  assign n1092 = pi086 & ~n916;
  assign n1093 = pi142 & n918;
  assign n1094 = pi086 & ~n918;
  assign n1095 = ~n1093 & ~n1094;
  assign n1096 = n916 & ~n1095;
  assign po101 = n1092 | n1096;
  assign n1098 = pi087 & ~n916;
  assign n1099 = pi143 & n918;
  assign n1100 = pi087 & ~n918;
  assign n1101 = ~n1099 & ~n1100;
  assign n1102 = n916 & ~n1101;
  assign po102 = n1098 | n1102;
  assign n1104 = pi088 & ~n916;
  assign n1105 = pi145 & n918;
  assign n1106 = pi088 & ~n918;
  assign n1107 = ~n1105 & ~n1106;
  assign n1108 = n916 & ~n1107;
  assign po103 = n1104 | n1108;
  assign n1110 = pi089 & ~n916;
  assign n1111 = pi147 & n918;
  assign n1112 = pi089 & ~n918;
  assign n1113 = ~n1111 & ~n1112;
  assign n1114 = n916 & ~n1113;
  assign po104 = n1110 | n1114;
  assign n1116 = pi090 & ~n916;
  assign n1117 = pi141 & n917;
  assign n1118 = pi090 & ~n917;
  assign n1119 = ~n1117 & ~n1118;
  assign n1120 = n916 & ~n1119;
  assign po105 = n1116 | n1120;
  assign n1122 = pi091 & ~n916;
  assign n1123 = pi142 & n917;
  assign n1124 = pi091 & ~n917;
  assign n1125 = ~n1123 & ~n1124;
  assign n1126 = n916 & ~n1125;
  assign po106 = n1122 | n1126;
  assign n1128 = pi092 & ~n916;
  assign n1129 = pi143 & n917;
  assign n1130 = pi092 & ~n917;
  assign n1131 = ~n1129 & ~n1130;
  assign n1132 = n916 & ~n1131;
  assign po107 = n1128 | n1132;
  assign n1134 = pi093 & ~n916;
  assign n1135 = pi145 & n917;
  assign n1136 = pi093 & ~n917;
  assign n1137 = ~n1135 & ~n1136;
  assign n1138 = n916 & ~n1137;
  assign po108 = n1134 | n1138;
  assign n1140 = pi094 & ~n916;
  assign n1141 = pi146 & n917;
  assign n1142 = pi094 & ~n917;
  assign n1143 = ~n1141 & ~n1142;
  assign n1144 = n916 & ~n1143;
  assign po109 = n1140 | n1144;
  assign n1146 = pi095 & ~n916;
  assign n1147 = pi147 & n917;
  assign n1148 = pi095 & ~n917;
  assign n1149 = ~n1147 & ~n1148;
  assign n1150 = n916 & ~n1149;
  assign po110 = n1146 | n1150;
  assign n1152 = pi096 & ~n916;
  assign n1153 = ~pi082 & ~pi083;
  assign n1154 = pi096 & ~n1153;
  assign n1155 = pi144 & n1153;
  assign n1156 = ~n1154 & ~n1155;
  assign n1157 = n916 & ~n1156;
  assign po111 = n1152 | n1157;
  assign n1159 = pi097 & ~n916;
  assign n1160 = pi082 & pi083;
  assign n1161 = pi144 & n1160;
  assign n1162 = pi097 & ~n1160;
  assign n1163 = ~n1161 & ~n1162;
  assign n1164 = n916 & ~n1163;
  assign po112 = n1159 | n1164;
  assign n1166 = pi098 & ~n916;
  assign n1167 = pi140 & n1160;
  assign n1168 = pi098 & ~n1160;
  assign n1169 = ~n1167 & ~n1168;
  assign n1170 = n916 & ~n1169;
  assign po113 = n1166 | n1170;
  assign n1172 = pi099 & ~n916;
  assign n1173 = pi099 & ~n1153;
  assign n1174 = pi147 & n1153;
  assign n1175 = ~n1173 & ~n1174;
  assign n1176 = n916 & ~n1175;
  assign po114 = n1172 | n1176;
  assign n1178 = pi100 & ~n916;
  assign n1179 = pi100 & ~n1153;
  assign n1180 = pi140 & n1153;
  assign n1181 = ~n1179 & ~n1180;
  assign n1182 = n916 & ~n1181;
  assign po115 = n1178 | n1182;
  assign n1184 = pi101 & ~n916;
  assign n1185 = pi101 & ~n1153;
  assign n1186 = pi141 & n1153;
  assign n1187 = ~n1185 & ~n1186;
  assign n1188 = n916 & ~n1187;
  assign po116 = n1184 | n1188;
  assign n1190 = pi102 & ~n916;
  assign n1191 = pi102 & ~n1153;
  assign n1192 = pi142 & n1153;
  assign n1193 = ~n1191 & ~n1192;
  assign n1194 = n916 & ~n1193;
  assign po117 = n1190 | n1194;
  assign n1196 = pi103 & ~n916;
  assign n1197 = pi103 & ~n1153;
  assign n1198 = pi143 & n1153;
  assign n1199 = ~n1197 & ~n1198;
  assign n1200 = n916 & ~n1199;
  assign po118 = n1196 | n1200;
  assign n1202 = pi104 & ~n916;
  assign n1203 = pi104 & ~n1153;
  assign n1204 = pi146 & n1153;
  assign n1205 = ~n1203 & ~n1204;
  assign n1206 = n916 & ~n1205;
  assign po119 = n1202 | n1206;
  assign n1208 = pi105 & ~n916;
  assign n1209 = pi105 & ~n1153;
  assign n1210 = pi145 & n1153;
  assign n1211 = ~n1209 & ~n1210;
  assign n1212 = n916 & ~n1211;
  assign po120 = n1208 | n1212;
  assign n1214 = pi106 & ~n916;
  assign n1215 = pi141 & n1160;
  assign n1216 = pi106 & ~n1160;
  assign n1217 = ~n1215 & ~n1216;
  assign n1218 = n916 & ~n1217;
  assign po121 = n1214 | n1218;
  assign n1220 = pi107 & ~n916;
  assign n1221 = pi142 & n1160;
  assign n1222 = pi107 & ~n1160;
  assign n1223 = ~n1221 & ~n1222;
  assign n1224 = n916 & ~n1223;
  assign po122 = n1220 | n1224;
  assign n1226 = pi108 & ~n916;
  assign n1227 = pi143 & n1160;
  assign n1228 = pi108 & ~n1160;
  assign n1229 = ~n1227 & ~n1228;
  assign n1230 = n916 & ~n1229;
  assign po123 = n1226 | n1230;
  assign n1232 = pi109 & ~n916;
  assign n1233 = pi145 & n1160;
  assign n1234 = pi109 & ~n1160;
  assign n1235 = ~n1233 & ~n1234;
  assign n1236 = n916 & ~n1235;
  assign po124 = n1232 | n1236;
  assign n1238 = pi110 & ~n916;
  assign n1239 = pi146 & n1160;
  assign n1240 = pi110 & ~n1160;
  assign n1241 = ~n1239 & ~n1240;
  assign n1242 = n916 & ~n1241;
  assign po125 = n1238 | n1242;
  assign n1244 = pi111 & ~n916;
  assign n1245 = pi147 & n1160;
  assign n1246 = pi111 & ~n1160;
  assign n1247 = ~n1245 & ~n1246;
  assign n1248 = n916 & ~n1247;
  assign po126 = n1244 | n1248;
  assign n1250 = pi112 & ~n910;
  assign n1251 = pi145 & n910;
  assign n1252 = ~n1250 & ~n1251;
  assign n1253 = n340 & ~n1252;
  assign n1254 = pi112 & ~n340;
  assign po127 = n1253 | n1254;
  assign n1256 = pi128 & n567;
  assign po128 = ~n558 & n1256;
  assign n1258 = pi114 & ~n910;
  assign n1259 = pi140 & n910;
  assign n1260 = ~n1258 & ~n1259;
  assign n1261 = n340 & ~n1260;
  assign n1262 = pi114 & ~n340;
  assign po129 = n1261 | n1262;
  assign n1264 = pi115 & ~n910;
  assign n1265 = pi141 & n910;
  assign n1266 = ~n1264 & ~n1265;
  assign n1267 = n340 & ~n1266;
  assign n1268 = pi115 & ~n340;
  assign po130 = n1267 | n1268;
  assign n1270 = pi116 & ~n910;
  assign n1271 = pi142 & n910;
  assign n1272 = ~n1270 & ~n1271;
  assign n1273 = n340 & ~n1272;
  assign n1274 = pi116 & ~n340;
  assign po131 = n1273 | n1274;
  assign n1276 = pi117 & ~n910;
  assign n1277 = pi143 & n910;
  assign n1278 = ~n1276 & ~n1277;
  assign n1279 = n340 & ~n1278;
  assign n1280 = pi117 & ~n340;
  assign po132 = n1279 | n1280;
  assign n1282 = pi118 & ~n910;
  assign n1283 = pi144 & n910;
  assign n1284 = ~n1282 & ~n1283;
  assign n1285 = n340 & ~n1284;
  assign n1286 = pi118 & ~n340;
  assign po133 = n1285 | n1286;
  assign n1288 = pi119 & ~n910;
  assign n1289 = pi146 & n910;
  assign n1290 = ~n1288 & ~n1289;
  assign n1291 = n340 & ~n1290;
  assign n1292 = pi119 & ~n340;
  assign po134 = n1291 | n1292;
  assign n1294 = pi120 & ~n910;
  assign n1295 = pi147 & n910;
  assign n1296 = ~n1294 & ~n1295;
  assign n1297 = n340 & ~n1296;
  assign n1298 = pi120 & ~n340;
  assign po135 = n1297 | n1298;
  assign n1300 = pi121 & ~n907;
  assign n1301 = pi147 & n907;
  assign n1302 = ~n1300 & ~n1301;
  assign n1303 = n340 & ~n1302;
  assign n1304 = pi121 & ~n340;
  assign po136 = n1303 | n1304;
  assign n1306 = pi122 & ~n907;
  assign n1307 = pi145 & n907;
  assign n1308 = ~n1306 & ~n1307;
  assign n1309 = n340 & ~n1308;
  assign n1310 = pi122 & ~n340;
  assign po137 = n1309 | n1310;
  assign n1312 = pi140 & n907;
  assign n1313 = pi123 & ~n907;
  assign n1314 = ~n1312 & ~n1313;
  assign n1315 = n340 & ~n1314;
  assign n1316 = pi123 & ~n340;
  assign po138 = n1315 | n1316;
  assign n1318 = pi124 & ~n907;
  assign n1319 = pi142 & n907;
  assign n1320 = ~n1318 & ~n1319;
  assign n1321 = n340 & ~n1320;
  assign n1322 = pi124 & ~n340;
  assign po139 = n1321 | n1322;
  assign n1324 = n340 & n907;
  assign po140 = pi125 | n1324;
  assign n1326 = pi126 & ~n907;
  assign n1327 = pi141 & n907;
  assign n1328 = ~n1326 & ~n1327;
  assign n1329 = n340 & ~n1328;
  assign n1330 = pi126 & ~n340;
  assign po141 = n1329 | n1330;
  assign n1332 = pi127 & ~n907;
  assign n1333 = pi143 & n907;
  assign n1334 = ~n1332 & ~n1333;
  assign n1335 = n340 & ~n1334;
  assign n1336 = pi127 & ~n340;
  assign po142 = n1335 | n1336;
  assign n1338 = pi146 & n907;
  assign n1339 = pi128 & ~n907;
  assign n1340 = ~n1338 & ~n1339;
  assign n1341 = n340 & ~n1340;
  assign n1342 = pi128 & ~n340;
  assign po143 = n1341 | n1342;
  assign n1344 = pi113 & ~pi129;
  assign n1345 = ~pi113 & pi129;
  assign n1346 = ~n1344 & ~n1345;
  assign po144 = pi128 & ~n1346;
  assign po145 = ~pi130 & n313;
  assign po146 = pi003 & pi121;
  assign po012 = 1'b1;
  assign po000 = pi071;
  assign po001 = pi069;
  assign po002 = pi068;
  assign po003 = pi067;
  assign po004 = pi074;
  assign po005 = pi070;
  assign po006 = pi065;
  assign po007 = pi073;
  assign po008 = pi130;
  assign po009 = pi131;
  assign po010 = pi038;
  assign po011 = pi043;
  assign po013 = pi132;
  assign po018 = pi133;
endmodule


