// Benchmark "div16" written by ABC on Wed Apr 29 17:28:58 2015

module div16 ( 
    pi00, pi01, pi02, pi03, pi04, pi05, pi06, pi07, pi08, pi09, pi10, pi11,
    pi12, pi13, pi14, pi15, pi16, pi17, pi18, pi19, pi20, pi21, pi22, pi23,
    pi24, pi25, pi26, pi27, pi28, pi29, pi30, pi31,
    po00, po01, po02, po03, po04, po05, po06, po07, po08, po09, po10, po11,
    po12, po13, po14, po15, po16, po17, po18, po19, po20, po21, po22, po23,
    po24, po25, po26, po27, po28, po29, po30, po31  );
  input  pi00, pi01, pi02, pi03, pi04, pi05, pi06, pi07, pi08, pi09,
    pi10, pi11, pi12, pi13, pi14, pi15, pi16, pi17, pi18, pi19, pi20, pi21,
    pi22, pi23, pi24, pi25, pi26, pi27, pi28, pi29, pi30, pi31;
  output po00, po01, po02, po03, po04, po05, po06, po07, po08, po09, po10,
    po11, po12, po13, po14, po15, po16, po17, po18, po19, po20, po21, po22,
    po23, po24, po25, po26, po27, po28, po29, po30, po31;
  wire n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78,
    n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92,
    n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105,
    n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116, n117,
    n118, n119, n120, n121, n122, n123, n124, n125, n126, n127, n128, n129,
    n130, n131, n132, n133, n134, n135, n136, n137, n138, n139, n140, n141,
    n142, n143, n144, n145, n146, n147, n148, n149, n150, n151, n152, n153,
    n154, n155, n156, n157, n158, n159, n160, n161, n162, n163, n164, n165,
    n166, n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
    n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188, n189,
    n190, n191, n192, n193, n194, n195, n196, n197, n198, n199, n200, n201,
    n202, n203, n204, n205, n206, n207, n208, n209, n210, n211, n212, n213,
    n214, n215, n216, n217, n218, n219, n220, n221, n222, n223, n224, n225,
    n226, n227, n228, n229, n230, n231, n232, n233, n234, n235, n236, n237,
    n238, n239, n240, n241, n242, n243, n244, n245, n246, n247, n248, n249,
    n250, n251, n252, n253, n254, n255, n256, n257, n258, n259, n260, n261,
    n262, n263, n264, n265, n266, n267, n268, n269, n270, n271, n272, n273,
    n274, n275, n276, n277, n278, n279, n280, n281, n282, n283, n284, n285,
    n286, n287, n288, n289, n290, n291, n292, n293, n294, n295, n296, n297,
    n298, n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
    n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320, n321,
    n322, n323, n324, n325, n326, n327, n328, n329, n330, n331, n332, n333,
    n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345,
    n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357,
    n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369,
    n371, n373, n374, n375, n376, n377, n378, n379, n380, n381, n382, n383,
    n384, n385, n386, n387, n388, n389, n390, n391, n392, n393, n394, n395,
    n396, n397, n398, n399, n400, n401, n402, n403, n404, n405, n406, n407,
    n408, n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
    n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431,
    n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443,
    n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455,
    n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467,
    n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, n479,
    n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, n490, n491,
    n492, n493, n494, n495, n496, n497, n498, n499, n500, n501, n502, n503,
    n504, n505, n506, n507, n508, n509, n510, n511, n512, n513, n514, n515,
    n516, n517, n518, n519, n520, n521, n522, n523, n524, n525, n526, n527,
    n528, n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539,
    n540, n541, n542, n543, n544, n545, n546, n547, n548, n550, n551, n552,
    n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
    n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
    n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588,
    n589, n590, n591, n592, n593, n594, n595, n596, n597, n598, n599, n600,
    n601, n602, n603, n604, n605, n606, n607, n608, n609, n610, n611, n612,
    n613, n614, n615, n616, n617, n618, n619, n620, n621, n622, n623, n624,
    n625, n626, n627, n628, n629, n630, n631, n632, n633, n634, n635, n636,
    n637, n638, n639, n640, n641, n642, n643, n644, n645, n646, n647, n648,
    n649, n650, n651, n652, n653, n654, n655, n656, n657, n658, n659, n660,
    n661, n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
    n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684,
    n685, n686, n687, n688, n689, n690, n691, n692, n693, n694, n695, n696,
    n697, n698, n699, n700, n701, n702, n703, n704, n705, n706, n707, n708,
    n709, n710, n711, n712, n713, n714, n715, n716, n717, n718, n719, n720,
    n721, n722, n723, n724, n725, n726, n727, n728, n729, n730, n731, n732,
    n733, n734, n735, n736, n737, n738, n739, n740, n741, n742, n743, n744,
    n746, n747, n748, n749, n750, n751, n752, n753, n754, n755, n756, n757,
    n758, n759, n760, n761, n762, n763, n764, n765, n766, n767, n768, n769,
    n770, n771, n772, n773, n774, n775, n776, n777, n778, n779, n780, n781,
    n782, n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793,
    n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804, n805,
    n806, n807, n808, n809, n810, n811, n812, n813, n814, n815, n816, n817,
    n818, n819, n820, n821, n822, n823, n824, n825, n826, n827, n828, n829,
    n830, n831, n832, n833, n834, n835, n836, n837, n838, n839, n840, n841,
    n842, n843, n844, n845, n846, n847, n848, n849, n850, n851, n852, n853,
    n854, n855, n856, n857, n858, n859, n860, n861, n862, n863, n864, n865,
    n866, n867, n868, n869, n870, n871, n872, n873, n874, n875, n876, n877,
    n878, n879, n880, n881, n882, n883, n884, n885, n886, n887, n888, n889,
    n890, n891, n892, n893, n894, n895, n896, n897, n898, n899, n900, n901,
    n902, n903, n904, n905, n906, n907, n908, n909, n910, n911, n912, n913,
    n914, n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925,
    n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936, n937,
    n938, n939, n940, n941, n942, n943, n944, n945, n946, n947, n948, n949,
    n950, n951, n952, n953, n954, n955, n956, n957, n958, n959, n960, n961,
    n962, n963, n964, n965, n966, n967, n968, n969, n970, n971, n972, n973,
    n974, n975, n976, n977, n979, n980, n981, n982, n983, n984, n985, n986,
    n987, n988, n989, n990, n991, n992, n993, n994, n995, n996, n997, n998,
    n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008,
    n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018,
    n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028,
    n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038,
    n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048,
    n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058,
    n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068,
    n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078,
    n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088,
    n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098,
    n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108,
    n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118,
    n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128,
    n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138,
    n1139, n1140, n1141, n1142, n1143, n1145, n1146, n1147, n1148, n1149,
    n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159,
    n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169,
    n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179,
    n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189,
    n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199,
    n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209,
    n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219,
    n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229,
    n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239,
    n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249,
    n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259,
    n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269,
    n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279,
    n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289,
    n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299,
    n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309,
    n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319,
    n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329,
    n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339,
    n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349,
    n1350, n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1358, n1359,
    n1360, n1361, n1362, n1363, n1364, n1365, n1366, n1367, n1368, n1369,
    n1370, n1371, n1372, n1373, n1374, n1375, n1376, n1377, n1378, n1379,
    n1380, n1381, n1382, n1383, n1384, n1385, n1386, n1387, n1388, n1389,
    n1390, n1391, n1392, n1393, n1394, n1395, n1396, n1397, n1398, n1399,
    n1400, n1401, n1402, n1403, n1404, n1405, n1406, n1407, n1408, n1409,
    n1410, n1411, n1412, n1413, n1414, n1415, n1416, n1417, n1418, n1419,
    n1420, n1421, n1422, n1423, n1424, n1425, n1426, n1427, n1428, n1429,
    n1430, n1432, n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440,
    n1441, n1442, n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450,
    n1451, n1452, n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460,
    n1461, n1462, n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470,
    n1471, n1472, n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480,
    n1481, n1482, n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1490,
    n1491, n1492, n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500,
    n1501, n1502, n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510,
    n1511, n1512, n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1520,
    n1521, n1522, n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530,
    n1531, n1532, n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540,
    n1541, n1542, n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550,
    n1551, n1552, n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560,
    n1561, n1562, n1563, n1564, n1565, n1566, n1567, n1568, n1569, n1570,
    n1571, n1572, n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1580,
    n1581, n1582, n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590,
    n1591, n1592, n1593, n1594, n1595, n1596, n1597, n1598, n1599, n1600,
    n1601, n1602, n1603, n1604, n1605, n1606, n1607, n1608, n1609, n1610,
    n1611, n1612, n1613, n1614, n1615, n1616, n1617, n1618, n1619, n1620,
    n1621, n1622, n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630,
    n1631, n1632, n1633, n1634, n1635, n1636, n1637, n1638, n1639, n1640,
    n1641, n1642, n1643, n1644, n1645, n1646, n1647, n1648, n1649, n1650,
    n1651, n1652, n1653, n1654, n1655, n1656, n1657, n1658, n1659, n1660,
    n1661, n1662, n1663, n1664, n1665, n1666, n1667, n1668, n1669, n1670,
    n1671, n1672, n1673, n1674, n1675, n1676, n1677, n1678, n1679, n1680,
    n1681, n1682, n1683, n1684, n1685, n1686, n1687, n1688, n1689, n1690,
    n1691, n1692, n1693, n1694, n1695, n1696, n1697, n1698, n1699, n1700,
    n1701, n1702, n1703, n1704, n1705, n1706, n1707, n1708, n1709, n1710,
    n1711, n1712, n1713, n1714, n1715, n1716, n1717, n1718, n1719, n1720,
    n1721, n1722, n1723, n1724, n1725, n1726, n1727, n1728, n1729, n1730,
    n1731, n1732, n1733, n1734, n1735, n1736, n1737, n1738, n1739, n1740,
    n1741, n1742, n1743, n1744, n1745, n1746, n1747, n1748, n1749, n1750,
    n1751, n1752, n1753, n1754, n1755, n1756, n1757, n1758, n1759, n1760,
    n1761, n1762, n1763, n1764, n1765, n1766, n1767, n1768, n1769, n1770,
    n1771, n1772, n1773, n1774, n1775, n1776, n1777, n1778, n1779, n1780,
    n1781, n1782, n1783, n1784, n1785, n1786, n1787, n1788, n1789, n1790,
    n1791, n1792, n1793, n1794, n1795, n1796, n1797, n1798, n1799, n1800,
    n1801, n1802, n1803, n1804, n1805, n1806, n1807, n1808, n1809, n1810,
    n1811, n1812, n1813, n1814, n1815, n1816, n1817, n1818, n1819, n1820,
    n1821, n1822, n1823, n1824, n1825, n1826, n1827, n1828, n1830, n1831,
    n1832, n1833, n1834, n1835, n1836, n1837, n1838, n1839, n1840, n1841,
    n1842, n1843, n1844, n1845, n1846, n1847, n1848, n1849, n1850, n1851,
    n1852, n1853, n1854, n1855, n1856, n1857, n1858, n1859, n1860, n1861,
    n1862, n1863, n1864, n1865, n1866, n1867, n1868, n1869, n1870, n1871,
    n1872, n1873, n1874, n1875, n1876, n1877, n1878, n1879, n1880, n1881,
    n1882, n1883, n1884, n1885, n1886, n1887, n1888, n1889, n1890, n1891,
    n1892, n1893, n1894, n1895, n1896, n1897, n1898, n1899, n1900, n1901,
    n1902, n1903, n1904, n1905, n1906, n1907, n1908, n1909, n1910, n1911,
    n1912, n1913, n1914, n1915, n1916, n1917, n1918, n1919, n1920, n1921,
    n1922, n1923, n1924, n1925, n1926, n1927, n1928, n1929, n1930, n1931,
    n1932, n1933, n1934, n1935, n1936, n1937, n1938, n1939, n1940, n1941,
    n1942, n1943, n1944, n1945, n1946, n1947, n1948, n1949, n1950, n1951,
    n1952, n1953, n1954, n1955, n1956, n1957, n1958, n1959, n1960, n1961,
    n1962, n1963, n1964, n1965, n1966, n1967, n1968, n1969, n1970, n1971,
    n1972, n1973, n1974, n1975, n1976, n1977, n1978, n1979, n1980, n1981,
    n1982, n1983, n1984, n1985, n1986, n1987, n1988, n1989, n1990, n1991,
    n1992, n1993, n1994, n1995, n1996, n1997, n1998, n1999, n2000, n2001,
    n2002, n2003, n2004, n2005, n2006, n2007, n2008, n2009, n2010, n2011,
    n2012, n2013, n2014, n2015, n2016, n2017, n2018, n2019, n2020, n2021,
    n2022, n2023, n2024, n2025, n2026, n2027, n2028, n2029, n2030, n2031,
    n2032, n2033, n2034, n2035, n2036, n2037, n2038, n2039, n2040, n2041,
    n2042, n2043, n2044, n2045, n2046, n2047, n2048, n2049, n2050, n2051,
    n2052, n2053, n2054, n2055, n2056, n2057, n2058, n2059, n2060, n2061,
    n2062, n2063, n2064, n2065, n2066, n2067, n2068, n2069, n2070, n2071,
    n2072, n2073, n2074, n2075, n2076, n2077, n2078, n2079, n2080, n2081,
    n2082, n2083, n2084, n2085, n2086, n2087, n2088, n2089, n2090, n2091,
    n2092, n2093, n2094, n2095, n2096, n2097, n2098, n2099, n2100, n2102,
    n2103, n2104, n2105, n2106, n2107, n2108, n2109, n2110, n2111, n2112,
    n2113, n2114, n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122,
    n2123, n2124, n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132,
    n2133, n2134, n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142,
    n2143, n2144, n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152,
    n2153, n2154, n2155, n2156, n2157, n2158, n2159, n2160, n2161, n2162,
    n2163, n2164, n2165, n2166, n2167, n2168, n2169, n2170, n2171, n2172,
    n2173, n2174, n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2182,
    n2183, n2184, n2185, n2186, n2187, n2188, n2189, n2190, n2191, n2192,
    n2193, n2194, n2195, n2196, n2197, n2198, n2199, n2200, n2201, n2202,
    n2203, n2204, n2205, n2206, n2207, n2208, n2209, n2210, n2211, n2212,
    n2213, n2214, n2215, n2216, n2217, n2218, n2219, n2220, n2221, n2222,
    n2223, n2224, n2225, n2226, n2227, n2228, n2229, n2230, n2231, n2232,
    n2233, n2234, n2235, n2236, n2237, n2238, n2239, n2240, n2241, n2242,
    n2243, n2244, n2245, n2246, n2247, n2248, n2249, n2250, n2251, n2252,
    n2253, n2254, n2255, n2256, n2257, n2258, n2259, n2260, n2261, n2262,
    n2263, n2264, n2265, n2266, n2267, n2268, n2269, n2270, n2271, n2272,
    n2273, n2274, n2275, n2276, n2277, n2278, n2279, n2280, n2281, n2282,
    n2283, n2284, n2285, n2286, n2287, n2288, n2289, n2290, n2291, n2292,
    n2293, n2294, n2295, n2296, n2297, n2298, n2299, n2300, n2301, n2302,
    n2303, n2304, n2305, n2306, n2307, n2308, n2309, n2310, n2311, n2312,
    n2313, n2314, n2315, n2316, n2317, n2318, n2319, n2320, n2321, n2322,
    n2323, n2324, n2325, n2326, n2327, n2328, n2329, n2330, n2331, n2332,
    n2333, n2334, n2335, n2336, n2337, n2338, n2339, n2340, n2341, n2342,
    n2343, n2344, n2345, n2346, n2347, n2348, n2349, n2350, n2351, n2352,
    n2353, n2354, n2355, n2356, n2357, n2358, n2359, n2360, n2361, n2362,
    n2363, n2364, n2365, n2366, n2367, n2368, n2369, n2370, n2371, n2372,
    n2373, n2374, n2375, n2376, n2377, n2378, n2379, n2380, n2381, n2382,
    n2383, n2384, n2385, n2386, n2387, n2388, n2389, n2390, n2391, n2392,
    n2393, n2394, n2395, n2396, n2397, n2398, n2399, n2400, n2401, n2402,
    n2403, n2404, n2405, n2406, n2407, n2408, n2409, n2410, n2411, n2412,
    n2413, n2414, n2415, n2416, n2417, n2418, n2419, n2420, n2421, n2422,
    n2423, n2424, n2425, n2426, n2427, n2428, n2429, n2430, n2431, n2432,
    n2433, n2434, n2435, n2436, n2437, n2438, n2439, n2440, n2441, n2442,
    n2443, n2444, n2445, n2446, n2447, n2448, n2449, n2450, n2451, n2452,
    n2453, n2454, n2455, n2456, n2457, n2458, n2459, n2461, n2462, n2463,
    n2464, n2465, n2466, n2467, n2468, n2469, n2470, n2471, n2472, n2473,
    n2474, n2475, n2476, n2477, n2478, n2479, n2480, n2481, n2482, n2483,
    n2484, n2485, n2486, n2487, n2488, n2489, n2490, n2491, n2492, n2493,
    n2494, n2495, n2496, n2497, n2498, n2499, n2500, n2501, n2502, n2503,
    n2504, n2505, n2506, n2507, n2508, n2509, n2510, n2511, n2512, n2513,
    n2514, n2515, n2516, n2517, n2518, n2519, n2520, n2521, n2522, n2523,
    n2524, n2525, n2526, n2527, n2528, n2529, n2530, n2531, n2532, n2533,
    n2534, n2535, n2536, n2537, n2538, n2539, n2540, n2541, n2542, n2543,
    n2544, n2545, n2546, n2547, n2548, n2549, n2550, n2551, n2552, n2553,
    n2554, n2555, n2556, n2557, n2558, n2559, n2560, n2561, n2562, n2563,
    n2564, n2565, n2566, n2567, n2568, n2569, n2570, n2571, n2572, n2573,
    n2574, n2575, n2576, n2577, n2578, n2579, n2580, n2581, n2582, n2583,
    n2584, n2585, n2586, n2587, n2588, n2589, n2590, n2591, n2592, n2593,
    n2594, n2595, n2596, n2597, n2598, n2599, n2600, n2601, n2602, n2603,
    n2604, n2605, n2606, n2607, n2608, n2609, n2610, n2611, n2612, n2613,
    n2614, n2615, n2616, n2617, n2618, n2619, n2620, n2621, n2622, n2623,
    n2624, n2625, n2626, n2627, n2628, n2629, n2630, n2631, n2632, n2633,
    n2634, n2635, n2636, n2637, n2638, n2639, n2640, n2641, n2642, n2643,
    n2644, n2645, n2646, n2647, n2648, n2649, n2650, n2651, n2652, n2653,
    n2654, n2655, n2656, n2657, n2658, n2659, n2660, n2661, n2662, n2663,
    n2664, n2665, n2666, n2667, n2668, n2669, n2670, n2671, n2672, n2673,
    n2674, n2675, n2676, n2677, n2678, n2679, n2680, n2681, n2682, n2683,
    n2684, n2685, n2686, n2687, n2688, n2689, n2690, n2691, n2692, n2693,
    n2694, n2695, n2696, n2697, n2698, n2699, n2700, n2701, n2702, n2703,
    n2704, n2705, n2706, n2707, n2708, n2709, n2710, n2711, n2712, n2713,
    n2714, n2715, n2716, n2717, n2718, n2719, n2720, n2721, n2722, n2723,
    n2724, n2725, n2726, n2727, n2728, n2729, n2730, n2731, n2732, n2733,
    n2734, n2735, n2736, n2737, n2738, n2739, n2740, n2741, n2742, n2743,
    n2744, n2745, n2746, n2747, n2748, n2749, n2750, n2751, n2752, n2753,
    n2754, n2755, n2756, n2757, n2758, n2759, n2760, n2761, n2762, n2763,
    n2764, n2765, n2766, n2767, n2768, n2769, n2770, n2771, n2772, n2773,
    n2774, n2775, n2776, n2777, n2778, n2779, n2780, n2781, n2782, n2783,
    n2784, n2785, n2786, n2787, n2788, n2789, n2790, n2791, n2792, n2793,
    n2794, n2795, n2796, n2797, n2798, n2799, n2800, n2801, n2802, n2803,
    n2804, n2805, n2806, n2807, n2808, n2809, n2810, n2811, n2812, n2813,
    n2814, n2815, n2816, n2817, n2818, n2819, n2820, n2821, n2822, n2823,
    n2824, n2825, n2826, n2827, n2828, n2829, n2830, n2831, n2832, n2833,
    n2834, n2835, n2836, n2837, n2838, n2839, n2840, n2841, n2842, n2843,
    n2844, n2845, n2846, n2847, n2848, n2849, n2850, n2851, n2852, n2853,
    n2854, n2855, n2856, n2857, n2858, n2859, n2860, n2861, n2862, n2863,
    n2864, n2865, n2866, n2867, n2868, n2869, n2870, n2871, n2872, n2873,
    n2874, n2875, n2876, n2877, n2878, n2879, n2880, n2881, n2882, n2883,
    n2884, n2885, n2886, n2887, n2888, n2889, n2890, n2891, n2892, n2893,
    n2894, n2895, n2896, n2897, n2898, n2899, n2900, n2901, n2902, n2903,
    n2904, n2905, n2906, n2907, n2908, n2909, n2910, n2911, n2912, n2913,
    n2914, n2915, n2916, n2917, n2918, n2920, n2921, n2922, n2923, n2924,
    n2925, n2926, n2927, n2928, n2929, n2930, n2931, n2932, n2933, n2934,
    n2935, n2936, n2937, n2938, n2939, n2940, n2941, n2942, n2943, n2944,
    n2945, n2946, n2947, n2948, n2949, n2950, n2951, n2952, n2953, n2954,
    n2955, n2956, n2957, n2958, n2959, n2960, n2961, n2962, n2963, n2964,
    n2965, n2966, n2967, n2968, n2969, n2970, n2971, n2972, n2973, n2974,
    n2975, n2976, n2977, n2978, n2979, n2980, n2981, n2982, n2983, n2984,
    n2985, n2986, n2987, n2988, n2989, n2990, n2991, n2992, n2993, n2994,
    n2995, n2996, n2997, n2998, n2999, n3000, n3001, n3002, n3003, n3004,
    n3005, n3006, n3007, n3008, n3009, n3010, n3011, n3012, n3013, n3014,
    n3015, n3016, n3017, n3018, n3019, n3020, n3021, n3022, n3023, n3024,
    n3025, n3026, n3027, n3028, n3029, n3030, n3031, n3032, n3033, n3034,
    n3035, n3036, n3037, n3038, n3039, n3040, n3041, n3042, n3043, n3044,
    n3045, n3046, n3047, n3048, n3049, n3050, n3051, n3052, n3053, n3054,
    n3055, n3056, n3057, n3058, n3059, n3060, n3061, n3062, n3063, n3064,
    n3065, n3066, n3067, n3068, n3069, n3070, n3071, n3072, n3073, n3074,
    n3075, n3076, n3077, n3078, n3079, n3080, n3081, n3082, n3083, n3084,
    n3085, n3086, n3087, n3088, n3089, n3090, n3091, n3092, n3093, n3094,
    n3095, n3096, n3097, n3098, n3099, n3100, n3101, n3102, n3103, n3104,
    n3105, n3106, n3107, n3108, n3109, n3110, n3111, n3112, n3113, n3114,
    n3115, n3116, n3117, n3118, n3119, n3120, n3121, n3122, n3123, n3124,
    n3125, n3126, n3127, n3128, n3129, n3130, n3131, n3132, n3133, n3134,
    n3135, n3136, n3137, n3138, n3139, n3140, n3141, n3142, n3143, n3144,
    n3145, n3146, n3147, n3148, n3149, n3150, n3151, n3152, n3153, n3154,
    n3155, n3156, n3157, n3158, n3159, n3160, n3161, n3162, n3163, n3164,
    n3165, n3166, n3167, n3168, n3169, n3170, n3171, n3172, n3173, n3174,
    n3175, n3176, n3177, n3178, n3179, n3180, n3181, n3182, n3183, n3184,
    n3185, n3186, n3187, n3188, n3189, n3190, n3191, n3192, n3193, n3194,
    n3195, n3196, n3197, n3198, n3199, n3200, n3201, n3202, n3203, n3204,
    n3205, n3206, n3207, n3208, n3209, n3210, n3211, n3212, n3213, n3214,
    n3215, n3216, n3217, n3218, n3219, n3220, n3221, n3222, n3223, n3224,
    n3225, n3226, n3227, n3228, n3229, n3230, n3231, n3232, n3233, n3234,
    n3235, n3236, n3237, n3238, n3239, n3240, n3241, n3242, n3243, n3244,
    n3245, n3246, n3247, n3248, n3249, n3250, n3251, n3252, n3253, n3254,
    n3255, n3256, n3257, n3258, n3259, n3260, n3261, n3262, n3263, n3264,
    n3265, n3266, n3267, n3268, n3269, n3270, n3271, n3272, n3273, n3274,
    n3275, n3276, n3277, n3278, n3279, n3280, n3281, n3282, n3283, n3284,
    n3285, n3286, n3287, n3288, n3289, n3290, n3291, n3292, n3293, n3294,
    n3295, n3296, n3297, n3298, n3299, n3300, n3301, n3302, n3303, n3304,
    n3305, n3306, n3307, n3308, n3309, n3310, n3311, n3312, n3313, n3314,
    n3315, n3316, n3317, n3318, n3319, n3320, n3321, n3322, n3323, n3324,
    n3325, n3326, n3327, n3328, n3329, n3330, n3331, n3332, n3333, n3334,
    n3335, n3336, n3337, n3338, n3339, n3340, n3341, n3342, n3343, n3344,
    n3345, n3346, n3347, n3348, n3349, n3350, n3351, n3352, n3353, n3354,
    n3355, n3356, n3357, n3358, n3359, n3360, n3361, n3362, n3363, n3364,
    n3365, n3366, n3367, n3368, n3369, n3370, n3371, n3372, n3373, n3374,
    n3375, n3376, n3377, n3378, n3379, n3380, n3381, n3382, n3383, n3384,
    n3385, n3386, n3387, n3388, n3389, n3390, n3391, n3392, n3393, n3394,
    n3395, n3396, n3397, n3398, n3399, n3400, n3401, n3402, n3403, n3404,
    n3405, n3406, n3407, n3408, n3409, n3410, n3411, n3412, n3413, n3414,
    n3415, n3416, n3417, n3418, n3419, n3420, n3421, n3422, n3423, n3424,
    n3425, n3426, n3427, n3428, n3429, n3430, n3431, n3432, n3433, n3434,
    n3435, n3436, n3437, n3438, n3439, n3440, n3441, n3443, n3444, n3445,
    n3446, n3447, n3448, n3449, n3450, n3451, n3452, n3453, n3454, n3455,
    n3456, n3457, n3458, n3459, n3460, n3461, n3462, n3463, n3464, n3465,
    n3466, n3467, n3468, n3469, n3470, n3471, n3472, n3473, n3474, n3475,
    n3476, n3477, n3478, n3479, n3480, n3481, n3482, n3483, n3484, n3485,
    n3486, n3487, n3488, n3489, n3490, n3491, n3492, n3493, n3494, n3495,
    n3496, n3497, n3498, n3499, n3500, n3501, n3502, n3503, n3504, n3505,
    n3506, n3507, n3508, n3509, n3510, n3511, n3512, n3513, n3514, n3515,
    n3516, n3517, n3518, n3519, n3520, n3521, n3522, n3523, n3524, n3525,
    n3526, n3527, n3528, n3529, n3530, n3531, n3532, n3533, n3534, n3535,
    n3536, n3537, n3538, n3539, n3540, n3541, n3542, n3543, n3544, n3545,
    n3546, n3547, n3548, n3549, n3550, n3551, n3552, n3553, n3554, n3555,
    n3556, n3557, n3558, n3559, n3560, n3561, n3562, n3563, n3564, n3565,
    n3566, n3567, n3568, n3569, n3570, n3571, n3572, n3573, n3574, n3575,
    n3576, n3577, n3578, n3579, n3580, n3581, n3582, n3583, n3584, n3585,
    n3586, n3587, n3588, n3589, n3590, n3591, n3592, n3593, n3594, n3595,
    n3596, n3597, n3598, n3599, n3600, n3601, n3602, n3603, n3604, n3605,
    n3606, n3607, n3608, n3609, n3610, n3611, n3612, n3613, n3614, n3615,
    n3616, n3617, n3618, n3619, n3620, n3621, n3622, n3623, n3624, n3625,
    n3626, n3627, n3628, n3629, n3630, n3631, n3632, n3633, n3634, n3635,
    n3636, n3637, n3638, n3639, n3640, n3641, n3642, n3643, n3644, n3645,
    n3646, n3647, n3648, n3649, n3650, n3651, n3652, n3653, n3654, n3655,
    n3656, n3657, n3658, n3659, n3660, n3661, n3662, n3663, n3664, n3665,
    n3666, n3667, n3668, n3669, n3670, n3671, n3672, n3673, n3674, n3675,
    n3676, n3677, n3678, n3679, n3680, n3681, n3682, n3683, n3684, n3685,
    n3686, n3687, n3688, n3689, n3690, n3691, n3692, n3693, n3694, n3695,
    n3696, n3697, n3698, n3699, n3700, n3701, n3702, n3703, n3704, n3705,
    n3706, n3707, n3708, n3709, n3710, n3711, n3712, n3713, n3714, n3715,
    n3716, n3717, n3718, n3720, n3721, n3722, n3723, n3724, n3725, n3726,
    n3727, n3728, n3729, n3730, n3731, n3732, n3733, n3734, n3735, n3736,
    n3737, n3738, n3739, n3740, n3741, n3742, n3743, n3744, n3745, n3746,
    n3747, n3748, n3749, n3750, n3751, n3752, n3753, n3754, n3755, n3756,
    n3757, n3758, n3759, n3760, n3761, n3762, n3763, n3764, n3765, n3766,
    n3767, n3768, n3769, n3770, n3771, n3772, n3773, n3774, n3775, n3776,
    n3777, n3778, n3779, n3780, n3781, n3782, n3783, n3784, n3785, n3786,
    n3787, n3788, n3789, n3790, n3791, n3792, n3793, n3794, n3795, n3796,
    n3797, n3798, n3799, n3800, n3801, n3802, n3803, n3804, n3805, n3806,
    n3807, n3808, n3809, n3810, n3811, n3812, n3813, n3814, n3815, n3816,
    n3817, n3818, n3819, n3820, n3821, n3822, n3823, n3824, n3825, n3826,
    n3827, n3828, n3829, n3830, n3831, n3832, n3833, n3834, n3835, n3836,
    n3837, n3838, n3839, n3840, n3841, n3842, n3843, n3844, n3845, n3846,
    n3847, n3848, n3849, n3850, n3851, n3852, n3853, n3854, n3855, n3856,
    n3857, n3858, n3859, n3860, n3861, n3862, n3863, n3864, n3865, n3866,
    n3867, n3868, n3869, n3870, n3871, n3872, n3873, n3874, n3875, n3876,
    n3877, n3878, n3879, n3880, n3881, n3882, n3883, n3884, n3885, n3886,
    n3887, n3888, n3889, n3890, n3891, n3892, n3893, n3894, n3895, n3896,
    n3897, n3898, n3899, n3900, n3901, n3902, n3903, n3904, n3905, n3906,
    n3907, n3908, n3909, n3910, n3911, n3912, n3913, n3914, n3915, n3916,
    n3917, n3918, n3919, n3920, n3921, n3922, n3923, n3924, n3925, n3926,
    n3927, n3928, n3929, n3930, n3931, n3932, n3933, n3934, n3935, n3936,
    n3937, n3938, n3939, n3940, n3941, n3942, n3943, n3944, n3945, n3946,
    n3947, n3948, n3949, n3950, n3951, n3952, n3953, n3954, n3955, n3956,
    n3957, n3958, n3959, n3960, n3961, n3962, n3963, n3964, n3965, n3966,
    n3967, n3968, n3969, n3970, n3971, n3972, n3973, n3974, n3975, n3976,
    n3977, n3978, n3979, n3980, n3981, n3982, n3983, n3984, n3985, n3986,
    n3987, n3988, n3989, n3990, n3991, n3992, n3993, n3994, n3995, n3996,
    n3997, n3998, n3999, n4000, n4001, n4002, n4003, n4004, n4005, n4006,
    n4007, n4008, n4009, n4010, n4011, n4012, n4013, n4014, n4015, n4016,
    n4017, n4018, n4019, n4020, n4021, n4022, n4023, n4024, n4025, n4026,
    n4027, n4028, n4029, n4030, n4031, n4032, n4033, n4034, n4035, n4036,
    n4037, n4038, n4039, n4040, n4041, n4042, n4043, n4044, n4045, n4046,
    n4047, n4048, n4049, n4050, n4051, n4052, n4053, n4054, n4055, n4056,
    n4057, n4058, n4059, n4060, n4061, n4062, n4063, n4064, n4065, n4066,
    n4067, n4068, n4069, n4070, n4071, n4072, n4073, n4074, n4075, n4076,
    n4077, n4078, n4079, n4080, n4081, n4082, n4083, n4084, n4085, n4086,
    n4087, n4088, n4089, n4090, n4091, n4092, n4093, n4094, n4095, n4096,
    n4097, n4098, n4099, n4100, n4101, n4102, n4103, n4104, n4105, n4106,
    n4107, n4108, n4109, n4110, n4111, n4112, n4113, n4114, n4115, n4116,
    n4117, n4118, n4119, n4120, n4121, n4122, n4123, n4124, n4125, n4126,
    n4127, n4128, n4129, n4130, n4131, n4132, n4133, n4134, n4135, n4136,
    n4137, n4138, n4139, n4140, n4141, n4142, n4143, n4144, n4145, n4146,
    n4147, n4148, n4149, n4150, n4151, n4152, n4153, n4154, n4155, n4156,
    n4157, n4158, n4159, n4160, n4161, n4162, n4163, n4164, n4165, n4166,
    n4167, n4168, n4169, n4170, n4171, n4172, n4173, n4174, n4175, n4176,
    n4177, n4178, n4179, n4180, n4181, n4182, n4183, n4184, n4185, n4186,
    n4187, n4188, n4189, n4190, n4191, n4192, n4193, n4194, n4195, n4196,
    n4197, n4198, n4199, n4200, n4201, n4202, n4203, n4204, n4205, n4206,
    n4207, n4208, n4209, n4210, n4211, n4212, n4213, n4214, n4215, n4216,
    n4217, n4218, n4219, n4220, n4221, n4222, n4223, n4224, n4225, n4226,
    n4227, n4228, n4229, n4230, n4231, n4232, n4233, n4234, n4235, n4236,
    n4237, n4238, n4239, n4240, n4241, n4242, n4243, n4244, n4245, n4246,
    n4247, n4248, n4249, n4250, n4251, n4252, n4253, n4254, n4255, n4256,
    n4257, n4258, n4259, n4260, n4261, n4262, n4263, n4264, n4265, n4266,
    n4267, n4268, n4269, n4270, n4271, n4272, n4273, n4274, n4275, n4276,
    n4277, n4278, n4279, n4280, n4281, n4282, n4283, n4284, n4285, n4286,
    n4287, n4288, n4289, n4290, n4291, n4292, n4293, n4294, n4295, n4296,
    n4297, n4298, n4299, n4300, n4301, n4302, n4303, n4304, n4305, n4306,
    n4307, n4308, n4309, n4310, n4311, n4312, n4313, n4314, n4315, n4316,
    n4317, n4318, n4319, n4320, n4321, n4322, n4323, n4324, n4325, n4326,
    n4327, n4328, n4329, n4330, n4331, n4332, n4333, n4334, n4335, n4336,
    n4337, n4338, n4339, n4340, n4341, n4342, n4343, n4344, n4345, n4346,
    n4347, n4348, n4349, n4350, n4351, n4352, n4353, n4354, n4355, n4356,
    n4357, n4358, n4359, n4360, n4361, n4362, n4363, n4364, n4365, n4366,
    n4367, n4368, n4369, n4370, n4371, n4372, n4373, n4374, n4375, n4376,
    n4377, n4378, n4379, n4380, n4381, n4382, n4383, n4384, n4385, n4386,
    n4387, n4388, n4389, n4390, n4391, n4392, n4393, n4394, n4395, n4396,
    n4397, n4398, n4399, n4400, n4401, n4402, n4403, n4404, n4405, n4406,
    n4407, n4408, n4409, n4410, n4411, n4412, n4413, n4414, n4415, n4416,
    n4417, n4418, n4419, n4420, n4421, n4422, n4423, n4424, n4425, n4426,
    n4427, n4428, n4429, n4430, n4431, n4432, n4433, n4434, n4435, n4436,
    n4437, n4438, n4439, n4440, n4441, n4442, n4443, n4444, n4445, n4446,
    n4447, n4448, n4449, n4450, n4451, n4452, n4453, n4454, n4455, n4456,
    n4457, n4458, n4459, n4460, n4461, n4462, n4463, n4464, n4465, n4466,
    n4467, n4468, n4469, n4470, n4471, n4472, n4473, n4474, n4475, n4476,
    n4477, n4478, n4479, n4480, n4481, n4482, n4483, n4484, n4485, n4486,
    n4487, n4488, n4489, n4490, n4491, n4492, n4493, n4494, n4495, n4496,
    n4497, n4498, n4499, n4500, n4501, n4502, n4503, n4504, n4505, n4506,
    n4507, n4508, n4509, n4510, n4511, n4512, n4513, n4514, n4515, n4516,
    n4517, n4518, n4519, n4520, n4521, n4522, n4523, n4524, n4525, n4526,
    n4527, n4528, n4529, n4530, n4531, n4532, n4533, n4534, n4535, n4536,
    n4537, n4538, n4539, n4540, n4541, n4542, n4543, n4544, n4545, n4546,
    n4547, n4548, n4549, n4550, n4551, n4552, n4553, n4554, n4555, n4556,
    n4557, n4558, n4559, n4560, n4561, n4562, n4563, n4564, n4565, n4566,
    n4567, n4568, n4569, n4570, n4571, n4572, n4573, n4574, n4575, n4576,
    n4577, n4578, n4579, n4580, n4581, n4582, n4583, n4584, n4585, n4586,
    n4587, n4588, n4589, n4590, n4591, n4592, n4593, n4594, n4595, n4596,
    n4597, n4598, n4599, n4600, n4601, n4602, n4603, n4604, n4605, n4606,
    n4607, n4608, n4609, n4610, n4611, n4612, n4613, n4614, n4615, n4616,
    n4617, n4618, n4619, n4620, n4621, n4622, n4623, n4624, n4625, n4626,
    n4627, n4628, n4629, n4630, n4631, n4632, n4633, n4634, n4635, n4636,
    n4637, n4638, n4639, n4640, n4641, n4642, n4643, n4644, n4645, n4646,
    n4647, n4648, n4649, n4650, n4651, n4652, n4653, n4654, n4655, n4656,
    n4657, n4658, n4659, n4660, n4661, n4662, n4663, n4664, n4665, n4666,
    n4667, n4668, n4669, n4670, n4671, n4672, n4673, n4674, n4675, n4676,
    n4677, n4678, n4679, n4680, n4681, n4682, n4683, n4684, n4685, n4686,
    n4687, n4688, n4689, n4690, n4691, n4692, n4693, n4694, n4695, n4696,
    n4697, n4698, n4699, n4700, n4701, n4702, n4703, n4704, n4705, n4706,
    n4707, n4708, n4709, n4710, n4711, n4712, n4713, n4714, n4715, n4716,
    n4717, n4718, n4719, n4720, n4721, n4722, n4723, n4724, n4725, n4726,
    n4727, n4728, n4729, n4730, n4731, n4732, n4733, n4734, n4735, n4736,
    n4737, n4738, n4739, n4740, n4741, n4742, n4743, n4744, n4745, n4746,
    n4747, n4748, n4749, n4750, n4751, n4752, n4753, n4754, n4755, n4756,
    n4757, n4758, n4759, n4760, n4761, n4762, n4763, n4764, n4765, n4766,
    n4767, n4768, n4769, n4770, n4771, n4772, n4773, n4774, n4775, n4776,
    n4777, n4778, n4779, n4780, n4781, n4782, n4783, n4784, n4785, n4786,
    n4787, n4788, n4789, n4790, n4791, n4792, n4793, n4794, n4795, n4796,
    n4797, n4798, n4799, n4800, n4801, n4802, n4803, n4804, n4805, n4806,
    n4807, n4808, n4809, n4810, n4811, n4812, n4813, n4814, n4815, n4816,
    n4817, n4818, n4819, n4820, n4821, n4822, n4823, n4824, n4825, n4826,
    n4827, n4828, n4829, n4830, n4831, n4832, n4833, n4834, n4835, n4836,
    n4837, n4838, n4839, n4840, n4841, n4842, n4843, n4844, n4845, n4846,
    n4847, n4848, n4849, n4850, n4851, n4852, n4853, n4854, n4855, n4856,
    n4857, n4858, n4859, n4860, n4861, n4862, n4863, n4864, n4865, n4866,
    n4867, n4868, n4869, n4870, n4871, n4872, n4873, n4874, n4875, n4876,
    n4877, n4878, n4879, n4880, n4881, n4882, n4883, n4884, n4885, n4886,
    n4887, n4888, n4889, n4890, n4891, n4892, n4893, n4894, n4895, n4896,
    n4897, n4898, n4899, n4900, n4901, n4902, n4903, n4904, n4905, n4906,
    n4907, n4908, n4909, n4910, n4911, n4912, n4913, n4914, n4915, n4916,
    n4917, n4918, n4919, n4920, n4921, n4922, n4923, n4924, n4925, n4926,
    n4927, n4928, n4929, n4930, n4931, n4932, n4933, n4934, n4935, n4936,
    n4937, n4938, n4939, n4940, n4941, n4942, n4943, n4944, n4945, n4946,
    n4947, n4948, n4949, n4950, n4951, n4952, n4953, n4954, n4955, n4956,
    n4957, n4958, n4959, n4960, n4961, n4962, n4963, n4964, n4965, n4966,
    n4967, n4968, n4969, n4970, n4971, n4972, n4973, n4974, n4975, n4976,
    n4977, n4978, n4979, n4980, n4981, n4982, n4983, n4984, n4985, n4986,
    n4987, n4988, n4989, n4990, n4991, n4992, n4993, n4994, n4995, n4996,
    n4997, n4998, n4999, n5000, n5001, n5002, n5003, n5004, n5005, n5006,
    n5007, n5008, n5009, n5010, n5011, n5012, n5013, n5014, n5015, n5016,
    n5017, n5018, n5019, n5020, n5021, n5022, n5023, n5024, n5025, n5026,
    n5027, n5028, n5029, n5030, n5031, n5032, n5033, n5034, n5035, n5036,
    n5037, n5038, n5039, n5040, n5041, n5042, n5043, n5044, n5045, n5046,
    n5047, n5048, n5049, n5050, n5051, n5052, n5053, n5054, n5055, n5056,
    n5057, n5058, n5059, n5060, n5061, n5062, n5063, n5064, n5065, n5066,
    n5067, n5068, n5069, n5070, n5071, n5072, n5073, n5074, n5075, n5076,
    n5077, n5078, n5079, n5080, n5081, n5082, n5083, n5084, n5085, n5086,
    n5087, n5088, n5089, n5090, n5091, n5092, n5093, n5094, n5095, n5096,
    n5097, n5098, n5099, n5100, n5101, n5102, n5103, n5104, n5105, n5106,
    n5107, n5108, n5109, n5110, n5111, n5112, n5113, n5114, n5115, n5116,
    n5117, n5118, n5119, n5120, n5121, n5122, n5123, n5124, n5125, n5126,
    n5127, n5128, n5129, n5130, n5131, n5132, n5133, n5134, n5135, n5136,
    n5137, n5138, n5139, n5140, n5141, n5142, n5143, n5144, n5145, n5146,
    n5147, n5148, n5149, n5150, n5151, n5152, n5153, n5154, n5155, n5156,
    n5157, n5158, n5159, n5160, n5161, n5162, n5163, n5164, n5165, n5166,
    n5167, n5168, n5169, n5170, n5171, n5172, n5173, n5174, n5175, n5176,
    n5177, n5178, n5179, n5180, n5181, n5182, n5183, n5184, n5185, n5186,
    n5187, n5188, n5189, n5190, n5191, n5192, n5193, n5194, n5195, n5196,
    n5197, n5198, n5199, n5200, n5201, n5202, n5203, n5204, n5205, n5206,
    n5207, n5208, n5209, n5210, n5211, n5212, n5213, n5214, n5215, n5216,
    n5217, n5218, n5219, n5220, n5221, n5222, n5223, n5224, n5225, n5226,
    n5227, n5228, n5229, n5230, n5231, n5232, n5233, n5234, n5235, n5236,
    n5237, n5238, n5239, n5240, n5241, n5242, n5243, n5244, n5245, n5246,
    n5247, n5248, n5249, n5250, n5251, n5252, n5253, n5254, n5255, n5256,
    n5257, n5258, n5259, n5260, n5261, n5262, n5263, n5264, n5265, n5266,
    n5267, n5268, n5269, n5270, n5271, n5272, n5273, n5274, n5275, n5276,
    n5277, n5278, n5279, n5280, n5281, n5282, n5283, n5284, n5285, n5286,
    n5287, n5288, n5289, n5290, n5291, n5292, n5293, n5294, n5295, n5296,
    n5297, n5298, n5299, n5300, n5301, n5302, n5303, n5304, n5305, n5306,
    n5307, n5308, n5309, n5310, n5311, n5312, n5313, n5314, n5315, n5316,
    n5317, n5318, n5319, n5320, n5321, n5322, n5323, n5324, n5325, n5326,
    n5327, n5328, n5329, n5330, n5331, n5332, n5333, n5334, n5335, n5336,
    n5337, n5338, n5339, n5340, n5341, n5342, n5343, n5344, n5345, n5346,
    n5347, n5348, n5349, n5350, n5351, n5352, n5353, n5354, n5355, n5356,
    n5357, n5358, n5359, n5360, n5361, n5362, n5363, n5364, n5365, n5366,
    n5367, n5368, n5369, n5370, n5371, n5372, n5373, n5374, n5375, n5376,
    n5377, n5378, n5379, n5380, n5381, n5382, n5383, n5384, n5385, n5386,
    n5387, n5388, n5389, n5390, n5391, n5392, n5393, n5394, n5395, n5396,
    n5397, n5398, n5399, n5400, n5401, n5402, n5403, n5404, n5405, n5406,
    n5407, n5408, n5409, n5410, n5411, n5412, n5413, n5414, n5415, n5416,
    n5417, n5418, n5419, n5420, n5421, n5422, n5423, n5424, n5425, n5426,
    n5427, n5428, n5429, n5430, n5431, n5432, n5433, n5434, n5435, n5436,
    n5437, n5438, n5439, n5440, n5441, n5442, n5443, n5444, n5445, n5446,
    n5447, n5448, n5449, n5450, n5451, n5452, n5453, n5454, n5455, n5456,
    n5457, n5458, n5459, n5460, n5461, n5462, n5463, n5464, n5465, n5466,
    n5467, n5468, n5469, n5470, n5471, n5472, n5473, n5474, n5475, n5476,
    n5477, n5478, n5479, n5480, n5481, n5482, n5483, n5484, n5485, n5486,
    n5487, n5488, n5489, n5490, n5491, n5492, n5493, n5494, n5495, n5496,
    n5497, n5498, n5499, n5500, n5501, n5502, n5503, n5504, n5505, n5506,
    n5507, n5508, n5509, n5510, n5511, n5512, n5513, n5514, n5515, n5516,
    n5517, n5518, n5519, n5520, n5521, n5522, n5523, n5524, n5525, n5526,
    n5527, n5528, n5529, n5530, n5531, n5532, n5533, n5534, n5535, n5536,
    n5537, n5538, n5539, n5540, n5541, n5542, n5543, n5544, n5545, n5546,
    n5547, n5548, n5549, n5550, n5551, n5552, n5553, n5554, n5555, n5556,
    n5557, n5558, n5559, n5560, n5561, n5562, n5563, n5564, n5565, n5566,
    n5567, n5568, n5569, n5570, n5571, n5572, n5573, n5574, n5575, n5576,
    n5577, n5578, n5579, n5580, n5581, n5582, n5583, n5584, n5585, n5586,
    n5587, n5588, n5589, n5590, n5591, n5592, n5593, n5594, n5595, n5596,
    n5597, n5598, n5599, n5600, n5601, n5602, n5603, n5604, n5605, n5606,
    n5607, n5608, n5609, n5610, n5611, n5612, n5613, n5614, n5615, n5616,
    n5617, n5618, n5619, n5620, n5621, n5622, n5623, n5624, n5625, n5626,
    n5627, n5628, n5629, n5630, n5631, n5632, n5633, n5634, n5635, n5636,
    n5637, n5638, n5639, n5640, n5641, n5642, n5643, n5644, n5645, n5646,
    n5647, n5648, n5649, n5650, n5651, n5652, n5653, n5654, n5655, n5656,
    n5657, n5658, n5659, n5660, n5661, n5662, n5663, n5664, n5665, n5666,
    n5667, n5668, n5669, n5670, n5671, n5672, n5673, n5674, n5675, n5676,
    n5677, n5678, n5679, n5680, n5681, n5682, n5683, n5684, n5685, n5686,
    n5687, n5688, n5689, n5690, n5691, n5692, n5693, n5694, n5695, n5696,
    n5697, n5698, n5699, n5700, n5701, n5702, n5703, n5704, n5705, n5706,
    n5707, n5708, n5709, n5710, n5711, n5712, n5713, n5714, n5715, n5716,
    n5717, n5718, n5719, n5720, n5721, n5722, n5723, n5724, n5725, n5726,
    n5727, n5728, n5729, n5730, n5731, n5732, n5733, n5734, n5735, n5736,
    n5737, n5738, n5739, n5740, n5741, n5742, n5743, n5744, n5745, n5746,
    n5747, n5748, n5749, n5750, n5751, n5752, n5753, n5754, n5755, n5756,
    n5757, n5758, n5759, n5760, n5761, n5762, n5763, n5764, n5765, n5766,
    n5767, n5768, n5769, n5770, n5771, n5772, n5773, n5774, n5775, n5776,
    n5777, n5778, n5779, n5780, n5781, n5782, n5783, n5784, n5785, n5786,
    n5787, n5788, n5789, n5790, n5791, n5792, n5793, n5794, n5795, n5796,
    n5797, n5798, n5799, n5800, n5801, n5802, n5803, n5804, n5805, n5806,
    n5807, n5808, n5809, n5810, n5811, n5812, n5813, n5814, n5815, n5816,
    n5817, n5818, n5819, n5820, n5821, n5822, n5823, n5824, n5825, n5826,
    n5827, n5828, n5829, n5830, n5831, n5832, n5833, n5834, n5835, n5836,
    n5837, n5838, n5839, n5840, n5841, n5842, n5843, n5844, n5845, n5846,
    n5847, n5848, n5849, n5850, n5851, n5852, n5853, n5854, n5855, n5856,
    n5857, n5858, n5859, n5860, n5861, n5862, n5863, n5864, n5865, n5866,
    n5867, n5868, n5869, n5870, n5871, n5872, n5873, n5874, n5875, n5876,
    n5877, n5878, n5879, n5880, n5881, n5882, n5883, n5884, n5885, n5886,
    n5887, n5888, n5889, n5890, n5891, n5892, n5893, n5894, n5895, n5896,
    n5897, n5898, n5899, n5900, n5901, n5902, n5903, n5904, n5905, n5906,
    n5907, n5908, n5909, n5910, n5911, n5912, n5913, n5914, n5915, n5916,
    n5917, n5918, n5919, n5920, n5921, n5922, n5923, n5924, n5925, n5926,
    n5927, n5928, n5929, n5930, n5931, n5932, n5933, n5934, n5935, n5936,
    n5937, n5938, n5939, n5940, n5941, n5942, n5943, n5944, n5945, n5946,
    n5947, n5948, n5949, n5950, n5951, n5952, n5953, n5954, n5955, n5956,
    n5957, n5958, n5959, n5960, n5961, n5962, n5963, n5964, n5965, n5966,
    n5967, n5968, n5969, n5970, n5971, n5972, n5973, n5974, n5975, n5976,
    n5977, n5978, n5979, n5980, n5981, n5982, n5983, n5984, n5985, n5986,
    n5987, n5988, n5989, n5990, n5991, n5992, n5993, n5994, n5995, n5996,
    n5997, n5998, n5999, n6000, n6001, n6002, n6003, n6004, n6005, n6006,
    n6007, n6008, n6009, n6010, n6011, n6012, n6013, n6014, n6015, n6016,
    n6017, n6018, n6019, n6020, n6021, n6022, n6023, n6024, n6025, n6026,
    n6027, n6028, n6029, n6030, n6031, n6032, n6033, n6034, n6035, n6036,
    n6037, n6038, n6039, n6040, n6041, n6042, n6043, n6044, n6045, n6046,
    n6047, n6048, n6049, n6050, n6051, n6052, n6053, n6054, n6055, n6056,
    n6057, n6058, n6059, n6060, n6061, n6062, n6063, n6064, n6065, n6066,
    n6067, n6068, n6069, n6070, n6071, n6072, n6073, n6074, n6075, n6076,
    n6077, n6078, n6079, n6080, n6081, n6082, n6083, n6084, n6085, n6086,
    n6087, n6088, n6089, n6090, n6091, n6092, n6093, n6094, n6095, n6096,
    n6097, n6098, n6099, n6100, n6101, n6102, n6103, n6104, n6105, n6106,
    n6107, n6108, n6109, n6110, n6111, n6112, n6113, n6114, n6115, n6116,
    n6117, n6118, n6119, n6120, n6121, n6122, n6123, n6124, n6125, n6126,
    n6127, n6128, n6129, n6130, n6131, n6132, n6133, n6134, n6135, n6136,
    n6137, n6138, n6139, n6140, n6141, n6142, n6143, n6144, n6145, n6146,
    n6147, n6148, n6149, n6150, n6151, n6152, n6153, n6154, n6155, n6156,
    n6157, n6158, n6159, n6160, n6161, n6162, n6163, n6164, n6165, n6166,
    n6167, n6168, n6169, n6170, n6171, n6172, n6173, n6174, n6175, n6176,
    n6177, n6178, n6179, n6180, n6181, n6182, n6183, n6184, n6185, n6186,
    n6187, n6188, n6189, n6190, n6191, n6192, n6193, n6194, n6195, n6196,
    n6197, n6198, n6199, n6200, n6201, n6202, n6203, n6204, n6205, n6206,
    n6207, n6208, n6209, n6210, n6211, n6212, n6213, n6214, n6215, n6216,
    n6217, n6218, n6219, n6220, n6221, n6222, n6223, n6224, n6225, n6226,
    n6227, n6228, n6229, n6230, n6231, n6232, n6233, n6234, n6235, n6236,
    n6237, n6238, n6239, n6240, n6241, n6242, n6243, n6244, n6245, n6246,
    n6247, n6248, n6249, n6250, n6251, n6252, n6253, n6254, n6255, n6256,
    n6257, n6258, n6259, n6260, n6261, n6262, n6263, n6264, n6265, n6266,
    n6267, n6268, n6269, n6270, n6271, n6272, n6273, n6274, n6275, n6276,
    n6277, n6278, n6279, n6280, n6281, n6282, n6283, n6284, n6285, n6286,
    n6287, n6288, n6289, n6290, n6291, n6292, n6293, n6294, n6295, n6296,
    n6297, n6298, n6299, n6300, n6301, n6302, n6303, n6304, n6305, n6306,
    n6307, n6308, n6309, n6310, n6311, n6312, n6313, n6314, n6315, n6316,
    n6317, n6318, n6319, n6320, n6321, n6322, n6323, n6324, n6325, n6326,
    n6327, n6328, n6329, n6330, n6331, n6332, n6333, n6334, n6335, n6336,
    n6337, n6338, n6339, n6340, n6341, n6342, n6343, n6344, n6345, n6346,
    n6347, n6348, n6349, n6350, n6351, n6352, n6353, n6354, n6355, n6356,
    n6357, n6358, n6359, n6360, n6361, n6362, n6363, n6364, n6365, n6366,
    n6367, n6368, n6369, n6370, n6371, n6372, n6373, n6374, n6375, n6376,
    n6377, n6378, n6379, n6380, n6381, n6382, n6383, n6384, n6385, n6386,
    n6387, n6388, n6389, n6390, n6391, n6392, n6393, n6394, n6395, n6396,
    n6397, n6398, n6399, n6400, n6401, n6402, n6403, n6404, n6405, n6406,
    n6407, n6408, n6409, n6410, n6411, n6412, n6413, n6414, n6415, n6416,
    n6417, n6418, n6419, n6420, n6421, n6422, n6423, n6424, n6425, n6426,
    n6427, n6428, n6429, n6430, n6431, n6432, n6433, n6434, n6435, n6436,
    n6437, n6438, n6439, n6440, n6441, n6442, n6443, n6444, n6445, n6446,
    n6447, n6448, n6449, n6450, n6451, n6452, n6453, n6454, n6455, n6456,
    n6457, n6458, n6459, n6460, n6461, n6462, n6463, n6464, n6465, n6466,
    n6467, n6468, n6469, n6470, n6471, n6472, n6473, n6474, n6475, n6476,
    n6477, n6478, n6479, n6480, n6481, n6482, n6483, n6484, n6485, n6486,
    n6487, n6488, n6489, n6490, n6491, n6492, n6493, n6494, n6495, n6496,
    n6497, n6498, n6499, n6500, n6501, n6502, n6503, n6504, n6505, n6506,
    n6507, n6508, n6509, n6510, n6511, n6512, n6513, n6514, n6515, n6516,
    n6517, n6518, n6519, n6520, n6521, n6522, n6523, n6524, n6525, n6526,
    n6527, n6528, n6529, n6530, n6531, n6532, n6533, n6534, n6535, n6536,
    n6537, n6538, n6539, n6540, n6541, n6542, n6543, n6544, n6545, n6546,
    n6547, n6548, n6549, n6550, n6551, n6552, n6553, n6554, n6555, n6556,
    n6557, n6558, n6559, n6560, n6561, n6562, n6563, n6564, n6565, n6566,
    n6567, n6568, n6569, n6570, n6571, n6572, n6573, n6574, n6575, n6576,
    n6577, n6578, n6579, n6580, n6581, n6582, n6583, n6584, n6585, n6586,
    n6587, n6588, n6589, n6590, n6591, n6592, n6593, n6594, n6595, n6596,
    n6597, n6598, n6599, n6600, n6601, n6602, n6603, n6604, n6605, n6606,
    n6607, n6608, n6609, n6610, n6611, n6612, n6613, n6614, n6615, n6616,
    n6617, n6618, n6619, n6620, n6621, n6622, n6623, n6624, n6625, n6626,
    n6627, n6628, n6629, n6630, n6631, n6632, n6633, n6634, n6635, n6636,
    n6637, n6638, n6639, n6640, n6641, n6642, n6643, n6644, n6645, n6646,
    n6647, n6648, n6649, n6650, n6651, n6652, n6653, n6654, n6655, n6656,
    n6657, n6658, n6659, n6660, n6661, n6662, n6663, n6664, n6665, n6666,
    n6667, n6668, n6669, n6670, n6671, n6672, n6673, n6674, n6675, n6676,
    n6677, n6678, n6679, n6680, n6681, n6682, n6683, n6684, n6685, n6686,
    n6687, n6688, n6689, n6690, n6691, n6692, n6693, n6694, n6695, n6696,
    n6697, n6698, n6699, n6700, n6701, n6702, n6703, n6704, n6705, n6706,
    n6707, n6708, n6709, n6710, n6711, n6712, n6713, n6714, n6715, n6716,
    n6717, n6718, n6719, n6720, n6721, n6722, n6723, n6724, n6725, n6726,
    n6727, n6728, n6729, n6730, n6731, n6732, n6733, n6734, n6735, n6736,
    n6737, n6738, n6739, n6740, n6741, n6742, n6743, n6744, n6745, n6746,
    n6747, n6748, n6749, n6750, n6751, n6752, n6753, n6754, n6755, n6756,
    n6757, n6758, n6759, n6760, n6761, n6762, n6763, n6764, n6765, n6766,
    n6767, n6768, n6769, n6770, n6771, n6772, n6773, n6774, n6775, n6776,
    n6777, n6778, n6779, n6780, n6781, n6782, n6783, n6784, n6785, n6786,
    n6787, n6788, n6789, n6790, n6791, n6792, n6793, n6794, n6795, n6796,
    n6797, n6798, n6799, n6800, n6801, n6802, n6803, n6804, n6805, n6806,
    n6807, n6808, n6809, n6810, n6811, n6812, n6813, n6814, n6815, n6816,
    n6817, n6818, n6819, n6820, n6821, n6822, n6823, n6824, n6825, n6826,
    n6827, n6828, n6829, n6830, n6831, n6832, n6833, n6834, n6835, n6836,
    n6837, n6838, n6839, n6840, n6841, n6842, n6843, n6844, n6845, n6846,
    n6847, n6848, n6849, n6850, n6851, n6852, n6853, n6854, n6855, n6856,
    n6857, n6858, n6859, n6860, n6861, n6862, n6863, n6864, n6865, n6866,
    n6867, n6868, n6869, n6870, n6871, n6872, n6873, n6874, n6875, n6876,
    n6877, n6878, n6879, n6880, n6881, n6882, n6883, n6884, n6885, n6886,
    n6887, n6888, n6889, n6890, n6891, n6892, n6893, n6894, n6895, n6896,
    n6897, n6898, n6899, n6900, n6901, n6902, n6903, n6904, n6905, n6906,
    n6907, n6908, n6909, n6910, n6911, n6912, n6913, n6914, n6915, n6916,
    n6917, n6918, n6919, n6920, n6921, n6922, n6923, n6924, n6925, n6926,
    n6927, n6928, n6929, n6930, n6931, n6932, n6933, n6934, n6935, n6936,
    n6937, n6938, n6939, n6940, n6941, n6942, n6943, n6944, n6945, n6946,
    n6947, n6948, n6949, n6950, n6951, n6952, n6953, n6954, n6955, n6956,
    n6957, n6958, n6959, n6960, n6961, n6962, n6963, n6964, n6965, n6966,
    n6967, n6968, n6969, n6970, n6971, n6972, n6973, n6974, n6975, n6976,
    n6977, n6978, n6979, n6980, n6981, n6982, n6983, n6984, n6985, n6986,
    n6987, n6988, n6989, n6990, n6991, n6992, n6993, n6994, n6995, n6997,
    n6998, n6999, n7000, n7001, n7002, n7003, n7004, n7005, n7006, n7007,
    n7008, n7010, n7011, n7012, n7013, n7014, n7015, n7016, n7017, n7018,
    n7019, n7020, n7021, n7022, n7023, n7024, n7025, n7026, n7027, n7028,
    n7030, n7031, n7032, n7033, n7034, n7035, n7036, n7037, n7038, n7039,
    n7040, n7041, n7042, n7043, n7044, n7045, n7046, n7048, n7049, n7050,
    n7051, n7052, n7053, n7054, n7055, n7056, n7057, n7058, n7059, n7060,
    n7061, n7063, n7064, n7065, n7066, n7067, n7068, n7069, n7070, n7071,
    n7072, n7073, n7074, n7075, n7076, n7078, n7079, n7080, n7081, n7082,
    n7083, n7084, n7085, n7086, n7087, n7088, n7089, n7090, n7091, n7092,
    n7094, n7095, n7096, n7097, n7098, n7099, n7100, n7101, n7102, n7103,
    n7104, n7105, n7106, n7107, n7108, n7109, n7110, n7111, n7112, n7113,
    n7115, n7116, n7117, n7118, n7119, n7120, n7121, n7122, n7123, n7124,
    n7125, n7126, n7127, n7128, n7130, n7131, n7132, n7133, n7134, n7135,
    n7136, n7137, n7138, n7139, n7140, n7141, n7142, n7144, n7145, n7146,
    n7147, n7148, n7149, n7150, n7151, n7152, n7153, n7154, n7155, n7156,
    n7157, n7158, n7159, n7161, n7162, n7163, n7164, n7165, n7166, n7167,
    n7168, n7169, n7170, n7171, n7172, n7174, n7175, n7176, n7177, n7178,
    n7179, n7180, n7181, n7182, n7183, n7184, n7185, n7186, n7187, n7188,
    n7189, n7190, n7192, n7193, n7194, n7195, n7197, n7198, n7199, n7200,
    n7201, n7202, n7203, n7204, n7205, n7206, n7207, n7208, n7209, n7210,
    n7211, n7212, n7213, n7214, n7215, n7217, n7219, n7220, n7221, n7222,
    n7223, n7224, n7225, n7226, n7227, n7228, n7230, n7231, n7232, n7234,
    n7235, n7236, n7237, n7238;
  assign n65 = ~pi29 & ~pi31;
  assign n66 = ~pi27 & ~pi29;
  assign n67 = ~pi31 & n66;
  assign n68 = ~pi25 & ~pi27;
  assign n69 = n65 & n68;
  assign n70 = pi01 & ~pi14;
  assign n71 = ~pi13 & ~pi15;
  assign n72 = ~pi17 & ~pi19;
  assign n73 = ~pi21 & ~pi23;
  assign n74 = n72 & n73;
  assign n75 = n71 & n74;
  assign n76 = n69 & n75;
  assign n77 = pi01 & ~pi03;
  assign n78 = ~pi09 & ~pi11;
  assign n79 = ~pi05 & ~pi07;
  assign n80 = n78 & n79;
  assign n81 = n77 & n80;
  assign n82 = n68 & n73;
  assign n83 = n71 & n72;
  assign n84 = n82 & n83;
  assign n85 = pi01 & ~pi28;
  assign n86 = ~pi03 & ~n85;
  assign n87 = pi30 & n65;
  assign n88 = ~n86 & n87;
  assign n89 = n84 & n88;
  assign n90 = n81 & n89;
  assign n91 = pi01 & ~pi05;
  assign n92 = ~pi07 & ~pi09;
  assign n93 = n91 & n92;
  assign n94 = pi03 & ~pi30;
  assign n95 = ~n85 & ~n94;
  assign n96 = n93 & n95;
  assign n97 = ~pi19 & ~pi21;
  assign n98 = ~pi23 & ~pi25;
  assign n99 = n97 & n98;
  assign n100 = ~pi11 & ~pi13;
  assign n101 = ~pi15 & ~pi17;
  assign n102 = n100 & n101;
  assign n103 = n99 & n102;
  assign n104 = pi01 & ~pi26;
  assign n105 = ~pi03 & ~n104;
  assign n106 = pi26 & ~pi27;
  assign n107 = n65 & n106;
  assign n108 = ~n105 & n107;
  assign n109 = n103 & n108;
  assign n110 = n96 & n109;
  assign n111 = ~n90 & n110;
  assign n112 = ~pi01 & pi26;
  assign n113 = pi01 & pi03;
  assign n114 = ~pi26 & n113;
  assign n115 = pi28 & ~n114;
  assign n116 = ~n105 & ~n115;
  assign n117 = n71 & n78;
  assign n118 = n79 & n117;
  assign n119 = n69 & n74;
  assign n120 = n118 & n119;
  assign n121 = ~n116 & n120;
  assign n122 = pi26 & ~n121;
  assign n123 = ~n112 & ~n122;
  assign n124 = ~n111 & n123;
  assign n125 = ~pi05 & pi30;
  assign n126 = n77 & n125;
  assign n127 = ~n86 & n126;
  assign n128 = ~n85 & n91;
  assign n129 = ~n94 & n128;
  assign n130 = ~n127 & n129;
  assign n131 = n115 & ~n130;
  assign n132 = pi05 & ~n105;
  assign n133 = ~n131 & n132;
  assign n134 = n79 & ~n85;
  assign n135 = ~n94 & n134;
  assign n136 = n74 & n117;
  assign n137 = n69 & ~n86;
  assign n138 = n136 & n137;
  assign n139 = n135 & n138;
  assign n140 = ~n90 & n139;
  assign n141 = n84 & n87;
  assign n142 = n81 & n141;
  assign n143 = n92 & ~n112;
  assign n144 = n102 & n143;
  assign n145 = pi30 & ~pi31;
  assign n146 = n66 & n145;
  assign n147 = n99 & n146;
  assign n148 = n144 & n147;
  assign n149 = ~n142 & n148;
  assign n150 = ~n140 & n149;
  assign n151 = ~n133 & n150;
  assign n152 = ~n124 & ~n151;
  assign n153 = n78 & n104;
  assign n154 = n83 & n153;
  assign n155 = ~pi07 & ~pi29;
  assign n156 = n145 & n155;
  assign n157 = n82 & n156;
  assign n158 = n154 & n157;
  assign n159 = ~n142 & n158;
  assign n160 = ~n140 & n159;
  assign n161 = ~n133 & n160;
  assign n162 = n67 & ~n105;
  assign n163 = n103 & n162;
  assign n164 = n96 & n163;
  assign n165 = ~n90 & n164;
  assign n166 = n93 & n102;
  assign n167 = ~pi26 & ~pi27;
  assign n168 = n65 & n167;
  assign n169 = n99 & n168;
  assign n170 = n166 & n169;
  assign n171 = ~n116 & n170;
  assign n172 = ~n165 & n171;
  assign n173 = ~n161 & ~n172;
  assign n174 = ~n152 & n173;
  assign n175 = ~n116 & n125;
  assign n176 = ~n142 & n175;
  assign n177 = ~n140 & n176;
  assign n178 = ~n165 & n177;
  assign n179 = n92 & n102;
  assign n180 = n67 & n99;
  assign n181 = n179 & n180;
  assign n182 = ~n133 & n181;
  assign n183 = pi30 & ~n142;
  assign n184 = ~n140 & n183;
  assign n185 = ~n182 & n184;
  assign n186 = pi07 & ~n185;
  assign n187 = ~n178 & n186;
  assign n188 = pi01 & ~pi24;
  assign n189 = ~pi03 & ~n188;
  assign n190 = ~n172 & ~n189;
  assign n191 = ~n161 & n190;
  assign n192 = ~n152 & n191;
  assign n193 = pi03 & ~pi07;
  assign n194 = n78 & n193;
  assign n195 = ~n104 & n194;
  assign n196 = n141 & n195;
  assign n197 = ~n142 & n196;
  assign n198 = ~n140 & n197;
  assign n199 = ~n133 & n198;
  assign n200 = ~pi05 & ~pi09;
  assign n201 = n193 & n200;
  assign n202 = ~n104 & n201;
  assign n203 = n67 & n103;
  assign n204 = n202 & n203;
  assign n205 = ~n116 & n204;
  assign n206 = ~n165 & n205;
  assign n207 = n96 & ~n127;
  assign n208 = n203 & n207;
  assign n209 = pi28 & ~n208;
  assign n210 = pi05 & ~n209;
  assign n211 = ~n206 & n210;
  assign n212 = ~n199 & n211;
  assign n213 = pi05 & ~pi07;
  assign n214 = n78 & n213;
  assign n215 = n83 & n214;
  assign n216 = pi28 & ~pi29;
  assign n217 = n145 & n216;
  assign n218 = n82 & n217;
  assign n219 = ~n105 & n218;
  assign n220 = n215 & n219;
  assign n221 = ~n142 & n220;
  assign n222 = ~n208 & n221;
  assign n223 = ~n133 & ~n140;
  assign n224 = n222 & n223;
  assign n225 = ~pi24 & n113;
  assign n226 = ~n224 & ~n225;
  assign n227 = ~n212 & n226;
  assign n228 = ~n192 & n227;
  assign n229 = ~n187 & n228;
  assign n230 = ~n178 & ~n185;
  assign n231 = n181 & ~n230;
  assign n232 = ~n206 & ~n209;
  assign n233 = ~n199 & n232;
  assign n234 = n97 & n101;
  assign n235 = n92 & n100;
  assign n236 = n234 & n235;
  assign n237 = pi28 & pi30;
  assign n238 = n98 & n237;
  assign n239 = n67 & n238;
  assign n240 = ~n105 & n239;
  assign n241 = n236 & n240;
  assign n242 = ~n142 & n241;
  assign n243 = ~n208 & n242;
  assign n244 = n223 & n243;
  assign n245 = n80 & n83;
  assign n246 = ~pi31 & n216;
  assign n247 = n82 & n246;
  assign n248 = ~n105 & ~n114;
  assign n249 = n247 & n248;
  assign n250 = n245 & n249;
  assign n251 = ~n208 & n250;
  assign n252 = ~n165 & n251;
  assign n253 = ~pi05 & ~n252;
  assign n254 = ~n244 & n253;
  assign n255 = ~n233 & n254;
  assign n256 = ~n187 & n255;
  assign n257 = ~n231 & ~n256;
  assign n258 = ~n229 & n257;
  assign n259 = n69 & n136;
  assign n260 = ~n231 & ~n259;
  assign n261 = ~pi24 & n77;
  assign n262 = pi03 & ~n188;
  assign n263 = ~n261 & ~n262;
  assign n264 = ~n260 & ~n263;
  assign n265 = ~n258 & n264;
  assign n266 = ~n174 & ~n265;
  assign n267 = ~n189 & ~n225;
  assign n268 = ~n172 & n267;
  assign n269 = ~n161 & n268;
  assign n270 = ~n152 & n269;
  assign n271 = ~n260 & n270;
  assign n272 = ~n258 & n271;
  assign n273 = pi05 & ~n272;
  assign n274 = ~n266 & n273;
  assign n275 = ~pi22 & n113;
  assign n276 = n188 & ~n260;
  assign n277 = pi01 & ~pi22;
  assign n278 = ~pi03 & ~n277;
  assign n279 = ~pi01 & pi24;
  assign n280 = ~n278 & ~n279;
  assign n281 = ~n276 & n280;
  assign n282 = n78 & n188;
  assign n283 = n83 & n282;
  assign n284 = ~pi31 & n68;
  assign n285 = n73 & n155;
  assign n286 = n284 & n285;
  assign n287 = n283 & n286;
  assign n288 = ~n230 & n287;
  assign n289 = n280 & ~n288;
  assign n290 = ~n256 & n289;
  assign n291 = ~n229 & n290;
  assign n292 = ~n281 & ~n291;
  assign n293 = pi24 & ~n259;
  assign n294 = ~n231 & n293;
  assign n295 = pi24 & ~n231;
  assign n296 = ~n256 & n295;
  assign n297 = ~n229 & n296;
  assign n298 = ~n294 & ~n297;
  assign n299 = ~n292 & n298;
  assign n300 = ~n275 & ~n299;
  assign n301 = ~n274 & n300;
  assign n302 = ~n229 & ~n256;
  assign n303 = ~pi05 & ~n225;
  assign n304 = ~n252 & n303;
  assign n305 = ~n244 & n304;
  assign n306 = ~n233 & n305;
  assign n307 = ~n192 & n306;
  assign n308 = n259 & ~n307;
  assign n309 = ~n302 & n308;
  assign n310 = ~n244 & ~n252;
  assign n311 = ~n233 & n310;
  assign n312 = ~n231 & n311;
  assign n313 = ~n307 & ~n312;
  assign n314 = ~pi07 & ~n313;
  assign n315 = ~n309 & n314;
  assign n316 = ~n189 & n303;
  assign n317 = ~n172 & n316;
  assign n318 = ~n161 & n317;
  assign n319 = ~n152 & n318;
  assign n320 = ~n260 & n319;
  assign n321 = ~n258 & n320;
  assign n322 = ~n228 & ~n255;
  assign n323 = n231 & ~n322;
  assign n324 = ~n181 & n259;
  assign n325 = ~n230 & n324;
  assign n326 = ~n256 & n325;
  assign n327 = ~n229 & n326;
  assign n328 = ~n323 & ~n327;
  assign n329 = ~n321 & n328;
  assign n330 = ~n315 & n329;
  assign n331 = ~n192 & ~n225;
  assign n332 = pi05 & ~n224;
  assign n333 = ~n212 & n332;
  assign n334 = ~n331 & ~n333;
  assign n335 = ~pi07 & ~n228;
  assign n336 = ~n260 & n335;
  assign n337 = ~n334 & n336;
  assign n338 = ~n258 & n337;
  assign n339 = ~pi05 & ~n174;
  assign n340 = ~n265 & n339;
  assign n341 = ~n338 & ~n340;
  assign n342 = n330 & n341;
  assign n343 = ~n301 & n342;
  assign n344 = n203 & ~n259;
  assign n345 = ~n230 & n344;
  assign n346 = ~n231 & n345;
  assign n347 = ~n323 & ~n346;
  assign n348 = n203 & ~n230;
  assign n349 = ~n231 & n348;
  assign n350 = ~n256 & n349;
  assign n351 = ~n229 & n350;
  assign n352 = pi09 & ~n255;
  assign n353 = ~n228 & n352;
  assign n354 = ~pi07 & ~n230;
  assign n355 = pi09 & ~n354;
  assign n356 = n203 & ~n355;
  assign n357 = ~n353 & n356;
  assign n358 = ~n327 & ~n357;
  assign n359 = ~n351 & n358;
  assign n360 = n347 & n359;
  assign n361 = ~n309 & ~n313;
  assign n362 = ~n228 & ~n260;
  assign n363 = ~n334 & n362;
  assign n364 = ~n258 & n363;
  assign n365 = pi07 & ~n323;
  assign n366 = ~n327 & n365;
  assign n367 = ~n364 & n366;
  assign n368 = ~n361 & n367;
  assign n369 = ~n360 & ~n368;
  assign po22 = ~n343 & n369;
  assign n371 = ~n322 & n354;
  assign po24 = ~n258 & ~n260;
  assign n373 = ~n230 & ~po24;
  assign n374 = ~n371 & ~n373;
  assign n375 = ~po22 & ~n374;
  assign n376 = ~n315 & ~n321;
  assign n377 = n341 & n376;
  assign n378 = ~n301 & n377;
  assign n379 = pi07 & ~n364;
  assign n380 = ~n361 & n379;
  assign n381 = ~pi09 & ~n374;
  assign n382 = ~n380 & n381;
  assign n383 = ~n378 & n382;
  assign n384 = ~n375 & ~n383;
  assign n385 = ~n321 & ~n340;
  assign n386 = ~n301 & n385;
  assign n387 = ~n315 & ~n338;
  assign n388 = ~n380 & n387;
  assign n389 = ~n386 & ~n388;
  assign n390 = n377 & ~n380;
  assign n391 = ~n301 & n390;
  assign n392 = ~n389 & ~n391;
  assign n393 = po22 & ~n392;
  assign n394 = ~n361 & ~n364;
  assign n395 = ~po22 & ~n394;
  assign n396 = pi09 & ~n395;
  assign n397 = ~n393 & n396;
  assign n398 = ~pi11 & ~n384;
  assign n399 = pi11 & ~n383;
  assign n400 = ~n375 & n399;
  assign n401 = n76 & ~n400;
  assign n402 = ~n398 & n401;
  assign n403 = ~n397 & n402;
  assign n404 = n259 & ~n374;
  assign n405 = ~n380 & n404;
  assign n406 = ~n378 & n405;
  assign n407 = n203 & ~n374;
  assign n408 = ~po22 & n407;
  assign n409 = ~n406 & ~n408;
  assign n410 = ~n403 & n409;
  assign n411 = ~n393 & ~n395;
  assign n412 = ~pi09 & ~n411;
  assign n413 = ~n274 & n385;
  assign n414 = ~n300 & ~n413;
  assign n415 = ~n266 & ~n272;
  assign n416 = ~pi05 & ~n415;
  assign n417 = ~n414 & n416;
  assign n418 = ~n346 & ~n357;
  assign n419 = ~n351 & n418;
  assign n420 = ~n380 & ~n419;
  assign n421 = ~n378 & n420;
  assign n422 = n328 & ~n415;
  assign n423 = ~n421 & n422;
  assign n424 = ~n417 & ~n423;
  assign n425 = ~n301 & ~n414;
  assign n426 = po22 & n425;
  assign n427 = n424 & ~n426;
  assign n428 = ~pi07 & ~n427;
  assign n429 = n409 & ~n428;
  assign n430 = ~n412 & n429;
  assign n431 = ~pi07 & ~n425;
  assign n432 = ~pi07 & ~n323;
  assign n433 = ~n327 & n432;
  assign n434 = ~n421 & n433;
  assign n435 = ~n431 & ~n434;
  assign n436 = n424 & ~n435;
  assign n437 = pi07 & ~n360;
  assign n438 = ~n301 & n437;
  assign n439 = ~n368 & n438;
  assign n440 = ~n343 & ~n414;
  assign n441 = n439 & n440;
  assign n442 = pi07 & ~n174;
  assign n443 = ~n265 & n442;
  assign n444 = pi07 & ~n189;
  assign n445 = ~n225 & n444;
  assign n446 = ~n172 & n445;
  assign n447 = ~n161 & n446;
  assign n448 = ~n152 & n447;
  assign n449 = ~n260 & n448;
  assign n450 = ~n258 & n449;
  assign n451 = ~n443 & ~n450;
  assign n452 = ~pi05 & ~n451;
  assign n453 = ~n414 & n452;
  assign n454 = n328 & ~n451;
  assign n455 = ~n421 & n454;
  assign n456 = ~n453 & ~n455;
  assign n457 = ~n441 & n456;
  assign n458 = ~n436 & n457;
  assign n459 = ~pi22 & n77;
  assign n460 = pi03 & ~n277;
  assign n461 = ~n459 & ~n460;
  assign n462 = ~n360 & ~n461;
  assign n463 = ~n368 & n462;
  assign n464 = ~n343 & n463;
  assign n465 = ~n256 & ~n288;
  assign n466 = ~n229 & n465;
  assign n467 = n276 & ~n466;
  assign n468 = ~n279 & ~n294;
  assign n469 = ~n297 & n468;
  assign n470 = ~n467 & n469;
  assign n471 = ~n464 & n470;
  assign n472 = ~n461 & ~n470;
  assign n473 = ~n360 & n472;
  assign n474 = ~n368 & n473;
  assign n475 = ~n343 & n474;
  assign n476 = ~pi05 & ~n475;
  assign n477 = ~n471 & n476;
  assign n478 = ~n458 & n477;
  assign n479 = ~pi05 & ~n279;
  assign n480 = ~n294 & n479;
  assign n481 = ~n297 & n480;
  assign n482 = n328 & n481;
  assign n483 = ~n467 & n482;
  assign n484 = ~n275 & ~n278;
  assign n485 = n479 & ~n484;
  assign n486 = ~n294 & n485;
  assign n487 = ~n297 & n486;
  assign n488 = ~n467 & n487;
  assign n489 = ~n483 & ~n488;
  assign n490 = ~n419 & ~n488;
  assign n491 = ~n380 & n490;
  assign n492 = ~n378 & n491;
  assign n493 = ~n489 & ~n492;
  assign n494 = pi05 & ~n459;
  assign n495 = ~n460 & n494;
  assign n496 = ~n470 & n495;
  assign n497 = pi05 & ~n323;
  assign n498 = ~n327 & n497;
  assign n499 = ~n470 & n498;
  assign n500 = ~n496 & ~n499;
  assign n501 = n420 & ~n496;
  assign n502 = ~n378 & n501;
  assign n503 = ~n500 & ~n502;
  assign n504 = ~pi05 & ~n461;
  assign n505 = ~n470 & n504;
  assign n506 = ~n360 & n505;
  assign n507 = ~n368 & n506;
  assign n508 = ~n343 & n507;
  assign n509 = pi05 & ~n279;
  assign n510 = ~n275 & n509;
  assign n511 = ~n278 & n510;
  assign n512 = ~n294 & n511;
  assign n513 = ~n297 & n512;
  assign n514 = ~n467 & n513;
  assign n515 = ~n360 & n514;
  assign n516 = ~n368 & n515;
  assign n517 = ~n343 & n516;
  assign n518 = ~n508 & ~n517;
  assign n519 = ~n503 & n518;
  assign n520 = ~n493 & n519;
  assign n521 = pi01 & ~n360;
  assign n522 = ~n368 & n521;
  assign n523 = ~n343 & n522;
  assign n524 = ~pi20 & n113;
  assign n525 = pi22 & ~n524;
  assign n526 = ~n523 & n525;
  assign n527 = pi01 & ~pi20;
  assign n528 = n277 & ~n527;
  assign n529 = pi03 & ~n528;
  assign n530 = pi03 & ~n323;
  assign n531 = ~n327 & n530;
  assign n532 = ~n529 & ~n531;
  assign n533 = ~n419 & ~n529;
  assign n534 = ~n380 & n533;
  assign n535 = ~n378 & n534;
  assign n536 = ~n532 & ~n535;
  assign n537 = ~n526 & n536;
  assign n538 = pi22 & ~n523;
  assign n539 = n277 & ~n360;
  assign n540 = ~n368 & n539;
  assign n541 = ~n343 & n540;
  assign n542 = n527 & ~n541;
  assign n543 = ~n538 & n542;
  assign n544 = ~n537 & ~n543;
  assign n545 = ~n520 & n544;
  assign n546 = ~n458 & n545;
  assign n547 = ~n478 & ~n546;
  assign n548 = n430 & n547;
  assign po20 = ~n410 & ~n548;
  assign n550 = ~n384 & ~po20;
  assign n551 = ~n412 & ~n428;
  assign n552 = ~n478 & n551;
  assign n553 = ~n546 & n552;
  assign n554 = ~n398 & ~n400;
  assign n555 = ~n397 & ~n554;
  assign n556 = ~n410 & n555;
  assign n557 = ~n548 & n556;
  assign n558 = ~n553 & n557;
  assign n559 = ~n550 & ~n558;
  assign n560 = n76 & ~n559;
  assign n561 = ~pi20 & ~n406;
  assign n562 = ~n408 & n561;
  assign n563 = ~pi01 & pi20;
  assign n564 = ~n527 & ~n563;
  assign n565 = ~n409 & n564;
  assign n566 = ~n562 & ~n565;
  assign n567 = pi01 & ~pi18;
  assign n568 = ~pi03 & ~n567;
  assign n569 = ~n566 & ~n568;
  assign n570 = ~n546 & n569;
  assign n571 = n552 & n570;
  assign n572 = pi03 & ~n567;
  assign n573 = ~n562 & ~n572;
  assign n574 = ~n565 & n573;
  assign n575 = ~n428 & n574;
  assign n576 = ~n412 & n575;
  assign n577 = n547 & n576;
  assign n578 = ~n403 & n574;
  assign n579 = ~n403 & n569;
  assign n580 = ~n578 & ~n579;
  assign n581 = ~n577 & n580;
  assign n582 = ~n571 & n581;
  assign n583 = n69 & ~n564;
  assign n584 = ~n572 & n583;
  assign n585 = n75 & n584;
  assign n586 = ~n400 & n585;
  assign n587 = ~n398 & n586;
  assign n588 = ~n397 & n587;
  assign n589 = ~n553 & n588;
  assign n590 = n71 & ~n527;
  assign n591 = ~n563 & n590;
  assign n592 = n119 & ~n568;
  assign n593 = n591 & n592;
  assign n594 = ~n400 & n593;
  assign n595 = ~n398 & n594;
  assign n596 = ~n397 & n595;
  assign n597 = ~n553 & n596;
  assign n598 = ~n589 & ~n597;
  assign n599 = n582 & n598;
  assign n600 = ~n538 & ~n541;
  assign n601 = ~pi05 & ~n406;
  assign n602 = ~n408 & n601;
  assign n603 = ~n600 & n602;
  assign n604 = ~n428 & n603;
  assign n605 = ~n412 & n604;
  assign n606 = n547 & n605;
  assign n607 = ~pi03 & ~n562;
  assign n608 = ~n565 & n607;
  assign n609 = ~n428 & n608;
  assign n610 = ~n412 & n609;
  assign n611 = n547 & n610;
  assign n612 = ~n403 & n608;
  assign n613 = ~n403 & n603;
  assign n614 = ~n612 & ~n613;
  assign n615 = ~n611 & n614;
  assign n616 = ~n606 & n615;
  assign n617 = ~pi03 & ~pi13;
  assign n618 = n101 & n617;
  assign n619 = n99 & n618;
  assign n620 = n67 & ~n564;
  assign n621 = n619 & n620;
  assign n622 = ~n400 & n621;
  assign n623 = ~n398 & n622;
  assign n624 = ~n397 & n623;
  assign n625 = ~n553 & n624;
  assign n626 = pi03 & ~pi05;
  assign n627 = n527 & ~n626;
  assign n628 = ~pi03 & ~pi05;
  assign n629 = ~n527 & ~n628;
  assign n630 = ~n627 & ~n629;
  assign n631 = ~n600 & ~n630;
  assign n632 = ~n527 & ~n626;
  assign n633 = n527 & ~n628;
  assign n634 = ~n632 & ~n633;
  assign n635 = ~n541 & ~n634;
  assign n636 = ~n538 & n635;
  assign n637 = ~n409 & ~n636;
  assign n638 = ~n631 & n637;
  assign n639 = n551 & ~n638;
  assign n640 = n547 & n639;
  assign n641 = ~n631 & ~n636;
  assign n642 = ~n410 & n641;
  assign n643 = ~n640 & n642;
  assign n644 = ~n625 & ~n643;
  assign n645 = n616 & n644;
  assign n646 = ~n599 & n645;
  assign n647 = n457 & ~n477;
  assign n648 = ~n436 & n647;
  assign n649 = ~n545 & n648;
  assign n650 = n547 & ~n649;
  assign n651 = pi09 & ~n410;
  assign n652 = ~n548 & n651;
  assign n653 = ~n650 & n652;
  assign n654 = pi05 & ~n541;
  assign n655 = ~n538 & n654;
  assign n656 = ~po20 & n655;
  assign n657 = ~n653 & ~n656;
  assign n658 = ~pi07 & ~n475;
  assign n659 = ~n471 & n658;
  assign n660 = ~n471 & ~n475;
  assign n661 = pi07 & ~n660;
  assign n662 = ~n659 & ~n661;
  assign n663 = ~po20 & ~n662;
  assign n664 = n520 & ~n544;
  assign n665 = ~pi07 & ~n545;
  assign n666 = ~n664 & n665;
  assign n667 = ~n545 & ~n664;
  assign n668 = pi07 & ~n667;
  assign n669 = ~n666 & ~n668;
  assign n670 = po20 & ~n669;
  assign n671 = ~n663 & ~n670;
  assign n672 = n657 & n671;
  assign n673 = ~pi09 & ~n478;
  assign n674 = ~n546 & n673;
  assign n675 = ~n410 & ~n649;
  assign n676 = n674 & n675;
  assign n677 = ~n548 & n676;
  assign n678 = ~pi03 & ~n600;
  assign n679 = pi03 & ~n541;
  assign n680 = ~n538 & n679;
  assign n681 = ~n678 & ~n680;
  assign n682 = ~n527 & ~n681;
  assign n683 = n527 & ~n680;
  assign n684 = ~n678 & n683;
  assign n685 = pi05 & ~n684;
  assign n686 = ~n682 & n685;
  assign n687 = ~n410 & n686;
  assign n688 = ~n548 & n687;
  assign n689 = ~n677 & ~n688;
  assign n690 = ~pi09 & ~n427;
  assign n691 = ~po20 & n690;
  assign n692 = pi09 & ~n417;
  assign n693 = ~n423 & n692;
  assign n694 = ~n426 & n693;
  assign n695 = ~po20 & n694;
  assign n696 = ~n691 & ~n695;
  assign n697 = n689 & n696;
  assign n698 = n672 & n697;
  assign n699 = ~n646 & n698;
  assign n700 = ~po20 & n659;
  assign n701 = ~n410 & n666;
  assign n702 = ~n548 & n701;
  assign n703 = ~n700 & ~n702;
  assign n704 = ~n653 & ~n695;
  assign n705 = ~n703 & n704;
  assign n706 = ~n397 & ~n412;
  assign n707 = ~n428 & ~n478;
  assign n708 = ~n546 & n707;
  assign n709 = n706 & ~n708;
  assign n710 = ~n546 & ~n706;
  assign n711 = n707 & n710;
  assign n712 = ~pi11 & ~n410;
  assign n713 = ~n548 & n712;
  assign n714 = ~n711 & n713;
  assign n715 = ~n709 & n714;
  assign n716 = n403 & ~n553;
  assign n717 = ~pi11 & ~n406;
  assign n718 = ~n408 & n717;
  assign n719 = ~n411 & n718;
  assign n720 = ~n716 & n719;
  assign n721 = ~n677 & ~n720;
  assign n722 = ~n691 & n721;
  assign n723 = ~n715 & n722;
  assign n724 = ~n705 & n723;
  assign n725 = ~n699 & n724;
  assign n726 = pi13 & ~n550;
  assign n727 = ~pi13 & ~n384;
  assign n728 = ~po20 & n727;
  assign n729 = ~n726 & ~n728;
  assign n730 = ~n558 & ~n729;
  assign n731 = n558 & ~n728;
  assign n732 = ~n726 & n731;
  assign n733 = po20 & ~n711;
  assign n734 = ~n709 & n733;
  assign n735 = n409 & ~n411;
  assign n736 = ~n716 & n735;
  assign n737 = pi11 & ~n736;
  assign n738 = ~n734 & n737;
  assign n739 = n99 & n101;
  assign n740 = n67 & n739;
  assign n741 = ~n738 & n740;
  assign n742 = ~n732 & n741;
  assign n743 = ~n730 & n742;
  assign n744 = ~n725 & n743;
  assign po18 = n560 | n744;
  assign n746 = ~n611 & ~n612;
  assign n747 = ~n625 & n746;
  assign n748 = ~n599 & n747;
  assign n749 = ~po20 & n600;
  assign n750 = ~n682 & ~n684;
  assign n751 = ~n410 & n750;
  assign n752 = ~n548 & n751;
  assign n753 = ~n749 & ~n752;
  assign n754 = ~pi05 & ~n753;
  assign n755 = pi05 & ~n752;
  assign n756 = ~n749 & n755;
  assign n757 = ~n754 & ~n756;
  assign n758 = ~n748 & ~n757;
  assign n759 = n748 & ~n756;
  assign n760 = ~n754 & n759;
  assign n761 = ~pi07 & ~n760;
  assign n762 = ~n758 & n761;
  assign n763 = ~n758 & ~n760;
  assign n764 = pi07 & ~n763;
  assign n765 = ~n762 & ~n764;
  assign n766 = po18 & ~n765;
  assign n767 = pi01 & ~pi16;
  assign n768 = pi18 & n767;
  assign n769 = po18 & n768;
  assign n770 = ~pi16 & n567;
  assign n771 = ~n560 & n770;
  assign n772 = ~n744 & n771;
  assign n773 = ~pi07 & ~n752;
  assign n774 = ~n749 & n773;
  assign n775 = pi07 & ~n753;
  assign n776 = ~n774 & ~n775;
  assign n777 = ~n560 & ~n776;
  assign n778 = ~n744 & n777;
  assign n779 = ~n772 & ~n778;
  assign n780 = ~n769 & n779;
  assign n781 = ~n766 & n780;
  assign n782 = pi03 & ~n560;
  assign n783 = ~n744 & n782;
  assign n784 = ~pi16 & n113;
  assign n785 = ~n572 & ~n784;
  assign n786 = ~n783 & n785;
  assign n787 = ~pi01 & pi18;
  assign n788 = pi18 & ~n784;
  assign n789 = ~n560 & n788;
  assign n790 = ~n744 & n789;
  assign n791 = ~n787 & ~n790;
  assign n792 = ~n786 & n791;
  assign n793 = n119 & n591;
  assign n794 = ~n400 & n793;
  assign n795 = ~n398 & n794;
  assign n796 = ~n397 & n795;
  assign n797 = ~n553 & n796;
  assign n798 = ~n566 & ~n716;
  assign n799 = ~n797 & ~n798;
  assign n800 = pi05 & ~n799;
  assign n801 = ~pi05 & ~n797;
  assign n802 = ~n798 & n801;
  assign n803 = ~n560 & ~n802;
  assign n804 = ~n800 & n803;
  assign n805 = ~n744 & n804;
  assign n806 = ~pi03 & pi05;
  assign n807 = ~n626 & ~n806;
  assign n808 = ~n567 & ~n807;
  assign n809 = n567 & ~n626;
  assign n810 = ~n806 & n809;
  assign n811 = ~n808 & ~n810;
  assign n812 = ~n797 & n811;
  assign n813 = ~n798 & n812;
  assign n814 = ~n799 & ~n811;
  assign n815 = ~n813 & ~n814;
  assign n816 = po18 & n815;
  assign n817 = ~n805 & ~n816;
  assign n818 = ~n792 & ~n817;
  assign n819 = n781 & n818;
  assign n820 = ~n560 & n802;
  assign n821 = ~n744 & n820;
  assign n822 = ~pi18 & n77;
  assign n823 = ~n572 & ~n822;
  assign n824 = ~n797 & n823;
  assign n825 = ~n798 & n824;
  assign n826 = ~n799 & ~n823;
  assign n827 = ~n825 & ~n826;
  assign n828 = ~pi05 & ~n827;
  assign n829 = po18 & n828;
  assign n830 = ~n821 & ~n829;
  assign n831 = ~n766 & ~n778;
  assign n832 = ~n830 & n831;
  assign n833 = po18 & n762;
  assign n834 = ~n656 & ~n688;
  assign n835 = ~n646 & n834;
  assign n836 = ~n671 & ~n835;
  assign n837 = n671 & n834;
  assign n838 = ~n646 & n837;
  assign n839 = ~pi09 & ~n838;
  assign n840 = ~n836 & n839;
  assign n841 = po18 & n840;
  assign n842 = ~po20 & ~n660;
  assign n843 = ~n410 & ~n667;
  assign n844 = ~n548 & n843;
  assign n845 = ~pi09 & ~n844;
  assign n846 = ~n842 & n845;
  assign n847 = ~n560 & n846;
  assign n848 = ~n744 & n847;
  assign n849 = ~n560 & n774;
  assign n850 = ~n744 & n849;
  assign n851 = ~n848 & ~n850;
  assign n852 = ~n841 & n851;
  assign n853 = ~n833 & n852;
  assign n854 = ~n832 & n853;
  assign n855 = ~n819 & n854;
  assign n856 = ~n734 & ~n736;
  assign n857 = ~n560 & n856;
  assign n858 = ~n744 & n857;
  assign n859 = ~n677 & ~n691;
  assign n860 = ~n705 & n859;
  assign n861 = ~n699 & n860;
  assign n862 = ~n715 & ~n720;
  assign n863 = ~n738 & n862;
  assign n864 = ~n861 & n863;
  assign n865 = n860 & ~n863;
  assign n866 = ~n699 & n865;
  assign n867 = ~n864 & ~n866;
  assign n868 = po18 & ~n867;
  assign n869 = ~n858 & ~n868;
  assign n870 = pi13 & ~n869;
  assign n871 = ~n836 & ~n838;
  assign n872 = pi09 & ~n871;
  assign n873 = po18 & n872;
  assign n874 = n704 & n859;
  assign n875 = ~n671 & n703;
  assign n876 = ~n874 & n875;
  assign n877 = n705 & n859;
  assign n878 = ~pi11 & ~n877;
  assign n879 = ~n876 & n878;
  assign n880 = n703 & ~n874;
  assign n881 = ~n835 & n880;
  assign n882 = ~n699 & ~n881;
  assign n883 = n879 & n882;
  assign n884 = po18 & n883;
  assign n885 = po20 & ~n650;
  assign n886 = n427 & ~po20;
  assign n887 = ~pi11 & ~n886;
  assign n888 = ~n885 & n887;
  assign n889 = ~n560 & n888;
  assign n890 = ~n744 & n889;
  assign n891 = ~n842 & ~n844;
  assign n892 = pi09 & ~n891;
  assign n893 = ~n560 & n892;
  assign n894 = ~n744 & n893;
  assign n895 = ~n890 & ~n894;
  assign n896 = ~n884 & n895;
  assign n897 = ~n873 & n896;
  assign n898 = ~pi13 & ~n858;
  assign n899 = ~n868 & n898;
  assign n900 = ~n876 & ~n877;
  assign n901 = ~n699 & n900;
  assign n902 = ~n881 & n901;
  assign n903 = po18 & n902;
  assign n904 = ~n885 & ~n886;
  assign n905 = ~n560 & n904;
  assign n906 = ~n744 & n905;
  assign n907 = pi11 & ~n906;
  assign n908 = ~n903 & n907;
  assign n909 = ~n899 & ~n908;
  assign n910 = n897 & n909;
  assign n911 = ~n870 & n910;
  assign n912 = ~n855 & n911;
  assign n913 = ~n884 & ~n890;
  assign n914 = ~n899 & n913;
  assign n915 = ~n870 & ~n914;
  assign n916 = ~n912 & ~n915;
  assign n917 = ~n730 & ~n732;
  assign n918 = ~n738 & ~n917;
  assign n919 = ~n725 & n918;
  assign n920 = po18 & n919;
  assign n921 = ~n559 & ~n560;
  assign n922 = ~n744 & n921;
  assign n923 = ~pi15 & ~n922;
  assign n924 = ~n920 & n923;
  assign n925 = ~n920 & ~n922;
  assign n926 = pi15 & ~n925;
  assign n927 = ~n924 & ~n926;
  assign n928 = ~pi01 & pi16;
  assign n929 = ~n767 & ~n928;
  assign n930 = n119 & ~n929;
  assign n931 = ~n927 & n930;
  assign n932 = ~n916 & n931;
  assign n933 = n740 & ~n925;
  assign n934 = ~pi16 & ~n933;
  assign n935 = n101 & ~n767;
  assign n936 = ~n928 & n935;
  assign n937 = n180 & n936;
  assign n938 = ~n925 & n937;
  assign n939 = ~n915 & ~n938;
  assign n940 = ~n934 & n939;
  assign n941 = ~n912 & n940;
  assign n942 = n119 & ~n927;
  assign n943 = ~n934 & ~n938;
  assign n944 = ~n942 & n943;
  assign n945 = ~n941 & ~n944;
  assign n946 = ~n932 & n945;
  assign n947 = ~pi03 & ~n946;
  assign n948 = pi03 & ~n944;
  assign n949 = ~n941 & n948;
  assign n950 = ~n932 & n949;
  assign n951 = ~n947 & ~n950;
  assign n952 = ~n70 & ~n951;
  assign n953 = n70 & ~n950;
  assign n954 = ~n947 & n953;
  assign n955 = ~n952 & ~n954;
  assign n956 = pi01 & po18;
  assign n957 = pi18 & ~n956;
  assign n958 = n567 & po18;
  assign n959 = ~n957 & ~n958;
  assign n960 = ~pi03 & ~n959;
  assign n961 = pi03 & ~n958;
  assign n962 = ~n957 & n961;
  assign n963 = ~n960 & ~n962;
  assign n964 = ~n767 & ~n963;
  assign n965 = n767 & ~n962;
  assign n966 = ~n960 & n965;
  assign n967 = ~n964 & ~n966;
  assign n968 = ~n915 & ~n933;
  assign n969 = ~n912 & n968;
  assign n970 = ~n933 & ~n942;
  assign n971 = ~pi05 & ~n970;
  assign n972 = ~n969 & n971;
  assign n973 = ~n967 & n972;
  assign n974 = ~pi03 & ~n70;
  assign n975 = ~n944 & n974;
  assign n976 = ~n941 & n975;
  assign n977 = ~n932 & n976;
  assign po16 = ~n969 & ~n970;
  assign n979 = ~pi05 & ~n959;
  assign n980 = ~po16 & n979;
  assign n981 = ~n977 & ~n980;
  assign n982 = ~n973 & n981;
  assign n983 = pi03 & ~n70;
  assign n984 = ~n946 & n983;
  assign n985 = ~n947 & ~n984;
  assign n986 = n982 & n985;
  assign n987 = pi05 & ~n958;
  assign n988 = ~n957 & n987;
  assign n989 = ~po16 & n988;
  assign n990 = pi05 & ~n966;
  assign n991 = ~n970 & n990;
  assign n992 = ~n964 & n991;
  assign n993 = ~n969 & n992;
  assign n994 = ~n989 & ~n993;
  assign n995 = po18 & ~n763;
  assign n996 = ~n560 & ~n753;
  assign n997 = ~n744 & n996;
  assign n998 = ~pi09 & ~n997;
  assign n999 = ~n995 & n998;
  assign n1000 = ~n995 & ~n997;
  assign n1001 = pi09 & ~n1000;
  assign n1002 = ~n999 & ~n1001;
  assign n1003 = ~po16 & ~n1002;
  assign n1004 = ~n769 & ~n772;
  assign n1005 = ~n792 & n1004;
  assign n1006 = ~n817 & n1005;
  assign n1007 = n830 & ~n831;
  assign n1008 = ~n1006 & n1007;
  assign n1009 = ~pi09 & ~n832;
  assign n1010 = ~n819 & n1009;
  assign n1011 = ~n1008 & n1010;
  assign n1012 = ~n819 & ~n832;
  assign n1013 = ~n1008 & n1012;
  assign n1014 = pi09 & ~n1013;
  assign n1015 = ~n1011 & ~n1014;
  assign n1016 = po16 & ~n1015;
  assign n1017 = ~n1003 & ~n1016;
  assign n1018 = po18 & n827;
  assign n1019 = ~n560 & ~n799;
  assign n1020 = ~n744 & n1019;
  assign n1021 = ~pi07 & ~n1020;
  assign n1022 = ~n1018 & n1021;
  assign n1023 = ~n1018 & ~n1020;
  assign n1024 = pi07 & ~n1023;
  assign n1025 = ~n1022 & ~n1024;
  assign n1026 = ~po16 & ~n1025;
  assign n1027 = n817 & ~n1005;
  assign n1028 = ~pi07 & ~n1006;
  assign n1029 = ~n1027 & n1028;
  assign n1030 = ~n1006 & ~n1027;
  assign n1031 = pi07 & ~n1030;
  assign n1032 = ~n1029 & ~n1031;
  assign n1033 = po16 & ~n1032;
  assign n1034 = ~n1026 & ~n1033;
  assign n1035 = n1017 & n1034;
  assign n1036 = n994 & n1035;
  assign n1037 = ~n986 & n1036;
  assign n1038 = n869 & ~n933;
  assign n1039 = ~n942 & n1038;
  assign n1040 = ~n915 & n1038;
  assign n1041 = ~n912 & n1040;
  assign n1042 = ~n1039 & ~n1041;
  assign n1043 = ~pi15 & ~n1042;
  assign n1044 = ~n970 & n1011;
  assign n1045 = ~n969 & n1044;
  assign n1046 = ~n1043 & ~n1045;
  assign n1047 = n897 & ~n908;
  assign n1048 = ~n855 & n1047;
  assign n1049 = ~n870 & ~n899;
  assign n1050 = ~n913 & ~n1049;
  assign n1051 = ~n870 & n914;
  assign n1052 = ~n1050 & ~n1051;
  assign n1053 = ~n1048 & ~n1052;
  assign n1054 = n1047 & ~n1051;
  assign n1055 = ~n855 & n1054;
  assign n1056 = ~n1050 & n1055;
  assign n1057 = ~n1053 & ~n1056;
  assign n1058 = n740 & ~n969;
  assign n1059 = ~n1057 & n1058;
  assign n1060 = ~po16 & n999;
  assign n1061 = ~n1059 & ~n1060;
  assign n1062 = po18 & ~n871;
  assign n1063 = ~n560 & ~n891;
  assign n1064 = ~n744 & n1063;
  assign n1065 = ~pi11 & ~n1064;
  assign n1066 = ~n1062 & n1065;
  assign n1067 = ~po16 & n1066;
  assign n1068 = ~n848 & ~n894;
  assign n1069 = ~n841 & n1068;
  assign n1070 = ~n873 & n1069;
  assign n1071 = ~n833 & ~n850;
  assign n1072 = ~n832 & n1071;
  assign n1073 = ~n1070 & n1072;
  assign n1074 = ~n819 & n1073;
  assign n1075 = ~n819 & n1072;
  assign n1076 = n1070 & ~n1075;
  assign n1077 = ~n1074 & ~n1076;
  assign n1078 = ~pi11 & ~n970;
  assign n1079 = n1077 & n1078;
  assign n1080 = ~n969 & n1079;
  assign n1081 = ~n1067 & ~n1080;
  assign n1082 = n1061 & n1081;
  assign n1083 = n1046 & n1082;
  assign n1084 = po16 & ~n1057;
  assign n1085 = pi15 & ~n1039;
  assign n1086 = ~n1041 & n1085;
  assign n1087 = ~n1084 & n1086;
  assign n1088 = ~n908 & n913;
  assign n1089 = ~n873 & ~n894;
  assign n1090 = ~n855 & n1089;
  assign n1091 = ~n1088 & ~n1090;
  assign n1092 = ~n1048 & ~n1091;
  assign n1093 = po16 & ~n1092;
  assign n1094 = ~n903 & ~n906;
  assign n1095 = ~n933 & n1094;
  assign n1096 = ~n915 & n1095;
  assign n1097 = ~n912 & n1096;
  assign n1098 = ~n942 & n1095;
  assign n1099 = ~pi13 & ~n1098;
  assign n1100 = ~n1097 & n1099;
  assign n1101 = ~n1093 & n1100;
  assign n1102 = ~n1087 & n1101;
  assign n1103 = ~po16 & n1022;
  assign n1104 = ~n970 & n1029;
  assign n1105 = ~n969 & n1104;
  assign n1106 = ~n1103 & ~n1105;
  assign n1107 = n1017 & ~n1106;
  assign n1108 = ~n1102 & ~n1107;
  assign n1109 = n1083 & n1108;
  assign n1110 = ~n1037 & n1109;
  assign n1111 = ~n1097 & ~n1098;
  assign n1112 = ~n1093 & n1111;
  assign n1113 = ~pi13 & ~n1112;
  assign n1114 = pi13 & ~n1098;
  assign n1115 = ~n1097 & n1114;
  assign n1116 = ~n1093 & n1115;
  assign n1117 = ~n1113 & ~n1116;
  assign n1118 = ~n1043 & ~n1059;
  assign n1119 = ~n1062 & ~n1064;
  assign n1120 = pi11 & ~n1119;
  assign n1121 = ~po16 & n1120;
  assign n1122 = pi11 & ~n970;
  assign n1123 = ~n969 & n1122;
  assign n1124 = ~n1077 & n1123;
  assign n1125 = ~n1121 & ~n1124;
  assign n1126 = n1118 & n1125;
  assign n1127 = ~n1087 & n1126;
  assign n1128 = ~n1117 & n1127;
  assign n1129 = ~n1102 & n1118;
  assign n1130 = ~n1128 & n1129;
  assign n1131 = n927 & ~n970;
  assign n1132 = ~n969 & n1131;
  assign n1133 = ~n916 & n1132;
  assign n1134 = ~n925 & ~po16;
  assign n1135 = ~pi17 & ~n1134;
  assign n1136 = ~n1133 & n1135;
  assign n1137 = ~n1133 & ~n1134;
  assign n1138 = pi17 & ~n1137;
  assign n1139 = ~n1136 & ~n1138;
  assign n1140 = n180 & ~n1139;
  assign n1141 = ~n1130 & n1140;
  assign n1142 = ~n1110 & n1141;
  assign n1143 = n119 & ~n1137;
  assign po14 = n1142 | n1143;
  assign n1145 = n955 & po14;
  assign n1146 = n946 & ~n1143;
  assign n1147 = ~n1142 & n1146;
  assign n1148 = ~n1145 & ~n1147;
  assign n1149 = pi05 & ~n1148;
  assign n1150 = pi01 & ~pi17;
  assign n1151 = n99 & n1150;
  assign n1152 = n67 & n1151;
  assign n1153 = ~n1137 & n1152;
  assign n1154 = ~pi14 & ~n1153;
  assign n1155 = pi14 & ~pi19;
  assign n1156 = n73 & n1155;
  assign n1157 = n1150 & n1156;
  assign n1158 = n69 & n1157;
  assign n1159 = ~n1137 & n1158;
  assign n1160 = ~n1154 & ~n1159;
  assign n1161 = pi01 & ~pi12;
  assign n1162 = ~pi03 & ~n1161;
  assign n1163 = ~n1160 & ~n1162;
  assign n1164 = ~n1142 & n1163;
  assign n1165 = pi03 & ~n1161;
  assign n1166 = ~n1159 & ~n1165;
  assign n1167 = ~n1154 & n1166;
  assign n1168 = ~n1142 & n1167;
  assign n1169 = ~pi01 & pi14;
  assign n1170 = ~n70 & ~n1169;
  assign n1171 = ~n1165 & ~n1170;
  assign n1172 = n180 & n1171;
  assign n1173 = ~n1139 & n1172;
  assign n1174 = ~n1130 & n1173;
  assign n1175 = ~n1110 & n1174;
  assign n1176 = n99 & n1170;
  assign n1177 = n67 & ~n1162;
  assign n1178 = n1176 & n1177;
  assign n1179 = ~n1139 & n1178;
  assign n1180 = ~n1130 & n1179;
  assign n1181 = ~n1110 & n1180;
  assign n1182 = ~n1175 & ~n1181;
  assign n1183 = ~n1168 & n1182;
  assign n1184 = ~n1164 & n1183;
  assign n1185 = ~pi05 & ~pi19;
  assign n1186 = n73 & n1185;
  assign n1187 = n69 & n1186;
  assign n1188 = ~n1139 & n1187;
  assign n1189 = ~n955 & n1188;
  assign n1190 = ~n1130 & n1189;
  assign n1191 = ~n1110 & n1190;
  assign n1192 = ~pi03 & ~pi19;
  assign n1193 = n73 & n1192;
  assign n1194 = n69 & n1193;
  assign n1195 = ~n1170 & n1194;
  assign n1196 = ~n1139 & n1195;
  assign n1197 = ~n1130 & n1196;
  assign n1198 = ~n1110 & n1197;
  assign n1199 = ~pi05 & ~pi17;
  assign n1200 = n99 & n1199;
  assign n1201 = n67 & n1200;
  assign n1202 = ~n1137 & n1201;
  assign n1203 = ~n955 & n1202;
  assign n1204 = ~n1198 & ~n1203;
  assign n1205 = ~n1191 & n1204;
  assign n1206 = ~pi03 & ~n1159;
  assign n1207 = ~n1154 & n1206;
  assign n1208 = ~n1142 & n1207;
  assign n1209 = ~pi05 & ~n946;
  assign n1210 = ~n1143 & n1209;
  assign n1211 = ~n1142 & n1210;
  assign n1212 = ~n1208 & ~n1211;
  assign n1213 = n1205 & n1212;
  assign n1214 = ~n1184 & n1213;
  assign n1215 = ~n977 & ~n984;
  assign n1216 = ~n947 & n1215;
  assign n1217 = n959 & ~po16;
  assign n1218 = n967 & po16;
  assign n1219 = ~n1217 & ~n1218;
  assign n1220 = ~pi05 & ~n1219;
  assign n1221 = pi05 & ~n1217;
  assign n1222 = ~n1218 & n1221;
  assign n1223 = ~n1220 & ~n1222;
  assign n1224 = ~n1216 & ~n1223;
  assign n1225 = n1216 & n1223;
  assign n1226 = ~pi07 & ~n1225;
  assign n1227 = ~n1224 & n1226;
  assign n1228 = ~n1224 & ~n1225;
  assign n1229 = pi07 & ~n1228;
  assign n1230 = ~n1227 & ~n1229;
  assign n1231 = po14 & ~n1230;
  assign n1232 = ~n986 & n994;
  assign n1233 = ~n1034 & ~n1232;
  assign n1234 = n994 & n1034;
  assign n1235 = ~n986 & n1234;
  assign n1236 = ~pi09 & ~n1235;
  assign n1237 = ~n1233 & n1236;
  assign n1238 = ~n1233 & ~n1235;
  assign n1239 = pi09 & ~n1238;
  assign n1240 = ~n1237 & ~n1239;
  assign n1241 = po14 & ~n1240;
  assign n1242 = ~po16 & ~n1023;
  assign n1243 = ~n970 & ~n1030;
  assign n1244 = ~n969 & n1243;
  assign n1245 = ~pi09 & ~n1244;
  assign n1246 = ~n1242 & n1245;
  assign n1247 = ~n1242 & ~n1244;
  assign n1248 = pi09 & ~n1247;
  assign n1249 = ~n1246 & ~n1248;
  assign n1250 = ~n1143 & ~n1249;
  assign n1251 = ~n1142 & n1250;
  assign n1252 = ~pi07 & ~n1217;
  assign n1253 = ~n1218 & n1252;
  assign n1254 = pi07 & ~n1219;
  assign n1255 = ~n1253 & ~n1254;
  assign n1256 = ~n1143 & ~n1255;
  assign n1257 = ~n1142 & n1256;
  assign n1258 = ~n1251 & ~n1257;
  assign n1259 = ~n1241 & n1258;
  assign n1260 = ~n1231 & n1259;
  assign n1261 = ~n1214 & n1260;
  assign n1262 = ~n1149 & n1261;
  assign n1263 = ~n1143 & n1253;
  assign n1264 = ~n1142 & n1263;
  assign n1265 = po14 & n1227;
  assign n1266 = ~n1264 & ~n1265;
  assign n1267 = ~n1241 & ~n1251;
  assign n1268 = ~n1266 & n1267;
  assign n1269 = n1106 & ~n1235;
  assign n1270 = n1017 & ~n1269;
  assign n1271 = ~n1017 & n1106;
  assign n1272 = ~n1235 & n1271;
  assign n1273 = ~pi11 & ~n1272;
  assign n1274 = ~n1270 & n1273;
  assign n1275 = po14 & n1274;
  assign n1276 = po14 & n1237;
  assign n1277 = ~n1143 & n1246;
  assign n1278 = ~n1142 & n1277;
  assign n1279 = ~po16 & ~n1000;
  assign n1280 = ~n970 & ~n1013;
  assign n1281 = ~n969 & n1280;
  assign n1282 = ~pi11 & ~n1281;
  assign n1283 = ~n1279 & n1282;
  assign n1284 = ~n1143 & n1283;
  assign n1285 = ~n1142 & n1284;
  assign n1286 = ~n1278 & ~n1285;
  assign n1287 = ~n1276 & n1286;
  assign n1288 = ~n1275 & n1287;
  assign n1289 = ~n1268 & n1288;
  assign n1290 = ~n1262 & n1289;
  assign n1291 = n994 & n1125;
  assign n1292 = n1035 & n1291;
  assign n1293 = ~n986 & n1292;
  assign n1294 = ~n1045 & ~n1060;
  assign n1295 = n1081 & n1294;
  assign n1296 = ~n1107 & n1295;
  assign n1297 = n1125 & ~n1296;
  assign n1298 = ~n1293 & ~n1297;
  assign n1299 = ~n1117 & ~n1298;
  assign n1300 = n1117 & ~n1293;
  assign n1301 = ~n1297 & n1300;
  assign n1302 = ~n1299 & ~n1301;
  assign n1303 = pi15 & ~n1302;
  assign n1304 = po14 & n1303;
  assign n1305 = ~pi15 & ~n1299;
  assign n1306 = ~n1301 & n1305;
  assign n1307 = po14 & n1306;
  assign n1308 = ~pi15 & ~n1098;
  assign n1309 = ~n1097 & n1308;
  assign n1310 = ~n1093 & n1309;
  assign n1311 = ~n1143 & n1310;
  assign n1312 = ~n1142 & n1311;
  assign n1313 = pi15 & ~n1112;
  assign n1314 = ~n1143 & n1313;
  assign n1315 = ~n1142 & n1314;
  assign n1316 = ~n1312 & ~n1315;
  assign n1317 = ~n1307 & n1316;
  assign n1318 = ~n1304 & n1317;
  assign n1319 = ~n1107 & n1294;
  assign n1320 = ~n1037 & n1319;
  assign n1321 = ~po16 & ~n1119;
  assign n1322 = po16 & ~n1077;
  assign n1323 = ~n1321 & ~n1322;
  assign n1324 = ~pi11 & ~n1323;
  assign n1325 = pi11 & ~n1321;
  assign n1326 = ~n1322 & n1325;
  assign n1327 = ~n1324 & ~n1326;
  assign n1328 = ~pi13 & ~n1327;
  assign n1329 = pi13 & ~n1324;
  assign n1330 = ~n1326 & n1329;
  assign n1331 = ~n1328 & ~n1330;
  assign n1332 = ~n1320 & ~n1331;
  assign n1333 = n1320 & n1331;
  assign n1334 = ~n1332 & ~n1333;
  assign n1335 = po14 & n1334;
  assign n1336 = ~n1270 & ~n1272;
  assign n1337 = pi11 & ~n1336;
  assign n1338 = po14 & n1337;
  assign n1339 = ~n1279 & ~n1281;
  assign n1340 = pi11 & ~n1339;
  assign n1341 = ~n1143 & n1340;
  assign n1342 = ~n1142 & n1341;
  assign n1343 = ~pi13 & ~n1321;
  assign n1344 = ~n1322 & n1343;
  assign n1345 = pi13 & ~n1323;
  assign n1346 = ~n1344 & ~n1345;
  assign n1347 = ~n1143 & ~n1346;
  assign n1348 = ~n1142 & n1347;
  assign n1349 = ~n1342 & ~n1348;
  assign n1350 = ~n1338 & n1349;
  assign n1351 = ~n1335 & n1350;
  assign n1352 = ~n1318 & n1351;
  assign n1353 = ~n1290 & n1352;
  assign n1354 = ~n1275 & ~n1307;
  assign n1355 = ~n1304 & n1316;
  assign n1356 = n1354 & n1355;
  assign n1357 = ~n1143 & n1344;
  assign n1358 = ~n1142 & n1357;
  assign n1359 = ~n1320 & ~n1327;
  assign n1360 = n1319 & n1327;
  assign n1361 = ~n1037 & n1360;
  assign n1362 = ~pi13 & ~n1361;
  assign n1363 = ~n1359 & n1362;
  assign n1364 = po14 & n1363;
  assign n1365 = ~n1358 & ~n1364;
  assign n1366 = n1287 & n1365;
  assign n1367 = n1356 & n1366;
  assign n1368 = ~n1268 & n1367;
  assign n1369 = ~n1262 & n1368;
  assign n1370 = ~n1318 & ~n1365;
  assign n1371 = ~n1304 & ~n1307;
  assign n1372 = n1316 & n1371;
  assign n1373 = n1365 & n1372;
  assign n1374 = ~n1351 & n1373;
  assign n1375 = ~n1370 & ~n1374;
  assign n1376 = ~n1369 & n1375;
  assign n1377 = ~n1353 & n1376;
  assign n1378 = pi17 & ~pi19;
  assign n1379 = n73 & n1378;
  assign n1380 = n69 & n1379;
  assign n1381 = ~n1130 & n1380;
  assign n1382 = ~n1110 & n1381;
  assign n1383 = ~n1110 & ~n1130;
  assign n1384 = n119 & ~n1383;
  assign n1385 = ~n1137 & ~n1384;
  assign n1386 = ~n1382 & n1385;
  assign n1387 = ~n180 & ~n1386;
  assign n1388 = n1316 & n1349;
  assign n1389 = pi19 & ~pi21;
  assign n1390 = n98 & n1389;
  assign n1391 = n67 & n1390;
  assign n1392 = ~n1137 & ~n1391;
  assign n1393 = ~n1384 & n1392;
  assign n1394 = ~n1382 & n1393;
  assign n1395 = ~n1307 & ~n1394;
  assign n1396 = n1388 & n1395;
  assign n1397 = ~n1387 & n1396;
  assign n1398 = n1042 & ~n1084;
  assign n1399 = ~n1143 & n1398;
  assign n1400 = ~n1142 & n1399;
  assign n1401 = ~n1087 & n1118;
  assign n1402 = ~n1101 & ~n1401;
  assign n1403 = n1101 & n1401;
  assign n1404 = ~n1402 & ~n1403;
  assign n1405 = ~n1299 & n1404;
  assign n1406 = ~n1117 & ~n1401;
  assign n1407 = ~n1298 & n1406;
  assign n1408 = ~n1405 & ~n1407;
  assign n1409 = po14 & n1408;
  assign n1410 = ~n1400 & ~n1409;
  assign n1411 = pi17 & ~n1410;
  assign n1412 = ~n1304 & ~n1338;
  assign n1413 = ~n1335 & n1412;
  assign n1414 = ~n1411 & n1413;
  assign n1415 = n1397 & n1414;
  assign n1416 = ~n1290 & n1415;
  assign n1417 = ~n1387 & ~n1394;
  assign n1418 = ~n1411 & n1417;
  assign n1419 = n180 & ~n1137;
  assign n1420 = ~n1384 & n1419;
  assign n1421 = ~n1382 & n1420;
  assign n1422 = ~n1418 & ~n1421;
  assign n1423 = n1318 & ~n1365;
  assign n1424 = ~pi17 & ~n1400;
  assign n1425 = ~n1409 & n1424;
  assign n1426 = ~n1307 & ~n1312;
  assign n1427 = ~n1421 & n1426;
  assign n1428 = ~n1425 & n1427;
  assign n1429 = ~n1423 & n1428;
  assign n1430 = ~n1422 & ~n1429;
  assign po12 = n1416 | n1430;
  assign n1432 = pi17 & po12;
  assign n1433 = ~n1377 & n1432;
  assign n1434 = ~pi17 & ~n1422;
  assign n1435 = ~n1429 & n1434;
  assign n1436 = ~n1315 & ~n1342;
  assign n1437 = ~n1348 & n1436;
  assign n1438 = ~pi17 & ~n1312;
  assign n1439 = ~n1394 & n1438;
  assign n1440 = n1437 & n1439;
  assign n1441 = ~n1387 & n1440;
  assign n1442 = ~n1335 & ~n1338;
  assign n1443 = n1371 & n1442;
  assign n1444 = ~n1411 & n1443;
  assign n1445 = n1441 & n1444;
  assign n1446 = ~n1290 & n1445;
  assign n1447 = ~n1435 & ~n1446;
  assign n1448 = n1377 & ~n1447;
  assign n1449 = po14 & ~n1302;
  assign n1450 = ~n1112 & ~n1143;
  assign n1451 = ~n1142 & n1450;
  assign n1452 = ~pi17 & ~n1451;
  assign n1453 = ~n1449 & n1452;
  assign n1454 = ~n1449 & ~n1451;
  assign n1455 = pi17 & ~n1454;
  assign n1456 = ~n1453 & ~n1455;
  assign n1457 = ~n1430 & n1456;
  assign n1458 = ~n1416 & n1457;
  assign n1459 = ~n1448 & ~n1458;
  assign n1460 = ~n1433 & n1459;
  assign n1461 = ~n1143 & n1323;
  assign n1462 = ~n1142 & n1461;
  assign n1463 = ~n1359 & ~n1361;
  assign n1464 = po14 & n1463;
  assign n1465 = ~n1462 & ~n1464;
  assign n1466 = ~n1430 & n1465;
  assign n1467 = ~n1416 & n1466;
  assign n1468 = ~n1338 & ~n1342;
  assign n1469 = ~n1289 & n1468;
  assign n1470 = n1260 & n1468;
  assign n1471 = ~n1149 & ~n1214;
  assign n1472 = n1470 & n1471;
  assign n1473 = ~n1469 & ~n1472;
  assign n1474 = ~n1335 & ~n1348;
  assign n1475 = ~n1473 & n1474;
  assign n1476 = ~n1469 & ~n1474;
  assign n1477 = ~n1472 & n1476;
  assign n1478 = ~n1475 & ~n1477;
  assign n1479 = po12 & ~n1478;
  assign n1480 = ~n1467 & ~n1479;
  assign n1481 = pi15 & ~n1480;
  assign n1482 = ~n1460 & ~n1481;
  assign n1483 = ~n1304 & ~n1315;
  assign n1484 = ~n1365 & n1483;
  assign n1485 = n1388 & n1443;
  assign n1486 = ~n1484 & n1485;
  assign n1487 = ~n1290 & n1486;
  assign n1488 = n1426 & ~n1484;
  assign n1489 = ~n1411 & ~n1425;
  assign n1490 = ~n1488 & ~n1489;
  assign n1491 = ~n1425 & n1426;
  assign n1492 = ~n1411 & n1491;
  assign n1493 = ~n1484 & n1492;
  assign n1494 = ~n1490 & ~n1493;
  assign n1495 = ~n1487 & ~n1494;
  assign n1496 = n1486 & ~n1490;
  assign n1497 = ~n1493 & n1496;
  assign n1498 = ~n1290 & n1497;
  assign n1499 = ~n1495 & ~n1498;
  assign n1500 = ~n1423 & n1491;
  assign n1501 = n1418 & ~n1500;
  assign n1502 = n1410 & ~n1421;
  assign n1503 = ~n1501 & n1502;
  assign n1504 = ~n1416 & n1503;
  assign n1505 = po12 & ~n1504;
  assign n1506 = ~n1499 & n1505;
  assign n1507 = pi19 & ~n1504;
  assign n1508 = ~pi19 & ~n1400;
  assign n1509 = ~n1409 & n1508;
  assign n1510 = ~n1421 & n1509;
  assign n1511 = ~n1501 & n1510;
  assign n1512 = ~n1416 & n1511;
  assign n1513 = ~n1507 & ~n1512;
  assign n1514 = ~n1506 & ~n1513;
  assign n1515 = n1506 & n1513;
  assign n1516 = ~n1514 & ~n1515;
  assign n1517 = n1482 & n1516;
  assign n1518 = po12 & ~n1499;
  assign n1519 = ~n1504 & ~n1518;
  assign n1520 = ~pi19 & ~n1519;
  assign n1521 = ~n1447 & ~n1499;
  assign n1522 = ~pi17 & ~n1507;
  assign n1523 = ~n1521 & ~n1522;
  assign n1524 = ~n1430 & ~n1454;
  assign n1525 = ~n1416 & n1524;
  assign n1526 = n1377 & po12;
  assign n1527 = ~n1525 & ~n1526;
  assign n1528 = ~n1523 & n1527;
  assign n1529 = ~n1520 & ~n1528;
  assign n1530 = ~n1517 & n1529;
  assign n1531 = ~n1142 & ~n1160;
  assign n1532 = n67 & n1176;
  assign n1533 = ~n1139 & n1532;
  assign n1534 = ~n1130 & n1533;
  assign n1535 = ~n1110 & n1534;
  assign n1536 = ~pi12 & n77;
  assign n1537 = ~n1165 & ~n1536;
  assign n1538 = ~n1535 & n1537;
  assign n1539 = ~n1531 & n1538;
  assign n1540 = ~n1531 & ~n1535;
  assign n1541 = ~n1537 & ~n1540;
  assign n1542 = ~n1539 & ~n1541;
  assign n1543 = ~pi05 & ~n1542;
  assign n1544 = pi05 & ~n1539;
  assign n1545 = ~n1541 & n1544;
  assign n1546 = ~n1543 & ~n1545;
  assign n1547 = po12 & ~n1546;
  assign n1548 = pi01 & ~pi10;
  assign n1549 = pi12 & n1548;
  assign n1550 = po12 & n1549;
  assign n1551 = ~pi05 & ~n1147;
  assign n1552 = ~n1145 & n1551;
  assign n1553 = ~n1198 & ~n1208;
  assign n1554 = ~n1184 & n1553;
  assign n1555 = ~n1552 & n1554;
  assign n1556 = ~n1149 & n1555;
  assign n1557 = ~n1149 & ~n1552;
  assign n1558 = ~n1554 & ~n1557;
  assign n1559 = ~n1556 & ~n1558;
  assign n1560 = ~pi07 & ~n1559;
  assign n1561 = pi07 & ~n1556;
  assign n1562 = ~n1558 & n1561;
  assign n1563 = ~n1560 & ~n1562;
  assign n1564 = po12 & ~n1563;
  assign n1565 = ~n1550 & ~n1564;
  assign n1566 = ~n1547 & n1565;
  assign n1567 = pi03 & ~n1421;
  assign n1568 = ~n1501 & n1567;
  assign n1569 = ~n1416 & n1568;
  assign n1570 = ~pi10 & n113;
  assign n1571 = ~n1165 & ~n1570;
  assign n1572 = ~n1569 & n1571;
  assign n1573 = ~pi01 & pi12;
  assign n1574 = pi12 & ~n1570;
  assign n1575 = ~n1421 & n1574;
  assign n1576 = ~n1501 & n1575;
  assign n1577 = ~n1416 & n1576;
  assign n1578 = ~n1573 & ~n1577;
  assign n1579 = ~n1572 & n1578;
  assign n1580 = ~pi05 & ~n1535;
  assign n1581 = ~n1531 & n1580;
  assign n1582 = pi05 & ~n1540;
  assign n1583 = ~n1581 & ~n1582;
  assign n1584 = ~n1430 & ~n1583;
  assign n1585 = ~n1416 & n1584;
  assign n1586 = ~pi10 & n1161;
  assign n1587 = ~n1430 & n1586;
  assign n1588 = ~n1416 & n1587;
  assign n1589 = ~pi07 & ~n1147;
  assign n1590 = ~n1145 & n1589;
  assign n1591 = pi07 & ~n1148;
  assign n1592 = ~n1590 & ~n1591;
  assign n1593 = ~n1430 & ~n1592;
  assign n1594 = ~n1416 & n1593;
  assign n1595 = ~n1588 & ~n1594;
  assign n1596 = ~n1585 & n1595;
  assign n1597 = ~n1579 & n1596;
  assign n1598 = n1566 & n1597;
  assign n1599 = ~n1430 & n1581;
  assign n1600 = ~n1416 & n1599;
  assign n1601 = po12 & n1543;
  assign n1602 = ~n1600 & ~n1601;
  assign n1603 = ~n1564 & ~n1594;
  assign n1604 = ~n1602 & n1603;
  assign n1605 = po12 & n1560;
  assign n1606 = ~n1231 & ~n1257;
  assign n1607 = ~n1214 & n1606;
  assign n1608 = ~n1149 & n1607;
  assign n1609 = ~n1471 & ~n1606;
  assign n1610 = ~pi09 & ~n1609;
  assign n1611 = ~n1608 & n1610;
  assign n1612 = po12 & n1611;
  assign n1613 = po14 & ~n1228;
  assign n1614 = ~n1143 & ~n1219;
  assign n1615 = ~n1142 & n1614;
  assign n1616 = ~pi09 & ~n1615;
  assign n1617 = ~n1613 & n1616;
  assign n1618 = ~n1430 & n1617;
  assign n1619 = ~n1416 & n1618;
  assign n1620 = ~n1430 & n1590;
  assign n1621 = ~n1416 & n1620;
  assign n1622 = ~n1619 & ~n1621;
  assign n1623 = ~n1612 & n1622;
  assign n1624 = ~n1605 & n1623;
  assign n1625 = ~n1604 & n1624;
  assign n1626 = ~n1598 & n1625;
  assign n1627 = ~n1276 & ~n1278;
  assign n1628 = ~n1268 & n1627;
  assign n1629 = ~n1283 & ~n1340;
  assign n1630 = ~n1143 & ~n1629;
  assign n1631 = ~n1142 & n1630;
  assign n1632 = ~n1275 & ~n1631;
  assign n1633 = ~n1338 & n1632;
  assign n1634 = n1628 & ~n1633;
  assign n1635 = ~n1262 & n1634;
  assign n1636 = ~n1628 & n1633;
  assign n1637 = n1258 & ~n1631;
  assign n1638 = ~n1231 & ~n1241;
  assign n1639 = ~n1275 & ~n1338;
  assign n1640 = n1638 & n1639;
  assign n1641 = n1637 & n1640;
  assign n1642 = n1471 & n1641;
  assign n1643 = ~pi13 & ~n1642;
  assign n1644 = ~n1636 & n1643;
  assign n1645 = ~n1635 & n1644;
  assign n1646 = ~n1636 & ~n1642;
  assign n1647 = ~n1635 & n1646;
  assign n1648 = pi13 & ~n1647;
  assign n1649 = ~n1645 & ~n1648;
  assign n1650 = po12 & ~n1649;
  assign n1651 = po14 & ~n1238;
  assign n1652 = ~n1143 & ~n1247;
  assign n1653 = ~n1142 & n1652;
  assign n1654 = ~pi11 & ~n1653;
  assign n1655 = ~n1651 & n1654;
  assign n1656 = ~n1651 & ~n1653;
  assign n1657 = pi11 & ~n1656;
  assign n1658 = ~n1655 & ~n1657;
  assign n1659 = ~n1430 & ~n1658;
  assign n1660 = ~n1416 & n1659;
  assign n1661 = po14 & ~n1336;
  assign n1662 = ~n1143 & ~n1339;
  assign n1663 = ~n1142 & n1662;
  assign n1664 = ~pi13 & ~n1663;
  assign n1665 = ~n1661 & n1664;
  assign n1666 = ~n1661 & ~n1663;
  assign n1667 = pi13 & ~n1666;
  assign n1668 = ~n1665 & ~n1667;
  assign n1669 = ~n1430 & ~n1668;
  assign n1670 = ~n1416 & n1669;
  assign n1671 = ~n1613 & ~n1615;
  assign n1672 = pi09 & ~n1671;
  assign n1673 = ~n1430 & n1672;
  assign n1674 = ~n1416 & n1673;
  assign n1675 = ~n1670 & ~n1674;
  assign n1676 = ~n1660 & n1675;
  assign n1677 = ~n1608 & ~n1609;
  assign n1678 = pi09 & ~n1677;
  assign n1679 = po12 & n1678;
  assign n1680 = pi11 & ~n1267;
  assign n1681 = ~pi11 & ~n1251;
  assign n1682 = ~n1241 & n1681;
  assign n1683 = n1266 & ~n1682;
  assign n1684 = ~n1680 & n1683;
  assign n1685 = ~n1608 & n1684;
  assign n1686 = n1266 & ~n1608;
  assign n1687 = ~n1680 & ~n1682;
  assign n1688 = ~n1686 & ~n1687;
  assign n1689 = ~n1685 & ~n1688;
  assign n1690 = po12 & n1689;
  assign n1691 = ~n1679 & ~n1690;
  assign n1692 = n1676 & n1691;
  assign n1693 = ~n1650 & n1692;
  assign n1694 = ~n1626 & n1693;
  assign n1695 = ~pi15 & ~n1467;
  assign n1696 = ~n1479 & n1695;
  assign n1697 = ~n1430 & n1665;
  assign n1698 = ~n1416 & n1697;
  assign n1699 = po12 & n1645;
  assign n1700 = ~n1698 & ~n1699;
  assign n1701 = ~n1696 & n1700;
  assign n1702 = ~n1520 & n1701;
  assign n1703 = n1267 & ~n1686;
  assign n1704 = n1266 & ~n1267;
  assign n1705 = ~n1608 & n1704;
  assign n1706 = ~n1703 & ~n1705;
  assign n1707 = po12 & ~n1706;
  assign n1708 = ~n1430 & ~n1656;
  assign n1709 = ~n1416 & n1708;
  assign n1710 = ~pi11 & ~n1670;
  assign n1711 = ~n1709 & n1710;
  assign n1712 = ~n1707 & n1711;
  assign n1713 = ~n1650 & n1712;
  assign n1714 = ~n1528 & ~n1713;
  assign n1715 = n1702 & n1714;
  assign n1716 = ~n1694 & n1715;
  assign n1717 = ~n1530 & ~n1716;
  assign n1718 = n69 & n73;
  assign n1719 = ~n1717 & n1718;
  assign n1720 = n1386 & ~n1430;
  assign n1721 = ~n1416 & n1720;
  assign n1722 = ~n1290 & n1485;
  assign n1723 = n1500 & ~n1722;
  assign n1724 = ~pi19 & ~n1386;
  assign n1725 = pi19 & ~n1137;
  assign n1726 = ~n1384 & n1725;
  assign n1727 = ~n1382 & n1726;
  assign n1728 = ~n1724 & ~n1727;
  assign n1729 = ~n1411 & n1728;
  assign n1730 = po12 & n1729;
  assign n1731 = ~n1723 & n1730;
  assign n1732 = ~n1721 & ~n1731;
  assign n1733 = pi21 & ~pi23;
  assign n1734 = n69 & n1733;
  assign n1735 = ~n1530 & n1734;
  assign n1736 = ~n1716 & n1735;
  assign n1737 = ~n1732 & ~n1736;
  assign n1738 = ~n1719 & n1737;
  assign n1739 = ~pi23 & ~n1738;
  assign n1740 = pi23 & ~n1732;
  assign n1741 = ~n1736 & n1740;
  assign n1742 = ~n1719 & n1741;
  assign n1743 = ~n1739 & ~n1742;
  assign n1744 = n69 & ~n1743;
  assign n1745 = n67 & n98;
  assign n1746 = ~n1732 & n1745;
  assign n1747 = ~n1736 & n1746;
  assign n1748 = ~n1719 & n1747;
  assign n1749 = ~n1744 & ~n1748;
  assign n1750 = n1718 & ~n1721;
  assign n1751 = ~n1731 & n1750;
  assign n1752 = ~n1732 & n1734;
  assign n1753 = ~n1751 & ~n1752;
  assign n1754 = ~n1530 & ~n1753;
  assign n1755 = ~n1716 & n1754;
  assign n1756 = pi01 & ~pi21;
  assign n1757 = n98 & n1756;
  assign n1758 = n67 & n1757;
  assign n1759 = ~n1732 & n1758;
  assign n1760 = ~pi10 & ~n1759;
  assign n1761 = pi10 & ~pi23;
  assign n1762 = n1756 & n1761;
  assign n1763 = n69 & n1762;
  assign n1764 = ~n1732 & n1763;
  assign n1765 = ~n1760 & ~n1764;
  assign n1766 = pi01 & ~pi08;
  assign n1767 = ~pi03 & ~n1766;
  assign n1768 = ~n1765 & ~n1767;
  assign n1769 = ~n1755 & n1768;
  assign n1770 = pi03 & ~n1766;
  assign n1771 = ~n1764 & ~n1770;
  assign n1772 = ~n1760 & n1771;
  assign n1773 = ~n1755 & n1772;
  assign n1774 = ~pi01 & pi10;
  assign n1775 = ~n1548 & ~n1774;
  assign n1776 = ~n1770 & ~n1775;
  assign n1777 = ~n1753 & n1776;
  assign n1778 = ~n1530 & n1777;
  assign n1779 = ~n1716 & n1778;
  assign n1780 = ~n1767 & n1775;
  assign n1781 = ~n1753 & n1780;
  assign n1782 = ~n1530 & n1781;
  assign n1783 = ~n1716 & n1782;
  assign n1784 = ~n1779 & ~n1783;
  assign n1785 = ~n1773 & n1784;
  assign n1786 = ~n1769 & n1785;
  assign n1787 = ~pi12 & ~n1430;
  assign n1788 = ~n1416 & n1787;
  assign n1789 = pi01 & ~n1430;
  assign n1790 = ~n1416 & n1789;
  assign n1791 = ~n1161 & ~n1573;
  assign n1792 = ~n1790 & n1791;
  assign n1793 = ~n1788 & ~n1792;
  assign n1794 = ~pi03 & ~n1548;
  assign n1795 = ~n1570 & ~n1794;
  assign n1796 = ~n1793 & ~n1795;
  assign n1797 = ~n1788 & n1795;
  assign n1798 = ~n1792 & n1797;
  assign n1799 = ~pi05 & ~n1798;
  assign n1800 = ~n1796 & n1799;
  assign n1801 = ~n1753 & n1800;
  assign n1802 = ~n1530 & n1801;
  assign n1803 = ~n1716 & n1802;
  assign n1804 = ~pi03 & ~n1775;
  assign n1805 = ~n1753 & n1804;
  assign n1806 = ~n1530 & n1805;
  assign n1807 = ~n1716 & n1806;
  assign n1808 = ~pi05 & ~pi21;
  assign n1809 = n98 & n1808;
  assign n1810 = n67 & n1809;
  assign n1811 = ~n1798 & n1810;
  assign n1812 = ~n1732 & n1811;
  assign n1813 = ~n1796 & n1812;
  assign n1814 = ~n1807 & ~n1813;
  assign n1815 = ~n1803 & n1814;
  assign n1816 = ~pi03 & ~n1764;
  assign n1817 = ~n1760 & n1816;
  assign n1818 = ~n1755 & n1817;
  assign n1819 = n1718 & ~n1732;
  assign n1820 = ~pi05 & ~n1788;
  assign n1821 = ~n1792 & n1820;
  assign n1822 = ~n1819 & n1821;
  assign n1823 = ~n1755 & n1822;
  assign n1824 = ~n1818 & ~n1823;
  assign n1825 = n1815 & n1824;
  assign n1826 = ~n1786 & n1825;
  assign n1827 = ~n1793 & ~n1819;
  assign n1828 = ~n1755 & n1827;
  assign po10 = n1755 | n1819;
  assign n1830 = ~pi03 & ~n1788;
  assign n1831 = ~n1792 & n1830;
  assign n1832 = pi03 & ~n1793;
  assign n1833 = ~n1831 & ~n1832;
  assign n1834 = ~n1548 & ~n1833;
  assign n1835 = n1548 & ~n1831;
  assign n1836 = ~n1832 & n1835;
  assign n1837 = ~n1834 & ~n1836;
  assign n1838 = po10 & n1837;
  assign n1839 = ~n1828 & ~n1838;
  assign n1840 = pi05 & ~n1839;
  assign n1841 = ~n1550 & ~n1588;
  assign n1842 = ~n1579 & n1841;
  assign n1843 = ~n1547 & ~n1585;
  assign n1844 = ~n1842 & ~n1843;
  assign n1845 = ~n1585 & ~n1588;
  assign n1846 = ~n1550 & n1845;
  assign n1847 = ~n1547 & n1846;
  assign n1848 = ~n1579 & n1847;
  assign n1849 = ~pi07 & ~n1848;
  assign n1850 = ~n1844 & n1849;
  assign n1851 = ~n1844 & ~n1848;
  assign n1852 = pi07 & ~n1851;
  assign n1853 = ~n1850 & ~n1852;
  assign n1854 = po10 & ~n1853;
  assign n1855 = n1602 & ~n1848;
  assign n1856 = n1603 & ~n1855;
  assign n1857 = n1602 & ~n1603;
  assign n1858 = ~n1848 & n1857;
  assign n1859 = ~pi09 & ~n1858;
  assign n1860 = ~n1856 & n1859;
  assign n1861 = ~n1856 & ~n1858;
  assign n1862 = pi09 & ~n1861;
  assign n1863 = ~n1860 & ~n1862;
  assign n1864 = po10 & ~n1863;
  assign n1865 = po12 & n1559;
  assign n1866 = ~n1148 & ~n1430;
  assign n1867 = ~n1416 & n1866;
  assign n1868 = ~pi09 & ~n1867;
  assign n1869 = ~n1865 & n1868;
  assign n1870 = ~n1865 & ~n1867;
  assign n1871 = pi09 & ~n1870;
  assign n1872 = ~n1869 & ~n1871;
  assign n1873 = ~n1819 & ~n1872;
  assign n1874 = ~n1755 & n1873;
  assign n1875 = po12 & n1542;
  assign n1876 = ~n1430 & ~n1540;
  assign n1877 = ~n1416 & n1876;
  assign n1878 = ~pi07 & ~n1877;
  assign n1879 = ~n1875 & n1878;
  assign n1880 = ~n1875 & ~n1877;
  assign n1881 = pi07 & ~n1880;
  assign n1882 = ~n1879 & ~n1881;
  assign n1883 = ~n1819 & ~n1882;
  assign n1884 = ~n1755 & n1883;
  assign n1885 = ~n1874 & ~n1884;
  assign n1886 = ~n1864 & n1885;
  assign n1887 = ~n1854 & n1886;
  assign n1888 = ~n1840 & n1887;
  assign n1889 = ~n1826 & n1888;
  assign n1890 = ~n1819 & n1879;
  assign n1891 = ~n1755 & n1890;
  assign n1892 = po10 & n1850;
  assign n1893 = ~n1891 & ~n1892;
  assign n1894 = ~n1864 & ~n1874;
  assign n1895 = ~n1893 & n1894;
  assign n1896 = ~n1619 & ~n1674;
  assign n1897 = ~n1612 & n1896;
  assign n1898 = ~n1679 & n1897;
  assign n1899 = ~n1605 & ~n1621;
  assign n1900 = ~n1604 & n1899;
  assign n1901 = ~n1898 & n1900;
  assign n1902 = ~n1598 & n1901;
  assign n1903 = ~n1598 & n1900;
  assign n1904 = n1898 & ~n1903;
  assign n1905 = ~n1902 & ~n1904;
  assign n1906 = po10 & ~n1905;
  assign n1907 = ~n1430 & ~n1671;
  assign n1908 = ~n1416 & n1907;
  assign n1909 = po12 & ~n1677;
  assign n1910 = ~n1908 & ~n1909;
  assign n1911 = ~n1819 & ~n1910;
  assign n1912 = ~n1755 & n1911;
  assign n1913 = ~pi11 & ~n1912;
  assign n1914 = ~n1906 & n1913;
  assign n1915 = ~n1819 & n1869;
  assign n1916 = ~n1755 & n1915;
  assign n1917 = po10 & n1860;
  assign n1918 = ~n1916 & ~n1917;
  assign n1919 = ~n1914 & n1918;
  assign n1920 = ~n1895 & n1919;
  assign n1921 = ~n1889 & n1920;
  assign n1922 = ~n1460 & n1701;
  assign n1923 = ~n1713 & n1922;
  assign n1924 = ~n1694 & n1923;
  assign n1925 = ~n1458 & ~n1698;
  assign n1926 = ~n1448 & n1925;
  assign n1927 = ~n1699 & n1926;
  assign n1928 = ~n1433 & ~n1696;
  assign n1929 = n1927 & n1928;
  assign n1930 = ~n1713 & n1929;
  assign n1931 = pi15 & ~n1458;
  assign n1932 = ~n1448 & n1931;
  assign n1933 = ~n1433 & n1932;
  assign n1934 = ~n1480 & n1933;
  assign n1935 = ~n1482 & ~n1934;
  assign n1936 = ~n1930 & n1935;
  assign n1937 = ~n1458 & ~n1670;
  assign n1938 = ~n1660 & ~n1674;
  assign n1939 = n1937 & n1938;
  assign n1940 = ~n1433 & n1939;
  assign n1941 = ~n1650 & n1940;
  assign n1942 = ~n1448 & ~n1679;
  assign n1943 = ~n1690 & n1942;
  assign n1944 = ~n1481 & n1943;
  assign n1945 = n1941 & n1944;
  assign n1946 = ~n1626 & n1945;
  assign n1947 = ~n1936 & ~n1946;
  assign n1948 = ~n1924 & n1947;
  assign n1949 = ~pi19 & ~n1948;
  assign n1950 = pi19 & ~n1936;
  assign n1951 = ~n1946 & n1950;
  assign n1952 = ~n1924 & n1951;
  assign n1953 = ~n1949 & ~n1952;
  assign n1954 = po10 & ~n1953;
  assign n1955 = ~pi13 & ~n1709;
  assign n1956 = ~n1707 & n1955;
  assign n1957 = ~n1707 & ~n1709;
  assign n1958 = pi13 & ~n1957;
  assign n1959 = ~n1956 & ~n1958;
  assign n1960 = ~n1819 & ~n1959;
  assign n1961 = ~n1755 & n1960;
  assign n1962 = ~pi19 & ~n1525;
  assign n1963 = ~n1526 & n1962;
  assign n1964 = pi19 & ~n1527;
  assign n1965 = ~n1963 & ~n1964;
  assign n1966 = ~n1819 & ~n1965;
  assign n1967 = ~n1755 & n1966;
  assign n1968 = po12 & ~n1647;
  assign n1969 = ~n1430 & ~n1666;
  assign n1970 = ~n1416 & n1969;
  assign n1971 = ~pi15 & ~n1970;
  assign n1972 = ~n1968 & n1971;
  assign n1973 = ~n1968 & ~n1970;
  assign n1974 = pi15 & ~n1973;
  assign n1975 = ~n1972 & ~n1974;
  assign n1976 = ~n1819 & ~n1975;
  assign n1977 = ~n1755 & n1976;
  assign n1978 = ~n1967 & ~n1977;
  assign n1979 = ~n1961 & n1978;
  assign n1980 = ~n1954 & n1979;
  assign n1981 = ~pi11 & ~n1709;
  assign n1982 = ~n1707 & n1981;
  assign n1983 = n1624 & ~n1982;
  assign n1984 = ~n1650 & ~n1670;
  assign n1985 = ~n1604 & ~n1984;
  assign n1986 = n1983 & n1985;
  assign n1987 = ~n1598 & n1986;
  assign n1988 = ~n1679 & n1938;
  assign n1989 = ~n1690 & n1988;
  assign n1990 = ~n1982 & ~n1989;
  assign n1991 = ~n1984 & n1990;
  assign n1992 = ~pi15 & ~n1713;
  assign n1993 = ~n1991 & n1992;
  assign n1994 = ~n1694 & n1993;
  assign n1995 = ~n1987 & n1994;
  assign n1996 = ~n1713 & ~n1991;
  assign n1997 = ~n1694 & n1996;
  assign n1998 = ~n1987 & n1997;
  assign n1999 = pi15 & ~n1998;
  assign n2000 = ~n1995 & ~n1999;
  assign n2001 = po10 & ~n2000;
  assign n2002 = ~n1660 & ~n1690;
  assign n2003 = ~n1674 & ~n1679;
  assign n2004 = ~n1626 & n2003;
  assign n2005 = ~n2002 & ~n2004;
  assign n2006 = ~n1626 & n1989;
  assign n2007 = ~pi13 & ~n2006;
  assign n2008 = ~n2005 & n2007;
  assign n2009 = ~n2005 & ~n2006;
  assign n2010 = pi13 & ~n2009;
  assign n2011 = ~n2008 & ~n2010;
  assign n2012 = po10 & ~n2011;
  assign n2013 = ~n2001 & ~n2012;
  assign n2014 = n1980 & n2013;
  assign n2015 = ~n1906 & ~n1912;
  assign n2016 = pi11 & ~n2015;
  assign n2017 = ~n1481 & n1693;
  assign n2018 = ~n1626 & n2017;
  assign n2019 = n1701 & ~n1713;
  assign n2020 = ~n1481 & ~n2019;
  assign n2021 = ~n2018 & ~n2020;
  assign n2022 = ~pi17 & ~n1525;
  assign n2023 = ~n1526 & n2022;
  assign n2024 = n1460 & ~n2023;
  assign n2025 = ~n1516 & n2024;
  assign n2026 = n1516 & ~n2024;
  assign n2027 = ~n2025 & ~n2026;
  assign n2028 = ~n2021 & n2027;
  assign n2029 = ~n1516 & n2023;
  assign n2030 = ~n1514 & ~n2023;
  assign n2031 = ~n1515 & n2030;
  assign n2032 = ~n2029 & ~n2031;
  assign n2033 = n2021 & ~n2032;
  assign n2034 = ~n2028 & ~n2033;
  assign n2035 = pi21 & po10;
  assign n2036 = ~n2034 & n2035;
  assign n2037 = ~pi21 & ~n1519;
  assign n2038 = pi21 & ~n1504;
  assign n2039 = ~n1518 & n2038;
  assign n2040 = ~n1819 & ~n2039;
  assign n2041 = ~n2037 & n2040;
  assign n2042 = ~n1755 & n2041;
  assign n2043 = ~n1530 & n1751;
  assign n2044 = ~n1716 & n2043;
  assign n2045 = ~n1819 & ~n2044;
  assign n2046 = n2034 & ~n2045;
  assign n2047 = ~n2042 & ~n2046;
  assign n2048 = ~n2036 & n2047;
  assign n2049 = ~n1481 & n1701;
  assign n2050 = ~n1713 & n2049;
  assign n2051 = ~n1694 & n2050;
  assign n2052 = n1700 & ~n1713;
  assign n2053 = ~n1694 & n2052;
  assign n2054 = ~n1481 & ~n1696;
  assign n2055 = ~n2053 & ~n2054;
  assign n2056 = ~n2051 & ~n2055;
  assign n2057 = po10 & n2056;
  assign n2058 = ~n1480 & ~n1819;
  assign n2059 = ~n1755 & n2058;
  assign n2060 = ~n2057 & ~n2059;
  assign n2061 = pi17 & ~n2060;
  assign n2062 = ~n2048 & ~n2061;
  assign n2063 = ~n2016 & n2062;
  assign n2064 = n2014 & n2063;
  assign n2065 = ~n1921 & n2064;
  assign n2066 = po10 & ~n2009;
  assign n2067 = ~n1819 & ~n1957;
  assign n2068 = ~n1755 & n2067;
  assign n2069 = ~pi13 & ~n1977;
  assign n2070 = ~n2068 & n2069;
  assign n2071 = ~n2066 & n2070;
  assign n2072 = ~n2001 & n2071;
  assign n2073 = po10 & ~n1998;
  assign n2074 = ~n1819 & ~n1973;
  assign n2075 = ~n1755 & n2074;
  assign n2076 = ~pi15 & ~n2075;
  assign n2077 = ~n2073 & n2076;
  assign n2078 = ~pi17 & ~n2059;
  assign n2079 = ~n2057 & n2078;
  assign n2080 = ~n2077 & ~n2079;
  assign n2081 = ~n2072 & n2080;
  assign n2082 = ~n1954 & ~n1967;
  assign n2083 = ~n2048 & n2082;
  assign n2084 = ~n2061 & n2083;
  assign n2085 = ~n2081 & n2084;
  assign n2086 = po10 & n1948;
  assign n2087 = ~n1527 & ~n1819;
  assign n2088 = ~n1755 & n2087;
  assign n2089 = ~pi19 & ~n2088;
  assign n2090 = ~n2086 & n2089;
  assign n2091 = ~n2048 & n2090;
  assign n2092 = po10 & n2034;
  assign n2093 = n1519 & ~n1819;
  assign n2094 = ~n1755 & n2093;
  assign n2095 = ~pi21 & ~n2094;
  assign n2096 = ~n2092 & n2095;
  assign n2097 = ~n1748 & ~n2096;
  assign n2098 = ~n2091 & n2097;
  assign n2099 = ~n2085 & n2098;
  assign n2100 = ~n2065 & n2099;
  assign po08 = ~n1749 & ~n2100;
  assign n2102 = ~n1755 & ~n1765;
  assign n2103 = ~n1753 & n1775;
  assign n2104 = ~n1530 & n2103;
  assign n2105 = ~n1716 & n2104;
  assign n2106 = ~pi05 & ~n2105;
  assign n2107 = ~n2102 & n2106;
  assign n2108 = ~po08 & n2107;
  assign n2109 = ~n2091 & ~n2096;
  assign n2110 = ~n2085 & n2109;
  assign n2111 = ~n2065 & n2110;
  assign n2112 = ~pi01 & pi08;
  assign n2113 = ~n1766 & ~n2112;
  assign n2114 = n69 & ~n2113;
  assign n2115 = ~n1743 & n2114;
  assign n2116 = ~n2111 & n2115;
  assign n2117 = pi01 & ~pi23;
  assign n2118 = n69 & n2117;
  assign n2119 = ~n1732 & n2118;
  assign n2120 = ~n1736 & n2119;
  assign n2121 = ~n1719 & n2120;
  assign n2122 = pi08 & ~n2121;
  assign n2123 = n98 & n1766;
  assign n2124 = n67 & n2123;
  assign n2125 = ~n1732 & n2124;
  assign n2126 = ~n1736 & n2125;
  assign n2127 = ~n1719 & n2126;
  assign n2128 = ~n2122 & ~n2127;
  assign n2129 = ~n2096 & ~n2128;
  assign n2130 = ~n2091 & n2129;
  assign n2131 = ~n2085 & n2130;
  assign n2132 = ~n2065 & n2131;
  assign n2133 = ~n1744 & ~n2128;
  assign n2134 = pi01 & ~pi06;
  assign n2135 = ~pi03 & ~n2134;
  assign n2136 = ~n2133 & n2135;
  assign n2137 = ~n2132 & n2136;
  assign n2138 = ~n2116 & n2137;
  assign n2139 = ~pi08 & n77;
  assign n2140 = ~n1770 & ~n2139;
  assign n2141 = ~n2105 & n2140;
  assign n2142 = ~n2102 & n2141;
  assign n2143 = ~n2102 & ~n2105;
  assign n2144 = ~n2140 & ~n2143;
  assign n2145 = ~n2142 & ~n2144;
  assign n2146 = ~pi05 & ~n2145;
  assign n2147 = ~n1749 & n2146;
  assign n2148 = ~n2100 & n2147;
  assign n2149 = ~n2138 & ~n2148;
  assign n2150 = ~n2108 & n2149;
  assign n2151 = ~n2132 & ~n2133;
  assign n2152 = ~n2116 & n2151;
  assign n2153 = pi03 & ~n2134;
  assign n2154 = ~n2152 & n2153;
  assign n2155 = ~pi03 & ~n2152;
  assign n2156 = ~n2154 & ~n2155;
  assign n2157 = n2150 & n2156;
  assign n2158 = po10 & ~n1851;
  assign n2159 = ~n1819 & ~n1880;
  assign n2160 = ~n1755 & n2159;
  assign n2161 = ~pi09 & ~n2160;
  assign n2162 = ~n2158 & n2161;
  assign n2163 = ~n2158 & ~n2160;
  assign n2164 = pi09 & ~n2163;
  assign n2165 = ~n2162 & ~n2164;
  assign n2166 = ~po08 & ~n2165;
  assign n2167 = pi05 & ~n2142;
  assign n2168 = ~n2144 & n2167;
  assign n2169 = ~n1749 & n2168;
  assign n2170 = ~n2100 & n2169;
  assign n2171 = ~n2166 & ~n2170;
  assign n2172 = ~n1854 & ~n1884;
  assign n2173 = ~n1826 & ~n1840;
  assign n2174 = ~n2172 & ~n2173;
  assign n2175 = ~n1840 & n2172;
  assign n2176 = ~n1826 & n2175;
  assign n2177 = ~pi09 & ~n2176;
  assign n2178 = ~n2174 & n2177;
  assign n2179 = ~n2174 & ~n2176;
  assign n2180 = pi09 & ~n2179;
  assign n2181 = ~n2178 & ~n2180;
  assign n2182 = po08 & ~n2181;
  assign n2183 = ~pi07 & ~n1828;
  assign n2184 = ~n1838 & n2183;
  assign n2185 = pi07 & ~n1839;
  assign n2186 = ~n2184 & ~n2185;
  assign n2187 = ~po08 & ~n2186;
  assign n2188 = ~n2182 & ~n2187;
  assign n2189 = ~pi05 & ~n1828;
  assign n2190 = ~n1838 & n2189;
  assign n2191 = ~n1840 & ~n2190;
  assign n2192 = ~n1807 & ~n1818;
  assign n2193 = ~n1786 & n2192;
  assign n2194 = n2191 & ~n2193;
  assign n2195 = ~n2191 & n2193;
  assign n2196 = ~pi07 & ~n2195;
  assign n2197 = ~n2194 & n2196;
  assign n2198 = ~n2194 & ~n2195;
  assign n2199 = pi07 & ~n2198;
  assign n2200 = ~n2197 & ~n2199;
  assign n2201 = po08 & ~n2200;
  assign n2202 = pi05 & ~n2143;
  assign n2203 = ~po08 & n2202;
  assign n2204 = ~n2201 & ~n2203;
  assign n2205 = n2188 & n2204;
  assign n2206 = n2171 & n2205;
  assign n2207 = ~n2157 & n2206;
  assign n2208 = po10 & ~n1861;
  assign n2209 = ~n1819 & ~n1870;
  assign n2210 = ~n1755 & n2209;
  assign n2211 = ~pi11 & ~n2210;
  assign n2212 = ~n2208 & n2211;
  assign n2213 = ~po08 & n2212;
  assign n2214 = ~n1961 & ~n2012;
  assign n2215 = ~n2016 & n2214;
  assign n2216 = ~n1977 & ~n2001;
  assign n2217 = n2215 & ~n2216;
  assign n2218 = ~n1921 & n2217;
  assign n2219 = ~n1916 & ~n1977;
  assign n2220 = ~n1917 & n2219;
  assign n2221 = ~n1914 & n2220;
  assign n2222 = ~pi13 & ~n2068;
  assign n2223 = ~n2066 & n2222;
  assign n2224 = ~n2001 & ~n2223;
  assign n2225 = n2221 & n2224;
  assign n2226 = ~n1895 & n2225;
  assign n2227 = ~n1889 & n2226;
  assign n2228 = n2216 & ~n2223;
  assign n2229 = ~n2215 & n2228;
  assign n2230 = ~n2216 & n2223;
  assign n2231 = ~n2229 & ~n2230;
  assign n2232 = ~n2227 & n2231;
  assign n2233 = ~n2218 & n2232;
  assign n2234 = ~pi17 & ~n1749;
  assign n2235 = ~n2100 & n2234;
  assign n2236 = ~n2233 & n2235;
  assign n2237 = ~po08 & n2162;
  assign n2238 = ~n2236 & ~n2237;
  assign n2239 = ~n2213 & n2238;
  assign n2240 = ~pi15 & ~n2068;
  assign n2241 = ~n2066 & n2240;
  assign n2242 = ~po08 & n2241;
  assign n2243 = ~n1749 & ~n2174;
  assign n2244 = n2177 & n2243;
  assign n2245 = ~n2100 & n2244;
  assign n2246 = n1893 & ~n2176;
  assign n2247 = n1894 & ~n2246;
  assign n2248 = n1893 & ~n1894;
  assign n2249 = ~n2176 & n2248;
  assign n2250 = ~pi11 & ~n1749;
  assign n2251 = ~n2249 & n2250;
  assign n2252 = ~n2247 & n2251;
  assign n2253 = ~n2100 & n2252;
  assign n2254 = ~n2245 & ~n2253;
  assign n2255 = ~n2242 & n2254;
  assign n2256 = ~n1826 & ~n2016;
  assign n2257 = n1888 & n2256;
  assign n2258 = ~n1920 & ~n2016;
  assign n2259 = ~n2214 & ~n2258;
  assign n2260 = ~n2257 & n2259;
  assign n2261 = ~n2257 & ~n2258;
  assign n2262 = n2214 & ~n2261;
  assign n2263 = ~pi15 & ~n1749;
  assign n2264 = ~n2262 & n2263;
  assign n2265 = ~n2260 & n2264;
  assign n2266 = ~n2100 & n2265;
  assign n2267 = ~pi17 & ~n2075;
  assign n2268 = ~n2073 & n2267;
  assign n2269 = ~po08 & n2268;
  assign n2270 = ~n2266 & ~n2269;
  assign n2271 = n2255 & n2270;
  assign n2272 = n2239 & n2271;
  assign n2273 = ~pi13 & ~n1912;
  assign n2274 = ~n1906 & n2273;
  assign n2275 = ~po08 & n2274;
  assign n2276 = ~n1914 & ~n2016;
  assign n2277 = ~n1895 & n1918;
  assign n2278 = ~n1889 & n2277;
  assign n2279 = n2276 & ~n2278;
  assign n2280 = ~n2276 & n2277;
  assign n2281 = ~n1889 & n2280;
  assign n2282 = ~pi13 & ~n1749;
  assign n2283 = ~n2281 & n2282;
  assign n2284 = ~n2279 & n2283;
  assign n2285 = ~n2100 & n2284;
  assign n2286 = ~n2275 & ~n2285;
  assign n2287 = ~n2066 & ~n2068;
  assign n2288 = pi15 & ~n2287;
  assign n2289 = ~n2241 & ~n2288;
  assign n2290 = ~po08 & ~n2289;
  assign n2291 = ~pi15 & ~n1961;
  assign n2292 = ~n2012 & n2291;
  assign n2293 = pi15 & ~n2214;
  assign n2294 = ~n2292 & ~n2293;
  assign n2295 = ~n2258 & n2294;
  assign n2296 = ~n2257 & n2295;
  assign n2297 = ~n2261 & ~n2294;
  assign n2298 = ~n1749 & ~n2297;
  assign n2299 = ~n2296 & n2298;
  assign n2300 = ~n2100 & n2299;
  assign n2301 = ~n2290 & ~n2300;
  assign n2302 = ~n2286 & n2301;
  assign n2303 = ~po08 & n2184;
  assign n2304 = ~n1749 & ~n2194;
  assign n2305 = n2196 & n2304;
  assign n2306 = ~n2100 & n2305;
  assign n2307 = ~n2303 & ~n2306;
  assign n2308 = ~n2166 & ~n2182;
  assign n2309 = ~n2307 & n2308;
  assign n2310 = ~n2302 & ~n2309;
  assign n2311 = n2272 & n2310;
  assign n2312 = ~n2207 & n2311;
  assign n2313 = ~n2247 & ~n2249;
  assign n2314 = pi11 & ~n1749;
  assign n2315 = ~n2100 & n2314;
  assign n2316 = ~n2313 & n2315;
  assign n2317 = ~n2208 & ~n2210;
  assign n2318 = pi11 & ~n2317;
  assign n2319 = ~po08 & n2318;
  assign n2320 = ~n2300 & ~n2319;
  assign n2321 = ~n2316 & n2320;
  assign n2322 = ~pi13 & ~n2281;
  assign n2323 = ~n2279 & n2322;
  assign n2324 = ~n2279 & ~n2281;
  assign n2325 = pi13 & ~n2324;
  assign n2326 = ~n2323 & ~n2325;
  assign n2327 = po08 & ~n2326;
  assign n2328 = pi13 & ~n2015;
  assign n2329 = ~n2274 & ~n2328;
  assign n2330 = ~po08 & ~n2329;
  assign n2331 = ~n2290 & ~n2330;
  assign n2332 = ~n2327 & n2331;
  assign n2333 = n2321 & n2332;
  assign n2334 = ~n2242 & ~n2266;
  assign n2335 = ~n2236 & ~n2269;
  assign n2336 = n2334 & n2335;
  assign n2337 = ~n2302 & n2336;
  assign n2338 = ~n2333 & n2337;
  assign n2339 = ~n2060 & ~po08;
  assign n2340 = ~n1961 & ~n1977;
  assign n2341 = ~n2001 & n2340;
  assign n2342 = ~n2012 & n2341;
  assign n2343 = ~n2016 & n2342;
  assign n2344 = ~n1921 & n2343;
  assign n2345 = ~n2072 & ~n2077;
  assign n2346 = ~n2061 & ~n2079;
  assign n2347 = n2345 & ~n2346;
  assign n2348 = ~n2344 & n2347;
  assign n2349 = ~n2016 & ~n2061;
  assign n2350 = ~n2012 & ~n2079;
  assign n2351 = n2341 & n2350;
  assign n2352 = n2349 & n2351;
  assign n2353 = ~n1921 & n2352;
  assign n2354 = ~n2345 & n2346;
  assign n2355 = ~n2353 & ~n2354;
  assign n2356 = ~n2348 & n2355;
  assign n2357 = po08 & ~n2356;
  assign n2358 = ~n2339 & ~n2357;
  assign n2359 = pi19 & ~n2358;
  assign n2360 = ~pi19 & ~n2339;
  assign n2361 = ~n2357 & n2360;
  assign n2362 = n2342 & n2349;
  assign n2363 = ~n1921 & n2362;
  assign n2364 = ~n2061 & ~n2081;
  assign n2365 = n2082 & ~n2364;
  assign n2366 = ~n2363 & n2365;
  assign n2367 = ~n2082 & n2349;
  assign n2368 = n2342 & n2367;
  assign n2369 = ~n1921 & n2368;
  assign n2370 = ~n2061 & ~n2082;
  assign n2371 = ~n2081 & n2370;
  assign n2372 = pi21 & ~n1749;
  assign n2373 = ~n2371 & n2372;
  assign n2374 = ~n2369 & n2373;
  assign n2375 = ~n2100 & n2374;
  assign n2376 = ~n2366 & n2375;
  assign n2377 = ~n2073 & ~n2075;
  assign n2378 = pi17 & ~n2377;
  assign n2379 = ~po08 & n2378;
  assign n2380 = pi17 & ~n2230;
  assign n2381 = ~n1749 & n2380;
  assign n2382 = ~n2229 & n2381;
  assign n2383 = ~n2227 & n2382;
  assign n2384 = ~n2218 & n2383;
  assign n2385 = ~n2100 & n2384;
  assign n2386 = ~n2379 & ~n2385;
  assign n2387 = ~n2376 & n2386;
  assign n2388 = ~n2361 & n2387;
  assign n2389 = ~n2359 & n2388;
  assign n2390 = n1743 & ~n1749;
  assign n2391 = ~n2100 & n2390;
  assign n2392 = ~n2111 & n2391;
  assign n2393 = n1738 & ~po08;
  assign n2394 = ~pi25 & ~n2393;
  assign n2395 = ~n2392 & n2394;
  assign n2396 = ~n2392 & ~n2393;
  assign n2397 = pi25 & ~n2396;
  assign n2398 = ~n2395 & ~n2397;
  assign n2399 = ~n2363 & ~n2364;
  assign n2400 = ~n2082 & ~n2090;
  assign n2401 = ~n2048 & ~n2400;
  assign n2402 = n2048 & n2400;
  assign n2403 = ~n2401 & ~n2402;
  assign n2404 = ~n2399 & n2403;
  assign n2405 = n2048 & ~n2090;
  assign n2406 = ~n2091 & ~n2405;
  assign n2407 = ~n2364 & n2406;
  assign n2408 = ~n2363 & n2407;
  assign n2409 = pi23 & ~n1749;
  assign n2410 = ~n2100 & n2409;
  assign n2411 = ~n2408 & n2410;
  assign n2412 = ~n2404 & n2411;
  assign n2413 = ~n2092 & ~n2094;
  assign n2414 = pi23 & ~n2413;
  assign n2415 = ~po08 & n2414;
  assign n2416 = n67 & ~n2415;
  assign n2417 = ~pi21 & ~n2088;
  assign n2418 = ~n2086 & n2417;
  assign n2419 = ~n2086 & ~n2088;
  assign n2420 = pi21 & ~n2419;
  assign n2421 = ~n2418 & ~n2420;
  assign n2422 = ~po08 & ~n2421;
  assign n2423 = ~n2369 & ~n2371;
  assign n2424 = ~n2366 & n2423;
  assign n2425 = ~pi21 & ~n1749;
  assign n2426 = ~n2100 & n2425;
  assign n2427 = ~n2424 & n2426;
  assign n2428 = ~n2422 & ~n2427;
  assign n2429 = n2416 & n2428;
  assign n2430 = ~n2412 & n2429;
  assign n2431 = ~n2398 & n2430;
  assign n2432 = n2389 & n2431;
  assign n2433 = ~n2338 & n2432;
  assign n2434 = ~n2312 & n2433;
  assign n2435 = ~n2357 & ~n2376;
  assign n2436 = n2428 & n2435;
  assign n2437 = n2360 & n2436;
  assign n2438 = ~po08 & ~n2419;
  assign n2439 = ~n1749 & ~n2371;
  assign n2440 = ~n2369 & n2439;
  assign n2441 = ~n2100 & n2440;
  assign n2442 = ~n2366 & n2441;
  assign n2443 = ~pi21 & ~n2442;
  assign n2444 = ~n2438 & n2443;
  assign n2445 = po08 & ~n2408;
  assign n2446 = ~n2404 & n2445;
  assign n2447 = ~po08 & ~n2413;
  assign n2448 = ~pi23 & ~n2447;
  assign n2449 = ~n2446 & n2448;
  assign n2450 = ~n2444 & ~n2449;
  assign n2451 = ~n2437 & n2450;
  assign n2452 = ~n2412 & n2416;
  assign n2453 = ~n2398 & n2452;
  assign n2454 = ~n2451 & n2453;
  assign n2455 = n69 & ~n2396;
  assign n2456 = ~n2396 & ~n2455;
  assign n2457 = ~n2454 & n2456;
  assign n2458 = ~n2434 & n2457;
  assign n2459 = ~n2454 & ~n2455;
  assign po06 = n2434 | ~n2459;
  assign n2461 = n2387 & n2428;
  assign n2462 = ~n2359 & ~n2361;
  assign n2463 = n2461 & n2462;
  assign n2464 = ~n2338 & n2463;
  assign n2465 = ~n2312 & n2464;
  assign n2466 = n2451 & ~n2465;
  assign n2467 = ~n2412 & ~n2415;
  assign n2468 = ~n2395 & n2467;
  assign n2469 = ~n2397 & n2468;
  assign n2470 = ~n2466 & n2469;
  assign n2471 = po06 & n2470;
  assign n2472 = ~n2458 & ~n2471;
  assign n2473 = n67 & ~n2472;
  assign n2474 = ~pi27 & ~n2458;
  assign n2475 = ~n2471 & n2474;
  assign n2476 = pi27 & ~n2472;
  assign n2477 = ~n2475 & ~n2476;
  assign n2478 = ~n2473 & n2477;
  assign n2479 = n2358 & ~n2455;
  assign n2480 = ~n2454 & n2479;
  assign n2481 = ~n2434 & n2480;
  assign n2482 = ~n2361 & n2386;
  assign n2483 = ~n2359 & n2482;
  assign n2484 = ~n2338 & n2483;
  assign n2485 = ~n2312 & n2484;
  assign n2486 = ~n2338 & n2386;
  assign n2487 = ~n2312 & n2486;
  assign n2488 = ~n2462 & ~n2487;
  assign n2489 = ~n2485 & ~n2488;
  assign n2490 = po06 & n2489;
  assign n2491 = ~n2481 & ~n2490;
  assign n2492 = ~pi21 & ~n2491;
  assign n2493 = pi21 & ~n2481;
  assign n2494 = ~n2490 & n2493;
  assign n2495 = n2335 & n2386;
  assign n2496 = ~n2302 & n2334;
  assign n2497 = ~n2333 & n2496;
  assign n2498 = ~n2237 & ~n2266;
  assign n2499 = ~n2213 & n2498;
  assign n2500 = n2255 & n2499;
  assign n2501 = n2310 & n2500;
  assign n2502 = ~n2207 & n2501;
  assign n2503 = ~n2497 & ~n2502;
  assign n2504 = ~n2495 & ~n2503;
  assign n2505 = n2495 & ~n2497;
  assign n2506 = ~n2502 & n2505;
  assign n2507 = ~n2504 & ~n2506;
  assign n2508 = po06 & ~n2507;
  assign n2509 = ~po08 & ~n2377;
  assign n2510 = ~n1749 & n2231;
  assign n2511 = ~n2227 & n2510;
  assign n2512 = ~n2218 & n2511;
  assign n2513 = ~n2100 & n2512;
  assign n2514 = ~n2509 & ~n2513;
  assign n2515 = ~n2455 & ~n2514;
  assign n2516 = ~n2454 & n2515;
  assign n2517 = ~n2434 & n2516;
  assign n2518 = ~pi19 & ~n2517;
  assign n2519 = ~n2508 & n2518;
  assign n2520 = ~n2494 & n2519;
  assign n2521 = ~n2492 & n2520;
  assign n2522 = ~pi23 & ~n2442;
  assign n2523 = ~n2438 & n2522;
  assign n2524 = ~n2455 & n2523;
  assign n2525 = ~n2454 & n2524;
  assign n2526 = ~n2434 & n2525;
  assign n2527 = ~n2376 & n2428;
  assign n2528 = ~n2361 & ~n2485;
  assign n2529 = n2527 & ~n2528;
  assign n2530 = ~n2361 & ~n2527;
  assign n2531 = ~n2485 & n2530;
  assign n2532 = ~pi23 & ~n2531;
  assign n2533 = po06 & n2532;
  assign n2534 = ~n2529 & n2533;
  assign n2535 = ~n2526 & ~n2534;
  assign n2536 = ~n2492 & n2535;
  assign n2537 = ~n2521 & n2536;
  assign n2538 = po06 & ~n2531;
  assign n2539 = ~n2529 & n2538;
  assign n2540 = ~n2438 & ~n2442;
  assign n2541 = ~n2455 & n2540;
  assign n2542 = ~n2454 & n2541;
  assign n2543 = ~n2434 & n2542;
  assign n2544 = pi23 & ~n2543;
  assign n2545 = ~n2539 & n2544;
  assign n2546 = ~n2437 & ~n2444;
  assign n2547 = ~n2465 & n2546;
  assign n2548 = ~n2446 & ~n2447;
  assign n2549 = pi23 & ~n2548;
  assign n2550 = ~n2449 & ~n2549;
  assign n2551 = ~n2547 & ~n2550;
  assign n2552 = n2451 & ~n2549;
  assign n2553 = ~n2465 & n2552;
  assign n2554 = pi25 & ~n2553;
  assign n2555 = po06 & n2554;
  assign n2556 = ~n2551 & n2555;
  assign n2557 = ~n2551 & ~n2553;
  assign n2558 = ~pi25 & po06;
  assign n2559 = ~n2557 & n2558;
  assign n2560 = ~pi25 & ~n2447;
  assign n2561 = ~n2446 & n2560;
  assign n2562 = pi25 & ~n2548;
  assign n2563 = ~n2561 & ~n2562;
  assign n2564 = ~n2455 & ~n2563;
  assign n2565 = ~n2454 & n2564;
  assign n2566 = ~n2434 & n2565;
  assign n2567 = n65 & ~n2566;
  assign n2568 = ~n2559 & n2567;
  assign n2569 = ~n2556 & n2568;
  assign n2570 = ~n2545 & n2569;
  assign n2571 = ~n2537 & n2570;
  assign n2572 = ~pi25 & ~pi29;
  assign n2573 = ~pi31 & n2572;
  assign n2574 = ~n2447 & n2573;
  assign n2575 = ~n2446 & n2574;
  assign n2576 = ~n2455 & n2575;
  assign n2577 = ~n2454 & n2576;
  assign n2578 = ~n2434 & n2577;
  assign n2579 = po06 & n2573;
  assign n2580 = ~n2557 & n2579;
  assign n2581 = ~n2578 & ~n2580;
  assign n2582 = ~n2473 & n2581;
  assign n2583 = ~n2571 & n2582;
  assign n2584 = ~n2478 & ~n2583;
  assign n2585 = pi03 & ~n2133;
  assign n2586 = ~n2132 & n2585;
  assign n2587 = ~n2116 & n2586;
  assign n2588 = ~n2155 & ~n2587;
  assign n2589 = ~n2134 & ~n2588;
  assign n2590 = n2134 & ~n2587;
  assign n2591 = ~n2155 & n2590;
  assign n2592 = ~n2589 & ~n2591;
  assign n2593 = ~pi05 & ~n2592;
  assign n2594 = po06 & n2593;
  assign n2595 = pi01 & ~pi25;
  assign n2596 = n67 & n2595;
  assign n2597 = ~n2396 & n2596;
  assign n2598 = ~pi06 & ~n2597;
  assign n2599 = pi06 & ~pi27;
  assign n2600 = n65 & n2599;
  assign n2601 = n2595 & n2600;
  assign n2602 = ~n2396 & n2601;
  assign n2603 = ~n2598 & ~n2602;
  assign n2604 = ~n2454 & n2603;
  assign n2605 = ~n2434 & n2604;
  assign n2606 = ~pi01 & pi06;
  assign n2607 = ~n2134 & ~n2606;
  assign n2608 = n67 & ~n2607;
  assign n2609 = ~n2415 & n2608;
  assign n2610 = n2428 & n2609;
  assign n2611 = ~n2412 & n2610;
  assign n2612 = ~n2398 & n2611;
  assign n2613 = n2389 & n2612;
  assign n2614 = ~n2338 & n2613;
  assign n2615 = ~n2312 & n2614;
  assign n2616 = ~n2412 & n2609;
  assign n2617 = ~n2398 & n2616;
  assign n2618 = ~n2451 & n2617;
  assign n2619 = pi01 & ~pi04;
  assign n2620 = ~pi03 & ~n2619;
  assign n2621 = ~n2618 & n2620;
  assign n2622 = ~n2615 & n2621;
  assign n2623 = ~n2605 & n2622;
  assign n2624 = ~pi05 & ~n2152;
  assign n2625 = ~n2455 & n2624;
  assign n2626 = ~n2454 & n2625;
  assign n2627 = ~n2434 & n2626;
  assign n2628 = ~n2623 & ~n2627;
  assign n2629 = ~n2594 & n2628;
  assign n2630 = ~n2615 & ~n2618;
  assign n2631 = ~n2605 & n2630;
  assign n2632 = pi03 & ~n2619;
  assign n2633 = ~n2631 & n2632;
  assign n2634 = ~pi03 & ~n2631;
  assign n2635 = ~n2633 & ~n2634;
  assign n2636 = n2629 & n2635;
  assign n2637 = ~n1839 & ~po08;
  assign n2638 = ~n1749 & ~n2198;
  assign n2639 = ~n2100 & n2638;
  assign n2640 = ~pi09 & ~n2639;
  assign n2641 = ~n2637 & n2640;
  assign n2642 = ~n2637 & ~n2639;
  assign n2643 = pi09 & ~n2642;
  assign n2644 = ~n2641 & ~n2643;
  assign n2645 = ~n2455 & ~n2644;
  assign n2646 = ~n2454 & n2645;
  assign n2647 = ~n2434 & n2646;
  assign n2648 = pi05 & ~n2133;
  assign n2649 = ~n2132 & n2648;
  assign n2650 = ~n2116 & n2649;
  assign n2651 = ~n2455 & n2650;
  assign n2652 = ~n2454 & n2651;
  assign n2653 = ~n2434 & n2652;
  assign n2654 = ~po08 & ~n2143;
  assign n2655 = ~n1749 & n2145;
  assign n2656 = ~n2100 & n2655;
  assign n2657 = ~pi07 & ~n2656;
  assign n2658 = ~n2654 & n2657;
  assign n2659 = ~n2654 & ~n2656;
  assign n2660 = pi07 & ~n2659;
  assign n2661 = ~n2658 & ~n2660;
  assign n2662 = ~n2455 & ~n2661;
  assign n2663 = ~n2454 & n2662;
  assign n2664 = ~n2434 & n2663;
  assign n2665 = ~n2653 & ~n2664;
  assign n2666 = ~n2647 & n2665;
  assign n2667 = ~n2187 & ~n2201;
  assign n2668 = ~n2170 & ~n2203;
  assign n2669 = ~n2157 & n2668;
  assign n2670 = ~n2667 & ~n2669;
  assign n2671 = ~n2170 & ~n2187;
  assign n2672 = n2204 & n2671;
  assign n2673 = ~n2157 & n2672;
  assign n2674 = ~pi09 & ~n2673;
  assign n2675 = ~n2670 & n2674;
  assign n2676 = ~n2670 & ~n2673;
  assign n2677 = pi09 & ~n2676;
  assign n2678 = ~n2675 & ~n2677;
  assign n2679 = po06 & ~n2678;
  assign n2680 = pi05 & ~n2591;
  assign n2681 = ~n2589 & n2680;
  assign n2682 = po06 & n2681;
  assign n2683 = ~pi05 & ~n2659;
  assign n2684 = pi05 & ~n2656;
  assign n2685 = ~n2654 & n2684;
  assign n2686 = ~n2683 & ~n2685;
  assign n2687 = ~n2138 & ~n2154;
  assign n2688 = ~n2155 & n2687;
  assign n2689 = ~n2686 & ~n2688;
  assign n2690 = ~n2155 & ~n2685;
  assign n2691 = n2687 & n2690;
  assign n2692 = ~n2683 & n2691;
  assign n2693 = ~pi07 & ~n2692;
  assign n2694 = ~n2689 & n2693;
  assign n2695 = ~n2689 & ~n2692;
  assign n2696 = pi07 & ~n2695;
  assign n2697 = ~n2694 & ~n2696;
  assign n2698 = po06 & ~n2697;
  assign n2699 = ~n2682 & ~n2698;
  assign n2700 = ~n2679 & n2699;
  assign n2701 = n2666 & n2700;
  assign n2702 = ~n2636 & n2701;
  assign n2703 = po08 & ~n2324;
  assign n2704 = ~n2015 & ~po08;
  assign n2705 = ~pi15 & ~n2704;
  assign n2706 = ~n2703 & n2705;
  assign n2707 = ~n2455 & n2706;
  assign n2708 = ~n2454 & n2707;
  assign n2709 = ~n2434 & n2708;
  assign n2710 = ~n2260 & ~n2262;
  assign n2711 = po08 & ~n2710;
  assign n2712 = ~po08 & ~n2287;
  assign n2713 = ~pi17 & ~n2712;
  assign n2714 = ~n2711 & n2713;
  assign n2715 = ~n2455 & n2714;
  assign n2716 = ~n2454 & n2715;
  assign n2717 = ~n2434 & n2716;
  assign n2718 = ~n2709 & ~n2717;
  assign n2719 = ~n2455 & n2641;
  assign n2720 = ~n2454 & n2719;
  assign n2721 = ~n2434 & n2720;
  assign n2722 = ~po08 & ~n2163;
  assign n2723 = ~n1749 & ~n2179;
  assign n2724 = ~n2100 & n2723;
  assign n2725 = ~pi11 & ~n2724;
  assign n2726 = ~n2722 & n2725;
  assign n2727 = ~n2455 & n2726;
  assign n2728 = ~n2454 & n2727;
  assign n2729 = ~n2434 & n2728;
  assign n2730 = ~n2721 & ~n2729;
  assign n2731 = n2718 & n2730;
  assign n2732 = ~n2237 & n2254;
  assign n2733 = ~n2213 & n2732;
  assign n2734 = ~n2309 & n2733;
  assign n2735 = ~n2207 & n2734;
  assign n2736 = ~n2327 & ~n2330;
  assign n2737 = ~pi15 & ~n2319;
  assign n2738 = ~n2316 & n2737;
  assign n2739 = ~n2736 & n2738;
  assign n2740 = ~n2735 & n2739;
  assign n2741 = ~n2316 & ~n2319;
  assign n2742 = ~n2735 & n2741;
  assign n2743 = ~pi15 & ~n2330;
  assign n2744 = ~n2327 & n2743;
  assign n2745 = ~n2742 & n2744;
  assign n2746 = ~n2740 & ~n2745;
  assign n2747 = po06 & ~n2746;
  assign n2748 = ~n2703 & ~n2704;
  assign n2749 = pi13 & ~n2748;
  assign n2750 = ~n2301 & n2749;
  assign n2751 = n2301 & ~n2749;
  assign n2752 = n2741 & ~n2751;
  assign n2753 = ~n2750 & n2752;
  assign n2754 = ~n2735 & n2753;
  assign n2755 = n2286 & n2301;
  assign n2756 = ~n2286 & ~n2301;
  assign n2757 = ~n2755 & ~n2756;
  assign n2758 = ~n2741 & ~n2757;
  assign n2759 = n2734 & ~n2757;
  assign n2760 = ~n2207 & n2759;
  assign n2761 = ~n2758 & ~n2760;
  assign n2762 = ~n2754 & n2761;
  assign n2763 = ~pi17 & ~n2762;
  assign n2764 = po06 & n2763;
  assign n2765 = ~n2747 & ~n2764;
  assign n2766 = po06 & n2675;
  assign n2767 = n2307 & ~n2673;
  assign n2768 = n2308 & ~n2767;
  assign n2769 = n2307 & ~n2308;
  assign n2770 = ~n2673 & n2769;
  assign n2771 = ~pi11 & ~n2770;
  assign n2772 = ~n2768 & n2771;
  assign n2773 = po06 & n2772;
  assign n2774 = ~n2766 & ~n2773;
  assign n2775 = n2765 & n2774;
  assign n2776 = n2731 & n2775;
  assign n2777 = po08 & ~n2313;
  assign n2778 = ~po08 & ~n2317;
  assign n2779 = ~pi13 & ~n2778;
  assign n2780 = ~n2777 & n2779;
  assign n2781 = ~n2455 & n2780;
  assign n2782 = ~n2454 & n2781;
  assign n2783 = ~n2434 & n2782;
  assign n2784 = ~n2253 & ~n2319;
  assign n2785 = ~n2213 & ~n2316;
  assign n2786 = n2784 & n2785;
  assign n2787 = ~n2237 & ~n2245;
  assign n2788 = ~n2309 & n2787;
  assign n2789 = ~n2207 & n2788;
  assign n2790 = n2786 & ~n2789;
  assign n2791 = ~n2786 & n2788;
  assign n2792 = ~n2207 & n2791;
  assign n2793 = ~pi13 & ~n2792;
  assign n2794 = ~n2790 & n2793;
  assign n2795 = po06 & n2794;
  assign n2796 = ~n2783 & ~n2795;
  assign n2797 = pi15 & ~n2748;
  assign n2798 = ~n2706 & ~n2797;
  assign n2799 = ~n2455 & ~n2798;
  assign n2800 = ~n2454 & n2799;
  assign n2801 = ~n2434 & n2800;
  assign n2802 = ~n2237 & ~n2330;
  assign n2803 = ~n2213 & n2802;
  assign n2804 = pi15 & ~n2245;
  assign n2805 = ~n2253 & n2804;
  assign n2806 = ~n2327 & n2805;
  assign n2807 = n2803 & n2806;
  assign n2808 = ~n2309 & n2807;
  assign n2809 = ~n2207 & n2808;
  assign n2810 = ~pi15 & ~n2245;
  assign n2811 = ~n2253 & n2810;
  assign n2812 = ~n2213 & ~n2237;
  assign n2813 = n2811 & n2812;
  assign n2814 = ~n2309 & n2813;
  assign n2815 = ~n2736 & n2814;
  assign n2816 = ~n2207 & n2815;
  assign n2817 = ~pi15 & ~n2741;
  assign n2818 = ~n2736 & n2817;
  assign n2819 = pi15 & ~n2330;
  assign n2820 = ~n2327 & n2819;
  assign n2821 = ~n2741 & n2820;
  assign n2822 = ~n2818 & ~n2821;
  assign n2823 = ~n2816 & n2822;
  assign n2824 = ~n2809 & n2823;
  assign n2825 = n2741 & n2743;
  assign n2826 = ~n2327 & n2825;
  assign n2827 = ~n2735 & n2826;
  assign n2828 = pi15 & ~n2319;
  assign n2829 = ~n2316 & n2828;
  assign n2830 = ~n2736 & n2829;
  assign n2831 = ~n2735 & n2830;
  assign n2832 = ~n2827 & ~n2831;
  assign n2833 = n2824 & n2832;
  assign n2834 = po06 & n2833;
  assign n2835 = ~n2801 & ~n2834;
  assign n2836 = ~n2796 & n2835;
  assign n2837 = ~n2455 & n2658;
  assign n2838 = ~n2454 & n2837;
  assign n2839 = ~n2434 & n2838;
  assign n2840 = po06 & n2694;
  assign n2841 = ~n2839 & ~n2840;
  assign n2842 = ~n2647 & ~n2679;
  assign n2843 = ~n2841 & n2842;
  assign n2844 = ~n2836 & ~n2843;
  assign n2845 = n2776 & n2844;
  assign n2846 = ~n2702 & n2845;
  assign n2847 = pi17 & ~n2758;
  assign n2848 = ~n2760 & n2847;
  assign n2849 = ~n2754 & n2848;
  assign n2850 = po06 & n2849;
  assign n2851 = ~n2711 & ~n2712;
  assign n2852 = pi17 & ~n2851;
  assign n2853 = ~n2455 & n2852;
  assign n2854 = ~n2454 & n2853;
  assign n2855 = ~n2434 & n2854;
  assign n2856 = n2567 & ~n2855;
  assign n2857 = ~n2850 & n2856;
  assign n2858 = ~n2545 & n2857;
  assign n2859 = ~n2492 & n2858;
  assign n2860 = ~n2508 & ~n2517;
  assign n2861 = ~pi19 & ~n2860;
  assign n2862 = pi19 & ~n2517;
  assign n2863 = ~n2508 & n2862;
  assign n2864 = ~n2861 & ~n2863;
  assign n2865 = ~n2556 & ~n2559;
  assign n2866 = ~n2494 & n2865;
  assign n2867 = ~n2864 & n2866;
  assign n2868 = n2859 & n2867;
  assign n2869 = ~n2790 & ~n2792;
  assign n2870 = pi13 & ~n2869;
  assign n2871 = ~n2794 & ~n2870;
  assign n2872 = po06 & ~n2871;
  assign n2873 = ~n2722 & ~n2724;
  assign n2874 = pi11 & ~n2873;
  assign n2875 = ~n2455 & n2874;
  assign n2876 = ~n2454 & n2875;
  assign n2877 = ~n2434 & n2876;
  assign n2878 = ~n2777 & ~n2778;
  assign n2879 = pi13 & ~n2878;
  assign n2880 = ~n2780 & ~n2879;
  assign n2881 = ~n2455 & ~n2880;
  assign n2882 = ~n2454 & n2881;
  assign n2883 = ~n2434 & n2882;
  assign n2884 = ~n2801 & ~n2883;
  assign n2885 = ~n2877 & n2884;
  assign n2886 = ~n2768 & ~n2770;
  assign n2887 = pi11 & ~n2886;
  assign n2888 = po06 & n2887;
  assign n2889 = ~n2834 & ~n2888;
  assign n2890 = n2885 & n2889;
  assign n2891 = ~n2872 & n2890;
  assign n2892 = n2718 & ~n2747;
  assign n2893 = ~n2764 & n2892;
  assign n2894 = ~n2836 & n2893;
  assign n2895 = ~n2891 & n2894;
  assign n2896 = ~n2478 & ~n2895;
  assign n2897 = n2868 & n2896;
  assign n2898 = ~n2846 & n2897;
  assign n2899 = ~n2472 & ~n2898;
  assign n2900 = ~n2584 & n2899;
  assign n2901 = po06 & n2557;
  assign n2902 = ~n2455 & ~n2548;
  assign n2903 = ~n2454 & n2902;
  assign n2904 = ~n2434 & n2903;
  assign n2905 = ~pi25 & ~n2904;
  assign n2906 = ~n2901 & n2905;
  assign n2907 = ~n2850 & ~n2855;
  assign n2908 = ~n2494 & n2907;
  assign n2909 = ~n2492 & n2908;
  assign n2910 = ~n2864 & n2909;
  assign n2911 = ~n2895 & n2910;
  assign n2912 = ~n2846 & n2911;
  assign n2913 = n2537 & ~n2912;
  assign n2914 = ~n2559 & ~n2566;
  assign n2915 = ~n2556 & n2914;
  assign n2916 = ~n2545 & n2915;
  assign n2917 = ~n2913 & n2916;
  assign n2918 = ~n2906 & ~n2917;
  assign po04 = n2584 | n2898;
  assign n2920 = n2477 & po04;
  assign n2921 = ~n2918 & n2920;
  assign n2922 = ~n2900 & ~n2921;
  assign n2923 = n65 & ~n2922;
  assign n2924 = ~pi23 & ~n2491;
  assign n2925 = ~n2898 & n2924;
  assign n2926 = ~n2584 & n2925;
  assign n2927 = ~n2492 & ~n2494;
  assign n2928 = ~n2864 & n2907;
  assign n2929 = ~n2895 & n2928;
  assign n2930 = ~n2846 & n2929;
  assign n2931 = ~n2519 & ~n2930;
  assign n2932 = n2927 & ~n2931;
  assign n2933 = ~n2519 & ~n2927;
  assign n2934 = ~n2930 & n2933;
  assign n2935 = ~pi23 & ~n2934;
  assign n2936 = po04 & n2935;
  assign n2937 = ~n2932 & n2936;
  assign n2938 = ~n2926 & ~n2937;
  assign n2939 = n2535 & ~n2545;
  assign n2940 = ~n2492 & ~n2521;
  assign n2941 = ~n2939 & n2940;
  assign n2942 = ~n2912 & n2941;
  assign n2943 = ~n2912 & n2940;
  assign n2944 = n2939 & ~n2943;
  assign n2945 = ~n2942 & ~n2944;
  assign n2946 = pi25 & po04;
  assign n2947 = ~n2945 & n2946;
  assign n2948 = ~pi25 & ~n2942;
  assign n2949 = po04 & n2948;
  assign n2950 = ~n2944 & n2949;
  assign n2951 = ~n2539 & ~n2543;
  assign n2952 = ~pi25 & ~n2951;
  assign n2953 = pi25 & ~n2543;
  assign n2954 = ~n2539 & n2953;
  assign n2955 = ~n2952 & ~n2954;
  assign n2956 = ~n2898 & ~n2955;
  assign n2957 = ~n2584 & n2956;
  assign n2958 = ~n2950 & ~n2957;
  assign n2959 = ~n2947 & n2958;
  assign n2960 = ~n2938 & n2959;
  assign n2961 = ~n2545 & ~n2913;
  assign n2962 = ~n2915 & ~n2961;
  assign n2963 = ~pi27 & ~n2917;
  assign n2964 = po04 & n2963;
  assign n2965 = ~n2962 & n2964;
  assign n2966 = po04 & ~n2945;
  assign n2967 = ~n2898 & n2951;
  assign n2968 = ~n2584 & n2967;
  assign n2969 = ~pi25 & ~n2968;
  assign n2970 = ~n2966 & n2969;
  assign n2971 = ~pi27 & ~n2904;
  assign n2972 = ~n2901 & n2971;
  assign n2973 = ~n2898 & n2972;
  assign n2974 = ~n2584 & n2973;
  assign n2975 = ~n2970 & ~n2974;
  assign n2976 = ~n2965 & n2975;
  assign n2977 = ~n2960 & n2976;
  assign n2978 = ~pi29 & ~n2900;
  assign n2979 = ~n2921 & n2978;
  assign n2980 = pi29 & ~n2922;
  assign n2981 = ~n2979 & ~n2980;
  assign n2982 = ~n2917 & po04;
  assign n2983 = ~n2962 & n2982;
  assign n2984 = ~n2901 & ~n2904;
  assign n2985 = ~n2898 & n2984;
  assign n2986 = ~n2584 & n2985;
  assign n2987 = pi27 & ~n2986;
  assign n2988 = ~n2983 & n2987;
  assign n2989 = ~pi31 & ~n2988;
  assign n2990 = ~n2981 & n2989;
  assign n2991 = ~n2977 & n2990;
  assign n2992 = ~n2923 & ~n2991;
  assign n2993 = ~pi00 & pi01;
  assign n2994 = pi02 & n2993;
  assign n2995 = ~pi03 & ~n2994;
  assign n2996 = ~n2992 & n2995;
  assign n2997 = ~pi01 & pi04;
  assign n2998 = ~n2477 & ~n2997;
  assign n2999 = pi01 & ~pi27;
  assign n3000 = n65 & n2999;
  assign n3001 = ~n2472 & n3000;
  assign n3002 = pi04 & ~n3001;
  assign n3003 = ~n2998 & n3002;
  assign n3004 = n2868 & ~n2895;
  assign n3005 = ~n2846 & n3004;
  assign n3006 = pi04 & ~n2578;
  assign n3007 = ~n2580 & n3006;
  assign n3008 = ~n3001 & n3007;
  assign n3009 = ~n2571 & n3008;
  assign n3010 = ~n3005 & n3009;
  assign n3011 = ~n3003 & ~n3010;
  assign n3012 = pi01 & ~pi02;
  assign n3013 = pi03 & n3012;
  assign n3014 = ~n3011 & ~n3013;
  assign n3015 = n67 & n2619;
  assign n3016 = ~n2472 & n3015;
  assign n3017 = pi03 & ~n2578;
  assign n3018 = ~n2580 & n3017;
  assign n3019 = ~n3016 & n3018;
  assign n3020 = ~n2571 & n3019;
  assign n3021 = ~n3005 & n3020;
  assign n3022 = ~n2578 & n3012;
  assign n3023 = ~n2580 & n3022;
  assign n3024 = ~n3016 & n3023;
  assign n3025 = ~n2571 & n3024;
  assign n3026 = ~n3005 & n3025;
  assign n3027 = ~n2478 & n2619;
  assign n3028 = n3012 & ~n3027;
  assign n3029 = n2619 & ~n3012;
  assign n3030 = ~n2478 & n3029;
  assign n3031 = pi03 & ~n3030;
  assign n3032 = ~n3028 & ~n3031;
  assign n3033 = ~n3026 & n3032;
  assign n3034 = ~n3021 & n3033;
  assign n3035 = ~n3014 & ~n3034;
  assign n3036 = po06 & n2592;
  assign n3037 = n2152 & ~n2455;
  assign n3038 = ~n2454 & n3037;
  assign n3039 = ~n2434 & n3038;
  assign n3040 = ~pi07 & ~n3039;
  assign n3041 = ~n3036 & n3040;
  assign n3042 = ~n3036 & ~n3039;
  assign n3043 = pi07 & ~n3042;
  assign n3044 = ~n3041 & ~n3043;
  assign n3045 = ~n2898 & ~n3044;
  assign n3046 = ~n2584 & n3045;
  assign n3047 = ~pi05 & ~n3042;
  assign n3048 = pi05 & ~n3039;
  assign n3049 = ~n3036 & n3048;
  assign n3050 = ~n3047 & ~n3049;
  assign n3051 = ~n2623 & ~n2633;
  assign n3052 = ~n2634 & n3051;
  assign n3053 = ~n3050 & ~n3052;
  assign n3054 = ~n2634 & ~n3049;
  assign n3055 = n3051 & n3054;
  assign n3056 = ~n3047 & n3055;
  assign n3057 = ~pi07 & ~n3056;
  assign n3058 = ~n3053 & n3057;
  assign n3059 = ~n3053 & ~n3056;
  assign n3060 = pi07 & ~n3059;
  assign n3061 = ~n3058 & ~n3060;
  assign n3062 = po04 & ~n3061;
  assign n3063 = ~n3046 & ~n3062;
  assign n3064 = ~pi05 & ~n2631;
  assign n3065 = pi05 & ~n2618;
  assign n3066 = ~n2615 & n3065;
  assign n3067 = ~n2605 & n3066;
  assign n3068 = ~n3064 & ~n3067;
  assign n3069 = ~n2898 & ~n3068;
  assign n3070 = ~n2584 & n3069;
  assign n3071 = pi03 & ~n2618;
  assign n3072 = ~n2615 & n3071;
  assign n3073 = ~n2605 & n3072;
  assign n3074 = ~n2634 & ~n3073;
  assign n3075 = ~n2619 & ~n3074;
  assign n3076 = n2619 & ~n3073;
  assign n3077 = ~n2634 & n3076;
  assign n3078 = ~n3075 & ~n3077;
  assign n3079 = ~pi05 & ~n3078;
  assign n3080 = pi05 & ~n3077;
  assign n3081 = ~n3075 & n3080;
  assign n3082 = ~n3079 & ~n3081;
  assign n3083 = po04 & ~n3082;
  assign n3084 = ~n3070 & ~n3083;
  assign n3085 = n3063 & n3084;
  assign n3086 = ~n3035 & n3085;
  assign n3087 = po04 & n3079;
  assign n3088 = ~n2898 & n3064;
  assign n3089 = ~n2584 & n3088;
  assign n3090 = ~n3087 & ~n3089;
  assign n3091 = n3063 & ~n3090;
  assign n3092 = po06 & ~n2695;
  assign n3093 = ~n2455 & ~n2659;
  assign n3094 = ~n2454 & n3093;
  assign n3095 = ~n2434 & n3094;
  assign n3096 = ~pi09 & ~n3095;
  assign n3097 = ~n3092 & n3096;
  assign n3098 = ~n2898 & n3097;
  assign n3099 = ~n2584 & n3098;
  assign n3100 = ~n2664 & ~n2698;
  assign n3101 = ~n2653 & ~n2682;
  assign n3102 = ~n2636 & n3101;
  assign n3103 = ~n3100 & ~n3102;
  assign n3104 = n2665 & ~n2682;
  assign n3105 = ~n2698 & n3104;
  assign n3106 = ~n2636 & n3105;
  assign n3107 = ~pi09 & ~n3106;
  assign n3108 = ~n3103 & n3107;
  assign n3109 = po04 & n3108;
  assign n3110 = ~n3099 & ~n3109;
  assign n3111 = ~n2898 & n3041;
  assign n3112 = ~n2584 & n3111;
  assign n3113 = po04 & n3058;
  assign n3114 = ~n3112 & ~n3113;
  assign n3115 = n3110 & n3114;
  assign n3116 = ~n3091 & n3115;
  assign n3117 = ~n3086 & n3116;
  assign n3118 = ~n3092 & ~n3095;
  assign n3119 = ~n2898 & ~n3118;
  assign n3120 = ~n2584 & n3119;
  assign n3121 = ~n3103 & ~n3106;
  assign n3122 = po04 & ~n3121;
  assign n3123 = ~n3120 & ~n3122;
  assign n3124 = pi09 & ~n3123;
  assign n3125 = po06 & ~n2886;
  assign n3126 = ~n2455 & ~n2873;
  assign n3127 = ~n2454 & n3126;
  assign n3128 = ~n2434 & n3127;
  assign n3129 = ~pi13 & ~n3128;
  assign n3130 = ~n3125 & n3129;
  assign n3131 = ~n3125 & ~n3128;
  assign n3132 = pi13 & ~n3131;
  assign n3133 = ~n3130 & ~n3132;
  assign n3134 = ~n2898 & ~n3133;
  assign n3135 = ~n2584 & n3134;
  assign n3136 = ~n2721 & ~n2766;
  assign n3137 = ~n2843 & n3136;
  assign n3138 = ~n2702 & n3137;
  assign n3139 = ~pi11 & ~n3131;
  assign n3140 = pi11 & ~n3128;
  assign n3141 = ~n3125 & n3140;
  assign n3142 = ~n3139 & ~n3141;
  assign n3143 = ~pi13 & ~n3142;
  assign n3144 = pi13 & ~n3141;
  assign n3145 = ~n3139 & n3144;
  assign n3146 = ~n3143 & ~n3145;
  assign n3147 = ~n3138 & ~n3146;
  assign n3148 = n3137 & ~n3145;
  assign n3149 = ~n2702 & n3148;
  assign n3150 = ~n3143 & n3149;
  assign n3151 = ~n3147 & ~n3150;
  assign n3152 = po04 & n3151;
  assign n3153 = ~n3135 & ~n3152;
  assign n3154 = po06 & ~n2676;
  assign n3155 = ~n2455 & ~n2642;
  assign n3156 = ~n2454 & n3155;
  assign n3157 = ~n2434 & n3156;
  assign n3158 = ~pi11 & ~n3157;
  assign n3159 = ~n3154 & n3158;
  assign n3160 = ~n3154 & ~n3157;
  assign n3161 = pi11 & ~n3160;
  assign n3162 = ~n3159 & ~n3161;
  assign n3163 = ~n2898 & ~n3162;
  assign n3164 = ~n2584 & n3163;
  assign n3165 = n2841 & ~n2842;
  assign n3166 = ~n3102 & n3165;
  assign n3167 = ~n3100 & n3165;
  assign n3168 = ~pi11 & ~n2843;
  assign n3169 = ~n3167 & n3168;
  assign n3170 = ~n2702 & n3169;
  assign n3171 = ~n3166 & n3170;
  assign n3172 = ~n2843 & ~n3167;
  assign n3173 = ~n2702 & n3172;
  assign n3174 = ~n3166 & n3173;
  assign n3175 = pi11 & ~n3174;
  assign n3176 = ~n3171 & ~n3175;
  assign n3177 = po04 & ~n3176;
  assign n3178 = ~n3164 & ~n3177;
  assign n3179 = n3153 & n3178;
  assign n3180 = ~n3124 & n3179;
  assign n3181 = ~n3117 & n3180;
  assign n3182 = n2583 & ~n3005;
  assign n3183 = ~n2709 & ~n2747;
  assign n3184 = ~n2836 & n3183;
  assign n3185 = ~n2891 & n3184;
  assign n3186 = ~n2709 & ~n2721;
  assign n3187 = ~n2729 & n3186;
  assign n3188 = ~n2747 & ~n2766;
  assign n3189 = ~n2773 & n3188;
  assign n3190 = n3187 & n3189;
  assign n3191 = n2844 & n3190;
  assign n3192 = ~n2702 & n3191;
  assign n3193 = ~n3185 & ~n3192;
  assign n3194 = ~n2455 & ~n2851;
  assign n3195 = ~n2454 & n3194;
  assign n3196 = ~n2434 & n3195;
  assign n3197 = po06 & n2762;
  assign n3198 = ~n3196 & ~n3197;
  assign n3199 = ~pi17 & ~n3198;
  assign n3200 = pi17 & ~n3196;
  assign n3201 = ~n3197 & n3200;
  assign n3202 = ~n3199 & ~n3201;
  assign n3203 = ~n2478 & ~n3202;
  assign n3204 = ~n3193 & n3203;
  assign n3205 = ~n2478 & n3202;
  assign n3206 = n3193 & n3205;
  assign n3207 = ~n3204 & ~n3206;
  assign n3208 = ~n3182 & ~n3207;
  assign n3209 = ~n2578 & ~n3196;
  assign n3210 = ~n3197 & n3209;
  assign n3211 = ~n2580 & n3210;
  assign n3212 = ~n2473 & n3211;
  assign n3213 = ~n2571 & n3212;
  assign n3214 = ~n3005 & n3213;
  assign n3215 = ~n2475 & n3198;
  assign n3216 = ~n2476 & n3215;
  assign n3217 = ~n2473 & n3216;
  assign n3218 = ~pi19 & ~n3217;
  assign n3219 = ~n3214 & n3218;
  assign n3220 = ~n3208 & n3219;
  assign n3221 = ~n3214 & ~n3217;
  assign n3222 = ~n3208 & n3221;
  assign n3223 = pi19 & ~n3222;
  assign n3224 = ~n3220 & ~n3223;
  assign n3225 = n2730 & ~n2766;
  assign n3226 = ~n2773 & n3225;
  assign n3227 = ~n2843 & n3226;
  assign n3228 = ~n2702 & n3227;
  assign n3229 = ~n2877 & ~n2883;
  assign n3230 = ~n2888 & n3229;
  assign n3231 = ~n2872 & n3230;
  assign n3232 = ~n3228 & n3231;
  assign n3233 = n2796 & ~n3232;
  assign n3234 = n2835 & ~n3233;
  assign n3235 = n2796 & ~n2835;
  assign n3236 = ~n3232 & n3235;
  assign n3237 = ~n3234 & ~n3236;
  assign n3238 = po04 & ~n3237;
  assign n3239 = ~n2455 & n2748;
  assign n3240 = ~n2454 & n3239;
  assign n3241 = ~n2434 & n3240;
  assign n3242 = ~n2319 & ~n2330;
  assign n3243 = ~n2316 & n3242;
  assign n3244 = ~n2327 & n3243;
  assign n3245 = ~n2735 & n3244;
  assign n3246 = ~n2736 & ~n2742;
  assign n3247 = ~n3245 & ~n3246;
  assign n3248 = po06 & n3247;
  assign n3249 = ~n3241 & ~n3248;
  assign n3250 = ~n2898 & n3249;
  assign n3251 = ~n2584 & n3250;
  assign n3252 = ~pi17 & ~n3251;
  assign n3253 = ~n3238 & n3252;
  assign n3254 = ~n3224 & n3253;
  assign n3255 = ~pi19 & ~n3222;
  assign n3256 = ~n2898 & n3130;
  assign n3257 = ~n2584 & n3256;
  assign n3258 = ~n3138 & ~n3142;
  assign n3259 = n3136 & ~n3141;
  assign n3260 = ~n2843 & n3259;
  assign n3261 = ~n3139 & n3260;
  assign n3262 = ~n2702 & n3261;
  assign n3263 = ~pi13 & ~n3262;
  assign n3264 = ~n3258 & n3263;
  assign n3265 = po04 & n3264;
  assign n3266 = ~n3257 & ~n3265;
  assign n3267 = po06 & ~n2869;
  assign n3268 = ~n2455 & ~n2878;
  assign n3269 = ~n2454 & n3268;
  assign n3270 = ~n2434 & n3269;
  assign n3271 = ~pi15 & ~n3270;
  assign n3272 = ~n3267 & n3271;
  assign n3273 = ~n2898 & n3272;
  assign n3274 = ~n2584 & n3273;
  assign n3275 = ~n2872 & ~n2883;
  assign n3276 = ~n2877 & ~n2888;
  assign n3277 = ~n3275 & ~n3276;
  assign n3278 = ~n3231 & ~n3277;
  assign n3279 = ~n3228 & n3278;
  assign n3280 = ~n2721 & ~n2883;
  assign n3281 = ~n2729 & n3280;
  assign n3282 = n2774 & n3281;
  assign n3283 = ~n2872 & n3282;
  assign n3284 = ~n2843 & n3283;
  assign n3285 = ~n2702 & n3284;
  assign n3286 = ~n3279 & ~n3285;
  assign n3287 = ~pi15 & ~n3286;
  assign n3288 = po04 & n3287;
  assign n3289 = ~n3274 & ~n3288;
  assign n3290 = n3266 & n3289;
  assign n3291 = ~n3255 & n3290;
  assign n3292 = ~n2895 & n2907;
  assign n3293 = ~n2846 & n3292;
  assign n3294 = n2864 & ~n3293;
  assign n3295 = ~n2930 & ~n3294;
  assign n3296 = po04 & ~n3295;
  assign n3297 = ~n2860 & ~n2898;
  assign n3298 = ~n2584 & n3297;
  assign n3299 = ~pi21 & ~n3298;
  assign n3300 = ~n3296 & n3299;
  assign n3301 = ~n2898 & n3159;
  assign n3302 = ~n2584 & n3301;
  assign n3303 = po04 & n3171;
  assign n3304 = ~n3302 & ~n3303;
  assign n3305 = n3153 & ~n3304;
  assign n3306 = ~n3300 & ~n3305;
  assign n3307 = n3291 & n3306;
  assign n3308 = ~n3254 & n3307;
  assign n3309 = ~n3181 & n3308;
  assign n3310 = ~n3238 & ~n3251;
  assign n3311 = ~pi17 & ~n3310;
  assign n3312 = pi17 & ~n3251;
  assign n3313 = ~n3238 & n3312;
  assign n3314 = ~n3311 & ~n3313;
  assign n3315 = ~n3267 & ~n3270;
  assign n3316 = ~n2898 & ~n3315;
  assign n3317 = ~n2584 & n3316;
  assign n3318 = po04 & n3286;
  assign n3319 = ~n3317 & ~n3318;
  assign n3320 = pi15 & ~n3319;
  assign n3321 = ~n3224 & ~n3320;
  assign n3322 = ~n3314 & n3321;
  assign n3323 = ~n3255 & ~n3300;
  assign n3324 = ~n3254 & n3323;
  assign n3325 = ~n3322 & n3324;
  assign n3326 = po04 & ~n2934;
  assign n3327 = ~n2932 & n3326;
  assign n3328 = ~n2491 & ~n2898;
  assign n3329 = ~n2584 & n3328;
  assign n3330 = pi23 & ~n3329;
  assign n3331 = ~n3327 & n3330;
  assign n3332 = ~n3296 & ~n3298;
  assign n3333 = pi21 & ~n3332;
  assign n3334 = ~n3331 & ~n3333;
  assign n3335 = ~pi03 & ~pi31;
  assign n3336 = ~n2994 & n3335;
  assign n3337 = ~n2926 & n3336;
  assign n3338 = ~n2937 & n3337;
  assign n3339 = ~n2988 & n3338;
  assign n3340 = n3334 & n3339;
  assign n3341 = n2959 & n3340;
  assign n3342 = ~n2981 & n3341;
  assign n3343 = ~n3325 & n3342;
  assign n3344 = ~n3309 & n3343;
  assign n3345 = ~n2996 & ~n3344;
  assign n3346 = ~n2993 & n3012;
  assign n3347 = ~n2992 & n3346;
  assign n3348 = ~pi31 & n3012;
  assign n3349 = ~n2993 & n3348;
  assign n3350 = ~n2926 & n3349;
  assign n3351 = ~n2937 & n3350;
  assign n3352 = ~n2988 & n3351;
  assign n3353 = n3334 & n3352;
  assign n3354 = n2959 & n3353;
  assign n3355 = ~n2981 & n3354;
  assign n3356 = ~n3325 & n3355;
  assign n3357 = ~n3309 & n3356;
  assign n3358 = ~n3347 & ~n3357;
  assign n3359 = n3345 & n3358;
  assign n3360 = ~pi31 & ~n2926;
  assign n3361 = ~n2937 & n3360;
  assign n3362 = ~n2988 & n3361;
  assign n3363 = n3334 & n3362;
  assign n3364 = n2959 & n3363;
  assign n3365 = ~n2981 & n3364;
  assign n3366 = ~n3325 & n3365;
  assign n3367 = ~n3309 & n3366;
  assign n3368 = n2581 & ~n3016;
  assign n3369 = ~n2571 & n3368;
  assign n3370 = ~n3005 & n3369;
  assign n3371 = n3027 & ~n3370;
  assign n3372 = n3011 & ~n3371;
  assign n3373 = ~n2923 & ~n3372;
  assign n3374 = ~n2991 & n3373;
  assign n3375 = ~n3367 & n3374;
  assign n3376 = ~pi03 & ~n3372;
  assign n3377 = pi03 & ~n3003;
  assign n3378 = ~n3010 & n3377;
  assign n3379 = ~n3371 & n3378;
  assign n3380 = ~n3376 & ~n3379;
  assign n3381 = ~n3012 & ~n3380;
  assign n3382 = n3012 & ~n3379;
  assign n3383 = ~n3376 & n3382;
  assign n3384 = ~n3381 & ~n3383;
  assign n3385 = ~n2992 & ~n3384;
  assign n3386 = n3365 & ~n3384;
  assign n3387 = ~n3309 & ~n3325;
  assign n3388 = n3386 & n3387;
  assign n3389 = ~n3385 & ~n3388;
  assign n3390 = ~n3375 & n3389;
  assign n3391 = ~pi02 & n2993;
  assign n3392 = ~pi03 & ~n3391;
  assign n3393 = ~n2923 & n3392;
  assign n3394 = ~n2991 & n3393;
  assign n3395 = ~n3367 & n3394;
  assign n3396 = ~pi01 & pi02;
  assign n3397 = ~pi31 & ~n3396;
  assign n3398 = ~n2926 & n3397;
  assign n3399 = ~n2937 & n3398;
  assign n3400 = ~n2988 & n3399;
  assign n3401 = n3334 & n3400;
  assign n3402 = n2959 & n3401;
  assign n3403 = ~n2981 & n3402;
  assign n3404 = ~n3325 & n3403;
  assign n3405 = ~n3309 & n3404;
  assign n3406 = pi02 & ~n2993;
  assign n3407 = ~n2923 & n3406;
  assign n3408 = ~n2991 & n3407;
  assign n3409 = ~n3396 & ~n3408;
  assign n3410 = ~n3405 & ~n3409;
  assign n3411 = ~n3395 & ~n3410;
  assign n3412 = n3390 & n3411;
  assign n3413 = n3359 & n3412;
  assign n3414 = n2631 & ~n2898;
  assign n3415 = ~n2584 & n3414;
  assign n3416 = po04 & n3078;
  assign n3417 = ~n3415 & ~n3416;
  assign n3418 = ~n2923 & n3417;
  assign n3419 = ~n2991 & n3418;
  assign n3420 = ~n3367 & n3419;
  assign n3421 = ~n3035 & n3084;
  assign n3422 = n3035 & ~n3084;
  assign n3423 = ~n3421 & ~n3422;
  assign n3424 = ~n2992 & n3423;
  assign n3425 = n2959 & ~n3421;
  assign n3426 = ~n3422 & n3425;
  assign n3427 = ~n2981 & n3363;
  assign n3428 = n3426 & n3427;
  assign n3429 = ~n3325 & n3428;
  assign n3430 = ~n3309 & n3429;
  assign n3431 = ~n3424 & ~n3430;
  assign n3432 = ~n3420 & n3431;
  assign n3433 = ~pi05 & ~n3432;
  assign n3434 = ~n3413 & n3433;
  assign n3435 = ~n2898 & ~n3042;
  assign n3436 = ~n2584 & n3435;
  assign n3437 = po04 & ~n3059;
  assign n3438 = ~n3436 & ~n3437;
  assign n3439 = ~n2923 & ~n3438;
  assign n3440 = ~n2991 & n3439;
  assign n3441 = ~n3367 & n3440;
  assign po02 = ~n2992 | n3367;
  assign n3443 = n3090 & ~n3421;
  assign n3444 = n3063 & ~n3443;
  assign n3445 = ~n3063 & n3090;
  assign n3446 = ~n3421 & n3445;
  assign n3447 = ~n3444 & ~n3446;
  assign n3448 = po02 & ~n3447;
  assign n3449 = ~n3441 & ~n3448;
  assign n3450 = n3359 & n3411;
  assign n3451 = ~n3390 & ~n3432;
  assign n3452 = ~n3450 & n3451;
  assign n3453 = ~n3449 & ~n3452;
  assign n3454 = ~n3434 & n3453;
  assign n3455 = ~pi09 & ~n3454;
  assign n3456 = ~pi05 & ~n3441;
  assign n3457 = ~n3432 & n3456;
  assign n3458 = ~n3448 & n3457;
  assign n3459 = ~n3413 & n3458;
  assign n3460 = ~n2923 & ~n3123;
  assign n3461 = ~n2991 & n3460;
  assign n3462 = ~n3367 & n3461;
  assign n3463 = n3110 & ~n3124;
  assign n3464 = ~n3091 & n3114;
  assign n3465 = ~n3086 & n3464;
  assign n3466 = ~n3463 & n3465;
  assign n3467 = n3463 & ~n3465;
  assign n3468 = ~n3466 & ~n3467;
  assign n3469 = po02 & ~n3468;
  assign n3470 = ~n3462 & ~n3469;
  assign n3471 = n3449 & n3452;
  assign n3472 = ~n3470 & ~n3471;
  assign n3473 = ~n3459 & n3472;
  assign n3474 = ~n3455 & n3473;
  assign n3475 = ~pi05 & ~n3413;
  assign n3476 = ~n3390 & ~n3450;
  assign n3477 = n3432 & ~n3476;
  assign n3478 = ~n3475 & n3477;
  assign n3479 = n92 & ~n3478;
  assign n3480 = ~pi07 & ~n3441;
  assign n3481 = ~n3448 & n3480;
  assign n3482 = ~n3478 & n3481;
  assign n3483 = ~n3479 & ~n3482;
  assign n3484 = n3474 & n3483;
  assign n3485 = ~pi11 & ~n3484;
  assign n3486 = ~n2898 & ~n3160;
  assign n3487 = ~n2584 & n3486;
  assign n3488 = po04 & ~n3174;
  assign n3489 = ~n3487 & ~n3488;
  assign n3490 = ~n2923 & ~n3489;
  assign n3491 = ~n2991 & n3490;
  assign n3492 = ~n3367 & n3491;
  assign n3493 = ~n3124 & n3178;
  assign n3494 = ~n3117 & n3493;
  assign n3495 = ~n3117 & ~n3124;
  assign n3496 = ~n3178 & ~n3495;
  assign n3497 = ~n3494 & ~n3496;
  assign n3498 = po02 & ~n3497;
  assign n3499 = ~n3492 & ~n3498;
  assign n3500 = ~n3459 & ~n3471;
  assign n3501 = n3470 & ~n3500;
  assign n3502 = ~n3499 & ~n3501;
  assign n3503 = n92 & ~n3462;
  assign n3504 = ~n3469 & n3503;
  assign n3505 = ~n3478 & n3504;
  assign n3506 = n3470 & n3481;
  assign n3507 = ~n3478 & n3506;
  assign n3508 = ~pi09 & ~n3462;
  assign n3509 = ~n3469 & n3508;
  assign n3510 = ~n3454 & n3509;
  assign n3511 = ~n3507 & ~n3510;
  assign n3512 = ~n3505 & n3511;
  assign n3513 = n3502 & n3512;
  assign n3514 = ~n3485 & n3513;
  assign n3515 = ~pi13 & ~n3514;
  assign n3516 = ~pi11 & ~n3492;
  assign n3517 = ~n3498 & n3516;
  assign n3518 = ~n3484 & n3517;
  assign n3519 = ~n2898 & ~n3131;
  assign n3520 = ~n2584 & n3519;
  assign n3521 = ~n3258 & ~n3262;
  assign n3522 = po04 & ~n3521;
  assign n3523 = ~n3520 & ~n3522;
  assign n3524 = ~n2923 & ~n3523;
  assign n3525 = ~n2991 & n3524;
  assign n3526 = ~n3367 & n3525;
  assign n3527 = n3304 & ~n3494;
  assign n3528 = n3153 & ~n3527;
  assign n3529 = ~n3153 & n3304;
  assign n3530 = ~n3494 & n3529;
  assign n3531 = ~n3528 & ~n3530;
  assign n3532 = po02 & ~n3531;
  assign n3533 = ~n3526 & ~n3532;
  assign n3534 = ~n3501 & ~n3507;
  assign n3535 = ~n3505 & ~n3510;
  assign n3536 = n3534 & n3535;
  assign n3537 = n3499 & ~n3536;
  assign n3538 = ~n3533 & ~n3537;
  assign n3539 = ~n3518 & n3538;
  assign n3540 = ~n3515 & n3539;
  assign n3541 = ~pi15 & ~n3540;
  assign n3542 = ~pi13 & ~n3526;
  assign n3543 = ~n3532 & n3542;
  assign n3544 = ~n3514 & n3543;
  assign n3545 = ~n2923 & ~n3319;
  assign n3546 = ~n2991 & n3545;
  assign n3547 = ~n3367 & n3546;
  assign n3548 = n3289 & ~n3320;
  assign n3549 = n3266 & ~n3305;
  assign n3550 = ~n3548 & n3549;
  assign n3551 = ~n3181 & n3550;
  assign n3552 = ~n3181 & n3549;
  assign n3553 = n3548 & ~n3552;
  assign n3554 = ~n3551 & ~n3553;
  assign n3555 = po02 & ~n3554;
  assign n3556 = ~n3547 & ~n3555;
  assign n3557 = ~n3518 & ~n3537;
  assign n3558 = n3533 & ~n3557;
  assign n3559 = ~n3556 & ~n3558;
  assign n3560 = ~n3544 & n3559;
  assign n3561 = ~n3541 & n3560;
  assign n3562 = ~pi17 & ~n3561;
  assign n3563 = ~pi15 & ~n3547;
  assign n3564 = ~n3555 & n3563;
  assign n3565 = ~n3540 & n3564;
  assign n3566 = ~n2923 & ~n3310;
  assign n3567 = ~n2991 & n3566;
  assign n3568 = ~n3367 & n3567;
  assign n3569 = n3290 & ~n3305;
  assign n3570 = ~n3181 & n3569;
  assign n3571 = ~n3320 & ~n3570;
  assign n3572 = n3314 & ~n3571;
  assign n3573 = ~n3314 & ~n3320;
  assign n3574 = ~n3570 & n3573;
  assign n3575 = ~n3572 & ~n3574;
  assign n3576 = po02 & ~n3575;
  assign n3577 = ~n3568 & ~n3576;
  assign n3578 = ~n3544 & ~n3558;
  assign n3579 = n3556 & ~n3578;
  assign n3580 = ~n3577 & ~n3579;
  assign n3581 = ~n3565 & n3580;
  assign n3582 = ~n3562 & n3581;
  assign n3583 = ~pi19 & ~n3582;
  assign n3584 = ~pi17 & ~n3568;
  assign n3585 = ~n3576 & n3584;
  assign n3586 = ~n3561 & n3585;
  assign n3587 = ~n2923 & n3222;
  assign n3588 = ~n2991 & n3587;
  assign n3589 = ~n3367 & n3588;
  assign n3590 = n3224 & ~n3253;
  assign n3591 = ~n3574 & n3590;
  assign n3592 = ~n3253 & ~n3574;
  assign n3593 = ~n3224 & ~n3592;
  assign n3594 = ~n3591 & ~n3593;
  assign n3595 = po02 & ~n3594;
  assign n3596 = ~n3589 & ~n3595;
  assign n3597 = ~n3565 & ~n3579;
  assign n3598 = n3577 & ~n3597;
  assign n3599 = ~n3596 & ~n3598;
  assign n3600 = ~n3586 & n3599;
  assign n3601 = ~n3583 & n3600;
  assign n3602 = ~pi21 & ~n3601;
  assign n3603 = ~pi19 & ~n3589;
  assign n3604 = ~n3595 & n3603;
  assign n3605 = ~n3582 & n3604;
  assign n3606 = ~n2923 & ~n3332;
  assign n3607 = ~n2991 & n3606;
  assign n3608 = ~n3367 & n3607;
  assign n3609 = n3322 & ~n3570;
  assign n3610 = ~n3300 & ~n3333;
  assign n3611 = ~n3255 & ~n3610;
  assign n3612 = ~n3254 & n3611;
  assign n3613 = ~n3609 & n3612;
  assign n3614 = ~n3254 & ~n3255;
  assign n3615 = ~n3609 & n3614;
  assign n3616 = n3610 & ~n3615;
  assign n3617 = ~n3613 & ~n3616;
  assign n3618 = po02 & ~n3617;
  assign n3619 = ~n3608 & ~n3618;
  assign n3620 = ~n3586 & ~n3598;
  assign n3621 = n3596 & ~n3620;
  assign n3622 = ~n3619 & ~n3621;
  assign n3623 = ~n3605 & n3622;
  assign n3624 = ~n3602 & n3623;
  assign n3625 = ~pi23 & ~n3624;
  assign n3626 = ~pi21 & ~n3608;
  assign n3627 = ~n3618 & n3626;
  assign n3628 = ~n3601 & n3627;
  assign n3629 = ~n3327 & ~n3329;
  assign n3630 = ~n2923 & n3629;
  assign n3631 = ~n2991 & n3630;
  assign n3632 = ~n3367 & n3631;
  assign n3633 = n2938 & ~n3331;
  assign n3634 = ~n3325 & ~n3333;
  assign n3635 = ~n3309 & n3634;
  assign n3636 = ~n3633 & ~n3635;
  assign n3637 = ~n3333 & n3633;
  assign n3638 = ~n3325 & n3637;
  assign n3639 = ~n3309 & n3638;
  assign n3640 = ~n3636 & ~n3639;
  assign n3641 = po02 & ~n3640;
  assign n3642 = ~n3632 & ~n3641;
  assign n3643 = ~n3605 & ~n3621;
  assign n3644 = n3619 & ~n3643;
  assign n3645 = ~n3642 & ~n3644;
  assign n3646 = ~n3628 & n3645;
  assign n3647 = ~n3625 & n3646;
  assign n3648 = ~pi25 & ~n3647;
  assign n3649 = ~n3628 & ~n3644;
  assign n3650 = n3642 & ~n3649;
  assign n3651 = ~n2966 & ~n2968;
  assign n3652 = ~n2923 & ~n3651;
  assign n3653 = ~n2991 & n3652;
  assign n3654 = ~n3367 & n3653;
  assign n3655 = n2938 & ~n3639;
  assign n3656 = n2959 & ~n3655;
  assign n3657 = n2938 & ~n2959;
  assign n3658 = ~n3639 & n3657;
  assign n3659 = ~n3656 & ~n3658;
  assign n3660 = po02 & ~n3659;
  assign n3661 = ~n3654 & ~n3660;
  assign n3662 = ~pi23 & ~n3632;
  assign n3663 = ~n3641 & n3662;
  assign n3664 = ~n3624 & n3663;
  assign n3665 = ~n3661 & ~n3664;
  assign n3666 = ~n3650 & n3665;
  assign n3667 = ~n3648 & n3666;
  assign n3668 = ~pi27 & ~n3667;
  assign n3669 = ~pi25 & ~n3654;
  assign n3670 = ~n3660 & n3669;
  assign n3671 = ~n3647 & n3670;
  assign n3672 = ~n2983 & ~n2986;
  assign n3673 = ~n2923 & n3672;
  assign n3674 = ~n2991 & n3673;
  assign n3675 = ~n3367 & n3674;
  assign n3676 = ~n2926 & ~n2957;
  assign n3677 = ~n2937 & n3676;
  assign n3678 = ~n2947 & ~n2950;
  assign n3679 = n3677 & n3678;
  assign n3680 = n3334 & n3679;
  assign n3681 = ~n3325 & n3680;
  assign n3682 = ~n3309 & n3681;
  assign n3683 = ~n2974 & ~n2988;
  assign n3684 = ~n2965 & n3683;
  assign n3685 = ~n2960 & ~n2970;
  assign n3686 = ~n3684 & n3685;
  assign n3687 = ~n3682 & n3686;
  assign n3688 = ~n3682 & n3685;
  assign n3689 = n3684 & ~n3688;
  assign n3690 = ~n3687 & ~n3689;
  assign n3691 = po02 & ~n3690;
  assign n3692 = ~n3675 & ~n3691;
  assign n3693 = ~n3650 & ~n3664;
  assign n3694 = n3661 & ~n3693;
  assign n3695 = ~n3692 & ~n3694;
  assign n3696 = ~n3671 & n3695;
  assign n3697 = ~n3668 & n3696;
  assign n3698 = ~pi29 & ~n3697;
  assign n3699 = ~pi27 & ~n3675;
  assign n3700 = ~n3691 & n3699;
  assign n3701 = ~n3667 & n3700;
  assign n3702 = ~n3671 & ~n3694;
  assign n3703 = n3692 & ~n3702;
  assign n3704 = ~n3701 & ~n3703;
  assign n3705 = ~n3698 & n3704;
  assign n3706 = n2977 & ~n3682;
  assign n3707 = ~n2979 & ~n2988;
  assign n3708 = ~n2980 & n3707;
  assign n3709 = po02 & n3708;
  assign n3710 = ~n3706 & n3709;
  assign n3711 = ~n2922 & ~n2923;
  assign n3712 = ~n2991 & n3711;
  assign n3713 = ~n3367 & n3712;
  assign n3714 = pi31 & ~n3713;
  assign n3715 = ~n3710 & n3714;
  assign n3716 = ~n3705 & ~n3715;
  assign n3717 = ~n3710 & ~n3713;
  assign n3718 = ~pi31 & ~n3717;
  assign po00 = n3716 | n3718;
  assign n3720 = n93 & ~n94;
  assign n3721 = n203 & n3720;
  assign n3722 = n115 & ~n3721;
  assign n3723 = ~n105 & ~n3722;
  assign n3724 = ~pi05 & ~n3723;
  assign n3725 = pi03 & ~n85;
  assign n3726 = ~n77 & ~n3725;
  assign n3727 = n120 & ~n3726;
  assign n3728 = pi30 & ~n3727;
  assign n3729 = ~n3724 & ~n3728;
  assign n3730 = n132 & ~n3722;
  assign n3731 = n181 & ~n3730;
  assign n3732 = ~n3724 & n3731;
  assign n3733 = ~n3729 & n3732;
  assign n3734 = n147 & n179;
  assign n3735 = ~n3727 & n3734;
  assign n3736 = ~n3733 & n3735;
  assign n3737 = n117 & n1150;
  assign n3738 = ~pi19 & ~pi31;
  assign n3739 = n68 & n3738;
  assign n3740 = n285 & n3739;
  assign n3741 = n3737 & n3740;
  assign n3742 = ~n3730 & n3741;
  assign n3743 = ~n3729 & n3742;
  assign n3744 = pi26 & ~n3743;
  assign n3745 = n71 & n155;
  assign n3746 = n78 & n1150;
  assign n3747 = n3745 & n3746;
  assign n3748 = ~pi19 & ~pi26;
  assign n3749 = n73 & n3748;
  assign n3750 = n284 & n3749;
  assign n3751 = n3747 & n3750;
  assign n3752 = ~n3730 & n3751;
  assign n3753 = ~n3729 & n3752;
  assign n3754 = ~n3744 & ~n3753;
  assign n3755 = ~n225 & ~n3754;
  assign n3756 = ~n189 & ~n3755;
  assign n3757 = pi28 & ~pi31;
  assign n3758 = n66 & n3757;
  assign n3759 = n99 & n3758;
  assign n3760 = ~n105 & n3759;
  assign n3761 = n179 & n3760;
  assign n3762 = ~n3721 & n3761;
  assign n3763 = ~n3730 & n3762;
  assign n3764 = ~n3729 & n3763;
  assign n3765 = pi28 & ~n3721;
  assign n3766 = ~n104 & n193;
  assign n3767 = n117 & n3766;
  assign n3768 = n119 & n3767;
  assign n3769 = ~n3730 & n3768;
  assign n3770 = ~n3729 & n3769;
  assign n3771 = ~n3765 & ~n3770;
  assign n3772 = ~n3764 & ~n3771;
  assign n3773 = pi05 & ~n3772;
  assign n3774 = ~n3756 & ~n3773;
  assign n3775 = ~pi05 & ~n3764;
  assign n3776 = ~n3771 & n3775;
  assign n3777 = ~n3774 & ~n3776;
  assign n3778 = n3728 & ~n3733;
  assign n3779 = pi07 & ~n3778;
  assign n3780 = n259 & ~n3779;
  assign n3781 = ~n3777 & n3780;
  assign n3782 = ~n3736 & ~n3781;
  assign n3783 = ~pi07 & ~n3777;
  assign n3784 = ~n3782 & ~n3783;
  assign n3785 = ~pi09 & pi30;
  assign n3786 = ~n3727 & n3785;
  assign n3787 = ~n3733 & n3786;
  assign n3788 = ~n3784 & n3787;
  assign n3789 = pi05 & ~n3764;
  assign n3790 = ~n3771 & n3789;
  assign n3791 = ~n189 & ~n3790;
  assign n3792 = ~n3755 & n3791;
  assign n3793 = ~pi05 & ~n3792;
  assign n3794 = ~n3782 & ~n3793;
  assign n3795 = n3772 & ~n3794;
  assign n3796 = ~n3774 & ~n3792;
  assign n3797 = ~n3782 & n3796;
  assign n3798 = pi07 & ~n3797;
  assign n3799 = ~n3795 & n3798;
  assign n3800 = ~n263 & ~n3782;
  assign n3801 = ~n3754 & ~n3800;
  assign n3802 = ~n263 & ~n3753;
  assign n3803 = ~n3744 & n3802;
  assign n3804 = ~n3782 & n3803;
  assign n3805 = pi05 & ~n3804;
  assign n3806 = ~n3801 & n3805;
  assign n3807 = pi01 & ~n3782;
  assign n3808 = pi24 & ~n3807;
  assign n3809 = n188 & ~n3782;
  assign n3810 = ~n3808 & ~n3809;
  assign n3811 = ~n275 & ~n3810;
  assign n3812 = ~n278 & ~n3811;
  assign n3813 = ~n3806 & ~n3812;
  assign n3814 = ~n3795 & ~n3797;
  assign n3815 = ~pi07 & ~n3814;
  assign n3816 = ~n3801 & ~n3804;
  assign n3817 = ~pi05 & ~n3816;
  assign n3818 = ~n3815 & ~n3817;
  assign n3819 = ~n3813 & n3818;
  assign n3820 = ~n3799 & ~n3819;
  assign n3821 = ~n3788 & ~n3820;
  assign n3822 = n3778 & ~n3784;
  assign n3823 = pi09 & ~n3822;
  assign n3824 = ~pi11 & ~pi19;
  assign n3825 = n73 & n3824;
  assign n3826 = n71 & n1150;
  assign n3827 = n3825 & n3826;
  assign n3828 = n69 & n3827;
  assign n3829 = ~n3823 & n3828;
  assign n3830 = ~n3821 & n3829;
  assign n3831 = pi22 & ~n3830;
  assign n3832 = n71 & n3824;
  assign n3833 = n1150 & n3832;
  assign n3834 = ~pi22 & ~pi25;
  assign n3835 = n73 & n3834;
  assign n3836 = n67 & n3835;
  assign n3837 = n3833 & n3836;
  assign n3838 = ~n3823 & n3837;
  assign n3839 = ~n3821 & n3838;
  assign n3840 = ~n3831 & ~n3839;
  assign n3841 = ~n524 & ~n3840;
  assign n3842 = ~pi03 & ~n527;
  assign n3843 = ~n3841 & ~n3842;
  assign n3844 = n203 & ~n3823;
  assign n3845 = ~n3806 & ~n3817;
  assign n3846 = n3812 & ~n3845;
  assign n3847 = ~pi05 & ~n3846;
  assign n3848 = n3844 & ~n3847;
  assign n3849 = ~n3821 & n3848;
  assign n3850 = ~n3816 & ~n3849;
  assign n3851 = ~n3813 & n3844;
  assign n3852 = ~n3846 & n3851;
  assign n3853 = ~n3821 & n3852;
  assign n3854 = ~pi07 & ~n3853;
  assign n3855 = ~n3850 & n3854;
  assign n3856 = pi07 & ~pi11;
  assign n3857 = n71 & n3856;
  assign n3858 = n74 & n3857;
  assign n3859 = n69 & n3858;
  assign n3860 = ~n3823 & n3859;
  assign n3861 = ~n3813 & n3860;
  assign n3862 = ~n3846 & n3861;
  assign n3863 = ~n3821 & n3862;
  assign n3864 = pi07 & ~n3816;
  assign n3865 = ~n3849 & n3864;
  assign n3866 = ~n3863 & ~n3865;
  assign n3867 = ~n3855 & n3866;
  assign n3868 = pi05 & ~n3810;
  assign n3869 = n67 & ~n275;
  assign n3870 = ~n278 & n3869;
  assign n3871 = n103 & n3870;
  assign n3872 = ~n3823 & n3871;
  assign n3873 = ~pi05 & ~n3809;
  assign n3874 = ~n3808 & n3873;
  assign n3875 = n3872 & ~n3874;
  assign n3876 = ~n3868 & n3875;
  assign n3877 = ~n3821 & n3876;
  assign n3878 = ~n3821 & n3872;
  assign n3879 = ~n3868 & ~n3874;
  assign n3880 = ~n3878 & ~n3879;
  assign n3881 = ~n3877 & ~n3880;
  assign n3882 = ~n3867 & ~n3881;
  assign n3883 = ~n3843 & n3882;
  assign n3884 = n3810 & ~n3878;
  assign n3885 = ~n3810 & n3872;
  assign n3886 = ~n3821 & n3885;
  assign n3887 = ~pi05 & ~n3886;
  assign n3888 = ~n3884 & n3887;
  assign n3889 = ~n3867 & n3888;
  assign n3890 = ~n3821 & n3844;
  assign n3891 = n3814 & ~n3890;
  assign n3892 = ~n3799 & ~n3815;
  assign n3893 = ~n3813 & ~n3817;
  assign n3894 = ~n3892 & ~n3893;
  assign n3895 = ~n3817 & n3892;
  assign n3896 = ~n3813 & n3895;
  assign n3897 = n3844 & ~n3896;
  assign n3898 = ~n3894 & n3897;
  assign n3899 = ~n3821 & n3898;
  assign n3900 = ~pi09 & ~n3899;
  assign n3901 = ~n3891 & n3900;
  assign n3902 = ~n3850 & ~n3853;
  assign n3903 = ~pi07 & ~n3902;
  assign n3904 = ~n3901 & ~n3903;
  assign n3905 = ~n3889 & n3904;
  assign n3906 = ~n3883 & n3905;
  assign n3907 = ~n3891 & ~n3899;
  assign n3908 = ~pi09 & ~n3907;
  assign n3909 = pi09 & ~n3899;
  assign n3910 = ~n3891 & n3909;
  assign n3911 = ~n3901 & ~n3910;
  assign n3912 = ~n3908 & n3911;
  assign n3913 = n3822 & ~n3890;
  assign n3914 = n3788 & ~n3799;
  assign n3915 = ~n3819 & n3914;
  assign n3916 = ~n3913 & ~n3915;
  assign n3917 = ~pi11 & ~n3916;
  assign n3918 = pi11 & ~n3915;
  assign n3919 = ~n3913 & n3918;
  assign n3920 = n76 & ~n3919;
  assign n3921 = ~n3917 & n3920;
  assign n3922 = ~n3912 & n3921;
  assign n3923 = ~n3906 & n3922;
  assign n3924 = n203 & ~n3916;
  assign n3925 = ~n3923 & ~n3924;
  assign n3926 = ~n3843 & ~n3881;
  assign n3927 = ~n3842 & ~n3877;
  assign n3928 = ~n3880 & n3927;
  assign n3929 = ~n3841 & n3928;
  assign n3930 = ~n3926 & ~n3929;
  assign n3931 = ~n3925 & ~n3930;
  assign n3932 = ~n3884 & ~n3886;
  assign n3933 = ~n3924 & ~n3932;
  assign n3934 = ~n3923 & n3933;
  assign n3935 = ~pi07 & ~n3934;
  assign n3936 = ~n3931 & n3935;
  assign n3937 = n3840 & ~n3924;
  assign n3938 = ~n3923 & n3937;
  assign n3939 = ~n524 & ~n3842;
  assign n3940 = ~n3839 & n3939;
  assign n3941 = ~n3831 & n3940;
  assign n3942 = ~n3840 & ~n3939;
  assign n3943 = ~n3941 & ~n3942;
  assign n3944 = ~n3925 & n3943;
  assign n3945 = ~n3938 & ~n3944;
  assign n3946 = ~pi05 & ~n3945;
  assign n3947 = ~pi05 & ~n3938;
  assign n3948 = ~n3944 & n3947;
  assign n3949 = pi05 & ~n3938;
  assign n3950 = ~n3944 & n3949;
  assign n3951 = ~n3948 & ~n3950;
  assign n3952 = ~n3946 & n3951;
  assign n3953 = ~pi01 & ~pi20;
  assign n3954 = ~n3924 & ~n3953;
  assign n3955 = ~n3923 & n3954;
  assign n3956 = n564 & ~n3955;
  assign n3957 = ~pi20 & ~n3924;
  assign n3958 = ~n3923 & n3957;
  assign n3959 = ~n3956 & ~n3958;
  assign n3960 = n568 & ~n3959;
  assign n3961 = ~pi03 & ~n3958;
  assign n3962 = ~n3956 & n3961;
  assign n3963 = n572 & ~n3958;
  assign n3964 = ~n3956 & n3963;
  assign n3965 = ~n3948 & ~n3964;
  assign n3966 = ~n3962 & n3965;
  assign n3967 = ~n3960 & n3966;
  assign n3968 = ~n3952 & ~n3967;
  assign n3969 = ~n3936 & ~n3968;
  assign n3970 = n3867 & ~n3888;
  assign n3971 = ~n3926 & n3970;
  assign n3972 = ~n3883 & ~n3889;
  assign n3973 = ~n3971 & n3972;
  assign n3974 = ~n3925 & n3973;
  assign n3975 = ~n3902 & ~n3924;
  assign n3976 = ~n3923 & n3975;
  assign n3977 = ~pi09 & ~n3976;
  assign n3978 = ~n3974 & n3977;
  assign n3979 = ~n3974 & ~n3976;
  assign n3980 = pi09 & ~n3979;
  assign n3981 = ~n3978 & ~n3980;
  assign n3982 = ~n3931 & ~n3934;
  assign n3983 = pi07 & ~n3982;
  assign n3984 = ~n3981 & ~n3983;
  assign n3985 = ~n3969 & n3984;
  assign n3986 = ~n3908 & ~n3910;
  assign n3987 = ~n3903 & n3986;
  assign n3988 = ~n3889 & n3987;
  assign n3989 = ~n3883 & n3988;
  assign n3990 = ~n3889 & ~n3903;
  assign n3991 = ~n3883 & n3990;
  assign n3992 = ~n3986 & ~n3991;
  assign n3993 = ~n3989 & ~n3992;
  assign n3994 = ~n3925 & ~n3993;
  assign n3995 = ~n3907 & ~n3924;
  assign n3996 = ~n3923 & n3995;
  assign n3997 = ~pi11 & ~n3996;
  assign n3998 = ~n3994 & n3997;
  assign n3999 = ~pi09 & ~n3979;
  assign n4000 = ~n3998 & ~n3999;
  assign n4001 = ~n3985 & n4000;
  assign n4002 = ~n3994 & ~n3996;
  assign n4003 = pi11 & ~n4002;
  assign n4004 = ~n3916 & ~n3924;
  assign n4005 = ~n3923 & n4004;
  assign n4006 = ~n3912 & n3924;
  assign n4007 = ~n3906 & n4006;
  assign n4008 = pi13 & ~n4007;
  assign n4009 = ~n4005 & n4008;
  assign n4010 = n740 & ~n4009;
  assign n4011 = ~n4003 & n4010;
  assign n4012 = ~n4001 & n4011;
  assign n4013 = ~n4005 & ~n4007;
  assign n4014 = n76 & ~n4013;
  assign n4015 = ~n4013 & ~n4014;
  assign n4016 = ~n4012 & n4015;
  assign n4017 = ~n4003 & n4014;
  assign n4018 = ~n4001 & n4017;
  assign n4019 = ~pi15 & ~n4018;
  assign n4020 = ~n4016 & n4019;
  assign n4021 = ~n4016 & ~n4018;
  assign n4022 = pi15 & ~n4021;
  assign n4023 = ~n4020 & ~n4022;
  assign n4024 = pi16 & ~pi19;
  assign n4025 = n73 & n4024;
  assign n4026 = n1150 & n4025;
  assign n4027 = n69 & n4026;
  assign n4028 = ~n4023 & n4027;
  assign n4029 = ~pi01 & ~pi16;
  assign n4030 = ~pi15 & pi16;
  assign n4031 = n1150 & n4030;
  assign n4032 = n99 & n4031;
  assign n4033 = n67 & n4032;
  assign n4034 = ~n4021 & n4033;
  assign n4035 = ~n4029 & ~n4034;
  assign n4036 = ~n4028 & n4035;
  assign n4037 = ~n4012 & ~n4014;
  assign n4038 = n823 & ~n3958;
  assign n4039 = ~n3956 & n4038;
  assign n4040 = ~n823 & ~n3959;
  assign n4041 = ~n4039 & ~n4040;
  assign n4042 = ~pi05 & ~n4041;
  assign n4043 = pi05 & ~n4039;
  assign n4044 = ~n4040 & n4043;
  assign n4045 = ~n4042 & ~n4044;
  assign n4046 = ~n4037 & ~n4045;
  assign n4047 = n768 & ~n4037;
  assign n4048 = ~n3946 & ~n3950;
  assign n4049 = ~n3962 & ~n3964;
  assign n4050 = ~n3960 & n4049;
  assign n4051 = ~n4048 & ~n4050;
  assign n4052 = ~n3950 & ~n3964;
  assign n4053 = ~n3962 & n4052;
  assign n4054 = ~n3946 & ~n3960;
  assign n4055 = n4053 & n4054;
  assign n4056 = ~pi07 & ~n4055;
  assign n4057 = ~n4051 & n4056;
  assign n4058 = ~n4051 & ~n4055;
  assign n4059 = pi07 & ~n4058;
  assign n4060 = ~n4057 & ~n4059;
  assign n4061 = ~n4037 & ~n4060;
  assign n4062 = ~n4047 & ~n4061;
  assign n4063 = ~n4046 & n4062;
  assign n4064 = pi03 & ~n4014;
  assign n4065 = ~n4012 & n4064;
  assign n4066 = n785 & ~n4065;
  assign n4067 = n788 & ~n4014;
  assign n4068 = ~n4012 & n4067;
  assign n4069 = ~n787 & ~n4068;
  assign n4070 = ~n4066 & n4069;
  assign n4071 = ~pi05 & ~n3958;
  assign n4072 = ~n3956 & n4071;
  assign n4073 = pi05 & ~n3959;
  assign n4074 = ~n4072 & ~n4073;
  assign n4075 = ~n4014 & ~n4074;
  assign n4076 = ~n4012 & n4075;
  assign n4077 = ~pi18 & n767;
  assign n4078 = ~n4014 & n4077;
  assign n4079 = ~n4012 & n4078;
  assign n4080 = ~pi07 & ~n3938;
  assign n4081 = ~n3944 & n4080;
  assign n4082 = pi07 & ~n3945;
  assign n4083 = ~n4081 & ~n4082;
  assign n4084 = ~n4014 & ~n4083;
  assign n4085 = ~n4012 & n4084;
  assign n4086 = ~n4079 & ~n4085;
  assign n4087 = ~n4076 & n4086;
  assign n4088 = ~n4070 & n4087;
  assign n4089 = n4063 & n4088;
  assign n4090 = ~n4014 & n4072;
  assign n4091 = ~n4012 & n4090;
  assign n4092 = ~n4037 & n4042;
  assign n4093 = ~n4091 & ~n4092;
  assign n4094 = ~n4061 & ~n4085;
  assign n4095 = ~n4093 & n4094;
  assign n4096 = ~n4037 & n4057;
  assign n4097 = ~n3936 & ~n3983;
  assign n4098 = ~n3968 & ~n4097;
  assign n4099 = ~n3952 & n4097;
  assign n4100 = ~n3967 & n4099;
  assign n4101 = ~pi09 & ~n4100;
  assign n4102 = ~n4098 & n4101;
  assign n4103 = ~n4037 & n4102;
  assign n4104 = ~pi09 & ~n3934;
  assign n4105 = ~n3931 & n4104;
  assign n4106 = ~n4014 & n4105;
  assign n4107 = ~n4012 & n4106;
  assign n4108 = ~n4014 & n4081;
  assign n4109 = ~n4012 & n4108;
  assign n4110 = ~n4107 & ~n4109;
  assign n4111 = ~n4103 & n4110;
  assign n4112 = ~n4096 & n4111;
  assign n4113 = ~n4095 & n4112;
  assign n4114 = ~n4089 & n4113;
  assign n4115 = ~n4002 & ~n4014;
  assign n4116 = ~n4012 & n4115;
  assign n4117 = ~n3998 & ~n4003;
  assign n4118 = ~n3999 & ~n4117;
  assign n4119 = ~n3985 & n4118;
  assign n4120 = ~n3985 & ~n3999;
  assign n4121 = n4117 & ~n4120;
  assign n4122 = ~n4119 & ~n4121;
  assign n4123 = ~n4037 & ~n4122;
  assign n4124 = ~n4116 & ~n4123;
  assign n4125 = ~pi13 & ~n4124;
  assign n4126 = pi13 & ~n4116;
  assign n4127 = ~n4123 & n4126;
  assign n4128 = ~n4125 & ~n4127;
  assign n4129 = ~n3982 & ~n4014;
  assign n4130 = ~n4012 & n4129;
  assign n4131 = ~n4098 & ~n4100;
  assign n4132 = ~n4037 & ~n4131;
  assign n4133 = ~n4130 & ~n4132;
  assign n4134 = pi09 & ~n4133;
  assign n4135 = ~pi11 & ~n3979;
  assign n4136 = pi11 & ~n3976;
  assign n4137 = ~n3974 & n4136;
  assign n4138 = ~n4135 & ~n4137;
  assign n4139 = ~n4014 & ~n4138;
  assign n4140 = ~n4012 & n4139;
  assign n4141 = ~n3936 & ~n3978;
  assign n4142 = ~n3980 & n4141;
  assign n4143 = ~n4100 & n4142;
  assign n4144 = ~pi11 & ~n4143;
  assign n4145 = ~n3985 & n4144;
  assign n4146 = ~n3985 & ~n4143;
  assign n4147 = pi11 & ~n4146;
  assign n4148 = ~n4145 & ~n4147;
  assign n4149 = ~n4037 & ~n4148;
  assign n4150 = ~n4140 & ~n4149;
  assign n4151 = ~n4134 & n4150;
  assign n4152 = ~n4128 & n4151;
  assign n4153 = ~n4114 & n4152;
  assign n4154 = ~n4014 & n4135;
  assign n4155 = ~n4012 & n4154;
  assign n4156 = ~n4037 & n4145;
  assign n4157 = ~n4155 & ~n4156;
  assign n4158 = ~n4124 & n4157;
  assign n4159 = ~pi13 & ~n4158;
  assign n4160 = n4124 & ~n4157;
  assign n4161 = n4035 & ~n4160;
  assign n4162 = ~n4159 & n4161;
  assign n4163 = ~n4153 & n4162;
  assign n4164 = ~n4036 & ~n4163;
  assign n4165 = n119 & ~n4023;
  assign n4166 = n740 & ~n4021;
  assign n4167 = ~pi16 & ~n4166;
  assign n4168 = ~n4165 & n4167;
  assign n4169 = ~n4160 & n4167;
  assign n4170 = ~n4159 & n4169;
  assign n4171 = ~n4153 & n4170;
  assign n4172 = ~n4168 & ~n4171;
  assign n4173 = ~n4164 & n4172;
  assign n4174 = n974 & ~n4173;
  assign n4175 = n983 & ~n4168;
  assign n4176 = ~n4171 & n4175;
  assign n4177 = ~n4164 & n4176;
  assign n4178 = ~n4165 & ~n4166;
  assign n4179 = ~n4160 & ~n4166;
  assign n4180 = ~n4159 & n4179;
  assign n4181 = ~n4153 & n4180;
  assign n4182 = ~n4178 & ~n4181;
  assign n4183 = pi01 & ~n4037;
  assign n4184 = pi18 & ~n4183;
  assign n4185 = n567 & ~n4037;
  assign n4186 = ~n4184 & ~n4185;
  assign n4187 = ~pi05 & ~n4186;
  assign n4188 = ~n4182 & n4187;
  assign n4189 = ~n4177 & ~n4188;
  assign n4190 = ~pi03 & ~n4186;
  assign n4191 = pi03 & ~n4185;
  assign n4192 = ~n4184 & n4191;
  assign n4193 = ~n4190 & ~n4192;
  assign n4194 = ~n767 & ~n4193;
  assign n4195 = n767 & ~n4192;
  assign n4196 = ~n4190 & n4195;
  assign n4197 = ~n4194 & ~n4196;
  assign n4198 = ~pi05 & ~n4178;
  assign n4199 = ~n4181 & n4198;
  assign n4200 = ~n4197 & n4199;
  assign n4201 = ~pi03 & ~n4168;
  assign n4202 = ~n4171 & n4201;
  assign n4203 = ~n4164 & n4202;
  assign n4204 = ~n4200 & ~n4203;
  assign n4205 = n4189 & n4204;
  assign n4206 = ~n4174 & n4205;
  assign n4207 = pi05 & ~n4185;
  assign n4208 = ~n4184 & n4207;
  assign n4209 = ~n4182 & n4208;
  assign n4210 = pi05 & ~n4178;
  assign n4211 = n4197 & n4210;
  assign n4212 = ~n4181 & n4211;
  assign n4213 = ~n4209 & ~n4212;
  assign n4214 = ~n4037 & ~n4058;
  assign n4215 = ~n3945 & ~n4014;
  assign n4216 = ~n4012 & n4215;
  assign n4217 = ~pi09 & ~n4216;
  assign n4218 = ~n4214 & n4217;
  assign n4219 = ~n4214 & ~n4216;
  assign n4220 = pi09 & ~n4219;
  assign n4221 = ~n4218 & ~n4220;
  assign n4222 = ~n4182 & ~n4221;
  assign n4223 = ~n4076 & ~n4079;
  assign n4224 = ~n4047 & n4223;
  assign n4225 = ~n4046 & n4224;
  assign n4226 = ~n4070 & n4225;
  assign n4227 = n4093 & ~n4094;
  assign n4228 = ~n4226 & n4227;
  assign n4229 = ~pi09 & ~n4095;
  assign n4230 = ~n4089 & n4229;
  assign n4231 = ~n4228 & n4230;
  assign n4232 = ~n4089 & ~n4095;
  assign n4233 = ~n4228 & n4232;
  assign n4234 = pi09 & ~n4233;
  assign n4235 = ~n4231 & ~n4234;
  assign n4236 = n4182 & ~n4235;
  assign n4237 = ~n4222 & ~n4236;
  assign n4238 = ~n4037 & n4041;
  assign n4239 = ~n3959 & ~n4014;
  assign n4240 = ~n4012 & n4239;
  assign n4241 = ~pi07 & ~n4240;
  assign n4242 = ~n4238 & n4241;
  assign n4243 = ~n4238 & ~n4240;
  assign n4244 = pi07 & ~n4243;
  assign n4245 = ~n4242 & ~n4244;
  assign n4246 = ~n4182 & ~n4245;
  assign n4247 = ~n4047 & ~n4079;
  assign n4248 = ~n4070 & n4247;
  assign n4249 = ~n4046 & ~n4076;
  assign n4250 = ~n4248 & ~n4249;
  assign n4251 = ~pi07 & ~n4226;
  assign n4252 = ~n4250 & n4251;
  assign n4253 = ~n4226 & ~n4250;
  assign n4254 = pi07 & ~n4253;
  assign n4255 = ~n4252 & ~n4254;
  assign n4256 = n4182 & ~n4255;
  assign n4257 = ~n4246 & ~n4256;
  assign n4258 = n4237 & n4257;
  assign n4259 = n4213 & n4258;
  assign n4260 = ~n4206 & n4259;
  assign n4261 = ~n4127 & n4150;
  assign n4262 = ~n4125 & n4261;
  assign n4263 = ~n4134 & n4262;
  assign n4264 = ~n4114 & n4263;
  assign n4265 = ~n4127 & ~n4157;
  assign n4266 = ~n4125 & n4265;
  assign n4267 = ~n4128 & n4157;
  assign n4268 = ~n4266 & ~n4267;
  assign n4269 = ~n4264 & n4268;
  assign n4270 = ~n4153 & ~n4178;
  assign n4271 = ~n4181 & n4270;
  assign n4272 = ~n4269 & n4271;
  assign n4273 = n4124 & ~n4166;
  assign n4274 = ~n4160 & n4273;
  assign n4275 = ~n4159 & n4274;
  assign n4276 = ~n4153 & n4275;
  assign n4277 = ~n4165 & n4273;
  assign n4278 = pi15 & ~n4277;
  assign n4279 = ~n4276 & n4278;
  assign n4280 = ~n4272 & n4279;
  assign n4281 = ~n4114 & n4151;
  assign n4282 = ~n4114 & ~n4134;
  assign n4283 = ~n4150 & ~n4282;
  assign n4284 = ~n4281 & ~n4283;
  assign n4285 = n4182 & ~n4284;
  assign n4286 = n3979 & ~n4014;
  assign n4287 = ~n4012 & n4286;
  assign n4288 = ~n4037 & ~n4146;
  assign n4289 = ~n4287 & ~n4288;
  assign n4290 = ~n4182 & ~n4289;
  assign n4291 = ~pi13 & ~n4290;
  assign n4292 = ~n4285 & n4291;
  assign n4293 = ~n4280 & n4292;
  assign n4294 = ~n4182 & n4242;
  assign n4295 = ~n4178 & n4252;
  assign n4296 = ~n4181 & n4295;
  assign n4297 = ~n4294 & ~n4296;
  assign n4298 = n4237 & ~n4297;
  assign n4299 = ~n4276 & ~n4277;
  assign n4300 = ~pi15 & ~n4299;
  assign n4301 = ~n4178 & n4231;
  assign n4302 = ~n4181 & n4301;
  assign n4303 = ~n4300 & ~n4302;
  assign n4304 = n740 & ~n4153;
  assign n4305 = ~n4181 & n4304;
  assign n4306 = ~n4269 & n4305;
  assign n4307 = ~n4182 & n4218;
  assign n4308 = ~n4306 & ~n4307;
  assign n4309 = ~pi11 & ~n4130;
  assign n4310 = ~n4132 & n4309;
  assign n4311 = ~n4182 & n4310;
  assign n4312 = ~n4103 & ~n4107;
  assign n4313 = ~n4134 & n4312;
  assign n4314 = ~n4096 & ~n4109;
  assign n4315 = ~n4095 & n4314;
  assign n4316 = ~n4089 & n4315;
  assign n4317 = n4313 & ~n4316;
  assign n4318 = ~n4313 & n4316;
  assign n4319 = ~pi11 & ~n4178;
  assign n4320 = ~n4318 & n4319;
  assign n4321 = ~n4317 & n4320;
  assign n4322 = ~n4181 & n4321;
  assign n4323 = ~n4311 & ~n4322;
  assign n4324 = n4308 & n4323;
  assign n4325 = n4303 & n4324;
  assign n4326 = ~n4298 & n4325;
  assign n4327 = ~n4293 & n4326;
  assign n4328 = ~n4260 & n4327;
  assign n4329 = ~n4300 & ~n4306;
  assign n4330 = pi11 & ~n4133;
  assign n4331 = ~n4182 & n4330;
  assign n4332 = ~n4317 & ~n4318;
  assign n4333 = pi11 & ~n4178;
  assign n4334 = ~n4181 & n4333;
  assign n4335 = ~n4332 & n4334;
  assign n4336 = ~n4331 & ~n4335;
  assign n4337 = n4329 & n4336;
  assign n4338 = ~n4280 & n4337;
  assign n4339 = ~n4285 & ~n4290;
  assign n4340 = pi13 & ~n4339;
  assign n4341 = ~n4292 & ~n4340;
  assign n4342 = n4338 & n4341;
  assign n4343 = ~n4293 & n4329;
  assign n4344 = ~n4342 & n4343;
  assign n4345 = ~n4159 & ~n4160;
  assign n4346 = ~n4153 & n4345;
  assign n4347 = n4023 & ~n4178;
  assign n4348 = ~n4181 & n4347;
  assign n4349 = ~n4346 & n4348;
  assign n4350 = ~n4021 & ~n4182;
  assign n4351 = ~pi17 & ~n4350;
  assign n4352 = ~n4349 & n4351;
  assign n4353 = ~n4349 & ~n4350;
  assign n4354 = pi17 & ~n4353;
  assign n4355 = ~n4352 & ~n4354;
  assign n4356 = n180 & ~n4355;
  assign n4357 = ~n4344 & n4356;
  assign n4358 = ~n4328 & n4357;
  assign n4359 = n119 & ~n4353;
  assign n4360 = ~n4358 & ~n4359;
  assign n4361 = pi03 & ~n4173;
  assign n4362 = ~n4203 & ~n4361;
  assign n4363 = ~n70 & ~n4362;
  assign n4364 = n70 & ~n4203;
  assign n4365 = ~n4361 & n4364;
  assign n4366 = ~n4363 & ~n4365;
  assign n4367 = ~n4360 & n4366;
  assign n4368 = ~n4173 & ~n4359;
  assign n4369 = ~n4358 & n4368;
  assign n4370 = ~n4367 & ~n4369;
  assign n4371 = pi05 & ~n4370;
  assign n4372 = pi14 & ~n4359;
  assign n4373 = n70 & n74;
  assign n4374 = n69 & n4373;
  assign n4375 = ~n4353 & n4374;
  assign n4376 = ~n1169 & ~n4375;
  assign n4377 = ~n4372 & n4376;
  assign n4378 = ~n1165 & ~n4377;
  assign n4379 = ~n4358 & n4378;
  assign n4380 = ~n1162 & ~n1169;
  assign n4381 = ~n4375 & n4380;
  assign n4382 = ~n4372 & n4381;
  assign n4383 = ~n4358 & n4382;
  assign n4384 = n1178 & ~n4355;
  assign n4385 = ~n4344 & n4384;
  assign n4386 = ~n4328 & n4385;
  assign n4387 = n1172 & ~n4355;
  assign n4388 = ~n4344 & n4387;
  assign n4389 = ~n4328 & n4388;
  assign n4390 = ~n4386 & ~n4389;
  assign n4391 = ~n4383 & n4390;
  assign n4392 = ~n4379 & n4391;
  assign n4393 = ~pi05 & ~n70;
  assign n4394 = ~n4362 & n4393;
  assign n4395 = ~pi14 & n91;
  assign n4396 = ~n4203 & n4395;
  assign n4397 = ~n4361 & n4396;
  assign n4398 = ~n4394 & ~n4397;
  assign n4399 = n4356 & ~n4398;
  assign n4400 = ~n4344 & n4399;
  assign n4401 = ~n4328 & n4400;
  assign n4402 = n1195 & ~n4355;
  assign n4403 = ~n4344 & n4402;
  assign n4404 = ~n4328 & n4403;
  assign n4405 = n1201 & ~n4353;
  assign n4406 = ~n4366 & n4405;
  assign n4407 = ~n4404 & ~n4406;
  assign n4408 = ~n4401 & n4407;
  assign n4409 = ~pi03 & ~n4377;
  assign n4410 = ~n4358 & n4409;
  assign n4411 = ~pi05 & ~n4168;
  assign n4412 = ~n4171 & n4411;
  assign n4413 = ~n4164 & n4412;
  assign n4414 = ~n4359 & n4413;
  assign n4415 = ~n4358 & n4414;
  assign n4416 = ~n4410 & ~n4415;
  assign n4417 = n4408 & n4416;
  assign n4418 = ~n4392 & n4417;
  assign n4419 = ~n4177 & ~n4203;
  assign n4420 = ~n4174 & n4419;
  assign n4421 = ~n4182 & n4186;
  assign n4422 = ~n4178 & ~n4196;
  assign n4423 = ~n4194 & n4422;
  assign n4424 = ~n4181 & n4423;
  assign n4425 = ~n4421 & ~n4424;
  assign n4426 = ~pi05 & ~n4425;
  assign n4427 = pi05 & ~n4424;
  assign n4428 = ~n4421 & n4427;
  assign n4429 = ~n4426 & ~n4428;
  assign n4430 = ~n4420 & ~n4429;
  assign n4431 = n4420 & ~n4428;
  assign n4432 = ~n4426 & n4431;
  assign n4433 = ~pi07 & ~n4432;
  assign n4434 = ~n4430 & n4433;
  assign n4435 = ~n4430 & ~n4432;
  assign n4436 = pi07 & ~n4435;
  assign n4437 = ~n4434 & ~n4436;
  assign n4438 = ~n4360 & ~n4437;
  assign n4439 = ~n4206 & n4213;
  assign n4440 = ~n4257 & ~n4439;
  assign n4441 = n4213 & n4257;
  assign n4442 = ~n4206 & n4441;
  assign n4443 = ~pi09 & ~n4442;
  assign n4444 = ~n4440 & n4443;
  assign n4445 = ~n4440 & ~n4442;
  assign n4446 = pi09 & ~n4445;
  assign n4447 = ~n4444 & ~n4446;
  assign n4448 = ~n4360 & ~n4447;
  assign n4449 = ~n4182 & ~n4243;
  assign n4450 = ~n4178 & ~n4253;
  assign n4451 = ~n4181 & n4450;
  assign n4452 = ~pi09 & ~n4451;
  assign n4453 = ~n4449 & n4452;
  assign n4454 = ~n4449 & ~n4451;
  assign n4455 = pi09 & ~n4454;
  assign n4456 = ~n4453 & ~n4455;
  assign n4457 = ~n4359 & ~n4456;
  assign n4458 = ~n4358 & n4457;
  assign n4459 = ~pi07 & ~n4424;
  assign n4460 = ~n4421 & n4459;
  assign n4461 = pi07 & ~n4425;
  assign n4462 = ~n4460 & ~n4461;
  assign n4463 = ~n4359 & ~n4462;
  assign n4464 = ~n4358 & n4463;
  assign n4465 = ~n4458 & ~n4464;
  assign n4466 = ~n4448 & n4465;
  assign n4467 = ~n4438 & n4466;
  assign n4468 = ~n4418 & n4467;
  assign n4469 = ~n4371 & n4468;
  assign n4470 = ~n4360 & n4434;
  assign n4471 = ~n4359 & n4460;
  assign n4472 = ~n4358 & n4471;
  assign n4473 = ~n4470 & ~n4472;
  assign n4474 = ~n4448 & ~n4458;
  assign n4475 = ~n4473 & n4474;
  assign n4476 = ~n4237 & n4297;
  assign n4477 = ~n4439 & n4476;
  assign n4478 = ~n4257 & n4476;
  assign n4479 = ~pi11 & ~n4298;
  assign n4480 = ~n4478 & n4479;
  assign n4481 = ~n4260 & n4480;
  assign n4482 = ~n4477 & n4481;
  assign n4483 = ~n4360 & n4482;
  assign n4484 = ~n4360 & n4444;
  assign n4485 = ~n4359 & n4453;
  assign n4486 = ~n4358 & n4485;
  assign n4487 = ~n4182 & ~n4219;
  assign n4488 = ~n4178 & ~n4233;
  assign n4489 = ~n4181 & n4488;
  assign n4490 = ~pi11 & ~n4489;
  assign n4491 = ~n4487 & n4490;
  assign n4492 = ~n4359 & n4491;
  assign n4493 = ~n4358 & n4492;
  assign n4494 = ~n4486 & ~n4493;
  assign n4495 = ~n4484 & n4494;
  assign n4496 = ~n4483 & n4495;
  assign n4497 = ~n4475 & n4496;
  assign n4498 = ~n4469 & n4497;
  assign n4499 = ~n4344 & n4355;
  assign n4500 = ~n4328 & n4499;
  assign n4501 = ~n4360 & n4500;
  assign n4502 = ~n4353 & ~n4359;
  assign n4503 = ~n4358 & n4502;
  assign n4504 = ~pi19 & ~n4503;
  assign n4505 = ~n4501 & n4504;
  assign n4506 = ~n4501 & ~n4503;
  assign n4507 = pi19 & ~n4506;
  assign n4508 = ~n4505 & ~n4507;
  assign n4509 = n4323 & n4336;
  assign n4510 = ~n4302 & ~n4307;
  assign n4511 = ~n4298 & n4510;
  assign n4512 = ~n4260 & n4511;
  assign n4513 = n4509 & ~n4512;
  assign n4514 = ~n4509 & n4511;
  assign n4515 = ~n4260 & n4514;
  assign n4516 = ~pi13 & ~n4515;
  assign n4517 = ~n4513 & n4516;
  assign n4518 = ~n4513 & ~n4515;
  assign n4519 = pi13 & ~n4518;
  assign n4520 = ~n4517 & ~n4519;
  assign n4521 = ~n4360 & ~n4520;
  assign n4522 = ~pi15 & ~n4290;
  assign n4523 = ~n4285 & n4522;
  assign n4524 = ~n4359 & n4523;
  assign n4525 = ~n4358 & n4524;
  assign n4526 = n1718 & ~n4525;
  assign n4527 = pi15 & ~n4339;
  assign n4528 = ~n4359 & n4527;
  assign n4529 = ~n4358 & n4528;
  assign n4530 = n4182 & ~n4332;
  assign n4531 = ~n4133 & ~n4182;
  assign n4532 = ~pi13 & ~n4531;
  assign n4533 = ~n4530 & n4532;
  assign n4534 = ~n4530 & ~n4531;
  assign n4535 = pi13 & ~n4534;
  assign n4536 = ~n4533 & ~n4535;
  assign n4537 = ~n4359 & ~n4536;
  assign n4538 = ~n4358 & n4537;
  assign n4539 = ~n4529 & ~n4538;
  assign n4540 = n4526 & n4539;
  assign n4541 = n4257 & n4336;
  assign n4542 = n4213 & n4237;
  assign n4543 = n4541 & n4542;
  assign n4544 = ~n4206 & n4543;
  assign n4545 = n4323 & n4510;
  assign n4546 = ~n4298 & n4545;
  assign n4547 = n4336 & ~n4546;
  assign n4548 = ~n4544 & ~n4547;
  assign n4549 = n4341 & ~n4548;
  assign n4550 = ~n4341 & ~n4544;
  assign n4551 = ~n4547 & n4550;
  assign n4552 = ~pi15 & ~n4551;
  assign n4553 = ~n4549 & n4552;
  assign n4554 = ~n4360 & n4553;
  assign n4555 = ~n4549 & ~n4551;
  assign n4556 = pi15 & ~n4555;
  assign n4557 = ~n4360 & n4556;
  assign n4558 = ~n4554 & ~n4557;
  assign n4559 = n4540 & n4558;
  assign n4560 = ~n4521 & n4559;
  assign n4561 = ~n4487 & ~n4489;
  assign n4562 = ~n4359 & ~n4561;
  assign n4563 = ~n4358 & n4562;
  assign n4564 = ~n4298 & ~n4478;
  assign n4565 = ~n4260 & n4564;
  assign n4566 = ~n4477 & n4565;
  assign n4567 = ~n4360 & ~n4566;
  assign n4568 = ~n4563 & ~n4567;
  assign n4569 = pi11 & ~n4568;
  assign n4570 = ~n4280 & n4329;
  assign n4571 = ~n4292 & ~n4570;
  assign n4572 = n4292 & n4570;
  assign n4573 = ~n4571 & ~n4572;
  assign n4574 = ~n4549 & n4573;
  assign n4575 = n4341 & ~n4570;
  assign n4576 = ~n4548 & n4575;
  assign n4577 = ~n4574 & ~n4576;
  assign n4578 = ~n4360 & n4577;
  assign n4579 = ~n4272 & n4299;
  assign n4580 = ~n4359 & n4579;
  assign n4581 = ~n4358 & n4580;
  assign n4582 = ~n4578 & ~n4581;
  assign n4583 = pi17 & ~n4582;
  assign n4584 = ~n4569 & ~n4583;
  assign n4585 = n4560 & n4584;
  assign n4586 = ~n4508 & n4585;
  assign n4587 = ~n4498 & n4586;
  assign n4588 = n180 & ~n4506;
  assign n4589 = ~n4360 & n4517;
  assign n4590 = ~n4359 & n4533;
  assign n4591 = ~n4358 & n4590;
  assign n4592 = ~n4589 & ~n4591;
  assign n4593 = ~n4529 & ~n4557;
  assign n4594 = ~n4592 & n4593;
  assign n4595 = ~pi17 & ~n4581;
  assign n4596 = ~n4578 & n4595;
  assign n4597 = ~n4525 & ~n4554;
  assign n4598 = ~n4596 & n4597;
  assign n4599 = ~n4594 & n4598;
  assign n4600 = n1718 & ~n4583;
  assign n4601 = ~n4508 & n4600;
  assign n4602 = ~n4599 & n4601;
  assign n4603 = ~n4588 & ~n4602;
  assign n4604 = ~n4587 & n4603;
  assign n4605 = ~n4358 & n4377;
  assign n4606 = n1532 & ~n4355;
  assign n4607 = ~n4344 & n4606;
  assign n4608 = ~n4328 & n4607;
  assign n4609 = n1537 & ~n4608;
  assign n4610 = ~n4605 & n4609;
  assign n4611 = ~n4605 & ~n4608;
  assign n4612 = ~n1537 & ~n4611;
  assign n4613 = ~n4610 & ~n4612;
  assign n4614 = ~pi05 & ~n4613;
  assign n4615 = pi05 & ~n4610;
  assign n4616 = ~n4612 & n4615;
  assign n4617 = ~n4614 & ~n4616;
  assign n4618 = ~n4604 & ~n4617;
  assign n4619 = n1549 & ~n4604;
  assign n4620 = ~pi05 & ~n4369;
  assign n4621 = ~n4367 & n4620;
  assign n4622 = ~n4371 & ~n4621;
  assign n4623 = ~n4404 & ~n4410;
  assign n4624 = ~n4392 & n4623;
  assign n4625 = n4622 & ~n4624;
  assign n4626 = ~n4622 & n4624;
  assign n4627 = ~pi07 & ~n4626;
  assign n4628 = ~n4625 & n4627;
  assign n4629 = ~n4625 & ~n4626;
  assign n4630 = pi07 & ~n4629;
  assign n4631 = ~n4628 & ~n4630;
  assign n4632 = ~n4604 & ~n4631;
  assign n4633 = ~n4619 & ~n4632;
  assign n4634 = ~n4618 & n4633;
  assign n4635 = pi03 & ~n4588;
  assign n4636 = ~n4602 & n4635;
  assign n4637 = ~n4587 & n4636;
  assign n4638 = n1571 & ~n4637;
  assign n4639 = n1574 & ~n4588;
  assign n4640 = ~n4602 & n4639;
  assign n4641 = ~n4587 & n4640;
  assign n4642 = ~n1573 & ~n4641;
  assign n4643 = ~n4638 & n4642;
  assign n4644 = ~pi05 & ~n4608;
  assign n4645 = ~n4605 & n4644;
  assign n4646 = pi05 & ~n4611;
  assign n4647 = ~n4645 & ~n4646;
  assign n4648 = ~n4588 & ~n4647;
  assign n4649 = ~n4602 & n4648;
  assign n4650 = ~n4587 & n4649;
  assign n4651 = ~pi12 & n1548;
  assign n4652 = ~n4588 & n4651;
  assign n4653 = ~n4602 & n4652;
  assign n4654 = ~n4587 & n4653;
  assign n4655 = ~pi07 & ~n4369;
  assign n4656 = ~n4367 & n4655;
  assign n4657 = pi07 & ~n4370;
  assign n4658 = ~n4656 & ~n4657;
  assign n4659 = ~n4588 & ~n4658;
  assign n4660 = ~n4602 & n4659;
  assign n4661 = ~n4587 & n4660;
  assign n4662 = ~n4654 & ~n4661;
  assign n4663 = ~n4650 & n4662;
  assign n4664 = ~n4643 & n4663;
  assign n4665 = n4634 & n4664;
  assign n4666 = ~n4588 & n4645;
  assign n4667 = ~n4602 & n4666;
  assign n4668 = ~n4587 & n4667;
  assign n4669 = ~n4604 & n4614;
  assign n4670 = ~n4668 & ~n4669;
  assign n4671 = ~n4632 & ~n4661;
  assign n4672 = ~n4670 & n4671;
  assign n4673 = ~n4604 & n4628;
  assign n4674 = ~n4438 & ~n4464;
  assign n4675 = ~n4418 & n4674;
  assign n4676 = ~n4371 & n4675;
  assign n4677 = ~n4371 & ~n4418;
  assign n4678 = ~n4674 & ~n4677;
  assign n4679 = ~pi09 & ~n4678;
  assign n4680 = ~n4676 & n4679;
  assign n4681 = ~n4604 & n4680;
  assign n4682 = ~n4360 & ~n4435;
  assign n4683 = ~n4359 & ~n4425;
  assign n4684 = ~n4358 & n4683;
  assign n4685 = ~pi09 & ~n4684;
  assign n4686 = ~n4682 & n4685;
  assign n4687 = ~n4588 & n4686;
  assign n4688 = ~n4602 & n4687;
  assign n4689 = ~n4587 & n4688;
  assign n4690 = ~n4588 & n4656;
  assign n4691 = ~n4602 & n4690;
  assign n4692 = ~n4587 & n4691;
  assign n4693 = ~n4689 & ~n4692;
  assign n4694 = ~n4681 & n4693;
  assign n4695 = ~n4673 & n4694;
  assign n4696 = ~n4672 & n4695;
  assign n4697 = ~n4665 & n4696;
  assign n4698 = ~n4676 & ~n4678;
  assign n4699 = ~n4604 & ~n4698;
  assign n4700 = ~n4682 & ~n4684;
  assign n4701 = ~n4588 & ~n4700;
  assign n4702 = ~n4602 & n4701;
  assign n4703 = ~n4587 & n4702;
  assign n4704 = ~n4699 & ~n4703;
  assign n4705 = pi09 & ~n4704;
  assign n4706 = pi11 & ~n4474;
  assign n4707 = ~pi11 & ~n4458;
  assign n4708 = ~n4448 & n4707;
  assign n4709 = n4473 & ~n4708;
  assign n4710 = ~n4706 & n4709;
  assign n4711 = ~n4676 & n4710;
  assign n4712 = n4473 & ~n4676;
  assign n4713 = ~n4706 & ~n4708;
  assign n4714 = ~n4712 & ~n4713;
  assign n4715 = ~n4711 & ~n4714;
  assign n4716 = ~n4604 & n4715;
  assign n4717 = ~n4484 & ~n4486;
  assign n4718 = ~n4475 & n4717;
  assign n4719 = ~n4469 & n4718;
  assign n4720 = ~pi13 & ~n4493;
  assign n4721 = ~n4483 & n4720;
  assign n4722 = ~n4569 & n4721;
  assign n4723 = ~n4483 & ~n4493;
  assign n4724 = ~n4569 & n4723;
  assign n4725 = pi13 & ~n4724;
  assign n4726 = ~n4722 & ~n4725;
  assign n4727 = ~n4719 & ~n4726;
  assign n4728 = n4718 & ~n4722;
  assign n4729 = ~n4469 & n4728;
  assign n4730 = ~n4725 & n4729;
  assign n4731 = ~n4727 & ~n4730;
  assign n4732 = ~n4604 & n4731;
  assign n4733 = ~pi13 & ~n4563;
  assign n4734 = ~n4567 & n4733;
  assign n4735 = pi13 & ~n4568;
  assign n4736 = ~n4734 & ~n4735;
  assign n4737 = ~n4588 & ~n4736;
  assign n4738 = ~n4602 & n4737;
  assign n4739 = ~n4587 & n4738;
  assign n4740 = ~n4360 & ~n4445;
  assign n4741 = ~n4359 & ~n4454;
  assign n4742 = ~n4358 & n4741;
  assign n4743 = ~pi11 & ~n4742;
  assign n4744 = ~n4740 & n4743;
  assign n4745 = ~n4740 & ~n4742;
  assign n4746 = pi11 & ~n4745;
  assign n4747 = ~n4744 & ~n4746;
  assign n4748 = ~n4588 & ~n4747;
  assign n4749 = ~n4602 & n4748;
  assign n4750 = ~n4587 & n4749;
  assign n4751 = ~n4739 & ~n4750;
  assign n4752 = ~n4732 & n4751;
  assign n4753 = ~n4716 & n4752;
  assign n4754 = ~n4705 & n4753;
  assign n4755 = ~n4697 & n4754;
  assign n4756 = ~pi17 & ~n4604;
  assign n4757 = ~n4525 & ~n4529;
  assign n4758 = ~n4538 & n4757;
  assign n4759 = n4558 & n4758;
  assign n4760 = ~n4521 & n4759;
  assign n4761 = ~n4569 & ~n4594;
  assign n4762 = n4760 & n4761;
  assign n4763 = ~n4498 & n4762;
  assign n4764 = ~pi17 & ~n4582;
  assign n4765 = pi17 & ~n4581;
  assign n4766 = ~n4578 & n4765;
  assign n4767 = n4597 & ~n4766;
  assign n4768 = ~n4594 & n4767;
  assign n4769 = ~n4764 & n4768;
  assign n4770 = ~n4594 & n4597;
  assign n4771 = ~n4764 & ~n4766;
  assign n4772 = ~n4770 & ~n4771;
  assign n4773 = ~n4769 & ~n4772;
  assign n4774 = ~n4763 & ~n4773;
  assign n4775 = n4762 & ~n4769;
  assign n4776 = ~n4772 & n4775;
  assign n4777 = ~n4498 & n4776;
  assign n4778 = ~n4774 & ~n4777;
  assign n4779 = n4756 & n4778;
  assign n4780 = n4582 & ~n4588;
  assign n4781 = ~n4602 & n4780;
  assign n4782 = ~n4587 & n4781;
  assign n4783 = pi19 & ~n4782;
  assign n4784 = ~pi17 & ~n4783;
  assign n4785 = ~n4779 & ~n4784;
  assign n4786 = ~n4569 & n4760;
  assign n4787 = ~n4498 & n4786;
  assign n4788 = n4496 & n4592;
  assign n4789 = ~n4554 & n4757;
  assign n4790 = ~n4557 & n4789;
  assign n4791 = ~n4475 & ~n4790;
  assign n4792 = n4788 & n4791;
  assign n4793 = ~n4469 & n4792;
  assign n4794 = ~n4592 & n4790;
  assign n4795 = ~n4521 & ~n4538;
  assign n4796 = ~n4569 & n4795;
  assign n4797 = n4592 & ~n4790;
  assign n4798 = ~n4796 & n4797;
  assign n4799 = ~n4794 & ~n4798;
  assign n4800 = ~n4793 & n4799;
  assign n4801 = ~n4787 & n4800;
  assign n4802 = ~n4604 & ~n4801;
  assign n4803 = ~n4339 & ~n4359;
  assign n4804 = ~n4358 & n4803;
  assign n4805 = ~n4360 & ~n4555;
  assign n4806 = ~n4804 & ~n4805;
  assign n4807 = ~n4588 & ~n4806;
  assign n4808 = ~n4602 & n4807;
  assign n4809 = ~n4587 & n4808;
  assign n4810 = ~n4802 & ~n4809;
  assign n4811 = ~n4785 & n4810;
  assign n4812 = ~n4604 & ~n4774;
  assign n4813 = ~n4777 & n4812;
  assign n4814 = ~n4782 & ~n4813;
  assign n4815 = ~pi19 & ~n4814;
  assign n4816 = ~n4588 & ~n4745;
  assign n4817 = ~n4602 & n4816;
  assign n4818 = ~n4587 & n4817;
  assign n4819 = ~pi11 & ~n4739;
  assign n4820 = ~n4818 & n4819;
  assign n4821 = n4474 & ~n4712;
  assign n4822 = n4473 & ~n4474;
  assign n4823 = ~n4676 & n4822;
  assign n4824 = ~n4821 & ~n4823;
  assign n4825 = ~n4604 & ~n4824;
  assign n4826 = ~n4732 & ~n4825;
  assign n4827 = n4820 & n4826;
  assign n4828 = ~n4719 & n4724;
  assign n4829 = n4718 & ~n4724;
  assign n4830 = ~n4469 & n4829;
  assign n4831 = ~n4828 & ~n4830;
  assign n4832 = ~n4604 & ~n4831;
  assign n4833 = ~n4568 & ~n4588;
  assign n4834 = ~n4602 & n4833;
  assign n4835 = ~n4587 & n4834;
  assign n4836 = ~pi13 & ~n4835;
  assign n4837 = ~n4832 & n4836;
  assign n4838 = ~n4497 & ~n4569;
  assign n4839 = ~n4371 & ~n4569;
  assign n4840 = n4468 & n4839;
  assign n4841 = ~n4838 & ~n4840;
  assign n4842 = n4795 & ~n4841;
  assign n4843 = ~n4795 & ~n4838;
  assign n4844 = ~n4840 & n4843;
  assign n4845 = ~n4842 & ~n4844;
  assign n4846 = ~n4604 & ~n4845;
  assign n4847 = ~n4359 & ~n4534;
  assign n4848 = ~n4358 & n4847;
  assign n4849 = ~n4360 & ~n4518;
  assign n4850 = ~n4848 & ~n4849;
  assign n4851 = ~n4588 & ~n4850;
  assign n4852 = ~n4602 & n4851;
  assign n4853 = ~n4587 & n4852;
  assign n4854 = ~pi15 & ~n4853;
  assign n4855 = ~n4846 & n4854;
  assign n4856 = ~n4837 & ~n4855;
  assign n4857 = ~n4827 & n4856;
  assign n4858 = ~n4815 & n4857;
  assign n4859 = ~n4811 & n4858;
  assign n4860 = ~n4755 & n4859;
  assign n4861 = ~n4846 & ~n4853;
  assign n4862 = pi15 & ~n4861;
  assign n4863 = pi17 & ~n4604;
  assign n4864 = ~n4801 & n4863;
  assign n4865 = ~pi17 & ~n4794;
  assign n4866 = ~n4798 & n4865;
  assign n4867 = ~n4793 & n4866;
  assign n4868 = ~n4787 & n4867;
  assign n4869 = ~n4604 & n4868;
  assign n4870 = ~pi17 & ~n4804;
  assign n4871 = ~n4805 & n4870;
  assign n4872 = pi17 & ~n4806;
  assign n4873 = ~n4871 & ~n4872;
  assign n4874 = ~n4588 & ~n4873;
  assign n4875 = ~n4602 & n4874;
  assign n4876 = ~n4587 & n4875;
  assign n4877 = ~n4869 & ~n4876;
  assign n4878 = ~n4864 & n4877;
  assign n4879 = ~n4862 & n4878;
  assign n4880 = ~n4777 & ~n4782;
  assign n4881 = n4812 & n4880;
  assign n4882 = ~pi19 & ~n4581;
  assign n4883 = ~n4578 & n4882;
  assign n4884 = ~n4588 & n4883;
  assign n4885 = ~n4602 & n4884;
  assign n4886 = ~n4587 & n4885;
  assign n4887 = ~n4783 & ~n4886;
  assign n4888 = ~n4881 & ~n4887;
  assign n4889 = n4881 & n4887;
  assign n4890 = ~n4888 & ~n4889;
  assign n4891 = n4879 & n4890;
  assign n4892 = ~n4811 & ~n4815;
  assign n4893 = ~n4891 & n4892;
  assign n4894 = n4599 & ~n4787;
  assign n4895 = n4508 & ~n4583;
  assign n4896 = ~n4894 & n4895;
  assign n4897 = ~n4604 & n4896;
  assign n4898 = ~n4506 & ~n4588;
  assign n4899 = ~n4602 & n4898;
  assign n4900 = ~n4587 & n4899;
  assign n4901 = ~pi21 & ~n4900;
  assign n4902 = ~n4897 & n4901;
  assign n4903 = ~n4897 & ~n4900;
  assign n4904 = pi21 & ~n4903;
  assign n4905 = ~n4902 & ~n4904;
  assign n4906 = n1745 & ~n4905;
  assign n4907 = ~n4893 & n4906;
  assign n4908 = ~n4860 & n4907;
  assign n4909 = n1718 & ~n4903;
  assign n4910 = ~n4903 & ~n4909;
  assign n4911 = ~n4908 & n4910;
  assign n4912 = ~n4893 & n4909;
  assign n4913 = ~n4860 & n4912;
  assign n4914 = ~pi23 & ~n4913;
  assign n4915 = ~n4911 & n4914;
  assign n4916 = ~n4911 & ~n4913;
  assign n4917 = pi23 & ~n4916;
  assign n4918 = ~n4915 & ~n4917;
  assign n4919 = n69 & ~n4918;
  assign n4920 = n1745 & ~n4916;
  assign n4921 = ~n4919 & ~n4920;
  assign n4922 = ~pi13 & ~n4818;
  assign n4923 = ~n4825 & n4922;
  assign n4924 = ~n4909 & n4923;
  assign n4925 = ~n4908 & n4924;
  assign n4926 = ~n4908 & ~n4909;
  assign n4927 = ~n4716 & ~n4750;
  assign n4928 = ~n4697 & ~n4705;
  assign n4929 = ~n4927 & ~n4928;
  assign n4930 = ~n4705 & n4927;
  assign n4931 = ~n4697 & n4930;
  assign n4932 = ~pi13 & ~n4931;
  assign n4933 = ~n4929 & n4932;
  assign n4934 = ~n4926 & n4933;
  assign n4935 = ~n4925 & ~n4934;
  assign n4936 = ~pi15 & ~n4835;
  assign n4937 = ~n4832 & n4936;
  assign n4938 = ~n4832 & ~n4835;
  assign n4939 = pi15 & ~n4938;
  assign n4940 = ~n4937 & ~n4939;
  assign n4941 = ~n4909 & ~n4940;
  assign n4942 = ~n4908 & n4941;
  assign n4943 = ~n4732 & ~n4739;
  assign n4944 = ~pi11 & ~n4818;
  assign n4945 = ~n4825 & n4944;
  assign n4946 = ~n4943 & ~n4945;
  assign n4947 = ~n4827 & ~n4946;
  assign n4948 = ~n4827 & n4930;
  assign n4949 = ~n4697 & n4948;
  assign n4950 = ~n4947 & ~n4949;
  assign n4951 = ~pi15 & ~n4755;
  assign n4952 = ~n4950 & n4951;
  assign n4953 = ~n4755 & ~n4950;
  assign n4954 = pi15 & ~n4953;
  assign n4955 = ~n4952 & ~n4954;
  assign n4956 = ~n4926 & ~n4955;
  assign n4957 = ~n4942 & ~n4956;
  assign n4958 = ~n4935 & n4957;
  assign n4959 = ~n4926 & ~n4953;
  assign n4960 = ~n4909 & ~n4938;
  assign n4961 = ~n4908 & n4960;
  assign n4962 = ~pi15 & ~n4961;
  assign n4963 = ~n4959 & n4962;
  assign n4964 = ~n4855 & ~n4862;
  assign n4965 = ~n4827 & ~n4837;
  assign n4966 = ~n4964 & n4965;
  assign n4967 = ~n4755 & n4966;
  assign n4968 = ~n4755 & n4965;
  assign n4969 = n4964 & ~n4968;
  assign n4970 = ~n4967 & ~n4969;
  assign n4971 = ~n4926 & ~n4970;
  assign n4972 = ~n4861 & ~n4909;
  assign n4973 = ~n4908 & n4972;
  assign n4974 = ~pi17 & ~n4973;
  assign n4975 = ~n4971 & n4974;
  assign n4976 = ~n4963 & ~n4975;
  assign n4977 = ~n4958 & n4976;
  assign n4978 = ~pi17 & ~n4809;
  assign n4979 = ~n4802 & n4978;
  assign n4980 = ~n4879 & ~n4979;
  assign n4981 = n4856 & ~n4979;
  assign n4982 = ~n4827 & n4981;
  assign n4983 = ~n4755 & n4982;
  assign n4984 = ~n4980 & ~n4983;
  assign n4985 = ~n4890 & ~n4984;
  assign n4986 = n4890 & ~n4980;
  assign n4987 = ~n4983 & n4986;
  assign n4988 = pi21 & ~n4987;
  assign n4989 = ~n4926 & n4988;
  assign n4990 = ~n4985 & n4989;
  assign n4991 = ~pi21 & ~n4814;
  assign n4992 = pi21 & ~n4782;
  assign n4993 = ~n4813 & n4992;
  assign n4994 = ~n4909 & ~n4993;
  assign n4995 = ~n4991 & n4994;
  assign n4996 = ~n4908 & n4995;
  assign n4997 = ~n4985 & ~n4987;
  assign n4998 = ~n4860 & ~n4893;
  assign n4999 = n4903 & ~n4998;
  assign n5000 = n1718 & ~n4999;
  assign n5001 = ~n4997 & n5000;
  assign n5002 = ~n4996 & ~n5001;
  assign n5003 = ~n4990 & n5002;
  assign n5004 = n4857 & ~n4862;
  assign n5005 = ~n4755 & n5004;
  assign n5006 = n4862 & ~n4878;
  assign n5007 = ~n4879 & ~n5006;
  assign n5008 = ~n5005 & ~n5007;
  assign n5009 = n5004 & n5007;
  assign n5010 = ~n4755 & n5009;
  assign n5011 = ~pi19 & ~n5010;
  assign n5012 = ~n5008 & n5011;
  assign n5013 = ~n5008 & ~n5010;
  assign n5014 = pi19 & ~n5013;
  assign n5015 = ~n5012 & ~n5014;
  assign n5016 = ~n4926 & ~n5015;
  assign n5017 = ~n4971 & ~n4973;
  assign n5018 = pi17 & ~n5017;
  assign n5019 = ~pi19 & ~n4809;
  assign n5020 = ~n4802 & n5019;
  assign n5021 = pi19 & ~n4810;
  assign n5022 = ~n5020 & ~n5021;
  assign n5023 = ~n4909 & ~n5022;
  assign n5024 = ~n4908 & n5023;
  assign n5025 = ~n5018 & ~n5024;
  assign n5026 = ~n5016 & n5025;
  assign n5027 = ~n5003 & n5026;
  assign n5028 = ~n4977 & n5027;
  assign n5029 = pi10 & ~n4909;
  assign n5030 = n73 & n1548;
  assign n5031 = n69 & n5030;
  assign n5032 = ~n4903 & n5031;
  assign n5033 = ~n1774 & ~n5032;
  assign n5034 = ~n5029 & n5033;
  assign n5035 = ~n1770 & ~n5034;
  assign n5036 = ~n4908 & n5035;
  assign n5037 = ~n1767 & ~n1774;
  assign n5038 = ~n5032 & n5037;
  assign n5039 = ~n5029 & n5038;
  assign n5040 = ~n4908 & n5039;
  assign n5041 = n98 & ~n1548;
  assign n5042 = ~n1774 & n5041;
  assign n5043 = n67 & ~n1767;
  assign n5044 = n5042 & n5043;
  assign n5045 = ~n4905 & n5044;
  assign n5046 = ~n4893 & n5045;
  assign n5047 = ~n4860 & n5046;
  assign n5048 = n1745 & n1776;
  assign n5049 = ~n4905 & n5048;
  assign n5050 = ~n4893 & n5049;
  assign n5051 = ~n4860 & n5050;
  assign n5052 = ~n5047 & ~n5051;
  assign n5053 = ~n5040 & n5052;
  assign n5054 = ~n5036 & n5053;
  assign n5055 = ~pi03 & ~n5034;
  assign n5056 = ~n4908 & n5055;
  assign n5057 = ~pi23 & ~pi29;
  assign n5058 = n68 & n5057;
  assign n5059 = n3335 & n5058;
  assign n5060 = ~n1775 & n5059;
  assign n5061 = ~n4905 & n5060;
  assign n5062 = ~n4893 & n5061;
  assign n5063 = ~n4860 & n5062;
  assign n5064 = pi01 & ~n4604;
  assign n5065 = pi12 & ~n5064;
  assign n5066 = n1161 & ~n4604;
  assign n5067 = ~n5065 & ~n5066;
  assign n5068 = ~pi03 & ~n5067;
  assign n5069 = pi03 & ~n5066;
  assign n5070 = ~n5065 & n5069;
  assign n5071 = ~n5068 & ~n5070;
  assign n5072 = ~pi05 & ~n1548;
  assign n5073 = ~n5071 & n5072;
  assign n5074 = ~pi10 & n91;
  assign n5075 = ~n5070 & n5074;
  assign n5076 = ~n5068 & n5075;
  assign n5077 = ~n5073 & ~n5076;
  assign n5078 = n4909 & ~n5077;
  assign n5079 = ~n5063 & ~n5078;
  assign n5080 = ~n5056 & n5079;
  assign n5081 = ~pi05 & ~n5067;
  assign n5082 = ~n4909 & n5081;
  assign n5083 = ~n4908 & n5082;
  assign n5084 = n4908 & ~n5077;
  assign n5085 = ~n5083 & ~n5084;
  assign n5086 = n5080 & n5085;
  assign n5087 = ~n5054 & n5086;
  assign n5088 = ~n4909 & n5067;
  assign n5089 = ~n4908 & n5088;
  assign n5090 = ~n1548 & ~n5071;
  assign n5091 = n1548 & ~n5070;
  assign n5092 = ~n5068 & n5091;
  assign n5093 = ~n5090 & ~n5092;
  assign n5094 = ~n4926 & n5093;
  assign n5095 = ~n5089 & ~n5094;
  assign n5096 = pi05 & ~n5095;
  assign n5097 = ~n4619 & ~n4654;
  assign n5098 = ~n4643 & n5097;
  assign n5099 = ~n4618 & ~n4650;
  assign n5100 = ~n5098 & ~n5099;
  assign n5101 = ~n4650 & ~n4654;
  assign n5102 = ~n4619 & n5101;
  assign n5103 = ~n4618 & n5102;
  assign n5104 = ~n4643 & n5103;
  assign n5105 = ~pi07 & ~n5104;
  assign n5106 = ~n5100 & n5105;
  assign n5107 = ~n5100 & ~n5104;
  assign n5108 = pi07 & ~n5107;
  assign n5109 = ~n5106 & ~n5108;
  assign n5110 = ~n4926 & ~n5109;
  assign n5111 = n4670 & ~n5104;
  assign n5112 = n4671 & ~n5111;
  assign n5113 = n4670 & ~n4671;
  assign n5114 = ~n5104 & n5113;
  assign n5115 = ~pi09 & ~n5114;
  assign n5116 = ~n5112 & n5115;
  assign n5117 = ~n5112 & ~n5114;
  assign n5118 = pi09 & ~n5117;
  assign n5119 = ~n5116 & ~n5118;
  assign n5120 = ~n4926 & ~n5119;
  assign n5121 = ~n4604 & ~n4629;
  assign n5122 = ~n4370 & ~n4588;
  assign n5123 = ~n4602 & n5122;
  assign n5124 = ~n4587 & n5123;
  assign n5125 = ~pi09 & ~n5124;
  assign n5126 = ~n5121 & n5125;
  assign n5127 = ~n5121 & ~n5124;
  assign n5128 = pi09 & ~n5127;
  assign n5129 = ~n5126 & ~n5128;
  assign n5130 = ~n4909 & ~n5129;
  assign n5131 = ~n4908 & n5130;
  assign n5132 = ~n4604 & n4613;
  assign n5133 = ~n4588 & ~n4611;
  assign n5134 = ~n4602 & n5133;
  assign n5135 = ~n4587 & n5134;
  assign n5136 = ~pi07 & ~n5135;
  assign n5137 = ~n5132 & n5136;
  assign n5138 = ~n5132 & ~n5135;
  assign n5139 = pi07 & ~n5138;
  assign n5140 = ~n5137 & ~n5139;
  assign n5141 = ~n4909 & ~n5140;
  assign n5142 = ~n4908 & n5141;
  assign n5143 = ~n5131 & ~n5142;
  assign n5144 = ~n5120 & n5143;
  assign n5145 = ~n5110 & n5144;
  assign n5146 = ~n5096 & n5145;
  assign n5147 = ~n5087 & n5146;
  assign n5148 = ~n4926 & n5106;
  assign n5149 = ~n4909 & n5137;
  assign n5150 = ~n4908 & n5149;
  assign n5151 = ~n5148 & ~n5150;
  assign n5152 = ~n5120 & ~n5131;
  assign n5153 = ~n5151 & n5152;
  assign n5154 = ~n4704 & ~n4909;
  assign n5155 = ~n4908 & n5154;
  assign n5156 = ~n4681 & ~n4689;
  assign n5157 = ~n4705 & n5156;
  assign n5158 = ~n4673 & ~n4692;
  assign n5159 = ~n4672 & n5158;
  assign n5160 = ~n4665 & n5159;
  assign n5161 = ~n5157 & n5160;
  assign n5162 = n5157 & ~n5160;
  assign n5163 = ~n5161 & ~n5162;
  assign n5164 = n4908 & ~n5163;
  assign n5165 = n4909 & ~n5163;
  assign n5166 = ~pi11 & ~n5165;
  assign n5167 = ~n5164 & n5166;
  assign n5168 = ~n5155 & n5167;
  assign n5169 = ~n4926 & n5116;
  assign n5170 = ~n4909 & n5126;
  assign n5171 = ~n4908 & n5170;
  assign n5172 = ~n5169 & ~n5171;
  assign n5173 = ~n5168 & n5172;
  assign n5174 = ~n5153 & n5173;
  assign n5175 = ~n5147 & n5174;
  assign n5176 = ~n5164 & ~n5165;
  assign n5177 = ~n5155 & n5176;
  assign n5178 = pi11 & ~n5177;
  assign n5179 = ~n5016 & ~n5018;
  assign n5180 = ~n5178 & n5179;
  assign n5181 = ~n4929 & ~n4931;
  assign n5182 = pi13 & ~n5181;
  assign n5183 = ~n4933 & ~n5182;
  assign n5184 = ~n4926 & ~n5183;
  assign n5185 = ~n4818 & ~n4825;
  assign n5186 = pi13 & ~n5185;
  assign n5187 = ~n4923 & ~n5186;
  assign n5188 = ~n4909 & ~n5187;
  assign n5189 = ~n4908 & n5188;
  assign n5190 = ~n4942 & ~n5024;
  assign n5191 = ~n5189 & n5190;
  assign n5192 = ~n4956 & n5191;
  assign n5193 = ~n5184 & n5192;
  assign n5194 = ~n5003 & n5193;
  assign n5195 = n5180 & n5194;
  assign n5196 = ~n5175 & n5195;
  assign n5197 = ~n4926 & ~n5013;
  assign n5198 = ~n4810 & ~n4909;
  assign n5199 = ~n4908 & n5198;
  assign n5200 = ~pi19 & ~n5199;
  assign n5201 = ~n5197 & n5200;
  assign n5202 = ~n5003 & n5201;
  assign n5203 = ~n4926 & ~n4997;
  assign n5204 = n4814 & ~n4909;
  assign n5205 = ~n4908 & n5204;
  assign n5206 = ~pi21 & ~n5205;
  assign n5207 = ~n5203 & n5206;
  assign n5208 = ~n4920 & ~n5207;
  assign n5209 = ~n5202 & n5208;
  assign n5210 = ~n5196 & n5209;
  assign n5211 = ~n5028 & n5210;
  assign n5212 = ~n4921 & ~n5211;
  assign n5213 = ~n4908 & n5034;
  assign n5214 = n67 & n5042;
  assign n5215 = ~n4905 & n5214;
  assign n5216 = ~n4893 & n5215;
  assign n5217 = ~n4860 & n5216;
  assign n5218 = ~pi05 & ~n5217;
  assign n5219 = ~n5213 & n5218;
  assign n5220 = ~n5212 & n5219;
  assign n5221 = ~n5202 & ~n5207;
  assign n5222 = ~n5196 & n5221;
  assign n5223 = ~n5028 & n5222;
  assign n5224 = n2114 & ~n4918;
  assign n5225 = ~n5223 & n5224;
  assign n5226 = pi08 & ~n4920;
  assign n5227 = n2124 & ~n4916;
  assign n5228 = ~n2112 & ~n5227;
  assign n5229 = ~n5226 & n5228;
  assign n5230 = ~n5207 & ~n5229;
  assign n5231 = ~n5202 & n5230;
  assign n5232 = ~n5196 & n5231;
  assign n5233 = ~n5028 & n5232;
  assign n5234 = ~n4919 & ~n5229;
  assign n5235 = n2135 & ~n5234;
  assign n5236 = ~n5233 & n5235;
  assign n5237 = ~n5225 & n5236;
  assign n5238 = n2140 & ~n5217;
  assign n5239 = ~n5213 & n5238;
  assign n5240 = ~n5213 & ~n5217;
  assign n5241 = ~n2140 & ~n5240;
  assign n5242 = ~n5239 & ~n5241;
  assign n5243 = ~pi05 & ~n5242;
  assign n5244 = ~n4921 & n5243;
  assign n5245 = ~n5211 & n5244;
  assign n5246 = ~n5237 & ~n5245;
  assign n5247 = ~n5220 & n5246;
  assign n5248 = ~n5233 & ~n5234;
  assign n5249 = ~n5225 & n5248;
  assign n5250 = n2153 & ~n5249;
  assign n5251 = ~pi03 & ~n5249;
  assign n5252 = ~n5250 & ~n5251;
  assign n5253 = n5247 & n5252;
  assign n5254 = pi05 & ~n5239;
  assign n5255 = ~n5241 & n5254;
  assign n5256 = ~n4921 & n5255;
  assign n5257 = ~n5211 & n5256;
  assign n5258 = ~n5110 & ~n5142;
  assign n5259 = ~n5087 & ~n5096;
  assign n5260 = ~n5258 & ~n5259;
  assign n5261 = ~n5096 & n5258;
  assign n5262 = ~n5087 & n5261;
  assign n5263 = ~pi09 & ~n5262;
  assign n5264 = ~n5260 & n5263;
  assign n5265 = ~n5260 & ~n5262;
  assign n5266 = pi09 & ~n5265;
  assign n5267 = ~n5264 & ~n5266;
  assign n5268 = ~n4921 & ~n5267;
  assign n5269 = ~n5211 & n5268;
  assign n5270 = ~pi05 & ~n5089;
  assign n5271 = ~n5094 & n5270;
  assign n5272 = ~n5056 & ~n5063;
  assign n5273 = ~n5054 & n5272;
  assign n5274 = ~n5271 & n5273;
  assign n5275 = ~n5096 & n5274;
  assign n5276 = ~n5096 & ~n5271;
  assign n5277 = ~n5273 & ~n5276;
  assign n5278 = ~n5275 & ~n5277;
  assign n5279 = ~pi07 & ~n5278;
  assign n5280 = pi07 & ~n5275;
  assign n5281 = ~n5277 & n5280;
  assign n5282 = ~n5279 & ~n5281;
  assign n5283 = ~n4921 & ~n5282;
  assign n5284 = ~n5211 & n5283;
  assign n5285 = ~n5269 & ~n5284;
  assign n5286 = ~n5257 & n5285;
  assign n5287 = pi05 & ~n5240;
  assign n5288 = ~n5212 & n5287;
  assign n5289 = ~n4926 & ~n5107;
  assign n5290 = ~n4909 & ~n5138;
  assign n5291 = ~n4908 & n5290;
  assign n5292 = ~pi09 & ~n5291;
  assign n5293 = ~n5289 & n5292;
  assign n5294 = ~n5289 & ~n5291;
  assign n5295 = pi09 & ~n5294;
  assign n5296 = ~n5293 & ~n5295;
  assign n5297 = ~n5212 & ~n5296;
  assign n5298 = ~pi07 & ~n5089;
  assign n5299 = ~n5094 & n5298;
  assign n5300 = pi07 & ~n5095;
  assign n5301 = ~n5299 & ~n5300;
  assign n5302 = ~n5212 & ~n5301;
  assign n5303 = ~n5297 & ~n5302;
  assign n5304 = ~n5288 & n5303;
  assign n5305 = n5286 & n5304;
  assign n5306 = ~n5253 & n5305;
  assign n5307 = ~n4926 & ~n5117;
  assign n5308 = ~n4909 & ~n5127;
  assign n5309 = ~n4908 & n5308;
  assign n5310 = ~pi11 & ~n5309;
  assign n5311 = ~n5307 & n5310;
  assign n5312 = ~n5212 & n5311;
  assign n5313 = n4935 & ~n4957;
  assign n5314 = ~n4958 & n5174;
  assign n5315 = ~n5313 & n5314;
  assign n5316 = ~n5147 & n5315;
  assign n5317 = ~n5184 & ~n5189;
  assign n5318 = ~n5178 & n5317;
  assign n5319 = n5313 & ~n5318;
  assign n5320 = ~n4942 & ~n5189;
  assign n5321 = ~n4956 & n5320;
  assign n5322 = ~n5184 & n5321;
  assign n5323 = ~n5178 & n5322;
  assign n5324 = ~n4958 & ~n5323;
  assign n5325 = ~n5319 & n5324;
  assign n5326 = ~n5175 & n5325;
  assign n5327 = ~n5316 & ~n5326;
  assign n5328 = ~pi17 & ~n4921;
  assign n5329 = ~n5211 & n5328;
  assign n5330 = ~n5327 & n5329;
  assign n5331 = ~n5212 & n5293;
  assign n5332 = ~n5330 & ~n5331;
  assign n5333 = ~n5312 & n5332;
  assign n5334 = n5151 & ~n5262;
  assign n5335 = n5152 & ~n5334;
  assign n5336 = n5151 & ~n5152;
  assign n5337 = ~n5262 & n5336;
  assign n5338 = ~pi11 & ~n4921;
  assign n5339 = ~n5337 & n5338;
  assign n5340 = ~n5335 & n5339;
  assign n5341 = ~n5211 & n5340;
  assign n5342 = ~n5087 & ~n5178;
  assign n5343 = n5146 & n5342;
  assign n5344 = ~n5174 & ~n5178;
  assign n5345 = ~n5317 & ~n5344;
  assign n5346 = ~n5343 & n5345;
  assign n5347 = ~n5343 & ~n5344;
  assign n5348 = n5317 & ~n5347;
  assign n5349 = ~pi15 & ~n4921;
  assign n5350 = ~n5348 & n5349;
  assign n5351 = ~n5346 & n5350;
  assign n5352 = ~n5211 & n5351;
  assign n5353 = ~n4921 & ~n5260;
  assign n5354 = n5263 & n5353;
  assign n5355 = ~n5211 & n5354;
  assign n5356 = ~n5352 & ~n5355;
  assign n5357 = ~n5341 & n5356;
  assign n5358 = ~n4926 & ~n5181;
  assign n5359 = ~n4909 & ~n5185;
  assign n5360 = ~n4908 & n5359;
  assign n5361 = ~pi15 & ~n5360;
  assign n5362 = ~n5358 & n5361;
  assign n5363 = ~n5212 & n5362;
  assign n5364 = ~pi17 & ~n4961;
  assign n5365 = ~n4959 & n5364;
  assign n5366 = ~n5212 & n5365;
  assign n5367 = ~n5363 & ~n5366;
  assign n5368 = n5357 & n5367;
  assign n5369 = n5333 & n5368;
  assign n5370 = ~pi13 & ~n5165;
  assign n5371 = ~n5164 & n5370;
  assign n5372 = ~n5155 & n5371;
  assign n5373 = ~n5212 & n5372;
  assign n5374 = n5174 & ~n5178;
  assign n5375 = ~n5147 & n5374;
  assign n5376 = ~n5153 & n5172;
  assign n5377 = ~n5147 & n5376;
  assign n5378 = ~n5168 & ~n5178;
  assign n5379 = ~n5377 & ~n5378;
  assign n5380 = ~n5375 & ~n5379;
  assign n5381 = ~pi13 & ~n4921;
  assign n5382 = ~n5380 & n5381;
  assign n5383 = ~n5211 & n5382;
  assign n5384 = ~n5373 & ~n5383;
  assign n5385 = ~n5358 & ~n5360;
  assign n5386 = pi15 & ~n5385;
  assign n5387 = ~n5362 & ~n5386;
  assign n5388 = ~n5212 & ~n5387;
  assign n5389 = ~pi15 & ~n5189;
  assign n5390 = ~n5184 & n5389;
  assign n5391 = pi15 & ~n5317;
  assign n5392 = ~n5390 & ~n5391;
  assign n5393 = ~n5344 & n5392;
  assign n5394 = ~n5343 & n5393;
  assign n5395 = ~n5347 & ~n5392;
  assign n5396 = ~n4921 & ~n5395;
  assign n5397 = ~n5394 & n5396;
  assign n5398 = ~n5211 & n5397;
  assign n5399 = ~n5388 & ~n5398;
  assign n5400 = ~n5384 & n5399;
  assign n5401 = ~n5212 & n5299;
  assign n5402 = ~pi07 & ~n4921;
  assign n5403 = ~n5278 & n5402;
  assign n5404 = ~n5211 & n5403;
  assign n5405 = ~n5401 & ~n5404;
  assign n5406 = ~n5269 & ~n5297;
  assign n5407 = ~n5405 & n5406;
  assign n5408 = ~n5400 & ~n5407;
  assign n5409 = n5369 & n5408;
  assign n5410 = ~n5306 & n5409;
  assign n5411 = pi13 & ~n5177;
  assign n5412 = ~n5372 & ~n5411;
  assign n5413 = ~n5212 & ~n5412;
  assign n5414 = ~n5335 & ~n5337;
  assign n5415 = pi11 & ~n4921;
  assign n5416 = ~n5414 & n5415;
  assign n5417 = ~n5211 & n5416;
  assign n5418 = ~n5398 & ~n5417;
  assign n5419 = ~n5413 & n5418;
  assign n5420 = ~n5307 & ~n5309;
  assign n5421 = pi11 & ~n5420;
  assign n5422 = ~n5212 & n5421;
  assign n5423 = ~pi13 & ~n5380;
  assign n5424 = pi13 & ~n5375;
  assign n5425 = ~n5379 & n5424;
  assign n5426 = ~n5423 & ~n5425;
  assign n5427 = n5212 & ~n5426;
  assign n5428 = ~n5388 & ~n5427;
  assign n5429 = ~n5422 & n5428;
  assign n5430 = n5419 & n5429;
  assign n5431 = ~n5352 & ~n5363;
  assign n5432 = ~n5330 & ~n5366;
  assign n5433 = n5431 & n5432;
  assign n5434 = ~n5400 & n5433;
  assign n5435 = ~n5430 & n5434;
  assign n5436 = ~n5203 & ~n5205;
  assign n5437 = ~n5212 & ~n5436;
  assign n5438 = ~n5018 & ~n5178;
  assign n5439 = n5322 & n5438;
  assign n5440 = ~n5175 & n5439;
  assign n5441 = ~n4977 & ~n5018;
  assign n5442 = ~n4990 & ~n5201;
  assign n5443 = n5002 & n5442;
  assign n5444 = ~n5202 & ~n5443;
  assign n5445 = ~n5441 & n5444;
  assign n5446 = ~n5440 & n5445;
  assign n5447 = ~n5197 & ~n5199;
  assign n5448 = pi19 & ~n5447;
  assign n5449 = ~n5003 & ~n5448;
  assign n5450 = pi19 & ~n4996;
  assign n5451 = ~n5001 & n5450;
  assign n5452 = ~n4990 & ~n5447;
  assign n5453 = n5451 & n5452;
  assign n5454 = n5439 & ~n5453;
  assign n5455 = ~n5449 & n5454;
  assign n5456 = ~n5175 & n5455;
  assign n5457 = ~n5018 & ~n5453;
  assign n5458 = ~n4977 & n5457;
  assign n5459 = ~n5449 & n5458;
  assign n5460 = ~n4921 & ~n5459;
  assign n5461 = ~n5456 & n5460;
  assign n5462 = ~n5446 & n5461;
  assign n5463 = ~n5211 & n5462;
  assign n5464 = ~n5437 & ~n5463;
  assign n5465 = pi23 & ~n5464;
  assign n5466 = ~n5016 & ~n5024;
  assign n5467 = ~n5441 & n5466;
  assign n5468 = ~n5440 & n5467;
  assign n5469 = n5439 & ~n5466;
  assign n5470 = ~n5175 & n5469;
  assign n5471 = ~n5018 & ~n5466;
  assign n5472 = ~n4977 & n5471;
  assign n5473 = pi21 & ~n4921;
  assign n5474 = ~n5472 & n5473;
  assign n5475 = ~n5470 & n5474;
  assign n5476 = ~n5468 & n5475;
  assign n5477 = ~n5211 & n5476;
  assign n5478 = pi17 & ~n4921;
  assign n5479 = ~n5316 & n5478;
  assign n5480 = ~n5326 & n5479;
  assign n5481 = ~n5211 & n5480;
  assign n5482 = n67 & ~n5481;
  assign n5483 = ~n5477 & n5482;
  assign n5484 = ~n5470 & ~n5472;
  assign n5485 = ~n5468 & n5484;
  assign n5486 = ~pi21 & ~n4921;
  assign n5487 = ~n5211 & n5486;
  assign n5488 = ~n5485 & n5487;
  assign n5489 = ~n4959 & ~n4961;
  assign n5490 = pi17 & ~n5489;
  assign n5491 = ~n5212 & n5490;
  assign n5492 = ~pi21 & ~n5199;
  assign n5493 = ~n5197 & n5492;
  assign n5494 = pi21 & ~n5447;
  assign n5495 = ~n5493 & ~n5494;
  assign n5496 = ~n5212 & ~n5495;
  assign n5497 = ~n5491 & ~n5496;
  assign n5498 = ~n5488 & n5497;
  assign n5499 = n5483 & n5498;
  assign n5500 = ~n5465 & n5499;
  assign n5501 = n4918 & ~n4921;
  assign n5502 = ~n5211 & n5501;
  assign n5503 = ~n5223 & n5502;
  assign n5504 = ~n4916 & ~n5212;
  assign n5505 = ~pi25 & ~n5504;
  assign n5506 = ~n5503 & n5505;
  assign n5507 = ~n5503 & ~n5504;
  assign n5508 = pi25 & ~n5507;
  assign n5509 = ~n5506 & ~n5508;
  assign n5510 = ~n5017 & ~n5212;
  assign n5511 = ~n4963 & ~n5184;
  assign n5512 = n5321 & n5511;
  assign n5513 = ~n5178 & n5512;
  assign n5514 = ~n4958 & n5513;
  assign n5515 = ~n5175 & n5514;
  assign n5516 = n4976 & ~n5018;
  assign n5517 = ~n4958 & n5516;
  assign n5518 = ~n4958 & ~n4963;
  assign n5519 = ~n4975 & ~n5018;
  assign n5520 = ~n5518 & ~n5519;
  assign n5521 = ~n5517 & ~n5520;
  assign n5522 = n5515 & n5521;
  assign n5523 = ~n5515 & ~n5521;
  assign n5524 = ~n4921 & ~n5523;
  assign n5525 = ~n5522 & n5524;
  assign n5526 = ~n5211 & n5525;
  assign n5527 = ~n5510 & ~n5526;
  assign n5528 = ~pi19 & ~n5527;
  assign n5529 = pi19 & ~n5510;
  assign n5530 = ~n5526 & n5529;
  assign n5531 = ~n5528 & ~n5530;
  assign n5532 = ~n5509 & ~n5531;
  assign n5533 = n5500 & n5532;
  assign n5534 = ~n5435 & n5533;
  assign n5535 = ~n5410 & n5534;
  assign n5536 = ~pi19 & ~n5477;
  assign n5537 = ~n5510 & n5536;
  assign n5538 = ~n5496 & ~n5526;
  assign n5539 = ~n5488 & n5538;
  assign n5540 = n5537 & n5539;
  assign n5541 = ~n5212 & ~n5447;
  assign n5542 = ~n4921 & ~n5472;
  assign n5543 = ~n5470 & n5542;
  assign n5544 = ~n5468 & n5543;
  assign n5545 = ~n5211 & n5544;
  assign n5546 = ~pi21 & ~n5545;
  assign n5547 = ~n5541 & n5546;
  assign n5548 = ~pi23 & ~n5437;
  assign n5549 = ~n5463 & n5548;
  assign n5550 = ~n5547 & ~n5549;
  assign n5551 = ~n5540 & n5550;
  assign n5552 = n67 & ~n5465;
  assign n5553 = ~n5509 & n5552;
  assign n5554 = ~n5551 & n5553;
  assign n5555 = n69 & ~n5507;
  assign n5556 = ~n5554 & ~n5555;
  assign n5557 = ~n5535 & n5556;
  assign n5558 = ~n5477 & ~n5481;
  assign n5559 = ~n5491 & n5558;
  assign n5560 = ~n5488 & ~n5496;
  assign n5561 = n5559 & n5560;
  assign n5562 = ~n5531 & n5561;
  assign n5563 = ~n5435 & n5562;
  assign n5564 = ~n5410 & n5563;
  assign n5565 = n5551 & ~n5564;
  assign n5566 = ~n5465 & n5509;
  assign n5567 = ~n5565 & n5566;
  assign n5568 = ~n5557 & n5567;
  assign n5569 = ~n5507 & ~n5555;
  assign n5570 = ~n5554 & n5569;
  assign n5571 = ~n5535 & n5570;
  assign n5572 = ~pi27 & ~n5571;
  assign n5573 = ~n5568 & n5572;
  assign n5574 = ~n5568 & ~n5571;
  assign n5575 = pi27 & ~n5574;
  assign n5576 = ~n5573 & ~n5575;
  assign n5577 = ~n2997 & ~n5576;
  assign n5578 = n3000 & ~n5574;
  assign n5579 = pi04 & ~n5578;
  assign n5580 = ~n5577 & n5579;
  assign n5581 = pi03 & ~n5234;
  assign n5582 = ~n5233 & n5581;
  assign n5583 = ~n5225 & n5582;
  assign n5584 = ~n5251 & ~n5583;
  assign n5585 = ~n2134 & ~n5584;
  assign n5586 = n2134 & ~n5583;
  assign n5587 = ~n5251 & n5586;
  assign n5588 = ~n5585 & ~n5587;
  assign n5589 = ~pi05 & ~n5588;
  assign n5590 = ~n5557 & n5589;
  assign n5591 = pi06 & ~n5555;
  assign n5592 = n69 & n2134;
  assign n5593 = ~n5507 & n5592;
  assign n5594 = ~n2606 & ~n5593;
  assign n5595 = ~n5591 & n5594;
  assign n5596 = ~n5554 & ~n5595;
  assign n5597 = ~n5535 & n5596;
  assign n5598 = n2608 & ~n5481;
  assign n5599 = ~n5477 & n5598;
  assign n5600 = n5498 & n5599;
  assign n5601 = ~n5465 & n5600;
  assign n5602 = n5532 & n5601;
  assign n5603 = ~n5435 & n5602;
  assign n5604 = ~n5410 & n5603;
  assign n5605 = n2608 & ~n5465;
  assign n5606 = ~n5509 & n5605;
  assign n5607 = ~n5551 & n5606;
  assign n5608 = n2620 & ~n5607;
  assign n5609 = ~n5604 & n5608;
  assign n5610 = ~n5597 & n5609;
  assign n5611 = ~pi05 & ~n5249;
  assign n5612 = ~n5555 & n5611;
  assign n5613 = ~n5554 & n5612;
  assign n5614 = ~n5535 & n5613;
  assign n5615 = ~n5610 & ~n5614;
  assign n5616 = ~n5590 & n5615;
  assign n5617 = ~n5604 & ~n5607;
  assign n5618 = ~n5597 & n5617;
  assign n5619 = n2632 & ~n5618;
  assign n5620 = ~pi03 & ~n5618;
  assign n5621 = ~n5619 & ~n5620;
  assign n5622 = n5616 & n5621;
  assign n5623 = pi05 & ~n5234;
  assign n5624 = ~n5233 & n5623;
  assign n5625 = ~n5225 & n5624;
  assign n5626 = ~n5555 & n5625;
  assign n5627 = ~n5554 & n5626;
  assign n5628 = ~n5535 & n5627;
  assign n5629 = ~n5095 & ~n5212;
  assign n5630 = ~n4921 & ~n5275;
  assign n5631 = ~n5277 & n5630;
  assign n5632 = ~n5211 & n5631;
  assign n5633 = ~pi09 & ~n5632;
  assign n5634 = ~n5629 & n5633;
  assign n5635 = ~n5629 & ~n5632;
  assign n5636 = pi09 & ~n5635;
  assign n5637 = ~n5634 & ~n5636;
  assign n5638 = ~n5555 & ~n5637;
  assign n5639 = ~n5554 & n5638;
  assign n5640 = ~n5535 & n5639;
  assign n5641 = ~n5212 & ~n5240;
  assign n5642 = ~n4921 & n5242;
  assign n5643 = ~n5211 & n5642;
  assign n5644 = ~pi07 & ~n5643;
  assign n5645 = ~n5641 & n5644;
  assign n5646 = ~n5641 & ~n5643;
  assign n5647 = pi07 & ~n5646;
  assign n5648 = ~n5645 & ~n5647;
  assign n5649 = ~n5555 & ~n5648;
  assign n5650 = ~n5554 & n5649;
  assign n5651 = ~n5535 & n5650;
  assign n5652 = ~n5640 & ~n5651;
  assign n5653 = ~n5628 & n5652;
  assign n5654 = pi05 & ~n5587;
  assign n5655 = ~n5585 & n5654;
  assign n5656 = ~n5557 & n5655;
  assign n5657 = ~n5284 & ~n5302;
  assign n5658 = ~n5257 & ~n5288;
  assign n5659 = ~n5253 & n5658;
  assign n5660 = ~n5657 & ~n5659;
  assign n5661 = ~n5257 & ~n5284;
  assign n5662 = ~n5302 & n5661;
  assign n5663 = ~n5288 & n5662;
  assign n5664 = ~n5253 & n5663;
  assign n5665 = ~pi09 & ~n5664;
  assign n5666 = ~n5660 & n5665;
  assign n5667 = ~n5660 & ~n5664;
  assign n5668 = pi09 & ~n5667;
  assign n5669 = ~n5666 & ~n5668;
  assign n5670 = ~n5557 & ~n5669;
  assign n5671 = ~pi05 & ~n5646;
  assign n5672 = pi05 & ~n5643;
  assign n5673 = ~n5641 & n5672;
  assign n5674 = ~n5671 & ~n5673;
  assign n5675 = ~n5237 & ~n5250;
  assign n5676 = ~n5251 & n5675;
  assign n5677 = ~n5674 & ~n5676;
  assign n5678 = ~n5251 & ~n5673;
  assign n5679 = n5675 & n5678;
  assign n5680 = ~n5671 & n5679;
  assign n5681 = ~pi07 & ~n5680;
  assign n5682 = ~n5677 & n5681;
  assign n5683 = ~n5677 & ~n5680;
  assign n5684 = pi07 & ~n5683;
  assign n5685 = ~n5682 & ~n5684;
  assign n5686 = ~n5557 & ~n5685;
  assign n5687 = ~n5670 & ~n5686;
  assign n5688 = ~n5656 & n5687;
  assign n5689 = n5653 & n5688;
  assign n5690 = ~n5622 & n5689;
  assign n5691 = ~n5177 & ~n5212;
  assign n5692 = ~n4921 & ~n5375;
  assign n5693 = ~n5379 & n5692;
  assign n5694 = ~n5211 & n5693;
  assign n5695 = ~pi15 & ~n5694;
  assign n5696 = ~n5691 & n5695;
  assign n5697 = ~n5555 & n5696;
  assign n5698 = ~n5554 & n5697;
  assign n5699 = ~n5535 & n5698;
  assign n5700 = ~n5212 & ~n5385;
  assign n5701 = ~n5346 & ~n5348;
  assign n5702 = ~n4921 & ~n5701;
  assign n5703 = ~n5211 & n5702;
  assign n5704 = ~pi17 & ~n5703;
  assign n5705 = ~n5700 & n5704;
  assign n5706 = ~n5555 & n5705;
  assign n5707 = ~n5554 & n5706;
  assign n5708 = ~n5535 & n5707;
  assign n5709 = ~n5699 & ~n5708;
  assign n5710 = ~n5555 & n5634;
  assign n5711 = ~n5554 & n5710;
  assign n5712 = ~n5535 & n5711;
  assign n5713 = ~n5212 & ~n5294;
  assign n5714 = ~n4921 & ~n5265;
  assign n5715 = ~n5211 & n5714;
  assign n5716 = ~pi11 & ~n5715;
  assign n5717 = ~n5713 & n5716;
  assign n5718 = ~n5555 & n5717;
  assign n5719 = ~n5554 & n5718;
  assign n5720 = ~n5535 & n5719;
  assign n5721 = ~n5712 & ~n5720;
  assign n5722 = n5709 & n5721;
  assign n5723 = ~n5341 & ~n5355;
  assign n5724 = ~n5331 & n5723;
  assign n5725 = ~n5312 & n5724;
  assign n5726 = ~n5407 & n5725;
  assign n5727 = ~n5306 & n5726;
  assign n5728 = ~n5413 & ~n5427;
  assign n5729 = ~pi15 & ~n5417;
  assign n5730 = ~n5422 & n5729;
  assign n5731 = ~n5728 & n5730;
  assign n5732 = ~n5727 & n5731;
  assign n5733 = ~n5417 & ~n5422;
  assign n5734 = ~n5727 & n5733;
  assign n5735 = ~pi15 & ~n5413;
  assign n5736 = ~n5427 & n5735;
  assign n5737 = ~n5734 & n5736;
  assign n5738 = ~n5732 & ~n5737;
  assign n5739 = ~n5557 & ~n5738;
  assign n5740 = ~n5691 & ~n5694;
  assign n5741 = pi13 & ~n5740;
  assign n5742 = ~n5399 & n5741;
  assign n5743 = n5399 & ~n5741;
  assign n5744 = n5733 & ~n5743;
  assign n5745 = ~n5742 & n5744;
  assign n5746 = ~n5727 & n5745;
  assign n5747 = ~n5383 & ~n5398;
  assign n5748 = ~n5388 & n5747;
  assign n5749 = ~n5373 & n5748;
  assign n5750 = ~n5384 & ~n5399;
  assign n5751 = ~n5749 & ~n5750;
  assign n5752 = ~n5733 & ~n5751;
  assign n5753 = n5726 & ~n5751;
  assign n5754 = ~n5306 & n5753;
  assign n5755 = ~n5752 & ~n5754;
  assign n5756 = ~n5746 & n5755;
  assign n5757 = ~pi17 & ~n5756;
  assign n5758 = ~n5557 & n5757;
  assign n5759 = ~n5739 & ~n5758;
  assign n5760 = ~n5557 & n5666;
  assign n5761 = n5405 & ~n5664;
  assign n5762 = n5406 & ~n5761;
  assign n5763 = n5405 & ~n5406;
  assign n5764 = ~n5664 & n5763;
  assign n5765 = ~pi11 & ~n5764;
  assign n5766 = ~n5762 & n5765;
  assign n5767 = ~n5557 & n5766;
  assign n5768 = ~n5760 & ~n5767;
  assign n5769 = n5759 & n5768;
  assign n5770 = n5722 & n5769;
  assign n5771 = ~n5341 & ~n5417;
  assign n5772 = ~n5422 & n5771;
  assign n5773 = ~n5312 & n5772;
  assign n5774 = ~n5331 & ~n5355;
  assign n5775 = ~n5407 & n5774;
  assign n5776 = ~n5306 & n5775;
  assign n5777 = n5773 & ~n5776;
  assign n5778 = ~n5773 & n5775;
  assign n5779 = ~n5306 & n5778;
  assign n5780 = ~pi13 & ~n5779;
  assign n5781 = ~n5777 & n5780;
  assign n5782 = ~n5557 & n5781;
  assign n5783 = ~n5212 & ~n5420;
  assign n5784 = ~n4921 & ~n5414;
  assign n5785 = ~n5211 & n5784;
  assign n5786 = ~pi13 & ~n5785;
  assign n5787 = ~n5783 & n5786;
  assign n5788 = ~n5555 & n5787;
  assign n5789 = ~n5554 & n5788;
  assign n5790 = ~n5535 & n5789;
  assign n5791 = ~n5782 & ~n5790;
  assign n5792 = pi15 & ~n5740;
  assign n5793 = ~n5696 & ~n5792;
  assign n5794 = ~n5555 & ~n5793;
  assign n5795 = ~n5554 & n5794;
  assign n5796 = ~n5535 & n5795;
  assign n5797 = pi15 & ~n5355;
  assign n5798 = ~n5341 & n5797;
  assign n5799 = ~n5312 & ~n5331;
  assign n5800 = n5728 & n5799;
  assign n5801 = n5798 & n5800;
  assign n5802 = ~n5407 & n5801;
  assign n5803 = ~n5306 & n5802;
  assign n5804 = ~pi15 & ~n5355;
  assign n5805 = ~n5341 & n5804;
  assign n5806 = n5799 & n5805;
  assign n5807 = ~n5728 & n5806;
  assign n5808 = ~n5407 & n5807;
  assign n5809 = ~n5306 & n5808;
  assign n5810 = ~pi15 & ~n5733;
  assign n5811 = ~n5728 & n5810;
  assign n5812 = pi15 & ~n5413;
  assign n5813 = ~n5427 & n5812;
  assign n5814 = ~n5733 & n5813;
  assign n5815 = ~n5811 & ~n5814;
  assign n5816 = ~n5809 & n5815;
  assign n5817 = ~n5803 & n5816;
  assign n5818 = ~n5413 & n5729;
  assign n5819 = ~n5422 & ~n5427;
  assign n5820 = n5818 & n5819;
  assign n5821 = ~n5727 & n5820;
  assign n5822 = pi15 & ~n5417;
  assign n5823 = ~n5422 & n5822;
  assign n5824 = ~n5728 & n5823;
  assign n5825 = ~n5727 & n5824;
  assign n5826 = ~n5821 & ~n5825;
  assign n5827 = n5817 & n5826;
  assign n5828 = ~n5557 & n5827;
  assign n5829 = ~n5796 & ~n5828;
  assign n5830 = ~n5791 & n5829;
  assign n5831 = ~n5557 & n5682;
  assign n5832 = ~n5555 & n5645;
  assign n5833 = ~n5554 & n5832;
  assign n5834 = ~n5535 & n5833;
  assign n5835 = ~n5831 & ~n5834;
  assign n5836 = ~n5640 & ~n5670;
  assign n5837 = ~n5835 & n5836;
  assign n5838 = ~n5830 & ~n5837;
  assign n5839 = n5770 & n5838;
  assign n5840 = ~n5690 & n5839;
  assign n5841 = ~n5777 & ~n5779;
  assign n5842 = pi13 & ~n5841;
  assign n5843 = ~n5781 & ~n5842;
  assign n5844 = ~n5557 & ~n5843;
  assign n5845 = ~n5713 & ~n5715;
  assign n5846 = pi11 & ~n5845;
  assign n5847 = ~n5555 & n5846;
  assign n5848 = ~n5554 & n5847;
  assign n5849 = ~n5535 & n5848;
  assign n5850 = ~n5783 & ~n5785;
  assign n5851 = pi13 & ~n5850;
  assign n5852 = ~n5787 & ~n5851;
  assign n5853 = ~n5555 & ~n5852;
  assign n5854 = ~n5554 & n5853;
  assign n5855 = ~n5535 & n5854;
  assign n5856 = ~n5796 & ~n5855;
  assign n5857 = ~n5849 & n5856;
  assign n5858 = ~n5762 & ~n5764;
  assign n5859 = pi11 & ~n5858;
  assign n5860 = ~n5557 & n5859;
  assign n5861 = ~n5828 & ~n5860;
  assign n5862 = n5857 & n5861;
  assign n5863 = ~n5844 & n5862;
  assign n5864 = n5709 & ~n5739;
  assign n5865 = ~n5758 & n5864;
  assign n5866 = ~n5830 & n5865;
  assign n5867 = ~n5863 & n5866;
  assign n5868 = ~n5481 & ~n5491;
  assign n5869 = ~n5531 & n5868;
  assign n5870 = ~n5435 & n5869;
  assign n5871 = ~n5410 & n5870;
  assign n5872 = ~n5435 & n5868;
  assign n5873 = ~n5410 & n5872;
  assign n5874 = n5531 & ~n5873;
  assign n5875 = ~n5871 & ~n5874;
  assign n5876 = ~n5557 & ~n5875;
  assign n5877 = ~n5527 & ~n5555;
  assign n5878 = ~n5554 & n5877;
  assign n5879 = ~n5535 & n5878;
  assign n5880 = ~pi21 & ~n5879;
  assign n5881 = ~n5876 & n5880;
  assign n5882 = ~n5366 & ~n5481;
  assign n5883 = ~n5330 & ~n5491;
  assign n5884 = n5882 & n5883;
  assign n5885 = ~n5400 & n5431;
  assign n5886 = ~n5430 & n5885;
  assign n5887 = ~n5331 & ~n5363;
  assign n5888 = ~n5312 & n5887;
  assign n5889 = n5357 & n5888;
  assign n5890 = n5408 & n5889;
  assign n5891 = ~n5306 & n5890;
  assign n5892 = ~n5886 & ~n5891;
  assign n5893 = ~n5884 & ~n5892;
  assign n5894 = n5884 & ~n5886;
  assign n5895 = ~n5891 & n5894;
  assign n5896 = ~n5893 & ~n5895;
  assign n5897 = ~n5557 & n5896;
  assign n5898 = ~n5212 & ~n5489;
  assign n5899 = ~n4921 & ~n5316;
  assign n5900 = ~n5326 & n5899;
  assign n5901 = ~n5211 & n5900;
  assign n5902 = ~n5898 & ~n5901;
  assign n5903 = ~n5555 & n5902;
  assign n5904 = ~n5554 & n5903;
  assign n5905 = ~n5535 & n5904;
  assign n5906 = pi19 & ~n5905;
  assign n5907 = ~n5897 & n5906;
  assign n5908 = pi17 & ~n5752;
  assign n5909 = ~n5754 & n5908;
  assign n5910 = ~n5746 & n5909;
  assign n5911 = ~n5557 & n5910;
  assign n5912 = ~n5700 & ~n5703;
  assign n5913 = pi17 & ~n5912;
  assign n5914 = ~n5555 & n5913;
  assign n5915 = ~n5554 & n5914;
  assign n5916 = ~n5535 & n5915;
  assign n5917 = ~n5911 & ~n5916;
  assign n5918 = ~n5907 & n5917;
  assign n5919 = ~n5881 & n5918;
  assign n5920 = ~n5897 & ~n5905;
  assign n5921 = ~pi19 & ~n5920;
  assign n5922 = ~n5876 & ~n5879;
  assign n5923 = pi21 & ~n5922;
  assign n5924 = ~n5921 & ~n5923;
  assign n5925 = ~n5465 & n5550;
  assign n5926 = ~n5540 & n5925;
  assign n5927 = ~n5564 & n5926;
  assign n5928 = pi25 & ~n5556;
  assign n5929 = pi25 & ~pi27;
  assign n5930 = n65 & n5929;
  assign n5931 = ~n5481 & n5930;
  assign n5932 = ~n5477 & n5931;
  assign n5933 = n5498 & n5932;
  assign n5934 = ~n5465 & n5933;
  assign n5935 = n5532 & n5934;
  assign n5936 = ~n5435 & n5935;
  assign n5937 = ~n5410 & n5936;
  assign n5938 = ~n5928 & ~n5937;
  assign n5939 = ~n5927 & n5938;
  assign n5940 = ~pi25 & ~n5437;
  assign n5941 = ~n5463 & n5940;
  assign n5942 = pi25 & ~n5464;
  assign n5943 = ~n5941 & ~n5942;
  assign n5944 = ~n5555 & ~n5943;
  assign n5945 = ~n5554 & n5944;
  assign n5946 = ~n5535 & n5945;
  assign n5947 = ~n5540 & ~n5547;
  assign n5948 = ~n5564 & n5947;
  assign n5949 = ~n5465 & ~n5549;
  assign n5950 = ~n5948 & ~n5949;
  assign n5951 = ~n5946 & ~n5950;
  assign n5952 = n5939 & n5951;
  assign n5953 = ~n5927 & ~n5950;
  assign n5954 = n69 & ~n5481;
  assign n5955 = ~n5477 & n5954;
  assign n5956 = n5498 & n5955;
  assign n5957 = ~n5465 & n5956;
  assign n5958 = n5532 & n5957;
  assign n5959 = ~n5435 & n5958;
  assign n5960 = ~n5410 & n5959;
  assign n5961 = ~pi25 & ~n5556;
  assign n5962 = ~n5960 & ~n5961;
  assign n5963 = ~n5946 & n5962;
  assign n5964 = ~n5953 & n5963;
  assign n5965 = ~n5952 & ~n5964;
  assign n5966 = ~n5541 & ~n5545;
  assign n5967 = ~n5555 & n5966;
  assign n5968 = ~n5554 & n5967;
  assign n5969 = ~n5535 & n5968;
  assign n5970 = pi23 & ~n5969;
  assign n5971 = n65 & ~n5970;
  assign n5972 = ~n5477 & ~n5496;
  assign n5973 = ~n5488 & n5972;
  assign n5974 = ~pi19 & ~n5510;
  assign n5975 = ~n5526 & n5974;
  assign n5976 = ~n5871 & ~n5975;
  assign n5977 = n5973 & ~n5976;
  assign n5978 = ~n5973 & ~n5975;
  assign n5979 = ~n5871 & n5978;
  assign n5980 = n65 & ~n5979;
  assign n5981 = ~n5557 & n5980;
  assign n5982 = ~n5977 & n5981;
  assign n5983 = ~n5971 & ~n5982;
  assign n5984 = ~n5965 & ~n5983;
  assign n5985 = n5924 & n5984;
  assign n5986 = n5919 & n5985;
  assign n5987 = ~n5867 & n5986;
  assign n5988 = ~n5840 & n5987;
  assign n5989 = ~n5881 & n5921;
  assign n5990 = ~n5923 & n5989;
  assign n5991 = ~pi23 & ~n5979;
  assign n5992 = ~n5557 & n5991;
  assign n5993 = ~n5977 & n5992;
  assign n5994 = ~pi23 & ~n5545;
  assign n5995 = ~n5541 & n5994;
  assign n5996 = ~n5555 & n5995;
  assign n5997 = ~n5554 & n5996;
  assign n5998 = ~n5535 & n5997;
  assign n5999 = ~n5881 & ~n5998;
  assign n6000 = ~n5993 & n5999;
  assign n6001 = ~n5990 & n6000;
  assign n6002 = n5984 & ~n6001;
  assign n6003 = ~n5557 & n5953;
  assign n6004 = ~n5464 & ~n5555;
  assign n6005 = ~n5554 & n6004;
  assign n6006 = ~n5535 & n6005;
  assign n6007 = n2573 & ~n6006;
  assign n6008 = ~n6003 & n6007;
  assign n6009 = n5579 & ~n6008;
  assign n6010 = ~n6002 & n6009;
  assign n6011 = ~n5988 & n6010;
  assign n6012 = ~n5580 & ~n6011;
  assign n6013 = ~n3013 & ~n6012;
  assign n6014 = n3015 & ~n5574;
  assign n6015 = pi03 & ~n6008;
  assign n6016 = ~n6014 & n6015;
  assign n6017 = ~n6002 & n6016;
  assign n6018 = ~n5988 & n6017;
  assign n6019 = n3012 & ~n6008;
  assign n6020 = ~n6014 & n6019;
  assign n6021 = ~n6002 & n6020;
  assign n6022 = ~n5988 & n6021;
  assign n6023 = ~pi27 & ~n65;
  assign n6024 = ~n5574 & ~n6023;
  assign n6025 = ~n5573 & ~n6024;
  assign n6026 = n2619 & ~n6025;
  assign n6027 = n3012 & ~n6026;
  assign n6028 = n3029 & ~n6025;
  assign n6029 = pi03 & ~n6028;
  assign n6030 = ~n6027 & ~n6029;
  assign n6031 = ~n6022 & n6030;
  assign n6032 = ~n6018 & n6031;
  assign n6033 = ~n6013 & ~n6032;
  assign n6034 = n5919 & ~n6025;
  assign n6035 = n5985 & n6034;
  assign n6036 = ~n5867 & n6035;
  assign n6037 = ~n5840 & n6036;
  assign n6038 = n67 & ~n5574;
  assign n6039 = ~n6008 & ~n6038;
  assign n6040 = n6000 & n6039;
  assign n6041 = ~n5990 & n6040;
  assign n6042 = ~n5984 & n6039;
  assign n6043 = ~n6025 & ~n6042;
  assign n6044 = ~n6041 & n6043;
  assign n6045 = ~n6037 & ~n6044;
  assign n6046 = pi03 & ~n5607;
  assign n6047 = ~n5604 & n6046;
  assign n6048 = ~n5597 & n6047;
  assign n6049 = ~n5620 & ~n6048;
  assign n6050 = ~n2619 & ~n6049;
  assign n6051 = n2619 & ~n6048;
  assign n6052 = ~n5620 & n6051;
  assign n6053 = ~n6050 & ~n6052;
  assign n6054 = ~pi05 & ~n6053;
  assign n6055 = pi05 & ~n6052;
  assign n6056 = ~n6050 & n6055;
  assign n6057 = ~n6054 & ~n6056;
  assign n6058 = ~n6045 & ~n6057;
  assign n6059 = ~n5557 & n5588;
  assign n6060 = n5249 & ~n5555;
  assign n6061 = ~n5554 & n6060;
  assign n6062 = ~n5535 & n6061;
  assign n6063 = ~n6059 & ~n6062;
  assign n6064 = ~pi05 & ~n6063;
  assign n6065 = pi05 & ~n6062;
  assign n6066 = ~n6059 & n6065;
  assign n6067 = ~n6064 & ~n6066;
  assign n6068 = ~n5610 & ~n5619;
  assign n6069 = ~n5620 & n6068;
  assign n6070 = ~n6067 & ~n6069;
  assign n6071 = ~n5620 & ~n6066;
  assign n6072 = n6068 & n6071;
  assign n6073 = ~n6064 & n6072;
  assign n6074 = ~pi07 & ~n6073;
  assign n6075 = ~n6070 & n6074;
  assign n6076 = ~n6070 & ~n6073;
  assign n6077 = pi07 & ~n6076;
  assign n6078 = ~n6075 & ~n6077;
  assign n6079 = ~n6045 & ~n6078;
  assign n6080 = ~pi07 & ~n6062;
  assign n6081 = ~n6059 & n6080;
  assign n6082 = pi07 & ~n6063;
  assign n6083 = ~n6081 & ~n6082;
  assign n6084 = ~n6044 & ~n6083;
  assign n6085 = ~n6037 & n6084;
  assign n6086 = ~pi05 & ~n5618;
  assign n6087 = pi05 & ~n5607;
  assign n6088 = ~n5604 & n6087;
  assign n6089 = ~n5597 & n6088;
  assign n6090 = ~n6086 & ~n6089;
  assign n6091 = ~n6044 & ~n6090;
  assign n6092 = ~n6037 & n6091;
  assign n6093 = ~n6085 & ~n6092;
  assign n6094 = ~n6079 & n6093;
  assign n6095 = ~n6058 & n6094;
  assign n6096 = ~n6033 & n6095;
  assign n6097 = ~n6044 & n6086;
  assign n6098 = ~n6037 & n6097;
  assign n6099 = ~n6045 & n6054;
  assign n6100 = ~n6098 & ~n6099;
  assign n6101 = ~n6079 & ~n6085;
  assign n6102 = ~n6100 & n6101;
  assign n6103 = ~n6045 & n6075;
  assign n6104 = ~n5651 & ~n5686;
  assign n6105 = ~n5628 & ~n5656;
  assign n6106 = ~n5622 & n6105;
  assign n6107 = ~n6104 & ~n6106;
  assign n6108 = ~n5628 & ~n5651;
  assign n6109 = ~n5686 & n6108;
  assign n6110 = ~n5656 & n6109;
  assign n6111 = ~n5622 & n6110;
  assign n6112 = ~pi09 & ~n6111;
  assign n6113 = ~n6107 & n6112;
  assign n6114 = ~n6045 & n6113;
  assign n6115 = ~n5557 & ~n5683;
  assign n6116 = ~n5555 & ~n5646;
  assign n6117 = ~n5554 & n6116;
  assign n6118 = ~n5535 & n6117;
  assign n6119 = ~pi09 & ~n6118;
  assign n6120 = ~n6115 & n6119;
  assign n6121 = ~n6044 & n6120;
  assign n6122 = ~n6037 & n6121;
  assign n6123 = ~n6044 & n6081;
  assign n6124 = ~n6037 & n6123;
  assign n6125 = ~n6122 & ~n6124;
  assign n6126 = ~n6114 & n6125;
  assign n6127 = ~n6103 & n6126;
  assign n6128 = ~n6102 & n6127;
  assign n6129 = ~n6096 & n6128;
  assign n6130 = ~n5557 & ~n5667;
  assign n6131 = ~n5555 & ~n5635;
  assign n6132 = ~n5554 & n6131;
  assign n6133 = ~n5535 & n6132;
  assign n6134 = ~pi11 & ~n6133;
  assign n6135 = ~n6130 & n6134;
  assign n6136 = ~n6130 & ~n6133;
  assign n6137 = pi11 & ~n6136;
  assign n6138 = ~n6135 & ~n6137;
  assign n6139 = ~n6044 & ~n6138;
  assign n6140 = ~n6037 & n6139;
  assign n6141 = ~n5557 & ~n5858;
  assign n6142 = ~n5555 & ~n5845;
  assign n6143 = ~n5554 & n6142;
  assign n6144 = ~n5535 & n6143;
  assign n6145 = ~pi13 & ~n6144;
  assign n6146 = ~n6141 & n6145;
  assign n6147 = ~n6141 & ~n6144;
  assign n6148 = pi13 & ~n6147;
  assign n6149 = ~n6146 & ~n6148;
  assign n6150 = ~n6044 & ~n6149;
  assign n6151 = ~n6037 & n6150;
  assign n6152 = ~n6115 & ~n6118;
  assign n6153 = pi09 & ~n6152;
  assign n6154 = ~n6044 & n6153;
  assign n6155 = ~n6037 & n6154;
  assign n6156 = ~n6151 & ~n6155;
  assign n6157 = ~n6140 & n6156;
  assign n6158 = n5835 & ~n5836;
  assign n6159 = ~n5837 & ~n6158;
  assign n6160 = ~n6111 & n6159;
  assign n6161 = ~n5836 & n6110;
  assign n6162 = ~n5622 & n6161;
  assign n6163 = ~n6160 & ~n6162;
  assign n6164 = ~pi11 & ~n6163;
  assign n6165 = pi11 & ~n6162;
  assign n6166 = ~n6160 & n6165;
  assign n6167 = ~n6164 & ~n6166;
  assign n6168 = ~n6045 & ~n6167;
  assign n6169 = ~n5712 & ~n5760;
  assign n6170 = ~n5837 & n6169;
  assign n6171 = ~n5690 & n6170;
  assign n6172 = ~pi11 & ~n6147;
  assign n6173 = pi11 & ~n6144;
  assign n6174 = ~n6141 & n6173;
  assign n6175 = ~n6172 & ~n6174;
  assign n6176 = ~pi13 & ~n6175;
  assign n6177 = pi13 & ~n6174;
  assign n6178 = ~n6172 & n6177;
  assign n6179 = ~n6176 & ~n6178;
  assign n6180 = ~n6171 & ~n6179;
  assign n6181 = n6170 & ~n6178;
  assign n6182 = ~n5690 & n6181;
  assign n6183 = ~n6176 & n6182;
  assign n6184 = ~n6180 & ~n6183;
  assign n6185 = ~n6045 & n6184;
  assign n6186 = ~n6107 & ~n6111;
  assign n6187 = pi09 & ~n6186;
  assign n6188 = ~n6045 & n6187;
  assign n6189 = ~n6185 & ~n6188;
  assign n6190 = ~n6168 & n6189;
  assign n6191 = n6157 & n6190;
  assign n6192 = ~n6129 & n6191;
  assign n6193 = ~n6041 & ~n6042;
  assign n6194 = ~n5988 & ~n6193;
  assign n6195 = ~n5699 & ~n5739;
  assign n6196 = ~n5830 & n6195;
  assign n6197 = ~n5863 & n6196;
  assign n6198 = ~n5699 & ~n5712;
  assign n6199 = ~n5720 & n6198;
  assign n6200 = ~n5739 & ~n5760;
  assign n6201 = ~n5767 & n6200;
  assign n6202 = n6199 & n6201;
  assign n6203 = n5838 & n6202;
  assign n6204 = ~n5690 & n6203;
  assign n6205 = ~n6197 & ~n6204;
  assign n6206 = ~n5557 & n5756;
  assign n6207 = ~n5555 & ~n5912;
  assign n6208 = ~n5554 & n6207;
  assign n6209 = ~n5535 & n6208;
  assign n6210 = ~n6206 & ~n6209;
  assign n6211 = ~pi17 & ~n6210;
  assign n6212 = pi17 & ~n6209;
  assign n6213 = ~n6206 & n6212;
  assign n6214 = ~n6211 & ~n6213;
  assign n6215 = ~n6025 & ~n6214;
  assign n6216 = ~n6205 & n6215;
  assign n6217 = ~n6025 & n6214;
  assign n6218 = ~n6197 & n6217;
  assign n6219 = ~n6204 & n6218;
  assign n6220 = ~n6216 & ~n6219;
  assign n6221 = ~n6194 & ~n6220;
  assign n6222 = ~n5573 & n6210;
  assign n6223 = ~n6024 & n6222;
  assign n6224 = ~n6038 & n6210;
  assign n6225 = ~n6008 & n6224;
  assign n6226 = ~n6002 & n6225;
  assign n6227 = ~n5988 & n6226;
  assign n6228 = ~n6223 & ~n6227;
  assign n6229 = ~n6221 & n6228;
  assign n6230 = ~pi19 & ~n6229;
  assign n6231 = pi19 & ~n6223;
  assign n6232 = ~n6227 & n6231;
  assign n6233 = ~n6221 & n6232;
  assign n6234 = ~n5712 & ~n5790;
  assign n6235 = ~n5720 & n6234;
  assign n6236 = ~n5760 & ~n5782;
  assign n6237 = ~n5767 & n6236;
  assign n6238 = n6235 & n6237;
  assign n6239 = ~n5837 & n6238;
  assign n6240 = ~n5690 & n6239;
  assign n6241 = ~n5849 & ~n5855;
  assign n6242 = ~n5860 & n6241;
  assign n6243 = ~n5844 & n6242;
  assign n6244 = n5791 & ~n6243;
  assign n6245 = n5829 & ~n6244;
  assign n6246 = ~n6240 & n6245;
  assign n6247 = ~n6240 & ~n6244;
  assign n6248 = ~n5829 & ~n6247;
  assign n6249 = ~n6246 & ~n6248;
  assign n6250 = ~n6045 & ~n6249;
  assign n6251 = ~n5555 & n5740;
  assign n6252 = ~n5554 & n6251;
  assign n6253 = ~n5535 & n6252;
  assign n6254 = n5728 & n5733;
  assign n6255 = ~n5727 & n6254;
  assign n6256 = ~n5728 & ~n5734;
  assign n6257 = ~n6255 & ~n6256;
  assign n6258 = ~n5557 & n6257;
  assign n6259 = ~n6253 & ~n6258;
  assign n6260 = ~n6044 & n6259;
  assign n6261 = ~n6037 & n6260;
  assign n6262 = ~pi17 & ~n6261;
  assign n6263 = ~n6250 & n6262;
  assign n6264 = ~n6233 & n6263;
  assign n6265 = ~n6230 & n6264;
  assign n6266 = ~n5867 & n5917;
  assign n6267 = ~n5840 & n6266;
  assign n6268 = ~n5907 & ~n5921;
  assign n6269 = ~n6267 & n6268;
  assign n6270 = n5917 & ~n6268;
  assign n6271 = ~n5867 & n6270;
  assign n6272 = ~n5840 & n6271;
  assign n6273 = ~n6269 & ~n6272;
  assign n6274 = ~n6045 & n6273;
  assign n6275 = n5920 & ~n6044;
  assign n6276 = ~n6037 & n6275;
  assign n6277 = ~pi21 & ~n6276;
  assign n6278 = ~n6274 & n6277;
  assign n6279 = ~n5844 & ~n5855;
  assign n6280 = ~n5849 & ~n5860;
  assign n6281 = ~n6279 & ~n6280;
  assign n6282 = ~n5712 & ~n5849;
  assign n6283 = ~n5720 & n6282;
  assign n6284 = ~n5760 & ~n5860;
  assign n6285 = ~n5767 & n6284;
  assign n6286 = n6283 & n6285;
  assign n6287 = ~n5837 & ~n6243;
  assign n6288 = n6286 & n6287;
  assign n6289 = ~n6281 & n6288;
  assign n6290 = ~n5690 & n6289;
  assign n6291 = ~n6243 & ~n6281;
  assign n6292 = ~n5837 & n6286;
  assign n6293 = ~n5690 & n6292;
  assign n6294 = ~n6291 & ~n6293;
  assign n6295 = ~pi15 & ~n6294;
  assign n6296 = ~n6290 & n6295;
  assign n6297 = ~n6045 & n6296;
  assign n6298 = ~n6171 & ~n6175;
  assign n6299 = n6169 & ~n6174;
  assign n6300 = ~n5837 & n6299;
  assign n6301 = ~n6172 & n6300;
  assign n6302 = ~n5690 & n6301;
  assign n6303 = ~pi13 & ~n6302;
  assign n6304 = ~n6298 & n6303;
  assign n6305 = ~n6045 & n6304;
  assign n6306 = ~n6044 & n6146;
  assign n6307 = ~n6037 & n6306;
  assign n6308 = ~n5557 & ~n5841;
  assign n6309 = ~n5555 & ~n5850;
  assign n6310 = ~n5554 & n6309;
  assign n6311 = ~n5535 & n6310;
  assign n6312 = ~pi15 & ~n6311;
  assign n6313 = ~n6308 & n6312;
  assign n6314 = ~n6044 & n6313;
  assign n6315 = ~n6037 & n6314;
  assign n6316 = ~n6307 & ~n6315;
  assign n6317 = ~n6305 & n6316;
  assign n6318 = ~n6297 & n6317;
  assign n6319 = ~n6278 & n6318;
  assign n6320 = ~n6044 & n6135;
  assign n6321 = ~n6037 & n6320;
  assign n6322 = ~n6045 & n6164;
  assign n6323 = ~n6321 & ~n6322;
  assign n6324 = ~n6151 & ~n6185;
  assign n6325 = ~n6323 & n6324;
  assign n6326 = ~n6230 & ~n6325;
  assign n6327 = n6319 & n6326;
  assign n6328 = ~n6265 & n6327;
  assign n6329 = ~n6192 & n6328;
  assign n6330 = ~n6250 & ~n6261;
  assign n6331 = ~pi17 & ~n6330;
  assign n6332 = pi17 & ~n6261;
  assign n6333 = ~n6250 & n6332;
  assign n6334 = ~n6331 & ~n6333;
  assign n6335 = ~n6308 & ~n6311;
  assign n6336 = pi15 & ~n6335;
  assign n6337 = ~n6044 & n6336;
  assign n6338 = ~n6037 & n6337;
  assign n6339 = ~n6290 & ~n6294;
  assign n6340 = pi15 & ~n6339;
  assign n6341 = ~n6045 & n6340;
  assign n6342 = ~n6338 & ~n6341;
  assign n6343 = ~n6233 & n6342;
  assign n6344 = ~n6230 & n6343;
  assign n6345 = ~n6334 & n6344;
  assign n6346 = ~n6230 & ~n6278;
  assign n6347 = ~n6265 & n6346;
  assign n6348 = ~n6345 & n6347;
  assign n6349 = ~n6274 & ~n6276;
  assign n6350 = pi21 & ~n6349;
  assign n6351 = n5919 & n5924;
  assign n6352 = ~n5867 & n6351;
  assign n6353 = ~n5840 & n6352;
  assign n6354 = n6001 & ~n6353;
  assign n6355 = ~n5557 & ~n5979;
  assign n6356 = ~n5977 & n6355;
  assign n6357 = n5970 & ~n6356;
  assign n6358 = ~n5965 & ~n6357;
  assign n6359 = n5965 & n6357;
  assign n6360 = ~n6358 & ~n6359;
  assign n6361 = ~n6354 & n6360;
  assign n6362 = ~n5965 & n6000;
  assign n6363 = ~n5990 & n6362;
  assign n6364 = ~n6353 & n6363;
  assign n6365 = ~n6361 & ~n6364;
  assign n6366 = ~n6045 & ~n6365;
  assign n6367 = ~n6003 & ~n6006;
  assign n6368 = ~n6044 & n6367;
  assign n6369 = ~n6037 & n6368;
  assign n6370 = pi27 & ~n6369;
  assign n6371 = ~n6366 & n6370;
  assign n6372 = ~n5993 & ~n5998;
  assign n6373 = ~n6357 & n6372;
  assign n6374 = ~n5881 & ~n6373;
  assign n6375 = ~n5990 & n6374;
  assign n6376 = ~n6353 & n6375;
  assign n6377 = ~n5881 & ~n5990;
  assign n6378 = ~n6353 & n6377;
  assign n6379 = n6373 & ~n6378;
  assign n6380 = ~n6376 & ~n6379;
  assign n6381 = ~n5969 & ~n6356;
  assign n6382 = ~pi25 & ~n6381;
  assign n6383 = pi25 & ~n5969;
  assign n6384 = ~n6356 & n6383;
  assign n6385 = ~n6382 & ~n6384;
  assign n6386 = ~n6044 & n6385;
  assign n6387 = ~n6037 & n6386;
  assign n6388 = ~pi25 & ~n6025;
  assign n6389 = ~n6042 & n6388;
  assign n6390 = ~n6041 & n6389;
  assign n6391 = ~pi25 & ~n5916;
  assign n6392 = ~n5911 & n6391;
  assign n6393 = ~n5907 & n6392;
  assign n6394 = ~n5881 & n6393;
  assign n6395 = ~n6025 & n6394;
  assign n6396 = n5985 & n6395;
  assign n6397 = ~n5867 & n6396;
  assign n6398 = ~n5840 & n6397;
  assign n6399 = ~n6390 & ~n6398;
  assign n6400 = ~n6387 & n6399;
  assign n6401 = ~n6380 & n6400;
  assign n6402 = ~pi31 & ~n6401;
  assign n6403 = ~n6371 & n6402;
  assign n6404 = ~n6350 & n6403;
  assign n6405 = ~pi25 & ~n6006;
  assign n6406 = ~n6003 & n6405;
  assign n6407 = ~n6358 & ~n6406;
  assign n6408 = n6000 & ~n6406;
  assign n6409 = ~n5990 & n6408;
  assign n6410 = ~n6353 & n6409;
  assign n6411 = ~n6407 & ~n6410;
  assign n6412 = ~n5574 & ~n6044;
  assign n6413 = ~n6037 & n6412;
  assign n6414 = ~pi29 & ~n6413;
  assign n6415 = ~n6411 & n6414;
  assign n6416 = ~n5573 & ~n5881;
  assign n6417 = n5918 & n6416;
  assign n6418 = n5924 & n6417;
  assign n6419 = ~n6025 & n6418;
  assign n6420 = ~n5575 & n5984;
  assign n6421 = ~n5867 & n6420;
  assign n6422 = n6419 & n6421;
  assign n6423 = ~n5840 & n6422;
  assign n6424 = n5576 & ~n6025;
  assign n6425 = ~n6042 & n6424;
  assign n6426 = ~n6041 & n6425;
  assign n6427 = ~n6423 & ~n6426;
  assign n6428 = pi29 & ~n6407;
  assign n6429 = ~n6410 & n6428;
  assign n6430 = ~n6427 & n6429;
  assign n6431 = pi29 & ~n5574;
  assign n6432 = ~n6044 & n6431;
  assign n6433 = ~n6037 & n6432;
  assign n6434 = ~pi29 & ~n6426;
  assign n6435 = ~n6423 & n6434;
  assign n6436 = ~n6413 & n6435;
  assign n6437 = ~n6433 & ~n6436;
  assign n6438 = ~n6430 & n6437;
  assign n6439 = ~n6415 & n6438;
  assign n6440 = ~n5881 & ~n5923;
  assign n6441 = ~n6025 & n6440;
  assign n6442 = pi23 & ~n5916;
  assign n6443 = ~n5911 & n6442;
  assign n6444 = ~n5907 & n6443;
  assign n6445 = ~n5921 & n6444;
  assign n6446 = n5984 & n6445;
  assign n6447 = n6441 & n6446;
  assign n6448 = ~n5867 & n6447;
  assign n6449 = ~n5840 & n6448;
  assign n6450 = n5918 & ~n5921;
  assign n6451 = ~n5867 & n6450;
  assign n6452 = ~n5840 & n6451;
  assign n6453 = ~n5921 & ~n6440;
  assign n6454 = ~n6452 & n6453;
  assign n6455 = pi23 & ~n6025;
  assign n6456 = ~n6042 & n6455;
  assign n6457 = ~n6041 & n6456;
  assign n6458 = ~n6454 & ~n6457;
  assign n6459 = ~n6449 & n6458;
  assign n6460 = ~n5921 & ~n6452;
  assign n6461 = n6440 & ~n6460;
  assign n6462 = ~pi23 & ~n5879;
  assign n6463 = ~n5876 & n6462;
  assign n6464 = pi23 & ~n5922;
  assign n6465 = ~n6463 & ~n6464;
  assign n6466 = ~n6044 & n6465;
  assign n6467 = ~n6037 & n6466;
  assign n6468 = ~n6461 & ~n6467;
  assign n6469 = n6459 & n6468;
  assign n6470 = pi25 & ~n5916;
  assign n6471 = ~n5911 & n6470;
  assign n6472 = ~n5907 & n6471;
  assign n6473 = ~n5881 & n6472;
  assign n6474 = ~n6025 & n6473;
  assign n6475 = n5985 & n6474;
  assign n6476 = ~n5867 & n6475;
  assign n6477 = ~n5840 & n6476;
  assign n6478 = pi25 & ~n6025;
  assign n6479 = ~n6042 & n6478;
  assign n6480 = ~n6041 & n6479;
  assign n6481 = ~n6376 & ~n6480;
  assign n6482 = ~n6477 & n6481;
  assign n6483 = ~n6379 & ~n6387;
  assign n6484 = n6482 & n6483;
  assign n6485 = ~n6454 & ~n6461;
  assign n6486 = ~pi23 & ~n6025;
  assign n6487 = ~n6042 & n6486;
  assign n6488 = ~n6041 & n6487;
  assign n6489 = ~pi23 & ~n5916;
  assign n6490 = ~n5911 & n6489;
  assign n6491 = ~n5907 & n6490;
  assign n6492 = ~n5921 & n6491;
  assign n6493 = n5984 & n6492;
  assign n6494 = n6441 & n6493;
  assign n6495 = ~n5867 & n6494;
  assign n6496 = ~n5840 & n6495;
  assign n6497 = ~n6488 & ~n6496;
  assign n6498 = ~n6467 & n6497;
  assign n6499 = ~n6485 & n6498;
  assign n6500 = ~n6484 & ~n6499;
  assign n6501 = ~n6469 & n6500;
  assign n6502 = ~n6439 & n6501;
  assign n6503 = n6404 & n6502;
  assign n6504 = ~n6348 & n6503;
  assign n6505 = ~n6329 & n6504;
  assign n6506 = ~n6366 & ~n6369;
  assign n6507 = ~pi27 & ~n6506;
  assign n6508 = ~n5922 & ~n6044;
  assign n6509 = ~n6037 & n6508;
  assign n6510 = ~pi23 & ~n6509;
  assign n6511 = ~n6401 & n6510;
  assign n6512 = ~n6045 & ~n6485;
  assign n6513 = ~n6484 & ~n6512;
  assign n6514 = n6511 & n6513;
  assign n6515 = ~n6045 & ~n6380;
  assign n6516 = ~n6044 & n6381;
  assign n6517 = ~n6037 & n6516;
  assign n6518 = ~pi25 & ~n6517;
  assign n6519 = ~n6515 & n6518;
  assign n6520 = ~n6514 & ~n6519;
  assign n6521 = ~n6507 & n6520;
  assign n6522 = ~pi31 & ~n6371;
  assign n6523 = ~n6439 & n6522;
  assign n6524 = ~n6521 & n6523;
  assign n6525 = n6411 & ~n6427;
  assign n6526 = ~n6413 & ~n6525;
  assign n6527 = n65 & ~n6526;
  assign n6528 = ~n6524 & ~n6527;
  assign n6529 = ~n6505 & n6528;
  assign n6530 = ~n6469 & ~n6499;
  assign n6531 = ~n6350 & n6530;
  assign n6532 = ~n6348 & n6531;
  assign n6533 = ~n6329 & n6532;
  assign n6534 = ~n6348 & ~n6350;
  assign n6535 = ~n6329 & n6534;
  assign n6536 = ~n6530 & ~n6535;
  assign n6537 = ~n6533 & ~n6536;
  assign n6538 = ~n6529 & ~n6537;
  assign n6539 = ~n6509 & ~n6512;
  assign n6540 = ~n6527 & ~n6539;
  assign n6541 = ~n6524 & n6540;
  assign n6542 = ~n6505 & n6541;
  assign n6543 = ~n6538 & ~n6542;
  assign n6544 = ~n6264 & n6318;
  assign n6545 = n6326 & n6544;
  assign n6546 = ~n6192 & n6545;
  assign n6547 = ~pi21 & ~n6349;
  assign n6548 = pi21 & ~n6276;
  assign n6549 = ~n6274 & n6548;
  assign n6550 = ~n6547 & ~n6549;
  assign n6551 = ~n6230 & ~n6264;
  assign n6552 = ~n6345 & n6551;
  assign n6553 = ~n6550 & ~n6552;
  assign n6554 = ~n6546 & n6553;
  assign n6555 = ~n6230 & ~n6549;
  assign n6556 = ~n6264 & ~n6547;
  assign n6557 = n6555 & n6556;
  assign n6558 = ~n6345 & n6557;
  assign n6559 = ~n6325 & ~n6547;
  assign n6560 = n6544 & n6559;
  assign n6561 = n6555 & n6560;
  assign n6562 = ~n6192 & n6561;
  assign n6563 = ~n6558 & ~n6562;
  assign n6564 = ~n6554 & n6563;
  assign n6565 = ~n6529 & n6564;
  assign n6566 = n6349 & ~n6527;
  assign n6567 = ~n6524 & n6566;
  assign n6568 = ~n6505 & n6567;
  assign n6569 = pi23 & ~n6568;
  assign n6570 = ~n6565 & n6569;
  assign n6571 = ~pi25 & ~n6570;
  assign n6572 = ~n6543 & n6571;
  assign n6573 = pi25 & ~n6542;
  assign n6574 = ~n6538 & n6573;
  assign n6575 = ~n6570 & n6574;
  assign n6576 = ~n6572 & ~n6575;
  assign n6577 = ~n6330 & ~n6527;
  assign n6578 = ~n6524 & n6577;
  assign n6579 = ~n6505 & n6578;
  assign n6580 = ~n6140 & ~n6338;
  assign n6581 = n6156 & n6580;
  assign n6582 = ~n6168 & ~n6341;
  assign n6583 = n6189 & n6582;
  assign n6584 = n6581 & n6583;
  assign n6585 = ~n6129 & n6584;
  assign n6586 = n6318 & ~n6325;
  assign n6587 = n6342 & ~n6586;
  assign n6588 = n6334 & ~n6587;
  assign n6589 = ~n6585 & n6588;
  assign n6590 = ~n6585 & ~n6587;
  assign n6591 = ~n6334 & ~n6590;
  assign n6592 = ~n6589 & ~n6591;
  assign n6593 = ~n6529 & ~n6592;
  assign n6594 = ~n6579 & ~n6593;
  assign n6595 = pi19 & ~n6594;
  assign n6596 = ~n6401 & ~n6484;
  assign n6597 = n6510 & ~n6512;
  assign n6598 = ~n6533 & ~n6597;
  assign n6599 = n6596 & ~n6598;
  assign n6600 = ~n6596 & ~n6597;
  assign n6601 = ~n6533 & n6600;
  assign n6602 = ~pi27 & ~n6529;
  assign n6603 = ~n6601 & n6602;
  assign n6604 = ~n6599 & n6603;
  assign n6605 = ~n6305 & ~n6307;
  assign n6606 = ~n6325 & n6605;
  assign n6607 = ~n6315 & ~n6338;
  assign n6608 = ~n6297 & n6607;
  assign n6609 = ~n6341 & n6608;
  assign n6610 = n6606 & ~n6609;
  assign n6611 = ~n6192 & n6610;
  assign n6612 = ~n6192 & n6606;
  assign n6613 = n6609 & ~n6612;
  assign n6614 = ~n6611 & ~n6613;
  assign n6615 = ~n6529 & ~n6614;
  assign n6616 = ~n6044 & ~n6335;
  assign n6617 = ~n6037 & n6616;
  assign n6618 = ~n6045 & ~n6339;
  assign n6619 = ~n6617 & ~n6618;
  assign n6620 = ~n6527 & ~n6619;
  assign n6621 = ~n6524 & n6620;
  assign n6622 = ~n6505 & n6621;
  assign n6623 = ~n6615 & ~n6622;
  assign n6624 = pi17 & ~n6623;
  assign n6625 = ~n6604 & ~n6624;
  assign n6626 = ~n6595 & n6625;
  assign n6627 = ~n6229 & ~n6527;
  assign n6628 = ~n6524 & n6627;
  assign n6629 = ~n6505 & n6628;
  assign n6630 = ~n6263 & ~n6333;
  assign n6631 = ~n6331 & n6630;
  assign n6632 = ~n6230 & ~n6233;
  assign n6633 = ~n6631 & n6632;
  assign n6634 = n6631 & ~n6632;
  assign n6635 = ~n6633 & ~n6634;
  assign n6636 = ~n6590 & n6635;
  assign n6637 = ~n6233 & ~n6263;
  assign n6638 = ~n6230 & n6637;
  assign n6639 = n6263 & ~n6632;
  assign n6640 = ~n6638 & ~n6639;
  assign n6641 = n6590 & ~n6640;
  assign n6642 = ~n6636 & ~n6641;
  assign n6643 = ~n6529 & ~n6642;
  assign n6644 = ~n6629 & ~n6643;
  assign n6645 = pi21 & ~n6644;
  assign n6646 = ~pi21 & ~n6629;
  assign n6647 = ~n6643 & n6646;
  assign n6648 = ~n6645 & ~n6647;
  assign n6649 = pi27 & ~n6401;
  assign n6650 = ~n6484 & n6649;
  assign n6651 = ~n6598 & n6650;
  assign n6652 = pi27 & ~n6596;
  assign n6653 = ~n6597 & n6652;
  assign n6654 = ~n6533 & n6653;
  assign n6655 = ~n6529 & ~n6654;
  assign n6656 = ~n6651 & n6655;
  assign n6657 = ~n6515 & ~n6517;
  assign n6658 = pi27 & ~n6657;
  assign n6659 = ~pi27 & ~n6517;
  assign n6660 = ~n6515 & n6659;
  assign n6661 = ~n6527 & ~n6660;
  assign n6662 = ~n6658 & n6661;
  assign n6663 = ~n6524 & n6662;
  assign n6664 = ~n6505 & n6663;
  assign n6665 = ~n6656 & ~n6664;
  assign n6666 = ~pi19 & ~n6579;
  assign n6667 = ~n6593 & n6666;
  assign n6668 = ~n6665 & ~n6667;
  assign n6669 = ~n6648 & n6668;
  assign n6670 = n6626 & n6669;
  assign n6671 = ~n6576 & n6670;
  assign n6672 = ~n6044 & ~n6136;
  assign n6673 = ~n6037 & n6672;
  assign n6674 = ~n6045 & n6163;
  assign n6675 = ~n6673 & ~n6674;
  assign n6676 = ~n6527 & ~n6675;
  assign n6677 = ~n6524 & n6676;
  assign n6678 = ~n6505 & n6677;
  assign n6679 = ~n6140 & ~n6155;
  assign n6680 = ~n6188 & n6679;
  assign n6681 = ~n6168 & n6680;
  assign n6682 = ~n6129 & n6681;
  assign n6683 = ~n6140 & ~n6168;
  assign n6684 = ~n6155 & ~n6188;
  assign n6685 = ~n6129 & n6684;
  assign n6686 = ~n6683 & ~n6685;
  assign n6687 = ~n6682 & ~n6686;
  assign n6688 = ~n6529 & ~n6687;
  assign n6689 = ~n6678 & ~n6688;
  assign n6690 = pi13 & ~n6689;
  assign n6691 = ~n6045 & ~n6186;
  assign n6692 = ~n6044 & ~n6152;
  assign n6693 = ~n6037 & n6692;
  assign n6694 = ~n6691 & ~n6693;
  assign n6695 = ~n6527 & ~n6694;
  assign n6696 = ~n6524 & n6695;
  assign n6697 = ~n6505 & n6696;
  assign n6698 = ~n6122 & ~n6155;
  assign n6699 = ~n6114 & n6698;
  assign n6700 = ~n6188 & n6699;
  assign n6701 = ~n6103 & ~n6124;
  assign n6702 = ~n6102 & n6701;
  assign n6703 = ~n6700 & n6702;
  assign n6704 = ~n6096 & n6703;
  assign n6705 = ~n6096 & n6702;
  assign n6706 = n6700 & ~n6705;
  assign n6707 = ~n6704 & ~n6706;
  assign n6708 = ~n6529 & ~n6707;
  assign n6709 = ~n6697 & ~n6708;
  assign n6710 = pi11 & ~n6709;
  assign n6711 = ~pi13 & ~n6678;
  assign n6712 = ~n6688 & n6711;
  assign n6713 = ~n6298 & ~n6302;
  assign n6714 = ~n6045 & ~n6713;
  assign n6715 = ~n6044 & ~n6147;
  assign n6716 = ~n6037 & n6715;
  assign n6717 = ~pi15 & ~n6716;
  assign n6718 = ~n6714 & n6717;
  assign n6719 = ~n6714 & ~n6716;
  assign n6720 = pi15 & ~n6719;
  assign n6721 = ~n6718 & ~n6720;
  assign n6722 = ~n6527 & ~n6721;
  assign n6723 = ~n6524 & n6722;
  assign n6724 = ~n6505 & n6723;
  assign n6725 = pi15 & ~n6324;
  assign n6726 = ~pi15 & ~n6151;
  assign n6727 = ~n6185 & n6726;
  assign n6728 = n6323 & ~n6727;
  assign n6729 = ~n6725 & n6728;
  assign n6730 = ~n6682 & n6729;
  assign n6731 = n6323 & ~n6682;
  assign n6732 = ~n6725 & ~n6727;
  assign n6733 = ~n6731 & ~n6732;
  assign n6734 = ~n6730 & ~n6733;
  assign n6735 = ~n6529 & n6734;
  assign n6736 = ~n6724 & ~n6735;
  assign n6737 = ~n6712 & n6736;
  assign n6738 = ~n6710 & n6737;
  assign n6739 = ~n6690 & n6738;
  assign n6740 = ~pi13 & ~n6682;
  assign n6741 = ~n6686 & n6740;
  assign n6742 = ~n6529 & n6741;
  assign n6743 = ~pi13 & ~n6673;
  assign n6744 = ~n6674 & n6743;
  assign n6745 = ~n6527 & n6744;
  assign n6746 = ~n6524 & n6745;
  assign n6747 = ~n6505 & n6746;
  assign n6748 = ~n6742 & ~n6747;
  assign n6749 = n6736 & ~n6748;
  assign n6750 = ~pi17 & ~n6307;
  assign n6751 = n6607 & n6750;
  assign n6752 = ~n6297 & ~n6305;
  assign n6753 = ~n6341 & n6752;
  assign n6754 = n6751 & n6753;
  assign n6755 = ~n6325 & n6754;
  assign n6756 = ~n6192 & n6755;
  assign n6757 = ~pi17 & ~n6609;
  assign n6758 = ~n6612 & n6757;
  assign n6759 = ~n6756 & ~n6758;
  assign n6760 = ~n6529 & ~n6759;
  assign n6761 = n6323 & n6727;
  assign n6762 = ~n6682 & n6761;
  assign n6763 = ~pi15 & ~n6324;
  assign n6764 = ~n6731 & n6763;
  assign n6765 = ~n6762 & ~n6764;
  assign n6766 = ~n6529 & ~n6765;
  assign n6767 = ~n6527 & n6718;
  assign n6768 = ~n6524 & n6767;
  assign n6769 = ~n6505 & n6768;
  assign n6770 = ~pi17 & ~n6617;
  assign n6771 = ~n6618 & n6770;
  assign n6772 = ~n6527 & n6771;
  assign n6773 = ~n6524 & n6772;
  assign n6774 = ~n6505 & n6773;
  assign n6775 = ~n6769 & ~n6774;
  assign n6776 = ~n6766 & n6775;
  assign n6777 = ~n6760 & n6776;
  assign n6778 = ~n6749 & n6777;
  assign n6779 = ~n6739 & n6778;
  assign n6780 = pi02 & ~n6527;
  assign n6781 = n65 & n3012;
  assign n6782 = ~n6526 & n6781;
  assign n6783 = ~n3396 & ~n6782;
  assign n6784 = ~n6780 & n6783;
  assign n6785 = ~n6524 & n6784;
  assign n6786 = ~n6505 & n6785;
  assign n6787 = ~n3012 & n3397;
  assign n6788 = ~n6371 & n6787;
  assign n6789 = ~n6439 & n6788;
  assign n6790 = ~n6521 & n6789;
  assign n6791 = ~n6401 & n6787;
  assign n6792 = ~n6371 & n6791;
  assign n6793 = ~n6350 & n6792;
  assign n6794 = n6502 & n6793;
  assign n6795 = ~n6348 & n6794;
  assign n6796 = ~n6329 & n6795;
  assign n6797 = ~n6790 & ~n6796;
  assign n6798 = ~n6786 & n6797;
  assign n6799 = ~pi03 & ~n2993;
  assign n6800 = ~n6798 & n6799;
  assign n6801 = pi03 & ~n2993;
  assign n6802 = ~n6790 & n6801;
  assign n6803 = ~n6796 & n6802;
  assign n6804 = ~n6786 & n6803;
  assign n6805 = ~n6008 & ~n6014;
  assign n6806 = ~n6002 & n6805;
  assign n6807 = ~n5988 & n6806;
  assign n6808 = n6026 & ~n6807;
  assign n6809 = n6012 & ~n6808;
  assign n6810 = ~pi05 & ~n6809;
  assign n6811 = ~n6527 & n6810;
  assign n6812 = ~n6524 & n6811;
  assign n6813 = ~n6505 & n6812;
  assign n6814 = ~n6804 & ~n6813;
  assign n6815 = ~pi03 & ~n6809;
  assign n6816 = pi03 & ~n5580;
  assign n6817 = ~n6011 & n6816;
  assign n6818 = ~n6808 & n6817;
  assign n6819 = ~n6815 & ~n6818;
  assign n6820 = ~n3012 & ~n6819;
  assign n6821 = n3012 & ~n6818;
  assign n6822 = ~n6815 & n6821;
  assign n6823 = ~n6820 & ~n6822;
  assign n6824 = ~pi05 & ~n6823;
  assign n6825 = ~n6529 & n6824;
  assign n6826 = ~pi03 & ~n6790;
  assign n6827 = ~n6796 & n6826;
  assign n6828 = ~n6786 & n6827;
  assign n6829 = ~n6825 & ~n6828;
  assign n6830 = n6814 & n6829;
  assign n6831 = ~n6800 & n6830;
  assign n6832 = ~n6045 & ~n6076;
  assign n6833 = ~n6044 & ~n6063;
  assign n6834 = ~n6037 & n6833;
  assign n6835 = ~pi09 & ~n6834;
  assign n6836 = ~n6832 & n6835;
  assign n6837 = ~n6832 & ~n6834;
  assign n6838 = pi09 & ~n6837;
  assign n6839 = ~n6836 & ~n6838;
  assign n6840 = ~n6527 & ~n6839;
  assign n6841 = ~n6524 & n6840;
  assign n6842 = ~n6505 & n6841;
  assign n6843 = ~n6045 & n6053;
  assign n6844 = n5618 & ~n6044;
  assign n6845 = ~n6037 & n6844;
  assign n6846 = ~pi07 & ~n6845;
  assign n6847 = ~n6843 & n6846;
  assign n6848 = ~n6843 & ~n6845;
  assign n6849 = pi07 & ~n6848;
  assign n6850 = ~n6847 & ~n6849;
  assign n6851 = ~n6527 & ~n6850;
  assign n6852 = ~n6524 & n6851;
  assign n6853 = ~n6505 & n6852;
  assign n6854 = pi05 & ~n5580;
  assign n6855 = ~n6011 & n6854;
  assign n6856 = ~n6808 & n6855;
  assign n6857 = ~n6527 & n6856;
  assign n6858 = ~n6524 & n6857;
  assign n6859 = ~n6505 & n6858;
  assign n6860 = ~n6853 & ~n6859;
  assign n6861 = ~n6842 & n6860;
  assign n6862 = ~n6058 & ~n6092;
  assign n6863 = ~n6033 & n6862;
  assign n6864 = n6100 & ~n6863;
  assign n6865 = n6101 & ~n6864;
  assign n6866 = n6100 & ~n6101;
  assign n6867 = ~n6863 & n6866;
  assign n6868 = ~pi09 & ~n6867;
  assign n6869 = ~n6865 & n6868;
  assign n6870 = ~n6865 & ~n6867;
  assign n6871 = pi09 & ~n6870;
  assign n6872 = ~n6869 & ~n6871;
  assign n6873 = ~n6529 & ~n6872;
  assign n6874 = n6033 & ~n6862;
  assign n6875 = ~pi07 & ~n6863;
  assign n6876 = ~n6874 & n6875;
  assign n6877 = ~n6863 & ~n6874;
  assign n6878 = pi07 & ~n6877;
  assign n6879 = ~n6876 & ~n6878;
  assign n6880 = ~n6529 & ~n6879;
  assign n6881 = pi05 & ~n6822;
  assign n6882 = ~n6820 & n6881;
  assign n6883 = ~n6529 & n6882;
  assign n6884 = ~n6880 & ~n6883;
  assign n6885 = ~n6873 & n6884;
  assign n6886 = n6861 & n6885;
  assign n6887 = ~n6831 & n6886;
  assign n6888 = ~n6527 & n6836;
  assign n6889 = ~n6524 & n6888;
  assign n6890 = ~n6505 & n6889;
  assign n6891 = ~pi11 & ~n6693;
  assign n6892 = ~n6691 & n6891;
  assign n6893 = ~n6527 & n6892;
  assign n6894 = ~n6524 & n6893;
  assign n6895 = ~n6505 & n6894;
  assign n6896 = ~n6890 & ~n6895;
  assign n6897 = n6775 & n6896;
  assign n6898 = ~n6760 & ~n6766;
  assign n6899 = ~n6529 & n6869;
  assign n6900 = ~pi11 & ~n6704;
  assign n6901 = ~n6706 & n6900;
  assign n6902 = ~n6529 & n6901;
  assign n6903 = ~n6899 & ~n6902;
  assign n6904 = n6898 & n6903;
  assign n6905 = n6897 & n6904;
  assign n6906 = ~n6529 & n6876;
  assign n6907 = ~n6527 & n6847;
  assign n6908 = ~n6524 & n6907;
  assign n6909 = ~n6505 & n6908;
  assign n6910 = ~n6906 & ~n6909;
  assign n6911 = ~n6842 & ~n6873;
  assign n6912 = ~n6910 & n6911;
  assign n6913 = ~n6749 & ~n6912;
  assign n6914 = n6905 & n6913;
  assign n6915 = ~n6887 & n6914;
  assign n6916 = ~n6779 & ~n6915;
  assign n6917 = n6671 & n6916;
  assign n6918 = ~n6648 & n6667;
  assign n6919 = ~pi21 & ~n6644;
  assign n6920 = ~n6565 & ~n6568;
  assign n6921 = ~pi23 & ~n6920;
  assign n6922 = ~n6919 & ~n6921;
  assign n6923 = ~n6918 & n6922;
  assign n6924 = ~n6604 & ~n6665;
  assign n6925 = ~n6576 & n6924;
  assign n6926 = ~n6923 & n6925;
  assign n6927 = ~pi25 & ~n6542;
  assign n6928 = ~n6538 & n6927;
  assign n6929 = ~n6665 & n6928;
  assign n6930 = ~n6604 & n6929;
  assign n6931 = ~n6599 & ~n6601;
  assign n6932 = ~n6529 & ~n6931;
  assign n6933 = ~n6527 & ~n6657;
  assign n6934 = ~n6524 & n6933;
  assign n6935 = ~n6505 & n6934;
  assign n6936 = ~pi27 & ~n6935;
  assign n6937 = ~n6932 & n6936;
  assign n6938 = ~n6930 & ~n6937;
  assign n6939 = ~n6926 & n6938;
  assign n6940 = ~n6917 & n6939;
  assign n6941 = n6530 & n6596;
  assign n6942 = ~n6350 & n6941;
  assign n6943 = ~n6348 & n6942;
  assign n6944 = ~n6329 & n6943;
  assign n6945 = n6521 & ~n6944;
  assign n6946 = ~n6371 & n6439;
  assign n6947 = ~n6945 & n6946;
  assign n6948 = ~n6529 & n6947;
  assign n6949 = ~n6526 & ~n6527;
  assign n6950 = ~n6524 & n6949;
  assign n6951 = ~n6505 & n6950;
  assign n6952 = ~pi31 & ~n6951;
  assign n6953 = ~n6948 & n6952;
  assign n6954 = ~n6948 & ~n6951;
  assign n6955 = pi31 & ~n6954;
  assign n6956 = ~n6953 & ~n6955;
  assign n6957 = ~n6371 & ~n6507;
  assign n6958 = n6520 & ~n6957;
  assign n6959 = ~n6944 & n6958;
  assign n6960 = n6520 & ~n6944;
  assign n6961 = n6957 & ~n6960;
  assign n6962 = ~n6959 & ~n6961;
  assign n6963 = n6506 & ~n6527;
  assign n6964 = ~n6524 & n6963;
  assign n6965 = ~n6505 & n6964;
  assign n6966 = pi29 & ~n6965;
  assign n6967 = ~pi29 & ~n6369;
  assign n6968 = ~n6366 & n6967;
  assign n6969 = ~n6527 & n6968;
  assign n6970 = ~n6524 & n6969;
  assign n6971 = ~n6505 & n6970;
  assign n6972 = ~n6529 & ~n6971;
  assign n6973 = ~n6966 & n6972;
  assign n6974 = ~n6962 & n6973;
  assign n6975 = ~n6529 & ~n6962;
  assign n6976 = ~n6966 & ~n6971;
  assign n6977 = ~n6975 & ~n6976;
  assign n6978 = ~n6974 & ~n6977;
  assign n6979 = ~n6956 & ~n6978;
  assign n6980 = ~n6940 & n6979;
  assign n6981 = ~pi29 & ~n6965;
  assign n6982 = ~n6975 & n6981;
  assign n6983 = ~n6956 & n6982;
  assign n6984 = ~pi31 & ~n6954;
  assign n6985 = pi00 & ~n6984;
  assign n6986 = pi00 & ~pi01;
  assign n6987 = ~pi31 & n2993;
  assign n6988 = ~n6954 & n6987;
  assign n6989 = ~n6986 & ~n6988;
  assign n6990 = ~n6985 & n6989;
  assign n6991 = ~n6983 & n6990;
  assign n6992 = ~n6980 & n6991;
  assign n6993 = ~n6980 & ~n6983;
  assign n6994 = ~n2993 & ~n6986;
  assign n6995 = ~n6993 & n6994;
  assign po01 = ~n6992 & ~n6995;
  assign n6997 = ~n6798 & ~n6984;
  assign n6998 = ~n6983 & n6997;
  assign n6999 = ~n6980 & n6998;
  assign n7000 = ~n6983 & ~n6984;
  assign n7001 = ~n6980 & n7000;
  assign n7002 = pi03 & ~n6798;
  assign n7003 = ~n6828 & ~n7002;
  assign n7004 = ~n2993 & ~n7003;
  assign n7005 = n2993 & ~n6828;
  assign n7006 = ~n7002 & n7005;
  assign n7007 = ~n7004 & ~n7006;
  assign n7008 = ~n7001 & n7007;
  assign po03 = ~n6999 & ~n7008;
  assign n7010 = ~n6527 & n6809;
  assign n7011 = ~n6524 & n7010;
  assign n7012 = ~n6505 & n7011;
  assign n7013 = ~n6529 & n6823;
  assign n7014 = ~n7012 & ~n7013;
  assign n7015 = ~n6984 & ~n7014;
  assign n7016 = ~n6983 & n7015;
  assign n7017 = ~n6980 & n7016;
  assign n7018 = ~pi05 & ~n7014;
  assign n7019 = pi05 & ~n7012;
  assign n7020 = ~n7013 & n7019;
  assign n7021 = ~n6804 & ~n6828;
  assign n7022 = ~n6800 & n7021;
  assign n7023 = ~n7020 & n7022;
  assign n7024 = ~n7018 & n7023;
  assign n7025 = ~n7018 & ~n7020;
  assign n7026 = ~n7022 & ~n7025;
  assign n7027 = ~n7024 & ~n7026;
  assign n7028 = ~n7001 & ~n7027;
  assign po05 = ~n7017 & ~n7028;
  assign n7030 = ~n6527 & ~n6848;
  assign n7031 = ~n6524 & n7030;
  assign n7032 = ~n6505 & n7031;
  assign n7033 = ~n6529 & ~n6877;
  assign n7034 = ~n7032 & ~n7033;
  assign n7035 = ~n6984 & ~n7034;
  assign n7036 = ~n6983 & n7035;
  assign n7037 = ~n6980 & n7036;
  assign n7038 = n6860 & ~n6880;
  assign n7039 = ~n6883 & n7038;
  assign n7040 = ~n6831 & n7039;
  assign n7041 = ~n6853 & ~n6880;
  assign n7042 = ~n6859 & ~n6883;
  assign n7043 = ~n6831 & n7042;
  assign n7044 = ~n7041 & ~n7043;
  assign n7045 = ~n7040 & ~n7044;
  assign n7046 = ~n7001 & ~n7045;
  assign po07 = ~n7037 & ~n7046;
  assign n7048 = ~n6527 & ~n6837;
  assign n7049 = ~n6524 & n7048;
  assign n7050 = ~n6505 & n7049;
  assign n7051 = ~n6529 & ~n6870;
  assign n7052 = ~n7050 & ~n7051;
  assign n7053 = ~n6984 & ~n7052;
  assign n7054 = ~n6983 & n7053;
  assign n7055 = ~n6980 & n7054;
  assign n7056 = n6910 & ~n7040;
  assign n7057 = n6911 & ~n7056;
  assign n7058 = n6910 & ~n6911;
  assign n7059 = ~n7040 & n7058;
  assign n7060 = ~n7057 & ~n7059;
  assign n7061 = ~n7001 & ~n7060;
  assign po09 = ~n7055 & ~n7061;
  assign n7063 = ~n6709 & ~n6984;
  assign n7064 = ~n6983 & n7063;
  assign n7065 = ~n6980 & n7064;
  assign n7066 = ~pi11 & ~n6697;
  assign n7067 = ~n6708 & n7066;
  assign n7068 = ~n6710 & ~n7067;
  assign n7069 = ~n6890 & ~n6899;
  assign n7070 = ~n6912 & n7069;
  assign n7071 = ~n7068 & n7070;
  assign n7072 = ~n6887 & n7071;
  assign n7073 = ~n6887 & n7070;
  assign n7074 = n7068 & ~n7073;
  assign n7075 = ~n7072 & ~n7074;
  assign n7076 = ~n7001 & ~n7075;
  assign po11 = ~n7065 & ~n7076;
  assign n7078 = ~n6689 & ~n6984;
  assign n7079 = ~n6983 & n7078;
  assign n7080 = ~n6980 & n7079;
  assign n7081 = n6896 & ~n6899;
  assign n7082 = ~n6902 & n7081;
  assign n7083 = ~n6912 & n7082;
  assign n7084 = ~n6887 & n7083;
  assign n7085 = ~n6710 & ~n6712;
  assign n7086 = ~n6690 & n7085;
  assign n7087 = ~n7084 & n7086;
  assign n7088 = ~n6690 & ~n6712;
  assign n7089 = ~n6710 & ~n7084;
  assign n7090 = ~n7088 & ~n7089;
  assign n7091 = ~n7087 & ~n7090;
  assign n7092 = ~n7001 & ~n7091;
  assign po13 = ~n7080 & ~n7092;
  assign n7094 = ~n6527 & n6719;
  assign n7095 = ~n6524 & n7094;
  assign n7096 = ~n6505 & n7095;
  assign n7097 = n6324 & ~n6731;
  assign n7098 = n6323 & ~n6324;
  assign n7099 = ~n6682 & n7098;
  assign n7100 = ~n7097 & ~n7099;
  assign n7101 = ~n6529 & n7100;
  assign n7102 = ~n7096 & ~n7101;
  assign n7103 = ~n6984 & n7102;
  assign n7104 = ~n6983 & n7103;
  assign n7105 = ~n6980 & n7104;
  assign n7106 = ~n6736 & n6748;
  assign n7107 = ~n7089 & n7106;
  assign n7108 = n6739 & ~n7084;
  assign n7109 = ~n7088 & n7106;
  assign n7110 = ~n6749 & ~n7109;
  assign n7111 = ~n7108 & n7110;
  assign n7112 = ~n7107 & n7111;
  assign n7113 = ~n7001 & ~n7112;
  assign po15 = ~n7105 & ~n7113;
  assign n7115 = ~n6623 & ~n6984;
  assign n7116 = ~n6983 & n7115;
  assign n7117 = ~n6980 & n7116;
  assign n7118 = ~pi17 & ~n6622;
  assign n7119 = ~n6615 & n7118;
  assign n7120 = ~n6624 & ~n7119;
  assign n7121 = ~n6766 & ~n6769;
  assign n7122 = ~n6749 & n7121;
  assign n7123 = ~n7120 & n7122;
  assign n7124 = ~n7108 & n7123;
  assign n7125 = ~n7108 & n7122;
  assign n7126 = n7120 & ~n7125;
  assign n7127 = ~n7124 & ~n7126;
  assign n7128 = ~n7001 & ~n7127;
  assign po17 = ~n7117 & ~n7128;
  assign n7130 = ~n6594 & ~n6984;
  assign n7131 = ~n6983 & n7130;
  assign n7132 = ~n6980 & n7131;
  assign n7133 = ~n6624 & ~n6667;
  assign n7134 = ~n6595 & n7133;
  assign n7135 = ~n6779 & n7134;
  assign n7136 = ~n6915 & n7135;
  assign n7137 = ~n6595 & ~n6667;
  assign n7138 = ~n6624 & ~n6779;
  assign n7139 = ~n6915 & n7138;
  assign n7140 = ~n7137 & ~n7139;
  assign n7141 = ~n7136 & ~n7140;
  assign n7142 = ~n7001 & ~n7141;
  assign po19 = ~n7132 & ~n7142;
  assign n7144 = n6644 & ~n6984;
  assign n7145 = ~n6983 & n7144;
  assign n7146 = ~n6980 & n7145;
  assign n7147 = ~n6648 & n7134;
  assign n7148 = ~n6779 & n7147;
  assign n7149 = ~n6915 & n7148;
  assign n7150 = ~n6647 & ~n6667;
  assign n7151 = ~n6645 & n7150;
  assign n7152 = ~n6918 & ~n7151;
  assign n7153 = ~n7149 & n7152;
  assign n7154 = ~n6595 & ~n6624;
  assign n7155 = n7151 & n7154;
  assign n7156 = ~n6779 & n7155;
  assign n7157 = ~n6915 & n7156;
  assign n7158 = ~n7153 & ~n7157;
  assign n7159 = ~n7001 & n7158;
  assign po21 = ~n7146 & ~n7159;
  assign n7161 = n6920 & ~n6984;
  assign n7162 = ~n6983 & n7161;
  assign n7163 = ~n6980 & n7162;
  assign n7164 = ~n6570 & ~n6921;
  assign n7165 = ~n6919 & ~n7164;
  assign n7166 = ~n6918 & n7165;
  assign n7167 = ~n7149 & n7166;
  assign n7168 = ~n6918 & ~n6919;
  assign n7169 = ~n7149 & n7168;
  assign n7170 = n7164 & ~n7169;
  assign n7171 = ~n7167 & ~n7170;
  assign n7172 = ~n7001 & ~n7171;
  assign po23 = ~n7163 & ~n7172;
  assign n7174 = n6543 & ~n6984;
  assign n7175 = ~n6983 & n7174;
  assign n7176 = ~n6980 & n7175;
  assign n7177 = pi25 & ~n6543;
  assign n7178 = ~n6570 & ~n6928;
  assign n7179 = ~n7177 & n7178;
  assign n7180 = ~n6928 & ~n7177;
  assign n7181 = n6570 & ~n7180;
  assign n7182 = ~n7179 & ~n7181;
  assign n7183 = ~n6919 & n7164;
  assign n7184 = ~n6918 & n7183;
  assign n7185 = ~n7149 & n7184;
  assign n7186 = ~n7182 & ~n7185;
  assign n7187 = n7182 & n7184;
  assign n7188 = ~n7149 & n7187;
  assign n7189 = ~n7186 & ~n7188;
  assign n7190 = ~n7001 & n7189;
  assign po25 = n7176 | n7190;
  assign n7192 = ~n142 & n3734;
  assign n7193 = ~n140 & n7192;
  assign n7194 = ~n133 & n7193;
  assign n7195 = n121 & ~n165;
  assign po26 = n7194 | n7195;
  assign n7197 = n6922 & ~n6928;
  assign n7198 = ~n6918 & n7197;
  assign n7199 = ~n7149 & n7198;
  assign n7200 = ~n6572 & ~n6928;
  assign n7201 = ~n6575 & ~n6924;
  assign n7202 = n7200 & n7201;
  assign n7203 = ~n6575 & n7200;
  assign n7204 = n6924 & ~n7203;
  assign n7205 = ~n7202 & ~n7204;
  assign n7206 = ~n7199 & n7205;
  assign n7207 = n6924 & n7197;
  assign n7208 = ~n6918 & n7207;
  assign n7209 = ~n7149 & n7208;
  assign n7210 = ~n7206 & ~n7209;
  assign n7211 = ~n7001 & n7210;
  assign n7212 = ~n6932 & ~n6935;
  assign n7213 = ~n6984 & ~n7212;
  assign n7214 = ~n6983 & n7213;
  assign n7215 = ~n6980 & n7214;
  assign po27 = ~n7211 & ~n7215;
  assign n7217 = n135 & n259;
  assign po28 = ~n90 & n7217;
  assign n7219 = ~n6965 & ~n6975;
  assign n7220 = ~n6984 & n7219;
  assign n7221 = ~n6983 & n7220;
  assign n7222 = ~n6980 & n7221;
  assign n7223 = ~n6940 & ~n6978;
  assign n7224 = n6938 & n6978;
  assign n7225 = ~n6926 & n7224;
  assign n7226 = ~n6917 & n7225;
  assign n7227 = ~n7223 & ~n7226;
  assign n7228 = ~n7001 & n7227;
  assign po29 = n7222 | n7228;
  assign n7230 = pi01 & ~pi30;
  assign n7231 = n92 & n628;
  assign n7232 = ~n7230 & n7231;
  assign po30 = n203 & n7232;
  assign n7234 = ~n6954 & ~n6984;
  assign n7235 = ~n6983 & n7234;
  assign n7236 = ~n6980 & n7235;
  assign n7237 = ~n6982 & ~n7223;
  assign n7238 = n6984 & ~n7237;
  assign po31 = n7236 | n7238;
endmodule


