//Written by the Majority Logic Package Thu Apr 30 23:01:05 2015
module top (
            pi000, pi001, pi002, pi003, pi004, pi005, pi006, pi007, pi008, pi009, pi010, pi011, pi012, pi013, pi014, pi015, pi016, pi017, pi018, pi019, pi020, pi021, pi022, pi023, pi024, pi025, pi026, pi027, pi028, pi029, pi030, pi031, pi032, pi033, pi034, pi035, pi036, pi037, pi038, pi039, pi040, pi041, pi042, pi043, pi044, pi045, pi046, pi047, pi048, pi049, pi050, pi051, pi052, pi053, pi054, pi055, pi056, pi057, pi058, pi059, pi060, pi061, pi062, pi063, pi064, pi065, pi066, pi067, pi068, pi069, pi070, pi071, pi072, pi073, pi074, pi075, pi076, pi077, pi078, pi079, pi080, pi081, pi082, pi083, pi084, pi085, pi086, pi087, pi088, pi089, pi090, pi091, pi092, pi093, pi094, pi095, pi096, pi097, pi098, pi099, pi100, pi101, pi102, pi103, pi104, pi105, pi106, pi107, pi108, pi109, pi110, pi111, pi112, pi113, pi114, pi115, pi116, pi117, pi118, pi119, pi120, pi121, pi122, pi123, pi124, pi125, pi126, pi127, pi128, pi129, pi130, pi131, pi132, pi133, pi134, pi135, pi136, pi137, pi138, pi139, pi140, pi141, pi142, pi143, pi144, pi145, pi146, pi147, pi148, pi149, pi150, pi151, pi152, pi153, pi154, pi155, pi156, pi157, pi158, pi159, pi160, pi161, pi162, pi163, pi164, pi165, pi166, pi167, pi168, pi169, pi170, pi171, pi172, pi173, pi174, pi175, pi176, pi177, pi178, pi179, pi180, pi181, pi182, pi183, pi184, pi185, pi186, pi187, pi188, pi189, pi190, pi191, pi192, pi193, pi194, pi195, pi196, pi197, pi198, pi199, 
            po0, po1, po2, po3, po4, po5, po6);
input pi000, pi001, pi002, pi003, pi004, pi005, pi006, pi007, pi008, pi009, pi010, pi011, pi012, pi013, pi014, pi015, pi016, pi017, pi018, pi019, pi020, pi021, pi022, pi023, pi024, pi025, pi026, pi027, pi028, pi029, pi030, pi031, pi032, pi033, pi034, pi035, pi036, pi037, pi038, pi039, pi040, pi041, pi042, pi043, pi044, pi045, pi046, pi047, pi048, pi049, pi050, pi051, pi052, pi053, pi054, pi055, pi056, pi057, pi058, pi059, pi060, pi061, pi062, pi063, pi064, pi065, pi066, pi067, pi068, pi069, pi070, pi071, pi072, pi073, pi074, pi075, pi076, pi077, pi078, pi079, pi080, pi081, pi082, pi083, pi084, pi085, pi086, pi087, pi088, pi089, pi090, pi091, pi092, pi093, pi094, pi095, pi096, pi097, pi098, pi099, pi100, pi101, pi102, pi103, pi104, pi105, pi106, pi107, pi108, pi109, pi110, pi111, pi112, pi113, pi114, pi115, pi116, pi117, pi118, pi119, pi120, pi121, pi122, pi123, pi124, pi125, pi126, pi127, pi128, pi129, pi130, pi131, pi132, pi133, pi134, pi135, pi136, pi137, pi138, pi139, pi140, pi141, pi142, pi143, pi144, pi145, pi146, pi147, pi148, pi149, pi150, pi151, pi152, pi153, pi154, pi155, pi156, pi157, pi158, pi159, pi160, pi161, pi162, pi163, pi164, pi165, pi166, pi167, pi168, pi169, pi170, pi171, pi172, pi173, pi174, pi175, pi176, pi177, pi178, pi179, pi180, pi181, pi182, pi183, pi184, pi185, pi186, pi187, pi188, pi189, pi190, pi191, pi192, pi193, pi194, pi195, pi196, pi197, pi198, pi199;
output po0, po1, po2, po3, po4, po5, po6;
wire one, v0, v1, v2, v3, v4, v5, v6, v7, v8, v9, v10, v11, v12, v13, v14, v15, v16, v17, v18, v19, v20, v21, v22, v23, v24, v25, v26, v27, v28, v29, v30, v31, v32, v33, v34, v35, v36, v37, v38, v39, v40, v41, v42, v43, v44, v45, v46, v47, v48, v49, v50, v51, v52, v53, v54, v55, v56, v57, v58, v59, v60, v61, v62, v63, v64, v65, v66, v67, v68, v69, v70, v71, v72, v73, v74, v75, v76, v77, v78, v79, v80, v81, v82, v83, v84, v85, v86, v87, v88, v89, v90, v91, v92, v93, v94, v95, v96, v97, v98, v99, v100, v101, v102, v103, v104, v105, v106, v107, v108, v109, v110, v111, v112, v113, v114, v115, v116, v117, v118, v119, v120, v121, v122, v123, v124, v125, v126, v127, v128, v129, v130, v131, v132, v133, v134, v135, v136, v137, v138, v139, v140, v141, v142, v143, v144, v145, v146, v147, v148, v149, v150, v151, v152, v153, v154, v155, v156, v157, v158, v159, v160, v161, v162, v163, v164, v165, v166, v167, v168, v169, v170, v171, v172, v173, v174, v175, v176, v177, v178, v179, v180, v181, v182, v183, v184, v185, v186, v187, v188, v189, v190, v191, v192, v193, v194, v195, v196, v197, v198, v199, v200, v201, v202, v203, v204, v205, v206, v207, v208, v209, v210, v211, v212, v213, v214, v215, v216, v217, v218, v219, v220, v221, v222, v223, v224, v225, v226, v227, v228, v229, v230, v231, v232, v233, v234, v235, v236, v237, v238, v239, v240, v241, v242, v243, v244, v245, v246, v247, v248, v249, v250, v251, v252, v253, v254, v255, v256, v257, v258, v259, v260, v261, v262, v263, v264, v265, v266, v267, v268, v269, v270, v271, v272, v273, v274, v275, v276, v277, v278, v279, v280, v281, v282, v283, v284, v285, v286, v287, v288, v289, v290, v291, v292, v293, v294, v295, v296, v297, v298, v299, v300, v301, v302, v303, v304, v305, v306, v307, v308, v309, v310, v311, v312, v313, v314, v315, v316, v317, v318, v319, v320, v321, v322, v323, v324, v325, v326, v327, v328, v329, v330, v331, v332, v333, v334, v335, v336, v337, v338, v339, v340, v341, v342, v343, v344, v345, v346, v347, v348, v349, v350, v351, v352, v353, v354, v355, v356, v357, v358, v359, v360, v361, v362, v363, v364, v365, v366, v367, v368, v369, v370, v371, v372, v373, v374, v375, v376, v377, v378, v379, v380, v381, v382, v383, v384, v385, v386, v387, v388, v389, v390, v391, v392, v393, v394, v395, v396, v397, v398, v399, v400, v401, v402, v403, v404, v405, v406, v407, v408, v409, v410, v411, v412, v413, v414, v415, v416, v417, v418, v419, v420, v421, v422, v423, v424, v425, v426, v427, v428, v429, v430, v431, v432, v433, v434, v435, v436, v437, v438, v439, v440, v441, v442, v443, v444, v445, v446, v447, v448, v449, v450, v451, v452, v453, v454, v455, v456, v457, v458, v459, v460, v461, v462, v463, v464, v465, v466, v467, v468, v469, v470, v471, v472, v473, v474, v475, v476, v477, v478, v479, v480, v481, v482, v483, v484, v485, v486, v487, v488, v489, v490, v491, v492, v493, v494, v495, v496, v497, v498, v499, v500, v501, v502, v503, v504, v505, v506, v507, v508, v509, v510, v511, v512, v513, v514, v515, v516, v517, v518, v519, v520, v521, v522, v523, v524, v525, v526, v527, v528, v529, v530, v531, v532, v533, v534, v535, v536, v537, v538, v539, v540, v541, v542, v543, v544, v545, v546, v547, v548, v549, v550, v551, v552, v553, v554, v555, v556, v557, v558, v559, v560, v561, v562, v563, v564, v565, v566, v567, v568, v569, v570, v571, v572, v573, v574, v575, v576, v577, v578, v579, v580, v581, v582, v583, v584, v585, v586, v587, v588, v589, v590, v591, v592, v593, v594, v595, v596, v597, v598, v599, v600, v601, v602, v603, v604, v605, v606, v607, v608, v609, v610, v611, v612, v613, v614, v615, v616, v617, v618, v619, v620, v621, v622, v623, v624, v625, v626, v627, v628, v629, v630, v631, v632, v633, v634, v635, v636, v637, v638, v639, v640, v641, v642, v643, v644, v645, v646, v647, v648, v649, v650, v651, v652, v653, v654, v655, v656, v657, v658, v659, v660, v661, v662, v663, v664, v665, v666, v667, v668, v669, v670, v671, v672, v673, v674, v675, v676, v677, v678, v679, v680, v681, v682, v683, v684, v685, v686, v687, v688, v689, v690, v691, v692, v693, v694, v695, v696, v697, v698, v699, v700, v701, v702, v703, v704, v705, v706, v707, v708, v709, v710, v711, v712, v713, v714, v715, v716, v717, v718, v719, v720, v721, v722, v723, v724, v725, v726, v727, v728, v729, v730, v731, v732, v733, v734, 
w0, w1, w2, w3, w4, w5, w6, w7, w8, w9, w10, w11, w12, w13, w14, w15, w16, w17, w18, w19, w20, w21, w22, w23, w24, w25, w26, w27, w28, w29, w30, w31, w32, w33, w34, w35, w36, w37, w38, w39, w40, w41, w42, w43, w44, w45, w46, w47, w48, w49, w50, w51, w52, w53, w54, w55, w56, w57, w58, w59, w60, w61, w62, w63, w64, w65, w66, w67, w68, w69, w70, w71, w72, w73, w74, w75, w76, w77, w78, w79, w80, w81, w82, w83, w84, w85, w86, w87, w88, w89, w90, w91, w92, w93, w94, w95, w96, w97, w98, w99, w100, w101, w102, w103, w104, w105, w106, w107, w108, w109, w110, w111, w112, w113, w114, w115, w116, w117, w118, w119, w120, w121, w122, w123, w124, w125, w126, w127, w128, w129, w130, w131, w132, w133, w134, w135, w136, w137, w138, w139, w140, w141, w142, w143, w144, w145, w146, w147, w148, w149, w150, w151, w152, w153, w154, w155, w156, w157, w158, w159, w160, w161, w162, w163, w164, w165, w166, w167, w168, w169, w170, w171, w172, w173, w174, w175, w176, w177, w178, w179, w180, w181, w182, w183, w184, w185, w186, w187, w188, w189, w190, w191, w192, w193, w194, w195, w196, w197, w198, w199, w200, w201, w202, w203, w204, w205, w206, w207, w208, w209, w210, w211, w212, w213, w214, w215, w216, w217, w218, w219, w220, w221, w222, w223, w224, w225, w226, w227, w228, w229, w230, w231, w232, w233, w234, w235, w236, w237, w238, w239, w240, w241, w242, w243, w244, w245, w246, w247, w248, w249, w250, w251, w252, w253, w254, w255, w256, w257, w258, w259, w260, w261, w262, w263, w264, w265, w266, w267, w268, w269, w270, w271, w272, w273, w274, w275, w276, w277, w278, w279, w280, w281, w282, w283, w284, w285, w286, w287, w288, w289, w290, w291, w292, w293, w294, w295, w296, w297, w298, w299, w300, w301, w302, w303, w304, w305, w306, w307, w308, w309, w310, w311, w312, w313, w314, w315, w316, w317, w318, w319, w320, w321, w322, w323, w324, w325, w326, w327, w328, w329, w330, w331, w332, w333, w334, w335, w336, w337, w338, w339, w340, w341, w342, w343, w344, w345, w346, w347, w348, w349, w350, w351, w352, w353, w354, w355, w356, w357, w358, w359, w360, w361, w362, w363, w364, w365, w366, w367, w368, w369, w370, w371, w372, w373, w374, w375, w376, w377, w378, w379, w380, w381, w382, w383, w384, w385, w386, w387, w388, w389, w390, w391, w392, w393, w394, w395, w396, w397, w398, w399, w400, w401, w402, w403, w404, w405, w406, w407, w408, w409, w410, w411, w412, w413, w414, w415, w416, w417, w418, w419, w420, w421, w422, w423, w424, w425, w426, w427, w428, w429, w430, w431, w432, w433, w434, w435, w436, w437, w438, w439, w440, w441, w442, w443, w444, w445, w446, w447, w448, w449, w450, w451, w452, w453, w454, w455, w456, w457, w458, w459, w460, w461, w462, w463, w464, w465, w466, w467, w468, w469, w470, w471, w472, w473, w474, w475, w476, w477, w478, w479, w480, w481, w482, w483, w484, w485, w486, w487, w488, w489, w490, w491, w492, w493, w494, w495, w496, w497, w498, w499, w500, w501, w502, w503, w504, w505, w506, w507, w508, w509, w510, w511, w512, w513, w514, w515, w516, w517, w518, w519, w520, w521, w522, w523, w524, w525, w526, w527, w528, w529, w530, w531, w532, w533, w534, w535, w536, w537, w538, w539, w540, w541, w542, w543, w544, w545, w546, w547, w548, w549, w550, w551, w552, w553, w554, w555, w556, w557, w558, w559, w560, w561, w562, w563, w564, w565, w566, w567, w568, w569, w570, w571, w572, w573, w574, w575, w576, w577, w578, w579, w580, w581, w582, w583, w584, w585, w586, w587, w588, w589, w590, w591, w592, w593, w594, w595, w596, w597, w598, w599, w600, w601, w602, w603, w604, w605, w606, w607, w608, w609, w610, w611, w612, w613, w614, w615, w616, w617, w618, w619, w620, w621, w622, w623, w624, w625, w626, w627, w628, w629, w630, w631, w632, w633, w634, w635, w636, w637, w638, w639, w640, w641, w642, w643, w644, w645, w646, w647, w648, w649, w650, w651, w652, w653, w654, w655, w656, w657, w658, w659, w660, w661, w662, w663, w664, w665, w666, w667, w668, w669, w670, w671, w672, w673, w674, w675, w676, w677, w678, w679, w680, w681, w682, w683, w684, w685, w686, w687, w688, w689, w690, w691, w692, w693, w694, w695, w696, w697, w698, w699, w700, w701, w702, w703, w704, w705, w706, w707, w708, w709, w710, w711, w712, w713, w714, w715, w716, w717, w718, w719, w720, w721, w722, w723, w724, w725, w726, w727, w728, w729, w730, w731, w732, w733, w734, w735, w736, w737, w738, w739, w740, w741, w742, w743, w744, w745, w746, w747, w748, w749, w750, w751, w752, w753, w754, w755, w756, w757, w758, w759, w760, w761, w762, w763, w764, w765, w766, w767, w768, w769, w770, w771, w772, w773, w774, w775, w776, w777, w778, w779, w780, w781, w782, w783, w784, w785, w786, w787, w788, w789, w790, w791, w792, w793, w794, w795, w796, w797, w798, w799, w800, w801, w802, w803, w804, w805, w806, w807, w808, w809, w810, w811, w812, w813, w814, w815, w816, w817, w818, w819, w820, w821, w822, w823, w824, w825, w826, w827, w828, w829, w830, w831, w832, w833, w834, w835, w836, w837, w838, w839, w840, w841, w842, w843, w844, w845, w846, w847, w848, w849, w850, w851, w852, w853, w854, w855, w856, w857, w858, w859, w860, w861, w862, w863, w864, w865, w866, w867, w868, w869, w870, w871, w872, w873, w874, w875, w876, w877, w878, w879, w880, w881, w882, w883, w884, w885, w886, w887, w888, w889, w890, w891, w892, w893, w894, w895, w896, w897, w898, w899, w900, w901, w902, w903, w904, w905, w906, w907, w908, w909, w910, w911, w912, w913, w914, w915, w916, w917, w918, w919, w920, w921, w922, w923, w924, w925, w926, w927, w928, w929, w930, w931, w932, w933, w934, w935, w936, w937, w938, w939, w940, w941, w942, w943, w944, w945, w946, w947, w948, w949, w950, w951, w952, w953, w954, w955, w956, w957, w958, w959, w960, w961, w962, w963, w964, w965, w966, w967, w968, w969, w970, w971, w972, w973, w974, w975, w976, w977, w978, w979, w980, w981, w982, w983, w984, w985, w986, w987, w988, w989, w990, w991, w992, w993, w994, w995, w996, w997, w998, w999, w1000, w1001, w1002, w1003, w1004, w1005, w1006, w1007, w1008, w1009, w1010, w1011, w1012, w1013, w1014, w1015, w1016, w1017, w1018, w1019, w1020, w1021, w1022, w1023, w1024, w1025, w1026, w1027, w1028, w1029, w1030, w1031, w1032, w1033, w1034, w1035, w1036, w1037, w1038, w1039, w1040, w1041, w1042, w1043, w1044, w1045, w1046, w1047, w1048, w1049, w1050, w1051, w1052, w1053, w1054, w1055, w1056, w1057, w1058, w1059, w1060, w1061, w1062, w1063, w1064, w1065, w1066, w1067, w1068, w1069, w1070, w1071, w1072, w1073, w1074, w1075, w1076, w1077, w1078, w1079, w1080, w1081, w1082, w1083, w1084, w1085, w1086, w1087, w1088, w1089, w1090, w1091, w1092, w1093, w1094, w1095, w1096, w1097, w1098, w1099, w1100, w1101, w1102, w1103, w1104, w1105, w1106, w1107, w1108, w1109, w1110, w1111, w1112, w1113, w1114, w1115, w1116, w1117, w1118, w1119, w1120, w1121, w1122, w1123, w1124, w1125, w1126, w1127, w1128, w1129, w1130, w1131, w1132, w1133, w1134, w1135, w1136, w1137, w1138, w1139, w1140, w1141, w1142, w1143, w1144, w1145, w1146, w1147, w1148, w1149, w1150, w1151, w1152, w1153, w1154, w1155, w1156, w1157, w1158, w1159, w1160, w1161, w1162, w1163, w1164, w1165, w1166, w1167, w1168, w1169, w1170, w1171, w1172, w1173, w1174, w1175, w1176, w1177, w1178, w1179, w1180, w1181, w1182, w1183, w1184, w1185, w1186, w1187, w1188, w1189, w1190, w1191, w1192, w1193, w1194, w1195, w1196, w1197, w1198, w1199, w1200, w1201, w1202, w1203, w1204, w1205, w1206, w1207, w1208, w1209, w1210, w1211, w1212, w1213, w1214, w1215, w1216, w1217, w1218, w1219, w1220, w1221, w1222, w1223, w1224, w1225, w1226, w1227, w1228, w1229, w1230, w1231, w1232, w1233, w1234, w1235, w1236, w1237, w1238, w1239, w1240, w1241, w1242, w1243, w1244, w1245, w1246, w1247, w1248, w1249, w1250, w1251, w1252, w1253, w1254, w1255, w1256, w1257, w1258, w1259, w1260, w1261, w1262, w1263, w1264, w1265, w1266, w1267, w1268, w1269, w1270, w1271, w1272, w1273, w1274, w1275, w1276, w1277, w1278, w1279, w1280, w1281, w1282, w1283, w1284, w1285, w1286, w1287, w1288, w1289, w1290, w1291, w1292, w1293, w1294, w1295, w1296, w1297, w1298, w1299, w1300, w1301, w1302, w1303, w1304, w1305, w1306, w1307, w1308, w1309, w1310, w1311, w1312, w1313, w1314, w1315, w1316, w1317, w1318, w1319, w1320, w1321, w1322, w1323, w1324, w1325, w1326, w1327, w1328, w1329, w1330, w1331, w1332, w1333, w1334, w1335, w1336, w1337, w1338, w1339, w1340, w1341, w1342, w1343, w1344, w1345, w1346, w1347, w1348, w1349, w1350, w1351, w1352, w1353, w1354, w1355, w1356, w1357, w1358, w1359, w1360, w1361, w1362, w1363, w1364, w1365, w1366, w1367, w1368, w1369, w1370, w1371, w1372, w1373, w1374, w1375, w1376, w1377, w1378, w1379, w1380, w1381, w1382, w1383, w1384, w1385, w1386, w1387, w1388, w1389, w1390, w1391, w1392, w1393, w1394, w1395, w1396, w1397, w1398, w1399, w1400, w1401, w1402, w1403, w1404, w1405, w1406, w1407, w1408, w1409, w1410, w1411, w1412, w1413, w1414, w1415, w1416, w1417, w1418, w1419, w1420, w1421, w1422, w1423, w1424, w1425, w1426, w1427, w1428, w1429, w1430, w1431, w1432, w1433, w1434, w1435, w1436, w1437, w1438, w1439, w1440, w1441, w1442, w1443, w1444, w1445, w1446, w1447, w1448, w1449, w1450, w1451, w1452, w1453, w1454, w1455, w1456, w1457, w1458, w1459, w1460, w1461, w1462, w1463, w1464, w1465, w1466, w1467, w1468, w1469, w1470, w1471, w1472, w1473, w1474, w1475, w1476, w1477, w1478, w1479, w1480, w1481, w1482, w1483, w1484, w1485, w1486, w1487, w1488, w1489, w1490, w1491, w1492, w1493, w1494, w1495, w1496, w1497, w1498, w1499, w1500, w1501, w1502, w1503, w1504, w1505, w1506, w1507, w1508, w1509, w1510, w1511, w1512, w1513, w1514, w1515, w1516, w1517, w1518, w1519, w1520, w1521, w1522, w1523, w1524, w1525, w1526, w1527, w1528, w1529, w1530, w1531, w1532, w1533, w1534, w1535, w1536, w1537, w1538, w1539, w1540, w1541, w1542, w1543, w1544, w1545, w1546, w1547, w1548, w1549, w1550, w1551, w1552, w1553, w1554, w1555, w1556, w1557, w1558, w1559, w1560, w1561, w1562, w1563, w1564, w1565, w1566, w1567, w1568, w1569, w1570, w1571, w1572, w1573, w1574, w1575, w1576, w1577, w1578, w1579, w1580, w1581, w1582, w1583, w1584, w1585, w1586, w1587, w1588, w1589, w1590, w1591, w1592, w1593, w1594, w1595, w1596, w1597, w1598, w1599, w1600, w1601, w1602, w1603, w1604, w1605, w1606, w1607, w1608, w1609, w1610, w1611, w1612, w1613, w1614, w1615, w1616, w1617, w1618, w1619, w1620, w1621, w1622, w1623, w1624, w1625, w1626, w1627, w1628, w1629, w1630, w1631, w1632, w1633, w1634, w1635, w1636, w1637, w1638, w1639, w1640, w1641, w1642, w1643, w1644, w1645, w1646, w1647, w1648, w1649, w1650, w1651, w1652, w1653, w1654, w1655, w1656, w1657, w1658, w1659, w1660, w1661, w1662, w1663, w1664, w1665, w1666, w1667, w1668, w1669, w1670, w1671, w1672, w1673, w1674, w1675, w1676, w1677, w1678, w1679, w1680, w1681, w1682, w1683, w1684, w1685, w1686, w1687, w1688, w1689, w1690, w1691, w1692, w1693, w1694, w1695, w1696, w1697, w1698, w1699, w1700, w1701, w1702, w1703, w1704, w1705, w1706, w1707, w1708, w1709, w1710, w1711, w1712, w1713, w1714, w1715, w1716, w1717, w1718, w1719, w1720, w1721, w1722, w1723, w1724, w1725, w1726, w1727, w1728, w1729, w1730, w1731, w1732, w1733, w1734, w1735, w1736, w1737, w1738, w1739, w1740, w1741, w1742, w1743, w1744, w1745, w1746, w1747, w1748, w1749, w1750, w1751, w1752, w1753, w1754, w1755, w1756, w1757, w1758, w1759, w1760, w1761, w1762, w1763, w1764, w1765, w1766, w1767, w1768, w1769, w1770, w1771, w1772, w1773, w1774, w1775, w1776, w1777, w1778, w1779, w1780, w1781, w1782, w1783, w1784, w1785, w1786, w1787, w1788, w1789, w1790, w1791, w1792, w1793, w1794, w1795, w1796, w1797, w1798, w1799, w1800, w1801, w1802, w1803, w1804, w1805, w1806, w1807, w1808, w1809, w1810, w1811, w1812, w1813, w1814, w1815, w1816, w1817, w1818, w1819, w1820, w1821, w1822, w1823, w1824, w1825, w1826, w1827, w1828, w1829, w1830, w1831, w1832, w1833, w1834, w1835, w1836, w1837, w1838, w1839, w1840, w1841, w1842, w1843, w1844, w1845, w1846, w1847, w1848, w1849, w1850, w1851, w1852, w1853, w1854, w1855, w1856, w1857, w1858, w1859, w1860, w1861, w1862, w1863, w1864, w1865, w1866, w1867, w1868, w1869, w1870, w1871, w1872, w1873, w1874, w1875, w1876, w1877, w1878, w1879, w1880, w1881, w1882, w1883, w1884, w1885, w1886, w1887, w1888, w1889, w1890, w1891, w1892, w1893, w1894, w1895, w1896, w1897, w1898, w1899, w1900, w1901, w1902, w1903, w1904, w1905, w1906, w1907, w1908, w1909, w1910, w1911, w1912, w1913, w1914, w1915, w1916, w1917, w1918, w1919, w1920, w1921, w1922, w1923, w1924, w1925, w1926, w1927, w1928, w1929, w1930, w1931, w1932, w1933, w1934, w1935, w1936, w1937, w1938, w1939, w1940, w1941, w1942, w1943, w1944, w1945, w1946, w1947, w1948, w1949, w1950, w1951, w1952, w1953, w1954, w1955, w1956, w1957, w1958, w1959, w1960, w1961, w1962, w1963, w1964, w1965, w1966, w1967, w1968, w1969, w1970, w1971, w1972, w1973, w1974, w1975, w1976, w1977, w1978, w1979, w1980, w1981, w1982, w1983, w1984, w1985, w1986, w1987, w1988, w1989, w1990, w1991, w1992, w1993, w1994, w1995, w1996, w1997, w1998, w1999, w2000, w2001, w2002, w2003, w2004, w2005, w2006, w2007, w2008, w2009, w2010, w2011, w2012, w2013, w2014, w2015, w2016, w2017, w2018, w2019, w2020, w2021, w2022, w2023, w2024, w2025, w2026, w2027, w2028, w2029, w2030, w2031, w2032, w2033, w2034, w2035, w2036, w2037, w2038, w2039, w2040, w2041, w2042, w2043, w2044, w2045, w2046, w2047, w2048, w2049, w2050, w2051, w2052, w2053, w2054, w2055, w2056, w2057, w2058, w2059, w2060, w2061, w2062, w2063, w2064, w2065, w2066, w2067, w2068, w2069, w2070;
assign w0 = pi093 & ~pi193;
assign w1 = ~pi093 & pi193;
assign v0 = ~(w0 | w1);
assign w2 = v0;
assign w3 = pi087 & ~pi187;
assign w4 = ~pi087 & pi187;
assign v1 = ~(w3 | w4);
assign w5 = v1;
assign w6 = pi088 & ~pi188;
assign w7 = ~pi088 & pi188;
assign v2 = ~(w6 | w7);
assign w8 = v2;
assign w9 = w5 & w8;
assign v3 = ~(w5 | w8);
assign w10 = v3;
assign v4 = ~(w9 | w10);
assign w11 = v4;
assign w12 = pi086 & ~pi186;
assign w13 = ~pi086 & pi186;
assign v5 = ~(w12 | w13);
assign w14 = v5;
assign w15 = pi085 & ~pi185;
assign w16 = ~pi085 & pi185;
assign v6 = ~(w15 | w16);
assign w17 = v6;
assign v7 = ~(w14 | w17);
assign w18 = v7;
assign w19 = w14 & w17;
assign v8 = ~(w18 | w19);
assign w20 = v8;
assign w21 = pi082 & ~pi182;
assign w22 = ~pi082 & pi182;
assign v9 = ~(w21 | w22);
assign w23 = v9;
assign w24 = pi081 & ~pi181;
assign w25 = ~pi081 & pi181;
assign v10 = ~(w24 | w25);
assign w26 = v10;
assign w27 = w23 & w26;
assign v11 = ~(w23 | w26);
assign w28 = v11;
assign v12 = ~(w27 | w28);
assign w29 = v12;
assign w30 = pi074 & ~pi174;
assign w31 = ~pi074 & pi174;
assign v13 = ~(w30 | w31);
assign w32 = v13;
assign w33 = pi073 & ~pi173;
assign w34 = ~pi073 & pi173;
assign v14 = ~(w33 | w34);
assign w35 = v14;
assign w36 = w32 & w35;
assign v15 = ~(w32 | w35);
assign w37 = v15;
assign v16 = ~(w36 | w37);
assign w38 = v16;
assign w39 = pi067 & ~pi167;
assign w40 = ~pi067 & pi167;
assign v17 = ~(w39 | w40);
assign w41 = v17;
assign w42 = pi068 & ~pi168;
assign w43 = ~pi068 & pi168;
assign v18 = ~(w42 | w43);
assign w44 = v18;
assign v19 = ~(w41 | w44);
assign w45 = v19;
assign w46 = w41 & w44;
assign v20 = ~(w45 | w46);
assign w47 = v20;
assign w48 = pi069 & ~pi169;
assign w49 = ~pi069 & pi169;
assign v21 = ~(w48 | w49);
assign w50 = v21;
assign w51 = w47 & ~w50;
assign w52 = ~w47 & w50;
assign v22 = ~(w51 | w52);
assign w53 = v22;
assign w54 = pi052 & ~pi152;
assign w55 = ~pi052 & pi152;
assign v23 = ~(w54 | w55);
assign w56 = v23;
assign w57 = pi047 & ~pi147;
assign w58 = ~pi047 & pi147;
assign v24 = ~(w57 | w58);
assign w59 = v24;
assign w60 = pi048 & ~pi148;
assign w61 = ~pi048 & pi148;
assign v25 = ~(w60 | w61);
assign w62 = v25;
assign w63 = w59 & w62;
assign v26 = ~(w59 | w62);
assign w64 = v26;
assign v27 = ~(w63 | w64);
assign w65 = v27;
assign w66 = pi049 & ~pi149;
assign w67 = ~pi049 & pi149;
assign v28 = ~(w66 | w67);
assign w68 = v28;
assign w69 = pi050 & ~pi150;
assign w70 = ~pi050 & pi150;
assign v29 = ~(w69 | w70);
assign w71 = v29;
assign v30 = ~(w68 | w71);
assign w72 = v30;
assign w73 = w68 & w71;
assign v31 = ~(w72 | w73);
assign w74 = v31;
assign w75 = w65 & ~w74;
assign w76 = ~w65 & w74;
assign v32 = ~(w75 | w76);
assign w77 = v32;
assign w78 = pi051 & ~pi151;
assign w79 = ~pi051 & pi151;
assign v33 = ~(w78 | w79);
assign w80 = v33;
assign w81 = pi043 & ~pi143;
assign w82 = ~pi043 & pi143;
assign v34 = ~(w81 | w82);
assign w83 = v34;
assign w84 = pi044 & ~pi144;
assign w85 = ~pi044 & pi144;
assign v35 = ~(w84 | w85);
assign w86 = v35;
assign w87 = w83 & w86;
assign v36 = ~(w83 | w86);
assign w88 = v36;
assign v37 = ~(w87 | w88);
assign w89 = v37;
assign w90 = pi042 & ~pi142;
assign w91 = ~pi042 & pi142;
assign v38 = ~(w90 | w91);
assign w92 = v38;
assign w93 = w89 & ~w92;
assign w94 = ~w89 & w92;
assign v39 = ~(w93 | w94);
assign w95 = v39;
assign w96 = pi046 & ~pi146;
assign w97 = ~pi046 & pi146;
assign v40 = ~(w96 | w97);
assign w98 = v40;
assign w99 = pi045 & ~pi145;
assign w100 = ~pi045 & pi145;
assign v41 = ~(w99 | w100);
assign w101 = v41;
assign w102 = w98 & ~w101;
assign w103 = ~w98 & w101;
assign v42 = ~(w102 | w103);
assign w104 = v42;
assign w105 = w95 & w104;
assign v43 = ~(w95 | w104);
assign w106 = v43;
assign v44 = ~(w105 | w106);
assign w107 = v44;
assign w108 = w80 & ~w107;
assign w109 = ~w80 & w107;
assign v45 = ~(w108 | w109);
assign w110 = v45;
assign w111 = w77 & w110;
assign v46 = ~(w77 | w110);
assign w112 = v46;
assign v47 = ~(w111 | w112);
assign w113 = v47;
assign v48 = ~(w56 | w113);
assign w114 = v48;
assign w115 = w56 & w113;
assign v49 = ~(w114 | w115);
assign w116 = v49;
assign w117 = pi010 & ~pi110;
assign w118 = ~pi010 & pi110;
assign v50 = ~(w117 | w118);
assign w119 = v50;
assign w120 = pi009 & ~pi109;
assign w121 = ~pi009 & pi109;
assign v51 = ~(w120 | w121);
assign w122 = v51;
assign v52 = ~(w119 | w122);
assign w123 = v52;
assign w124 = w119 & w122;
assign v53 = ~(w123 | w124);
assign w125 = v53;
assign w126 = pi007 & ~pi107;
assign w127 = ~pi007 & pi107;
assign v54 = ~(w126 | w127);
assign w128 = v54;
assign w129 = pi008 & ~pi108;
assign w130 = ~pi008 & pi108;
assign v55 = ~(w129 | w130);
assign w131 = v55;
assign w132 = w128 & w131;
assign v56 = ~(w128 | w131);
assign w133 = v56;
assign v57 = ~(w132 | w133);
assign w134 = v57;
assign w135 = w125 & ~w134;
assign w136 = ~w125 & w134;
assign v58 = ~(w135 | w136);
assign w137 = v58;
assign w138 = pi002 & ~pi102;
assign w139 = ~pi002 & pi102;
assign v59 = ~(w138 | w139);
assign w140 = v59;
assign w141 = pi003 & ~pi103;
assign w142 = ~pi003 & pi103;
assign v60 = ~(w141 | w142);
assign w143 = v60;
assign w144 = w140 & w143;
assign v61 = ~(w140 | w143);
assign w145 = v61;
assign v62 = ~(w144 | w145);
assign w146 = v62;
assign w147 = pi000 & ~pi100;
assign w148 = ~pi000 & pi100;
assign v63 = ~(w147 | w148);
assign w149 = v63;
assign w150 = pi001 & ~pi101;
assign w151 = ~pi001 & pi101;
assign v64 = ~(w150 | w151);
assign w152 = v64;
assign w153 = w149 & w152;
assign v65 = ~(w149 | w152);
assign w154 = v65;
assign v66 = ~(w153 | w154);
assign w155 = v66;
assign w156 = w146 & w155;
assign v67 = ~(w146 | w155);
assign w157 = v67;
assign v68 = ~(w156 | w157);
assign w158 = v68;
assign w159 = pi005 & ~pi105;
assign w160 = ~pi005 & pi105;
assign v69 = ~(w159 | w160);
assign w161 = v69;
assign w162 = pi006 & ~pi106;
assign w163 = ~pi006 & pi106;
assign v70 = ~(w162 | w163);
assign w164 = v70;
assign w165 = w161 & w164;
assign v71 = ~(w161 | w164);
assign w166 = v71;
assign v72 = ~(w165 | w166);
assign w167 = v72;
assign w168 = pi004 & ~pi104;
assign w169 = ~pi004 & pi104;
assign v73 = ~(w168 | w169);
assign w170 = v73;
assign w171 = w167 & ~w170;
assign w172 = ~w167 & w170;
assign v74 = ~(w171 | w172);
assign w173 = v74;
assign w174 = w158 & w173;
assign v75 = ~(w158 | w173);
assign w175 = v75;
assign v76 = ~(w174 | w175);
assign w176 = v76;
assign w177 = ~w137 & w176;
assign w178 = w137 & ~w176;
assign v77 = ~(w177 | w178);
assign w179 = v77;
assign w180 = pi014 & ~pi114;
assign w181 = ~pi014 & pi114;
assign v78 = ~(w180 | w181);
assign w182 = v78;
assign w183 = pi013 & ~pi113;
assign w184 = ~pi013 & pi113;
assign v79 = ~(w183 | w184);
assign w185 = v79;
assign v80 = ~(w182 | w185);
assign w186 = v80;
assign w187 = w182 & w185;
assign v81 = ~(w186 | w187);
assign w188 = v81;
assign w189 = pi011 & ~pi111;
assign w190 = ~pi011 & pi111;
assign v82 = ~(w189 | w190);
assign w191 = v82;
assign w192 = pi012 & ~pi112;
assign w193 = ~pi012 & pi112;
assign v83 = ~(w192 | w193);
assign w194 = v83;
assign w195 = w191 & w194;
assign v84 = ~(w191 | w194);
assign w196 = v84;
assign v85 = ~(w195 | w196);
assign w197 = v85;
assign w198 = ~w188 & w197;
assign w199 = w188 & ~w197;
assign v86 = ~(w198 | w199);
assign w200 = v86;
assign w201 = pi015 & ~pi115;
assign w202 = ~pi015 & pi115;
assign v87 = ~(w201 | w202);
assign w203 = v87;
assign w204 = w200 & w203;
assign v88 = ~(w200 | w203);
assign w205 = v88;
assign v89 = ~(w204 | w205);
assign w206 = v89;
assign w207 = pi035 & ~pi135;
assign w208 = ~pi035 & pi135;
assign v90 = ~(w207 | w208);
assign w209 = v90;
assign w210 = pi036 & ~pi136;
assign w211 = ~pi036 & pi136;
assign v91 = ~(w210 | w211);
assign w212 = v91;
assign v92 = ~(w209 | w212);
assign w213 = v92;
assign w214 = w209 & w212;
assign v93 = ~(w213 | w214);
assign w215 = v93;
assign w216 = pi034 & ~pi134;
assign w217 = ~pi034 & pi134;
assign v94 = ~(w216 | w217);
assign w218 = v94;
assign w219 = pi016 & ~pi116;
assign w220 = ~pi016 & pi116;
assign v95 = ~(w219 | w220);
assign w221 = v95;
assign w222 = w218 & w221;
assign v96 = ~(w218 | w221);
assign w223 = v96;
assign v97 = ~(w222 | w223);
assign w224 = v97;
assign w225 = w215 & w224;
assign v98 = ~(w215 | w224);
assign w226 = v98;
assign v99 = ~(w225 | w226);
assign w227 = v99;
assign w228 = pi031 & ~pi131;
assign w229 = ~pi031 & pi131;
assign v100 = ~(w228 | w229);
assign w230 = v100;
assign w231 = pi032 & ~pi132;
assign w232 = ~pi032 & pi132;
assign v101 = ~(w231 | w232);
assign w233 = v101;
assign w234 = w230 & w233;
assign v102 = ~(w230 | w233);
assign w235 = v102;
assign v103 = ~(w234 | w235);
assign w236 = v103;
assign w237 = pi033 & ~pi133;
assign w238 = ~pi033 & pi133;
assign v104 = ~(w237 | w238);
assign w239 = v104;
assign w240 = ~w236 & w239;
assign w241 = w236 & ~w239;
assign v105 = ~(w240 | w241);
assign w242 = v105;
assign w243 = w227 & ~w242;
assign w244 = ~w227 & w242;
assign v106 = ~(w243 | w244);
assign w245 = v106;
assign w246 = w206 & ~w245;
assign w247 = ~w206 & w245;
assign v107 = ~(w246 | w247);
assign w248 = v107;
assign w249 = w179 & w248;
assign v108 = ~(w179 | w248);
assign w250 = v108;
assign v109 = ~(w249 | w250);
assign w251 = v109;
assign w252 = pi023 & ~pi123;
assign w253 = ~pi023 & pi123;
assign v110 = ~(w252 | w253);
assign w254 = v110;
assign w255 = pi024 & ~pi124;
assign w256 = ~pi024 & pi124;
assign v111 = ~(w255 | w256);
assign w257 = v111;
assign w258 = w254 & w257;
assign v112 = ~(w254 | w257);
assign w259 = v112;
assign v113 = ~(w258 | w259);
assign w260 = v113;
assign w261 = pi022 & ~pi122;
assign w262 = ~pi022 & pi122;
assign v114 = ~(w261 | w262);
assign w263 = v114;
assign w264 = w260 & ~w263;
assign w265 = ~w260 & w263;
assign v115 = ~(w264 | w265);
assign w266 = v115;
assign w267 = pi025 & ~pi125;
assign w268 = ~pi025 & pi125;
assign v116 = ~(w267 | w268);
assign w269 = v116;
assign w270 = pi026 & ~pi126;
assign w271 = ~pi026 & pi126;
assign v117 = ~(w270 | w271);
assign w272 = v117;
assign v118 = ~(w269 | w272);
assign w273 = v118;
assign w274 = w269 & w272;
assign v119 = ~(w273 | w274);
assign w275 = v119;
assign w276 = pi027 & ~pi127;
assign w277 = ~pi027 & pi127;
assign v120 = ~(w276 | w277);
assign w278 = v120;
assign w279 = w275 & ~w278;
assign w280 = ~w275 & w278;
assign v121 = ~(w279 | w280);
assign w281 = v121;
assign w282 = w266 & w281;
assign v122 = ~(w266 | w281);
assign w283 = v122;
assign v123 = ~(w282 | w283);
assign w284 = v123;
assign w285 = pi021 & ~pi121;
assign w286 = ~pi021 & pi121;
assign v124 = ~(w285 | w286);
assign w287 = v124;
assign w288 = pi019 & ~pi119;
assign w289 = ~pi019 & pi119;
assign v125 = ~(w288 | w289);
assign w290 = v125;
assign w291 = pi020 & ~pi120;
assign w292 = ~pi020 & pi120;
assign v126 = ~(w291 | w292);
assign w293 = v126;
assign v127 = ~(w290 | w293);
assign w294 = v127;
assign w295 = w290 & w293;
assign v128 = ~(w294 | w295);
assign w296 = v128;
assign w297 = pi017 & ~pi117;
assign w298 = ~pi017 & pi117;
assign v129 = ~(w297 | w298);
assign w299 = v129;
assign w300 = pi018 & ~pi118;
assign w301 = ~pi018 & pi118;
assign v130 = ~(w300 | w301);
assign w302 = v130;
assign w303 = w299 & w302;
assign v131 = ~(w299 | w302);
assign w304 = v131;
assign v132 = ~(w303 | w304);
assign w305 = v132;
assign w306 = w296 & w305;
assign v133 = ~(w296 | w305);
assign w307 = v133;
assign v134 = ~(w306 | w307);
assign w308 = v134;
assign w309 = w287 & w308;
assign v135 = ~(w287 | w308);
assign w310 = v135;
assign v136 = ~(w309 | w310);
assign w311 = v136;
assign w312 = w284 & w311;
assign v137 = ~(w284 | w311);
assign w313 = v137;
assign v138 = ~(w312 | w313);
assign w314 = v138;
assign w315 = pi039 & ~pi139;
assign w316 = ~pi039 & pi139;
assign v139 = ~(w315 | w316);
assign w317 = v139;
assign w318 = pi040 & ~pi140;
assign w319 = ~pi040 & pi140;
assign v140 = ~(w318 | w319);
assign w320 = v140;
assign v141 = ~(w317 | w320);
assign w321 = v141;
assign w322 = w317 & w320;
assign v142 = ~(w321 | w322);
assign w323 = v142;
assign w324 = pi037 & ~pi137;
assign w325 = ~pi037 & pi137;
assign v143 = ~(w324 | w325);
assign w326 = v143;
assign w327 = pi038 & ~pi138;
assign w328 = ~pi038 & pi138;
assign v144 = ~(w327 | w328);
assign w329 = v144;
assign w330 = w326 & w329;
assign v145 = ~(w326 | w329);
assign w331 = v145;
assign v146 = ~(w330 | w331);
assign w332 = v146;
assign w333 = w323 & ~w332;
assign w334 = ~w323 & w332;
assign v147 = ~(w333 | w334);
assign w335 = v147;
assign w336 = pi041 & ~pi141;
assign w337 = ~pi041 & pi141;
assign v148 = ~(w336 | w337);
assign w338 = v148;
assign w339 = pi028 & ~pi128;
assign w340 = ~pi028 & pi128;
assign v149 = ~(w339 | w340);
assign w341 = v149;
assign w342 = pi029 & ~pi129;
assign w343 = ~pi029 & pi129;
assign v150 = ~(w342 | w343);
assign w344 = v150;
assign w345 = pi030 & ~pi130;
assign w346 = ~pi030 & pi130;
assign v151 = ~(w345 | w346);
assign w347 = v151;
assign w348 = w344 & ~w347;
assign w349 = ~w344 & w347;
assign v152 = ~(w348 | w349);
assign w350 = v152;
assign w351 = w341 & w350;
assign v153 = ~(w341 | w350);
assign w352 = v153;
assign v154 = ~(w351 | w352);
assign w353 = v154;
assign w354 = w338 & ~w353;
assign w355 = ~w338 & w353;
assign v155 = ~(w354 | w355);
assign w356 = v155;
assign w357 = w335 & ~w356;
assign w358 = ~w335 & w356;
assign v156 = ~(w357 | w358);
assign w359 = v156;
assign w360 = w314 & ~w359;
assign w361 = ~w314 & w359;
assign v157 = ~(w360 | w361);
assign w362 = v157;
assign w363 = w251 & w362;
assign v158 = ~(w251 | w362);
assign w364 = v158;
assign v159 = ~(w363 | w364);
assign w365 = v159;
assign w366 = w116 & w365;
assign v160 = ~(w116 | w365);
assign w367 = v160;
assign v161 = ~(w366 | w367);
assign w368 = v161;
assign w369 = pi058 & ~pi158;
assign w370 = ~pi058 & pi158;
assign v162 = ~(w369 | w370);
assign w371 = v162;
assign w372 = pi059 & ~pi159;
assign w373 = ~pi059 & pi159;
assign v163 = ~(w372 | w373);
assign w374 = v163;
assign w375 = pi060 & ~pi160;
assign w376 = ~pi060 & pi160;
assign v164 = ~(w375 | w376);
assign w377 = v164;
assign v165 = ~(w374 | w377);
assign w378 = v165;
assign w379 = w374 & w377;
assign v166 = ~(w378 | w379);
assign w380 = v166;
assign w381 = pi061 & ~pi161;
assign w382 = ~pi061 & pi161;
assign v167 = ~(w381 | w382);
assign w383 = v167;
assign w384 = pi053 & ~pi153;
assign w385 = ~pi053 & pi153;
assign v168 = ~(w384 | w385);
assign w386 = v168;
assign w387 = pi054 & ~pi154;
assign w388 = ~pi054 & pi154;
assign v169 = ~(w387 | w388);
assign w389 = v169;
assign w390 = w386 & w389;
assign v170 = ~(w386 | w389);
assign w391 = v170;
assign v171 = ~(w390 | w391);
assign w392 = v171;
assign w393 = pi055 & ~pi155;
assign w394 = ~pi055 & pi155;
assign v172 = ~(w393 | w394);
assign w395 = v172;
assign w396 = pi056 & ~pi156;
assign w397 = ~pi056 & pi156;
assign v173 = ~(w396 | w397);
assign w398 = v173;
assign v174 = ~(w395 | w398);
assign w399 = v174;
assign w400 = w395 & w398;
assign v175 = ~(w399 | w400);
assign w401 = v175;
assign w402 = pi057 & ~pi157;
assign w403 = ~pi057 & pi157;
assign v176 = ~(w402 | w403);
assign w404 = v176;
assign w405 = w401 & ~w404;
assign w406 = ~w401 & w404;
assign v177 = ~(w405 | w406);
assign w407 = v177;
assign w408 = w392 & w407;
assign v178 = ~(w392 | w407);
assign w409 = v178;
assign v179 = ~(w408 | w409);
assign w410 = v179;
assign v180 = ~(w383 | w410);
assign w411 = v180;
assign w412 = w383 & w410;
assign v181 = ~(w411 | w412);
assign w413 = v181;
assign w414 = w380 & ~w413;
assign w415 = ~w380 & w413;
assign v182 = ~(w414 | w415);
assign w416 = v182;
assign w417 = w371 & ~w416;
assign w418 = ~w371 & w416;
assign v183 = ~(w417 | w418);
assign w419 = v183;
assign w420 = w368 & w419;
assign v184 = ~(w368 | w419);
assign w421 = v184;
assign v185 = ~(w420 | w421);
assign w422 = v185;
assign w423 = pi064 & ~pi164;
assign w424 = ~pi064 & pi164;
assign v186 = ~(w423 | w424);
assign w425 = v186;
assign w426 = pi065 & ~pi165;
assign w427 = ~pi065 & pi165;
assign v187 = ~(w426 | w427);
assign w428 = v187;
assign w429 = pi066 & ~pi166;
assign w430 = ~pi066 & pi166;
assign v188 = ~(w429 | w430);
assign w431 = v188;
assign v189 = ~(w428 | w431);
assign w432 = v189;
assign w433 = w428 & w431;
assign v190 = ~(w432 | w433);
assign w434 = v190;
assign w435 = pi063 & ~pi163;
assign w436 = ~pi063 & pi163;
assign v191 = ~(w435 | w436);
assign w437 = v191;
assign w438 = pi062 & ~pi162;
assign w439 = ~pi062 & pi162;
assign v192 = ~(w438 | w439);
assign w440 = v192;
assign v193 = ~(w437 | w440);
assign w441 = v193;
assign w442 = w437 & w440;
assign v194 = ~(w441 | w442);
assign w443 = v194;
assign w444 = w434 & ~w443;
assign w445 = ~w434 & w443;
assign v195 = ~(w444 | w445);
assign w446 = v195;
assign w447 = w425 & ~w446;
assign w448 = ~w425 & w446;
assign v196 = ~(w447 | w448);
assign w449 = v196;
assign w450 = w422 & w449;
assign v197 = ~(w422 | w449);
assign w451 = v197;
assign v198 = ~(w450 | w451);
assign w452 = v198;
assign w453 = w53 & w452;
assign v199 = ~(w53 | w452);
assign w454 = v199;
assign v200 = ~(w453 | w454);
assign w455 = v200;
assign w456 = pi070 & ~pi170;
assign w457 = ~pi070 & pi170;
assign v201 = ~(w456 | w457);
assign w458 = v201;
assign w459 = pi071 & ~pi171;
assign w460 = ~pi071 & pi171;
assign v202 = ~(w459 | w460);
assign w461 = v202;
assign w462 = pi072 & ~pi172;
assign w463 = ~pi072 & pi172;
assign v203 = ~(w462 | w463);
assign w464 = v203;
assign w465 = w461 & ~w464;
assign w466 = ~w461 & w464;
assign v204 = ~(w465 | w466);
assign w467 = v204;
assign w468 = w458 & ~w467;
assign w469 = ~w458 & w467;
assign v205 = ~(w468 | w469);
assign w470 = v205;
assign w471 = w455 & w470;
assign v206 = ~(w455 | w470);
assign w472 = v206;
assign v207 = ~(w471 | w472);
assign w473 = v207;
assign w474 = w38 & ~w473;
assign w475 = ~w38 & w473;
assign v208 = ~(w474 | w475);
assign w476 = v208;
assign w477 = pi075 & ~pi175;
assign w478 = ~pi075 & pi175;
assign v209 = ~(w477 | w478);
assign w479 = v209;
assign w480 = pi076 & ~pi176;
assign w481 = ~pi076 & pi176;
assign v210 = ~(w480 | w481);
assign w482 = v210;
assign w483 = w479 & w482;
assign v211 = ~(w479 | w482);
assign w484 = v211;
assign v212 = ~(w483 | w484);
assign w485 = v212;
assign w486 = w476 & ~w485;
assign w487 = ~w476 & w485;
assign v213 = ~(w486 | w487);
assign w488 = v213;
assign w489 = pi079 & ~pi179;
assign w490 = ~pi079 & pi179;
assign v214 = ~(w489 | w490);
assign w491 = v214;
assign w492 = pi080 & ~pi180;
assign w493 = ~pi080 & pi180;
assign v215 = ~(w492 | w493);
assign w494 = v215;
assign v216 = ~(w491 | w494);
assign w495 = v216;
assign w496 = w491 & w494;
assign v217 = ~(w495 | w496);
assign w497 = v217;
assign w498 = pi077 & ~pi177;
assign w499 = ~pi077 & pi177;
assign v218 = ~(w498 | w499);
assign w500 = v218;
assign w501 = pi078 & ~pi178;
assign w502 = ~pi078 & pi178;
assign v219 = ~(w501 | w502);
assign w503 = v219;
assign w504 = w500 & w503;
assign v220 = ~(w500 | w503);
assign w505 = v220;
assign v221 = ~(w504 | w505);
assign w506 = v221;
assign w507 = w497 & ~w506;
assign w508 = ~w497 & w506;
assign v222 = ~(w507 | w508);
assign w509 = v222;
assign w510 = w488 & w509;
assign v223 = ~(w488 | w509);
assign w511 = v223;
assign v224 = ~(w510 | w511);
assign w512 = v224;
assign w513 = w29 & ~w512;
assign w514 = ~w29 & w512;
assign v225 = ~(w513 | w514);
assign w515 = v225;
assign w516 = pi083 & ~pi183;
assign w517 = ~pi083 & pi183;
assign v226 = ~(w516 | w517);
assign w518 = v226;
assign w519 = pi084 & ~pi184;
assign w520 = ~pi084 & pi184;
assign v227 = ~(w519 | w520);
assign w521 = v227;
assign w522 = w518 & w521;
assign v228 = ~(w518 | w521);
assign w523 = v228;
assign v229 = ~(w522 | w523);
assign w524 = v229;
assign w525 = w515 & w524;
assign v230 = ~(w515 | w524);
assign w526 = v230;
assign v231 = ~(w525 | w526);
assign w527 = v231;
assign w528 = w20 & ~w527;
assign w529 = ~w20 & w527;
assign v232 = ~(w528 | w529);
assign w530 = v232;
assign w531 = w11 & ~w530;
assign w532 = ~w11 & w530;
assign v233 = ~(w531 | w532);
assign w533 = v233;
assign w534 = pi089 & ~pi189;
assign w535 = ~pi089 & pi189;
assign v234 = ~(w534 | w535);
assign w536 = v234;
assign w537 = pi090 & ~pi190;
assign w538 = ~pi090 & pi190;
assign v235 = ~(w537 | w538);
assign w539 = v235;
assign w540 = w536 & w539;
assign v236 = ~(w536 | w539);
assign w541 = v236;
assign v237 = ~(w540 | w541);
assign w542 = v237;
assign w543 = w533 & w542;
assign v238 = ~(w533 | w542);
assign w544 = v238;
assign v239 = ~(w543 | w544);
assign w545 = v239;
assign w546 = pi091 & ~pi191;
assign w547 = ~pi091 & pi191;
assign v240 = ~(w546 | w547);
assign w548 = v240;
assign w549 = pi092 & ~pi192;
assign w550 = ~pi092 & pi192;
assign v241 = ~(w549 | w550);
assign w551 = v241;
assign w552 = w548 & w551;
assign v242 = ~(w548 | w551);
assign w553 = v242;
assign v243 = ~(w552 | w553);
assign w554 = v243;
assign w555 = w545 & w554;
assign v244 = ~(w545 | w554);
assign w556 = v244;
assign v245 = ~(w555 | w556);
assign w557 = v245;
assign v246 = ~(w2 | w557);
assign w558 = v246;
assign w559 = w2 & w557;
assign v247 = ~(w558 | w559);
assign w560 = v247;
assign w561 = pi094 & ~pi194;
assign w562 = ~pi094 & pi194;
assign v248 = ~(w561 | w562);
assign w563 = v248;
assign w564 = pi095 & ~pi195;
assign w565 = ~pi095 & pi195;
assign v249 = ~(w564 | w565);
assign w566 = v249;
assign w567 = w563 & w566;
assign v250 = ~(w563 | w566);
assign w568 = v250;
assign v251 = ~(w567 | w568);
assign w569 = v251;
assign w570 = w560 & ~w569;
assign w571 = ~w560 & w569;
assign v252 = ~(w570 | w571);
assign w572 = v252;
assign w573 = pi096 & ~pi196;
assign w574 = ~pi096 & pi196;
assign v253 = ~(w573 | w574);
assign w575 = v253;
assign w576 = w572 & w575;
assign v254 = ~(w572 | w575);
assign w577 = v254;
assign v255 = ~(w576 | w577);
assign w578 = v255;
assign w579 = pi097 & ~pi197;
assign w580 = ~pi097 & pi197;
assign v256 = ~(w579 | w580);
assign w581 = v256;
assign w582 = ~w578 & w581;
assign w583 = w578 & ~w581;
assign v257 = ~(w582 | w583);
assign w584 = v257;
assign w585 = pi098 & ~pi198;
assign w586 = ~pi098 & pi198;
assign v258 = ~(w585 | w586);
assign w587 = v258;
assign w588 = w584 & w587;
assign v259 = ~(w584 | w587);
assign w589 = v259;
assign v260 = ~(w588 | w589);
assign w590 = v260;
assign w591 = pi099 & ~pi199;
assign w592 = ~pi099 & pi199;
assign v261 = ~(w591 | w592);
assign w593 = v261;
assign v262 = ~(w590 | w593);
assign w594 = v262;
assign w595 = w590 & w593;
assign v263 = ~(w594 | w595);
assign w596 = v263;
assign v264 = ~(w545 | w548);
assign w597 = v264;
assign w598 = ~w551 & w557;
assign w599 = (~w597 & ~w557) | (~w597 & w1841) | (~w557 & w1841);
assign w600 = ~w521 & w527;
assign w601 = (~w27 & w512) | (~w27 & w1842) | (w512 & w1842);
assign v265 = ~(w422 | w443);
assign w602 = v265;
assign w603 = w422 & w443;
assign v266 = ~(w602 | w603);
assign w604 = v266;
assign v267 = ~(w425 | w604);
assign w605 = v267;
assign w606 = ~w604 & w1843;
assign v268 = ~(w107 | w365);
assign w607 = v268;
assign w608 = w107 & w365;
assign v269 = ~(w607 | w608);
assign w609 = v269;
assign w610 = ~w98 & w609;
assign w611 = ~w95 & w365;
assign w612 = w95 & ~w365;
assign v270 = ~(w611 | w612);
assign w613 = v270;
assign v271 = ~(w101 | w613);
assign w614 = v271;
assign v272 = ~(w610 | w614);
assign w615 = v272;
assign w616 = (~w64 & w609) | (~w64 & w1767) | (w609 & w1767);
assign w617 = w615 & ~w616;
assign w618 = ~w615 & w616;
assign v273 = ~(w617 | w618);
assign w619 = v273;
assign w620 = ~w92 & w365;
assign v274 = ~(w338 | w365);
assign w621 = v274;
assign v275 = ~(w620 | w621);
assign w622 = v275;
assign w623 = w92 & ~w365;
assign v276 = ~(w620 | w623);
assign w624 = v276;
assign w625 = (~w88 & ~w624) | (~w88 & w1768) | (~w624 & w1768);
assign w626 = ~w622 & w625;
assign w627 = w622 & ~w625;
assign v277 = ~(w626 | w627);
assign w628 = v277;
assign w629 = w619 & w628;
assign v278 = ~(w619 | w628);
assign w630 = v278;
assign v279 = ~(w629 | w630);
assign w631 = v279;
assign w632 = w609 & w1769;
assign w633 = (~w73 & w609) | (~w73 & w1770) | (w609 & w1770);
assign w634 = ~w632 & w633;
assign w635 = w314 & w353;
assign v280 = ~(w314 | w353);
assign w636 = v280;
assign v281 = ~(w635 | w636);
assign w637 = v281;
assign w638 = w251 & w637;
assign v282 = ~(w251 | w637);
assign w639 = v282;
assign v283 = ~(w638 | w639);
assign w640 = v283;
assign w641 = w332 & ~w640;
assign w642 = (~w331 & w640) | (~w331 & w1844) | (w640 & w1844);
assign w643 = (~w214 & w640) | (~w214 & w1845) | (w640 & w1845);
assign w644 = w642 & ~w643;
assign w645 = ~w642 & w643;
assign v284 = ~(w644 | w645);
assign w646 = v284;
assign w647 = w634 & w646;
assign v285 = ~(w634 | w646);
assign w648 = v285;
assign v286 = ~(w647 | w648);
assign w649 = v286;
assign w650 = w631 & w649;
assign v287 = ~(w631 | w649);
assign w651 = v287;
assign v288 = ~(w650 | w651);
assign w652 = v288;
assign w653 = ~w206 & w221;
assign w654 = w206 & ~w221;
assign v289 = ~(w653 | w654);
assign w655 = v289;
assign w656 = w179 & w655;
assign v290 = ~(w179 | w655);
assign w657 = v290;
assign v291 = ~(w656 | w657);
assign w658 = v291;
assign w659 = w311 & w658;
assign v292 = ~(w311 | w658);
assign w660 = v292;
assign v293 = ~(w659 | w660);
assign w661 = v293;
assign v294 = ~(w263 | w661);
assign w662 = v294;
assign w663 = w263 & w661;
assign v295 = ~(w662 | w663);
assign w664 = v295;
assign w665 = (~w259 & ~w664) | (~w259 & w1804) | (~w664 & w1804);
assign w666 = w266 & w661;
assign v296 = ~(w266 | w661);
assign w667 = v296;
assign v297 = ~(w666 | w667);
assign w668 = v297;
assign w669 = (~w274 & ~w668) | (~w274 & w1805) | (~w668 & w1805);
assign w670 = ~w665 & w669;
assign w671 = w665 & ~w669;
assign v298 = ~(w670 | w671);
assign w672 = v298;
assign v299 = ~(w140 | w153);
assign w673 = v299;
assign w674 = ~w673 & w1846;
assign w675 = w144 & w153;
assign w676 = w145 & w154;
assign w677 = (~w170 & w673) | (~w170 & w1847) | (w673 & w1847);
assign w678 = (~w676 & ~w158) | (~w676 & w1848) | (~w158 & w1848);
assign w679 = (~w675 & ~w158) | (~w675 & w2028) | (~w158 & w2028);
assign w680 = w678 & w679;
assign w681 = (~w166 & w176) | (~w166 & w1806) | (w176 & w1806);
assign w682 = w680 & ~w681;
assign w683 = ~w680 & w681;
assign v300 = ~(w682 | w683);
assign w684 = v300;
assign w685 = ~w176 & w1771;
assign w686 = (~w123 & ~w176) | (~w123 & w1772) | (~w176 & w1772);
assign w687 = ~w685 & w686;
assign w688 = (~w132 & w176) | (~w132 & w1807) | (w176 & w1807);
assign w689 = ~w687 & w688;
assign w690 = w687 & ~w688;
assign v301 = ~(w689 | w690);
assign w691 = v301;
assign v302 = ~(w684 | w691);
assign w692 = v302;
assign w693 = w684 & w691;
assign v303 = ~(w692 | w693);
assign w694 = v303;
assign w695 = (~w186 & ~w179) | (~w186 & w1773) | (~w179 & w1773);
assign w696 = (~w196 & ~w179) | (~w196 & w1808) | (~w179 & w1808);
assign v304 = ~(w695 | w696);
assign w697 = v304;
assign v305 = ~(w187 | w195);
assign w698 = v305;
assign w699 = (~w179 & w1809) | (~w179 & w1810) | (w1809 & w1810);
assign w700 = w696 & w699;
assign v306 = ~(w697 | w700);
assign w701 = v306;
assign w702 = w694 & ~w701;
assign w703 = ~w694 & w701;
assign v307 = ~(w702 | w703);
assign w704 = v307;
assign w705 = w179 & w206;
assign v308 = ~(w179 | w206);
assign w706 = v308;
assign v309 = ~(w705 | w706);
assign w707 = v309;
assign w708 = ~w221 & w707;
assign v310 = ~(w203 | w707);
assign w709 = v310;
assign v311 = ~(w708 | w709);
assign w710 = v311;
assign w711 = w221 & ~w304;
assign w712 = (~w303 & w707) | (~w303 & w1774) | (w707 & w1774);
assign w713 = w710 & ~w712;
assign w714 = w707 & w1775;
assign w715 = w712 & ~w714;
assign w716 = ~w710 & w715;
assign v312 = ~(w713 | w716);
assign w717 = v312;
assign w718 = w704 & ~w717;
assign w719 = ~w704 & w717;
assign v313 = ~(w718 | w719);
assign w720 = v313;
assign v314 = ~(w308 | w658);
assign w721 = v314;
assign w722 = w308 & w658;
assign v315 = ~(w721 | w722);
assign w723 = v315;
assign w724 = ~w287 & w723;
assign v316 = ~(w662 | w724);
assign w725 = v316;
assign w726 = (~w295 & ~w723) | (~w295 & w1811) | (~w723 & w1811);
assign w727 = w725 & ~w726;
assign w728 = ~w725 & w726;
assign v317 = ~(w727 | w728);
assign w729 = v317;
assign w730 = ~w720 & w729;
assign w731 = w720 & ~w729;
assign v318 = ~(w730 | w731);
assign w732 = v318;
assign w733 = ~w672 & w732;
assign w734 = w672 & ~w732;
assign v319 = ~(w733 | w734);
assign w735 = v319;
assign w736 = w637 & w658;
assign v320 = ~(w637 | w658);
assign w737 = v320;
assign v321 = ~(w736 | w737);
assign w738 = v321;
assign w739 = w236 & w239;
assign w740 = ~w738 & w739;
assign w741 = w240 & w738;
assign v322 = ~(w740 | w741);
assign w742 = v322;
assign w743 = ~w218 & w742;
assign w744 = ~w236 & w738;
assign w745 = (~w239 & w738) | (~w239 & w1776) | (w738 & w1776);
assign w746 = ~w744 & w745;
assign v323 = ~(w743 | w746);
assign w747 = v323;
assign w748 = ~w332 & w640;
assign v324 = ~(w641 | w748);
assign w749 = v324;
assign w750 = (~w321 & ~w749) | (~w321 & w1777) | (~w749 & w1777);
assign w751 = ~w747 & w750;
assign w752 = w747 & ~w750;
assign v325 = ~(w751 | w752);
assign w753 = v325;
assign w754 = (~w235 & w738) | (~w235 & w1849) | (w738 & w1849);
assign w755 = ~w347 & w738;
assign w756 = ~w314 & w341;
assign w757 = w314 & ~w341;
assign v326 = ~(w756 | w757);
assign w758 = v326;
assign w759 = w658 & ~w758;
assign w760 = ~w658 & w758;
assign v327 = ~(w344 | w759);
assign w761 = v327;
assign w762 = ~w760 & w761;
assign v328 = ~(w755 | w762);
assign w763 = v328;
assign v329 = ~(w314 | w658);
assign w764 = v329;
assign w765 = w314 & w658;
assign v330 = ~(w764 | w765);
assign w766 = v330;
assign w767 = w341 & ~w766;
assign w768 = w278 & w766;
assign v331 = ~(w767 | w768);
assign w769 = v331;
assign w770 = w763 & ~w769;
assign w771 = ~w763 & w769;
assign v332 = ~(w770 | w771);
assign w772 = v332;
assign w773 = w754 & ~w772;
assign w774 = ~w754 & w772;
assign v333 = ~(w773 | w774);
assign w775 = v333;
assign w776 = w753 & ~w775;
assign w777 = ~w753 & w775;
assign v334 = ~(w776 | w777);
assign w778 = v334;
assign w779 = ~w735 & w778;
assign w780 = w735 & ~w778;
assign v335 = ~(w779 | w780);
assign w781 = v335;
assign w782 = w652 & w781;
assign v336 = ~(w652 | w781);
assign w783 = v336;
assign v337 = ~(w782 | w783);
assign w784 = v337;
assign v338 = ~(w422 | w440);
assign w785 = v338;
assign w786 = w368 & w410;
assign v339 = ~(w368 | w410);
assign w787 = v339;
assign v340 = ~(w786 | w787);
assign w788 = v340;
assign v341 = ~(w371 | w788);
assign w789 = v341;
assign w790 = ~w404 & w788;
assign v342 = ~(w789 | w790);
assign w791 = v342;
assign w792 = w371 & w788;
assign v343 = ~(w789 | w792);
assign w793 = v343;
assign w794 = (~w378 & ~w793) | (~w378 & w1778) | (~w793 & w1778);
assign v344 = ~(w791 | w794);
assign w795 = v344;
assign w796 = w791 & w794;
assign v345 = ~(w795 | w796);
assign w797 = v345;
assign w798 = w113 & w365;
assign v346 = ~(w113 | w365);
assign w799 = v346;
assign v347 = ~(w798 | w799);
assign w800 = v347;
assign v348 = ~(w80 | w800);
assign w801 = v348;
assign w802 = ~w56 & w800;
assign v349 = ~(w801 | w802);
assign w803 = v349;
assign w804 = ~w368 & w392;
assign w805 = (~w391 & w368) | (~w391 & w1850) | (w368 & w1850);
assign w806 = ~w803 & w805;
assign w807 = w803 & ~w805;
assign v350 = ~(w806 | w807);
assign w808 = v350;
assign w809 = w368 & ~w392;
assign v351 = ~(w804 | w809);
assign w810 = v351;
assign w811 = (~w399 & ~w810) | (~w399 & w1851) | (~w810 & w1851);
assign w812 = w808 & ~w811;
assign w813 = ~w808 & w811;
assign v352 = ~(w812 | w813);
assign w814 = v352;
assign w815 = w797 & w814;
assign v353 = ~(w797 | w814);
assign w816 = v353;
assign v354 = ~(w815 | w816);
assign w817 = v354;
assign w818 = w785 & w817;
assign w819 = ~w784 & w818;
assign w820 = w785 & ~w817;
assign w821 = w784 & w820;
assign v355 = ~(w819 | w821);
assign w822 = v355;
assign w823 = ~w383 & w422;
assign w824 = w817 & w823;
assign w825 = ~w784 & w824;
assign w826 = ~w817 & w823;
assign w827 = w784 & w826;
assign v356 = ~(w825 | w827);
assign w828 = v356;
assign v357 = ~(w785 | w823);
assign w829 = v357;
assign w830 = w817 & w829;
assign w831 = w784 & ~w830;
assign w832 = ~w817 & w829;
assign v358 = ~(w784 | w832);
assign w833 = v358;
assign v359 = ~(w831 | w833);
assign w834 = v359;
assign w835 = w828 & ~w834;
assign w836 = w605 & w822;
assign w837 = w835 & w836;
assign v360 = ~(w606 | w837);
assign w838 = v360;
assign w839 = w432 & w822;
assign w840 = w835 & w839;
assign v361 = ~(w838 | w840);
assign w841 = v361;
assign w842 = w422 & w1852;
assign w843 = (~w437 & ~w422) | (~w437 & w1812) | (~w422 & w1812);
assign w844 = (~w842 & ~w829) | (~w842 & w1853) | (~w829 & w1853);
assign w845 = (~w433 & ~w452) | (~w433 & w1813) | (~w452 & w1813);
assign w846 = ~w844 & w845;
assign w847 = w844 & ~w845;
assign v362 = ~(w846 | w847);
assign w848 = v362;
assign v363 = ~(w605 | w848);
assign w849 = v363;
assign w850 = ~w817 & w849;
assign w851 = w784 & ~w850;
assign w852 = ~w605 & w848;
assign w853 = ~w817 & w852;
assign v364 = ~(w784 | w853);
assign w854 = v364;
assign v365 = ~(w851 | w854);
assign w855 = v365;
assign w856 = w817 & w852;
assign w857 = w784 & ~w856;
assign w858 = w817 & w849;
assign v366 = ~(w784 | w858);
assign w859 = v366;
assign v367 = ~(w857 | w859);
assign w860 = v367;
assign v368 = ~(w855 | w860);
assign w861 = v368;
assign w862 = w455 & ~w458;
assign w863 = ~w455 & w458;
assign v369 = ~(w862 | w863);
assign w864 = v369;
assign w865 = ~w461 & w864;
assign w866 = (~w464 & w864) | (~w464 & w1854) | (w864 & w1854);
assign v370 = ~(w865 | w866);
assign w867 = v370;
assign w868 = (~w46 & w452) | (~w46 & w1855) | (w452 & w1855);
assign w869 = w455 & w2029;
assign w870 = ~w455 & w1856;
assign w871 = (~w868 & w455) | (~w868 & w1857) | (w455 & w1857);
assign v371 = ~(w870 | w871);
assign w872 = v371;
assign w873 = (~w869 & ~w872) | (~w869 & w2030) | (~w872 & w2030);
assign w874 = w867 & ~w873;
assign w875 = ~w867 & w873;
assign v372 = ~(w874 | w875);
assign w876 = v372;
assign w877 = w861 & ~w876;
assign w878 = ~w861 & w876;
assign v373 = ~(w877 | w878);
assign w879 = v373;
assign w880 = w841 & w879;
assign v374 = ~(w841 | w879);
assign w881 = v374;
assign v375 = ~(w880 | w881);
assign w882 = v375;
assign w883 = w488 & w506;
assign v376 = ~(w488 | w506);
assign w884 = v376;
assign v377 = ~(w883 | w884);
assign w885 = v377;
assign w886 = (~w496 & ~w885) | (~w496 & w1814) | (~w885 & w1814);
assign w887 = (~w504 & ~w488) | (~w504 & w1840) | (~w488 & w1840);
assign w888 = (~w37 & w473) | (~w37 & w1858) | (w473 & w1858);
assign w889 = (w476 & w1859) | (w476 & w1860) | (w1859 & w1860);
assign w890 = (~w476 & w1861) | (~w476 & w1862) | (w1861 & w1862);
assign v378 = ~(w889 | w890);
assign w891 = v378;
assign w892 = w887 & ~w891;
assign w893 = ~w887 & w891;
assign v379 = ~(w892 | w893);
assign w894 = v379;
assign w895 = w886 & ~w894;
assign w896 = ~w886 & w894;
assign v380 = ~(w895 | w896);
assign w897 = v380;
assign w898 = w882 & w897;
assign v381 = ~(w882 | w897);
assign w899 = v381;
assign v382 = ~(w898 | w899);
assign w900 = v382;
assign w901 = w601 & w900;
assign v383 = ~(w601 | w900);
assign w902 = v383;
assign v384 = ~(w901 | w902);
assign w903 = v384;
assign v385 = ~(w515 | w518);
assign w904 = v385;
assign w905 = w903 & w904;
assign v386 = ~(w903 | w904);
assign w906 = v386;
assign v387 = ~(w905 | w906);
assign w907 = v387;
assign w908 = (~w18 & w527) | (~w18 & w1863) | (w527 & w1863);
assign w909 = w600 & w903;
assign w910 = (~w908 & ~w903) | (~w908 & w1864) | (~w903 & w1864);
assign w911 = (w910 & w907) | (w910 & w1865) | (w907 & w1865);
assign w912 = (w908 & w903) | (w908 & w1866) | (w903 & w1866);
assign w913 = (w912 & ~w907) | (w912 & w2031) | (~w907 & w2031);
assign w914 = (~w540 & ~w533) | (~w540 & w1867) | (~w533 & w1867);
assign w915 = (~w9 & w530) | (~w9 & w1868) | (w530 & w1868);
assign w916 = (w533 & w1869) | (w533 & w1870) | (w1869 & w1870);
assign w917 = (~w533 & w1871) | (~w533 & w1872) | (w1871 & w1872);
assign v388 = ~(w916 | w917);
assign w918 = v388;
assign w919 = ~w913 & w1873;
assign w920 = (~w918 & w913) | (~w918 & w1874) | (w913 & w1874);
assign v389 = ~(w919 | w920);
assign w921 = v389;
assign v390 = ~(w599 | w921);
assign w922 = v390;
assign w923 = w599 & w921;
assign v391 = ~(w922 | w923);
assign w924 = v391;
assign w925 = ~w557 & w1875;
assign w926 = (~w567 & w560) | (~w567 & w1779) | (w560 & w1779);
assign w927 = (~w560 & w2032) | (~w560 & w2033) | (w2032 & w2033);
assign w928 = w924 & ~w927;
assign w929 = ~w924 & w927;
assign v392 = ~(w928 | w929);
assign w930 = v392;
assign v393 = ~(w577 | w930);
assign w931 = v393;
assign w932 = w577 & w930;
assign v394 = ~(w931 | w932);
assign w933 = v394;
assign w934 = (~w582 & ~w584) | (~w582 & w1780) | (~w584 & w1780);
assign v395 = ~(w933 | w934);
assign w935 = v395;
assign w936 = (~w577 & ~w578) | (~w577 & w1878) | (~w578 & w1878);
assign w937 = w930 & ~w936;
assign w938 = (~w937 & w934) | (~w937 & w1879) | (w934 & w1879);
assign w939 = w594 & ~w938;
assign w940 = w933 & w934;
assign w941 = ~w594 & w1880;
assign v396 = ~(w939 | w941);
assign w942 = v396;
assign w943 = ~w913 & w1881;
assign w944 = ~w5 & w530;
assign w945 = w943 & ~w944;
assign w946 = (~w915 & w913) | (~w915 & w1882) | (w913 & w1882);
assign v397 = ~(w943 | w946);
assign w947 = v397;
assign w948 = w914 & w947;
assign v398 = ~(w945 | w948);
assign w949 = v398;
assign w950 = ~w26 & w512;
assign w951 = w900 & w1883;
assign w952 = (~w951 & ~w903) | (~w951 & w1884) | (~w903 & w1884);
assign v399 = ~(w882 | w891);
assign w953 = v399;
assign w954 = w882 & w891;
assign v400 = ~(w953 | w954);
assign w955 = v400;
assign w956 = w887 & w955;
assign w957 = ~w482 & w488;
assign w958 = ~w955 & w957;
assign v401 = ~(w956 | w958);
assign w959 = v401;
assign w960 = w900 & w950;
assign w961 = w882 & w894;
assign v402 = ~(w882 | w894);
assign w962 = v402;
assign v403 = ~(w961 | w962);
assign w963 = v403;
assign w964 = w886 & ~w963;
assign v404 = ~(w960 | w964);
assign w965 = v404;
assign w966 = w959 & ~w965;
assign w967 = ~w959 & w965;
assign v405 = ~(w966 | w967);
assign w968 = v405;
assign w969 = w784 & w817;
assign v406 = ~(w784 | w817);
assign w970 = v406;
assign v407 = ~(w969 | w970);
assign w971 = v407;
assign w972 = w844 & w971;
assign v408 = ~(w844 | w971);
assign w973 = v408;
assign v409 = ~(w972 | w973);
assign w974 = v409;
assign w975 = w845 & w974;
assign w976 = w838 & ~w975;
assign w977 = w840 & w861;
assign w978 = ~w606 & w861;
assign w979 = ~w837 & w978;
assign v410 = ~(w977 | w979);
assign w980 = v410;
assign w981 = (~w871 & ~w980) | (~w871 & w1816) | (~w980 & w1816);
assign w982 = ~w976 & w981;
assign w983 = w976 & ~w981;
assign v411 = ~(w982 | w983);
assign w984 = v411;
assign w985 = ~w395 & w810;
assign w986 = w790 & w985;
assign w987 = w649 & w807;
assign v412 = ~(w803 | w805);
assign w988 = v412;
assign w989 = ~w649 & w988;
assign v413 = ~(w987 | w989);
assign w990 = v413;
assign w991 = w631 & w990;
assign w992 = w649 & w988;
assign w993 = ~w649 & w807;
assign v414 = ~(w992 | w993);
assign w994 = v414;
assign w995 = ~w631 & w994;
assign v415 = ~(w991 | w995);
assign w996 = v415;
assign v416 = ~(w781 | w996);
assign w997 = v416;
assign w998 = w631 & w994;
assign w999 = ~w631 & w990;
assign v417 = ~(w998 | w999);
assign w1000 = v417;
assign w1001 = w781 & ~w1000;
assign v418 = ~(w997 | w1001);
assign w1002 = v418;
assign w1003 = ~w652 & w806;
assign w1004 = ~w790 & w811;
assign w1005 = w652 & w803;
assign v419 = ~(w781 | w1005);
assign w1006 = v419;
assign w1007 = w781 & w1005;
assign w1008 = (w805 & w652) | (w805 & w1781) | (w652 & w1781);
assign w1009 = ~w1006 & w1008;
assign w1010 = ~w1007 & w1009;
assign w1011 = (~w1004 & ~w1003) | (~w1004 & w1782) | (~w1003 & w1782);
assign w1012 = ~w1002 & w1011;
assign w1013 = (~w986 & w1010) | (~w986 & w1783) | (w1010 & w1783);
assign w1014 = ~w784 & w802;
assign v420 = ~(w1002 | w1014);
assign w1015 = v420;
assign v421 = ~(w1013 | w1015);
assign w1016 = v421;
assign w1017 = w1013 & w1015;
assign v422 = ~(w1016 | w1017);
assign w1018 = v422;
assign w1019 = (~w790 & ~w794) | (~w790 & w1885) | (~w794 & w1885);
assign w1020 = w784 & w814;
assign v423 = ~(w784 | w814);
assign w1021 = v423;
assign v424 = ~(w1020 | w1021);
assign w1022 = v424;
assign w1023 = ~w1019 & w1022;
assign v425 = ~(w795 | w1022);
assign w1024 = v425;
assign v426 = ~(w1023 | w1024);
assign w1025 = v426;
assign w1026 = w634 & w801;
assign w1027 = ~w646 & w778;
assign w1028 = w646 & ~w778;
assign v427 = ~(w1027 | w1028);
assign w1029 = v427;
assign w1030 = w735 & w1029;
assign v428 = ~(w735 | w1029);
assign w1031 = v428;
assign v429 = ~(w1030 | w1031);
assign w1032 = v429;
assign w1033 = w1032 & w1784;
assign v430 = ~(w634 | w801);
assign w1034 = v430;
assign w1035 = (~w1034 & w1032) | (~w1034 & w1785) | (w1032 & w1785);
assign w1036 = ~w1033 & w1035;
assign w1037 = ~w616 & w631;
assign w1038 = ~w1032 & w1037;
assign v431 = ~(w616 | w631);
assign w1039 = v431;
assign w1040 = w1032 & w1039;
assign v432 = ~(w1038 | w1040);
assign w1041 = v432;
assign w1042 = w610 & ~w628;
assign w1043 = w1032 & ~w1042;
assign w1044 = w610 & w628;
assign v433 = ~(w1032 | w1044);
assign w1045 = v433;
assign v434 = ~(w1043 | w1045);
assign w1046 = v434;
assign w1047 = w1041 & ~w1046;
assign w1048 = w1036 & w1047;
assign v435 = ~(w1036 | w1047);
assign w1049 = v435;
assign v436 = ~(w1048 | w1049);
assign w1050 = v436;
assign w1051 = w1025 & ~w1050;
assign w1052 = ~w1025 & w1050;
assign v437 = ~(w1051 | w1052);
assign w1053 = v437;
assign v438 = ~(w1018 | w1053);
assign w1054 = v438;
assign w1055 = w1018 & w1053;
assign v439 = ~(w1054 | w1055);
assign w1056 = v439;
assign w1057 = (~w842 & ~w971) | (~w842 & w1886) | (~w971 & w1886);
assign w1058 = ~w83 & w624;
assign w1059 = w614 & w1058;
assign w1060 = w622 & ~w735;
assign w1061 = ~w1029 & w1060;
assign w1062 = w622 & w735;
assign w1063 = w1029 & w1062;
assign v440 = ~(w1061 | w1063);
assign w1064 = v440;
assign w1065 = ~w614 & w625;
assign v441 = ~(w622 | w1065);
assign w1066 = v441;
assign w1067 = w1032 & w1066;
assign w1068 = (~w1059 & w1064) | (~w1059 & w1786) | (w1064 & w1786);
assign w1069 = ~w1067 & w1068;
assign w1070 = w747 & w775;
assign v442 = ~(w747 | w775);
assign w1071 = v442;
assign v443 = ~(w1070 | w1071);
assign w1072 = v443;
assign w1073 = ~w735 & w1072;
assign w1074 = w735 & ~w1072;
assign v444 = ~(w1073 | w1074);
assign w1075 = v444;
assign w1076 = w742 & ~w746;
assign w1077 = ~w218 & w1076;
assign v445 = ~(w1075 | w1077);
assign w1078 = v445;
assign w1079 = ~w643 & w1075;
assign v446 = ~(w1078 | w1079);
assign w1080 = v446;
assign w1081 = w330 & w640;
assign w1082 = (w640 & w1887) | (w640 & w1888) | (w1887 & w1888);
assign v447 = ~(w1081 | w1082);
assign w1083 = v447;
assign w1084 = w643 & w1083;
assign w1085 = w1073 & w1084;
assign w1086 = ~w1072 & w1084;
assign w1087 = ~w317 & w331;
assign w1088 = ~w640 & w1087;
assign w1089 = (~w1088 & ~w1086) | (~w1088 & w1787) | (~w1086 & w1787);
assign w1090 = ~w1085 & w1089;
assign w1091 = ~w643 & w1083;
assign w1092 = w1075 & w1091;
assign w1093 = w1090 & ~w1092;
assign v448 = ~(w1080 | w1093);
assign w1094 = v448;
assign w1095 = w1080 & w1090;
assign v449 = ~(w1094 | w1095);
assign w1096 = v449;
assign w1097 = ~w1069 & w1096;
assign w1098 = w1069 & ~w1096;
assign v450 = ~(w1097 | w1098);
assign w1099 = v450;
assign w1100 = (~w670 & w732) | (~w670 & w1889) | (w732 & w1889);
assign w1101 = (~w700 & w694) | (~w700 & w1817) | (w694 & w1817);
assign w1102 = (w678 & w681) | (w678 & w2034) | (w681 & w2034);
assign w1103 = (~w689 & ~w691) | (~w689 & w1818) | (~w691 & w1818);
assign w1104 = w1102 & w1103;
assign v451 = ~(w1102 | w1103);
assign w1105 = v451;
assign v452 = ~(w1104 | w1105);
assign w1106 = v452;
assign w1107 = ~w1101 & w1106;
assign w1108 = w1101 & ~w1106;
assign v453 = ~(w1107 | w1108);
assign w1109 = v453;
assign w1110 = ~w299 & w658;
assign w1111 = w710 & ~w1110;
assign w1112 = ~w710 & w1110;
assign w1113 = (~w1111 & ~w704) | (~w1111 & w1819) | (~w704 & w1819);
assign w1114 = ~w1109 & w1113;
assign w1115 = w1109 & ~w1113;
assign v454 = ~(w1114 | w1115);
assign w1116 = v454;
assign w1117 = w662 & w726;
assign w1118 = ~w720 & w1117;
assign w1119 = w662 & ~w726;
assign w1120 = w720 & w1119;
assign v455 = ~(w1118 | w1120);
assign w1121 = v455;
assign w1122 = w1116 & ~w1121;
assign w1123 = ~w1116 & w1121;
assign v456 = ~(w1122 | w1123);
assign w1124 = v456;
assign w1125 = w723 & w1890;
assign w1126 = w715 & ~w1110;
assign v457 = ~(w1125 | w1126);
assign w1127 = v457;
assign w1128 = ~w720 & w1127;
assign v458 = ~(w724 | w726);
assign w1129 = v458;
assign w1130 = w720 & w1129;
assign v459 = ~(w1128 | w1130);
assign w1131 = v459;
assign w1132 = w1124 & ~w1131;
assign w1133 = ~w1124 & w1131;
assign v460 = ~(w1132 | w1133);
assign w1134 = v460;
assign v461 = ~(w1100 | w1134);
assign w1135 = v461;
assign w1136 = w1100 & w1134;
assign v462 = ~(w1135 | w1136);
assign w1137 = v462;
assign w1138 = (~w770 & w735) | (~w770 & w1891) | (w735 & w1891);
assign w1139 = w235 & ~w239;
assign w1140 = ~w738 & w1139;
assign w1141 = ~w746 & w754;
assign w1142 = (~w1141 & w735) | (~w1141 & w1820) | (w735 & w1820);
assign w1143 = w772 & ~w1140;
assign w1144 = w735 & w1143;
assign w1145 = w1142 & ~w1144;
assign w1146 = w1138 & w1145;
assign v463 = ~(w1137 | w1146);
assign w1147 = v463;
assign w1148 = ~w1138 & w1142;
assign w1149 = w1137 & ~w1148;
assign v464 = ~(w1147 | w1149);
assign w1150 = v464;
assign v465 = ~(w1138 | w1142);
assign w1151 = v465;
assign v466 = ~(w1137 | w1151);
assign w1152 = v466;
assign w1153 = w1138 & ~w1145;
assign w1154 = w1137 & ~w1153;
assign v467 = ~(w1152 | w1154);
assign w1155 = v467;
assign v468 = ~(w1150 | w1155);
assign w1156 = v468;
assign w1157 = ~w317 & w749;
assign v469 = ~(w750 | w1157);
assign w1158 = v469;
assign v470 = ~(w735 | w1158);
assign w1159 = v470;
assign w1160 = w1029 & ~w1159;
assign w1161 = w735 & ~w1158;
assign v471 = ~(w1029 | w1161);
assign w1162 = v471;
assign v472 = ~(w1160 | w1162);
assign w1163 = v472;
assign w1164 = w1064 & ~w1163;
assign w1165 = w1156 & ~w1164;
assign w1166 = ~w1156 & w1164;
assign v473 = ~(w1165 | w1166);
assign w1167 = v473;
assign w1168 = w1099 & ~w1167;
assign w1169 = ~w1099 & w1167;
assign v474 = ~(w1168 | w1169);
assign w1170 = v474;
assign w1171 = w1057 & ~w1170;
assign w1172 = ~w1057 & w1170;
assign v475 = ~(w1171 | w1172);
assign w1173 = v475;
assign w1174 = w1056 & w1173;
assign v476 = ~(w1056 | w1173);
assign w1175 = v476;
assign v477 = ~(w1174 | w1175);
assign w1176 = v477;
assign v478 = ~(w984 | w1176);
assign w1177 = v478;
assign w1178 = w984 & w1176;
assign v479 = ~(w1177 | w1178);
assign w1179 = v479;
assign w1180 = w861 & ~w872;
assign w1181 = ~w861 & w872;
assign v480 = ~(w1180 | w1181);
assign w1182 = v480;
assign w1183 = w841 & ~w1182;
assign w1184 = ~w841 & w1182;
assign v481 = ~(w1183 | w1184);
assign w1185 = v481;
assign w1186 = w865 & w1185;
assign w1187 = w868 & ~w980;
assign w1188 = (w862 & ~w980) | (w862 & w1821) | (~w980 & w1821);
assign w1189 = ~w1187 & w1188;
assign v482 = ~(w1186 | w1189);
assign w1190 = v482;
assign w1191 = w37 & ~w479;
assign w1192 = ~w473 & w1191;
assign v483 = ~(w882 | w1192);
assign w1193 = v483;
assign w1194 = (~w479 & ~w473) | (~w479 & w1892) | (~w473 & w1892);
assign w1195 = w888 & ~w1194;
assign w1196 = w882 & w1195;
assign v484 = ~(w1193 | w1196);
assign w1197 = v484;
assign w1198 = ~w1190 & w1197;
assign w1199 = ~w865 & w866;
assign w1200 = (w1199 & w1185) | (w1199 & w1822) | (w1185 & w1822);
assign w1201 = w1190 & ~w1200;
assign w1202 = ~w1197 & w1201;
assign v485 = ~(w1198 | w1202);
assign w1203 = v485;
assign w1204 = w1179 & ~w1203;
assign w1205 = ~w1179 & w1203;
assign v486 = ~(w1204 | w1205);
assign w1206 = v486;
assign w1207 = ~w968 & w1206;
assign w1208 = w968 & ~w1206;
assign v487 = ~(w1207 | w1208);
assign w1209 = v487;
assign w1210 = w952 & ~w1209;
assign w1211 = ~w952 & w1209;
assign v488 = ~(w1210 | w1211);
assign w1212 = v488;
assign w1213 = (~w907 & w2035) | (~w907 & w2036) | (w2035 & w2036);
assign w1214 = (w907 & w2037) | (w907 & w2038) | (w2037 & w2038);
assign w1215 = w1213 & ~w1214;
assign w1216 = w1212 & ~w1215;
assign w1217 = ~w1212 & w1215;
assign v489 = ~(w1216 | w1217);
assign w1218 = v489;
assign w1219 = ~w949 & w1218;
assign w1220 = w949 & ~w1218;
assign v490 = ~(w1219 | w1220);
assign w1221 = v490;
assign w1222 = w558 & w924;
assign w1223 = (~w922 & ~w924) | (~w922 & w1823) | (~w924 & w1823);
assign w1224 = w1221 & w1223;
assign v491 = ~(w1221 | w1223);
assign w1225 = v491;
assign v492 = ~(w1224 | w1225);
assign w1226 = v492;
assign w1227 = w937 & ~w1226;
assign w1228 = (~w935 & w594) | (~w935 & w1788) | (w594 & w1788);
assign w1229 = w926 & ~w930;
assign w1230 = w1226 & ~w1229;
assign w1231 = ~w1226 & w1229;
assign v493 = ~(w1230 | w1231);
assign w1232 = v493;
assign w1233 = w1228 & w1232;
assign w1234 = (~w1227 & ~w1228) | (~w1227 & w1894) | (~w1228 & w1894);
assign v494 = ~(w937 | w1232);
assign w1235 = v494;
assign w1236 = ~w1228 & w1235;
assign w1237 = w1234 & ~w1236;
assign w1238 = w425 & w604;
assign w1239 = (~w428 & w604) | (~w428 & w1895) | (w604 & w1895);
assign w1240 = ~w1238 & w1239;
assign w1241 = w974 & w1240;
assign v495 = ~(w837 | w1241);
assign w1242 = v495;
assign w1243 = ~w976 & w1242;
assign w1244 = ~w41 & w452;
assign w1245 = ~w980 & w1244;
assign v496 = ~(w1243 | w1245);
assign w1246 = v496;
assign w1247 = (~w1246 & ~w1176) | (~w1246 & w1896) | (~w1176 & w1896);
assign w1248 = w976 & w1176;
assign v497 = ~(w976 | w1176);
assign w1249 = v497;
assign v498 = ~(w1248 | w1249);
assign w1250 = v498;
assign w1251 = w981 & ~w1245;
assign w1252 = (~w1247 & ~w1250) | (~w1247 & w1897) | (~w1250 & w1897);
assign w1253 = (~w789 & ~w793) | (~w789 & w2039) | (~w793 & w2039);
assign w1254 = w1022 & ~w1253;
assign w1255 = w793 & w1899;
assign w1256 = ~w1022 & w1255;
assign v499 = ~(w1254 | w1256);
assign w1257 = v499;
assign w1258 = w1025 & w1257;
assign w1259 = w828 & ~w1258;
assign v500 = ~(w1018 | w1050);
assign w1260 = v500;
assign w1261 = w1018 & w1050;
assign v501 = ~(w1260 | w1261);
assign w1262 = v501;
assign w1263 = w1170 & w1262;
assign v502 = ~(w1170 | w1262);
assign w1264 = v502;
assign v503 = ~(w1263 | w1264);
assign w1265 = v503;
assign w1266 = ~w1259 & w1265;
assign w1267 = w1050 & ~w1257;
assign w1268 = w1018 & ~w1267;
assign v504 = ~(w1050 | w1257);
assign w1269 = v504;
assign v505 = ~(w1018 | w1269);
assign w1270 = v505;
assign v506 = ~(w1268 | w1270);
assign w1271 = v506;
assign w1272 = w1170 & w1271;
assign w1273 = w1018 & w1269;
assign w1274 = ~w1018 & w1267;
assign v507 = ~(w1273 | w1274);
assign w1275 = v507;
assign v508 = ~(w1170 | w1275);
assign w1276 = v508;
assign v509 = ~(w1272 | w1276);
assign w1277 = v509;
assign w1278 = w784 & ~w803;
assign w1279 = (~w391 & w784) | (~w391 & w1900) | (w784 & w1900);
assign w1280 = ~w1278 & w1279;
assign w1281 = w985 & ~w1280;
assign w1282 = ~w1280 & w1901;
assign v510 = ~(w1013 | w1282);
assign w1283 = v510;
assign w1284 = w1015 & ~w1050;
assign w1285 = ~w1015 & w1050;
assign v511 = ~(w1284 | w1285);
assign w1286 = v511;
assign w1287 = w1283 & ~w1286;
assign w1288 = w1170 & ~w1287;
assign w1289 = w1283 & w1286;
assign v512 = ~(w1170 | w1289);
assign w1290 = v512;
assign v513 = ~(w1288 | w1290);
assign w1291 = v513;
assign w1292 = w1277 & ~w1291;
assign w1293 = ~w1266 & w1292;
assign w1294 = ~w785 & w843;
assign w1295 = w835 & w1294;
assign w1296 = (w822 & ~w835) | (w822 & w1902) | (~w835 & w1902);
assign w1297 = w1056 & w1170;
assign v514 = ~(w1056 | w1170);
assign w1298 = v514;
assign v515 = ~(w1297 | w1298);
assign w1299 = v515;
assign v516 = ~(w1296 | w1299);
assign w1300 = v516;
assign w1301 = w1293 & ~w1300;
assign w1302 = w218 & ~w1076;
assign w1303 = (~w209 & ~w1076) | (~w209 & w1903) | (~w1076 & w1903);
assign w1304 = w1075 & ~w1303;
assign w1305 = (~w1302 & w1075) | (~w1302 & w1824) | (w1075 & w1824);
assign w1306 = ~w1304 & w1305;
assign w1307 = w735 & w769;
assign v517 = ~(w735 | w769);
assign w1308 = v517;
assign w1309 = (w755 & ~w735) | (w755 & w1904) | (~w735 & w1904);
assign w1310 = ~w1308 & w1309;
assign w1311 = w1137 & w1310;
assign v518 = ~(w1306 | w1311);
assign w1312 = v518;
assign w1313 = ~w1150 & w1312;
assign w1314 = w1155 & ~w1311;
assign v519 = ~(w1313 | w1314);
assign w1315 = v519;
assign v520 = ~(w1104 | w1107);
assign w1316 = v520;
assign v521 = ~(w1114 | w1316);
assign w1317 = v521;
assign w1318 = w1105 & w1114;
assign v522 = ~(w1317 | w1318);
assign w1319 = v522;
assign w1320 = w1123 & ~w1131;
assign w1321 = ~w254 & w664;
assign w1322 = ~w732 & w1321;
assign w1323 = ~w1320 & w1322;
assign w1324 = ~w1123 & w1131;
assign v523 = ~(w1122 | w1324);
assign w1325 = v523;
assign w1326 = ~w1323 & w1325;
assign w1327 = ~w1319 & w1326;
assign w1328 = w1319 & ~w1326;
assign v524 = ~(w1327 | w1328);
assign w1329 = v524;
assign v525 = ~(w269 | w668);
assign w1330 = v525;
assign w1331 = (~w1330 & w732) | (~w1330 & w1905) | (w732 & w1905);
assign w1332 = w665 & w732;
assign v526 = ~(w1322 | w1332);
assign w1333 = v526;
assign w1334 = ~w1331 & w1333;
assign w1335 = ~w1134 & w1334;
assign w1336 = w1329 & ~w1335;
assign w1337 = ~w1329 & w1335;
assign v527 = ~(w1336 | w1337);
assign w1338 = v527;
assign w1339 = ~w1134 & w1906;
assign w1340 = (w762 & w735) | (w762 & w1907) | (w735 & w1907);
assign v528 = ~(w1307 | w1340);
assign w1341 = v528;
assign w1342 = (~w1339 & ~w1137) | (~w1339 & w1908) | (~w1137 & w1908);
assign w1343 = w1338 & ~w1342;
assign w1344 = ~w1338 & w1342;
assign v529 = ~(w1343 | w1344);
assign w1345 = v529;
assign w1346 = w1315 & ~w1345;
assign w1347 = ~w1315 & w1345;
assign v530 = ~(w1346 | w1347);
assign w1348 = v530;
assign w1349 = ~w1029 & w1062;
assign w1350 = (w1058 & ~w1029) | (w1058 & w1789) | (~w1029 & w1789);
assign w1351 = ~w1349 & w1350;
assign w1352 = ~w1164 & w1790;
assign w1353 = w1080 & ~w1352;
assign w1354 = ~w1156 & w1353;
assign w1355 = (~w1093 & w1164) | (~w1093 & w1791) | (w1164 & w1791);
assign w1356 = ~w212 & w640;
assign w1357 = w1072 & w1356;
assign w1358 = w735 & w1357;
assign w1359 = ~w1072 & w1356;
assign w1360 = ~w735 & w1359;
assign v531 = ~(w1358 | w1360);
assign w1361 = v531;
assign w1362 = ~w1361 & w1146;
assign w1363 = w1137 & w1362;
assign w1364 = ~w1361 & w1153;
assign w1365 = ~w1137 & w1364;
assign v532 = ~(w1137 | w1145);
assign w1366 = v532;
assign w1367 = w1137 & w1145;
assign v533 = ~(w1138 | w1361);
assign w1368 = v533;
assign w1369 = ~w1366 & w1368;
assign w1370 = ~w1367 & w1369;
assign v534 = ~(w1080 | w1352);
assign w1371 = v534;
assign w1372 = w1156 & w1371;
assign v535 = ~(w1363 | w1365);
assign w1373 = v535;
assign w1374 = ~w1355 & w1373;
assign w1375 = ~w1370 & w1374;
assign w1376 = w1375 & w1792;
assign w1377 = w1348 & ~w1376;
assign w1378 = ~w1348 & w1376;
assign v536 = ~(w1377 | w1378);
assign w1379 = v536;
assign v537 = ~(w622 | w1032);
assign w1380 = v537;
assign w1381 = w1351 & ~w1380;
assign v538 = ~(w1069 | w1381);
assign w1382 = v538;
assign w1383 = ~w1096 & w1382;
assign v539 = ~(w59 | w609);
assign w1384 = v539;
assign w1385 = ~w614 & w1384;
assign v540 = ~(w610 | w1385);
assign w1386 = v540;
assign w1387 = w628 & w1032;
assign v541 = ~(w628 | w1032);
assign w1388 = v541;
assign v542 = ~(w1387 | w1388);
assign w1389 = v542;
assign w1390 = ~w1386 & w1389;
assign w1391 = w614 & w1384;
assign w1392 = ~w1389 & w1391;
assign v543 = ~(w1390 | w1392);
assign w1393 = v543;
assign v544 = ~(w1099 | w1393);
assign w1394 = v544;
assign w1395 = w1167 & ~w1383;
assign w1396 = ~w1394 & w1395;
assign w1397 = w1096 & w1382;
assign w1398 = w1099 & ~w1393;
assign v545 = ~(w1167 | w1397);
assign w1399 = v545;
assign w1400 = ~w1398 & w1399;
assign v546 = ~(w1396 | w1400);
assign w1401 = v546;
assign w1402 = w1379 & ~w1401;
assign w1403 = ~w1379 & w1401;
assign v547 = ~(w1402 | w1403);
assign w1404 = v547;
assign v548 = ~(w1041 | w1384);
assign w1405 = v548;
assign w1406 = ~w609 & w65;
assign w1407 = w631 & ~w1032;
assign w1408 = (~w68 & ~w609) | (~w68 & w1909) | (~w609 & w1909);
assign w1409 = ~w1406 & w1408;
assign w1410 = (w1409 & ~w1032) | (w1409 & w1910) | (~w1032 & w1910);
assign w1411 = ~w1407 & w1410;
assign v549 = ~(w1405 | w1411);
assign w1412 = v549;
assign v550 = ~(w1170 | w1412);
assign w1413 = v550;
assign w1414 = w1047 & w1911;
assign v551 = ~(w1099 | w1414);
assign w1415 = v551;
assign w1416 = w1036 & ~w1047;
assign w1417 = w1099 & ~w1416;
assign w1418 = ~w1415 & w1793;
assign v552 = ~(w1099 | w1416);
assign w1419 = v552;
assign w1420 = w1099 & ~w1414;
assign v553 = ~(w1167 | w1419);
assign w1421 = v553;
assign w1422 = ~w1420 & w1421;
assign v554 = ~(w1418 | w1422);
assign w1423 = v554;
assign w1424 = ~w1413 & w1423;
assign w1425 = w1015 & ~w1281;
assign v555 = ~(w1050 | w1425);
assign w1426 = v555;
assign w1427 = w1170 & ~w1426;
assign w1428 = w1050 & ~w1425;
assign v556 = ~(w1170 | w1428);
assign w1429 = v556;
assign v557 = ~(w1427 | w1429);
assign w1430 = v557;
assign w1431 = w1424 & ~w1430;
assign w1432 = w1404 & ~w1431;
assign w1433 = ~w1404 & w1431;
assign v558 = ~(w1432 | w1433);
assign w1434 = v558;
assign w1435 = w1301 & w1434;
assign v559 = ~(w1301 | w1434);
assign w1436 = v559;
assign v560 = ~(w1435 | w1436);
assign w1437 = v560;
assign v561 = ~(w1176 | w1242);
assign w1438 = v561;
assign v562 = ~(w1437 | w1438);
assign w1439 = v562;
assign w1440 = w1295 & ~w1299;
assign v563 = ~(w1438 | w1440);
assign w1441 = v563;
assign w1442 = w1293 & w1434;
assign v564 = ~(w1293 | w1434);
assign w1443 = v564;
assign v565 = ~(w1441 | w1442);
assign w1444 = v565;
assign w1445 = ~w1443 & w1444;
assign w1446 = (w1252 & w1439) | (w1252 & w1794) | (w1439 & w1794);
assign w1447 = ~w1252 & w1437;
assign w1448 = w955 & w1912;
assign v566 = ~(w958 | w1448);
assign w1449 = v566;
assign w1450 = w1206 & ~w1449;
assign w1451 = ~w1447 & w1450;
assign w1452 = ~w1446 & w1451;
assign v567 = ~(w491 | w885);
assign w1453 = v567;
assign w1454 = ~w963 & w1453;
assign w1455 = (w1454 & w1206) | (w1454 & w1825) | (w1206 & w1825);
assign w1456 = w1206 & w1826;
assign v568 = ~(w1455 | w1456);
assign w1457 = v568;
assign w1458 = ~w1452 & w1457;
assign v569 = ~(w1446 | w1447);
assign w1459 = v569;
assign v570 = ~(w1179 | w1201);
assign w1460 = v570;
assign w1461 = ~w984 & w1190;
assign w1462 = w1176 & w1461;
assign w1463 = w984 & w1190;
assign w1464 = ~w1176 & w1463;
assign v571 = ~(w1462 | w1464);
assign w1465 = v571;
assign v572 = ~(w35 | w473);
assign w1466 = v572;
assign w1467 = w882 & w1466;
assign w1468 = w1465 & w1467;
assign v573 = ~(w1460 | w1468);
assign w1469 = v573;
assign w1470 = w1179 & w1201;
assign w1471 = w984 & ~w1190;
assign w1472 = w1176 & w1471;
assign v574 = ~(w984 | w1190);
assign w1473 = v574;
assign w1474 = ~w1176 & w1473;
assign v575 = ~(w1472 | w1474);
assign w1475 = v575;
assign w1476 = w882 & ~w888;
assign w1477 = w1197 & ~w1476;
assign w1478 = w1475 & w1477;
assign w1479 = ~w1470 & w1478;
assign w1480 = w1465 & w1475;
assign w1481 = w882 & w1913;
assign w1482 = w1480 & w1481;
assign v576 = ~(w1479 | w1482);
assign w1483 = v576;
assign w1484 = w1469 & w1483;
assign w1485 = w1459 & ~w1484;
assign w1486 = ~w1450 & w1484;
assign w1487 = ~w1459 & w1486;
assign v577 = ~(w1485 | w1487);
assign w1488 = v577;
assign w1489 = ~w1458 & w1488;
assign w1490 = w958 & w1206;
assign w1491 = w1206 & w1827;
assign v578 = ~(w1490 | w1491);
assign w1492 = v578;
assign w1493 = w1453 & ~w1492;
assign w1494 = w1457 & ~w1493;
assign w1495 = ~w1488 & w1494;
assign v579 = ~(w1489 | w1495);
assign w1496 = v579;
assign v580 = ~(w17 | w527);
assign w1497 = v580;
assign w1498 = w911 & w1212;
assign w1499 = w1212 & w1828;
assign w1500 = (~w909 & ~w907) | (~w909 & w1914) | (~w907 & w1914);
assign w1501 = (~w1500 & w1209) | (~w1500 & w1829) | (w1209 & w1829);
assign w1502 = w959 & w960;
assign w1503 = w1206 & w1502;
assign w1504 = ~w959 & w960;
assign w1505 = ~w1206 & w1504;
assign v581 = ~(w1503 | w1505);
assign w1506 = v581;
assign v582 = ~(w494 | w512);
assign w1507 = v582;
assign w1508 = ~w963 & w1507;
assign w1509 = w959 & w1508;
assign w1510 = w1206 & w1509;
assign w1511 = ~w959 & w1508;
assign w1512 = ~w1206 & w1511;
assign v583 = ~(w1510 | w1512);
assign w1513 = v583;
assign w1514 = w1506 & w1513;
assign w1515 = ~w1211 & w1514;
assign w1516 = ~w1501 & w1515;
assign w1517 = w1213 & w1214;
assign w1518 = w1212 & w1517;
assign w1519 = w1516 & ~w1518;
assign w1520 = ~w1499 & w1519;
assign w1521 = w1496 & ~w1520;
assign w1522 = ~w1496 & w1520;
assign v584 = ~(w1521 | w1522);
assign w1523 = v584;
assign w1524 = w1221 & w1222;
assign w1525 = w598 & ~w921;
assign w1526 = w1221 & w1525;
assign v585 = ~(w1524 | w1526);
assign w1527 = v585;
assign w1528 = w597 & ~w921;
assign w1529 = w1221 & w1528;
assign w1530 = (~w1219 & ~w1221) | (~w1219 & w1830) | (~w1221 & w1830);
assign w1531 = (w1523 & ~w1527) | (w1523 & w1831) | (~w1527 & w1831);
assign w1532 = w1527 & w1537;
assign v586 = ~(w1531 | w1532);
assign w1533 = v586;
assign w1534 = (w1533 & ~w1234) | (w1533 & w1915) | (~w1234 & w1915);
assign w1535 = w1234 & w1916;
assign v587 = ~(w1534 | w1535);
assign w1536 = v587;
assign w1537 = ~w1523 & w1530;
assign w1538 = ~w1496 & w1516;
assign w1539 = w1496 & ~w1516;
assign v588 = ~(w1538 | w1539);
assign w1540 = v588;
assign w1541 = w1529 & w1540;
assign v589 = ~(w1526 | w1541);
assign w1542 = v589;
assign v590 = ~(w1537 | w1542);
assign w1543 = v590;
assign v591 = ~(w533 | w536);
assign w1544 = v591;
assign w1545 = w947 & w1544;
assign v592 = ~(w945 | w1545);
assign w1546 = v592;
assign w1547 = w1219 & w1523;
assign w1548 = w1523 & w1917;
assign w1549 = (~w1548 & w1542) | (~w1548 & w1918) | (w1542 & w1918);
assign w1550 = (~w1524 & w1226) | (~w1524 & w1832) | (w1226 & w1832);
assign v593 = ~(w1537 | w1547);
assign w1551 = v593;
assign w1552 = ~w1550 & w1551;
assign w1553 = w1549 & ~w1552;
assign w1554 = w1523 & w1833;
assign w1555 = w1496 & w1498;
assign w1556 = (~w1555 & ~w1540) | (~w1555 & w1834) | (~w1540 & w1834);
assign w1557 = ~w1554 & w1556;
assign w1558 = w909 & w1209;
assign w1559 = w1496 & w1558;
assign w1560 = ~w1211 & w1506;
assign w1561 = w1496 & ~w1560;
assign v594 = ~(w1559 | w1561);
assign w1562 = v594;
assign v595 = ~(w1450 | w1479);
assign w1563 = v595;
assign w1564 = ~w1446 & w1835;
assign w1565 = (w1469 & w1446) | (w1469 & w1836) | (w1446 & w1836);
assign v596 = ~(w1564 | w1565);
assign w1566 = v596;
assign w1567 = ~w1563 & w1566;
assign w1568 = ~w1452 & w1837;
assign w1569 = w1488 & ~w1568;
assign v597 = ~(w1567 | w1569);
assign w1570 = v597;
assign v598 = ~(w1292 | w1434);
assign w1571 = v598;
assign w1572 = ~w1176 & w1243;
assign w1573 = (w1572 & ~w1301) | (w1572 & w1795) | (~w1301 & w1795);
assign w1574 = ~w1571 & w1573;
assign v599 = ~(w1445 | w1574);
assign w1575 = v599;
assign w1576 = w1266 & ~w1434;
assign v600 = ~(w822 | w1299);
assign w1577 = v600;
assign w1578 = ~w1442 & w1577;
assign v601 = ~(w1576 | w1578);
assign w1579 = v601;
assign w1580 = w1575 & w1579;
assign w1581 = (~w1378 & ~w1402) | (~w1378 & w1838) | (~w1402 & w1838);
assign w1582 = w1329 & w1919;
assign w1583 = w1116 & w1131;
assign v602 = ~(w1319 | w1583);
assign w1584 = v602;
assign v603 = ~(w1582 | w1584);
assign w1585 = v603;
assign w1586 = (~w1324 & w2040) | (~w1324 & w2041) | (w2040 & w2041);
assign w1587 = (w1586 & w1338) | (w1586 & w1921) | (w1338 & w1921);
assign w1588 = ~w1585 & w1587;
assign w1589 = ~w1346 & w1588;
assign v604 = ~(w1150 | w1306);
assign w1590 = v604;
assign w1591 = w1587 & w1922;
assign v605 = ~(w1155 | w1590);
assign w1592 = v605;
assign w1593 = ~w1345 & w1592;
assign w1594 = ~w1591 & w1593;
assign v606 = ~(w1589 | w1594);
assign w1595 = v606;
assign w1596 = ~w1581 & w1595;
assign w1597 = w1581 & ~w1595;
assign v607 = ~(w1596 | w1597);
assign w1598 = v607;
assign w1599 = w1050 & ~w1170;
assign w1600 = ~w1050 & w1170;
assign v608 = ~(w1599 | w1600);
assign w1601 = v608;
assign v609 = ~(w1015 | w1601);
assign w1602 = v609;
assign w1603 = (w1423 & w1601) | (w1423 & w1923) | (w1601 & w1923);
assign v610 = ~(w1404 | w1603);
assign w1604 = v610;
assign w1605 = w1598 & ~w1604;
assign w1606 = ~w1598 & w1604;
assign v611 = ~(w1605 | w1606);
assign w1607 = v611;
assign v612 = ~(w1404 | w1424);
assign w1608 = v612;
assign v613 = ~(w1013 | w1265);
assign w1609 = v613;
assign w1610 = w1277 & ~w1609;
assign w1611 = w1404 & w1424;
assign w1612 = ~w1602 & w1611;
assign v614 = ~(w1608 | w1610);
assign w1613 = v614;
assign w1614 = ~w1612 & w1613;
assign w1615 = w1607 & w1614;
assign v615 = ~(w1607 | w1614);
assign w1616 = v615;
assign v616 = ~(w1615 | w1616);
assign w1617 = v616;
assign w1618 = w1580 & ~w1617;
assign w1619 = ~w1580 & w1617;
assign v617 = ~(w1618 | w1619);
assign w1620 = v617;
assign w1621 = ~w1439 & w1796;
assign w1622 = w1187 & w1250;
assign w1623 = w1437 & w1622;
assign w1624 = (~w1623 & ~w1621) | (~w1623 & w1797) | (~w1621 & w1797);
assign w1625 = w1620 & w1624;
assign v618 = ~(w1620 | w1624);
assign w1626 = v618;
assign v619 = ~(w1625 | w1626);
assign w1627 = v619;
assign w1628 = w981 & w1250;
assign w1629 = (w1628 & w1437) | (w1628 & w1924) | (w1437 & w1924);
assign w1630 = (w1437 & w2042) | (w1437 & w2043) | (w2042 & w2043);
assign w1631 = ~w1189 & w1200;
assign v620 = ~(w1186 | w1631);
assign w1632 = v620;
assign w1633 = ~w1439 & w2044;
assign v621 = ~(w1630 | w1633);
assign w1634 = v621;
assign w1635 = w1476 & w1480;
assign w1636 = ~w1446 & w1925;
assign w1637 = w1634 & ~w1636;
assign w1638 = w1627 & w1637;
assign v622 = ~(w1627 | w1637);
assign w1639 = v622;
assign v623 = ~(w1638 | w1639);
assign w1640 = v623;
assign w1641 = w1570 & ~w1640;
assign v624 = ~(w1570 | w1627);
assign w1642 = v624;
assign v625 = ~(w1641 | w1642);
assign w1643 = v625;
assign w1644 = w1562 & ~w1643;
assign w1645 = ~w1562 & w1643;
assign v626 = ~(w1644 | w1645);
assign w1646 = v626;
assign w1647 = w1557 & w1646;
assign v627 = ~(w1557 | w1646);
assign w1648 = v627;
assign v628 = ~(w1647 | w1648);
assign w1649 = v628;
assign w1650 = ~w1553 & w1649;
assign w1651 = w1553 & ~w1649;
assign v629 = ~(w1650 | w1651);
assign w1652 = v629;
assign w1653 = w1228 & w1926;
assign w1654 = w1227 & w1533;
assign v630 = ~(w1653 | w1654);
assign w1655 = v630;
assign w1656 = w1652 & ~w1655;
assign w1657 = ~w1652 & w1655;
assign v631 = ~(w1656 | w1657);
assign w1658 = v631;
assign w1659 = w1548 & ~w1649;
assign w1660 = w10 & w18;
assign w1661 = w903 & w1927;
assign w1662 = (w943 & ~w1209) | (w943 & w2045) | (~w1209 & w2045);
assign w1663 = (w1662 & w1212) | (w1662 & w2046) | (w1212 & w2046);
assign w1664 = w1540 & w1663;
assign w1665 = (~w1555 & ~w1540) | (~w1555 & w1928) | (~w1540 & w1928);
assign w1666 = w1523 & w1929;
assign w1667 = (w1666 & w1646) | (w1666 & w2047) | (w1646 & w2047);
assign w1668 = (~w1667 & w1649) | (~w1667 & w2070) | (w1649 & w2070);
assign v632 = ~(w1555 | w1559);
assign w1669 = v632;
assign w1670 = ~w1664 & w1669;
assign w1671 = (~w1561 & w1641) | (~w1561 & w1798) | (w1641 & w1798);
assign v633 = ~(w1670 | w1671);
assign w1672 = v633;
assign v634 = ~(w1489 | w1567);
assign w1673 = v634;
assign w1674 = w1206 & w1448;
assign w1675 = (~w1674 & ~w1488) | (~w1674 & w1930) | (~w1488 & w1930);
assign v635 = ~(w1673 | w1675);
assign w1676 = v635;
assign w1677 = w1640 & w1676;
assign w1678 = (w1490 & w1566) | (w1490 & w1799) | (w1566 & w1799);
assign w1679 = w1488 & ~w1513;
assign v636 = ~(w1678 | w1679);
assign w1680 = v636;
assign w1681 = ~w1446 & w1931;
assign w1682 = (w1681 & ~w1627) | (w1681 & w1932) | (~w1627 & w1932);
assign w1683 = (~w1682 & ~w1640) | (~w1682 & w2048) | (~w1640 & w2048);
assign w1684 = ~w1677 & w1683;
assign w1685 = w1496 & ~w1642;
assign w1686 = ~w1641 & w1685;
assign w1687 = w905 & w1209;
assign w1688 = w1686 & w1687;
assign w1689 = w1684 & ~w1688;
assign w1690 = ~w1672 & w1689;
assign w1691 = w951 & w1209;
assign w1692 = w1506 & ~w1691;
assign w1693 = w1686 & ~w1692;
assign w1694 = ~w1439 & w2049;
assign w1695 = ~w1627 & w1694;
assign w1696 = ~w1446 & w1933;
assign w1697 = ~w1627 & w1696;
assign v637 = ~(w1695 | w1697);
assign w1698 = v637;
assign w1699 = w1620 & w1629;
assign w1700 = (~w1589 & w1581) | (~w1589 & w1934) | (w1581 & w1934);
assign w1701 = (~w1700 & w1598) | (~w1700 & w1935) | (w1598 & w1935);
assign w1702 = (w1701 & ~w1607) | (w1701 & w1936) | (~w1607 & w1936);
assign w1703 = (~w1702 & w1580) | (~w1702 & w1839) | (w1580 & w1839);
assign w1704 = (w1701 & w1607) | (w1701 & w1937) | (w1607 & w1937);
assign w1705 = (w1704 & ~w1575) | (w1704 & w1938) | (~w1575 & w1938);
assign v638 = ~(w1703 | w1705);
assign w1706 = v638;
assign w1707 = w1699 & ~w1706;
assign w1708 = ~w1699 & w1706;
assign v639 = ~(w1707 | w1708);
assign w1709 = v639;
assign w1710 = ~w1439 & w2050;
assign w1711 = w1620 & w1710;
assign w1712 = ~w1709 & w1711;
assign w1713 = w1709 & ~w1711;
assign v640 = ~(w1712 | w1713);
assign w1714 = v640;
assign w1715 = w1698 & ~w1714;
assign w1716 = ~w1698 & w1714;
assign v641 = ~(w1715 | w1716);
assign w1717 = v641;
assign w1718 = w1693 & w1717;
assign v642 = ~(w1693 | w1717);
assign w1719 = v642;
assign v643 = ~(w1718 | w1719);
assign w1720 = v643;
assign w1721 = w1690 & w1720;
assign v644 = ~(w1690 | w1720);
assign w1722 = v644;
assign v645 = ~(w1721 | w1722);
assign w1723 = v645;
assign w1724 = w1668 & ~w1723;
assign w1725 = ~w1668 & w1723;
assign v646 = ~(w1724 | w1725);
assign w1726 = v646;
assign w1727 = w1543 & ~w1649;
assign w1728 = w932 & ~w1226;
assign w1729 = w1533 & w1728;
assign v647 = ~(w1552 | w1729);
assign w1730 = v647;
assign w1731 = ~w1727 & w1730;
assign w1732 = w1549 & w1649;
assign v648 = ~(w1659 | w1732);
assign w1733 = v648;
assign w1734 = ~w1731 & w1733;
assign w1735 = ~w1652 & w1653;
assign v649 = ~(w1734 | w1735);
assign w1736 = v649;
assign w1737 = w1726 & w1736;
assign v650 = ~(w1726 | w1736);
assign w1738 = v650;
assign v651 = ~(w1737 | w1738);
assign w1739 = v651;
assign w1740 = (w1672 & ~w1720) | (w1672 & w1800) | (~w1720 & w1800);
assign w1741 = (w1683 & ~w1686) | (w1683 & w2051) | (~w1686 & w2051);
assign w1742 = ~w1677 & w1717;
assign v652 = ~(w1741 | w1742);
assign w1743 = v652;
assign w1744 = (~w1677 & ~w1686) | (~w1677 & w1939) | (~w1686 & w1939);
assign v653 = ~(w1717 | w1744);
assign w1745 = v653;
assign w1746 = (~w1711 & w1627) | (~w1711 & w1940) | (w1627 & w1940);
assign w1747 = w1579 & ~w1617;
assign w1748 = (w1620 & w2052) | (w1620 & w2053) | (w2052 & w2053);
assign w1749 = (~w1748 & w1746) | (~w1748 & w1942) | (w1746 & w1942);
assign w1750 = (w1749 & w1714) | (w1749 & w2054) | (w1714 & w2054);
assign w1751 = ~w1743 & w1943;
assign w1752 = ~w1740 & w1751;
assign v654 = ~(w1552 | w1654);
assign w1753 = v654;
assign v655 = ~(w1732 | w1753);
assign w1754 = v655;
assign w1755 = ~w1649 & w1801;
assign w1756 = w1541 & ~w1649;
assign w1757 = w1723 & w1756;
assign w1758 = w1233 & w1802;
assign w1759 = ~w1652 & w1758;
assign w1760 = w1752 & ~w1754;
assign v656 = ~(w1755 | w1757);
assign w1761 = v656;
assign w1762 = w1760 & w1761;
assign v657 = ~(w1725 | w1759);
assign w1763 = v657;
assign w1764 = w1762 & w1763;
assign w1765 = w1668 & w1944;
assign v658 = ~(w1764 | w1765);
assign w1766 = v658;
assign w1767 = w63 & ~w64;
assign w1768 = w87 & ~w88;
assign v659 = ~(w65 | w72);
assign w1769 = v659;
assign w1770 = (~w73 & ~w65) | (~w73 & w1945) | (~w65 & w1945);
assign w1771 = w137 & ~w124;
assign v660 = ~(w135 | w123);
assign w1772 = v660;
assign v661 = ~(w199 | w186);
assign w1773 = v661;
assign v662 = ~(w711 | w303);
assign w1774 = v662;
assign v663 = ~(w221 | w304);
assign w1775 = v663;
assign v664 = ~(w236 | w239);
assign w1776 = v664;
assign w1777 = w322 & ~w321;
assign w1778 = w379 & ~w378;
assign v665 = ~(w569 | w567);
assign w1779 = v665;
assign w1780 = (~w587 & w578) | (~w587 & w1946) | (w578 & w1946);
assign w1781 = w803 & w805;
assign w1782 = w781 & ~w1004;
assign v666 = ~(w1012 | w986);
assign w1783 = v666;
assign v667 = ~(w631 | w1026);
assign w1784 = v667;
assign w1785 = (~w1034 & ~w631) | (~w1034 & w1947) | (~w631 & w1947);
assign w1786 = w1065 & ~w1059;
assign v668 = ~(w735 | w1088);
assign w1787 = v668;
assign w1788 = w940 & ~w935;
assign w1789 = (w1058 & w735) | (w1058 & w1803) | (w735 & w1803);
assign w1790 = ~w1351 & w1093;
assign w1791 = w1351 & ~w1093;
assign v669 = ~(w1354 | w1372);
assign w1792 = v669;
assign w1793 = w1167 & ~w1417;
assign w1794 = w1445 & w1252;
assign w1795 = ~w1434 & w1572;
assign w1796 = (~w1179 & ~w1444) | (~w1179 & w1948) | (~w1444 & w1948);
assign w1797 = (~w1189 & ~w1437) | (~w1189 & w1949) | (~w1437 & w1949);
assign w1798 = w1642 & ~w1561;
assign w1799 = ~w1483 & w1490;
assign w1800 = ~w1670 & w2055;
assign w1801 = ~w1542 & w1950;
assign w1802 = w1533 & ~w937;
assign w1803 = ~w622 & w1058;
assign w1804 = w258 & ~w259;
assign w1805 = w273 & ~w274;
assign w1806 = w165 & ~w166;
assign w1807 = w133 & ~w132;
assign w1808 = w195 & ~w196;
assign v670 = ~(w698 | w186);
assign w1809 = v670;
assign w1810 = ~w199 & w1809;
assign w1811 = w294 & ~w295;
assign v671 = ~(w443 | w437);
assign w1812 = v671;
assign w1813 = w432 & ~w433;
assign w1814 = w495 & ~w496;
assign v672 = ~(w485 | w483);
assign w1815 = v672;
assign w1816 = w870 & ~w871;
assign v673 = ~(w701 | w700);
assign w1817 = v673;
assign v674 = ~(w684 | w689);
assign w1818 = v674;
assign w1819 = w1112 & ~w1111;
assign w1820 = (~w1141 & w772) | (~w1141 & w1951) | (w772 & w1951);
assign w1821 = w455 & w2056;
assign w1822 = w862 & w1199;
assign w1823 = (~w558 & w921) | (~w558 & w1952) | (w921 & w1952);
assign w1824 = w1077 & ~w1302;
assign w1825 = ~w959 & w1454;
assign w1826 = w955 & w1953;
assign w1827 = w955 & w2057;
assign w1828 = w911 & ~w1497;
assign w1829 = (w907 & w2058) | (w907 & w2059) | (w2058 & w2059);
assign w1830 = (~w1528 & ~w1218) | (~w1528 & w1954) | (~w1218 & w1954);
assign w1831 = ~w1530 & w1523;
assign v675 = ~(w1229 | w1524);
assign w1832 = v675;
assign w1833 = w1218 & ~w1546;
assign w1834 = (~w1518 & ~w1496) | (~w1518 & w1955) | (~w1496 & w1955);
assign v676 = ~(w1447 | w1469);
assign w1835 = v676;
assign w1836 = w1447 & w1469;
assign w1837 = w1457 & w1513;
assign w1838 = w1413 & ~w1378;
assign v677 = ~(w1617 | w1702);
assign w1839 = v677;
assign v678 = ~(w506 | w504);
assign w1840 = v678;
assign w1841 = (w551 & w545) | (w551 & w552) | (w545 & w552);
assign v679 = ~(w29 | w27);
assign w1842 = v679;
assign w1843 = ~w425 & w432;
assign v680 = ~(w332 | w331);
assign w1844 = v680;
assign w1845 = w213 & ~w214;
assign w1846 = ~w154 & w170;
assign w1847 = w154 & ~w170;
assign v681 = ~(w677 | w676);
assign w1848 = v681;
assign v682 = ~(w236 | w235);
assign w1849 = v682;
assign v683 = ~(w392 | w391);
assign w1850 = v683;
assign w1851 = w400 & ~w399;
assign w1852 = ~w383 & w441;
assign w1853 = w843 & ~w842;
assign v684 = ~(w461 | w464);
assign w1854 = v684;
assign w1855 = w45 & ~w46;
assign w1856 = (w452 & w1956) | (w452 & w1957) | (w1956 & w1957);
assign w1857 = (~w452 & w1958) | (~w452 & w1959) | (w1958 & w1959);
assign v685 = ~(w38 | w37);
assign w1858 = v685;
assign w1859 = (~w473 & w1960) | (~w473 & w1961) | (w1960 & w1961);
assign w1860 = (~w473 & w1962) | (~w473 & w1963) | (w1962 & w1963);
assign w1861 = (w473 & w1964) | (w473 & w1965) | (w1964 & w1965);
assign w1862 = (w473 & w1966) | (w473 & w1967) | (w1966 & w1967);
assign v686 = ~(w20 | w18);
assign w1863 = v686;
assign v687 = ~(w600 | w908);
assign w1864 = v687;
assign w1865 = (~w903 & w1968) | (~w903 & w1969) | (w1968 & w1969);
assign w1866 = ~w600 & w908;
assign v688 = ~(w542 | w540);
assign w1867 = v688;
assign v689 = ~(w11 | w9);
assign w1868 = v689;
assign w1869 = (w530 & w1970) | (w530 & w1971) | (w1970 & w1971);
assign w1870 = (w530 & w1972) | (w530 & w1973) | (w1972 & w1973);
assign w1871 = (~w530 & w1974) | (~w530 & w1975) | (w1974 & w1975);
assign w1872 = (~w530 & w1976) | (~w530 & w1977) | (w1976 & w1977);
assign w1873 = ~w911 & w918;
assign w1874 = w911 & ~w918;
assign v690 = ~(w2 | w568);
assign w1875 = v690;
assign w1876 = (~w567 & w557) | (~w567 & w1978) | (w557 & w1978);
assign w1877 = (w1779 & w557) | (w1779 & w1979) | (w557 & w1979);
assign w1878 = (w581 & w572) | (w581 & w1980) | (w572 & w1980);
assign w1879 = w933 & ~w937;
assign v691 = ~(w940 | w935);
assign w1880 = v691;
assign w1881 = (~w907 & w1981) | (~w907 & w1982) | (w1981 & w1982);
assign w1882 = (w907 & w1983) | (w907 & w1984) | (w1983 & w1984);
assign w1883 = w601 & ~w950;
assign w1884 = (~w904 & ~w900) | (~w904 & w1985) | (~w900 & w1985);
assign v692 = ~(w791 | w790);
assign w1885 = v692;
assign v693 = ~(w844 | w842);
assign w1886 = v693;
assign w1887 = w317 & ~w331;
assign w1888 = ~w332 & w1887;
assign v694 = ~(w672 | w670);
assign w1889 = v694;
assign w1890 = ~w287 & w294;
assign w1891 = w771 & ~w770;
assign w1892 = w38 & ~w479;
assign w1893 = (~w903 & w1986) | (~w903 & w1987) | (w1986 & w1987);
assign v695 = ~(w1232 | w1227);
assign w1894 = v695;
assign w1895 = w425 & ~w428;
assign v696 = ~(w1242 | w1246);
assign w1896 = v696;
assign w1897 = (w1176 & w1988) | (w1176 & w1989) | (w1988 & w1989);
assign w1898 = (~w374 & ~w788) | (~w374 & w1990) | (~w788 & w1990);
assign w1899 = w788 & w1991;
assign v697 = ~(w803 | w391);
assign w1900 = v697;
assign w1901 = w985 & ~w1002;
assign w1902 = ~w1294 & w822;
assign w1903 = w218 & ~w209;
assign w1904 = ~w769 & w755;
assign w1905 = w665 & ~w1330;
assign w1906 = ~w1100 & w1331;
assign w1907 = w769 & w762;
assign w1908 = w1341 & ~w1339;
assign w1909 = w65 & ~w68;
assign w1910 = w631 & w1409;
assign w1911 = w1036 & ~w1411;
assign v698 = ~(w488 | w500);
assign w1912 = v698;
assign v699 = ~(w888 | w1466);
assign w1913 = v699;
assign w1914 = (~w1497 & ~w903) | (~w1497 & w1992) | (~w903 & w1992);
assign w1915 = w1231 & w1533;
assign v700 = ~(w1231 | w1533);
assign w1916 = v700;
assign w1917 = w1218 & w1993;
assign w1918 = w1537 & ~w1548;
assign v701 = ~(w1335 | w1339);
assign w1919 = v701;
assign w1920 = ~w1121 & w1994;
assign w1921 = (w1586 & ~w1137) | (w1586 & w1995) | (~w1137 & w1995);
assign v702 = ~(w1585 | w1311);
assign w1922 = v702;
assign w1923 = w1015 & w1423;
assign w1924 = w1250 & w1996;
assign w1925 = ~w1447 & w1635;
assign w1926 = w1232 & w1533;
assign w1927 = w527 & w1997;
assign w1928 = (~w1663 & ~w1496) | (~w1663 & w1998) | (~w1496 & w1998);
assign w1929 = w1218 & w1545;
assign w1930 = w1452 & ~w1674;
assign v703 = ~(w1447 | w1483);
assign w1931 = v703;
assign w1932 = ~w1634 & w1681;
assign w1933 = (w1468 & ~w1437) | (w1468 & w1999) | (~w1437 & w1999);
assign v704 = ~(w1595 | w1589);
assign w1934 = v704;
assign v705 = ~(w1604 | w1700);
assign w1935 = v705;
assign w1936 = ~w1614 & w1701;
assign w1937 = w1614 & w1701;
assign w1938 = ~w1579 & w1704;
assign v706 = ~(w1211 | w1677);
assign w1939 = v706;
assign w1940 = (~w1694 & ~w1620) | (~w1694 & w2000) | (~w1620 & w2000);
assign w1941 = (~w1629 & w1747) | (~w1629 & w2001) | (w1747 & w2001);
assign w1942 = w1708 & ~w1748;
assign w1943 = w1750 & ~w1745;
assign w1944 = ~w1723 & w1752;
assign w1945 = w72 & ~w73;
assign v707 = ~(w581 | w587);
assign w1946 = v707;
assign w1947 = w1026 & ~w1034;
assign w1948 = w1443 & ~w1179;
assign w1949 = (~w1189 & ~w1250) | (~w1189 & w2002) | (~w1250 & w2002);
assign v708 = ~(w1537 | w1527);
assign w1950 = v708;
assign w1951 = (w1140 & w746) | (w1140 & w2003) | (w746 & w2003);
assign w1952 = w599 & ~w558;
assign w1953 = w885 & ~w503;
assign w1954 = w949 & ~w1528;
assign v709 = ~(w1498 | w1518);
assign w1955 = v709;
assign v710 = ~(w50 | w46);
assign w1956 = v710;
assign w1957 = ~w50 & w1855;
assign w1958 = w50 & w46;
assign w1959 = w50 & ~w1855;
assign w1960 = ~w483 & w37;
assign w1961 = (~w483 & w38) | (~w483 & w1960) | (w38 & w1960);
assign w1962 = ~w485 & w1960;
assign w1963 = w1815 & ~w1858;
assign w1964 = w483 & ~w37;
assign w1965 = ~w38 & w1964;
assign w1966 = (~w37 & w485) | (~w37 & w1964) | (w485 & w1964);
assign w1967 = ~w1815 & w1858;
assign w1968 = w600 & ~w908;
assign w1969 = w600 & w1864;
assign w1970 = w540 & ~w9;
assign w1971 = ~w11 & w1970;
assign w1972 = (~w9 & w542) | (~w9 & w1970) | (w542 & w1970);
assign w1973 = ~w1867 & w1868;
assign w1974 = ~w540 & w9;
assign w1975 = (~w540 & w11) | (~w540 & w1974) | (w11 & w1974);
assign w1976 = ~w542 & w1974;
assign w1977 = w1867 & ~w1868;
assign w1978 = w2 & ~w567;
assign w1979 = ~w569 & w1978;
assign w1980 = w575 & w581;
assign w1981 = (w903 & w2004) | (w903 & w2005) | (w2004 & w2005);
assign w1982 = (w903 & w2006) | (w903 & w2007) | (w2006 & w2007);
assign w1983 = (~w903 & w2008) | (~w903 & w2009) | (w2008 & w2009);
assign w1984 = (~w903 & w2010) | (~w903 & w2011) | (w2010 & w2011);
assign v711 = ~(w1883 | w904);
assign w1985 = v711;
assign w1986 = w530 & w2012;
assign w1987 = w944 & ~w1866;
assign w1988 = ~w1251 & w1246;
assign v712 = ~(w1251 | w1896);
assign w1989 = v712;
assign w1990 = w404 & ~w374;
assign v713 = ~(w404 | w374);
assign w1991 = v713;
assign v714 = ~(w600 | w1497);
assign w1992 = v714;
assign w1993 = ~w949 & w1546;
assign w1994 = w1116 & ~w1317;
assign w1995 = w1341 & w1586;
assign w1996 = ~w1176 & w2013;
assign w1997 = ~w521 & w1660;
assign v715 = ~(w1498 | w1663);
assign w1998 = v715;
assign w1999 = w1252 & w1468;
assign v716 = ~(w1710 | w1694);
assign w2000 = v716;
assign w2001 = w1575 & ~w1629;
assign v717 = ~(w1187 | w1189);
assign w2002 = v717;
assign w2003 = ~w754 & w1140;
assign w2004 = w915 & ~w1968;
assign w2005 = w915 & ~w1969;
assign w2006 = (w530 & w2014) | (w530 & w2015) | (w2014 & w2015);
assign w2007 = w915 & ~w1864;
assign w2008 = ~w915 & w1968;
assign w2009 = ~w915 & w1969;
assign w2010 = (~w530 & w2016) | (~w530 & w2017) | (w2016 & w2017);
assign w2011 = ~w915 & w1864;
assign w2012 = (~w527 & w2018) | (~w527 & w2019) | (w2018 & w2019);
assign w2013 = ~w1242 & w981;
assign w2014 = (w527 & w2020) | (w527 & w2021) | (w2020 & w2021);
assign w2015 = (w527 & w2022) | (w527 & w2023) | (w2022 & w2023);
assign w2016 = (~w527 & w2024) | (~w527 & w2025) | (w2024 & w2025);
assign w2017 = (~w527 & w2026) | (~w527 & w2027) | (w2026 & w2027);
assign w2018 = ~w5 & w18;
assign w2019 = (~w5 & w20) | (~w5 & w2018) | (w20 & w2018);
assign v718 = ~(w9 | w18);
assign w2020 = v718;
assign w2021 = ~w20 & w2020;
assign w2022 = ~w11 & w2020;
assign w2023 = w1868 & w1863;
assign w2024 = w9 & w18;
assign w2025 = (w9 & w20) | (w9 & w2024) | (w20 & w2024);
assign w2026 = (w18 & w11) | (w18 & w2024) | (w11 & w2024);
assign v719 = ~(w1868 | w1863);
assign w2027 = v719;
assign v720 = ~(w674 | w675);
assign w2028 = v720;
assign w2029 = (~w452 & w2060) | (~w452 & w2061) | (w2060 & w2061);
assign w2030 = w862 & ~w869;
assign w2031 = (w903 & w2062) | (w903 & w2063) | (w2062 & w2063);
assign v721 = ~(w925 | w1877);
assign w2032 = v721;
assign v722 = ~(w925 | w1876);
assign w2033 = v722;
assign w2034 = ~w680 & w678;
assign v723 = ~(w909 | w1865);
assign w2035 = v723;
assign v724 = ~(w909 | w910);
assign w2036 = v724;
assign w2037 = w1893 & w944;
assign w2038 = (w944 & w1893) | (w944 & ~w600) | (w1893 & ~w600);
assign v725 = ~(w1898 | w789);
assign w2039 = v725;
assign w2040 = ~w1318 & w1317;
assign v726 = ~(w1318 | w1920);
assign w2041 = v726;
assign w2042 = w1250 & w2064;
assign w2043 = w1250 & w2065;
assign w2044 = w1796 & ~w1632;
assign w2045 = ~w909 & w943;
assign w2046 = w1661 & w1662;
assign w2047 = ~w1665 & w1666;
assign w2048 = w1680 & ~w1682;
assign w2049 = w1796 & w1631;
assign w2050 = w1796 & ~w1190;
assign w2051 = w1506 & w1683;
assign v727 = ~(w1702 | w1941);
assign w2052 = v727;
assign w2053 = ~w1747 & w2066;
assign w2054 = ~w1697 & w1749;
assign v728 = ~(w1671 | w1684);
assign w2055 = v728;
assign w2056 = (w452 & w2067) | (w452 & w2068) | (w2067 & w2068);
assign v729 = ~(w488 | w503);
assign w2057 = v729;
assign v730 = ~(w952 | w1914);
assign w2058 = v730;
assign w2059 = ~w952 & w909;
assign w2060 = ~w458 & w46;
assign v731 = ~(w458 | w1855);
assign w2061 = v731;
assign w2062 = w600 & w908;
assign w2063 = w600 & w1866;
assign w2064 = ~w1176 & w2069;
assign w2065 = w981 & ~w1187;
assign v732 = ~(w1575 | w1702);
assign w2066 = v732;
assign v733 = ~(w458 | w46);
assign w2067 = v733;
assign w2068 = ~w458 & w1855;
assign w2069 = w2013 & ~w1187;
assign v734 = ~(w1548 | w1667);
assign w2070 = v734;
assign one = 1;
assign po0 = w596;// level 54
assign po1 = ~w942;// level 55
assign po2 = w1237;// level 56
assign po3 = w1536;// level 57
assign po4 = ~w1658;// level 59
assign po5 = ~w1739;// level 61
assign po6 = w1766;// level 61
endmodule
